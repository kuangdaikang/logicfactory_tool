// Benchmark "mem_ctrl" written by ABC on Fri Sep 15 11:26:50 2023

module mem_ctrl ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3291_, new_n3292_, new_n3293_, new_n3294_,
    new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_,
    new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_,
    new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_,
    new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_,
    new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_,
    new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_,
    new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_,
    new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_,
    new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_,
    new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_,
    new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_,
    new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_,
    new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_,
    new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_,
    new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_,
    new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_,
    new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_,
    new_n3475_, new_n3476_, new_n3477_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_,
    new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_,
    new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_,
    new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_,
    new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_,
    new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_,
    new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_,
    new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_,
    new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_,
    new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_,
    new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_,
    new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_,
    new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_,
    new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_,
    new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_,
    new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_,
    new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_,
    new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_,
    new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_,
    new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_,
    new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_,
    new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_,
    new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_,
    new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_,
    new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_,
    new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_,
    new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_,
    new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_,
    new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_,
    new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_,
    new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_,
    new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_,
    new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_,
    new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_,
    new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_,
    new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_,
    new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_,
    new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_,
    new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_,
    new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_,
    new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_,
    new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_,
    new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_,
    new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_,
    new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_,
    new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_,
    new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_,
    new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_,
    new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_,
    new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_,
    new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_,
    new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_,
    new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_,
    new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_,
    new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_,
    new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_,
    new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_,
    new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_,
    new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_,
    new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_,
    new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_,
    new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_,
    new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_,
    new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_,
    new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_,
    new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_,
    new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_,
    new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_,
    new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_,
    new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_,
    new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_,
    new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_,
    new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_,
    new_n4079_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_,
    new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_,
    new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_,
    new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_,
    new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_,
    new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_,
    new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_,
    new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_,
    new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_,
    new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_,
    new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_,
    new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_,
    new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_,
    new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_,
    new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_,
    new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_,
    new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_,
    new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_,
    new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_,
    new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_,
    new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_,
    new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_,
    new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_,
    new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_,
    new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_,
    new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_,
    new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_,
    new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_,
    new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_,
    new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_,
    new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_,
    new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_,
    new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_,
    new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_,
    new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_,
    new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_,
    new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_,
    new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_,
    new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_,
    new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_,
    new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_,
    new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_,
    new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_,
    new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_,
    new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_,
    new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_,
    new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_,
    new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_,
    new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_,
    new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_,
    new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_,
    new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_,
    new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_,
    new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_,
    new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_,
    new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_,
    new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_,
    new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_,
    new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_,
    new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_,
    new_n4882_, new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_,
    new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_,
    new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_,
    new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_,
    new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_,
    new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_,
    new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_,
    new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_,
    new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_,
    new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_,
    new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_,
    new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_,
    new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_,
    new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_,
    new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_,
    new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_,
    new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_,
    new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_,
    new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_,
    new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_,
    new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5327_, new_n5328_, new_n5329_, new_n5330_,
    new_n5331_, new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_,
    new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_,
    new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_,
    new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_,
    new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_,
    new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_,
    new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_,
    new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_,
    new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_,
    new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_,
    new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_,
    new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_,
    new_n5410_, new_n5411_, new_n5413_, new_n5414_, new_n5415_, new_n5416_,
    new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_,
    new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_,
    new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_,
    new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_,
    new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_,
    new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_,
    new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_,
    new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_,
    new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_,
    new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_,
    new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_,
    new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_,
    new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_,
    new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_,
    new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_,
    new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_,
    new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_,
    new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_,
    new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_,
    new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_,
    new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_,
    new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_,
    new_n5775_, new_n5776_, new_n5777_, new_n5779_, new_n5780_, new_n5781_,
    new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_,
    new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_,
    new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_,
    new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5805_,
    new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_,
    new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_,
    new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_,
    new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_,
    new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_,
    new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_,
    new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_,
    new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_,
    new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_,
    new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_,
    new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5871_, new_n5872_,
    new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_,
    new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_,
    new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_,
    new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_,
    new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_,
    new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_,
    new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_,
    new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_,
    new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_,
    new_n5927_, new_n5928_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_,
    new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_,
    new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_,
    new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_,
    new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_,
    new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_,
    new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_,
    new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_,
    new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_,
    new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_,
    new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_,
    new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_,
    new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_,
    new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_,
    new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_,
    new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_,
    new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6109_, new_n6110_,
    new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_,
    new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_,
    new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_,
    new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_,
    new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_,
    new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_,
    new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_,
    new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_,
    new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_,
    new_n6165_, new_n6166_, new_n6169_, new_n6170_, new_n6171_, new_n6172_,
    new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_,
    new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_,
    new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_,
    new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_,
    new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_,
    new_n6203_, new_n6205_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6245_, new_n6247_, new_n6249_, new_n6251_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_,
    new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_,
    new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_,
    new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_,
    new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_,
    new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_,
    new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_,
    new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_,
    new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_,
    new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_,
    new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_,
    new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_,
    new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_,
    new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_,
    new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_,
    new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_,
    new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_,
    new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_,
    new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_,
    new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_,
    new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_,
    new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_,
    new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_,
    new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_,
    new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_,
    new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_,
    new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_,
    new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_,
    new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_,
    new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_,
    new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_,
    new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_,
    new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_,
    new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_,
    new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_,
    new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_,
    new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_,
    new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_,
    new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_,
    new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_,
    new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_,
    new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_,
    new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_,
    new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_,
    new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_,
    new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_,
    new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_,
    new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_,
    new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_,
    new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_,
    new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_,
    new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_,
    new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_,
    new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_,
    new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_,
    new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_,
    new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_,
    new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_,
    new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_,
    new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_,
    new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_,
    new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_,
    new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_,
    new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_,
    new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_,
    new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_,
    new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_,
    new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_,
    new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_,
    new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_,
    new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_,
    new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_,
    new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_,
    new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_,
    new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_,
    new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_,
    new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_,
    new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_,
    new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_,
    new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_,
    new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_,
    new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_,
    new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_,
    new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_,
    new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_,
    new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_,
    new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_,
    new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_,
    new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_,
    new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_,
    new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_,
    new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_,
    new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_,
    new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_,
    new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_,
    new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_,
    new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_,
    new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_,
    new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_,
    new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_,
    new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_,
    new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_,
    new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_,
    new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_,
    new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_,
    new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_,
    new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_,
    new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_,
    new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_,
    new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_,
    new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_,
    new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_,
    new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_,
    new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_,
    new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_,
    new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_,
    new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_,
    new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_,
    new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_,
    new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_,
    new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_,
    new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_,
    new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_,
    new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_,
    new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_,
    new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_,
    new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_,
    new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_,
    new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_,
    new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_,
    new_n7261_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7290_, new_n7291_, new_n7292_,
    new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_,
    new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_,
    new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_,
    new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_,
    new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_,
    new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_,
    new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_,
    new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_,
    new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_,
    new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_,
    new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_,
    new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_,
    new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_,
    new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_,
    new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_,
    new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_,
    new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_,
    new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_,
    new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_,
    new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_,
    new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_,
    new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_,
    new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_,
    new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_,
    new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_,
    new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_,
    new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_,
    new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_,
    new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_,
    new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_,
    new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_,
    new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_,
    new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_,
    new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_,
    new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_,
    new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_,
    new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_,
    new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_,
    new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_,
    new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_,
    new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_,
    new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_,
    new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_,
    new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_,
    new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_,
    new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_,
    new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_,
    new_n7912_, new_n7913_, new_n7915_, new_n7916_, new_n7917_, new_n7918_,
    new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_,
    new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_,
    new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_,
    new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_,
    new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_,
    new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_,
    new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_,
    new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_,
    new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_,
    new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_,
    new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_,
    new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_,
    new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_,
    new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_,
    new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_,
    new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_,
    new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_,
    new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_,
    new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_,
    new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_,
    new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_,
    new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_,
    new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_,
    new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_,
    new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_,
    new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_,
    new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_,
    new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_,
    new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_,
    new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_,
    new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_,
    new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8241_, new_n8242_, new_n8243_, new_n8244_,
    new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_,
    new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_,
    new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_,
    new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_,
    new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_,
    new_n8276_, new_n8277_, new_n8278_, new_n8280_, new_n8281_, new_n8282_,
    new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_,
    new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_,
    new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_,
    new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_,
    new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_,
    new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_,
    new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_,
    new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_, new_n8330_,
    new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_,
    new_n8337_, new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_,
    new_n8344_, new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_,
    new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_,
    new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_,
    new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_,
    new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_,
    new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_,
    new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_,
    new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_,
    new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_,
    new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_,
    new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_,
    new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_,
    new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_,
    new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_,
    new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_,
    new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_,
    new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_,
    new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_,
    new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_,
    new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_,
    new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_,
    new_n8501_, new_n8502_, new_n8503_, new_n8505_, new_n8506_, new_n8507_,
    new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_,
    new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_,
    new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_,
    new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_,
    new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_,
    new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_,
    new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_,
    new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_,
    new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_,
    new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_,
    new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_,
    new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_,
    new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_,
    new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_,
    new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_,
    new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_,
    new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_,
    new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_,
    new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_,
    new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_,
    new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_,
    new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_,
    new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_,
    new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_,
    new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_,
    new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_,
    new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_,
    new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_,
    new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_,
    new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_,
    new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_,
    new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_,
    new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_,
    new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_,
    new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_,
    new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_,
    new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_,
    new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_,
    new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_,
    new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8896_, new_n8897_, new_n8898_, new_n8900_, new_n8901_,
    new_n8902_, new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_,
    new_n8908_, new_n8909_, new_n8910_, new_n8911_, new_n8913_, new_n8914_,
    new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_,
    new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_,
    new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_,
    new_n8933_, new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_,
    new_n8939_, new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_,
    new_n8946_, new_n8947_, new_n8948_, new_n8950_, new_n8951_, new_n8952_,
    new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_,
    new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_,
    new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_,
    new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_,
    new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_,
    new_n9004_, new_n9005_, new_n9006_, new_n9007_, new_n9008_, new_n9009_,
    new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_,
    new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_,
    new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_,
    new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_,
    new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_, new_n9039_,
    new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_, new_n9045_,
    new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_, new_n9051_,
    new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_,
    new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_, new_n9063_,
    new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_, new_n9069_,
    new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_, new_n9075_,
    new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_,
    new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_,
    new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_,
    new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_,
    new_n9101_, new_n9102_, new_n9103_, new_n9105_, new_n9106_, new_n9107_,
    new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_,
    new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9120_,
    new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_,
    new_n9127_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9134_,
    new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_,
    new_n9142_, new_n9143_, new_n9145_, new_n9146_, new_n9148_, new_n9149_,
    new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9155_, new_n9156_,
    new_n9158_, new_n9159_, new_n9161_, new_n9162_, new_n9164_, new_n9165_,
    new_n9166_, new_n9167_, new_n9169_, new_n9171_, new_n9172_, new_n9173_,
    new_n9174_, new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_,
    new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_,
    new_n9187_, new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_,
    new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_,
    new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_,
    new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_,
    new_n9214_, new_n9215_, new_n9217_, new_n9218_, new_n9219_, new_n9220_,
    new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_,
    new_n9227_, new_n9228_, new_n9229_, new_n9231_, new_n9232_, new_n9233_,
    new_n9234_, new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9240_,
    new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_,
    new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_,
    new_n9254_, new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_,
    new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_,
    new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_,
    new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_,
    new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_,
    new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_,
    new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_,
    new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_,
    new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_,
    new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_,
    new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_,
    new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_,
    new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_,
    new_n9383_, new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_,
    new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_,
    new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_,
    new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_,
    new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_,
    new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_,
    new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_,
    new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_,
    new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_,
    new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_,
    new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_,
    new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_,
    new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_,
    new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_,
    new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_,
    new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_,
    new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_,
    new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_,
    new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_,
    new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_,
    new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_,
    new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_,
    new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_,
    new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_,
    new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_,
    new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_,
    new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_,
    new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_,
    new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_,
    new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_,
    new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_,
    new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_,
    new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_,
    new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_,
    new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_,
    new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_,
    new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_,
    new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_,
    new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_,
    new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_,
    new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_,
    new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_,
    new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_,
    new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_,
    new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_,
    new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_,
    new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_,
    new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_,
    new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_,
    new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_,
    new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_,
    new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_,
    new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_,
    new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_,
    new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_,
    new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_,
    new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_,
    new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_,
    new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_,
    new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9745_,
    new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_,
    new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_,
    new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_,
    new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_,
    new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_,
    new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_,
    new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_,
    new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_,
    new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_, new_n9859_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_,
    new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_,
    new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_,
    new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10005_, new_n10006_, new_n10007_,
    new_n10008_, new_n10009_, new_n10010_, new_n10011_, new_n10012_,
    new_n10013_, new_n10014_, new_n10015_, new_n10016_, new_n10017_,
    new_n10018_, new_n10019_, new_n10020_, new_n10021_, new_n10022_,
    new_n10023_, new_n10024_, new_n10025_, new_n10026_, new_n10027_,
    new_n10028_, new_n10029_, new_n10030_, new_n10031_, new_n10032_,
    new_n10033_, new_n10034_, new_n10035_, new_n10036_, new_n10037_,
    new_n10038_, new_n10039_, new_n10040_, new_n10041_, new_n10042_,
    new_n10043_, new_n10044_, new_n10045_, new_n10046_, new_n10047_,
    new_n10048_, new_n10049_, new_n10050_, new_n10051_, new_n10052_,
    new_n10053_, new_n10054_, new_n10055_, new_n10056_, new_n10057_,
    new_n10058_, new_n10059_, new_n10060_, new_n10061_, new_n10062_,
    new_n10063_, new_n10064_, new_n10065_, new_n10066_, new_n10067_,
    new_n10068_, new_n10069_, new_n10070_, new_n10071_, new_n10072_,
    new_n10073_, new_n10074_, new_n10075_, new_n10076_, new_n10077_,
    new_n10078_, new_n10079_, new_n10080_, new_n10081_, new_n10082_,
    new_n10083_, new_n10084_, new_n10085_, new_n10086_, new_n10087_,
    new_n10088_, new_n10089_, new_n10090_, new_n10091_, new_n10092_,
    new_n10093_, new_n10094_, new_n10095_, new_n10096_, new_n10097_,
    new_n10098_, new_n10099_, new_n10100_, new_n10101_, new_n10102_,
    new_n10103_, new_n10104_, new_n10105_, new_n10106_, new_n10107_,
    new_n10108_, new_n10109_, new_n10110_, new_n10111_, new_n10112_,
    new_n10113_, new_n10114_, new_n10115_, new_n10116_, new_n10117_,
    new_n10118_, new_n10119_, new_n10120_, new_n10121_, new_n10122_,
    new_n10123_, new_n10124_, new_n10125_, new_n10126_, new_n10127_,
    new_n10128_, new_n10129_, new_n10130_, new_n10131_, new_n10132_,
    new_n10133_, new_n10134_, new_n10135_, new_n10136_, new_n10137_,
    new_n10138_, new_n10139_, new_n10140_, new_n10141_, new_n10142_,
    new_n10143_, new_n10144_, new_n10145_, new_n10146_, new_n10147_,
    new_n10148_, new_n10149_, new_n10150_, new_n10151_, new_n10152_,
    new_n10153_, new_n10154_, new_n10155_, new_n10156_, new_n10157_,
    new_n10158_, new_n10159_, new_n10160_, new_n10161_, new_n10162_,
    new_n10163_, new_n10164_, new_n10165_, new_n10166_, new_n10167_,
    new_n10168_, new_n10169_, new_n10170_, new_n10171_, new_n10172_,
    new_n10173_, new_n10174_, new_n10175_, new_n10176_, new_n10177_,
    new_n10178_, new_n10179_, new_n10180_, new_n10181_, new_n10182_,
    new_n10183_, new_n10184_, new_n10185_, new_n10186_, new_n10187_,
    new_n10188_, new_n10189_, new_n10190_, new_n10191_, new_n10192_,
    new_n10193_, new_n10194_, new_n10195_, new_n10196_, new_n10197_,
    new_n10198_, new_n10199_, new_n10200_, new_n10201_, new_n10202_,
    new_n10203_, new_n10204_, new_n10205_, new_n10206_, new_n10207_,
    new_n10208_, new_n10209_, new_n10210_, new_n10211_, new_n10212_,
    new_n10213_, new_n10214_, new_n10215_, new_n10216_, new_n10217_,
    new_n10218_, new_n10219_, new_n10220_, new_n10221_, new_n10222_,
    new_n10223_, new_n10224_, new_n10225_, new_n10226_, new_n10227_,
    new_n10228_, new_n10229_, new_n10230_, new_n10231_, new_n10232_,
    new_n10233_, new_n10234_, new_n10235_, new_n10236_, new_n10237_,
    new_n10238_, new_n10239_, new_n10240_, new_n10241_, new_n10242_,
    new_n10243_, new_n10244_, new_n10245_, new_n10246_, new_n10247_,
    new_n10248_, new_n10249_, new_n10250_, new_n10251_, new_n10252_,
    new_n10253_, new_n10254_, new_n10255_, new_n10256_, new_n10257_,
    new_n10258_, new_n10259_, new_n10260_, new_n10261_, new_n10262_,
    new_n10263_, new_n10264_, new_n10265_, new_n10266_, new_n10267_,
    new_n10268_, new_n10270_, new_n10271_, new_n10272_, new_n10273_,
    new_n10275_, new_n10276_, new_n10277_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10288_, new_n10289_, new_n10290_, new_n10292_,
    new_n10293_, new_n10294_, new_n10296_, new_n10297_, new_n10299_,
    new_n10300_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10314_, new_n10315_, new_n10316_,
    new_n10317_, new_n10319_, new_n10320_, new_n10322_, new_n10323_,
    new_n10324_, new_n10325_, new_n10326_, new_n10327_, new_n10328_,
    new_n10329_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10344_, new_n10345_, new_n10346_,
    new_n10347_, new_n10348_, new_n10349_, new_n10350_, new_n10351_,
    new_n10352_, new_n10353_, new_n10355_, new_n10356_, new_n10357_,
    new_n10358_, new_n10359_, new_n10360_, new_n10361_, new_n10362_,
    new_n10363_, new_n10364_, new_n10365_, new_n10367_, new_n10368_,
    new_n10369_, new_n10370_, new_n10371_, new_n10372_, new_n10373_,
    new_n10374_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10382_, new_n10384_, new_n10385_, new_n10386_,
    new_n10387_, new_n10388_, new_n10389_, new_n10390_, new_n10391_,
    new_n10392_, new_n10393_, new_n10394_, new_n10395_, new_n10396_,
    new_n10397_, new_n10398_, new_n10399_, new_n10400_, new_n10401_,
    new_n10402_, new_n10403_, new_n10404_, new_n10405_, new_n10406_,
    new_n10407_, new_n10408_, new_n10409_, new_n10410_, new_n10411_,
    new_n10412_, new_n10413_, new_n10414_, new_n10415_, new_n10416_,
    new_n10417_, new_n10418_, new_n10419_, new_n10420_, new_n10421_,
    new_n10422_, new_n10423_, new_n10424_, new_n10425_, new_n10426_,
    new_n10427_, new_n10428_, new_n10430_, new_n10431_, new_n10432_,
    new_n10433_, new_n10434_, new_n10435_, new_n10436_, new_n10437_,
    new_n10439_, new_n10440_, new_n10441_, new_n10442_, new_n10443_,
    new_n10444_, new_n10445_, new_n10446_, new_n10447_, new_n10448_,
    new_n10449_, new_n10450_, new_n10451_, new_n10452_, new_n10453_,
    new_n10454_, new_n10455_, new_n10456_, new_n10457_, new_n10458_,
    new_n10459_, new_n10460_, new_n10461_, new_n10462_, new_n10463_,
    new_n10464_, new_n10465_, new_n10466_, new_n10467_, new_n10468_,
    new_n10469_, new_n10470_, new_n10471_, new_n10472_, new_n10473_,
    new_n10474_, new_n10475_, new_n10476_, new_n10477_, new_n10478_,
    new_n10479_, new_n10480_, new_n10481_, new_n10482_, new_n10483_,
    new_n10484_, new_n10486_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10493_, new_n10494_, new_n10495_, new_n10496_,
    new_n10497_, new_n10498_, new_n10499_, new_n10500_, new_n10501_,
    new_n10502_, new_n10504_, new_n10505_, new_n10506_, new_n10507_,
    new_n10508_, new_n10510_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10524_, new_n10525_, new_n10526_,
    new_n10527_, new_n10528_, new_n10529_, new_n10531_, new_n10532_,
    new_n10534_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10592_, new_n10593_, new_n10594_, new_n10595_, new_n10596_,
    new_n10597_, new_n10598_, new_n10599_, new_n10600_, new_n10601_,
    new_n10602_, new_n10603_, new_n10604_, new_n10605_, new_n10606_,
    new_n10607_, new_n10608_, new_n10609_, new_n10610_, new_n10611_,
    new_n10612_, new_n10613_, new_n10614_, new_n10615_, new_n10616_,
    new_n10617_, new_n10618_, new_n10620_, new_n10621_, new_n10622_,
    new_n10623_, new_n10624_, new_n10625_, new_n10626_, new_n10627_,
    new_n10628_, new_n10629_, new_n10630_, new_n10631_, new_n10632_,
    new_n10633_, new_n10634_, new_n10635_, new_n10636_, new_n10637_,
    new_n10638_, new_n10639_, new_n10640_, new_n10641_, new_n10642_,
    new_n10643_, new_n10644_, new_n10645_, new_n10646_, new_n10647_,
    new_n10648_, new_n10649_, new_n10651_, new_n10652_, new_n10653_,
    new_n10654_, new_n10655_, new_n10656_, new_n10657_, new_n10658_,
    new_n10659_, new_n10660_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10846_, new_n10847_, new_n10848_, new_n10849_,
    new_n10850_, new_n10851_, new_n10852_, new_n10853_, new_n10854_,
    new_n10855_, new_n10856_, new_n10857_, new_n10858_, new_n10859_,
    new_n10860_, new_n10861_, new_n10862_, new_n10863_, new_n10864_,
    new_n10865_, new_n10866_, new_n10867_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10900_, new_n10901_,
    new_n10902_, new_n10903_, new_n10904_, new_n10905_, new_n10906_,
    new_n10907_, new_n10908_, new_n10909_, new_n10910_, new_n10911_,
    new_n10912_, new_n10913_, new_n10914_, new_n10915_, new_n10916_,
    new_n10917_, new_n10918_, new_n10919_, new_n10920_, new_n10921_,
    new_n10922_, new_n10923_, new_n10924_, new_n10925_, new_n10926_,
    new_n10927_, new_n10928_, new_n10929_, new_n10930_, new_n10931_,
    new_n10932_, new_n10933_, new_n10934_, new_n10935_, new_n10936_,
    new_n10937_, new_n10938_, new_n10939_, new_n10940_, new_n10941_,
    new_n10942_, new_n10943_, new_n10944_, new_n10945_, new_n10946_,
    new_n10947_, new_n10948_, new_n10949_, new_n10950_, new_n10951_,
    new_n10952_, new_n10953_, new_n10954_, new_n10955_, new_n10956_,
    new_n10957_, new_n10958_, new_n10959_, new_n10960_, new_n10961_,
    new_n10962_, new_n10963_, new_n10964_, new_n10965_, new_n10966_,
    new_n10967_, new_n10968_, new_n10969_, new_n10970_, new_n10971_,
    new_n10972_, new_n10973_, new_n10974_, new_n10975_, new_n10976_,
    new_n10977_, new_n10978_, new_n10979_, new_n10980_, new_n10981_,
    new_n10982_, new_n10983_, new_n10984_, new_n10985_, new_n10986_,
    new_n10987_, new_n10988_, new_n10989_, new_n10990_, new_n10991_,
    new_n10992_, new_n10993_, new_n10994_, new_n10995_, new_n10996_,
    new_n10997_, new_n10998_, new_n10999_, new_n11000_, new_n11001_,
    new_n11002_, new_n11003_, new_n11004_, new_n11005_, new_n11006_,
    new_n11007_, new_n11008_, new_n11009_, new_n11010_, new_n11011_,
    new_n11012_, new_n11013_, new_n11014_, new_n11015_, new_n11016_,
    new_n11017_, new_n11018_, new_n11019_, new_n11020_, new_n11021_,
    new_n11022_, new_n11023_, new_n11024_, new_n11025_, new_n11026_,
    new_n11027_, new_n11028_, new_n11029_, new_n11030_, new_n11031_,
    new_n11032_, new_n11033_, new_n11034_, new_n11035_, new_n11036_,
    new_n11037_, new_n11038_, new_n11039_, new_n11040_, new_n11041_,
    new_n11042_, new_n11043_, new_n11044_, new_n11045_, new_n11046_,
    new_n11047_, new_n11048_, new_n11049_, new_n11050_, new_n11051_,
    new_n11052_, new_n11053_, new_n11054_, new_n11055_, new_n11056_,
    new_n11057_, new_n11058_, new_n11059_, new_n11060_, new_n11061_,
    new_n11062_, new_n11063_, new_n11064_, new_n11065_, new_n11066_,
    new_n11067_, new_n11068_, new_n11069_, new_n11070_, new_n11071_,
    new_n11072_, new_n11073_, new_n11074_, new_n11075_, new_n11076_,
    new_n11077_, new_n11078_, new_n11079_, new_n11080_, new_n11081_,
    new_n11082_, new_n11083_, new_n11084_, new_n11085_, new_n11086_,
    new_n11087_, new_n11088_, new_n11089_, new_n11090_, new_n11091_,
    new_n11092_, new_n11093_, new_n11094_, new_n11095_, new_n11096_,
    new_n11097_, new_n11098_, new_n11099_, new_n11100_, new_n11101_,
    new_n11102_, new_n11103_, new_n11104_, new_n11105_, new_n11106_,
    new_n11107_, new_n11108_, new_n11109_, new_n11110_, new_n11111_,
    new_n11112_, new_n11113_, new_n11114_, new_n11115_, new_n11116_,
    new_n11117_, new_n11118_, new_n11119_, new_n11120_, new_n11121_,
    new_n11122_, new_n11123_, new_n11124_, new_n11125_, new_n11126_,
    new_n11127_, new_n11128_, new_n11129_, new_n11130_, new_n11131_,
    new_n11132_, new_n11133_, new_n11134_, new_n11135_, new_n11136_,
    new_n11137_, new_n11138_, new_n11139_, new_n11140_, new_n11141_,
    new_n11142_, new_n11143_, new_n11144_, new_n11145_, new_n11146_,
    new_n11147_, new_n11148_, new_n11149_, new_n11150_, new_n11151_,
    new_n11152_, new_n11153_, new_n11155_, new_n11156_, new_n11157_,
    new_n11158_, new_n11159_, new_n11160_, new_n11161_, new_n11162_,
    new_n11163_, new_n11164_, new_n11165_, new_n11166_, new_n11167_,
    new_n11168_, new_n11169_, new_n11170_, new_n11171_, new_n11172_,
    new_n11173_, new_n11174_, new_n11175_, new_n11176_, new_n11177_,
    new_n11178_, new_n11179_, new_n11180_, new_n11181_, new_n11182_,
    new_n11183_, new_n11184_, new_n11185_, new_n11186_, new_n11187_,
    new_n11188_, new_n11189_, new_n11190_, new_n11191_, new_n11192_,
    new_n11193_, new_n11194_, new_n11195_, new_n11196_, new_n11197_,
    new_n11198_, new_n11199_, new_n11200_, new_n11201_, new_n11202_,
    new_n11203_, new_n11204_, new_n11205_, new_n11206_, new_n11207_,
    new_n11208_, new_n11209_, new_n11210_, new_n11211_, new_n11212_,
    new_n11213_, new_n11214_, new_n11215_, new_n11216_, new_n11217_,
    new_n11218_, new_n11219_, new_n11220_, new_n11221_, new_n11222_,
    new_n11223_, new_n11224_, new_n11225_, new_n11226_, new_n11227_,
    new_n11228_, new_n11229_, new_n11230_, new_n11231_, new_n11232_,
    new_n11233_, new_n11234_, new_n11235_, new_n11236_, new_n11237_,
    new_n11238_, new_n11239_, new_n11240_, new_n11241_, new_n11242_,
    new_n11243_, new_n11244_, new_n11245_, new_n11246_, new_n11247_,
    new_n11248_, new_n11249_, new_n11250_, new_n11251_, new_n11252_,
    new_n11253_, new_n11254_, new_n11255_, new_n11256_, new_n11257_,
    new_n11258_, new_n11259_, new_n11260_, new_n11261_, new_n11262_,
    new_n11263_, new_n11264_, new_n11265_, new_n11266_, new_n11267_,
    new_n11268_, new_n11269_, new_n11270_, new_n11271_, new_n11272_,
    new_n11273_, new_n11274_, new_n11275_, new_n11276_, new_n11277_,
    new_n11278_, new_n11279_, new_n11280_, new_n11281_, new_n11282_,
    new_n11283_, new_n11284_, new_n11285_, new_n11286_, new_n11287_,
    new_n11288_, new_n11289_, new_n11290_, new_n11291_, new_n11292_,
    new_n11293_, new_n11294_, new_n11295_, new_n11296_, new_n11297_,
    new_n11298_, new_n11299_, new_n11300_, new_n11301_, new_n11302_,
    new_n11303_, new_n11304_, new_n11305_, new_n11306_, new_n11307_,
    new_n11308_, new_n11309_, new_n11310_, new_n11311_, new_n11312_,
    new_n11313_, new_n11314_, new_n11315_, new_n11316_, new_n11317_,
    new_n11318_, new_n11319_, new_n11320_, new_n11321_, new_n11322_,
    new_n11323_, new_n11324_, new_n11325_, new_n11326_, new_n11327_,
    new_n11328_, new_n11329_, new_n11330_, new_n11331_, new_n11332_,
    new_n11333_, new_n11334_, new_n11335_, new_n11336_, new_n11337_,
    new_n11338_, new_n11339_, new_n11340_, new_n11341_, new_n11342_,
    new_n11343_, new_n11344_, new_n11345_, new_n11346_, new_n11347_,
    new_n11348_, new_n11349_, new_n11350_, new_n11351_, new_n11352_,
    new_n11353_, new_n11354_, new_n11355_, new_n11356_, new_n11357_,
    new_n11358_, new_n11359_, new_n11360_, new_n11361_, new_n11362_,
    new_n11363_, new_n11364_, new_n11365_, new_n11366_, new_n11367_,
    new_n11368_, new_n11369_, new_n11370_, new_n11371_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11387_,
    new_n11388_, new_n11389_, new_n11390_, new_n11391_, new_n11392_,
    new_n11393_, new_n11394_, new_n11395_, new_n11396_, new_n11397_,
    new_n11398_, new_n11399_, new_n11400_, new_n11401_, new_n11402_,
    new_n11403_, new_n11404_, new_n11405_, new_n11406_, new_n11407_,
    new_n11408_, new_n11409_, new_n11410_, new_n11411_, new_n11412_,
    new_n11413_, new_n11414_, new_n11415_, new_n11416_, new_n11417_,
    new_n11418_, new_n11419_, new_n11420_, new_n11421_, new_n11422_,
    new_n11423_, new_n11424_, new_n11425_, new_n11426_, new_n11427_,
    new_n11428_, new_n11429_, new_n11430_, new_n11431_, new_n11432_,
    new_n11433_, new_n11434_, new_n11435_, new_n11436_, new_n11437_,
    new_n11438_, new_n11439_, new_n11440_, new_n11441_, new_n11442_,
    new_n11443_, new_n11444_, new_n11445_, new_n11446_, new_n11447_,
    new_n11448_, new_n11449_, new_n11450_, new_n11451_, new_n11452_,
    new_n11453_, new_n11454_, new_n11455_, new_n11456_, new_n11457_,
    new_n11458_, new_n11459_, new_n11460_, new_n11461_, new_n11462_,
    new_n11463_, new_n11464_, new_n11465_, new_n11466_, new_n11467_,
    new_n11468_, new_n11469_, new_n11470_, new_n11471_, new_n11472_,
    new_n11473_, new_n11474_, new_n11475_, new_n11476_, new_n11477_,
    new_n11478_, new_n11479_, new_n11480_, new_n11481_, new_n11482_,
    new_n11483_, new_n11484_, new_n11485_, new_n11486_, new_n11487_,
    new_n11488_, new_n11489_, new_n11490_, new_n11491_, new_n11492_,
    new_n11493_, new_n11494_, new_n11495_, new_n11496_, new_n11498_,
    new_n11499_, new_n11500_, new_n11501_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_,
    new_n11515_, new_n11516_, new_n11517_, new_n11518_, new_n11519_,
    new_n11520_, new_n11521_, new_n11522_, new_n11523_, new_n11524_,
    new_n11525_, new_n11526_, new_n11527_, new_n11528_, new_n11529_,
    new_n11530_, new_n11531_, new_n11532_, new_n11533_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11694_, new_n11695_,
    new_n11696_, new_n11697_, new_n11698_, new_n11699_, new_n11700_,
    new_n11701_, new_n11702_, new_n11703_, new_n11704_, new_n11705_,
    new_n11706_, new_n11707_, new_n11708_, new_n11709_, new_n11710_,
    new_n11711_, new_n11712_, new_n11713_, new_n11714_, new_n11715_,
    new_n11716_, new_n11717_, new_n11718_, new_n11719_, new_n11720_,
    new_n11721_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11730_,
    new_n11731_, new_n11732_, new_n11733_, new_n11734_, new_n11735_,
    new_n11736_, new_n11737_, new_n11738_, new_n11739_, new_n11740_,
    new_n11741_, new_n11742_, new_n11743_, new_n11744_, new_n11745_,
    new_n11746_, new_n11747_, new_n11748_, new_n11749_, new_n11750_,
    new_n11751_, new_n11752_, new_n11753_, new_n11754_, new_n11755_,
    new_n11756_, new_n11757_, new_n11758_, new_n11759_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11808_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11835_, new_n11836_,
    new_n11837_, new_n11838_, new_n11839_, new_n11840_, new_n11841_,
    new_n11842_, new_n11843_, new_n11844_, new_n11845_, new_n11846_,
    new_n11847_, new_n11848_, new_n11849_, new_n11850_, new_n11851_,
    new_n11852_, new_n11853_, new_n11854_, new_n11855_, new_n11856_,
    new_n11857_, new_n11858_, new_n11859_, new_n11860_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11866_,
    new_n11867_, new_n11868_, new_n11869_, new_n11870_, new_n11871_,
    new_n11872_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11880_, new_n11881_,
    new_n11882_, new_n11883_, new_n11884_, new_n11885_, new_n11886_,
    new_n11887_, new_n11888_, new_n11889_, new_n11890_, new_n11891_,
    new_n11892_, new_n11893_, new_n11894_, new_n11895_, new_n11896_,
    new_n11897_, new_n11898_, new_n11899_, new_n11900_, new_n11901_,
    new_n11902_, new_n11903_, new_n11904_, new_n11905_, new_n11906_,
    new_n11907_, new_n11908_, new_n11909_, new_n11910_, new_n11911_,
    new_n11912_, new_n11913_, new_n11914_, new_n11915_, new_n11916_,
    new_n11917_, new_n11918_, new_n11919_, new_n11920_, new_n11921_,
    new_n11922_, new_n11923_, new_n11924_, new_n11925_, new_n11926_,
    new_n11927_, new_n11928_, new_n11929_, new_n11930_, new_n11931_,
    new_n11932_, new_n11933_, new_n11934_, new_n11935_, new_n11936_,
    new_n11937_, new_n11938_, new_n11939_, new_n11940_, new_n11941_,
    new_n11942_, new_n11943_, new_n11944_, new_n11945_, new_n11946_,
    new_n11947_, new_n11948_, new_n11949_, new_n11950_, new_n11951_,
    new_n11952_, new_n11953_, new_n11954_, new_n11955_, new_n11956_,
    new_n11957_, new_n11958_, new_n11959_, new_n11960_, new_n11961_,
    new_n11962_, new_n11963_, new_n11964_, new_n11965_, new_n11966_,
    new_n11967_, new_n11968_, new_n11969_, new_n11970_, new_n11971_,
    new_n11972_, new_n11973_, new_n11974_, new_n11975_, new_n11976_,
    new_n11977_, new_n11978_, new_n11979_, new_n11980_, new_n11981_,
    new_n11982_, new_n11983_, new_n11984_, new_n11985_, new_n11986_,
    new_n11987_, new_n11988_, new_n11989_, new_n11990_, new_n11991_,
    new_n11992_, new_n11993_, new_n11994_, new_n11995_, new_n11996_,
    new_n11997_, new_n11998_, new_n11999_, new_n12000_, new_n12001_,
    new_n12002_, new_n12003_, new_n12004_, new_n12005_, new_n12006_,
    new_n12007_, new_n12008_, new_n12009_, new_n12010_, new_n12011_,
    new_n12012_, new_n12013_, new_n12014_, new_n12015_, new_n12016_,
    new_n12017_, new_n12018_, new_n12019_, new_n12020_, new_n12021_,
    new_n12022_, new_n12023_, new_n12024_, new_n12025_, new_n12026_,
    new_n12027_, new_n12028_, new_n12029_, new_n12030_, new_n12031_,
    new_n12032_, new_n12033_, new_n12034_, new_n12035_, new_n12036_,
    new_n12037_, new_n12038_, new_n12039_, new_n12041_, new_n12042_,
    new_n12043_, new_n12044_, new_n12045_, new_n12046_, new_n12047_,
    new_n12048_, new_n12049_, new_n12050_, new_n12051_, new_n12052_,
    new_n12053_, new_n12054_, new_n12055_, new_n12056_, new_n12057_,
    new_n12058_, new_n12059_, new_n12060_, new_n12061_, new_n12062_,
    new_n12063_, new_n12064_, new_n12065_, new_n12066_, new_n12067_,
    new_n12068_, new_n12069_, new_n12070_, new_n12071_, new_n12072_,
    new_n12073_, new_n12074_, new_n12075_, new_n12076_, new_n12077_,
    new_n12078_, new_n12079_, new_n12080_, new_n12081_, new_n12082_,
    new_n12083_, new_n12084_, new_n12085_, new_n12086_, new_n12087_,
    new_n12088_, new_n12089_, new_n12090_, new_n12091_, new_n12092_,
    new_n12093_, new_n12094_, new_n12095_, new_n12096_, new_n12097_,
    new_n12098_, new_n12099_, new_n12100_, new_n12102_, new_n12103_,
    new_n12104_, new_n12105_, new_n12106_, new_n12107_, new_n12108_,
    new_n12109_, new_n12110_, new_n12111_, new_n12112_, new_n12113_,
    new_n12114_, new_n12116_, new_n12117_, new_n12118_, new_n12119_,
    new_n12120_, new_n12121_, new_n12122_, new_n12123_, new_n12124_,
    new_n12125_, new_n12126_, new_n12127_, new_n12128_, new_n12129_,
    new_n12130_, new_n12131_, new_n12132_, new_n12133_, new_n12134_,
    new_n12135_, new_n12136_, new_n12137_, new_n12138_, new_n12139_,
    new_n12140_, new_n12141_, new_n12142_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12156_, new_n12157_, new_n12158_, new_n12159_,
    new_n12160_, new_n12161_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12171_, new_n12172_, new_n12173_, new_n12174_,
    new_n12175_, new_n12176_, new_n12177_, new_n12178_, new_n12179_,
    new_n12180_, new_n12181_, new_n12182_, new_n12183_, new_n12184_,
    new_n12185_, new_n12186_, new_n12187_, new_n12188_, new_n12189_,
    new_n12190_, new_n12191_, new_n12192_, new_n12193_, new_n12194_,
    new_n12195_, new_n12196_, new_n12197_, new_n12198_, new_n12199_,
    new_n12200_, new_n12201_, new_n12202_, new_n12203_, new_n12204_,
    new_n12205_, new_n12206_, new_n12207_, new_n12208_, new_n12209_,
    new_n12210_, new_n12211_, new_n12212_, new_n12213_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12220_, new_n12221_,
    new_n12222_, new_n12223_, new_n12224_, new_n12225_, new_n12226_,
    new_n12227_, new_n12228_, new_n12229_, new_n12230_, new_n12231_,
    new_n12232_, new_n12233_, new_n12234_, new_n12235_, new_n12236_,
    new_n12237_, new_n12238_, new_n12239_, new_n12240_, new_n12241_,
    new_n12242_, new_n12243_, new_n12244_, new_n12245_, new_n12246_,
    new_n12247_, new_n12248_, new_n12249_, new_n12250_, new_n12251_,
    new_n12252_, new_n12253_, new_n12254_, new_n12255_, new_n12256_,
    new_n12257_, new_n12258_, new_n12259_, new_n12260_, new_n12261_,
    new_n12262_, new_n12263_, new_n12264_, new_n12265_, new_n12266_,
    new_n12267_, new_n12268_, new_n12269_, new_n12270_, new_n12271_,
    new_n12272_, new_n12273_, new_n12274_, new_n12275_, new_n12276_,
    new_n12277_, new_n12278_, new_n12279_, new_n12280_, new_n12281_,
    new_n12282_, new_n12283_, new_n12284_, new_n12285_, new_n12286_,
    new_n12287_, new_n12288_, new_n12289_, new_n12290_, new_n12291_,
    new_n12292_, new_n12293_, new_n12294_, new_n12295_, new_n12296_,
    new_n12297_, new_n12298_, new_n12299_, new_n12300_, new_n12301_,
    new_n12302_, new_n12303_, new_n12304_, new_n12305_, new_n12306_,
    new_n12307_, new_n12308_, new_n12309_, new_n12310_, new_n12311_,
    new_n12312_, new_n12313_, new_n12314_, new_n12315_, new_n12316_,
    new_n12317_, new_n12318_, new_n12319_, new_n12320_, new_n12321_,
    new_n12322_, new_n12323_, new_n12324_, new_n12325_, new_n12326_,
    new_n12327_, new_n12328_, new_n12329_, new_n12330_, new_n12331_,
    new_n12332_, new_n12333_, new_n12334_, new_n12335_, new_n12336_,
    new_n12337_, new_n12338_, new_n12339_, new_n12340_, new_n12341_,
    new_n12342_, new_n12343_, new_n12344_, new_n12345_, new_n12346_,
    new_n12347_, new_n12348_, new_n12349_, new_n12350_, new_n12351_,
    new_n12352_, new_n12353_, new_n12354_, new_n12355_, new_n12356_,
    new_n12357_, new_n12358_, new_n12360_, new_n12361_, new_n12362_,
    new_n12363_, new_n12364_, new_n12365_, new_n12366_, new_n12367_,
    new_n12368_, new_n12369_, new_n12370_, new_n12371_, new_n12372_,
    new_n12373_, new_n12374_, new_n12375_, new_n12376_, new_n12377_,
    new_n12378_, new_n12379_, new_n12380_, new_n12381_, new_n12382_,
    new_n12383_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12389_, new_n12390_, new_n12391_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12396_, new_n12397_,
    new_n12398_, new_n12399_, new_n12401_, new_n12402_, new_n12403_,
    new_n12404_, new_n12405_, new_n12406_, new_n12407_, new_n12408_,
    new_n12409_, new_n12410_, new_n12411_, new_n12412_, new_n12413_,
    new_n12414_, new_n12415_, new_n12416_, new_n12417_, new_n12418_,
    new_n12419_, new_n12420_, new_n12421_, new_n12422_, new_n12423_,
    new_n12424_, new_n12425_, new_n12426_, new_n12427_, new_n12428_,
    new_n12429_, new_n12430_, new_n12431_, new_n12432_, new_n12433_,
    new_n12434_, new_n12435_, new_n12436_, new_n12437_, new_n12438_,
    new_n12439_, new_n12440_, new_n12441_, new_n12442_, new_n12443_,
    new_n12444_, new_n12445_, new_n12446_, new_n12447_, new_n12448_,
    new_n12449_, new_n12450_, new_n12451_, new_n12452_, new_n12453_,
    new_n12454_, new_n12455_, new_n12456_, new_n12457_, new_n12458_,
    new_n12459_, new_n12460_, new_n12461_, new_n12462_, new_n12463_,
    new_n12464_, new_n12465_, new_n12466_, new_n12467_, new_n12468_,
    new_n12469_, new_n12470_, new_n12471_, new_n12472_, new_n12473_,
    new_n12474_, new_n12475_, new_n12476_, new_n12477_, new_n12478_,
    new_n12479_, new_n12480_, new_n12481_, new_n12482_, new_n12484_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12491_, new_n12492_, new_n12493_, new_n12494_,
    new_n12495_, new_n12496_, new_n12497_, new_n12498_, new_n12499_,
    new_n12500_, new_n12501_, new_n12502_, new_n12503_, new_n12504_,
    new_n12505_, new_n12506_, new_n12507_, new_n12508_, new_n12509_,
    new_n12510_, new_n12511_, new_n12512_, new_n12513_, new_n12514_,
    new_n12515_, new_n12516_, new_n12517_, new_n12518_, new_n12519_,
    new_n12520_, new_n12521_, new_n12522_, new_n12523_, new_n12524_,
    new_n12525_, new_n12526_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12532_, new_n12533_, new_n12534_,
    new_n12535_, new_n12536_, new_n12537_, new_n12538_, new_n12539_,
    new_n12540_, new_n12541_, new_n12542_, new_n12543_, new_n12544_,
    new_n12545_, new_n12546_, new_n12547_, new_n12548_, new_n12549_,
    new_n12550_, new_n12551_, new_n12552_, new_n12553_, new_n12554_,
    new_n12555_, new_n12556_, new_n12557_, new_n12558_, new_n12559_,
    new_n12560_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12616_,
    new_n12617_, new_n12618_, new_n12619_, new_n12620_, new_n12621_,
    new_n12622_, new_n12624_, new_n12625_, new_n12626_, new_n12627_,
    new_n12628_, new_n12629_, new_n12630_, new_n12631_, new_n12632_,
    new_n12633_, new_n12634_, new_n12635_, new_n12636_, new_n12637_,
    new_n12638_, new_n12639_, new_n12640_, new_n12641_, new_n12642_,
    new_n12643_, new_n12644_, new_n12645_, new_n12646_, new_n12647_,
    new_n12648_, new_n12649_, new_n12650_, new_n12651_, new_n12652_,
    new_n12653_, new_n12654_, new_n12655_, new_n12656_, new_n12657_,
    new_n12658_, new_n12659_, new_n12660_, new_n12661_, new_n12662_,
    new_n12663_, new_n12664_, new_n12665_, new_n12666_, new_n12667_,
    new_n12668_, new_n12669_, new_n12670_, new_n12671_, new_n12672_,
    new_n12673_, new_n12674_, new_n12675_, new_n12676_, new_n12677_,
    new_n12678_, new_n12679_, new_n12680_, new_n12681_, new_n12682_,
    new_n12683_, new_n12684_, new_n12685_, new_n12686_, new_n12687_,
    new_n12688_, new_n12689_, new_n12690_, new_n12691_, new_n12692_,
    new_n12693_, new_n12695_, new_n12696_, new_n12697_, new_n12698_,
    new_n12699_, new_n12700_, new_n12701_, new_n12702_, new_n12703_,
    new_n12704_, new_n12705_, new_n12706_, new_n12707_, new_n12708_,
    new_n12709_, new_n12710_, new_n12711_, new_n12712_, new_n12713_,
    new_n12714_, new_n12715_, new_n12716_, new_n12717_, new_n12718_,
    new_n12719_, new_n12720_, new_n12721_, new_n12722_, new_n12723_,
    new_n12724_, new_n12725_, new_n12726_, new_n12727_, new_n12728_,
    new_n12729_, new_n12730_, new_n12731_, new_n12732_, new_n12733_,
    new_n12734_, new_n12735_, new_n12736_, new_n12738_, new_n12739_,
    new_n12740_, new_n12741_, new_n12742_, new_n12743_, new_n12744_,
    new_n12745_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12754_,
    new_n12755_, new_n12756_, new_n12757_, new_n12758_, new_n12759_,
    new_n12760_, new_n12761_, new_n12762_, new_n12763_, new_n12764_,
    new_n12765_, new_n12766_, new_n12767_, new_n12768_, new_n12769_,
    new_n12770_, new_n12771_, new_n12772_, new_n12773_, new_n12774_,
    new_n12775_, new_n12776_, new_n12777_, new_n12778_, new_n12779_,
    new_n12780_, new_n12781_, new_n12782_, new_n12783_, new_n12784_,
    new_n12785_, new_n12786_, new_n12787_, new_n12788_, new_n12789_,
    new_n12790_, new_n12791_, new_n12792_, new_n12793_, new_n12794_,
    new_n12795_, new_n12796_, new_n12797_, new_n12798_, new_n12799_,
    new_n12800_, new_n12801_, new_n12802_, new_n12803_, new_n12804_,
    new_n12805_, new_n12806_, new_n12807_, new_n12808_, new_n12809_,
    new_n12810_, new_n12811_, new_n12812_, new_n12813_, new_n12814_,
    new_n12815_, new_n12816_, new_n12817_, new_n12818_, new_n12819_,
    new_n12820_, new_n12821_, new_n12822_, new_n12823_, new_n12824_,
    new_n12825_, new_n12826_, new_n12827_, new_n12828_, new_n12829_,
    new_n12830_, new_n12831_, new_n12832_, new_n12833_, new_n12834_,
    new_n12835_, new_n12836_, new_n12837_, new_n12838_, new_n12839_,
    new_n12840_, new_n12841_, new_n12842_, new_n12843_, new_n12844_,
    new_n12845_, new_n12846_, new_n12847_, new_n12848_, new_n12849_,
    new_n12850_, new_n12851_, new_n12852_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12863_, new_n12864_,
    new_n12865_, new_n12866_, new_n12867_, new_n12868_, new_n12869_,
    new_n12870_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12875_, new_n12876_, new_n12877_, new_n12878_, new_n12879_,
    new_n12880_, new_n12881_, new_n12882_, new_n12883_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12889_,
    new_n12890_, new_n12891_, new_n12892_, new_n12893_, new_n12894_,
    new_n12895_, new_n12896_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13560_,
    new_n13561_, new_n13562_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13626_, new_n13627_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13638_, new_n13639_, new_n13640_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13655_,
    new_n13656_, new_n13657_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13668_, new_n13669_, new_n13670_,
    new_n13671_, new_n13672_, new_n13673_, new_n13674_, new_n13675_,
    new_n13676_, new_n13677_, new_n13678_, new_n13679_, new_n13680_,
    new_n13681_, new_n13682_, new_n13683_, new_n13684_, new_n13685_,
    new_n13686_, new_n13687_, new_n13688_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13750_,
    new_n13751_, new_n13752_, new_n13753_, new_n13754_, new_n13755_,
    new_n13756_, new_n13757_, new_n13758_, new_n13759_, new_n13760_,
    new_n13761_, new_n13762_, new_n13763_, new_n13764_, new_n13765_,
    new_n13766_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13776_, new_n13777_, new_n13778_, new_n13779_, new_n13780_,
    new_n13781_, new_n13782_, new_n13783_, new_n13784_, new_n13785_,
    new_n13786_, new_n13787_, new_n13788_, new_n13789_, new_n13790_,
    new_n13791_, new_n13792_, new_n13793_, new_n13794_, new_n13795_,
    new_n13796_, new_n13797_, new_n13798_, new_n13799_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13815_,
    new_n13816_, new_n13817_, new_n13818_, new_n13819_, new_n13820_,
    new_n13821_, new_n13822_, new_n13823_, new_n13824_, new_n13825_,
    new_n13826_, new_n13827_, new_n13828_, new_n13829_, new_n13830_,
    new_n13831_, new_n13832_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13898_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13968_, new_n13969_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13975_, new_n13976_,
    new_n13977_, new_n13978_, new_n13979_, new_n13980_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13985_, new_n13986_,
    new_n13987_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14194_, new_n14195_, new_n14196_,
    new_n14197_, new_n14198_, new_n14199_, new_n14200_, new_n14201_,
    new_n14202_, new_n14203_, new_n14204_, new_n14205_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14257_, new_n14258_, new_n14259_, new_n14260_, new_n14261_,
    new_n14262_, new_n14263_, new_n14264_, new_n14265_, new_n14266_,
    new_n14267_, new_n14268_, new_n14269_, new_n14270_, new_n14271_,
    new_n14272_, new_n14273_, new_n14274_, new_n14275_, new_n14276_,
    new_n14277_, new_n14278_, new_n14279_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14299_, new_n14300_, new_n14301_, new_n14302_,
    new_n14303_, new_n14304_, new_n14305_, new_n14306_, new_n14307_,
    new_n14308_, new_n14309_, new_n14310_, new_n14311_, new_n14312_,
    new_n14313_, new_n14314_, new_n14315_, new_n14316_, new_n14317_,
    new_n14318_, new_n14319_, new_n14320_, new_n14321_, new_n14322_,
    new_n14323_, new_n14324_, new_n14325_, new_n14326_, new_n14327_,
    new_n14328_, new_n14329_, new_n14330_, new_n14331_, new_n14332_,
    new_n14333_, new_n14334_, new_n14335_, new_n14336_, new_n14337_,
    new_n14338_, new_n14339_, new_n14340_, new_n14341_, new_n14342_,
    new_n14343_, new_n14344_, new_n14345_, new_n14346_, new_n14347_,
    new_n14348_, new_n14349_, new_n14350_, new_n14351_, new_n14352_,
    new_n14353_, new_n14354_, new_n14355_, new_n14356_, new_n14357_,
    new_n14358_, new_n14359_, new_n14360_, new_n14361_, new_n14362_,
    new_n14363_, new_n14364_, new_n14365_, new_n14366_, new_n14367_,
    new_n14368_, new_n14369_, new_n14370_, new_n14371_, new_n14372_,
    new_n14373_, new_n14374_, new_n14375_, new_n14376_, new_n14377_,
    new_n14378_, new_n14379_, new_n14380_, new_n14381_, new_n14382_,
    new_n14383_, new_n14384_, new_n14385_, new_n14386_, new_n14387_,
    new_n14388_, new_n14389_, new_n14390_, new_n14391_, new_n14392_,
    new_n14393_, new_n14394_, new_n14395_, new_n14396_, new_n14397_,
    new_n14398_, new_n14399_, new_n14400_, new_n14401_, new_n14402_,
    new_n14403_, new_n14404_, new_n14405_, new_n14406_, new_n14407_,
    new_n14408_, new_n14409_, new_n14410_, new_n14411_, new_n14412_,
    new_n14413_, new_n14414_, new_n14415_, new_n14416_, new_n14417_,
    new_n14418_, new_n14419_, new_n14420_, new_n14421_, new_n14422_,
    new_n14423_, new_n14424_, new_n14425_, new_n14426_, new_n14427_,
    new_n14428_, new_n14429_, new_n14430_, new_n14431_, new_n14432_,
    new_n14433_, new_n14434_, new_n14435_, new_n14436_, new_n14437_,
    new_n14438_, new_n14439_, new_n14440_, new_n14441_, new_n14442_,
    new_n14443_, new_n14444_, new_n14445_, new_n14446_, new_n14447_,
    new_n14448_, new_n14449_, new_n14450_, new_n14451_, new_n14452_,
    new_n14453_, new_n14454_, new_n14455_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14486_, new_n14487_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14496_, new_n14497_,
    new_n14498_, new_n14499_, new_n14500_, new_n14501_, new_n14502_,
    new_n14503_, new_n14504_, new_n14505_, new_n14506_, new_n14507_,
    new_n14508_, new_n14509_, new_n14510_, new_n14511_, new_n14512_,
    new_n14513_, new_n14514_, new_n14515_, new_n14516_, new_n14517_,
    new_n14518_, new_n14519_, new_n14520_, new_n14521_, new_n14522_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14539_, new_n14540_, new_n14541_, new_n14542_,
    new_n14543_, new_n14544_, new_n14545_, new_n14546_, new_n14547_,
    new_n14548_, new_n14549_, new_n14550_, new_n14551_, new_n14552_,
    new_n14553_, new_n14554_, new_n14555_, new_n14556_, new_n14557_,
    new_n14558_, new_n14559_, new_n14560_, new_n14561_, new_n14562_,
    new_n14563_, new_n14564_, new_n14565_, new_n14566_, new_n14567_,
    new_n14568_, new_n14569_, new_n14570_, new_n14571_, new_n14572_,
    new_n14573_, new_n14574_, new_n14575_, new_n14576_, new_n14577_,
    new_n14578_, new_n14579_, new_n14580_, new_n14581_, new_n14582_,
    new_n14583_, new_n14584_, new_n14585_, new_n14586_, new_n14587_,
    new_n14588_, new_n14589_, new_n14590_, new_n14591_, new_n14592_,
    new_n14593_, new_n14594_, new_n14595_, new_n14596_, new_n14597_,
    new_n14598_, new_n14599_, new_n14600_, new_n14601_, new_n14602_,
    new_n14603_, new_n14604_, new_n14605_, new_n14606_, new_n14607_,
    new_n14608_, new_n14609_, new_n14610_, new_n14611_, new_n14612_,
    new_n14613_, new_n14614_, new_n14615_, new_n14616_, new_n14617_,
    new_n14618_, new_n14619_, new_n14620_, new_n14621_, new_n14622_,
    new_n14623_, new_n14624_, new_n14625_, new_n14626_, new_n14627_,
    new_n14628_, new_n14629_, new_n14630_, new_n14631_, new_n14632_,
    new_n14633_, new_n14634_, new_n14635_, new_n14636_, new_n14637_,
    new_n14638_, new_n14639_, new_n14640_, new_n14641_, new_n14642_,
    new_n14643_, new_n14644_, new_n14645_, new_n14646_, new_n14647_,
    new_n14648_, new_n14649_, new_n14650_, new_n14651_, new_n14652_,
    new_n14653_, new_n14654_, new_n14655_, new_n14656_, new_n14657_,
    new_n14658_, new_n14659_, new_n14660_, new_n14661_, new_n14662_,
    new_n14663_, new_n14664_, new_n14665_, new_n14666_, new_n14667_,
    new_n14668_, new_n14669_, new_n14670_, new_n14671_, new_n14672_,
    new_n14673_, new_n14674_, new_n14675_, new_n14676_, new_n14677_,
    new_n14678_, new_n14679_, new_n14680_, new_n14681_, new_n14682_,
    new_n14683_, new_n14684_, new_n14685_, new_n14686_, new_n14687_,
    new_n14688_, new_n14689_, new_n14690_, new_n14691_, new_n14692_,
    new_n14693_, new_n14694_, new_n14695_, new_n14696_, new_n14697_,
    new_n14698_, new_n14699_, new_n14700_, new_n14701_, new_n14702_,
    new_n14703_, new_n14704_, new_n14705_, new_n14706_, new_n14707_,
    new_n14708_, new_n14709_, new_n14710_, new_n14711_, new_n14712_,
    new_n14713_, new_n14714_, new_n14715_, new_n14716_, new_n14717_,
    new_n14718_, new_n14719_, new_n14720_, new_n14721_, new_n14722_,
    new_n14723_, new_n14724_, new_n14725_, new_n14726_, new_n14727_,
    new_n14728_, new_n14729_, new_n14730_, new_n14731_, new_n14732_,
    new_n14733_, new_n14734_, new_n14735_, new_n14736_, new_n14737_,
    new_n14738_, new_n14739_, new_n14740_, new_n14741_, new_n14742_,
    new_n14743_, new_n14744_, new_n14745_, new_n14746_, new_n14747_,
    new_n14748_, new_n14749_, new_n14750_, new_n14751_, new_n14752_,
    new_n14753_, new_n14754_, new_n14755_, new_n14756_, new_n14757_,
    new_n14758_, new_n14759_, new_n14760_, new_n14761_, new_n14762_,
    new_n14763_, new_n14764_, new_n14765_, new_n14766_, new_n14767_,
    new_n14768_, new_n14769_, new_n14770_, new_n14771_, new_n14772_,
    new_n14773_, new_n14774_, new_n14775_, new_n14776_, new_n14777_,
    new_n14778_, new_n14779_, new_n14780_, new_n14781_, new_n14782_,
    new_n14783_, new_n14784_, new_n14785_, new_n14786_, new_n14787_,
    new_n14788_, new_n14789_, new_n14790_, new_n14791_, new_n14792_,
    new_n14793_, new_n14794_, new_n14795_, new_n14796_, new_n14797_,
    new_n14798_, new_n14799_, new_n14800_, new_n14801_, new_n14802_,
    new_n14803_, new_n14804_, new_n14805_, new_n14806_, new_n14807_,
    new_n14808_, new_n14809_, new_n14810_, new_n14811_, new_n14812_,
    new_n14813_, new_n14814_, new_n14815_, new_n14816_, new_n14817_,
    new_n14818_, new_n14819_, new_n14820_, new_n14821_, new_n14822_,
    new_n14823_, new_n14824_, new_n14825_, new_n14826_, new_n14827_,
    new_n14828_, new_n14829_, new_n14830_, new_n14831_, new_n14832_,
    new_n14833_, new_n14834_, new_n14835_, new_n14836_, new_n14837_,
    new_n14838_, new_n14839_, new_n14840_, new_n14841_, new_n14842_,
    new_n14843_, new_n14844_, new_n14845_, new_n14846_, new_n14847_,
    new_n14849_, new_n14850_, new_n14851_, new_n14852_, new_n14853_,
    new_n14854_, new_n14855_, new_n14856_, new_n14857_, new_n14858_,
    new_n14859_, new_n14860_, new_n14861_, new_n14862_, new_n14863_,
    new_n14864_, new_n14865_, new_n14866_, new_n14867_, new_n14868_,
    new_n14869_, new_n14870_, new_n14871_, new_n14872_, new_n14873_,
    new_n14874_, new_n14875_, new_n14876_, new_n14877_, new_n14878_,
    new_n14879_, new_n14880_, new_n14881_, new_n14882_, new_n14883_,
    new_n14884_, new_n14885_, new_n14886_, new_n14887_, new_n14888_,
    new_n14889_, new_n14890_, new_n14891_, new_n14892_, new_n14893_,
    new_n14894_, new_n14895_, new_n14896_, new_n14897_, new_n14898_,
    new_n14899_, new_n14900_, new_n14901_, new_n14902_, new_n14903_,
    new_n14904_, new_n14905_, new_n14906_, new_n14907_, new_n14908_,
    new_n14909_, new_n14910_, new_n14911_, new_n14912_, new_n14913_,
    new_n14914_, new_n14915_, new_n14916_, new_n14917_, new_n14918_,
    new_n14919_, new_n14920_, new_n14921_, new_n14922_, new_n14923_,
    new_n14924_, new_n14925_, new_n14926_, new_n14927_, new_n14928_,
    new_n14929_, new_n14930_, new_n14931_, new_n14932_, new_n14933_,
    new_n14934_, new_n14935_, new_n14936_, new_n14937_, new_n14938_,
    new_n14939_, new_n14940_, new_n14941_, new_n14942_, new_n14943_,
    new_n14944_, new_n14945_, new_n14946_, new_n14947_, new_n14948_,
    new_n14949_, new_n14950_, new_n14951_, new_n14952_, new_n14953_,
    new_n14954_, new_n14955_, new_n14956_, new_n14957_, new_n14958_,
    new_n14959_, new_n14960_, new_n14961_, new_n14962_, new_n14963_,
    new_n14964_, new_n14965_, new_n14966_, new_n14967_, new_n14968_,
    new_n14969_, new_n14970_, new_n14971_, new_n14972_, new_n14973_,
    new_n14974_, new_n14975_, new_n14976_, new_n14977_, new_n14978_,
    new_n14979_, new_n14980_, new_n14981_, new_n14982_, new_n14983_,
    new_n14984_, new_n14985_, new_n14986_, new_n14987_, new_n14988_,
    new_n14989_, new_n14990_, new_n14991_, new_n14992_, new_n14993_,
    new_n14994_, new_n14995_, new_n14996_, new_n14997_, new_n14998_,
    new_n14999_, new_n15000_, new_n15001_, new_n15002_, new_n15003_,
    new_n15004_, new_n15005_, new_n15006_, new_n15007_, new_n15008_,
    new_n15009_, new_n15010_, new_n15011_, new_n15012_, new_n15013_,
    new_n15014_, new_n15015_, new_n15016_, new_n15017_, new_n15018_,
    new_n15019_, new_n15020_, new_n15021_, new_n15022_, new_n15023_,
    new_n15024_, new_n15025_, new_n15026_, new_n15027_, new_n15028_,
    new_n15029_, new_n15030_, new_n15031_, new_n15032_, new_n15033_,
    new_n15034_, new_n15035_, new_n15036_, new_n15037_, new_n15038_,
    new_n15039_, new_n15040_, new_n15041_, new_n15042_, new_n15043_,
    new_n15044_, new_n15045_, new_n15046_, new_n15047_, new_n15048_,
    new_n15049_, new_n15050_, new_n15051_, new_n15052_, new_n15053_,
    new_n15054_, new_n15055_, new_n15056_, new_n15057_, new_n15058_,
    new_n15059_, new_n15060_, new_n15061_, new_n15062_, new_n15063_,
    new_n15064_, new_n15065_, new_n15066_, new_n15067_, new_n15068_,
    new_n15069_, new_n15070_, new_n15071_, new_n15072_, new_n15073_,
    new_n15074_, new_n15075_, new_n15076_, new_n15077_, new_n15078_,
    new_n15079_, new_n15080_, new_n15081_, new_n15082_, new_n15083_,
    new_n15084_, new_n15085_, new_n15086_, new_n15087_, new_n15088_,
    new_n15089_, new_n15090_, new_n15091_, new_n15092_, new_n15093_,
    new_n15094_, new_n15095_, new_n15096_, new_n15097_, new_n15098_,
    new_n15099_, new_n15100_, new_n15101_, new_n15102_, new_n15103_,
    new_n15104_, new_n15105_, new_n15106_, new_n15107_, new_n15108_,
    new_n15109_, new_n15110_, new_n15111_, new_n15112_, new_n15113_,
    new_n15114_, new_n15115_, new_n15116_, new_n15117_, new_n15118_,
    new_n15119_, new_n15120_, new_n15121_, new_n15122_, new_n15123_,
    new_n15124_, new_n15125_, new_n15126_, new_n15127_, new_n15128_,
    new_n15129_, new_n15130_, new_n15131_, new_n15132_, new_n15133_,
    new_n15134_, new_n15135_, new_n15136_, new_n15137_, new_n15138_,
    new_n15139_, new_n15140_, new_n15141_, new_n15142_, new_n15143_,
    new_n15144_, new_n15145_, new_n15146_, new_n15147_, new_n15148_,
    new_n15149_, new_n15150_, new_n15151_, new_n15152_, new_n15153_,
    new_n15154_, new_n15155_, new_n15156_, new_n15157_, new_n15158_,
    new_n15159_, new_n15160_, new_n15161_, new_n15162_, new_n15163_,
    new_n15164_, new_n15165_, new_n15166_, new_n15167_, new_n15168_,
    new_n15169_, new_n15170_, new_n15171_, new_n15172_, new_n15173_,
    new_n15174_, new_n15175_, new_n15176_, new_n15177_, new_n15178_,
    new_n15179_, new_n15180_, new_n15181_, new_n15182_, new_n15183_,
    new_n15184_, new_n15185_, new_n15186_, new_n15187_, new_n15188_,
    new_n15189_, new_n15190_, new_n15191_, new_n15192_, new_n15193_,
    new_n15194_, new_n15195_, new_n15196_, new_n15197_, new_n15198_,
    new_n15199_, new_n15200_, new_n15201_, new_n15202_, new_n15203_,
    new_n15204_, new_n15205_, new_n15206_, new_n15207_, new_n15208_,
    new_n15209_, new_n15210_, new_n15211_, new_n15212_, new_n15213_,
    new_n15215_, new_n15216_, new_n15217_, new_n15218_, new_n15219_,
    new_n15220_, new_n15221_, new_n15222_, new_n15223_, new_n15224_,
    new_n15225_, new_n15226_, new_n15227_, new_n15228_, new_n15229_,
    new_n15230_, new_n15231_, new_n15232_, new_n15233_, new_n15234_,
    new_n15235_, new_n15236_, new_n15237_, new_n15238_, new_n15239_,
    new_n15240_, new_n15241_, new_n15242_, new_n15243_, new_n15244_,
    new_n15245_, new_n15246_, new_n15247_, new_n15248_, new_n15249_,
    new_n15250_, new_n15251_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15267_, new_n15268_, new_n15269_,
    new_n15270_, new_n15271_, new_n15272_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15300_, new_n15301_, new_n15302_, new_n15303_, new_n15304_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15335_, new_n15336_, new_n15337_, new_n15338_, new_n15339_,
    new_n15340_, new_n15341_, new_n15342_, new_n15343_, new_n15344_,
    new_n15345_, new_n15346_, new_n15347_, new_n15348_, new_n15349_,
    new_n15350_, new_n15351_, new_n15352_, new_n15353_, new_n15354_,
    new_n15355_, new_n15356_, new_n15357_, new_n15358_, new_n15359_,
    new_n15360_, new_n15361_, new_n15362_, new_n15363_, new_n15364_,
    new_n15365_, new_n15366_, new_n15367_, new_n15368_, new_n15369_,
    new_n15370_, new_n15371_, new_n15372_, new_n15373_, new_n15374_,
    new_n15375_, new_n15376_, new_n15377_, new_n15378_, new_n15379_,
    new_n15380_, new_n15381_, new_n15382_, new_n15383_, new_n15384_,
    new_n15385_, new_n15386_, new_n15387_, new_n15388_, new_n15389_,
    new_n15390_, new_n15391_, new_n15392_, new_n15393_, new_n15394_,
    new_n15395_, new_n15396_, new_n15397_, new_n15398_, new_n15399_,
    new_n15400_, new_n15401_, new_n15402_, new_n15403_, new_n15404_,
    new_n15405_, new_n15406_, new_n15407_, new_n15408_, new_n15409_,
    new_n15410_, new_n15411_, new_n15412_, new_n15413_, new_n15414_,
    new_n15415_, new_n15416_, new_n15417_, new_n15418_, new_n15419_,
    new_n15420_, new_n15421_, new_n15422_, new_n15423_, new_n15424_,
    new_n15425_, new_n15426_, new_n15427_, new_n15428_, new_n15429_,
    new_n15430_, new_n15431_, new_n15432_, new_n15433_, new_n15434_,
    new_n15435_, new_n15436_, new_n15437_, new_n15438_, new_n15439_,
    new_n15440_, new_n15441_, new_n15442_, new_n15443_, new_n15444_,
    new_n15445_, new_n15446_, new_n15447_, new_n15448_, new_n15449_,
    new_n15450_, new_n15451_, new_n15452_, new_n15453_, new_n15454_,
    new_n15455_, new_n15456_, new_n15457_, new_n15458_, new_n15459_,
    new_n15460_, new_n15461_, new_n15462_, new_n15463_, new_n15464_,
    new_n15465_, new_n15466_, new_n15467_, new_n15468_, new_n15469_,
    new_n15470_, new_n15471_, new_n15472_, new_n15473_, new_n15474_,
    new_n15475_, new_n15476_, new_n15477_, new_n15478_, new_n15479_,
    new_n15480_, new_n15481_, new_n15482_, new_n15483_, new_n15484_,
    new_n15485_, new_n15486_, new_n15487_, new_n15488_, new_n15489_,
    new_n15490_, new_n15491_, new_n15492_, new_n15493_, new_n15494_,
    new_n15495_, new_n15496_, new_n15497_, new_n15498_, new_n15499_,
    new_n15500_, new_n15501_, new_n15502_, new_n15503_, new_n15504_,
    new_n15505_, new_n15506_, new_n15507_, new_n15508_, new_n15509_,
    new_n15510_, new_n15511_, new_n15512_, new_n15513_, new_n15514_,
    new_n15515_, new_n15516_, new_n15517_, new_n15518_, new_n15519_,
    new_n15520_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15526_, new_n15527_, new_n15528_, new_n15529_,
    new_n15530_, new_n15531_, new_n15532_, new_n15533_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15545_, new_n15546_, new_n15547_, new_n15548_, new_n15549_,
    new_n15550_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15562_, new_n15563_, new_n15564_,
    new_n15565_, new_n15566_, new_n15567_, new_n15568_, new_n15569_,
    new_n15570_, new_n15571_, new_n15572_, new_n15573_, new_n15574_,
    new_n15576_, new_n15577_, new_n15578_, new_n15579_, new_n15580_,
    new_n15581_, new_n15582_, new_n15583_, new_n15584_, new_n15585_,
    new_n15586_, new_n15587_, new_n15588_, new_n15589_, new_n15590_,
    new_n15591_, new_n15592_, new_n15593_, new_n15594_, new_n15595_,
    new_n15596_, new_n15597_, new_n15598_, new_n15599_, new_n15600_,
    new_n15601_, new_n15602_, new_n15603_, new_n15604_, new_n15605_,
    new_n15606_, new_n15607_, new_n15608_, new_n15609_, new_n15610_,
    new_n15611_, new_n15612_, new_n15613_, new_n15614_, new_n15615_,
    new_n15616_, new_n15617_, new_n15618_, new_n15619_, new_n15620_,
    new_n15621_, new_n15622_, new_n15623_, new_n15624_, new_n15625_,
    new_n15626_, new_n15627_, new_n15628_, new_n15629_, new_n15630_,
    new_n15631_, new_n15632_, new_n15633_, new_n15634_, new_n15635_,
    new_n15636_, new_n15637_, new_n15638_, new_n15639_, new_n15640_,
    new_n15641_, new_n15642_, new_n15643_, new_n15644_, new_n15645_,
    new_n15646_, new_n15647_, new_n15648_, new_n15649_, new_n15650_,
    new_n15651_, new_n15652_, new_n15653_, new_n15654_, new_n15655_,
    new_n15656_, new_n15657_, new_n15658_, new_n15659_, new_n15660_,
    new_n15661_, new_n15662_, new_n15663_, new_n15664_, new_n15665_,
    new_n15666_, new_n15667_, new_n15668_, new_n15669_, new_n15670_,
    new_n15671_, new_n15672_, new_n15673_, new_n15674_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15681_, new_n15682_, new_n15683_, new_n15684_, new_n15685_,
    new_n15686_, new_n15687_, new_n15688_, new_n15689_, new_n15690_,
    new_n15691_, new_n15692_, new_n15693_, new_n15694_, new_n15695_,
    new_n15696_, new_n15697_, new_n15698_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15840_,
    new_n15841_, new_n15842_, new_n15843_, new_n15844_, new_n15845_,
    new_n15846_, new_n15847_, new_n15848_, new_n15849_, new_n15850_,
    new_n15851_, new_n15852_, new_n15853_, new_n15854_, new_n15855_,
    new_n15856_, new_n15857_, new_n15858_, new_n15859_, new_n15860_,
    new_n15861_, new_n15862_, new_n15863_, new_n15864_, new_n15865_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15881_, new_n15882_, new_n15883_, new_n15884_, new_n15885_,
    new_n15886_, new_n15887_, new_n15888_, new_n15889_, new_n15890_,
    new_n15891_, new_n15892_, new_n15893_, new_n15894_, new_n15895_,
    new_n15896_, new_n15897_, new_n15898_, new_n15899_, new_n15900_,
    new_n15901_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15931_, new_n15932_, new_n15933_, new_n15934_, new_n15936_,
    new_n15937_, new_n15938_, new_n15939_, new_n15940_, new_n15941_,
    new_n15942_, new_n15943_, new_n15944_, new_n15945_, new_n15946_,
    new_n15947_, new_n15948_, new_n15949_, new_n15950_, new_n15951_,
    new_n15952_, new_n15953_, new_n15954_, new_n15955_, new_n15956_,
    new_n15957_, new_n15958_, new_n15959_, new_n15960_, new_n15961_,
    new_n15962_, new_n15963_, new_n15964_, new_n15965_, new_n15966_,
    new_n15967_, new_n15968_, new_n15969_, new_n15970_, new_n15971_,
    new_n15972_, new_n15973_, new_n15974_, new_n15975_, new_n15976_,
    new_n15977_, new_n15978_, new_n15979_, new_n15980_, new_n15981_,
    new_n15982_, new_n15983_, new_n15984_, new_n15985_, new_n15986_,
    new_n15987_, new_n15988_, new_n15989_, new_n15990_, new_n15991_,
    new_n15993_, new_n15994_, new_n15995_, new_n15996_, new_n15997_,
    new_n15998_, new_n15999_, new_n16000_, new_n16001_, new_n16002_,
    new_n16003_, new_n16004_, new_n16005_, new_n16006_, new_n16007_,
    new_n16008_, new_n16009_, new_n16010_, new_n16011_, new_n16012_,
    new_n16013_, new_n16014_, new_n16015_, new_n16016_, new_n16017_,
    new_n16018_, new_n16019_, new_n16020_, new_n16021_, new_n16022_,
    new_n16023_, new_n16024_, new_n16025_, new_n16026_, new_n16027_,
    new_n16028_, new_n16029_, new_n16030_, new_n16031_, new_n16032_,
    new_n16033_, new_n16034_, new_n16035_, new_n16036_, new_n16037_,
    new_n16038_, new_n16039_, new_n16040_, new_n16041_, new_n16042_,
    new_n16043_, new_n16044_, new_n16045_, new_n16046_, new_n16047_,
    new_n16048_, new_n16049_, new_n16050_, new_n16051_, new_n16052_,
    new_n16053_, new_n16054_, new_n16055_, new_n16056_, new_n16057_,
    new_n16058_, new_n16059_, new_n16060_, new_n16061_, new_n16062_,
    new_n16063_, new_n16064_, new_n16065_, new_n16066_, new_n16067_,
    new_n16068_, new_n16069_, new_n16070_, new_n16071_, new_n16072_,
    new_n16073_, new_n16074_, new_n16075_, new_n16076_, new_n16077_,
    new_n16078_, new_n16079_, new_n16080_, new_n16081_, new_n16082_,
    new_n16083_, new_n16084_, new_n16085_, new_n16086_, new_n16087_,
    new_n16088_, new_n16089_, new_n16090_, new_n16091_, new_n16092_,
    new_n16093_, new_n16094_, new_n16095_, new_n16096_, new_n16097_,
    new_n16098_, new_n16099_, new_n16100_, new_n16101_, new_n16102_,
    new_n16103_, new_n16104_, new_n16105_, new_n16106_, new_n16107_,
    new_n16108_, new_n16109_, new_n16110_, new_n16111_, new_n16112_,
    new_n16113_, new_n16114_, new_n16115_, new_n16116_, new_n16117_,
    new_n16118_, new_n16119_, new_n16120_, new_n16121_, new_n16122_,
    new_n16123_, new_n16124_, new_n16126_, new_n16127_, new_n16128_,
    new_n16129_, new_n16130_, new_n16131_, new_n16132_, new_n16133_,
    new_n16134_, new_n16135_, new_n16136_, new_n16137_, new_n16138_,
    new_n16139_, new_n16140_, new_n16141_, new_n16142_, new_n16143_,
    new_n16144_, new_n16145_, new_n16146_, new_n16147_, new_n16148_,
    new_n16149_, new_n16150_, new_n16151_, new_n16152_, new_n16153_,
    new_n16154_, new_n16155_, new_n16156_, new_n16157_, new_n16158_,
    new_n16159_, new_n16160_, new_n16161_, new_n16162_, new_n16163_,
    new_n16164_, new_n16165_, new_n16166_, new_n16168_, new_n16169_,
    new_n16170_, new_n16171_, new_n16172_, new_n16173_, new_n16174_,
    new_n16175_, new_n16176_, new_n16177_, new_n16178_, new_n16179_,
    new_n16180_, new_n16181_, new_n16182_, new_n16183_, new_n16184_,
    new_n16185_, new_n16186_, new_n16187_, new_n16188_, new_n16189_,
    new_n16190_, new_n16191_, new_n16192_, new_n16193_, new_n16194_,
    new_n16195_, new_n16196_, new_n16197_, new_n16198_, new_n16199_,
    new_n16200_, new_n16201_, new_n16202_, new_n16203_, new_n16204_,
    new_n16205_, new_n16206_, new_n16207_, new_n16208_, new_n16210_,
    new_n16211_, new_n16212_, new_n16213_, new_n16214_, new_n16215_,
    new_n16216_, new_n16217_, new_n16218_, new_n16219_, new_n16220_,
    new_n16221_, new_n16222_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16234_, new_n16235_,
    new_n16236_, new_n16237_, new_n16238_, new_n16239_, new_n16240_,
    new_n16241_, new_n16242_, new_n16243_, new_n16245_, new_n16246_,
    new_n16247_, new_n16248_, new_n16249_, new_n16250_, new_n16251_,
    new_n16252_, new_n16253_, new_n16254_, new_n16255_, new_n16256_,
    new_n16257_, new_n16258_, new_n16259_, new_n16260_, new_n16261_,
    new_n16262_, new_n16263_, new_n16264_, new_n16265_, new_n16266_,
    new_n16267_, new_n16268_, new_n16269_, new_n16270_, new_n16271_,
    new_n16272_, new_n16273_, new_n16274_, new_n16275_, new_n16276_,
    new_n16277_, new_n16278_, new_n16279_, new_n16280_, new_n16281_,
    new_n16282_, new_n16283_, new_n16284_, new_n16285_, new_n16286_,
    new_n16287_, new_n16288_, new_n16289_, new_n16290_, new_n16291_,
    new_n16292_, new_n16293_, new_n16294_, new_n16296_, new_n16297_,
    new_n16298_, new_n16299_, new_n16300_, new_n16301_, new_n16302_,
    new_n16303_, new_n16304_, new_n16305_, new_n16306_, new_n16307_,
    new_n16308_, new_n16309_, new_n16310_, new_n16311_, new_n16312_,
    new_n16313_, new_n16314_, new_n16315_, new_n16316_, new_n16317_,
    new_n16318_, new_n16319_, new_n16320_, new_n16321_, new_n16322_,
    new_n16323_, new_n16324_, new_n16325_, new_n16326_, new_n16327_,
    new_n16328_, new_n16329_, new_n16330_, new_n16331_, new_n16332_,
    new_n16333_, new_n16334_, new_n16335_, new_n16336_, new_n16337_,
    new_n16338_, new_n16339_, new_n16340_, new_n16341_, new_n16342_,
    new_n16343_, new_n16344_, new_n16345_, new_n16346_, new_n16347_,
    new_n16348_, new_n16349_, new_n16350_, new_n16351_, new_n16352_,
    new_n16353_, new_n16354_, new_n16355_, new_n16356_, new_n16357_,
    new_n16358_, new_n16359_, new_n16360_, new_n16361_, new_n16362_,
    new_n16363_, new_n16364_, new_n16365_, new_n16366_, new_n16367_,
    new_n16368_, new_n16369_, new_n16370_, new_n16372_, new_n16373_,
    new_n16374_, new_n16375_, new_n16376_, new_n16377_, new_n16378_,
    new_n16379_, new_n16380_, new_n16381_, new_n16382_, new_n16383_,
    new_n16384_, new_n16385_, new_n16386_, new_n16387_, new_n16388_,
    new_n16389_, new_n16390_, new_n16391_, new_n16392_, new_n16393_,
    new_n16394_, new_n16395_, new_n16396_, new_n16397_, new_n16398_,
    new_n16399_, new_n16400_, new_n16401_, new_n16402_, new_n16403_,
    new_n16404_, new_n16405_, new_n16406_, new_n16407_, new_n16408_,
    new_n16409_, new_n16410_, new_n16411_, new_n16412_, new_n16413_,
    new_n16414_, new_n16415_, new_n16416_, new_n16417_, new_n16418_,
    new_n16419_, new_n16420_, new_n16421_, new_n16422_, new_n16423_,
    new_n16425_, new_n16426_, new_n16427_, new_n16428_, new_n16429_,
    new_n16430_, new_n16431_, new_n16432_, new_n16433_, new_n16434_,
    new_n16435_, new_n16436_, new_n16437_, new_n16438_, new_n16439_,
    new_n16440_, new_n16441_, new_n16442_, new_n16443_, new_n16444_,
    new_n16445_, new_n16446_, new_n16447_, new_n16448_, new_n16449_,
    new_n16450_, new_n16451_, new_n16452_, new_n16453_, new_n16454_,
    new_n16455_, new_n16456_, new_n16457_, new_n16459_, new_n16460_,
    new_n16461_, new_n16462_, new_n16463_, new_n16464_, new_n16465_,
    new_n16466_, new_n16467_, new_n16468_, new_n16469_, new_n16470_,
    new_n16471_, new_n16472_, new_n16473_, new_n16474_, new_n16475_,
    new_n16476_, new_n16477_, new_n16478_, new_n16479_, new_n16480_,
    new_n16481_, new_n16482_, new_n16483_, new_n16484_, new_n16485_,
    new_n16486_, new_n16487_, new_n16488_, new_n16490_, new_n16491_,
    new_n16492_, new_n16493_, new_n16494_, new_n16495_, new_n16496_,
    new_n16497_, new_n16498_, new_n16499_, new_n16500_, new_n16501_,
    new_n16502_, new_n16503_, new_n16504_, new_n16505_, new_n16506_,
    new_n16507_, new_n16508_, new_n16510_, new_n16511_, new_n16512_,
    new_n16513_, new_n16514_, new_n16515_, new_n16516_, new_n16517_,
    new_n16518_, new_n16519_, new_n16520_, new_n16521_, new_n16522_,
    new_n16523_, new_n16524_, new_n16525_, new_n16526_, new_n16527_,
    new_n16528_, new_n16529_, new_n16530_, new_n16531_, new_n16532_,
    new_n16533_, new_n16534_, new_n16535_, new_n16536_, new_n16537_,
    new_n16538_, new_n16539_, new_n16540_, new_n16541_, new_n16542_,
    new_n16543_, new_n16544_, new_n16545_, new_n16546_, new_n16547_,
    new_n16548_, new_n16550_, new_n16551_, new_n16552_, new_n16553_,
    new_n16554_, new_n16555_, new_n16556_, new_n16557_, new_n16558_,
    new_n16559_, new_n16560_, new_n16561_, new_n16562_, new_n16563_,
    new_n16564_, new_n16565_, new_n16566_, new_n16567_, new_n16568_,
    new_n16569_, new_n16570_, new_n16571_, new_n16572_, new_n16573_,
    new_n16574_, new_n16575_, new_n16576_, new_n16577_, new_n16578_,
    new_n16579_, new_n16580_, new_n16581_, new_n16582_, new_n16583_,
    new_n16585_, new_n16586_, new_n16587_, new_n16588_, new_n16589_,
    new_n16590_, new_n16591_, new_n16592_, new_n16593_, new_n16594_,
    new_n16595_, new_n16596_, new_n16597_, new_n16598_, new_n16599_,
    new_n16600_, new_n16601_, new_n16602_, new_n16603_, new_n16604_,
    new_n16605_, new_n16606_, new_n16607_, new_n16608_, new_n16609_,
    new_n16610_, new_n16611_, new_n16612_, new_n16613_, new_n16614_,
    new_n16615_, new_n16616_, new_n16617_, new_n16618_, new_n16620_,
    new_n16621_, new_n16622_, new_n16623_, new_n16624_, new_n16625_,
    new_n16626_, new_n16627_, new_n16628_, new_n16629_, new_n16630_,
    new_n16631_, new_n16632_, new_n16633_, new_n16634_, new_n16635_,
    new_n16636_, new_n16637_, new_n16638_, new_n16639_, new_n16640_,
    new_n16641_, new_n16642_, new_n16643_, new_n16644_, new_n16645_,
    new_n16646_, new_n16647_, new_n16648_, new_n16649_, new_n16650_,
    new_n16651_, new_n16652_, new_n16653_, new_n16654_, new_n16655_,
    new_n16656_, new_n16657_, new_n16658_, new_n16659_, new_n16661_,
    new_n16662_, new_n16663_, new_n16664_, new_n16665_, new_n16666_,
    new_n16667_, new_n16668_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16722_,
    new_n16723_, new_n16724_, new_n16725_, new_n16726_, new_n16727_,
    new_n16728_, new_n16729_, new_n16730_, new_n16731_, new_n16732_,
    new_n16733_, new_n16734_, new_n16735_, new_n16736_, new_n16737_,
    new_n16738_, new_n16739_, new_n16740_, new_n16741_, new_n16742_,
    new_n16743_, new_n16744_, new_n16745_, new_n16746_, new_n16747_,
    new_n16748_, new_n16749_, new_n16750_, new_n16751_, new_n16752_,
    new_n16753_, new_n16754_, new_n16756_, new_n16757_, new_n16758_,
    new_n16759_, new_n16760_, new_n16761_, new_n16762_, new_n16763_,
    new_n16764_, new_n16765_, new_n16766_, new_n16767_, new_n16768_,
    new_n16769_, new_n16770_, new_n16771_, new_n16772_, new_n16773_,
    new_n16774_, new_n16775_, new_n16776_, new_n16777_, new_n16778_,
    new_n16779_, new_n16780_, new_n16781_, new_n16782_, new_n16783_,
    new_n16784_, new_n16785_, new_n16786_, new_n16787_, new_n16788_,
    new_n16789_, new_n16790_, new_n16791_, new_n16792_, new_n16793_,
    new_n16795_, new_n16796_, new_n16797_, new_n16798_, new_n16799_,
    new_n16800_, new_n16801_, new_n16802_, new_n16803_, new_n16804_,
    new_n16805_, new_n16806_, new_n16807_, new_n16808_, new_n16809_,
    new_n16810_, new_n16811_, new_n16812_, new_n16813_, new_n16814_,
    new_n16815_, new_n16816_, new_n16817_, new_n16818_, new_n16819_,
    new_n16821_, new_n16822_, new_n16823_, new_n16824_, new_n16825_,
    new_n16826_, new_n16827_, new_n16828_, new_n16829_, new_n16830_,
    new_n16831_, new_n16832_, new_n16833_, new_n16834_, new_n16835_,
    new_n16836_, new_n16837_, new_n16838_, new_n16839_, new_n16840_,
    new_n16841_, new_n16842_, new_n16844_, new_n16845_, new_n16846_,
    new_n16847_, new_n16848_, new_n16849_, new_n16850_, new_n16851_,
    new_n16852_, new_n16853_, new_n16854_, new_n16855_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16862_, new_n16863_, new_n16864_, new_n16865_, new_n16866_,
    new_n16867_, new_n16868_, new_n16869_, new_n16870_, new_n16871_,
    new_n16872_, new_n16873_, new_n16874_, new_n16875_, new_n16876_,
    new_n16877_, new_n16878_, new_n16879_, new_n16880_, new_n16881_,
    new_n16882_, new_n16883_, new_n16884_, new_n16885_, new_n16886_,
    new_n16887_, new_n16888_, new_n16889_, new_n16890_, new_n16891_,
    new_n16892_, new_n16893_, new_n16894_, new_n16895_, new_n16896_,
    new_n16897_, new_n16898_, new_n16899_, new_n16900_, new_n16901_,
    new_n16902_, new_n16903_, new_n16904_, new_n16906_, new_n16907_,
    new_n16908_, new_n16909_, new_n16910_, new_n16911_, new_n16912_,
    new_n16913_, new_n16914_, new_n16915_, new_n16916_, new_n16917_,
    new_n16918_, new_n16919_, new_n16920_, new_n16921_, new_n16922_,
    new_n16923_, new_n16924_, new_n16925_, new_n16926_, new_n16927_,
    new_n16928_, new_n16929_, new_n16930_, new_n16931_, new_n16933_,
    new_n16934_, new_n16935_, new_n16936_, new_n16937_, new_n16938_,
    new_n16939_, new_n16940_, new_n16941_, new_n16942_, new_n16943_,
    new_n16944_, new_n16945_, new_n16946_, new_n16947_, new_n16948_,
    new_n16949_, new_n16950_, new_n16951_, new_n16952_, new_n16953_,
    new_n16954_, new_n16955_, new_n16956_, new_n16957_, new_n16958_,
    new_n16959_, new_n16960_, new_n16961_, new_n16962_, new_n16963_,
    new_n16964_, new_n16965_, new_n16966_, new_n16967_, new_n16968_,
    new_n16969_, new_n16970_, new_n16971_, new_n16972_, new_n16973_,
    new_n16974_, new_n16975_, new_n16976_, new_n16977_, new_n16978_,
    new_n16979_, new_n16980_, new_n16981_, new_n16982_, new_n16984_,
    new_n16985_, new_n16986_, new_n16987_, new_n16988_, new_n16989_,
    new_n16990_, new_n16991_, new_n16992_, new_n16993_, new_n16994_,
    new_n16995_, new_n16996_, new_n16997_, new_n16998_, new_n16999_,
    new_n17000_, new_n17001_, new_n17002_, new_n17003_, new_n17004_,
    new_n17005_, new_n17006_, new_n17007_, new_n17008_, new_n17009_,
    new_n17010_, new_n17011_, new_n17012_, new_n17013_, new_n17014_,
    new_n17015_, new_n17016_, new_n17017_, new_n17018_, new_n17019_,
    new_n17020_, new_n17021_, new_n17022_, new_n17023_, new_n17024_,
    new_n17025_, new_n17026_, new_n17027_, new_n17028_, new_n17029_,
    new_n17030_, new_n17031_, new_n17032_, new_n17033_, new_n17035_,
    new_n17036_, new_n17037_, new_n17038_, new_n17039_, new_n17040_,
    new_n17041_, new_n17042_, new_n17043_, new_n17044_, new_n17045_,
    new_n17046_, new_n17047_, new_n17048_, new_n17049_, new_n17050_,
    new_n17051_, new_n17052_, new_n17053_, new_n17054_, new_n17055_,
    new_n17056_, new_n17057_, new_n17058_, new_n17059_, new_n17060_,
    new_n17061_, new_n17062_, new_n17063_, new_n17064_, new_n17065_,
    new_n17066_, new_n17067_, new_n17068_, new_n17069_, new_n17070_,
    new_n17071_, new_n17072_, new_n17073_, new_n17074_, new_n17075_,
    new_n17076_, new_n17077_, new_n17078_, new_n17079_, new_n17080_,
    new_n17081_, new_n17082_, new_n17084_, new_n17085_, new_n17086_,
    new_n17087_, new_n17088_, new_n17089_, new_n17090_, new_n17091_,
    new_n17092_, new_n17093_, new_n17094_, new_n17095_, new_n17096_,
    new_n17097_, new_n17098_, new_n17099_, new_n17100_, new_n17101_,
    new_n17102_, new_n17103_, new_n17104_, new_n17105_, new_n17106_,
    new_n17107_, new_n17108_, new_n17109_, new_n17110_, new_n17111_,
    new_n17112_, new_n17113_, new_n17114_, new_n17115_, new_n17116_,
    new_n17117_, new_n17118_, new_n17119_, new_n17120_, new_n17121_,
    new_n17122_, new_n17123_, new_n17124_, new_n17125_, new_n17126_,
    new_n17127_, new_n17128_, new_n17129_, new_n17130_, new_n17131_,
    new_n17132_, new_n17133_, new_n17135_, new_n17136_, new_n17137_,
    new_n17138_, new_n17139_, new_n17140_, new_n17141_, new_n17142_,
    new_n17143_, new_n17144_, new_n17145_, new_n17146_, new_n17147_,
    new_n17148_, new_n17149_, new_n17150_, new_n17151_, new_n17152_,
    new_n17153_, new_n17154_, new_n17155_, new_n17156_, new_n17157_,
    new_n17158_, new_n17159_, new_n17160_, new_n17161_, new_n17162_,
    new_n17163_, new_n17164_, new_n17165_, new_n17166_, new_n17167_,
    new_n17168_, new_n17169_, new_n17170_, new_n17171_, new_n17172_,
    new_n17173_, new_n17174_, new_n17175_, new_n17176_, new_n17177_,
    new_n17178_, new_n17179_, new_n17180_, new_n17181_, new_n17182_,
    new_n17183_, new_n17184_, new_n17185_, new_n17187_, new_n17188_,
    new_n17189_, new_n17190_, new_n17191_, new_n17192_, new_n17193_,
    new_n17194_, new_n17195_, new_n17196_, new_n17197_, new_n17198_,
    new_n17199_, new_n17200_, new_n17201_, new_n17202_, new_n17203_,
    new_n17204_, new_n17205_, new_n17206_, new_n17207_, new_n17208_,
    new_n17209_, new_n17210_, new_n17211_, new_n17212_, new_n17213_,
    new_n17214_, new_n17215_, new_n17216_, new_n17217_, new_n17218_,
    new_n17219_, new_n17220_, new_n17221_, new_n17222_, new_n17223_,
    new_n17224_, new_n17225_, new_n17226_, new_n17227_, new_n17228_,
    new_n17229_, new_n17230_, new_n17231_, new_n17232_, new_n17233_,
    new_n17234_, new_n17235_, new_n17236_, new_n17237_, new_n17238_,
    new_n17239_, new_n17240_, new_n17241_, new_n17242_, new_n17243_,
    new_n17244_, new_n17245_, new_n17246_, new_n17247_, new_n17248_,
    new_n17249_, new_n17250_, new_n17251_, new_n17252_, new_n17253_,
    new_n17254_, new_n17255_, new_n17256_, new_n17257_, new_n17258_,
    new_n17259_, new_n17260_, new_n17261_, new_n17262_, new_n17263_,
    new_n17264_, new_n17265_, new_n17266_, new_n17267_, new_n17268_,
    new_n17269_, new_n17270_, new_n17271_, new_n17272_, new_n17273_,
    new_n17274_, new_n17275_, new_n17276_, new_n17277_, new_n17278_,
    new_n17279_, new_n17280_, new_n17281_, new_n17282_, new_n17283_,
    new_n17284_, new_n17285_, new_n17286_, new_n17287_, new_n17288_,
    new_n17289_, new_n17290_, new_n17291_, new_n17292_, new_n17293_,
    new_n17294_, new_n17295_, new_n17296_, new_n17297_, new_n17298_,
    new_n17299_, new_n17300_, new_n17301_, new_n17302_, new_n17303_,
    new_n17304_, new_n17305_, new_n17306_, new_n17307_, new_n17308_,
    new_n17309_, new_n17310_, new_n17311_, new_n17312_, new_n17313_,
    new_n17314_, new_n17315_, new_n17316_, new_n17317_, new_n17318_,
    new_n17319_, new_n17320_, new_n17321_, new_n17322_, new_n17323_,
    new_n17324_, new_n17325_, new_n17326_, new_n17327_, new_n17328_,
    new_n17329_, new_n17330_, new_n17331_, new_n17332_, new_n17333_,
    new_n17334_, new_n17335_, new_n17336_, new_n17337_, new_n17338_,
    new_n17339_, new_n17340_, new_n17341_, new_n17342_, new_n17343_,
    new_n17344_, new_n17345_, new_n17346_, new_n17347_, new_n17348_,
    new_n17349_, new_n17350_, new_n17351_, new_n17352_, new_n17353_,
    new_n17354_, new_n17355_, new_n17356_, new_n17357_, new_n17358_,
    new_n17359_, new_n17360_, new_n17361_, new_n17362_, new_n17363_,
    new_n17364_, new_n17365_, new_n17366_, new_n17367_, new_n17368_,
    new_n17369_, new_n17370_, new_n17371_, new_n17372_, new_n17373_,
    new_n17374_, new_n17375_, new_n17376_, new_n17377_, new_n17378_,
    new_n17379_, new_n17380_, new_n17381_, new_n17382_, new_n17383_,
    new_n17384_, new_n17385_, new_n17386_, new_n17387_, new_n17388_,
    new_n17389_, new_n17390_, new_n17391_, new_n17392_, new_n17393_,
    new_n17394_, new_n17395_, new_n17396_, new_n17397_, new_n17398_,
    new_n17399_, new_n17400_, new_n17401_, new_n17402_, new_n17403_,
    new_n17404_, new_n17405_, new_n17406_, new_n17407_, new_n17408_,
    new_n17409_, new_n17410_, new_n17411_, new_n17412_, new_n17413_,
    new_n17414_, new_n17415_, new_n17416_, new_n17417_, new_n17418_,
    new_n17419_, new_n17420_, new_n17421_, new_n17422_, new_n17423_,
    new_n17424_, new_n17425_, new_n17426_, new_n17427_, new_n17428_,
    new_n17429_, new_n17430_, new_n17431_, new_n17432_, new_n17433_,
    new_n17434_, new_n17435_, new_n17436_, new_n17437_, new_n17438_,
    new_n17439_, new_n17440_, new_n17441_, new_n17442_, new_n17443_,
    new_n17444_, new_n17445_, new_n17446_, new_n17447_, new_n17448_,
    new_n17449_, new_n17450_, new_n17451_, new_n17452_, new_n17453_,
    new_n17454_, new_n17455_, new_n17456_, new_n17457_, new_n17458_,
    new_n17459_, new_n17460_, new_n17461_, new_n17462_, new_n17463_,
    new_n17464_, new_n17465_, new_n17466_, new_n17467_, new_n17468_,
    new_n17469_, new_n17470_, new_n17471_, new_n17472_, new_n17473_,
    new_n17474_, new_n17475_, new_n17476_, new_n17477_, new_n17478_,
    new_n17479_, new_n17480_, new_n17481_, new_n17482_, new_n17483_,
    new_n17484_, new_n17485_, new_n17486_, new_n17487_, new_n17488_,
    new_n17489_, new_n17490_, new_n17491_, new_n17492_, new_n17493_,
    new_n17494_, new_n17495_, new_n17496_, new_n17497_, new_n17498_,
    new_n17499_, new_n17500_, new_n17501_, new_n17503_, new_n17504_,
    new_n17505_, new_n17506_, new_n17507_, new_n17508_, new_n17509_,
    new_n17510_, new_n17511_, new_n17512_, new_n17513_, new_n17514_,
    new_n17515_, new_n17516_, new_n17517_, new_n17518_, new_n17519_,
    new_n17520_, new_n17521_, new_n17522_, new_n17523_, new_n17524_,
    new_n17525_, new_n17526_, new_n17527_, new_n17528_, new_n17529_,
    new_n17530_, new_n17531_, new_n17532_, new_n17533_, new_n17534_,
    new_n17535_, new_n17536_, new_n17537_, new_n17538_, new_n17539_,
    new_n17540_, new_n17541_, new_n17542_, new_n17543_, new_n17544_,
    new_n17545_, new_n17546_, new_n17547_, new_n17548_, new_n17549_,
    new_n17550_, new_n17551_, new_n17552_, new_n17553_, new_n17554_,
    new_n17555_, new_n17556_, new_n17557_, new_n17558_, new_n17559_,
    new_n17560_, new_n17561_, new_n17562_, new_n17563_, new_n17564_,
    new_n17565_, new_n17566_, new_n17567_, new_n17568_, new_n17569_,
    new_n17570_, new_n17571_, new_n17572_, new_n17573_, new_n17574_,
    new_n17575_, new_n17576_, new_n17577_, new_n17578_, new_n17579_,
    new_n17580_, new_n17581_, new_n17582_, new_n17583_, new_n17584_,
    new_n17585_, new_n17586_, new_n17587_, new_n17588_, new_n17589_,
    new_n17590_, new_n17591_, new_n17592_, new_n17593_, new_n17594_,
    new_n17595_, new_n17596_, new_n17597_, new_n17598_, new_n17599_,
    new_n17600_, new_n17601_, new_n17602_, new_n17603_, new_n17604_,
    new_n17605_, new_n17606_, new_n17607_, new_n17608_, new_n17609_,
    new_n17610_, new_n17611_, new_n17612_, new_n17613_, new_n17614_,
    new_n17615_, new_n17616_, new_n17617_, new_n17618_, new_n17619_,
    new_n17620_, new_n17621_, new_n17622_, new_n17623_, new_n17624_,
    new_n17625_, new_n17626_, new_n17627_, new_n17628_, new_n17629_,
    new_n17630_, new_n17631_, new_n17632_, new_n17633_, new_n17634_,
    new_n17635_, new_n17636_, new_n17637_, new_n17638_, new_n17639_,
    new_n17640_, new_n17641_, new_n17642_, new_n17643_, new_n17644_,
    new_n17645_, new_n17646_, new_n17647_, new_n17648_, new_n17649_,
    new_n17650_, new_n17651_, new_n17652_, new_n17653_, new_n17654_,
    new_n17655_, new_n17656_, new_n17657_, new_n17658_, new_n17659_,
    new_n17660_, new_n17661_, new_n17662_, new_n17663_, new_n17664_,
    new_n17665_, new_n17666_, new_n17667_, new_n17668_, new_n17669_,
    new_n17670_, new_n17671_, new_n17672_, new_n17673_, new_n17674_,
    new_n17675_, new_n17676_, new_n17677_, new_n17678_, new_n17679_,
    new_n17680_, new_n17681_, new_n17682_, new_n17683_, new_n17684_,
    new_n17685_, new_n17686_, new_n17687_, new_n17688_, new_n17689_,
    new_n17690_, new_n17691_, new_n17692_, new_n17693_, new_n17694_,
    new_n17695_, new_n17696_, new_n17697_, new_n17698_, new_n17699_,
    new_n17700_, new_n17701_, new_n17702_, new_n17703_, new_n17704_,
    new_n17705_, new_n17706_, new_n17707_, new_n17708_, new_n17709_,
    new_n17710_, new_n17711_, new_n17712_, new_n17713_, new_n17714_,
    new_n17715_, new_n17716_, new_n17717_, new_n17718_, new_n17719_,
    new_n17720_, new_n17721_, new_n17722_, new_n17723_, new_n17724_,
    new_n17725_, new_n17726_, new_n17727_, new_n17728_, new_n17729_,
    new_n17730_, new_n17731_, new_n17732_, new_n17733_, new_n17734_,
    new_n17735_, new_n17736_, new_n17737_, new_n17738_, new_n17739_,
    new_n17740_, new_n17741_, new_n17742_, new_n17743_, new_n17744_,
    new_n17745_, new_n17746_, new_n17747_, new_n17748_, new_n17749_,
    new_n17750_, new_n17751_, new_n17752_, new_n17753_, new_n17754_,
    new_n17755_, new_n17756_, new_n17757_, new_n17758_, new_n17759_,
    new_n17760_, new_n17761_, new_n17762_, new_n17763_, new_n17764_,
    new_n17765_, new_n17766_, new_n17767_, new_n17768_, new_n17769_,
    new_n17770_, new_n17771_, new_n17772_, new_n17773_, new_n17774_,
    new_n17775_, new_n17776_, new_n17777_, new_n17778_, new_n17779_,
    new_n17780_, new_n17781_, new_n17782_, new_n17783_, new_n17784_,
    new_n17785_, new_n17786_, new_n17787_, new_n17788_, new_n17789_,
    new_n17790_, new_n17791_, new_n17792_, new_n17793_, new_n17794_,
    new_n17795_, new_n17796_, new_n17797_, new_n17798_, new_n17799_,
    new_n17800_, new_n17801_, new_n17802_, new_n17803_, new_n17804_,
    new_n17805_, new_n17806_, new_n17807_, new_n17808_, new_n17809_,
    new_n17810_, new_n17811_, new_n17812_, new_n17813_, new_n17814_,
    new_n17815_, new_n17816_, new_n17817_, new_n17818_, new_n17819_,
    new_n17820_, new_n17821_, new_n17822_, new_n17823_, new_n17824_,
    new_n17825_, new_n17826_, new_n17827_, new_n17828_, new_n17829_,
    new_n17830_, new_n17831_, new_n17832_, new_n17833_, new_n17834_,
    new_n17835_, new_n17836_, new_n17837_, new_n17838_, new_n17839_,
    new_n17840_, new_n17841_, new_n17843_, new_n17844_, new_n17845_,
    new_n17846_, new_n17847_, new_n17848_, new_n17849_, new_n17850_,
    new_n17851_, new_n17852_, new_n17853_, new_n17854_, new_n17855_,
    new_n17856_, new_n17857_, new_n17858_, new_n17859_, new_n17860_,
    new_n17861_, new_n17862_, new_n17863_, new_n17864_, new_n17865_,
    new_n17866_, new_n17867_, new_n17868_, new_n17869_, new_n17870_,
    new_n17871_, new_n17872_, new_n17873_, new_n17874_, new_n17875_,
    new_n17876_, new_n17877_, new_n17878_, new_n17879_, new_n17880_,
    new_n17881_, new_n17882_, new_n17883_, new_n17884_, new_n17885_,
    new_n17886_, new_n17887_, new_n17888_, new_n17889_, new_n17890_,
    new_n17891_, new_n17892_, new_n17893_, new_n17894_, new_n17895_,
    new_n17896_, new_n17897_, new_n17898_, new_n17899_, new_n17900_,
    new_n17901_, new_n17902_, new_n17903_, new_n17904_, new_n17905_,
    new_n17906_, new_n17907_, new_n17908_, new_n17909_, new_n17910_,
    new_n17911_, new_n17912_, new_n17913_, new_n17914_, new_n17915_,
    new_n17916_, new_n17917_, new_n17918_, new_n17919_, new_n17920_,
    new_n17921_, new_n17922_, new_n17923_, new_n17924_, new_n17925_,
    new_n17926_, new_n17927_, new_n17928_, new_n17929_, new_n17930_,
    new_n17931_, new_n17932_, new_n17933_, new_n17934_, new_n17935_,
    new_n17936_, new_n17937_, new_n17938_, new_n17939_, new_n17940_,
    new_n17941_, new_n17942_, new_n17943_, new_n17944_, new_n17945_,
    new_n17946_, new_n17947_, new_n17948_, new_n17949_, new_n17950_,
    new_n17951_, new_n17952_, new_n17953_, new_n17954_, new_n17955_,
    new_n17956_, new_n17957_, new_n17958_, new_n17959_, new_n17960_,
    new_n17961_, new_n17962_, new_n17963_, new_n17964_, new_n17965_,
    new_n17966_, new_n17967_, new_n17968_, new_n17969_, new_n17970_,
    new_n17971_, new_n17972_, new_n17973_, new_n17974_, new_n17975_,
    new_n17976_, new_n17977_, new_n17978_, new_n17979_, new_n17980_,
    new_n17981_, new_n17982_, new_n17983_, new_n17984_, new_n17985_,
    new_n17986_, new_n17987_, new_n17988_, new_n17989_, new_n17990_,
    new_n17991_, new_n17992_, new_n17993_, new_n17994_, new_n17995_,
    new_n17996_, new_n17997_, new_n17998_, new_n17999_, new_n18000_,
    new_n18001_, new_n18002_, new_n18003_, new_n18004_, new_n18005_,
    new_n18006_, new_n18007_, new_n18008_, new_n18009_, new_n18010_,
    new_n18011_, new_n18012_, new_n18013_, new_n18014_, new_n18015_,
    new_n18016_, new_n18017_, new_n18018_, new_n18019_, new_n18020_,
    new_n18021_, new_n18022_, new_n18023_, new_n18024_, new_n18025_,
    new_n18026_, new_n18027_, new_n18028_, new_n18029_, new_n18030_,
    new_n18031_, new_n18032_, new_n18033_, new_n18034_, new_n18035_,
    new_n18036_, new_n18037_, new_n18038_, new_n18039_, new_n18040_,
    new_n18041_, new_n18042_, new_n18043_, new_n18044_, new_n18045_,
    new_n18046_, new_n18047_, new_n18048_, new_n18049_, new_n18050_,
    new_n18051_, new_n18052_, new_n18053_, new_n18054_, new_n18055_,
    new_n18056_, new_n18057_, new_n18058_, new_n18059_, new_n18060_,
    new_n18061_, new_n18062_, new_n18063_, new_n18064_, new_n18065_,
    new_n18066_, new_n18067_, new_n18068_, new_n18069_, new_n18070_,
    new_n18071_, new_n18072_, new_n18073_, new_n18074_, new_n18075_,
    new_n18076_, new_n18077_, new_n18078_, new_n18079_, new_n18080_,
    new_n18081_, new_n18082_, new_n18083_, new_n18084_, new_n18085_,
    new_n18086_, new_n18087_, new_n18088_, new_n18089_, new_n18090_,
    new_n18091_, new_n18092_, new_n18093_, new_n18094_, new_n18095_,
    new_n18096_, new_n18097_, new_n18098_, new_n18099_, new_n18100_,
    new_n18101_, new_n18102_, new_n18103_, new_n18104_, new_n18105_,
    new_n18106_, new_n18107_, new_n18108_, new_n18109_, new_n18110_,
    new_n18111_, new_n18112_, new_n18113_, new_n18114_, new_n18115_,
    new_n18116_, new_n18117_, new_n18118_, new_n18119_, new_n18120_,
    new_n18121_, new_n18122_, new_n18123_, new_n18124_, new_n18125_,
    new_n18126_, new_n18127_, new_n18128_, new_n18129_, new_n18130_,
    new_n18131_, new_n18132_, new_n18133_, new_n18134_, new_n18135_,
    new_n18136_, new_n18137_, new_n18138_, new_n18139_, new_n18140_,
    new_n18141_, new_n18142_, new_n18143_, new_n18144_, new_n18145_,
    new_n18146_, new_n18147_, new_n18148_, new_n18149_, new_n18150_,
    new_n18151_, new_n18152_, new_n18153_, new_n18154_, new_n18155_,
    new_n18156_, new_n18157_, new_n18158_, new_n18159_, new_n18160_,
    new_n18161_, new_n18162_, new_n18163_, new_n18164_, new_n18165_,
    new_n18166_, new_n18167_, new_n18168_, new_n18169_, new_n18170_,
    new_n18171_, new_n18172_, new_n18173_, new_n18174_, new_n18176_,
    new_n18177_, new_n18178_, new_n18179_, new_n18180_, new_n18181_,
    new_n18182_, new_n18183_, new_n18184_, new_n18185_, new_n18186_,
    new_n18187_, new_n18188_, new_n18189_, new_n18190_, new_n18191_,
    new_n18192_, new_n18193_, new_n18194_, new_n18195_, new_n18196_,
    new_n18197_, new_n18198_, new_n18199_, new_n18200_, new_n18201_,
    new_n18202_, new_n18203_, new_n18204_, new_n18205_, new_n18206_,
    new_n18207_, new_n18208_, new_n18209_, new_n18210_, new_n18211_,
    new_n18212_, new_n18213_, new_n18214_, new_n18215_, new_n18216_,
    new_n18217_, new_n18218_, new_n18219_, new_n18220_, new_n18221_,
    new_n18222_, new_n18223_, new_n18224_, new_n18225_, new_n18226_,
    new_n18227_, new_n18228_, new_n18229_, new_n18230_, new_n18231_,
    new_n18232_, new_n18233_, new_n18234_, new_n18235_, new_n18236_,
    new_n18237_, new_n18238_, new_n18239_, new_n18240_, new_n18241_,
    new_n18242_, new_n18243_, new_n18244_, new_n18245_, new_n18246_,
    new_n18247_, new_n18248_, new_n18249_, new_n18250_, new_n18251_,
    new_n18252_, new_n18253_, new_n18254_, new_n18255_, new_n18256_,
    new_n18257_, new_n18258_, new_n18259_, new_n18260_, new_n18261_,
    new_n18262_, new_n18263_, new_n18264_, new_n18265_, new_n18266_,
    new_n18267_, new_n18268_, new_n18269_, new_n18270_, new_n18271_,
    new_n18272_, new_n18273_, new_n18274_, new_n18275_, new_n18276_,
    new_n18277_, new_n18278_, new_n18279_, new_n18280_, new_n18281_,
    new_n18282_, new_n18283_, new_n18284_, new_n18285_, new_n18286_,
    new_n18287_, new_n18288_, new_n18289_, new_n18290_, new_n18291_,
    new_n18292_, new_n18293_, new_n18294_, new_n18295_, new_n18296_,
    new_n18297_, new_n18298_, new_n18299_, new_n18300_, new_n18301_,
    new_n18302_, new_n18303_, new_n18304_, new_n18305_, new_n18306_,
    new_n18307_, new_n18308_, new_n18309_, new_n18310_, new_n18311_,
    new_n18312_, new_n18313_, new_n18314_, new_n18315_, new_n18316_,
    new_n18317_, new_n18318_, new_n18319_, new_n18320_, new_n18321_,
    new_n18322_, new_n18323_, new_n18324_, new_n18325_, new_n18326_,
    new_n18327_, new_n18328_, new_n18329_, new_n18330_, new_n18331_,
    new_n18332_, new_n18333_, new_n18334_, new_n18335_, new_n18336_,
    new_n18337_, new_n18338_, new_n18339_, new_n18340_, new_n18341_,
    new_n18342_, new_n18343_, new_n18344_, new_n18345_, new_n18346_,
    new_n18347_, new_n18348_, new_n18349_, new_n18350_, new_n18351_,
    new_n18352_, new_n18353_, new_n18354_, new_n18355_, new_n18356_,
    new_n18357_, new_n18358_, new_n18359_, new_n18360_, new_n18361_,
    new_n18362_, new_n18363_, new_n18364_, new_n18365_, new_n18366_,
    new_n18367_, new_n18368_, new_n18369_, new_n18370_, new_n18371_,
    new_n18372_, new_n18373_, new_n18374_, new_n18375_, new_n18376_,
    new_n18377_, new_n18378_, new_n18379_, new_n18380_, new_n18381_,
    new_n18382_, new_n18383_, new_n18384_, new_n18385_, new_n18386_,
    new_n18387_, new_n18388_, new_n18389_, new_n18390_, new_n18391_,
    new_n18392_, new_n18393_, new_n18394_, new_n18395_, new_n18396_,
    new_n18397_, new_n18398_, new_n18399_, new_n18400_, new_n18401_,
    new_n18402_, new_n18403_, new_n18404_, new_n18405_, new_n18406_,
    new_n18407_, new_n18408_, new_n18409_, new_n18410_, new_n18411_,
    new_n18412_, new_n18413_, new_n18414_, new_n18415_, new_n18416_,
    new_n18417_, new_n18418_, new_n18419_, new_n18420_, new_n18421_,
    new_n18422_, new_n18423_, new_n18424_, new_n18425_, new_n18426_,
    new_n18427_, new_n18428_, new_n18429_, new_n18430_, new_n18431_,
    new_n18432_, new_n18433_, new_n18434_, new_n18435_, new_n18436_,
    new_n18437_, new_n18438_, new_n18439_, new_n18440_, new_n18441_,
    new_n18442_, new_n18443_, new_n18444_, new_n18445_, new_n18446_,
    new_n18447_, new_n18448_, new_n18449_, new_n18450_, new_n18451_,
    new_n18452_, new_n18453_, new_n18454_, new_n18455_, new_n18456_,
    new_n18457_, new_n18458_, new_n18459_, new_n18460_, new_n18461_,
    new_n18462_, new_n18463_, new_n18464_, new_n18465_, new_n18466_,
    new_n18467_, new_n18468_, new_n18469_, new_n18470_, new_n18471_,
    new_n18472_, new_n18473_, new_n18474_, new_n18475_, new_n18476_,
    new_n18477_, new_n18478_, new_n18479_, new_n18480_, new_n18481_,
    new_n18482_, new_n18483_, new_n18484_, new_n18485_, new_n18486_,
    new_n18487_, new_n18488_, new_n18489_, new_n18490_, new_n18491_,
    new_n18492_, new_n18493_, new_n18494_, new_n18495_, new_n18496_,
    new_n18497_, new_n18498_, new_n18499_, new_n18500_, new_n18501_,
    new_n18502_, new_n18503_, new_n18504_, new_n18505_, new_n18506_,
    new_n18507_, new_n18508_, new_n18509_, new_n18510_, new_n18512_,
    new_n18513_, new_n18514_, new_n18515_, new_n18516_, new_n18517_,
    new_n18518_, new_n18519_, new_n18520_, new_n18521_, new_n18522_,
    new_n18523_, new_n18524_, new_n18525_, new_n18526_, new_n18527_,
    new_n18528_, new_n18529_, new_n18530_, new_n18531_, new_n18532_,
    new_n18533_, new_n18534_, new_n18535_, new_n18536_, new_n18537_,
    new_n18538_, new_n18539_, new_n18540_, new_n18541_, new_n18542_,
    new_n18543_, new_n18544_, new_n18545_, new_n18546_, new_n18547_,
    new_n18548_, new_n18549_, new_n18550_, new_n18551_, new_n18552_,
    new_n18553_, new_n18554_, new_n18555_, new_n18556_, new_n18557_,
    new_n18558_, new_n18559_, new_n18560_, new_n18561_, new_n18562_,
    new_n18563_, new_n18564_, new_n18565_, new_n18566_, new_n18567_,
    new_n18568_, new_n18569_, new_n18570_, new_n18571_, new_n18572_,
    new_n18573_, new_n18574_, new_n18575_, new_n18576_, new_n18577_,
    new_n18578_, new_n18579_, new_n18580_, new_n18581_, new_n18582_,
    new_n18583_, new_n18584_, new_n18585_, new_n18586_, new_n18587_,
    new_n18588_, new_n18589_, new_n18590_, new_n18591_, new_n18592_,
    new_n18593_, new_n18594_, new_n18595_, new_n18596_, new_n18597_,
    new_n18598_, new_n18599_, new_n18600_, new_n18601_, new_n18602_,
    new_n18603_, new_n18604_, new_n18605_, new_n18606_, new_n18607_,
    new_n18608_, new_n18609_, new_n18610_, new_n18611_, new_n18612_,
    new_n18613_, new_n18614_, new_n18615_, new_n18616_, new_n18617_,
    new_n18618_, new_n18619_, new_n18620_, new_n18621_, new_n18622_,
    new_n18623_, new_n18624_, new_n18625_, new_n18626_, new_n18627_,
    new_n18628_, new_n18629_, new_n18630_, new_n18631_, new_n18632_,
    new_n18633_, new_n18634_, new_n18635_, new_n18636_, new_n18637_,
    new_n18638_, new_n18639_, new_n18640_, new_n18641_, new_n18642_,
    new_n18643_, new_n18644_, new_n18645_, new_n18646_, new_n18647_,
    new_n18648_, new_n18649_, new_n18650_, new_n18651_, new_n18652_,
    new_n18653_, new_n18654_, new_n18655_, new_n18656_, new_n18657_,
    new_n18658_, new_n18659_, new_n18660_, new_n18661_, new_n18662_,
    new_n18663_, new_n18664_, new_n18665_, new_n18666_, new_n18667_,
    new_n18668_, new_n18669_, new_n18670_, new_n18671_, new_n18672_,
    new_n18673_, new_n18674_, new_n18675_, new_n18676_, new_n18677_,
    new_n18678_, new_n18679_, new_n18680_, new_n18681_, new_n18682_,
    new_n18683_, new_n18684_, new_n18685_, new_n18686_, new_n18687_,
    new_n18688_, new_n18689_, new_n18690_, new_n18691_, new_n18692_,
    new_n18693_, new_n18694_, new_n18695_, new_n18696_, new_n18697_,
    new_n18698_, new_n18699_, new_n18700_, new_n18701_, new_n18702_,
    new_n18703_, new_n18704_, new_n18705_, new_n18706_, new_n18707_,
    new_n18708_, new_n18709_, new_n18710_, new_n18711_, new_n18712_,
    new_n18713_, new_n18714_, new_n18715_, new_n18716_, new_n18717_,
    new_n18718_, new_n18719_, new_n18720_, new_n18721_, new_n18722_,
    new_n18723_, new_n18724_, new_n18725_, new_n18726_, new_n18727_,
    new_n18728_, new_n18729_, new_n18730_, new_n18731_, new_n18732_,
    new_n18733_, new_n18734_, new_n18735_, new_n18736_, new_n18737_,
    new_n18738_, new_n18739_, new_n18740_, new_n18741_, new_n18742_,
    new_n18743_, new_n18744_, new_n18745_, new_n18746_, new_n18747_,
    new_n18748_, new_n18749_, new_n18750_, new_n18751_, new_n18752_,
    new_n18753_, new_n18754_, new_n18755_, new_n18756_, new_n18757_,
    new_n18758_, new_n18759_, new_n18760_, new_n18761_, new_n18762_,
    new_n18763_, new_n18764_, new_n18765_, new_n18766_, new_n18767_,
    new_n18768_, new_n18769_, new_n18770_, new_n18771_, new_n18772_,
    new_n18773_, new_n18774_, new_n18775_, new_n18776_, new_n18777_,
    new_n18778_, new_n18779_, new_n18780_, new_n18781_, new_n18782_,
    new_n18783_, new_n18784_, new_n18785_, new_n18786_, new_n18787_,
    new_n18788_, new_n18789_, new_n18790_, new_n18791_, new_n18792_,
    new_n18793_, new_n18794_, new_n18795_, new_n18796_, new_n18797_,
    new_n18798_, new_n18799_, new_n18800_, new_n18801_, new_n18802_,
    new_n18803_, new_n18804_, new_n18805_, new_n18806_, new_n18807_,
    new_n18808_, new_n18809_, new_n18810_, new_n18811_, new_n18812_,
    new_n18813_, new_n18814_, new_n18815_, new_n18816_, new_n18817_,
    new_n18818_, new_n18819_, new_n18820_, new_n18821_, new_n18822_,
    new_n18823_, new_n18824_, new_n18825_, new_n18826_, new_n18827_,
    new_n18828_, new_n18829_, new_n18830_, new_n18831_, new_n18832_,
    new_n18833_, new_n18834_, new_n18835_, new_n18836_, new_n18837_,
    new_n18838_, new_n18839_, new_n18840_, new_n18841_, new_n18842_,
    new_n18843_, new_n18844_, new_n18845_, new_n18846_, new_n18847_,
    new_n18848_, new_n18849_, new_n18850_, new_n18851_, new_n18852_,
    new_n18853_, new_n18854_, new_n18855_, new_n18856_, new_n18857_,
    new_n18859_, new_n18860_, new_n18861_, new_n18862_, new_n18863_,
    new_n18864_, new_n18865_, new_n18866_, new_n18867_, new_n18868_,
    new_n18869_, new_n18870_, new_n18871_, new_n18872_, new_n18873_,
    new_n18874_, new_n18875_, new_n18876_, new_n18877_, new_n18878_,
    new_n18879_, new_n18880_, new_n18881_, new_n18882_, new_n18883_,
    new_n18884_, new_n18885_, new_n18886_, new_n18887_, new_n18888_,
    new_n18889_, new_n18890_, new_n18891_, new_n18892_, new_n18893_,
    new_n18894_, new_n18895_, new_n18896_, new_n18897_, new_n18898_,
    new_n18899_, new_n18900_, new_n18901_, new_n18902_, new_n18903_,
    new_n18904_, new_n18905_, new_n18906_, new_n18907_, new_n18908_,
    new_n18909_, new_n18910_, new_n18911_, new_n18912_, new_n18913_,
    new_n18914_, new_n18915_, new_n18916_, new_n18917_, new_n18918_,
    new_n18919_, new_n18920_, new_n18921_, new_n18922_, new_n18923_,
    new_n18924_, new_n18925_, new_n18926_, new_n18927_, new_n18928_,
    new_n18929_, new_n18930_, new_n18931_, new_n18932_, new_n18933_,
    new_n18934_, new_n18935_, new_n18936_, new_n18937_, new_n18938_,
    new_n18939_, new_n18940_, new_n18941_, new_n18942_, new_n18943_,
    new_n18944_, new_n18945_, new_n18946_, new_n18947_, new_n18948_,
    new_n18949_, new_n18950_, new_n18951_, new_n18952_, new_n18953_,
    new_n18954_, new_n18955_, new_n18956_, new_n18957_, new_n18958_,
    new_n18959_, new_n18960_, new_n18961_, new_n18962_, new_n18963_,
    new_n18964_, new_n18965_, new_n18966_, new_n18967_, new_n18968_,
    new_n18969_, new_n18970_, new_n18971_, new_n18972_, new_n18973_,
    new_n18974_, new_n18975_, new_n18976_, new_n18977_, new_n18978_,
    new_n18979_, new_n18980_, new_n18981_, new_n18982_, new_n18983_,
    new_n18984_, new_n18985_, new_n18986_, new_n18987_, new_n18988_,
    new_n18989_, new_n18990_, new_n18991_, new_n18992_, new_n18993_,
    new_n18994_, new_n18995_, new_n18996_, new_n18997_, new_n18998_,
    new_n18999_, new_n19000_, new_n19001_, new_n19002_, new_n19003_,
    new_n19004_, new_n19005_, new_n19006_, new_n19007_, new_n19008_,
    new_n19009_, new_n19010_, new_n19011_, new_n19012_, new_n19013_,
    new_n19014_, new_n19015_, new_n19016_, new_n19017_, new_n19018_,
    new_n19019_, new_n19020_, new_n19021_, new_n19022_, new_n19023_,
    new_n19024_, new_n19025_, new_n19026_, new_n19027_, new_n19028_,
    new_n19029_, new_n19030_, new_n19031_, new_n19032_, new_n19033_,
    new_n19034_, new_n19035_, new_n19036_, new_n19037_, new_n19038_,
    new_n19039_, new_n19040_, new_n19041_, new_n19042_, new_n19043_,
    new_n19044_, new_n19045_, new_n19046_, new_n19047_, new_n19048_,
    new_n19049_, new_n19050_, new_n19051_, new_n19052_, new_n19053_,
    new_n19054_, new_n19055_, new_n19056_, new_n19057_, new_n19058_,
    new_n19059_, new_n19060_, new_n19061_, new_n19062_, new_n19063_,
    new_n19064_, new_n19065_, new_n19066_, new_n19067_, new_n19068_,
    new_n19069_, new_n19070_, new_n19071_, new_n19072_, new_n19073_,
    new_n19074_, new_n19075_, new_n19076_, new_n19077_, new_n19078_,
    new_n19079_, new_n19080_, new_n19081_, new_n19082_, new_n19083_,
    new_n19084_, new_n19085_, new_n19086_, new_n19087_, new_n19088_,
    new_n19089_, new_n19090_, new_n19091_, new_n19092_, new_n19093_,
    new_n19094_, new_n19095_, new_n19096_, new_n19097_, new_n19098_,
    new_n19099_, new_n19100_, new_n19101_, new_n19102_, new_n19103_,
    new_n19104_, new_n19105_, new_n19106_, new_n19107_, new_n19108_,
    new_n19109_, new_n19110_, new_n19111_, new_n19112_, new_n19113_,
    new_n19114_, new_n19115_, new_n19116_, new_n19117_, new_n19118_,
    new_n19119_, new_n19120_, new_n19121_, new_n19122_, new_n19123_,
    new_n19124_, new_n19125_, new_n19126_, new_n19127_, new_n19128_,
    new_n19129_, new_n19130_, new_n19131_, new_n19132_, new_n19133_,
    new_n19134_, new_n19135_, new_n19136_, new_n19137_, new_n19138_,
    new_n19139_, new_n19140_, new_n19141_, new_n19142_, new_n19143_,
    new_n19144_, new_n19145_, new_n19146_, new_n19147_, new_n19148_,
    new_n19149_, new_n19150_, new_n19151_, new_n19152_, new_n19153_,
    new_n19154_, new_n19155_, new_n19156_, new_n19157_, new_n19158_,
    new_n19159_, new_n19160_, new_n19161_, new_n19162_, new_n19163_,
    new_n19164_, new_n19165_, new_n19166_, new_n19167_, new_n19168_,
    new_n19169_, new_n19170_, new_n19171_, new_n19172_, new_n19173_,
    new_n19174_, new_n19176_, new_n19177_, new_n19178_, new_n19179_,
    new_n19180_, new_n19181_, new_n19182_, new_n19183_, new_n19184_,
    new_n19185_, new_n19186_, new_n19187_, new_n19188_, new_n19189_,
    new_n19190_, new_n19191_, new_n19192_, new_n19193_, new_n19194_,
    new_n19195_, new_n19196_, new_n19197_, new_n19198_, new_n19199_,
    new_n19200_, new_n19201_, new_n19202_, new_n19203_, new_n19204_,
    new_n19205_, new_n19206_, new_n19207_, new_n19208_, new_n19209_,
    new_n19210_, new_n19211_, new_n19212_, new_n19213_, new_n19214_,
    new_n19215_, new_n19216_, new_n19217_, new_n19218_, new_n19219_,
    new_n19220_, new_n19221_, new_n19222_, new_n19223_, new_n19224_,
    new_n19225_, new_n19226_, new_n19227_, new_n19228_, new_n19229_,
    new_n19230_, new_n19231_, new_n19232_, new_n19233_, new_n19234_,
    new_n19235_, new_n19236_, new_n19237_, new_n19238_, new_n19239_,
    new_n19240_, new_n19241_, new_n19242_, new_n19243_, new_n19244_,
    new_n19245_, new_n19246_, new_n19247_, new_n19248_, new_n19249_,
    new_n19250_, new_n19251_, new_n19252_, new_n19253_, new_n19254_,
    new_n19255_, new_n19256_, new_n19257_, new_n19258_, new_n19259_,
    new_n19260_, new_n19261_, new_n19262_, new_n19263_, new_n19264_,
    new_n19265_, new_n19266_, new_n19267_, new_n19268_, new_n19269_,
    new_n19270_, new_n19271_, new_n19272_, new_n19273_, new_n19274_,
    new_n19275_, new_n19276_, new_n19277_, new_n19278_, new_n19279_,
    new_n19280_, new_n19281_, new_n19282_, new_n19283_, new_n19284_,
    new_n19285_, new_n19286_, new_n19287_, new_n19288_, new_n19289_,
    new_n19290_, new_n19291_, new_n19292_, new_n19293_, new_n19294_,
    new_n19295_, new_n19296_, new_n19297_, new_n19298_, new_n19299_,
    new_n19300_, new_n19301_, new_n19302_, new_n19303_, new_n19304_,
    new_n19305_, new_n19306_, new_n19307_, new_n19308_, new_n19309_,
    new_n19310_, new_n19311_, new_n19312_, new_n19313_, new_n19314_,
    new_n19315_, new_n19316_, new_n19317_, new_n19318_, new_n19319_,
    new_n19320_, new_n19321_, new_n19322_, new_n19323_, new_n19324_,
    new_n19325_, new_n19326_, new_n19327_, new_n19328_, new_n19329_,
    new_n19330_, new_n19331_, new_n19332_, new_n19333_, new_n19334_,
    new_n19335_, new_n19336_, new_n19337_, new_n19338_, new_n19339_,
    new_n19340_, new_n19341_, new_n19342_, new_n19343_, new_n19344_,
    new_n19345_, new_n19346_, new_n19347_, new_n19348_, new_n19349_,
    new_n19350_, new_n19351_, new_n19352_, new_n19353_, new_n19354_,
    new_n19355_, new_n19356_, new_n19357_, new_n19358_, new_n19359_,
    new_n19360_, new_n19361_, new_n19362_, new_n19363_, new_n19364_,
    new_n19365_, new_n19366_, new_n19367_, new_n19368_, new_n19369_,
    new_n19370_, new_n19371_, new_n19372_, new_n19373_, new_n19374_,
    new_n19375_, new_n19376_, new_n19377_, new_n19378_, new_n19379_,
    new_n19380_, new_n19381_, new_n19382_, new_n19383_, new_n19384_,
    new_n19385_, new_n19386_, new_n19387_, new_n19388_, new_n19389_,
    new_n19390_, new_n19391_, new_n19392_, new_n19393_, new_n19394_,
    new_n19395_, new_n19396_, new_n19397_, new_n19398_, new_n19399_,
    new_n19400_, new_n19401_, new_n19402_, new_n19403_, new_n19404_,
    new_n19405_, new_n19406_, new_n19407_, new_n19408_, new_n19409_,
    new_n19410_, new_n19411_, new_n19412_, new_n19413_, new_n19414_,
    new_n19415_, new_n19416_, new_n19417_, new_n19418_, new_n19419_,
    new_n19420_, new_n19421_, new_n19422_, new_n19423_, new_n19424_,
    new_n19425_, new_n19426_, new_n19427_, new_n19428_, new_n19429_,
    new_n19430_, new_n19431_, new_n19432_, new_n19433_, new_n19434_,
    new_n19435_, new_n19436_, new_n19437_, new_n19438_, new_n19439_,
    new_n19440_, new_n19441_, new_n19442_, new_n19443_, new_n19444_,
    new_n19445_, new_n19446_, new_n19447_, new_n19448_, new_n19449_,
    new_n19450_, new_n19451_, new_n19452_, new_n19453_, new_n19454_,
    new_n19455_, new_n19456_, new_n19457_, new_n19458_, new_n19459_,
    new_n19460_, new_n19461_, new_n19462_, new_n19463_, new_n19464_,
    new_n19465_, new_n19466_, new_n19467_, new_n19468_, new_n19469_,
    new_n19470_, new_n19471_, new_n19472_, new_n19473_, new_n19474_,
    new_n19475_, new_n19476_, new_n19477_, new_n19478_, new_n19479_,
    new_n19480_, new_n19481_, new_n19482_, new_n19483_, new_n19484_,
    new_n19485_, new_n19486_, new_n19487_, new_n19488_, new_n19489_,
    new_n19490_, new_n19491_, new_n19492_, new_n19493_, new_n19494_,
    new_n19495_, new_n19496_, new_n19497_, new_n19498_, new_n19499_,
    new_n19500_, new_n19501_, new_n19502_, new_n19503_, new_n19504_,
    new_n19505_, new_n19506_, new_n19507_, new_n19508_, new_n19509_,
    new_n19510_, new_n19511_, new_n19512_, new_n19513_, new_n19515_,
    new_n19516_, new_n19517_, new_n19518_, new_n19519_, new_n19520_,
    new_n19521_, new_n19522_, new_n19523_, new_n19524_, new_n19525_,
    new_n19526_, new_n19527_, new_n19528_, new_n19529_, new_n19530_,
    new_n19531_, new_n19532_, new_n19533_, new_n19534_, new_n19535_,
    new_n19536_, new_n19537_, new_n19538_, new_n19539_, new_n19540_,
    new_n19541_, new_n19542_, new_n19543_, new_n19544_, new_n19545_,
    new_n19546_, new_n19547_, new_n19548_, new_n19549_, new_n19550_,
    new_n19551_, new_n19552_, new_n19553_, new_n19554_, new_n19555_,
    new_n19556_, new_n19557_, new_n19558_, new_n19559_, new_n19560_,
    new_n19561_, new_n19562_, new_n19563_, new_n19564_, new_n19565_,
    new_n19566_, new_n19567_, new_n19568_, new_n19569_, new_n19570_,
    new_n19571_, new_n19572_, new_n19573_, new_n19574_, new_n19575_,
    new_n19576_, new_n19577_, new_n19578_, new_n19579_, new_n19580_,
    new_n19581_, new_n19582_, new_n19583_, new_n19584_, new_n19585_,
    new_n19586_, new_n19587_, new_n19588_, new_n19589_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19639_, new_n19640_,
    new_n19641_, new_n19642_, new_n19643_, new_n19644_, new_n19645_,
    new_n19646_, new_n19647_, new_n19648_, new_n19649_, new_n19650_,
    new_n19651_, new_n19652_, new_n19653_, new_n19654_, new_n19655_,
    new_n19656_, new_n19657_, new_n19658_, new_n19659_, new_n19660_,
    new_n19661_, new_n19662_, new_n19663_, new_n19664_, new_n19665_,
    new_n19666_, new_n19667_, new_n19668_, new_n19669_, new_n19670_,
    new_n19671_, new_n19672_, new_n19673_, new_n19674_, new_n19675_,
    new_n19676_, new_n19677_, new_n19678_, new_n19679_, new_n19680_,
    new_n19681_, new_n19682_, new_n19683_, new_n19684_, new_n19685_,
    new_n19686_, new_n19687_, new_n19688_, new_n19689_, new_n19690_,
    new_n19691_, new_n19692_, new_n19693_, new_n19694_, new_n19695_,
    new_n19696_, new_n19697_, new_n19698_, new_n19699_, new_n19700_,
    new_n19701_, new_n19702_, new_n19703_, new_n19704_, new_n19705_,
    new_n19706_, new_n19707_, new_n19708_, new_n19709_, new_n19710_,
    new_n19711_, new_n19712_, new_n19713_, new_n19714_, new_n19715_,
    new_n19716_, new_n19717_, new_n19718_, new_n19719_, new_n19720_,
    new_n19721_, new_n19722_, new_n19723_, new_n19724_, new_n19725_,
    new_n19726_, new_n19727_, new_n19728_, new_n19729_, new_n19730_,
    new_n19731_, new_n19732_, new_n19733_, new_n19734_, new_n19735_,
    new_n19736_, new_n19737_, new_n19738_, new_n19739_, new_n19740_,
    new_n19741_, new_n19742_, new_n19743_, new_n19744_, new_n19745_,
    new_n19746_, new_n19747_, new_n19748_, new_n19749_, new_n19750_,
    new_n19751_, new_n19752_, new_n19753_, new_n19754_, new_n19755_,
    new_n19756_, new_n19757_, new_n19758_, new_n19759_, new_n19760_,
    new_n19761_, new_n19762_, new_n19763_, new_n19764_, new_n19765_,
    new_n19766_, new_n19767_, new_n19768_, new_n19769_, new_n19770_,
    new_n19771_, new_n19772_, new_n19773_, new_n19774_, new_n19775_,
    new_n19776_, new_n19777_, new_n19778_, new_n19779_, new_n19780_,
    new_n19781_, new_n19782_, new_n19783_, new_n19784_, new_n19785_,
    new_n19786_, new_n19787_, new_n19788_, new_n19789_, new_n19790_,
    new_n19791_, new_n19792_, new_n19793_, new_n19794_, new_n19795_,
    new_n19796_, new_n19797_, new_n19798_, new_n19799_, new_n19800_,
    new_n19801_, new_n19802_, new_n19803_, new_n19804_, new_n19805_,
    new_n19806_, new_n19807_, new_n19808_, new_n19809_, new_n19810_,
    new_n19811_, new_n19812_, new_n19813_, new_n19814_, new_n19815_,
    new_n19816_, new_n19817_, new_n19818_, new_n19819_, new_n19820_,
    new_n19821_, new_n19822_, new_n19823_, new_n19824_, new_n19825_,
    new_n19826_, new_n19827_, new_n19828_, new_n19829_, new_n19830_,
    new_n19831_, new_n19832_, new_n19833_, new_n19835_, new_n19836_,
    new_n19837_, new_n19838_, new_n19839_, new_n19840_, new_n19841_,
    new_n19842_, new_n19843_, new_n19844_, new_n19845_, new_n19846_,
    new_n19847_, new_n19848_, new_n19849_, new_n19850_, new_n19851_,
    new_n19852_, new_n19853_, new_n19854_, new_n19855_, new_n19856_,
    new_n19857_, new_n19858_, new_n19859_, new_n19860_, new_n19861_,
    new_n19862_, new_n19863_, new_n19864_, new_n19865_, new_n19866_,
    new_n19867_, new_n19868_, new_n19869_, new_n19870_, new_n19871_,
    new_n19872_, new_n19873_, new_n19874_, new_n19875_, new_n19876_,
    new_n19877_, new_n19878_, new_n19879_, new_n19880_, new_n19881_,
    new_n19882_, new_n19883_, new_n19884_, new_n19885_, new_n19886_,
    new_n19887_, new_n19888_, new_n19889_, new_n19890_, new_n19891_,
    new_n19892_, new_n19893_, new_n19894_, new_n19895_, new_n19896_,
    new_n19897_, new_n19898_, new_n19899_, new_n19900_, new_n19901_,
    new_n19902_, new_n19903_, new_n19904_, new_n19905_, new_n19906_,
    new_n19907_, new_n19908_, new_n19909_, new_n19910_, new_n19911_,
    new_n19912_, new_n19913_, new_n19914_, new_n19915_, new_n19916_,
    new_n19917_, new_n19918_, new_n19919_, new_n19920_, new_n19921_,
    new_n19922_, new_n19923_, new_n19924_, new_n19925_, new_n19926_,
    new_n19927_, new_n19928_, new_n19929_, new_n19930_, new_n19931_,
    new_n19932_, new_n19933_, new_n19934_, new_n19935_, new_n19936_,
    new_n19937_, new_n19938_, new_n19939_, new_n19940_, new_n19941_,
    new_n19942_, new_n19943_, new_n19944_, new_n19945_, new_n19946_,
    new_n19947_, new_n19948_, new_n19949_, new_n19950_, new_n19951_,
    new_n19952_, new_n19953_, new_n19954_, new_n19955_, new_n19956_,
    new_n19957_, new_n19958_, new_n19959_, new_n19960_, new_n19961_,
    new_n19962_, new_n19963_, new_n19964_, new_n19965_, new_n19966_,
    new_n19967_, new_n19968_, new_n19969_, new_n19970_, new_n19971_,
    new_n19972_, new_n19973_, new_n19974_, new_n19975_, new_n19976_,
    new_n19977_, new_n19978_, new_n19979_, new_n19980_, new_n19981_,
    new_n19982_, new_n19983_, new_n19984_, new_n19985_, new_n19986_,
    new_n19987_, new_n19988_, new_n19989_, new_n19990_, new_n19991_,
    new_n19992_, new_n19993_, new_n19994_, new_n19995_, new_n19996_,
    new_n19997_, new_n19998_, new_n19999_, new_n20000_, new_n20001_,
    new_n20002_, new_n20003_, new_n20004_, new_n20005_, new_n20006_,
    new_n20007_, new_n20008_, new_n20009_, new_n20010_, new_n20011_,
    new_n20012_, new_n20013_, new_n20014_, new_n20015_, new_n20016_,
    new_n20017_, new_n20018_, new_n20019_, new_n20020_, new_n20021_,
    new_n20022_, new_n20023_, new_n20024_, new_n20025_, new_n20026_,
    new_n20027_, new_n20028_, new_n20029_, new_n20030_, new_n20031_,
    new_n20032_, new_n20033_, new_n20034_, new_n20035_, new_n20036_,
    new_n20037_, new_n20038_, new_n20039_, new_n20040_, new_n20041_,
    new_n20042_, new_n20043_, new_n20044_, new_n20045_, new_n20046_,
    new_n20047_, new_n20048_, new_n20049_, new_n20050_, new_n20051_,
    new_n20052_, new_n20053_, new_n20054_, new_n20055_, new_n20056_,
    new_n20057_, new_n20058_, new_n20059_, new_n20060_, new_n20061_,
    new_n20062_, new_n20063_, new_n20064_, new_n20065_, new_n20066_,
    new_n20067_, new_n20068_, new_n20069_, new_n20070_, new_n20071_,
    new_n20072_, new_n20073_, new_n20074_, new_n20075_, new_n20076_,
    new_n20077_, new_n20078_, new_n20079_, new_n20080_, new_n20081_,
    new_n20082_, new_n20083_, new_n20084_, new_n20085_, new_n20086_,
    new_n20087_, new_n20088_, new_n20089_, new_n20090_, new_n20091_,
    new_n20092_, new_n20093_, new_n20094_, new_n20095_, new_n20096_,
    new_n20097_, new_n20098_, new_n20099_, new_n20100_, new_n20101_,
    new_n20102_, new_n20103_, new_n20104_, new_n20105_, new_n20106_,
    new_n20107_, new_n20108_, new_n20109_, new_n20110_, new_n20111_,
    new_n20112_, new_n20113_, new_n20114_, new_n20115_, new_n20116_,
    new_n20117_, new_n20118_, new_n20119_, new_n20120_, new_n20121_,
    new_n20122_, new_n20123_, new_n20124_, new_n20125_, new_n20126_,
    new_n20127_, new_n20128_, new_n20129_, new_n20130_, new_n20131_,
    new_n20132_, new_n20133_, new_n20134_, new_n20135_, new_n20136_,
    new_n20137_, new_n20138_, new_n20139_, new_n20140_, new_n20141_,
    new_n20142_, new_n20143_, new_n20144_, new_n20145_, new_n20146_,
    new_n20147_, new_n20148_, new_n20149_, new_n20150_, new_n20151_,
    new_n20152_, new_n20154_, new_n20155_, new_n20156_, new_n20157_,
    new_n20158_, new_n20159_, new_n20160_, new_n20161_, new_n20162_,
    new_n20163_, new_n20164_, new_n20165_, new_n20166_, new_n20167_,
    new_n20168_, new_n20169_, new_n20170_, new_n20171_, new_n20172_,
    new_n20173_, new_n20174_, new_n20175_, new_n20176_, new_n20177_,
    new_n20178_, new_n20179_, new_n20180_, new_n20181_, new_n20182_,
    new_n20183_, new_n20184_, new_n20185_, new_n20186_, new_n20187_,
    new_n20188_, new_n20189_, new_n20190_, new_n20191_, new_n20192_,
    new_n20193_, new_n20194_, new_n20195_, new_n20196_, new_n20197_,
    new_n20198_, new_n20199_, new_n20200_, new_n20201_, new_n20202_,
    new_n20203_, new_n20204_, new_n20205_, new_n20206_, new_n20207_,
    new_n20208_, new_n20209_, new_n20210_, new_n20211_, new_n20212_,
    new_n20213_, new_n20214_, new_n20215_, new_n20216_, new_n20217_,
    new_n20218_, new_n20219_, new_n20220_, new_n20221_, new_n20222_,
    new_n20223_, new_n20224_, new_n20225_, new_n20226_, new_n20227_,
    new_n20228_, new_n20229_, new_n20230_, new_n20231_, new_n20232_,
    new_n20233_, new_n20234_, new_n20235_, new_n20236_, new_n20237_,
    new_n20238_, new_n20239_, new_n20240_, new_n20241_, new_n20242_,
    new_n20243_, new_n20244_, new_n20245_, new_n20246_, new_n20247_,
    new_n20248_, new_n20249_, new_n20250_, new_n20251_, new_n20252_,
    new_n20253_, new_n20254_, new_n20255_, new_n20256_, new_n20257_,
    new_n20258_, new_n20259_, new_n20260_, new_n20261_, new_n20262_,
    new_n20263_, new_n20264_, new_n20265_, new_n20266_, new_n20267_,
    new_n20268_, new_n20269_, new_n20270_, new_n20271_, new_n20272_,
    new_n20273_, new_n20274_, new_n20275_, new_n20276_, new_n20277_,
    new_n20278_, new_n20279_, new_n20280_, new_n20281_, new_n20282_,
    new_n20283_, new_n20284_, new_n20285_, new_n20286_, new_n20287_,
    new_n20288_, new_n20289_, new_n20290_, new_n20291_, new_n20292_,
    new_n20293_, new_n20294_, new_n20295_, new_n20296_, new_n20297_,
    new_n20298_, new_n20299_, new_n20300_, new_n20301_, new_n20302_,
    new_n20303_, new_n20304_, new_n20305_, new_n20306_, new_n20307_,
    new_n20308_, new_n20309_, new_n20310_, new_n20311_, new_n20312_,
    new_n20313_, new_n20314_, new_n20315_, new_n20316_, new_n20317_,
    new_n20318_, new_n20319_, new_n20320_, new_n20321_, new_n20322_,
    new_n20323_, new_n20324_, new_n20325_, new_n20326_, new_n20327_,
    new_n20328_, new_n20329_, new_n20330_, new_n20331_, new_n20332_,
    new_n20333_, new_n20334_, new_n20335_, new_n20336_, new_n20337_,
    new_n20338_, new_n20339_, new_n20340_, new_n20341_, new_n20342_,
    new_n20343_, new_n20344_, new_n20345_, new_n20346_, new_n20347_,
    new_n20348_, new_n20349_, new_n20350_, new_n20351_, new_n20352_,
    new_n20353_, new_n20354_, new_n20355_, new_n20356_, new_n20357_,
    new_n20358_, new_n20359_, new_n20360_, new_n20361_, new_n20362_,
    new_n20363_, new_n20364_, new_n20365_, new_n20366_, new_n20367_,
    new_n20368_, new_n20369_, new_n20370_, new_n20371_, new_n20372_,
    new_n20373_, new_n20374_, new_n20375_, new_n20376_, new_n20377_,
    new_n20378_, new_n20379_, new_n20380_, new_n20381_, new_n20382_,
    new_n20383_, new_n20384_, new_n20385_, new_n20386_, new_n20387_,
    new_n20388_, new_n20389_, new_n20390_, new_n20391_, new_n20392_,
    new_n20393_, new_n20394_, new_n20395_, new_n20396_, new_n20397_,
    new_n20398_, new_n20399_, new_n20400_, new_n20401_, new_n20402_,
    new_n20403_, new_n20404_, new_n20405_, new_n20406_, new_n20407_,
    new_n20408_, new_n20409_, new_n20410_, new_n20411_, new_n20412_,
    new_n20413_, new_n20414_, new_n20415_, new_n20416_, new_n20417_,
    new_n20418_, new_n20419_, new_n20420_, new_n20421_, new_n20422_,
    new_n20423_, new_n20424_, new_n20425_, new_n20426_, new_n20427_,
    new_n20428_, new_n20429_, new_n20430_, new_n20431_, new_n20432_,
    new_n20433_, new_n20434_, new_n20435_, new_n20436_, new_n20437_,
    new_n20438_, new_n20439_, new_n20440_, new_n20441_, new_n20442_,
    new_n20443_, new_n20444_, new_n20445_, new_n20446_, new_n20447_,
    new_n20448_, new_n20449_, new_n20450_, new_n20451_, new_n20452_,
    new_n20453_, new_n20454_, new_n20455_, new_n20456_, new_n20457_,
    new_n20458_, new_n20459_, new_n20460_, new_n20461_, new_n20462_,
    new_n20463_, new_n20464_, new_n20465_, new_n20466_, new_n20467_,
    new_n20468_, new_n20470_, new_n20471_, new_n20472_, new_n20473_,
    new_n20474_, new_n20475_, new_n20476_, new_n20477_, new_n20478_,
    new_n20479_, new_n20480_, new_n20481_, new_n20482_, new_n20483_,
    new_n20484_, new_n20485_, new_n20486_, new_n20487_, new_n20488_,
    new_n20489_, new_n20490_, new_n20491_, new_n20492_, new_n20493_,
    new_n20494_, new_n20495_, new_n20496_, new_n20497_, new_n20498_,
    new_n20499_, new_n20500_, new_n20501_, new_n20502_, new_n20503_,
    new_n20504_, new_n20505_, new_n20506_, new_n20507_, new_n20508_,
    new_n20509_, new_n20510_, new_n20511_, new_n20512_, new_n20513_,
    new_n20514_, new_n20515_, new_n20516_, new_n20517_, new_n20518_,
    new_n20519_, new_n20520_, new_n20521_, new_n20522_, new_n20523_,
    new_n20524_, new_n20525_, new_n20526_, new_n20527_, new_n20528_,
    new_n20529_, new_n20530_, new_n20531_, new_n20532_, new_n20533_,
    new_n20534_, new_n20535_, new_n20536_, new_n20537_, new_n20538_,
    new_n20539_, new_n20540_, new_n20541_, new_n20542_, new_n20543_,
    new_n20544_, new_n20545_, new_n20546_, new_n20547_, new_n20548_,
    new_n20549_, new_n20550_, new_n20551_, new_n20552_, new_n20553_,
    new_n20554_, new_n20555_, new_n20556_, new_n20557_, new_n20558_,
    new_n20559_, new_n20560_, new_n20561_, new_n20562_, new_n20563_,
    new_n20564_, new_n20565_, new_n20566_, new_n20567_, new_n20568_,
    new_n20569_, new_n20570_, new_n20571_, new_n20572_, new_n20573_,
    new_n20574_, new_n20575_, new_n20576_, new_n20577_, new_n20578_,
    new_n20579_, new_n20580_, new_n20581_, new_n20582_, new_n20583_,
    new_n20584_, new_n20585_, new_n20586_, new_n20587_, new_n20588_,
    new_n20589_, new_n20590_, new_n20591_, new_n20592_, new_n20593_,
    new_n20594_, new_n20595_, new_n20596_, new_n20597_, new_n20598_,
    new_n20599_, new_n20600_, new_n20601_, new_n20602_, new_n20603_,
    new_n20604_, new_n20605_, new_n20606_, new_n20607_, new_n20608_,
    new_n20609_, new_n20610_, new_n20611_, new_n20612_, new_n20613_,
    new_n20614_, new_n20615_, new_n20616_, new_n20617_, new_n20618_,
    new_n20619_, new_n20620_, new_n20621_, new_n20622_, new_n20623_,
    new_n20624_, new_n20625_, new_n20626_, new_n20627_, new_n20628_,
    new_n20629_, new_n20630_, new_n20631_, new_n20632_, new_n20633_,
    new_n20634_, new_n20635_, new_n20636_, new_n20637_, new_n20638_,
    new_n20639_, new_n20640_, new_n20641_, new_n20642_, new_n20643_,
    new_n20644_, new_n20645_, new_n20646_, new_n20647_, new_n20648_,
    new_n20649_, new_n20650_, new_n20651_, new_n20652_, new_n20653_,
    new_n20654_, new_n20655_, new_n20656_, new_n20657_, new_n20658_,
    new_n20659_, new_n20660_, new_n20661_, new_n20662_, new_n20663_,
    new_n20664_, new_n20665_, new_n20666_, new_n20667_, new_n20668_,
    new_n20669_, new_n20670_, new_n20671_, new_n20672_, new_n20673_,
    new_n20674_, new_n20675_, new_n20676_, new_n20677_, new_n20678_,
    new_n20679_, new_n20680_, new_n20681_, new_n20682_, new_n20683_,
    new_n20684_, new_n20685_, new_n20686_, new_n20687_, new_n20688_,
    new_n20689_, new_n20690_, new_n20691_, new_n20692_, new_n20693_,
    new_n20694_, new_n20695_, new_n20696_, new_n20697_, new_n20698_,
    new_n20699_, new_n20700_, new_n20701_, new_n20702_, new_n20703_,
    new_n20704_, new_n20705_, new_n20706_, new_n20707_, new_n20708_,
    new_n20709_, new_n20710_, new_n20711_, new_n20712_, new_n20713_,
    new_n20714_, new_n20715_, new_n20716_, new_n20717_, new_n20718_,
    new_n20719_, new_n20720_, new_n20721_, new_n20722_, new_n20723_,
    new_n20724_, new_n20725_, new_n20726_, new_n20727_, new_n20728_,
    new_n20729_, new_n20730_, new_n20731_, new_n20732_, new_n20733_,
    new_n20734_, new_n20735_, new_n20736_, new_n20737_, new_n20738_,
    new_n20739_, new_n20740_, new_n20741_, new_n20742_, new_n20743_,
    new_n20744_, new_n20745_, new_n20746_, new_n20747_, new_n20748_,
    new_n20749_, new_n20750_, new_n20751_, new_n20752_, new_n20753_,
    new_n20754_, new_n20755_, new_n20756_, new_n20757_, new_n20758_,
    new_n20759_, new_n20760_, new_n20761_, new_n20762_, new_n20763_,
    new_n20764_, new_n20765_, new_n20766_, new_n20767_, new_n20768_,
    new_n20769_, new_n20770_, new_n20771_, new_n20772_, new_n20773_,
    new_n20774_, new_n20775_, new_n20776_, new_n20777_, new_n20778_,
    new_n20779_, new_n20780_, new_n20781_, new_n20782_, new_n20783_,
    new_n20784_, new_n20786_, new_n20787_, new_n20788_, new_n20789_,
    new_n20790_, new_n20791_, new_n20792_, new_n20793_, new_n20794_,
    new_n20795_, new_n20796_, new_n20797_, new_n20798_, new_n20799_,
    new_n20800_, new_n20801_, new_n20802_, new_n20803_, new_n20804_,
    new_n20805_, new_n20806_, new_n20807_, new_n20808_, new_n20809_,
    new_n20810_, new_n20811_, new_n20812_, new_n20813_, new_n20814_,
    new_n20815_, new_n20816_, new_n20817_, new_n20818_, new_n20819_,
    new_n20820_, new_n20821_, new_n20822_, new_n20823_, new_n20824_,
    new_n20825_, new_n20826_, new_n20827_, new_n20828_, new_n20829_,
    new_n20830_, new_n20831_, new_n20832_, new_n20833_, new_n20834_,
    new_n20835_, new_n20836_, new_n20837_, new_n20838_, new_n20839_,
    new_n20840_, new_n20841_, new_n20842_, new_n20843_, new_n20844_,
    new_n20845_, new_n20846_, new_n20847_, new_n20848_, new_n20849_,
    new_n20850_, new_n20851_, new_n20852_, new_n20853_, new_n20854_,
    new_n20855_, new_n20856_, new_n20857_, new_n20858_, new_n20859_,
    new_n20860_, new_n20861_, new_n20862_, new_n20863_, new_n20864_,
    new_n20865_, new_n20866_, new_n20867_, new_n20868_, new_n20869_,
    new_n20870_, new_n20871_, new_n20872_, new_n20873_, new_n20874_,
    new_n20875_, new_n20876_, new_n20877_, new_n20878_, new_n20879_,
    new_n20880_, new_n20881_, new_n20882_, new_n20883_, new_n20884_,
    new_n20885_, new_n20886_, new_n20887_, new_n20888_, new_n20889_,
    new_n20890_, new_n20891_, new_n20892_, new_n20893_, new_n20894_,
    new_n20895_, new_n20896_, new_n20897_, new_n20898_, new_n20899_,
    new_n20900_, new_n20901_, new_n20902_, new_n20903_, new_n20904_,
    new_n20905_, new_n20906_, new_n20907_, new_n20908_, new_n20909_,
    new_n20910_, new_n20911_, new_n20912_, new_n20913_, new_n20914_,
    new_n20915_, new_n20916_, new_n20917_, new_n20918_, new_n20919_,
    new_n20920_, new_n20921_, new_n20922_, new_n20923_, new_n20924_,
    new_n20925_, new_n20926_, new_n20927_, new_n20928_, new_n20929_,
    new_n20930_, new_n20931_, new_n20932_, new_n20933_, new_n20934_,
    new_n20935_, new_n20936_, new_n20937_, new_n20938_, new_n20939_,
    new_n20940_, new_n20941_, new_n20942_, new_n20943_, new_n20944_,
    new_n20945_, new_n20946_, new_n20947_, new_n20948_, new_n20949_,
    new_n20950_, new_n20951_, new_n20952_, new_n20953_, new_n20954_,
    new_n20955_, new_n20956_, new_n20957_, new_n20958_, new_n20959_,
    new_n20960_, new_n20961_, new_n20962_, new_n20963_, new_n20964_,
    new_n20965_, new_n20966_, new_n20967_, new_n20968_, new_n20969_,
    new_n20970_, new_n20971_, new_n20972_, new_n20973_, new_n20974_,
    new_n20975_, new_n20976_, new_n20977_, new_n20978_, new_n20979_,
    new_n20980_, new_n20981_, new_n20982_, new_n20983_, new_n20984_,
    new_n20985_, new_n20986_, new_n20987_, new_n20988_, new_n20989_,
    new_n20990_, new_n20991_, new_n20992_, new_n20993_, new_n20994_,
    new_n20995_, new_n20996_, new_n20997_, new_n20998_, new_n20999_,
    new_n21000_, new_n21001_, new_n21002_, new_n21003_, new_n21004_,
    new_n21005_, new_n21006_, new_n21007_, new_n21008_, new_n21009_,
    new_n21010_, new_n21011_, new_n21012_, new_n21013_, new_n21014_,
    new_n21015_, new_n21016_, new_n21017_, new_n21018_, new_n21019_,
    new_n21020_, new_n21021_, new_n21022_, new_n21023_, new_n21024_,
    new_n21025_, new_n21026_, new_n21027_, new_n21028_, new_n21029_,
    new_n21030_, new_n21031_, new_n21032_, new_n21033_, new_n21034_,
    new_n21035_, new_n21036_, new_n21037_, new_n21038_, new_n21039_,
    new_n21040_, new_n21041_, new_n21042_, new_n21043_, new_n21044_,
    new_n21045_, new_n21046_, new_n21047_, new_n21048_, new_n21049_,
    new_n21050_, new_n21051_, new_n21052_, new_n21053_, new_n21054_,
    new_n21055_, new_n21056_, new_n21057_, new_n21058_, new_n21059_,
    new_n21060_, new_n21061_, new_n21062_, new_n21063_, new_n21064_,
    new_n21065_, new_n21066_, new_n21067_, new_n21068_, new_n21069_,
    new_n21070_, new_n21071_, new_n21072_, new_n21073_, new_n21074_,
    new_n21075_, new_n21076_, new_n21077_, new_n21078_, new_n21079_,
    new_n21080_, new_n21081_, new_n21082_, new_n21083_, new_n21084_,
    new_n21085_, new_n21086_, new_n21087_, new_n21088_, new_n21089_,
    new_n21090_, new_n21091_, new_n21092_, new_n21093_, new_n21094_,
    new_n21095_, new_n21096_, new_n21097_, new_n21098_, new_n21099_,
    new_n21100_, new_n21102_, new_n21103_, new_n21104_, new_n21105_,
    new_n21106_, new_n21107_, new_n21108_, new_n21109_, new_n21110_,
    new_n21111_, new_n21112_, new_n21113_, new_n21114_, new_n21115_,
    new_n21116_, new_n21117_, new_n21118_, new_n21119_, new_n21120_,
    new_n21121_, new_n21122_, new_n21123_, new_n21124_, new_n21125_,
    new_n21126_, new_n21127_, new_n21128_, new_n21129_, new_n21130_,
    new_n21131_, new_n21132_, new_n21133_, new_n21134_, new_n21135_,
    new_n21136_, new_n21137_, new_n21138_, new_n21139_, new_n21140_,
    new_n21141_, new_n21142_, new_n21143_, new_n21144_, new_n21145_,
    new_n21146_, new_n21147_, new_n21148_, new_n21149_, new_n21150_,
    new_n21151_, new_n21152_, new_n21153_, new_n21154_, new_n21155_,
    new_n21156_, new_n21157_, new_n21158_, new_n21159_, new_n21160_,
    new_n21161_, new_n21162_, new_n21163_, new_n21164_, new_n21165_,
    new_n21166_, new_n21167_, new_n21168_, new_n21169_, new_n21170_,
    new_n21171_, new_n21172_, new_n21173_, new_n21174_, new_n21175_,
    new_n21176_, new_n21177_, new_n21178_, new_n21179_, new_n21180_,
    new_n21181_, new_n21182_, new_n21183_, new_n21184_, new_n21185_,
    new_n21186_, new_n21187_, new_n21188_, new_n21189_, new_n21190_,
    new_n21191_, new_n21192_, new_n21193_, new_n21194_, new_n21195_,
    new_n21196_, new_n21197_, new_n21198_, new_n21199_, new_n21200_,
    new_n21201_, new_n21202_, new_n21203_, new_n21204_, new_n21205_,
    new_n21206_, new_n21207_, new_n21208_, new_n21209_, new_n21210_,
    new_n21211_, new_n21212_, new_n21213_, new_n21214_, new_n21215_,
    new_n21216_, new_n21217_, new_n21218_, new_n21219_, new_n21220_,
    new_n21221_, new_n21222_, new_n21223_, new_n21224_, new_n21225_,
    new_n21226_, new_n21227_, new_n21228_, new_n21229_, new_n21230_,
    new_n21231_, new_n21232_, new_n21233_, new_n21234_, new_n21235_,
    new_n21236_, new_n21237_, new_n21238_, new_n21239_, new_n21240_,
    new_n21241_, new_n21242_, new_n21243_, new_n21244_, new_n21245_,
    new_n21246_, new_n21247_, new_n21248_, new_n21249_, new_n21250_,
    new_n21251_, new_n21252_, new_n21253_, new_n21254_, new_n21255_,
    new_n21256_, new_n21257_, new_n21258_, new_n21259_, new_n21260_,
    new_n21261_, new_n21262_, new_n21263_, new_n21264_, new_n21265_,
    new_n21266_, new_n21267_, new_n21268_, new_n21269_, new_n21270_,
    new_n21271_, new_n21272_, new_n21273_, new_n21274_, new_n21275_,
    new_n21276_, new_n21277_, new_n21278_, new_n21279_, new_n21280_,
    new_n21281_, new_n21282_, new_n21283_, new_n21284_, new_n21285_,
    new_n21286_, new_n21287_, new_n21288_, new_n21289_, new_n21290_,
    new_n21291_, new_n21292_, new_n21293_, new_n21294_, new_n21295_,
    new_n21296_, new_n21297_, new_n21298_, new_n21299_, new_n21300_,
    new_n21301_, new_n21302_, new_n21303_, new_n21304_, new_n21305_,
    new_n21306_, new_n21307_, new_n21308_, new_n21309_, new_n21310_,
    new_n21311_, new_n21312_, new_n21313_, new_n21314_, new_n21315_,
    new_n21316_, new_n21317_, new_n21318_, new_n21319_, new_n21320_,
    new_n21321_, new_n21322_, new_n21323_, new_n21324_, new_n21325_,
    new_n21326_, new_n21327_, new_n21328_, new_n21329_, new_n21330_,
    new_n21331_, new_n21332_, new_n21333_, new_n21334_, new_n21335_,
    new_n21336_, new_n21337_, new_n21338_, new_n21339_, new_n21340_,
    new_n21341_, new_n21342_, new_n21343_, new_n21344_, new_n21345_,
    new_n21346_, new_n21347_, new_n21348_, new_n21349_, new_n21350_,
    new_n21351_, new_n21352_, new_n21353_, new_n21354_, new_n21355_,
    new_n21356_, new_n21357_, new_n21358_, new_n21359_, new_n21360_,
    new_n21361_, new_n21362_, new_n21363_, new_n21364_, new_n21365_,
    new_n21366_, new_n21367_, new_n21368_, new_n21369_, new_n21370_,
    new_n21371_, new_n21372_, new_n21373_, new_n21374_, new_n21375_,
    new_n21376_, new_n21377_, new_n21378_, new_n21379_, new_n21380_,
    new_n21381_, new_n21382_, new_n21383_, new_n21384_, new_n21385_,
    new_n21386_, new_n21387_, new_n21388_, new_n21389_, new_n21390_,
    new_n21391_, new_n21392_, new_n21393_, new_n21394_, new_n21395_,
    new_n21396_, new_n21397_, new_n21398_, new_n21399_, new_n21400_,
    new_n21401_, new_n21402_, new_n21403_, new_n21404_, new_n21405_,
    new_n21406_, new_n21407_, new_n21408_, new_n21409_, new_n21410_,
    new_n21411_, new_n21412_, new_n21413_, new_n21414_, new_n21415_,
    new_n21416_, new_n21417_, new_n21418_, new_n21419_, new_n21421_,
    new_n21422_, new_n21423_, new_n21424_, new_n21425_, new_n21426_,
    new_n21427_, new_n21428_, new_n21429_, new_n21430_, new_n21431_,
    new_n21432_, new_n21433_, new_n21434_, new_n21435_, new_n21436_,
    new_n21437_, new_n21438_, new_n21439_, new_n21440_, new_n21441_,
    new_n21442_, new_n21443_, new_n21444_, new_n21445_, new_n21446_,
    new_n21447_, new_n21448_, new_n21449_, new_n21450_, new_n21451_,
    new_n21452_, new_n21453_, new_n21454_, new_n21455_, new_n21456_,
    new_n21457_, new_n21458_, new_n21459_, new_n21460_, new_n21461_,
    new_n21462_, new_n21463_, new_n21464_, new_n21465_, new_n21466_,
    new_n21467_, new_n21468_, new_n21469_, new_n21470_, new_n21471_,
    new_n21472_, new_n21473_, new_n21474_, new_n21475_, new_n21476_,
    new_n21477_, new_n21478_, new_n21479_, new_n21480_, new_n21481_,
    new_n21482_, new_n21483_, new_n21484_, new_n21485_, new_n21486_,
    new_n21487_, new_n21488_, new_n21489_, new_n21490_, new_n21491_,
    new_n21492_, new_n21493_, new_n21494_, new_n21495_, new_n21496_,
    new_n21497_, new_n21498_, new_n21499_, new_n21500_, new_n21501_,
    new_n21502_, new_n21503_, new_n21504_, new_n21505_, new_n21506_,
    new_n21507_, new_n21508_, new_n21509_, new_n21510_, new_n21511_,
    new_n21512_, new_n21513_, new_n21514_, new_n21515_, new_n21516_,
    new_n21517_, new_n21518_, new_n21519_, new_n21520_, new_n21521_,
    new_n21522_, new_n21523_, new_n21524_, new_n21525_, new_n21526_,
    new_n21527_, new_n21528_, new_n21529_, new_n21530_, new_n21531_,
    new_n21532_, new_n21533_, new_n21534_, new_n21535_, new_n21536_,
    new_n21537_, new_n21538_, new_n21539_, new_n21540_, new_n21541_,
    new_n21542_, new_n21543_, new_n21544_, new_n21545_, new_n21546_,
    new_n21547_, new_n21548_, new_n21549_, new_n21550_, new_n21551_,
    new_n21552_, new_n21553_, new_n21554_, new_n21555_, new_n21556_,
    new_n21557_, new_n21558_, new_n21559_, new_n21560_, new_n21561_,
    new_n21562_, new_n21563_, new_n21564_, new_n21565_, new_n21566_,
    new_n21567_, new_n21568_, new_n21569_, new_n21570_, new_n21571_,
    new_n21572_, new_n21573_, new_n21574_, new_n21575_, new_n21576_,
    new_n21577_, new_n21578_, new_n21579_, new_n21580_, new_n21581_,
    new_n21582_, new_n21583_, new_n21584_, new_n21585_, new_n21586_,
    new_n21587_, new_n21588_, new_n21589_, new_n21590_, new_n21591_,
    new_n21592_, new_n21593_, new_n21594_, new_n21595_, new_n21596_,
    new_n21597_, new_n21598_, new_n21599_, new_n21600_, new_n21601_,
    new_n21602_, new_n21603_, new_n21604_, new_n21605_, new_n21606_,
    new_n21607_, new_n21608_, new_n21609_, new_n21610_, new_n21611_,
    new_n21612_, new_n21613_, new_n21614_, new_n21615_, new_n21616_,
    new_n21617_, new_n21618_, new_n21619_, new_n21620_, new_n21621_,
    new_n21622_, new_n21623_, new_n21624_, new_n21625_, new_n21626_,
    new_n21627_, new_n21628_, new_n21629_, new_n21630_, new_n21631_,
    new_n21632_, new_n21633_, new_n21634_, new_n21635_, new_n21636_,
    new_n21637_, new_n21638_, new_n21639_, new_n21640_, new_n21641_,
    new_n21642_, new_n21643_, new_n21644_, new_n21645_, new_n21646_,
    new_n21647_, new_n21648_, new_n21649_, new_n21650_, new_n21651_,
    new_n21652_, new_n21653_, new_n21654_, new_n21655_, new_n21656_,
    new_n21657_, new_n21658_, new_n21659_, new_n21660_, new_n21661_,
    new_n21662_, new_n21663_, new_n21664_, new_n21665_, new_n21666_,
    new_n21667_, new_n21668_, new_n21669_, new_n21670_, new_n21671_,
    new_n21672_, new_n21673_, new_n21674_, new_n21675_, new_n21676_,
    new_n21677_, new_n21678_, new_n21679_, new_n21680_, new_n21681_,
    new_n21682_, new_n21683_, new_n21684_, new_n21685_, new_n21686_,
    new_n21687_, new_n21688_, new_n21689_, new_n21690_, new_n21691_,
    new_n21692_, new_n21693_, new_n21694_, new_n21695_, new_n21696_,
    new_n21697_, new_n21698_, new_n21699_, new_n21700_, new_n21701_,
    new_n21702_, new_n21703_, new_n21704_, new_n21705_, new_n21706_,
    new_n21707_, new_n21708_, new_n21709_, new_n21710_, new_n21711_,
    new_n21712_, new_n21713_, new_n21714_, new_n21715_, new_n21716_,
    new_n21717_, new_n21718_, new_n21719_, new_n21720_, new_n21721_,
    new_n21722_, new_n21723_, new_n21724_, new_n21725_, new_n21726_,
    new_n21727_, new_n21728_, new_n21729_, new_n21730_, new_n21731_,
    new_n21732_, new_n21733_, new_n21734_, new_n21735_, new_n21736_,
    new_n21737_, new_n21738_, new_n21739_, new_n21740_, new_n21741_,
    new_n21742_, new_n21743_, new_n21744_, new_n21745_, new_n21746_,
    new_n21747_, new_n21748_, new_n21750_, new_n21751_, new_n21752_,
    new_n21753_, new_n21754_, new_n21755_, new_n21756_, new_n21757_,
    new_n21758_, new_n21759_, new_n21760_, new_n21761_, new_n21762_,
    new_n21763_, new_n21764_, new_n21765_, new_n21766_, new_n21767_,
    new_n21768_, new_n21769_, new_n21770_, new_n21771_, new_n21772_,
    new_n21773_, new_n21774_, new_n21775_, new_n21776_, new_n21777_,
    new_n21778_, new_n21779_, new_n21780_, new_n21781_, new_n21782_,
    new_n21783_, new_n21784_, new_n21785_, new_n21786_, new_n21787_,
    new_n21788_, new_n21789_, new_n21790_, new_n21791_, new_n21792_,
    new_n21793_, new_n21794_, new_n21795_, new_n21796_, new_n21797_,
    new_n21798_, new_n21799_, new_n21800_, new_n21801_, new_n21802_,
    new_n21803_, new_n21804_, new_n21805_, new_n21806_, new_n21807_,
    new_n21808_, new_n21809_, new_n21810_, new_n21811_, new_n21812_,
    new_n21813_, new_n21814_, new_n21815_, new_n21816_, new_n21817_,
    new_n21818_, new_n21819_, new_n21820_, new_n21821_, new_n21822_,
    new_n21823_, new_n21824_, new_n21825_, new_n21826_, new_n21827_,
    new_n21828_, new_n21829_, new_n21830_, new_n21831_, new_n21832_,
    new_n21833_, new_n21834_, new_n21835_, new_n21836_, new_n21837_,
    new_n21838_, new_n21839_, new_n21840_, new_n21841_, new_n21842_,
    new_n21843_, new_n21844_, new_n21845_, new_n21846_, new_n21847_,
    new_n21848_, new_n21849_, new_n21850_, new_n21851_, new_n21852_,
    new_n21853_, new_n21854_, new_n21855_, new_n21856_, new_n21857_,
    new_n21858_, new_n21859_, new_n21860_, new_n21861_, new_n21862_,
    new_n21863_, new_n21864_, new_n21865_, new_n21866_, new_n21867_,
    new_n21868_, new_n21869_, new_n21870_, new_n21871_, new_n21872_,
    new_n21873_, new_n21874_, new_n21875_, new_n21876_, new_n21877_,
    new_n21878_, new_n21879_, new_n21880_, new_n21881_, new_n21882_,
    new_n21883_, new_n21884_, new_n21885_, new_n21886_, new_n21887_,
    new_n21888_, new_n21889_, new_n21890_, new_n21891_, new_n21892_,
    new_n21893_, new_n21894_, new_n21895_, new_n21896_, new_n21897_,
    new_n21898_, new_n21899_, new_n21900_, new_n21901_, new_n21902_,
    new_n21903_, new_n21904_, new_n21905_, new_n21906_, new_n21907_,
    new_n21908_, new_n21909_, new_n21910_, new_n21911_, new_n21912_,
    new_n21913_, new_n21914_, new_n21915_, new_n21916_, new_n21917_,
    new_n21918_, new_n21919_, new_n21920_, new_n21921_, new_n21922_,
    new_n21923_, new_n21924_, new_n21925_, new_n21926_, new_n21927_,
    new_n21928_, new_n21929_, new_n21930_, new_n21931_, new_n21932_,
    new_n21933_, new_n21934_, new_n21935_, new_n21936_, new_n21937_,
    new_n21938_, new_n21939_, new_n21940_, new_n21941_, new_n21942_,
    new_n21943_, new_n21944_, new_n21945_, new_n21946_, new_n21947_,
    new_n21948_, new_n21949_, new_n21950_, new_n21951_, new_n21952_,
    new_n21953_, new_n21954_, new_n21955_, new_n21956_, new_n21957_,
    new_n21958_, new_n21959_, new_n21960_, new_n21961_, new_n21962_,
    new_n21963_, new_n21964_, new_n21965_, new_n21966_, new_n21967_,
    new_n21968_, new_n21969_, new_n21970_, new_n21971_, new_n21972_,
    new_n21973_, new_n21974_, new_n21975_, new_n21976_, new_n21977_,
    new_n21978_, new_n21979_, new_n21980_, new_n21981_, new_n21982_,
    new_n21983_, new_n21984_, new_n21985_, new_n21986_, new_n21987_,
    new_n21988_, new_n21989_, new_n21990_, new_n21991_, new_n21992_,
    new_n21993_, new_n21994_, new_n21995_, new_n21996_, new_n21997_,
    new_n21998_, new_n21999_, new_n22000_, new_n22001_, new_n22002_,
    new_n22003_, new_n22004_, new_n22005_, new_n22006_, new_n22007_,
    new_n22008_, new_n22009_, new_n22010_, new_n22011_, new_n22012_,
    new_n22013_, new_n22014_, new_n22015_, new_n22016_, new_n22017_,
    new_n22018_, new_n22019_, new_n22020_, new_n22021_, new_n22022_,
    new_n22023_, new_n22024_, new_n22025_, new_n22026_, new_n22027_,
    new_n22028_, new_n22029_, new_n22030_, new_n22031_, new_n22032_,
    new_n22033_, new_n22034_, new_n22035_, new_n22036_, new_n22037_,
    new_n22038_, new_n22039_, new_n22040_, new_n22041_, new_n22042_,
    new_n22043_, new_n22044_, new_n22045_, new_n22046_, new_n22047_,
    new_n22048_, new_n22049_, new_n22050_, new_n22051_, new_n22052_,
    new_n22053_, new_n22054_, new_n22055_, new_n22056_, new_n22057_,
    new_n22058_, new_n22059_, new_n22060_, new_n22061_, new_n22062_,
    new_n22063_, new_n22064_, new_n22065_, new_n22066_, new_n22067_,
    new_n22068_, new_n22069_, new_n22070_, new_n22071_, new_n22072_,
    new_n22073_, new_n22074_, new_n22075_, new_n22077_, new_n22078_,
    new_n22079_, new_n22080_, new_n22081_, new_n22082_, new_n22083_,
    new_n22084_, new_n22085_, new_n22086_, new_n22087_, new_n22088_,
    new_n22089_, new_n22090_, new_n22091_, new_n22092_, new_n22093_,
    new_n22094_, new_n22095_, new_n22096_, new_n22097_, new_n22098_,
    new_n22099_, new_n22100_, new_n22101_, new_n22102_, new_n22103_,
    new_n22104_, new_n22105_, new_n22106_, new_n22107_, new_n22108_,
    new_n22109_, new_n22110_, new_n22111_, new_n22112_, new_n22113_,
    new_n22114_, new_n22115_, new_n22116_, new_n22117_, new_n22118_,
    new_n22119_, new_n22120_, new_n22121_, new_n22122_, new_n22123_,
    new_n22124_, new_n22125_, new_n22126_, new_n22127_, new_n22128_,
    new_n22129_, new_n22130_, new_n22131_, new_n22132_, new_n22133_,
    new_n22134_, new_n22135_, new_n22136_, new_n22137_, new_n22138_,
    new_n22139_, new_n22140_, new_n22141_, new_n22142_, new_n22143_,
    new_n22144_, new_n22145_, new_n22146_, new_n22147_, new_n22148_,
    new_n22149_, new_n22150_, new_n22151_, new_n22152_, new_n22153_,
    new_n22154_, new_n22155_, new_n22156_, new_n22157_, new_n22158_,
    new_n22159_, new_n22160_, new_n22161_, new_n22162_, new_n22163_,
    new_n22164_, new_n22165_, new_n22166_, new_n22167_, new_n22168_,
    new_n22169_, new_n22170_, new_n22171_, new_n22172_, new_n22173_,
    new_n22174_, new_n22175_, new_n22176_, new_n22177_, new_n22178_,
    new_n22179_, new_n22180_, new_n22181_, new_n22182_, new_n22183_,
    new_n22184_, new_n22185_, new_n22186_, new_n22187_, new_n22188_,
    new_n22189_, new_n22190_, new_n22191_, new_n22192_, new_n22193_,
    new_n22194_, new_n22195_, new_n22196_, new_n22197_, new_n22198_,
    new_n22199_, new_n22200_, new_n22201_, new_n22202_, new_n22203_,
    new_n22204_, new_n22205_, new_n22206_, new_n22207_, new_n22208_,
    new_n22209_, new_n22210_, new_n22211_, new_n22212_, new_n22213_,
    new_n22214_, new_n22215_, new_n22216_, new_n22217_, new_n22218_,
    new_n22219_, new_n22220_, new_n22221_, new_n22222_, new_n22223_,
    new_n22224_, new_n22225_, new_n22226_, new_n22227_, new_n22228_,
    new_n22229_, new_n22230_, new_n22231_, new_n22232_, new_n22233_,
    new_n22234_, new_n22235_, new_n22236_, new_n22237_, new_n22238_,
    new_n22239_, new_n22240_, new_n22241_, new_n22242_, new_n22243_,
    new_n22244_, new_n22245_, new_n22246_, new_n22247_, new_n22248_,
    new_n22249_, new_n22250_, new_n22251_, new_n22252_, new_n22253_,
    new_n22254_, new_n22255_, new_n22256_, new_n22257_, new_n22258_,
    new_n22259_, new_n22260_, new_n22261_, new_n22262_, new_n22263_,
    new_n22264_, new_n22265_, new_n22266_, new_n22267_, new_n22268_,
    new_n22269_, new_n22270_, new_n22271_, new_n22272_, new_n22273_,
    new_n22274_, new_n22275_, new_n22276_, new_n22277_, new_n22278_,
    new_n22279_, new_n22280_, new_n22281_, new_n22282_, new_n22283_,
    new_n22284_, new_n22285_, new_n22286_, new_n22287_, new_n22288_,
    new_n22289_, new_n22290_, new_n22291_, new_n22292_, new_n22293_,
    new_n22294_, new_n22295_, new_n22296_, new_n22297_, new_n22298_,
    new_n22299_, new_n22300_, new_n22301_, new_n22302_, new_n22303_,
    new_n22304_, new_n22305_, new_n22306_, new_n22307_, new_n22308_,
    new_n22309_, new_n22310_, new_n22311_, new_n22312_, new_n22313_,
    new_n22314_, new_n22315_, new_n22316_, new_n22317_, new_n22318_,
    new_n22319_, new_n22320_, new_n22321_, new_n22322_, new_n22323_,
    new_n22324_, new_n22325_, new_n22326_, new_n22327_, new_n22328_,
    new_n22329_, new_n22330_, new_n22331_, new_n22332_, new_n22333_,
    new_n22334_, new_n22335_, new_n22336_, new_n22337_, new_n22338_,
    new_n22339_, new_n22340_, new_n22341_, new_n22342_, new_n22343_,
    new_n22344_, new_n22345_, new_n22346_, new_n22347_, new_n22348_,
    new_n22349_, new_n22350_, new_n22351_, new_n22352_, new_n22353_,
    new_n22354_, new_n22355_, new_n22356_, new_n22357_, new_n22358_,
    new_n22359_, new_n22360_, new_n22361_, new_n22362_, new_n22363_,
    new_n22364_, new_n22365_, new_n22366_, new_n22367_, new_n22368_,
    new_n22369_, new_n22370_, new_n22371_, new_n22372_, new_n22373_,
    new_n22374_, new_n22375_, new_n22376_, new_n22377_, new_n22378_,
    new_n22379_, new_n22380_, new_n22381_, new_n22382_, new_n22383_,
    new_n22384_, new_n22385_, new_n22386_, new_n22387_, new_n22388_,
    new_n22389_, new_n22390_, new_n22391_, new_n22392_, new_n22393_,
    new_n22394_, new_n22395_, new_n22396_, new_n22397_, new_n22398_,
    new_n22399_, new_n22400_, new_n22401_, new_n22403_, new_n22404_,
    new_n22405_, new_n22406_, new_n22407_, new_n22408_, new_n22409_,
    new_n22410_, new_n22411_, new_n22412_, new_n22413_, new_n22414_,
    new_n22415_, new_n22416_, new_n22417_, new_n22418_, new_n22419_,
    new_n22420_, new_n22421_, new_n22422_, new_n22423_, new_n22424_,
    new_n22425_, new_n22426_, new_n22427_, new_n22428_, new_n22429_,
    new_n22430_, new_n22431_, new_n22432_, new_n22433_, new_n22434_,
    new_n22435_, new_n22436_, new_n22437_, new_n22438_, new_n22439_,
    new_n22440_, new_n22441_, new_n22442_, new_n22443_, new_n22444_,
    new_n22445_, new_n22446_, new_n22447_, new_n22448_, new_n22449_,
    new_n22450_, new_n22451_, new_n22452_, new_n22453_, new_n22454_,
    new_n22455_, new_n22456_, new_n22457_, new_n22458_, new_n22459_,
    new_n22460_, new_n22461_, new_n22462_, new_n22463_, new_n22464_,
    new_n22465_, new_n22466_, new_n22467_, new_n22468_, new_n22469_,
    new_n22470_, new_n22471_, new_n22472_, new_n22473_, new_n22474_,
    new_n22475_, new_n22476_, new_n22477_, new_n22478_, new_n22479_,
    new_n22480_, new_n22481_, new_n22482_, new_n22483_, new_n22484_,
    new_n22485_, new_n22486_, new_n22487_, new_n22488_, new_n22489_,
    new_n22490_, new_n22491_, new_n22492_, new_n22493_, new_n22494_,
    new_n22495_, new_n22496_, new_n22497_, new_n22498_, new_n22499_,
    new_n22500_, new_n22501_, new_n22502_, new_n22503_, new_n22504_,
    new_n22505_, new_n22506_, new_n22507_, new_n22508_, new_n22509_,
    new_n22510_, new_n22511_, new_n22512_, new_n22513_, new_n22514_,
    new_n22515_, new_n22516_, new_n22517_, new_n22518_, new_n22519_,
    new_n22520_, new_n22521_, new_n22522_, new_n22523_, new_n22524_,
    new_n22525_, new_n22526_, new_n22527_, new_n22528_, new_n22529_,
    new_n22530_, new_n22531_, new_n22532_, new_n22533_, new_n22534_,
    new_n22535_, new_n22536_, new_n22537_, new_n22538_, new_n22539_,
    new_n22540_, new_n22541_, new_n22542_, new_n22543_, new_n22544_,
    new_n22545_, new_n22546_, new_n22547_, new_n22548_, new_n22549_,
    new_n22550_, new_n22551_, new_n22552_, new_n22553_, new_n22554_,
    new_n22555_, new_n22556_, new_n22557_, new_n22558_, new_n22559_,
    new_n22560_, new_n22561_, new_n22562_, new_n22563_, new_n22564_,
    new_n22565_, new_n22566_, new_n22567_, new_n22568_, new_n22569_,
    new_n22570_, new_n22571_, new_n22572_, new_n22573_, new_n22574_,
    new_n22575_, new_n22576_, new_n22577_, new_n22578_, new_n22579_,
    new_n22580_, new_n22581_, new_n22582_, new_n22583_, new_n22584_,
    new_n22585_, new_n22586_, new_n22587_, new_n22588_, new_n22589_,
    new_n22590_, new_n22591_, new_n22592_, new_n22593_, new_n22594_,
    new_n22595_, new_n22596_, new_n22597_, new_n22598_, new_n22599_,
    new_n22600_, new_n22601_, new_n22602_, new_n22603_, new_n22604_,
    new_n22605_, new_n22606_, new_n22607_, new_n22608_, new_n22609_,
    new_n22610_, new_n22611_, new_n22612_, new_n22613_, new_n22614_,
    new_n22615_, new_n22616_, new_n22617_, new_n22618_, new_n22619_,
    new_n22620_, new_n22621_, new_n22622_, new_n22623_, new_n22624_,
    new_n22625_, new_n22626_, new_n22627_, new_n22628_, new_n22629_,
    new_n22630_, new_n22631_, new_n22632_, new_n22633_, new_n22634_,
    new_n22635_, new_n22636_, new_n22637_, new_n22638_, new_n22639_,
    new_n22640_, new_n22641_, new_n22642_, new_n22643_, new_n22644_,
    new_n22645_, new_n22646_, new_n22647_, new_n22648_, new_n22649_,
    new_n22650_, new_n22651_, new_n22652_, new_n22653_, new_n22654_,
    new_n22655_, new_n22656_, new_n22657_, new_n22658_, new_n22659_,
    new_n22660_, new_n22661_, new_n22662_, new_n22663_, new_n22664_,
    new_n22665_, new_n22666_, new_n22667_, new_n22668_, new_n22669_,
    new_n22670_, new_n22671_, new_n22672_, new_n22673_, new_n22674_,
    new_n22675_, new_n22676_, new_n22677_, new_n22678_, new_n22679_,
    new_n22680_, new_n22681_, new_n22682_, new_n22683_, new_n22684_,
    new_n22685_, new_n22686_, new_n22687_, new_n22688_, new_n22689_,
    new_n22690_, new_n22691_, new_n22692_, new_n22693_, new_n22694_,
    new_n22695_, new_n22696_, new_n22697_, new_n22698_, new_n22699_,
    new_n22700_, new_n22701_, new_n22702_, new_n22703_, new_n22704_,
    new_n22705_, new_n22706_, new_n22707_, new_n22708_, new_n22709_,
    new_n22710_, new_n22711_, new_n22712_, new_n22713_, new_n22714_,
    new_n22715_, new_n22716_, new_n22717_, new_n22718_, new_n22719_,
    new_n22720_, new_n22721_, new_n22722_, new_n22723_, new_n22724_,
    new_n22725_, new_n22726_, new_n22727_, new_n22728_, new_n22729_,
    new_n22730_, new_n22731_, new_n22732_, new_n22733_, new_n22735_,
    new_n22736_, new_n22737_, new_n22738_, new_n22739_, new_n22740_,
    new_n22741_, new_n22742_, new_n22743_, new_n22744_, new_n22745_,
    new_n22746_, new_n22747_, new_n22748_, new_n22749_, new_n22750_,
    new_n22751_, new_n22752_, new_n22753_, new_n22754_, new_n22755_,
    new_n22756_, new_n22757_, new_n22758_, new_n22759_, new_n22760_,
    new_n22761_, new_n22762_, new_n22763_, new_n22764_, new_n22765_,
    new_n22766_, new_n22767_, new_n22768_, new_n22769_, new_n22770_,
    new_n22771_, new_n22772_, new_n22773_, new_n22774_, new_n22775_,
    new_n22776_, new_n22777_, new_n22778_, new_n22779_, new_n22780_,
    new_n22781_, new_n22782_, new_n22783_, new_n22784_, new_n22785_,
    new_n22786_, new_n22787_, new_n22788_, new_n22789_, new_n22790_,
    new_n22791_, new_n22792_, new_n22793_, new_n22794_, new_n22795_,
    new_n22796_, new_n22797_, new_n22798_, new_n22799_, new_n22800_,
    new_n22801_, new_n22802_, new_n22803_, new_n22804_, new_n22805_,
    new_n22806_, new_n22807_, new_n22808_, new_n22809_, new_n22810_,
    new_n22811_, new_n22812_, new_n22813_, new_n22814_, new_n22815_,
    new_n22816_, new_n22817_, new_n22818_, new_n22819_, new_n22820_,
    new_n22821_, new_n22822_, new_n22823_, new_n22824_, new_n22825_,
    new_n22826_, new_n22827_, new_n22828_, new_n22829_, new_n22830_,
    new_n22831_, new_n22832_, new_n22833_, new_n22834_, new_n22835_,
    new_n22836_, new_n22837_, new_n22838_, new_n22839_, new_n22840_,
    new_n22841_, new_n22842_, new_n22843_, new_n22844_, new_n22845_,
    new_n22846_, new_n22847_, new_n22848_, new_n22849_, new_n22850_,
    new_n22851_, new_n22852_, new_n22853_, new_n22854_, new_n22855_,
    new_n22856_, new_n22857_, new_n22858_, new_n22859_, new_n22860_,
    new_n22861_, new_n22862_, new_n22863_, new_n22864_, new_n22865_,
    new_n22866_, new_n22867_, new_n22868_, new_n22869_, new_n22870_,
    new_n22871_, new_n22872_, new_n22873_, new_n22874_, new_n22875_,
    new_n22876_, new_n22877_, new_n22878_, new_n22879_, new_n22880_,
    new_n22881_, new_n22882_, new_n22883_, new_n22884_, new_n22885_,
    new_n22886_, new_n22887_, new_n22888_, new_n22889_, new_n22890_,
    new_n22891_, new_n22892_, new_n22893_, new_n22894_, new_n22895_,
    new_n22896_, new_n22897_, new_n22898_, new_n22899_, new_n22900_,
    new_n22901_, new_n22902_, new_n22903_, new_n22904_, new_n22905_,
    new_n22906_, new_n22907_, new_n22908_, new_n22909_, new_n22910_,
    new_n22911_, new_n22912_, new_n22913_, new_n22914_, new_n22915_,
    new_n22916_, new_n22917_, new_n22918_, new_n22919_, new_n22920_,
    new_n22921_, new_n22922_, new_n22923_, new_n22924_, new_n22925_,
    new_n22926_, new_n22927_, new_n22928_, new_n22929_, new_n22930_,
    new_n22931_, new_n22932_, new_n22933_, new_n22934_, new_n22935_,
    new_n22936_, new_n22937_, new_n22938_, new_n22939_, new_n22940_,
    new_n22941_, new_n22942_, new_n22943_, new_n22944_, new_n22945_,
    new_n22946_, new_n22947_, new_n22948_, new_n22949_, new_n22950_,
    new_n22951_, new_n22952_, new_n22953_, new_n22954_, new_n22955_,
    new_n22956_, new_n22957_, new_n22958_, new_n22959_, new_n22960_,
    new_n22961_, new_n22962_, new_n22963_, new_n22964_, new_n22965_,
    new_n22966_, new_n22967_, new_n22968_, new_n22969_, new_n22970_,
    new_n22971_, new_n22972_, new_n22973_, new_n22974_, new_n22975_,
    new_n22976_, new_n22977_, new_n22978_, new_n22979_, new_n22980_,
    new_n22981_, new_n22982_, new_n22983_, new_n22984_, new_n22985_,
    new_n22986_, new_n22987_, new_n22988_, new_n22989_, new_n22990_,
    new_n22991_, new_n22992_, new_n22993_, new_n22994_, new_n22995_,
    new_n22996_, new_n22997_, new_n22998_, new_n22999_, new_n23000_,
    new_n23001_, new_n23002_, new_n23003_, new_n23004_, new_n23005_,
    new_n23006_, new_n23007_, new_n23008_, new_n23009_, new_n23010_,
    new_n23011_, new_n23012_, new_n23013_, new_n23014_, new_n23015_,
    new_n23016_, new_n23017_, new_n23018_, new_n23019_, new_n23020_,
    new_n23021_, new_n23022_, new_n23023_, new_n23024_, new_n23025_,
    new_n23026_, new_n23027_, new_n23028_, new_n23029_, new_n23030_,
    new_n23031_, new_n23032_, new_n23033_, new_n23034_, new_n23035_,
    new_n23036_, new_n23037_, new_n23038_, new_n23039_, new_n23040_,
    new_n23041_, new_n23042_, new_n23043_, new_n23044_, new_n23045_,
    new_n23046_, new_n23047_, new_n23048_, new_n23049_, new_n23050_,
    new_n23051_, new_n23052_, new_n23053_, new_n23054_, new_n23055_,
    new_n23056_, new_n23057_, new_n23058_, new_n23060_, new_n23061_,
    new_n23062_, new_n23063_, new_n23064_, new_n23065_, new_n23066_,
    new_n23067_, new_n23068_, new_n23069_, new_n23070_, new_n23071_,
    new_n23072_, new_n23073_, new_n23074_, new_n23075_, new_n23076_,
    new_n23077_, new_n23078_, new_n23079_, new_n23080_, new_n23081_,
    new_n23082_, new_n23083_, new_n23084_, new_n23085_, new_n23086_,
    new_n23087_, new_n23088_, new_n23089_, new_n23090_, new_n23091_,
    new_n23092_, new_n23093_, new_n23094_, new_n23095_, new_n23096_,
    new_n23097_, new_n23098_, new_n23099_, new_n23100_, new_n23101_,
    new_n23102_, new_n23103_, new_n23104_, new_n23105_, new_n23106_,
    new_n23107_, new_n23108_, new_n23109_, new_n23110_, new_n23111_,
    new_n23112_, new_n23113_, new_n23114_, new_n23115_, new_n23116_,
    new_n23117_, new_n23118_, new_n23119_, new_n23120_, new_n23121_,
    new_n23122_, new_n23123_, new_n23124_, new_n23125_, new_n23126_,
    new_n23127_, new_n23128_, new_n23129_, new_n23130_, new_n23131_,
    new_n23132_, new_n23133_, new_n23134_, new_n23135_, new_n23136_,
    new_n23137_, new_n23138_, new_n23139_, new_n23140_, new_n23141_,
    new_n23142_, new_n23143_, new_n23144_, new_n23145_, new_n23146_,
    new_n23147_, new_n23148_, new_n23149_, new_n23150_, new_n23151_,
    new_n23152_, new_n23153_, new_n23154_, new_n23155_, new_n23156_,
    new_n23157_, new_n23158_, new_n23159_, new_n23160_, new_n23161_,
    new_n23162_, new_n23163_, new_n23164_, new_n23165_, new_n23166_,
    new_n23167_, new_n23168_, new_n23169_, new_n23170_, new_n23171_,
    new_n23172_, new_n23173_, new_n23174_, new_n23175_, new_n23176_,
    new_n23177_, new_n23178_, new_n23179_, new_n23180_, new_n23181_,
    new_n23182_, new_n23183_, new_n23184_, new_n23185_, new_n23186_,
    new_n23187_, new_n23188_, new_n23189_, new_n23190_, new_n23191_,
    new_n23192_, new_n23193_, new_n23194_, new_n23195_, new_n23196_,
    new_n23197_, new_n23198_, new_n23199_, new_n23200_, new_n23201_,
    new_n23202_, new_n23203_, new_n23204_, new_n23205_, new_n23206_,
    new_n23207_, new_n23208_, new_n23209_, new_n23210_, new_n23211_,
    new_n23212_, new_n23213_, new_n23214_, new_n23215_, new_n23216_,
    new_n23217_, new_n23218_, new_n23219_, new_n23220_, new_n23221_,
    new_n23222_, new_n23223_, new_n23224_, new_n23225_, new_n23226_,
    new_n23227_, new_n23228_, new_n23229_, new_n23230_, new_n23231_,
    new_n23232_, new_n23233_, new_n23234_, new_n23235_, new_n23236_,
    new_n23237_, new_n23238_, new_n23239_, new_n23240_, new_n23241_,
    new_n23242_, new_n23243_, new_n23244_, new_n23245_, new_n23246_,
    new_n23247_, new_n23248_, new_n23249_, new_n23250_, new_n23251_,
    new_n23252_, new_n23253_, new_n23254_, new_n23255_, new_n23256_,
    new_n23257_, new_n23258_, new_n23259_, new_n23260_, new_n23261_,
    new_n23262_, new_n23263_, new_n23264_, new_n23265_, new_n23266_,
    new_n23267_, new_n23268_, new_n23269_, new_n23270_, new_n23271_,
    new_n23272_, new_n23273_, new_n23274_, new_n23275_, new_n23276_,
    new_n23277_, new_n23278_, new_n23279_, new_n23280_, new_n23281_,
    new_n23282_, new_n23283_, new_n23284_, new_n23285_, new_n23286_,
    new_n23287_, new_n23288_, new_n23289_, new_n23290_, new_n23291_,
    new_n23292_, new_n23293_, new_n23294_, new_n23295_, new_n23296_,
    new_n23297_, new_n23298_, new_n23299_, new_n23300_, new_n23301_,
    new_n23302_, new_n23303_, new_n23304_, new_n23305_, new_n23306_,
    new_n23307_, new_n23308_, new_n23309_, new_n23310_, new_n23311_,
    new_n23312_, new_n23313_, new_n23314_, new_n23315_, new_n23316_,
    new_n23317_, new_n23318_, new_n23319_, new_n23320_, new_n23321_,
    new_n23322_, new_n23323_, new_n23324_, new_n23325_, new_n23326_,
    new_n23327_, new_n23328_, new_n23329_, new_n23330_, new_n23331_,
    new_n23332_, new_n23333_, new_n23334_, new_n23335_, new_n23336_,
    new_n23337_, new_n23338_, new_n23339_, new_n23340_, new_n23341_,
    new_n23342_, new_n23343_, new_n23344_, new_n23345_, new_n23346_,
    new_n23347_, new_n23348_, new_n23349_, new_n23350_, new_n23351_,
    new_n23352_, new_n23353_, new_n23354_, new_n23355_, new_n23356_,
    new_n23357_, new_n23358_, new_n23359_, new_n23360_, new_n23361_,
    new_n23362_, new_n23363_, new_n23364_, new_n23365_, new_n23366_,
    new_n23367_, new_n23368_, new_n23369_, new_n23370_, new_n23371_,
    new_n23372_, new_n23373_, new_n23374_, new_n23375_, new_n23376_,
    new_n23377_, new_n23378_, new_n23379_, new_n23380_, new_n23381_,
    new_n23382_, new_n23383_, new_n23385_, new_n23386_, new_n23387_,
    new_n23388_, new_n23389_, new_n23390_, new_n23391_, new_n23392_,
    new_n23393_, new_n23394_, new_n23395_, new_n23396_, new_n23397_,
    new_n23398_, new_n23399_, new_n23400_, new_n23401_, new_n23402_,
    new_n23403_, new_n23404_, new_n23405_, new_n23406_, new_n23407_,
    new_n23408_, new_n23409_, new_n23410_, new_n23411_, new_n23412_,
    new_n23413_, new_n23414_, new_n23415_, new_n23416_, new_n23417_,
    new_n23418_, new_n23419_, new_n23420_, new_n23421_, new_n23422_,
    new_n23423_, new_n23424_, new_n23425_, new_n23426_, new_n23427_,
    new_n23428_, new_n23429_, new_n23430_, new_n23431_, new_n23432_,
    new_n23433_, new_n23434_, new_n23435_, new_n23436_, new_n23437_,
    new_n23438_, new_n23439_, new_n23440_, new_n23441_, new_n23442_,
    new_n23443_, new_n23444_, new_n23445_, new_n23446_, new_n23447_,
    new_n23448_, new_n23449_, new_n23450_, new_n23451_, new_n23452_,
    new_n23453_, new_n23454_, new_n23455_, new_n23456_, new_n23457_,
    new_n23458_, new_n23459_, new_n23460_, new_n23461_, new_n23462_,
    new_n23463_, new_n23464_, new_n23465_, new_n23466_, new_n23467_,
    new_n23468_, new_n23469_, new_n23470_, new_n23471_, new_n23472_,
    new_n23473_, new_n23474_, new_n23475_, new_n23476_, new_n23477_,
    new_n23478_, new_n23479_, new_n23480_, new_n23481_, new_n23482_,
    new_n23483_, new_n23484_, new_n23485_, new_n23486_, new_n23487_,
    new_n23488_, new_n23489_, new_n23490_, new_n23491_, new_n23492_,
    new_n23493_, new_n23494_, new_n23495_, new_n23496_, new_n23497_,
    new_n23498_, new_n23499_, new_n23500_, new_n23501_, new_n23502_,
    new_n23503_, new_n23504_, new_n23505_, new_n23506_, new_n23507_,
    new_n23508_, new_n23509_, new_n23510_, new_n23511_, new_n23512_,
    new_n23513_, new_n23514_, new_n23515_, new_n23516_, new_n23517_,
    new_n23518_, new_n23519_, new_n23520_, new_n23521_, new_n23522_,
    new_n23523_, new_n23524_, new_n23525_, new_n23526_, new_n23527_,
    new_n23528_, new_n23529_, new_n23530_, new_n23531_, new_n23532_,
    new_n23533_, new_n23534_, new_n23535_, new_n23536_, new_n23537_,
    new_n23538_, new_n23539_, new_n23540_, new_n23541_, new_n23542_,
    new_n23543_, new_n23544_, new_n23545_, new_n23546_, new_n23547_,
    new_n23548_, new_n23549_, new_n23550_, new_n23551_, new_n23552_,
    new_n23553_, new_n23554_, new_n23555_, new_n23556_, new_n23557_,
    new_n23558_, new_n23559_, new_n23560_, new_n23561_, new_n23562_,
    new_n23563_, new_n23564_, new_n23565_, new_n23566_, new_n23567_,
    new_n23568_, new_n23569_, new_n23570_, new_n23571_, new_n23572_,
    new_n23573_, new_n23574_, new_n23575_, new_n23576_, new_n23577_,
    new_n23578_, new_n23579_, new_n23580_, new_n23581_, new_n23582_,
    new_n23583_, new_n23584_, new_n23585_, new_n23586_, new_n23587_,
    new_n23588_, new_n23589_, new_n23590_, new_n23591_, new_n23592_,
    new_n23593_, new_n23594_, new_n23595_, new_n23596_, new_n23597_,
    new_n23598_, new_n23599_, new_n23600_, new_n23601_, new_n23602_,
    new_n23603_, new_n23604_, new_n23605_, new_n23606_, new_n23607_,
    new_n23608_, new_n23609_, new_n23610_, new_n23611_, new_n23612_,
    new_n23613_, new_n23614_, new_n23615_, new_n23616_, new_n23617_,
    new_n23618_, new_n23619_, new_n23620_, new_n23621_, new_n23622_,
    new_n23623_, new_n23624_, new_n23625_, new_n23626_, new_n23627_,
    new_n23628_, new_n23629_, new_n23630_, new_n23631_, new_n23632_,
    new_n23633_, new_n23634_, new_n23635_, new_n23636_, new_n23637_,
    new_n23638_, new_n23639_, new_n23640_, new_n23641_, new_n23642_,
    new_n23643_, new_n23644_, new_n23645_, new_n23646_, new_n23647_,
    new_n23648_, new_n23649_, new_n23650_, new_n23651_, new_n23652_,
    new_n23653_, new_n23654_, new_n23655_, new_n23656_, new_n23657_,
    new_n23658_, new_n23659_, new_n23660_, new_n23661_, new_n23662_,
    new_n23663_, new_n23664_, new_n23665_, new_n23666_, new_n23667_,
    new_n23668_, new_n23669_, new_n23670_, new_n23671_, new_n23672_,
    new_n23673_, new_n23674_, new_n23675_, new_n23676_, new_n23677_,
    new_n23678_, new_n23679_, new_n23680_, new_n23681_, new_n23682_,
    new_n23683_, new_n23684_, new_n23685_, new_n23686_, new_n23687_,
    new_n23688_, new_n23689_, new_n23690_, new_n23691_, new_n23692_,
    new_n23693_, new_n23694_, new_n23695_, new_n23696_, new_n23697_,
    new_n23698_, new_n23699_, new_n23700_, new_n23701_, new_n23702_,
    new_n23703_, new_n23704_, new_n23705_, new_n23706_, new_n23707_,
    new_n23708_, new_n23710_, new_n23711_, new_n23712_, new_n23713_,
    new_n23714_, new_n23715_, new_n23716_, new_n23717_, new_n23718_,
    new_n23719_, new_n23720_, new_n23721_, new_n23722_, new_n23723_,
    new_n23724_, new_n23725_, new_n23726_, new_n23727_, new_n23728_,
    new_n23729_, new_n23730_, new_n23731_, new_n23732_, new_n23733_,
    new_n23734_, new_n23735_, new_n23736_, new_n23737_, new_n23738_,
    new_n23739_, new_n23740_, new_n23741_, new_n23742_, new_n23743_,
    new_n23744_, new_n23745_, new_n23746_, new_n23747_, new_n23748_,
    new_n23749_, new_n23750_, new_n23751_, new_n23752_, new_n23753_,
    new_n23754_, new_n23755_, new_n23756_, new_n23757_, new_n23758_,
    new_n23759_, new_n23760_, new_n23761_, new_n23762_, new_n23763_,
    new_n23764_, new_n23765_, new_n23766_, new_n23767_, new_n23768_,
    new_n23769_, new_n23770_, new_n23771_, new_n23772_, new_n23773_,
    new_n23774_, new_n23775_, new_n23776_, new_n23777_, new_n23778_,
    new_n23779_, new_n23780_, new_n23781_, new_n23782_, new_n23783_,
    new_n23784_, new_n23785_, new_n23786_, new_n23787_, new_n23788_,
    new_n23789_, new_n23790_, new_n23791_, new_n23792_, new_n23793_,
    new_n23794_, new_n23795_, new_n23796_, new_n23797_, new_n23798_,
    new_n23799_, new_n23800_, new_n23801_, new_n23802_, new_n23803_,
    new_n23804_, new_n23805_, new_n23806_, new_n23807_, new_n23808_,
    new_n23809_, new_n23810_, new_n23811_, new_n23812_, new_n23813_,
    new_n23814_, new_n23815_, new_n23816_, new_n23817_, new_n23818_,
    new_n23819_, new_n23820_, new_n23821_, new_n23822_, new_n23823_,
    new_n23824_, new_n23825_, new_n23826_, new_n23827_, new_n23828_,
    new_n23829_, new_n23830_, new_n23831_, new_n23832_, new_n23833_,
    new_n23834_, new_n23835_, new_n23836_, new_n23837_, new_n23838_,
    new_n23839_, new_n23840_, new_n23841_, new_n23842_, new_n23843_,
    new_n23844_, new_n23845_, new_n23846_, new_n23847_, new_n23848_,
    new_n23849_, new_n23850_, new_n23851_, new_n23852_, new_n23853_,
    new_n23854_, new_n23855_, new_n23856_, new_n23857_, new_n23858_,
    new_n23859_, new_n23860_, new_n23861_, new_n23862_, new_n23863_,
    new_n23864_, new_n23865_, new_n23866_, new_n23867_, new_n23868_,
    new_n23869_, new_n23870_, new_n23871_, new_n23872_, new_n23873_,
    new_n23874_, new_n23875_, new_n23876_, new_n23877_, new_n23878_,
    new_n23879_, new_n23880_, new_n23881_, new_n23882_, new_n23883_,
    new_n23884_, new_n23885_, new_n23886_, new_n23887_, new_n23888_,
    new_n23889_, new_n23890_, new_n23891_, new_n23892_, new_n23893_,
    new_n23894_, new_n23895_, new_n23896_, new_n23897_, new_n23898_,
    new_n23899_, new_n23900_, new_n23901_, new_n23902_, new_n23903_,
    new_n23904_, new_n23905_, new_n23906_, new_n23907_, new_n23908_,
    new_n23909_, new_n23910_, new_n23911_, new_n23912_, new_n23913_,
    new_n23914_, new_n23915_, new_n23916_, new_n23917_, new_n23918_,
    new_n23919_, new_n23920_, new_n23921_, new_n23922_, new_n23923_,
    new_n23924_, new_n23925_, new_n23926_, new_n23927_, new_n23928_,
    new_n23929_, new_n23930_, new_n23931_, new_n23932_, new_n23933_,
    new_n23934_, new_n23935_, new_n23936_, new_n23937_, new_n23938_,
    new_n23939_, new_n23940_, new_n23941_, new_n23942_, new_n23943_,
    new_n23944_, new_n23945_, new_n23946_, new_n23947_, new_n23948_,
    new_n23949_, new_n23950_, new_n23951_, new_n23952_, new_n23953_,
    new_n23954_, new_n23955_, new_n23956_, new_n23957_, new_n23958_,
    new_n23959_, new_n23960_, new_n23961_, new_n23962_, new_n23963_,
    new_n23964_, new_n23965_, new_n23966_, new_n23967_, new_n23968_,
    new_n23969_, new_n23970_, new_n23971_, new_n23972_, new_n23973_,
    new_n23974_, new_n23975_, new_n23976_, new_n23977_, new_n23978_,
    new_n23979_, new_n23980_, new_n23981_, new_n23982_, new_n23983_,
    new_n23984_, new_n23985_, new_n23986_, new_n23987_, new_n23988_,
    new_n23989_, new_n23990_, new_n23991_, new_n23992_, new_n23993_,
    new_n23994_, new_n23995_, new_n23996_, new_n23997_, new_n23998_,
    new_n23999_, new_n24000_, new_n24001_, new_n24002_, new_n24003_,
    new_n24004_, new_n24005_, new_n24006_, new_n24007_, new_n24008_,
    new_n24009_, new_n24010_, new_n24011_, new_n24012_, new_n24013_,
    new_n24014_, new_n24015_, new_n24016_, new_n24017_, new_n24018_,
    new_n24019_, new_n24020_, new_n24021_, new_n24022_, new_n24023_,
    new_n24024_, new_n24025_, new_n24027_, new_n24028_, new_n24029_,
    new_n24030_, new_n24031_, new_n24032_, new_n24033_, new_n24034_,
    new_n24035_, new_n24036_, new_n24037_, new_n24038_, new_n24039_,
    new_n24040_, new_n24041_, new_n24042_, new_n24043_, new_n24044_,
    new_n24045_, new_n24046_, new_n24047_, new_n24048_, new_n24049_,
    new_n24050_, new_n24051_, new_n24052_, new_n24053_, new_n24054_,
    new_n24055_, new_n24056_, new_n24057_, new_n24058_, new_n24059_,
    new_n24060_, new_n24061_, new_n24062_, new_n24063_, new_n24064_,
    new_n24065_, new_n24066_, new_n24067_, new_n24068_, new_n24069_,
    new_n24070_, new_n24071_, new_n24072_, new_n24073_, new_n24074_,
    new_n24075_, new_n24076_, new_n24077_, new_n24078_, new_n24079_,
    new_n24080_, new_n24081_, new_n24082_, new_n24083_, new_n24084_,
    new_n24085_, new_n24086_, new_n24087_, new_n24088_, new_n24089_,
    new_n24090_, new_n24091_, new_n24092_, new_n24093_, new_n24094_,
    new_n24095_, new_n24096_, new_n24097_, new_n24098_, new_n24099_,
    new_n24100_, new_n24101_, new_n24102_, new_n24103_, new_n24104_,
    new_n24105_, new_n24106_, new_n24107_, new_n24108_, new_n24109_,
    new_n24110_, new_n24111_, new_n24112_, new_n24113_, new_n24114_,
    new_n24115_, new_n24116_, new_n24117_, new_n24118_, new_n24119_,
    new_n24120_, new_n24121_, new_n24122_, new_n24123_, new_n24124_,
    new_n24125_, new_n24126_, new_n24127_, new_n24128_, new_n24129_,
    new_n24130_, new_n24131_, new_n24132_, new_n24133_, new_n24134_,
    new_n24135_, new_n24136_, new_n24137_, new_n24138_, new_n24139_,
    new_n24140_, new_n24141_, new_n24142_, new_n24143_, new_n24144_,
    new_n24145_, new_n24146_, new_n24147_, new_n24148_, new_n24149_,
    new_n24150_, new_n24151_, new_n24152_, new_n24153_, new_n24154_,
    new_n24155_, new_n24156_, new_n24157_, new_n24158_, new_n24159_,
    new_n24160_, new_n24161_, new_n24162_, new_n24163_, new_n24164_,
    new_n24165_, new_n24166_, new_n24167_, new_n24168_, new_n24169_,
    new_n24170_, new_n24171_, new_n24172_, new_n24173_, new_n24174_,
    new_n24175_, new_n24176_, new_n24177_, new_n24178_, new_n24179_,
    new_n24180_, new_n24181_, new_n24182_, new_n24183_, new_n24184_,
    new_n24185_, new_n24186_, new_n24187_, new_n24188_, new_n24189_,
    new_n24190_, new_n24191_, new_n24192_, new_n24193_, new_n24194_,
    new_n24195_, new_n24196_, new_n24197_, new_n24198_, new_n24199_,
    new_n24200_, new_n24201_, new_n24202_, new_n24203_, new_n24204_,
    new_n24205_, new_n24206_, new_n24207_, new_n24208_, new_n24209_,
    new_n24210_, new_n24211_, new_n24212_, new_n24213_, new_n24214_,
    new_n24215_, new_n24216_, new_n24217_, new_n24218_, new_n24219_,
    new_n24220_, new_n24221_, new_n24222_, new_n24223_, new_n24224_,
    new_n24225_, new_n24226_, new_n24227_, new_n24228_, new_n24229_,
    new_n24230_, new_n24231_, new_n24232_, new_n24233_, new_n24234_,
    new_n24235_, new_n24236_, new_n24237_, new_n24238_, new_n24239_,
    new_n24240_, new_n24241_, new_n24242_, new_n24243_, new_n24244_,
    new_n24245_, new_n24246_, new_n24247_, new_n24248_, new_n24249_,
    new_n24250_, new_n24251_, new_n24252_, new_n24253_, new_n24254_,
    new_n24255_, new_n24256_, new_n24257_, new_n24258_, new_n24259_,
    new_n24260_, new_n24261_, new_n24262_, new_n24263_, new_n24264_,
    new_n24265_, new_n24266_, new_n24267_, new_n24268_, new_n24269_,
    new_n24270_, new_n24271_, new_n24272_, new_n24273_, new_n24274_,
    new_n24275_, new_n24276_, new_n24277_, new_n24278_, new_n24279_,
    new_n24280_, new_n24281_, new_n24282_, new_n24283_, new_n24284_,
    new_n24285_, new_n24286_, new_n24287_, new_n24288_, new_n24289_,
    new_n24290_, new_n24291_, new_n24292_, new_n24293_, new_n24294_,
    new_n24295_, new_n24296_, new_n24297_, new_n24298_, new_n24299_,
    new_n24300_, new_n24301_, new_n24302_, new_n24303_, new_n24304_,
    new_n24305_, new_n24306_, new_n24307_, new_n24308_, new_n24309_,
    new_n24310_, new_n24311_, new_n24312_, new_n24313_, new_n24314_,
    new_n24315_, new_n24316_, new_n24317_, new_n24318_, new_n24319_,
    new_n24320_, new_n24321_, new_n24322_, new_n24323_, new_n24324_,
    new_n24325_, new_n24326_, new_n24327_, new_n24328_, new_n24329_,
    new_n24330_, new_n24331_, new_n24332_, new_n24333_, new_n24334_,
    new_n24335_, new_n24336_, new_n24337_, new_n24338_, new_n24339_,
    new_n24340_, new_n24341_, new_n24342_, new_n24343_, new_n24344_,
    new_n24345_, new_n24346_, new_n24347_, new_n24348_, new_n24349_,
    new_n24350_, new_n24351_, new_n24352_, new_n24354_, new_n24355_,
    new_n24356_, new_n24357_, new_n24358_, new_n24359_, new_n24360_,
    new_n24361_, new_n24362_, new_n24363_, new_n24364_, new_n24365_,
    new_n24366_, new_n24367_, new_n24368_, new_n24369_, new_n24370_,
    new_n24371_, new_n24372_, new_n24373_, new_n24374_, new_n24375_,
    new_n24376_, new_n24377_, new_n24378_, new_n24379_, new_n24380_,
    new_n24381_, new_n24383_, new_n24384_, new_n24385_, new_n24386_,
    new_n24387_, new_n24388_, new_n24389_, new_n24390_, new_n24391_,
    new_n24392_, new_n24393_, new_n24394_, new_n24395_, new_n24396_,
    new_n24397_, new_n24398_, new_n24399_, new_n24400_, new_n24401_,
    new_n24402_, new_n24403_, new_n24404_, new_n24405_, new_n24406_,
    new_n24407_, new_n24408_, new_n24409_, new_n24410_, new_n24411_,
    new_n24412_, new_n24413_, new_n24414_, new_n24415_, new_n24416_,
    new_n24417_, new_n24418_, new_n24419_, new_n24420_, new_n24421_,
    new_n24422_, new_n24423_, new_n24425_, new_n24426_, new_n24427_,
    new_n24428_, new_n24429_, new_n24430_, new_n24431_, new_n24432_,
    new_n24433_, new_n24434_, new_n24435_, new_n24436_, new_n24437_,
    new_n24438_, new_n24439_, new_n24440_, new_n24441_, new_n24442_,
    new_n24443_, new_n24444_, new_n24445_, new_n24446_, new_n24447_,
    new_n24448_, new_n24449_, new_n24450_, new_n24451_, new_n24452_,
    new_n24453_, new_n24454_, new_n24455_, new_n24456_, new_n24457_,
    new_n24458_, new_n24459_, new_n24460_, new_n24461_, new_n24462_,
    new_n24464_, new_n24465_, new_n24466_, new_n24467_, new_n24468_,
    new_n24469_, new_n24470_, new_n24471_, new_n24472_, new_n24473_,
    new_n24474_, new_n24475_, new_n24476_, new_n24477_, new_n24478_,
    new_n24479_, new_n24480_, new_n24481_, new_n24482_, new_n24483_,
    new_n24484_, new_n24485_, new_n24486_, new_n24487_, new_n24488_,
    new_n24489_, new_n24490_, new_n24491_, new_n24492_, new_n24493_,
    new_n24494_, new_n24495_, new_n24496_, new_n24497_, new_n24498_,
    new_n24499_, new_n24500_, new_n24501_, new_n24502_, new_n24503_,
    new_n24504_, new_n24505_, new_n24506_, new_n24507_, new_n24508_,
    new_n24509_, new_n24510_, new_n24511_, new_n24512_, new_n24513_,
    new_n24514_, new_n24515_, new_n24516_, new_n24517_, new_n24518_,
    new_n24519_, new_n24520_, new_n24521_, new_n24522_, new_n24523_,
    new_n24524_, new_n24525_, new_n24526_, new_n24527_, new_n24528_,
    new_n24529_, new_n24530_, new_n24531_, new_n24532_, new_n24533_,
    new_n24534_, new_n24535_, new_n24536_, new_n24537_, new_n24538_,
    new_n24539_, new_n24540_, new_n24541_, new_n24542_, new_n24543_,
    new_n24544_, new_n24545_, new_n24546_, new_n24547_, new_n24548_,
    new_n24549_, new_n24550_, new_n24551_, new_n24552_, new_n24553_,
    new_n24554_, new_n24555_, new_n24556_, new_n24557_, new_n24558_,
    new_n24559_, new_n24560_, new_n24561_, new_n24562_, new_n24563_,
    new_n24564_, new_n24565_, new_n24566_, new_n24567_, new_n24568_,
    new_n24569_, new_n24570_, new_n24571_, new_n24572_, new_n24573_,
    new_n24574_, new_n24575_, new_n24576_, new_n24577_, new_n24578_,
    new_n24579_, new_n24580_, new_n24581_, new_n24582_, new_n24583_,
    new_n24584_, new_n24585_, new_n24586_, new_n24587_, new_n24588_,
    new_n24589_, new_n24590_, new_n24591_, new_n24592_, new_n24593_,
    new_n24594_, new_n24595_, new_n24596_, new_n24597_, new_n24598_,
    new_n24599_, new_n24600_, new_n24601_, new_n24602_, new_n24603_,
    new_n24604_, new_n24605_, new_n24606_, new_n24607_, new_n24608_,
    new_n24609_, new_n24610_, new_n24611_, new_n24612_, new_n24613_,
    new_n24614_, new_n24615_, new_n24616_, new_n24617_, new_n24618_,
    new_n24619_, new_n24620_, new_n24621_, new_n24622_, new_n24623_,
    new_n24624_, new_n24625_, new_n24626_, new_n24627_, new_n24628_,
    new_n24629_, new_n24630_, new_n24631_, new_n24632_, new_n24633_,
    new_n24634_, new_n24635_, new_n24636_, new_n24637_, new_n24638_,
    new_n24639_, new_n24640_, new_n24641_, new_n24642_, new_n24643_,
    new_n24644_, new_n24645_, new_n24646_, new_n24647_, new_n24648_,
    new_n24649_, new_n24650_, new_n24651_, new_n24652_, new_n24653_,
    new_n24654_, new_n24655_, new_n24656_, new_n24657_, new_n24658_,
    new_n24659_, new_n24660_, new_n24661_, new_n24662_, new_n24663_,
    new_n24664_, new_n24665_, new_n24666_, new_n24667_, new_n24668_,
    new_n24669_, new_n24670_, new_n24671_, new_n24672_, new_n24673_,
    new_n24674_, new_n24675_, new_n24676_, new_n24677_, new_n24678_,
    new_n24679_, new_n24680_, new_n24681_, new_n24682_, new_n24683_,
    new_n24684_, new_n24685_, new_n24686_, new_n24687_, new_n24688_,
    new_n24689_, new_n24690_, new_n24691_, new_n24692_, new_n24693_,
    new_n24694_, new_n24695_, new_n24696_, new_n24697_, new_n24698_,
    new_n24699_, new_n24700_, new_n24701_, new_n24702_, new_n24703_,
    new_n24704_, new_n24705_, new_n24706_, new_n24707_, new_n24708_,
    new_n24709_, new_n24710_, new_n24711_, new_n24712_, new_n24713_,
    new_n24714_, new_n24715_, new_n24716_, new_n24717_, new_n24718_,
    new_n24719_, new_n24720_, new_n24721_, new_n24722_, new_n24723_,
    new_n24724_, new_n24725_, new_n24726_, new_n24727_, new_n24728_,
    new_n24729_, new_n24730_, new_n24731_, new_n24732_, new_n24733_,
    new_n24734_, new_n24735_, new_n24736_, new_n24737_, new_n24738_,
    new_n24739_, new_n24740_, new_n24741_, new_n24742_, new_n24743_,
    new_n24744_, new_n24745_, new_n24746_, new_n24747_, new_n24748_,
    new_n24749_, new_n24750_, new_n24751_, new_n24752_, new_n24753_,
    new_n24754_, new_n24755_, new_n24756_, new_n24757_, new_n24758_,
    new_n24759_, new_n24760_, new_n24761_, new_n24762_, new_n24763_,
    new_n24764_, new_n24765_, new_n24766_, new_n24767_, new_n24768_,
    new_n24769_, new_n24770_, new_n24771_, new_n24772_, new_n24773_,
    new_n24774_, new_n24775_, new_n24776_, new_n24777_, new_n24778_,
    new_n24779_, new_n24780_, new_n24781_, new_n24782_, new_n24783_,
    new_n24784_, new_n24785_, new_n24786_, new_n24787_, new_n24788_,
    new_n24789_, new_n24790_, new_n24791_, new_n24792_, new_n24793_,
    new_n24794_, new_n24795_, new_n24796_, new_n24797_, new_n24798_,
    new_n24799_, new_n24800_, new_n24801_, new_n24802_, new_n24803_,
    new_n24804_, new_n24805_, new_n24806_, new_n24807_, new_n24808_,
    new_n24809_, new_n24810_, new_n24811_, new_n24812_, new_n24813_,
    new_n24814_, new_n24815_, new_n24816_, new_n24817_, new_n24818_,
    new_n24819_, new_n24820_, new_n24821_, new_n24822_, new_n24823_,
    new_n24824_, new_n24825_, new_n24826_, new_n24827_, new_n24828_,
    new_n24829_, new_n24830_, new_n24831_, new_n24832_, new_n24833_,
    new_n24834_, new_n24835_, new_n24836_, new_n24837_, new_n24838_,
    new_n24839_, new_n24840_, new_n24841_, new_n24842_, new_n24843_,
    new_n24844_, new_n24845_, new_n24846_, new_n24847_, new_n24848_,
    new_n24849_, new_n24850_, new_n24851_, new_n24852_, new_n24853_,
    new_n24854_, new_n24855_, new_n24856_, new_n24857_, new_n24858_,
    new_n24859_, new_n24860_, new_n24861_, new_n24862_, new_n24863_,
    new_n24864_, new_n24865_, new_n24866_, new_n24867_, new_n24868_,
    new_n24869_, new_n24870_, new_n24871_, new_n24872_, new_n24873_,
    new_n24874_, new_n24875_, new_n24876_, new_n24877_, new_n24878_,
    new_n24879_, new_n24880_, new_n24881_, new_n24882_, new_n24883_,
    new_n24884_, new_n24885_, new_n24886_, new_n24887_, new_n24888_,
    new_n24889_, new_n24890_, new_n24891_, new_n24892_, new_n24893_,
    new_n24894_, new_n24895_, new_n24896_, new_n24897_, new_n24898_,
    new_n24899_, new_n24900_, new_n24901_, new_n24902_, new_n24903_,
    new_n24904_, new_n24905_, new_n24906_, new_n24907_, new_n24908_,
    new_n24909_, new_n24910_, new_n24911_, new_n24912_, new_n24913_,
    new_n24914_, new_n24915_, new_n24916_, new_n24917_, new_n24918_,
    new_n24919_, new_n24920_, new_n24921_, new_n24922_, new_n24923_,
    new_n24924_, new_n24925_, new_n24926_, new_n24927_, new_n24928_,
    new_n24930_, new_n24931_, new_n24932_, new_n24933_, new_n24934_,
    new_n24935_, new_n24936_, new_n24937_, new_n24938_, new_n24939_,
    new_n24940_, new_n24941_, new_n24942_, new_n24943_, new_n24944_,
    new_n24945_, new_n24946_, new_n24947_, new_n24948_, new_n24949_,
    new_n24950_, new_n24951_, new_n24952_, new_n24953_, new_n24954_,
    new_n24955_, new_n24956_, new_n24957_, new_n24958_, new_n24959_,
    new_n24960_, new_n24961_, new_n24962_, new_n24963_, new_n24964_,
    new_n24965_, new_n24966_, new_n24967_, new_n24968_, new_n24969_,
    new_n24970_, new_n24971_, new_n24972_, new_n24973_, new_n24974_,
    new_n24975_, new_n24976_, new_n24977_, new_n24978_, new_n24979_,
    new_n24980_, new_n24981_, new_n24982_, new_n24983_, new_n24984_,
    new_n24985_, new_n24986_, new_n24987_, new_n24988_, new_n24989_,
    new_n24990_, new_n24991_, new_n24992_, new_n24993_, new_n24994_,
    new_n24995_, new_n24996_, new_n24997_, new_n24998_, new_n24999_,
    new_n25000_, new_n25001_, new_n25002_, new_n25003_, new_n25004_,
    new_n25005_, new_n25006_, new_n25007_, new_n25008_, new_n25009_,
    new_n25010_, new_n25011_, new_n25012_, new_n25013_, new_n25014_,
    new_n25015_, new_n25016_, new_n25017_, new_n25018_, new_n25019_,
    new_n25020_, new_n25021_, new_n25022_, new_n25023_, new_n25024_,
    new_n25025_, new_n25026_, new_n25027_, new_n25028_, new_n25029_,
    new_n25030_, new_n25031_, new_n25032_, new_n25033_, new_n25034_,
    new_n25035_, new_n25036_, new_n25037_, new_n25038_, new_n25039_,
    new_n25040_, new_n25041_, new_n25042_, new_n25043_, new_n25044_,
    new_n25045_, new_n25046_, new_n25047_, new_n25048_, new_n25049_,
    new_n25050_, new_n25051_, new_n25052_, new_n25053_, new_n25054_,
    new_n25055_, new_n25056_, new_n25057_, new_n25058_, new_n25059_,
    new_n25060_, new_n25061_, new_n25062_, new_n25063_, new_n25064_,
    new_n25065_, new_n25066_, new_n25067_, new_n25068_, new_n25069_,
    new_n25070_, new_n25071_, new_n25072_, new_n25073_, new_n25074_,
    new_n25075_, new_n25076_, new_n25077_, new_n25078_, new_n25079_,
    new_n25080_, new_n25081_, new_n25082_, new_n25083_, new_n25084_,
    new_n25085_, new_n25086_, new_n25087_, new_n25088_, new_n25089_,
    new_n25090_, new_n25091_, new_n25092_, new_n25093_, new_n25094_,
    new_n25095_, new_n25096_, new_n25097_, new_n25098_, new_n25099_,
    new_n25100_, new_n25101_, new_n25102_, new_n25103_, new_n25104_,
    new_n25105_, new_n25106_, new_n25107_, new_n25108_, new_n25109_,
    new_n25110_, new_n25111_, new_n25112_, new_n25113_, new_n25114_,
    new_n25115_, new_n25116_, new_n25117_, new_n25118_, new_n25119_,
    new_n25120_, new_n25121_, new_n25122_, new_n25123_, new_n25124_,
    new_n25126_, new_n25127_, new_n25128_, new_n25129_, new_n25130_,
    new_n25131_, new_n25132_, new_n25133_, new_n25134_, new_n25135_,
    new_n25136_, new_n25137_, new_n25138_, new_n25139_, new_n25140_,
    new_n25141_, new_n25142_, new_n25143_, new_n25144_, new_n25145_,
    new_n25146_, new_n25147_, new_n25148_, new_n25149_, new_n25150_,
    new_n25151_, new_n25152_, new_n25153_, new_n25154_, new_n25155_,
    new_n25156_, new_n25157_, new_n25158_, new_n25159_, new_n25160_,
    new_n25161_, new_n25162_, new_n25163_, new_n25164_, new_n25165_,
    new_n25166_, new_n25167_, new_n25168_, new_n25169_, new_n25170_,
    new_n25171_, new_n25172_, new_n25173_, new_n25174_, new_n25175_,
    new_n25176_, new_n25177_, new_n25178_, new_n25179_, new_n25180_,
    new_n25181_, new_n25182_, new_n25183_, new_n25184_, new_n25185_,
    new_n25186_, new_n25187_, new_n25188_, new_n25189_, new_n25190_,
    new_n25191_, new_n25192_, new_n25193_, new_n25194_, new_n25195_,
    new_n25196_, new_n25197_, new_n25198_, new_n25199_, new_n25200_,
    new_n25201_, new_n25202_, new_n25203_, new_n25204_, new_n25205_,
    new_n25206_, new_n25207_, new_n25208_, new_n25209_, new_n25210_,
    new_n25211_, new_n25212_, new_n25213_, new_n25214_, new_n25215_,
    new_n25216_, new_n25217_, new_n25218_, new_n25219_, new_n25220_,
    new_n25221_, new_n25222_, new_n25223_, new_n25224_, new_n25225_,
    new_n25226_, new_n25227_, new_n25228_, new_n25229_, new_n25230_,
    new_n25231_, new_n25232_, new_n25233_, new_n25234_, new_n25235_,
    new_n25236_, new_n25237_, new_n25238_, new_n25239_, new_n25240_,
    new_n25241_, new_n25242_, new_n25243_, new_n25244_, new_n25245_,
    new_n25246_, new_n25247_, new_n25248_, new_n25249_, new_n25250_,
    new_n25251_, new_n25252_, new_n25253_, new_n25254_, new_n25255_,
    new_n25256_, new_n25257_, new_n25258_, new_n25259_, new_n25260_,
    new_n25261_, new_n25262_, new_n25263_, new_n25264_, new_n25265_,
    new_n25266_, new_n25267_, new_n25268_, new_n25269_, new_n25270_,
    new_n25271_, new_n25272_, new_n25273_, new_n25274_, new_n25275_,
    new_n25276_, new_n25277_, new_n25278_, new_n25279_, new_n25280_,
    new_n25281_, new_n25282_, new_n25283_, new_n25284_, new_n25285_,
    new_n25286_, new_n25287_, new_n25288_, new_n25289_, new_n25290_,
    new_n25291_, new_n25292_, new_n25293_, new_n25294_, new_n25295_,
    new_n25296_, new_n25297_, new_n25298_, new_n25299_, new_n25300_,
    new_n25301_, new_n25302_, new_n25303_, new_n25304_, new_n25305_,
    new_n25306_, new_n25307_, new_n25308_, new_n25309_, new_n25310_,
    new_n25311_, new_n25312_, new_n25313_, new_n25314_, new_n25315_,
    new_n25316_, new_n25317_, new_n25319_, new_n25320_, new_n25321_,
    new_n25322_, new_n25323_, new_n25324_, new_n25325_, new_n25326_,
    new_n25327_, new_n25328_, new_n25329_, new_n25330_, new_n25331_,
    new_n25332_, new_n25333_, new_n25334_, new_n25335_, new_n25336_,
    new_n25337_, new_n25338_, new_n25339_, new_n25340_, new_n25341_,
    new_n25342_, new_n25343_, new_n25344_, new_n25345_, new_n25346_,
    new_n25347_, new_n25348_, new_n25349_, new_n25350_, new_n25351_,
    new_n25352_, new_n25353_, new_n25354_, new_n25355_, new_n25356_,
    new_n25357_, new_n25358_, new_n25359_, new_n25360_, new_n25361_,
    new_n25362_, new_n25363_, new_n25364_, new_n25365_, new_n25366_,
    new_n25367_, new_n25368_, new_n25369_, new_n25370_, new_n25371_,
    new_n25372_, new_n25373_, new_n25374_, new_n25375_, new_n25376_,
    new_n25377_, new_n25378_, new_n25379_, new_n25380_, new_n25381_,
    new_n25382_, new_n25383_, new_n25384_, new_n25385_, new_n25386_,
    new_n25387_, new_n25388_, new_n25389_, new_n25390_, new_n25391_,
    new_n25392_, new_n25393_, new_n25394_, new_n25395_, new_n25396_,
    new_n25397_, new_n25398_, new_n25399_, new_n25400_, new_n25401_,
    new_n25402_, new_n25403_, new_n25404_, new_n25405_, new_n25406_,
    new_n25407_, new_n25408_, new_n25409_, new_n25410_, new_n25411_,
    new_n25412_, new_n25413_, new_n25414_, new_n25415_, new_n25416_,
    new_n25417_, new_n25418_, new_n25419_, new_n25420_, new_n25421_,
    new_n25422_, new_n25423_, new_n25424_, new_n25425_, new_n25426_,
    new_n25427_, new_n25428_, new_n25429_, new_n25430_, new_n25431_,
    new_n25432_, new_n25433_, new_n25434_, new_n25435_, new_n25436_,
    new_n25437_, new_n25438_, new_n25439_, new_n25440_, new_n25441_,
    new_n25442_, new_n25443_, new_n25444_, new_n25445_, new_n25446_,
    new_n25447_, new_n25448_, new_n25449_, new_n25450_, new_n25451_,
    new_n25452_, new_n25453_, new_n25454_, new_n25455_, new_n25456_,
    new_n25458_, new_n25459_, new_n25460_, new_n25461_, new_n25462_,
    new_n25463_, new_n25465_, new_n25466_, new_n25467_, new_n25468_,
    new_n25469_, new_n25470_, new_n25472_, new_n25473_, new_n25474_,
    new_n25475_, new_n25476_, new_n25477_, new_n25478_, new_n25479_,
    new_n25480_, new_n25481_, new_n25482_, new_n25483_, new_n25484_,
    new_n25485_, new_n25486_, new_n25487_, new_n25488_, new_n25489_,
    new_n25490_, new_n25491_, new_n25492_, new_n25493_, new_n25494_,
    new_n25495_, new_n25496_, new_n25497_, new_n25498_, new_n25499_,
    new_n25500_, new_n25501_, new_n25502_, new_n25503_, new_n25504_,
    new_n25505_, new_n25506_, new_n25507_, new_n25508_, new_n25509_,
    new_n25510_, new_n25511_, new_n25512_, new_n25513_, new_n25514_,
    new_n25515_, new_n25516_, new_n25517_, new_n25518_, new_n25519_,
    new_n25520_, new_n25521_, new_n25522_, new_n25523_, new_n25524_,
    new_n25525_, new_n25526_, new_n25527_, new_n25528_, new_n25529_,
    new_n25530_, new_n25531_, new_n25532_, new_n25533_, new_n25534_,
    new_n25535_, new_n25536_, new_n25537_, new_n25538_, new_n25539_,
    new_n25540_, new_n25541_, new_n25542_, new_n25543_, new_n25544_,
    new_n25545_, new_n25547_, new_n25548_, new_n25549_, new_n25550_,
    new_n25552_, new_n25553_, new_n25554_, new_n25555_, new_n25556_,
    new_n25557_, new_n25559_, new_n25560_, new_n25561_, new_n25562_,
    new_n25563_, new_n25564_, new_n25565_, new_n25566_, new_n25567_,
    new_n25568_, new_n25569_, new_n25570_, new_n25571_, new_n25572_,
    new_n25573_, new_n25574_, new_n25575_, new_n25576_, new_n25577_,
    new_n25578_, new_n25579_, new_n25580_, new_n25581_, new_n25582_,
    new_n25583_, new_n25584_, new_n25585_, new_n25586_, new_n25587_,
    new_n25588_, new_n25589_, new_n25590_, new_n25591_, new_n25592_,
    new_n25593_, new_n25594_, new_n25595_, new_n25596_, new_n25597_,
    new_n25598_, new_n25599_, new_n25600_, new_n25601_, new_n25602_,
    new_n25603_, new_n25604_, new_n25605_, new_n25606_, new_n25607_,
    new_n25608_, new_n25609_, new_n25610_, new_n25611_, new_n25612_,
    new_n25613_, new_n25614_, new_n25615_, new_n25616_, new_n25617_,
    new_n25618_, new_n25619_, new_n25620_, new_n25621_, new_n25622_,
    new_n25623_, new_n25624_, new_n25625_, new_n25626_, new_n25627_,
    new_n25628_, new_n25629_, new_n25630_, new_n25631_, new_n25632_,
    new_n25633_, new_n25634_, new_n25635_, new_n25636_, new_n25637_,
    new_n25638_, new_n25639_, new_n25640_, new_n25641_, new_n25642_,
    new_n25643_, new_n25644_, new_n25645_, new_n25646_, new_n25647_,
    new_n25648_, new_n25649_, new_n25650_, new_n25651_, new_n25652_,
    new_n25653_, new_n25654_, new_n25655_, new_n25656_, new_n25657_,
    new_n25658_, new_n25659_, new_n25660_, new_n25661_, new_n25662_,
    new_n25663_, new_n25664_, new_n25665_, new_n25666_, new_n25667_,
    new_n25668_, new_n25669_, new_n25670_, new_n25671_, new_n25672_,
    new_n25673_, new_n25674_, new_n25675_, new_n25676_, new_n25677_,
    new_n25678_, new_n25679_, new_n25680_, new_n25681_, new_n25682_,
    new_n25683_, new_n25684_, new_n25685_, new_n25686_, new_n25687_,
    new_n25688_, new_n25689_, new_n25690_, new_n25691_, new_n25692_,
    new_n25693_, new_n25694_, new_n25695_, new_n25696_, new_n25697_,
    new_n25698_, new_n25699_, new_n25700_, new_n25701_, new_n25702_,
    new_n25703_, new_n25704_, new_n25705_, new_n25706_, new_n25707_,
    new_n25708_, new_n25709_, new_n25710_, new_n25711_, new_n25712_,
    new_n25713_, new_n25714_, new_n25715_, new_n25716_, new_n25717_,
    new_n25718_, new_n25719_, new_n25720_, new_n25721_, new_n25722_,
    new_n25723_, new_n25724_, new_n25725_, new_n25726_, new_n25727_,
    new_n25728_, new_n25729_, new_n25730_, new_n25731_, new_n25732_,
    new_n25733_, new_n25734_, new_n25735_, new_n25736_, new_n25737_,
    new_n25738_, new_n25739_, new_n25740_, new_n25741_, new_n25742_,
    new_n25743_, new_n25744_, new_n25745_, new_n25746_, new_n25747_,
    new_n25748_, new_n25749_, new_n25750_, new_n25751_, new_n25752_,
    new_n25753_, new_n25754_, new_n25755_, new_n25756_, new_n25757_,
    new_n25758_, new_n25759_, new_n25760_, new_n25761_, new_n25762_,
    new_n25763_, new_n25764_, new_n25765_, new_n25766_, new_n25767_,
    new_n25768_, new_n25769_, new_n25770_, new_n25771_, new_n25772_,
    new_n25773_, new_n25774_, new_n25775_, new_n25776_, new_n25777_,
    new_n25778_, new_n25779_, new_n25780_, new_n25781_, new_n25782_,
    new_n25783_, new_n25784_, new_n25785_, new_n25786_, new_n25787_,
    new_n25788_, new_n25789_, new_n25790_, new_n25791_, new_n25792_,
    new_n25793_, new_n25794_, new_n25795_, new_n25796_, new_n25797_,
    new_n25798_, new_n25799_, new_n25800_, new_n25801_, new_n25802_,
    new_n25803_, new_n25804_, new_n25805_, new_n25806_, new_n25807_,
    new_n25808_, new_n25809_, new_n25810_, new_n25811_, new_n25812_,
    new_n25813_, new_n25814_, new_n25815_, new_n25816_, new_n25817_,
    new_n25818_, new_n25819_, new_n25820_, new_n25821_, new_n25822_,
    new_n25823_, new_n25824_, new_n25825_, new_n25826_, new_n25827_,
    new_n25828_, new_n25829_, new_n25830_, new_n25831_, new_n25832_,
    new_n25833_, new_n25834_, new_n25835_, new_n25836_, new_n25837_,
    new_n25838_, new_n25839_, new_n25840_, new_n25841_, new_n25842_,
    new_n25843_, new_n25844_, new_n25845_, new_n25846_, new_n25847_,
    new_n25848_, new_n25849_, new_n25850_, new_n25851_, new_n25852_,
    new_n25853_, new_n25854_, new_n25855_, new_n25856_, new_n25857_,
    new_n25858_, new_n25859_, new_n25860_, new_n25861_, new_n25862_,
    new_n25863_, new_n25864_, new_n25865_, new_n25866_, new_n25867_,
    new_n25868_, new_n25869_, new_n25870_, new_n25871_, new_n25872_,
    new_n25873_, new_n25874_, new_n25875_, new_n25876_, new_n25877_,
    new_n25878_, new_n25879_, new_n25880_, new_n25881_, new_n25882_,
    new_n25883_, new_n25884_, new_n25885_, new_n25886_, new_n25887_,
    new_n25888_, new_n25889_, new_n25890_, new_n25891_, new_n25892_,
    new_n25893_, new_n25894_, new_n25895_, new_n25896_, new_n25897_,
    new_n25898_, new_n25899_, new_n25900_, new_n25901_, new_n25902_,
    new_n25903_, new_n25904_, new_n25905_, new_n25906_, new_n25907_,
    new_n25908_, new_n25909_, new_n25910_, new_n25911_, new_n25912_,
    new_n25914_, new_n25915_, new_n25916_, new_n25917_, new_n25918_,
    new_n25919_, new_n25920_, new_n25921_, new_n25922_, new_n25923_,
    new_n25924_, new_n25925_, new_n25926_, new_n25927_, new_n25928_,
    new_n25929_, new_n25930_, new_n25931_, new_n25932_, new_n25933_,
    new_n25934_, new_n25935_, new_n25936_, new_n25937_, new_n25938_,
    new_n25939_, new_n25940_, new_n25941_, new_n25942_, new_n25943_,
    new_n25944_, new_n25945_, new_n25946_, new_n25947_, new_n25948_,
    new_n25949_, new_n25950_, new_n25951_, new_n25952_, new_n25953_,
    new_n25954_, new_n25955_, new_n25956_, new_n25957_, new_n25958_,
    new_n25959_, new_n25960_, new_n25961_, new_n25962_, new_n25963_,
    new_n25964_, new_n25966_, new_n25967_, new_n25968_, new_n25969_,
    new_n25970_, new_n25971_, new_n25972_, new_n25973_, new_n25974_,
    new_n25975_, new_n25976_, new_n25977_, new_n25978_, new_n25979_,
    new_n25980_, new_n25981_, new_n25982_, new_n25983_, new_n25984_,
    new_n25985_, new_n25986_, new_n25987_, new_n25988_, new_n25989_,
    new_n25990_, new_n25991_, new_n25992_, new_n25993_, new_n25994_,
    new_n25995_, new_n25996_, new_n25997_, new_n25998_, new_n25999_,
    new_n26000_, new_n26001_, new_n26002_, new_n26003_, new_n26004_,
    new_n26005_, new_n26006_, new_n26007_, new_n26008_, new_n26009_,
    new_n26010_, new_n26011_, new_n26012_, new_n26013_, new_n26014_,
    new_n26015_, new_n26016_, new_n26017_, new_n26018_, new_n26019_,
    new_n26020_, new_n26021_, new_n26022_, new_n26023_, new_n26024_,
    new_n26025_, new_n26026_, new_n26027_, new_n26028_, new_n26029_,
    new_n26030_, new_n26031_, new_n26032_, new_n26033_, new_n26034_,
    new_n26035_, new_n26036_, new_n26037_, new_n26038_, new_n26039_,
    new_n26040_, new_n26041_, new_n26042_, new_n26043_, new_n26044_,
    new_n26045_, new_n26046_, new_n26047_, new_n26048_, new_n26049_,
    new_n26050_, new_n26051_, new_n26052_, new_n26053_, new_n26054_,
    new_n26055_, new_n26056_, new_n26057_, new_n26058_, new_n26059_,
    new_n26060_, new_n26061_, new_n26062_, new_n26063_, new_n26064_,
    new_n26065_, new_n26066_, new_n26067_, new_n26068_, new_n26069_,
    new_n26071_, new_n26072_, new_n26073_, new_n26074_, new_n26075_,
    new_n26076_, new_n26077_, new_n26078_, new_n26079_, new_n26080_,
    new_n26081_, new_n26082_, new_n26083_, new_n26084_, new_n26085_,
    new_n26086_, new_n26087_, new_n26088_, new_n26089_, new_n26090_,
    new_n26091_, new_n26092_, new_n26093_, new_n26094_, new_n26095_,
    new_n26096_, new_n26097_, new_n26098_, new_n26099_, new_n26100_,
    new_n26101_, new_n26102_, new_n26103_, new_n26104_, new_n26105_,
    new_n26106_, new_n26107_, new_n26108_, new_n26109_, new_n26110_,
    new_n26111_, new_n26112_, new_n26113_, new_n26114_, new_n26115_,
    new_n26116_, new_n26117_, new_n26118_, new_n26119_, new_n26120_,
    new_n26121_, new_n26122_, new_n26123_, new_n26124_, new_n26125_,
    new_n26126_, new_n26127_, new_n26128_, new_n26129_, new_n26130_,
    new_n26131_, new_n26132_, new_n26133_, new_n26134_, new_n26135_,
    new_n26136_, new_n26137_, new_n26138_, new_n26139_, new_n26140_,
    new_n26141_, new_n26142_, new_n26143_, new_n26144_, new_n26145_,
    new_n26146_, new_n26147_, new_n26148_, new_n26149_, new_n26150_,
    new_n26151_, new_n26152_, new_n26153_, new_n26154_, new_n26155_,
    new_n26156_, new_n26157_, new_n26159_, new_n26160_, new_n26161_,
    new_n26162_, new_n26163_, new_n26164_, new_n26165_, new_n26166_,
    new_n26167_, new_n26168_, new_n26169_, new_n26170_, new_n26171_,
    new_n26172_, new_n26173_, new_n26174_, new_n26175_, new_n26176_,
    new_n26177_, new_n26179_, new_n26180_, new_n26181_, new_n26182_,
    new_n26183_, new_n26184_, new_n26185_, new_n26186_, new_n26187_,
    new_n26188_, new_n26189_, new_n26190_, new_n26191_, new_n26193_,
    new_n26194_, new_n26195_, new_n26196_, new_n26197_, new_n26198_,
    new_n26199_, new_n26200_, new_n26201_, new_n26202_, new_n26203_,
    new_n26204_, new_n26205_, new_n26206_, new_n26207_, new_n26209_,
    new_n26210_, new_n26211_, new_n26212_, new_n26213_, new_n26214_,
    new_n26215_, new_n26216_, new_n26217_, new_n26218_, new_n26219_,
    new_n26220_, new_n26221_, new_n26223_, new_n26224_, new_n26225_,
    new_n26226_, new_n26227_, new_n26228_, new_n26229_, new_n26230_,
    new_n26231_, new_n26232_, new_n26233_, new_n26234_, new_n26235_,
    new_n26236_, new_n26237_, new_n26238_, new_n26239_, new_n26240_,
    new_n26241_, new_n26242_, new_n26243_, new_n26244_, new_n26245_,
    new_n26246_, new_n26247_, new_n26248_, new_n26249_, new_n26250_,
    new_n26251_, new_n26252_, new_n26253_, new_n26254_, new_n26255_,
    new_n26256_, new_n26257_, new_n26258_, new_n26259_, new_n26260_,
    new_n26261_, new_n26262_, new_n26263_, new_n26264_, new_n26265_,
    new_n26266_, new_n26267_, new_n26268_, new_n26269_, new_n26270_,
    new_n26271_, new_n26272_, new_n26273_, new_n26274_, new_n26275_,
    new_n26276_, new_n26277_, new_n26278_, new_n26279_, new_n26280_,
    new_n26281_, new_n26282_, new_n26283_, new_n26284_, new_n26285_,
    new_n26286_, new_n26287_, new_n26288_, new_n26289_, new_n26290_,
    new_n26291_, new_n26292_, new_n26293_, new_n26294_, new_n26295_,
    new_n26296_, new_n26297_, new_n26298_, new_n26300_, new_n26301_,
    new_n26302_, new_n26303_, new_n26304_, new_n26305_, new_n26306_,
    new_n26307_, new_n26308_, new_n26309_, new_n26310_, new_n26311_,
    new_n26312_, new_n26313_, new_n26314_, new_n26315_, new_n26316_,
    new_n26317_, new_n26318_, new_n26319_, new_n26320_, new_n26321_,
    new_n26322_, new_n26323_, new_n26324_, new_n26325_, new_n26326_,
    new_n26327_, new_n26328_, new_n26329_, new_n26330_, new_n26331_,
    new_n26332_, new_n26333_, new_n26334_, new_n26335_, new_n26336_,
    new_n26337_, new_n26338_, new_n26339_, new_n26340_, new_n26341_,
    new_n26342_, new_n26343_, new_n26344_, new_n26345_, new_n26346_,
    new_n26347_, new_n26348_, new_n26349_, new_n26350_, new_n26351_,
    new_n26352_, new_n26353_, new_n26354_, new_n26355_, new_n26356_,
    new_n26357_, new_n26358_, new_n26359_, new_n26360_, new_n26361_,
    new_n26362_, new_n26363_, new_n26364_, new_n26365_, new_n26366_,
    new_n26367_, new_n26368_, new_n26369_, new_n26370_, new_n26371_,
    new_n26373_, new_n26374_, new_n26375_, new_n26376_, new_n26377_,
    new_n26378_, new_n26379_, new_n26380_, new_n26381_, new_n26382_,
    new_n26383_, new_n26384_, new_n26385_, new_n26386_, new_n26388_,
    new_n26389_, new_n26390_, new_n26391_, new_n26393_, new_n26394_,
    new_n26395_, new_n26396_, new_n26397_, new_n26398_, new_n26399_,
    new_n26400_, new_n26401_, new_n26402_, new_n26403_, new_n26404_,
    new_n26405_, new_n26407_, new_n26408_, new_n26409_, new_n26410_,
    new_n26412_, new_n26413_, new_n26414_, new_n26415_, new_n26416_,
    new_n26417_, new_n26418_, new_n26419_, new_n26420_, new_n26421_,
    new_n26422_, new_n26423_, new_n26424_, new_n26425_, new_n26426_,
    new_n26427_, new_n26428_, new_n26429_, new_n26430_, new_n26431_,
    new_n26432_, new_n26433_, new_n26434_, new_n26435_, new_n26436_,
    new_n26437_, new_n26438_, new_n26439_, new_n26440_, new_n26441_,
    new_n26442_, new_n26443_, new_n26444_, new_n26445_, new_n26446_,
    new_n26447_, new_n26448_, new_n26449_, new_n26450_, new_n26451_,
    new_n26452_, new_n26453_, new_n26454_, new_n26455_, new_n26456_,
    new_n26457_, new_n26458_, new_n26459_, new_n26460_, new_n26461_,
    new_n26462_, new_n26463_, new_n26464_, new_n26465_, new_n26466_,
    new_n26467_, new_n26468_, new_n26469_, new_n26470_, new_n26471_,
    new_n26472_, new_n26473_, new_n26474_, new_n26475_, new_n26476_,
    new_n26477_, new_n26478_, new_n26479_, new_n26480_, new_n26481_,
    new_n26482_, new_n26483_, new_n26484_, new_n26486_, new_n26487_,
    new_n26488_, new_n26489_, new_n26490_, new_n26491_, new_n26492_,
    new_n26493_, new_n26494_, new_n26495_, new_n26496_, new_n26497_,
    new_n26498_, new_n26499_, new_n26500_, new_n26501_, new_n26502_,
    new_n26503_, new_n26504_, new_n26505_, new_n26506_, new_n26507_,
    new_n26508_, new_n26509_, new_n26510_, new_n26511_, new_n26512_,
    new_n26513_, new_n26514_, new_n26515_, new_n26516_, new_n26517_,
    new_n26518_, new_n26519_, new_n26520_, new_n26521_, new_n26522_,
    new_n26523_, new_n26524_, new_n26525_, new_n26526_, new_n26527_,
    new_n26528_, new_n26529_, new_n26530_, new_n26531_, new_n26532_,
    new_n26533_, new_n26534_, new_n26535_, new_n26536_, new_n26537_,
    new_n26538_, new_n26539_, new_n26540_, new_n26541_, new_n26542_,
    new_n26543_, new_n26544_, new_n26545_, new_n26546_, new_n26547_,
    new_n26548_, new_n26549_, new_n26550_, new_n26551_, new_n26552_,
    new_n26553_, new_n26554_, new_n26555_, new_n26556_, new_n26557_,
    new_n26558_, new_n26559_, new_n26560_, new_n26561_, new_n26562_,
    new_n26563_, new_n26564_, new_n26565_, new_n26566_, new_n26567_,
    new_n26568_, new_n26569_, new_n26570_, new_n26571_, new_n26572_,
    new_n26573_, new_n26574_, new_n26575_, new_n26576_, new_n26577_,
    new_n26578_, new_n26579_, new_n26580_, new_n26581_, new_n26582_,
    new_n26583_, new_n26584_, new_n26585_, new_n26586_, new_n26587_,
    new_n26588_, new_n26589_, new_n26590_, new_n26591_, new_n26592_,
    new_n26593_, new_n26594_, new_n26595_, new_n26596_, new_n26597_,
    new_n26598_, new_n26599_, new_n26600_, new_n26601_, new_n26602_,
    new_n26603_, new_n26604_, new_n26605_, new_n26606_, new_n26607_,
    new_n26608_, new_n26609_, new_n26610_, new_n26611_, new_n26612_,
    new_n26613_, new_n26614_, new_n26615_, new_n26616_, new_n26617_,
    new_n26618_, new_n26619_, new_n26620_, new_n26621_, new_n26622_,
    new_n26623_, new_n26624_, new_n26625_, new_n26626_, new_n26627_,
    new_n26628_, new_n26629_, new_n26630_, new_n26631_, new_n26632_,
    new_n26633_, new_n26634_, new_n26635_, new_n26636_, new_n26637_,
    new_n26638_, new_n26639_, new_n26640_, new_n26641_, new_n26642_,
    new_n26643_, new_n26644_, new_n26645_, new_n26646_, new_n26647_,
    new_n26648_, new_n26649_, new_n26650_, new_n26651_, new_n26652_,
    new_n26653_, new_n26654_, new_n26655_, new_n26656_, new_n26657_,
    new_n26658_, new_n26659_, new_n26660_, new_n26661_, new_n26662_,
    new_n26663_, new_n26664_, new_n26665_, new_n26666_, new_n26667_,
    new_n26668_, new_n26669_, new_n26670_, new_n26671_, new_n26672_,
    new_n26673_, new_n26674_, new_n26675_, new_n26676_, new_n26677_,
    new_n26678_, new_n26679_, new_n26680_, new_n26681_, new_n26682_,
    new_n26683_, new_n26684_, new_n26685_, new_n26686_, new_n26687_,
    new_n26688_, new_n26689_, new_n26690_, new_n26691_, new_n26692_,
    new_n26693_, new_n26694_, new_n26695_, new_n26696_, new_n26697_,
    new_n26698_, new_n26699_, new_n26700_, new_n26701_, new_n26702_,
    new_n26703_, new_n26704_, new_n26705_, new_n26706_, new_n26707_,
    new_n26708_, new_n26709_, new_n26710_, new_n26711_, new_n26712_,
    new_n26713_, new_n26714_, new_n26715_, new_n26716_, new_n26717_,
    new_n26718_, new_n26719_, new_n26720_, new_n26721_, new_n26722_,
    new_n26723_, new_n26724_, new_n26725_, new_n26726_, new_n26727_,
    new_n26728_, new_n26729_, new_n26730_, new_n26731_, new_n26732_,
    new_n26733_, new_n26734_, new_n26735_, new_n26736_, new_n26737_,
    new_n26738_, new_n26739_, new_n26740_, new_n26741_, new_n26742_,
    new_n26743_, new_n26744_, new_n26745_, new_n26746_, new_n26747_,
    new_n26748_, new_n26749_, new_n26750_, new_n26751_, new_n26752_,
    new_n26753_, new_n26754_, new_n26755_, new_n26756_, new_n26757_,
    new_n26758_, new_n26759_, new_n26760_, new_n26761_, new_n26762_,
    new_n26763_, new_n26764_, new_n26765_, new_n26766_, new_n26767_,
    new_n26768_, new_n26769_, new_n26770_, new_n26771_, new_n26772_,
    new_n26773_, new_n26774_, new_n26775_, new_n26776_, new_n26777_,
    new_n26778_, new_n26779_, new_n26780_, new_n26781_, new_n26782_,
    new_n26783_, new_n26784_, new_n26785_, new_n26786_, new_n26787_,
    new_n26788_, new_n26789_, new_n26790_, new_n26791_, new_n26792_,
    new_n26793_, new_n26794_, new_n26795_, new_n26796_, new_n26797_,
    new_n26798_, new_n26799_, new_n26800_, new_n26801_, new_n26802_,
    new_n26803_, new_n26804_, new_n26805_, new_n26806_, new_n26807_,
    new_n26808_, new_n26809_, new_n26810_, new_n26811_, new_n26812_,
    new_n26813_, new_n26814_, new_n26815_, new_n26816_, new_n26817_,
    new_n26818_, new_n26819_, new_n26820_, new_n26821_, new_n26822_,
    new_n26823_, new_n26824_, new_n26825_, new_n26826_, new_n26827_,
    new_n26828_, new_n26829_, new_n26830_, new_n26831_, new_n26832_,
    new_n26833_, new_n26834_, new_n26835_, new_n26836_, new_n26837_,
    new_n26838_, new_n26839_, new_n26840_, new_n26841_, new_n26842_,
    new_n26843_, new_n26844_, new_n26845_, new_n26846_, new_n26847_,
    new_n26848_, new_n26849_, new_n26850_, new_n26851_, new_n26852_,
    new_n26853_, new_n26854_, new_n26855_, new_n26856_, new_n26857_,
    new_n26858_, new_n26859_, new_n26860_, new_n26861_, new_n26862_,
    new_n26863_, new_n26864_, new_n26865_, new_n26866_, new_n26867_,
    new_n26868_, new_n26869_, new_n26870_, new_n26871_, new_n26872_,
    new_n26873_, new_n26874_, new_n26875_, new_n26876_, new_n26877_,
    new_n26878_, new_n26879_, new_n26880_, new_n26881_, new_n26882_,
    new_n26883_, new_n26884_, new_n26885_, new_n26886_, new_n26887_,
    new_n26888_, new_n26889_, new_n26890_, new_n26891_, new_n26892_,
    new_n26893_, new_n26894_, new_n26895_, new_n26896_, new_n26897_,
    new_n26898_, new_n26899_, new_n26900_, new_n26901_, new_n26902_,
    new_n26903_, new_n26904_, new_n26905_, new_n26906_, new_n26907_,
    new_n26908_, new_n26909_, new_n26910_, new_n26911_, new_n26912_,
    new_n26913_, new_n26914_, new_n26915_, new_n26916_, new_n26917_,
    new_n26918_, new_n26919_, new_n26920_, new_n26921_, new_n26922_,
    new_n26923_, new_n26924_, new_n26925_, new_n26926_, new_n26928_,
    new_n26929_, new_n26930_, new_n26931_, new_n26932_, new_n26933_,
    new_n26934_, new_n26935_, new_n26936_, new_n26937_, new_n26938_,
    new_n26939_, new_n26940_, new_n26941_, new_n26942_, new_n26943_,
    new_n26944_, new_n26945_, new_n26946_, new_n26947_, new_n26948_,
    new_n26949_, new_n26950_, new_n26951_, new_n26952_, new_n26953_,
    new_n26954_, new_n26955_, new_n26956_, new_n26957_, new_n26958_,
    new_n26959_, new_n26960_, new_n26961_, new_n26962_, new_n26963_,
    new_n26964_, new_n26965_, new_n26966_, new_n26967_, new_n26968_,
    new_n26969_, new_n26970_, new_n26971_, new_n26972_, new_n26973_,
    new_n26974_, new_n26975_, new_n26976_, new_n26977_, new_n26978_,
    new_n26979_, new_n26980_, new_n26981_, new_n26982_, new_n26983_,
    new_n26984_, new_n26985_, new_n26986_, new_n26987_, new_n26988_,
    new_n26989_, new_n26990_, new_n26991_, new_n26992_, new_n26993_,
    new_n26994_, new_n26995_, new_n26996_, new_n26997_, new_n26998_,
    new_n26999_, new_n27000_, new_n27001_, new_n27002_, new_n27003_,
    new_n27004_, new_n27005_, new_n27006_, new_n27007_, new_n27008_,
    new_n27009_, new_n27010_, new_n27011_, new_n27012_, new_n27013_,
    new_n27014_, new_n27015_, new_n27016_, new_n27017_, new_n27018_,
    new_n27019_, new_n27020_, new_n27021_, new_n27022_, new_n27023_,
    new_n27024_, new_n27025_, new_n27026_, new_n27027_, new_n27028_,
    new_n27029_, new_n27030_, new_n27031_, new_n27032_, new_n27033_,
    new_n27034_, new_n27035_, new_n27036_, new_n27037_, new_n27038_,
    new_n27039_, new_n27040_, new_n27041_, new_n27042_, new_n27043_,
    new_n27044_, new_n27045_, new_n27046_, new_n27047_, new_n27048_,
    new_n27049_, new_n27050_, new_n27051_, new_n27052_, new_n27053_,
    new_n27054_, new_n27055_, new_n27056_, new_n27057_, new_n27058_,
    new_n27059_, new_n27060_, new_n27061_, new_n27062_, new_n27063_,
    new_n27064_, new_n27065_, new_n27066_, new_n27067_, new_n27068_,
    new_n27069_, new_n27070_, new_n27071_, new_n27072_, new_n27073_,
    new_n27074_, new_n27075_, new_n27076_, new_n27077_, new_n27078_,
    new_n27079_, new_n27080_, new_n27081_, new_n27082_, new_n27083_,
    new_n27084_, new_n27085_, new_n27086_, new_n27087_, new_n27088_,
    new_n27089_, new_n27090_, new_n27091_, new_n27092_, new_n27093_,
    new_n27094_, new_n27095_, new_n27096_, new_n27097_, new_n27098_,
    new_n27099_, new_n27100_, new_n27101_, new_n27102_, new_n27103_,
    new_n27104_, new_n27105_, new_n27106_, new_n27107_, new_n27108_,
    new_n27109_, new_n27110_, new_n27111_, new_n27112_, new_n27113_,
    new_n27114_, new_n27115_, new_n27116_, new_n27117_, new_n27118_,
    new_n27119_, new_n27120_, new_n27121_, new_n27122_, new_n27123_,
    new_n27124_, new_n27125_, new_n27126_, new_n27127_, new_n27128_,
    new_n27129_, new_n27130_, new_n27131_, new_n27132_, new_n27133_,
    new_n27134_, new_n27135_, new_n27136_, new_n27137_, new_n27138_,
    new_n27139_, new_n27140_, new_n27141_, new_n27142_, new_n27143_,
    new_n27144_, new_n27145_, new_n27146_, new_n27147_, new_n27148_,
    new_n27149_, new_n27150_, new_n27151_, new_n27152_, new_n27153_,
    new_n27154_, new_n27155_, new_n27156_, new_n27157_, new_n27158_,
    new_n27159_, new_n27160_, new_n27161_, new_n27162_, new_n27163_,
    new_n27164_, new_n27165_, new_n27166_, new_n27167_, new_n27168_,
    new_n27169_, new_n27170_, new_n27171_, new_n27172_, new_n27173_,
    new_n27174_, new_n27175_, new_n27176_, new_n27177_, new_n27178_,
    new_n27179_, new_n27180_, new_n27181_, new_n27182_, new_n27183_,
    new_n27184_, new_n27185_, new_n27186_, new_n27187_, new_n27188_,
    new_n27189_, new_n27190_, new_n27191_, new_n27192_, new_n27193_,
    new_n27194_, new_n27195_, new_n27196_, new_n27197_, new_n27198_,
    new_n27199_, new_n27200_, new_n27201_, new_n27202_, new_n27203_,
    new_n27204_, new_n27205_, new_n27206_, new_n27207_, new_n27208_,
    new_n27209_, new_n27210_, new_n27211_, new_n27212_, new_n27213_,
    new_n27214_, new_n27215_, new_n27216_, new_n27217_, new_n27218_,
    new_n27219_, new_n27220_, new_n27221_, new_n27222_, new_n27223_,
    new_n27224_, new_n27225_, new_n27226_, new_n27227_, new_n27228_,
    new_n27229_, new_n27230_, new_n27231_, new_n27232_, new_n27233_,
    new_n27234_, new_n27235_, new_n27236_, new_n27237_, new_n27238_,
    new_n27239_, new_n27240_, new_n27241_, new_n27242_, new_n27243_,
    new_n27244_, new_n27245_, new_n27246_, new_n27247_, new_n27248_,
    new_n27249_, new_n27250_, new_n27251_, new_n27252_, new_n27253_,
    new_n27254_, new_n27255_, new_n27256_, new_n27257_, new_n27258_,
    new_n27259_, new_n27260_, new_n27261_, new_n27262_, new_n27263_,
    new_n27264_, new_n27265_, new_n27266_, new_n27267_, new_n27268_,
    new_n27269_, new_n27270_, new_n27271_, new_n27272_, new_n27273_,
    new_n27274_, new_n27275_, new_n27276_, new_n27277_, new_n27278_,
    new_n27279_, new_n27280_, new_n27281_, new_n27282_, new_n27283_,
    new_n27284_, new_n27285_, new_n27286_, new_n27287_, new_n27288_,
    new_n27289_, new_n27290_, new_n27291_, new_n27292_, new_n27293_,
    new_n27294_, new_n27295_, new_n27296_, new_n27297_, new_n27298_,
    new_n27299_, new_n27300_, new_n27301_, new_n27302_, new_n27303_,
    new_n27304_, new_n27305_, new_n27306_, new_n27307_, new_n27308_,
    new_n27309_, new_n27310_, new_n27311_, new_n27312_, new_n27313_,
    new_n27314_, new_n27315_, new_n27316_, new_n27317_, new_n27318_,
    new_n27319_, new_n27320_, new_n27321_, new_n27322_, new_n27323_,
    new_n27324_, new_n27325_, new_n27326_, new_n27327_, new_n27328_,
    new_n27329_, new_n27330_, new_n27331_, new_n27332_, new_n27333_,
    new_n27334_, new_n27335_, new_n27336_, new_n27337_, new_n27338_,
    new_n27339_, new_n27340_, new_n27341_, new_n27342_, new_n27343_,
    new_n27344_, new_n27345_, new_n27346_, new_n27347_, new_n27348_,
    new_n27349_, new_n27350_, new_n27351_, new_n27352_, new_n27353_,
    new_n27355_, new_n27356_, new_n27357_, new_n27358_, new_n27359_,
    new_n27360_, new_n27361_, new_n27362_, new_n27363_, new_n27364_,
    new_n27365_, new_n27366_, new_n27367_, new_n27368_, new_n27369_,
    new_n27370_, new_n27371_, new_n27372_, new_n27373_, new_n27374_,
    new_n27375_, new_n27376_, new_n27377_, new_n27378_, new_n27379_,
    new_n27380_, new_n27381_, new_n27382_, new_n27383_, new_n27384_,
    new_n27385_, new_n27386_, new_n27387_, new_n27388_, new_n27389_,
    new_n27390_, new_n27391_, new_n27392_, new_n27393_, new_n27394_,
    new_n27395_, new_n27396_, new_n27397_, new_n27398_, new_n27399_,
    new_n27400_, new_n27401_, new_n27402_, new_n27403_, new_n27404_,
    new_n27405_, new_n27406_, new_n27407_, new_n27408_, new_n27409_,
    new_n27410_, new_n27411_, new_n27412_, new_n27413_, new_n27414_,
    new_n27415_, new_n27416_, new_n27417_, new_n27418_, new_n27419_,
    new_n27420_, new_n27421_, new_n27422_, new_n27423_, new_n27424_,
    new_n27425_, new_n27426_, new_n27427_, new_n27428_, new_n27429_,
    new_n27430_, new_n27431_, new_n27432_, new_n27433_, new_n27434_,
    new_n27435_, new_n27436_, new_n27437_, new_n27438_, new_n27439_,
    new_n27440_, new_n27441_, new_n27442_, new_n27443_, new_n27444_,
    new_n27445_, new_n27446_, new_n27447_, new_n27448_, new_n27449_,
    new_n27450_, new_n27451_, new_n27452_, new_n27453_, new_n27454_,
    new_n27455_, new_n27456_, new_n27457_, new_n27458_, new_n27459_,
    new_n27460_, new_n27461_, new_n27462_, new_n27463_, new_n27464_,
    new_n27465_, new_n27466_, new_n27467_, new_n27468_, new_n27469_,
    new_n27470_, new_n27471_, new_n27472_, new_n27473_, new_n27474_,
    new_n27475_, new_n27476_, new_n27477_, new_n27478_, new_n27479_,
    new_n27480_, new_n27481_, new_n27482_, new_n27483_, new_n27484_,
    new_n27485_, new_n27486_, new_n27487_, new_n27488_, new_n27489_,
    new_n27490_, new_n27491_, new_n27492_, new_n27493_, new_n27494_,
    new_n27495_, new_n27496_, new_n27497_, new_n27498_, new_n27499_,
    new_n27500_, new_n27501_, new_n27502_, new_n27503_, new_n27504_,
    new_n27505_, new_n27506_, new_n27507_, new_n27508_, new_n27509_,
    new_n27510_, new_n27511_, new_n27512_, new_n27513_, new_n27514_,
    new_n27515_, new_n27516_, new_n27517_, new_n27518_, new_n27519_,
    new_n27520_, new_n27521_, new_n27522_, new_n27523_, new_n27524_,
    new_n27525_, new_n27526_, new_n27527_, new_n27528_, new_n27529_,
    new_n27530_, new_n27531_, new_n27532_, new_n27533_, new_n27534_,
    new_n27535_, new_n27536_, new_n27537_, new_n27538_, new_n27539_,
    new_n27540_, new_n27541_, new_n27542_, new_n27543_, new_n27544_,
    new_n27545_, new_n27546_, new_n27547_, new_n27548_, new_n27549_,
    new_n27550_, new_n27551_, new_n27552_, new_n27553_, new_n27554_,
    new_n27555_, new_n27556_, new_n27557_, new_n27558_, new_n27559_,
    new_n27560_, new_n27561_, new_n27562_, new_n27563_, new_n27564_,
    new_n27565_, new_n27566_, new_n27567_, new_n27568_, new_n27569_,
    new_n27570_, new_n27571_, new_n27572_, new_n27573_, new_n27574_,
    new_n27575_, new_n27576_, new_n27577_, new_n27578_, new_n27579_,
    new_n27580_, new_n27581_, new_n27582_, new_n27583_, new_n27584_,
    new_n27585_, new_n27586_, new_n27587_, new_n27588_, new_n27589_,
    new_n27590_, new_n27591_, new_n27592_, new_n27593_, new_n27594_,
    new_n27595_, new_n27596_, new_n27597_, new_n27598_, new_n27599_,
    new_n27600_, new_n27601_, new_n27602_, new_n27603_, new_n27604_,
    new_n27605_, new_n27606_, new_n27607_, new_n27608_, new_n27609_,
    new_n27610_, new_n27611_, new_n27612_, new_n27613_, new_n27614_,
    new_n27615_, new_n27616_, new_n27617_, new_n27618_, new_n27619_,
    new_n27620_, new_n27621_, new_n27622_, new_n27623_, new_n27624_,
    new_n27625_, new_n27626_, new_n27627_, new_n27628_, new_n27629_,
    new_n27630_, new_n27631_, new_n27632_, new_n27633_, new_n27634_,
    new_n27635_, new_n27636_, new_n27637_, new_n27638_, new_n27639_,
    new_n27640_, new_n27641_, new_n27642_, new_n27643_, new_n27644_,
    new_n27645_, new_n27646_, new_n27647_, new_n27648_, new_n27649_,
    new_n27650_, new_n27651_, new_n27652_, new_n27653_, new_n27654_,
    new_n27655_, new_n27656_, new_n27657_, new_n27658_, new_n27659_,
    new_n27660_, new_n27661_, new_n27662_, new_n27663_, new_n27664_,
    new_n27665_, new_n27666_, new_n27667_, new_n27668_, new_n27669_,
    new_n27670_, new_n27671_, new_n27672_, new_n27673_, new_n27674_,
    new_n27675_, new_n27676_, new_n27677_, new_n27678_, new_n27679_,
    new_n27680_, new_n27681_, new_n27682_, new_n27683_, new_n27684_,
    new_n27685_, new_n27686_, new_n27687_, new_n27688_, new_n27689_,
    new_n27690_, new_n27691_, new_n27692_, new_n27693_, new_n27694_,
    new_n27695_, new_n27696_, new_n27697_, new_n27698_, new_n27699_,
    new_n27700_, new_n27701_, new_n27702_, new_n27703_, new_n27704_,
    new_n27705_, new_n27706_, new_n27707_, new_n27708_, new_n27709_,
    new_n27710_, new_n27711_, new_n27712_, new_n27713_, new_n27714_,
    new_n27715_, new_n27716_, new_n27717_, new_n27718_, new_n27719_,
    new_n27720_, new_n27721_, new_n27722_, new_n27723_, new_n27724_,
    new_n27725_, new_n27726_, new_n27727_, new_n27728_, new_n27729_,
    new_n27730_, new_n27731_, new_n27732_, new_n27733_, new_n27734_,
    new_n27735_, new_n27736_, new_n27737_, new_n27738_, new_n27739_,
    new_n27740_, new_n27741_, new_n27742_, new_n27743_, new_n27744_,
    new_n27745_, new_n27746_, new_n27747_, new_n27748_, new_n27749_,
    new_n27750_, new_n27751_, new_n27752_, new_n27753_, new_n27754_,
    new_n27755_, new_n27756_, new_n27757_, new_n27758_, new_n27759_,
    new_n27760_, new_n27761_, new_n27762_, new_n27763_, new_n27764_,
    new_n27765_, new_n27766_, new_n27768_, new_n27769_, new_n27770_,
    new_n27771_, new_n27772_, new_n27773_, new_n27774_, new_n27775_,
    new_n27776_, new_n27777_, new_n27778_, new_n27779_, new_n27780_,
    new_n27781_, new_n27782_, new_n27783_, new_n27784_, new_n27785_,
    new_n27786_, new_n27787_, new_n27788_, new_n27789_, new_n27790_,
    new_n27791_, new_n27792_, new_n27793_, new_n27794_, new_n27795_,
    new_n27796_, new_n27797_, new_n27798_, new_n27799_, new_n27800_,
    new_n27801_, new_n27802_, new_n27803_, new_n27804_, new_n27805_,
    new_n27806_, new_n27807_, new_n27808_, new_n27809_, new_n27810_,
    new_n27811_, new_n27812_, new_n27813_, new_n27814_, new_n27815_,
    new_n27816_, new_n27817_, new_n27818_, new_n27819_, new_n27820_,
    new_n27821_, new_n27822_, new_n27823_, new_n27824_, new_n27825_,
    new_n27826_, new_n27827_, new_n27828_, new_n27829_, new_n27830_,
    new_n27831_, new_n27832_, new_n27833_, new_n27834_, new_n27835_,
    new_n27836_, new_n27837_, new_n27838_, new_n27839_, new_n27840_,
    new_n27841_, new_n27842_, new_n27843_, new_n27844_, new_n27845_,
    new_n27847_, new_n27848_, new_n27849_, new_n27850_, new_n27851_,
    new_n27852_, new_n27853_, new_n27854_, new_n27855_, new_n27856_,
    new_n27857_, new_n27858_, new_n27859_, new_n27860_, new_n27861_,
    new_n27862_, new_n27863_, new_n27864_, new_n27865_, new_n27866_,
    new_n27867_, new_n27868_, new_n27869_, new_n27870_, new_n27871_,
    new_n27872_, new_n27873_, new_n27874_, new_n27875_, new_n27876_,
    new_n27877_, new_n27879_, new_n27880_, new_n27881_, new_n27882_,
    new_n27883_, new_n27884_, new_n27885_, new_n27886_, new_n27887_,
    new_n27888_, new_n27889_, new_n27890_, new_n27891_, new_n27892_,
    new_n27893_, new_n27894_, new_n27895_, new_n27896_, new_n27897_,
    new_n27898_, new_n27899_, new_n27901_, new_n27902_, new_n27903_,
    new_n27904_, new_n27905_, new_n27906_, new_n27908_, new_n27909_,
    new_n27910_, new_n27911_, new_n27912_, new_n27913_, new_n27914_,
    new_n27915_, new_n27916_, new_n27917_, new_n27918_, new_n27919_,
    new_n27920_, new_n27921_, new_n27922_, new_n27923_, new_n27924_,
    new_n27925_, new_n27926_, new_n27927_, new_n27928_, new_n27929_,
    new_n27930_, new_n27931_, new_n27932_, new_n27933_, new_n27934_,
    new_n27935_, new_n27936_, new_n27937_, new_n27938_, new_n27939_,
    new_n27940_, new_n27941_, new_n27942_, new_n27943_, new_n27944_,
    new_n27945_, new_n27946_, new_n27947_, new_n27948_, new_n27949_,
    new_n27950_, new_n27951_, new_n27952_, new_n27953_, new_n27954_,
    new_n27955_, new_n27956_, new_n27957_, new_n27958_, new_n27959_,
    new_n27960_, new_n27961_, new_n27962_, new_n27964_, new_n27965_,
    new_n27966_, new_n27967_, new_n27968_, new_n27969_, new_n27970_,
    new_n27971_, new_n27972_, new_n27973_, new_n27974_, new_n27975_,
    new_n27976_, new_n27977_, new_n27978_, new_n27979_, new_n27980_,
    new_n27981_, new_n27982_, new_n27983_, new_n27984_, new_n27985_,
    new_n27986_, new_n27987_, new_n27988_, new_n27989_, new_n27990_,
    new_n27991_, new_n27992_, new_n27993_, new_n27994_, new_n27995_,
    new_n27996_, new_n27997_, new_n27999_, new_n28000_, new_n28001_,
    new_n28002_, new_n28003_, new_n28004_, new_n28005_, new_n28006_,
    new_n28007_, new_n28008_, new_n28009_, new_n28010_, new_n28011_,
    new_n28012_, new_n28013_, new_n28014_, new_n28015_, new_n28016_,
    new_n28017_, new_n28018_, new_n28019_, new_n28020_, new_n28021_,
    new_n28022_, new_n28023_, new_n28024_, new_n28025_, new_n28026_,
    new_n28027_, new_n28028_, new_n28029_, new_n28030_, new_n28031_,
    new_n28032_, new_n28033_, new_n28034_, new_n28035_, new_n28036_,
    new_n28037_, new_n28038_, new_n28039_, new_n28040_, new_n28041_,
    new_n28042_, new_n28043_, new_n28044_, new_n28045_, new_n28046_,
    new_n28047_, new_n28048_, new_n28049_, new_n28050_, new_n28051_,
    new_n28052_, new_n28053_, new_n28054_, new_n28055_, new_n28056_,
    new_n28057_, new_n28058_, new_n28059_, new_n28060_, new_n28061_,
    new_n28062_, new_n28063_, new_n28064_, new_n28065_, new_n28066_,
    new_n28067_, new_n28068_, new_n28069_, new_n28070_, new_n28071_,
    new_n28072_, new_n28073_, new_n28074_, new_n28075_, new_n28076_,
    new_n28077_, new_n28078_, new_n28079_, new_n28080_, new_n28081_,
    new_n28082_, new_n28083_, new_n28084_, new_n28085_, new_n28086_,
    new_n28087_, new_n28088_, new_n28089_, new_n28090_, new_n28091_,
    new_n28092_, new_n28093_, new_n28094_, new_n28095_, new_n28096_,
    new_n28097_, new_n28098_, new_n28099_, new_n28100_, new_n28101_,
    new_n28102_, new_n28103_, new_n28104_, new_n28105_, new_n28106_,
    new_n28107_, new_n28108_, new_n28109_, new_n28110_, new_n28111_,
    new_n28112_, new_n28113_, new_n28114_, new_n28115_, new_n28116_,
    new_n28117_, new_n28118_, new_n28119_, new_n28120_, new_n28121_,
    new_n28122_, new_n28123_, new_n28124_, new_n28125_, new_n28126_,
    new_n28127_, new_n28128_, new_n28129_, new_n28130_, new_n28131_,
    new_n28132_, new_n28133_, new_n28134_, new_n28135_, new_n28136_,
    new_n28137_, new_n28138_, new_n28139_, new_n28140_, new_n28141_,
    new_n28142_, new_n28143_, new_n28144_, new_n28145_, new_n28146_,
    new_n28147_, new_n28148_, new_n28149_, new_n28150_, new_n28151_,
    new_n28152_, new_n28153_, new_n28154_, new_n28155_, new_n28156_,
    new_n28157_, new_n28158_, new_n28159_, new_n28160_, new_n28161_,
    new_n28162_, new_n28163_, new_n28164_, new_n28165_, new_n28166_,
    new_n28167_, new_n28168_, new_n28169_, new_n28170_, new_n28171_,
    new_n28172_, new_n28173_, new_n28174_, new_n28175_, new_n28176_,
    new_n28177_, new_n28178_, new_n28179_, new_n28180_, new_n28181_,
    new_n28182_, new_n28183_, new_n28184_, new_n28185_, new_n28186_,
    new_n28187_, new_n28188_, new_n28189_, new_n28190_, new_n28191_,
    new_n28192_, new_n28193_, new_n28194_, new_n28195_, new_n28196_,
    new_n28197_, new_n28198_, new_n28199_, new_n28200_, new_n28201_,
    new_n28202_, new_n28203_, new_n28204_, new_n28205_, new_n28206_,
    new_n28207_, new_n28208_, new_n28209_, new_n28210_, new_n28211_,
    new_n28212_, new_n28213_, new_n28214_, new_n28215_, new_n28216_,
    new_n28217_, new_n28218_, new_n28219_, new_n28220_, new_n28221_,
    new_n28222_, new_n28223_, new_n28224_, new_n28225_, new_n28226_,
    new_n28227_, new_n28228_, new_n28229_, new_n28230_, new_n28231_,
    new_n28232_, new_n28233_, new_n28234_, new_n28235_, new_n28236_,
    new_n28237_, new_n28238_, new_n28239_, new_n28240_, new_n28241_,
    new_n28242_, new_n28243_, new_n28244_, new_n28245_, new_n28246_,
    new_n28247_, new_n28248_, new_n28249_, new_n28250_, new_n28251_,
    new_n28252_, new_n28253_, new_n28254_, new_n28255_, new_n28256_,
    new_n28257_, new_n28258_, new_n28259_, new_n28260_, new_n28261_,
    new_n28262_, new_n28263_, new_n28264_, new_n28265_, new_n28266_,
    new_n28267_, new_n28268_, new_n28269_, new_n28270_, new_n28271_,
    new_n28272_, new_n28273_, new_n28274_, new_n28275_, new_n28276_,
    new_n28277_, new_n28278_, new_n28279_, new_n28280_, new_n28281_,
    new_n28282_, new_n28283_, new_n28284_, new_n28285_, new_n28286_,
    new_n28287_, new_n28288_, new_n28289_, new_n28290_, new_n28291_,
    new_n28292_, new_n28293_, new_n28294_, new_n28295_, new_n28296_,
    new_n28297_, new_n28298_, new_n28299_, new_n28300_, new_n28301_,
    new_n28302_, new_n28303_, new_n28304_, new_n28305_, new_n28306_,
    new_n28307_, new_n28308_, new_n28309_, new_n28310_, new_n28311_,
    new_n28312_, new_n28313_, new_n28314_, new_n28315_, new_n28316_,
    new_n28317_, new_n28318_, new_n28319_, new_n28320_, new_n28321_,
    new_n28322_, new_n28323_, new_n28324_, new_n28325_, new_n28326_,
    new_n28327_, new_n28328_, new_n28329_, new_n28330_, new_n28331_,
    new_n28332_, new_n28333_, new_n28334_, new_n28335_, new_n28336_,
    new_n28337_, new_n28338_, new_n28339_, new_n28340_, new_n28341_,
    new_n28342_, new_n28343_, new_n28344_, new_n28345_, new_n28346_,
    new_n28347_, new_n28348_, new_n28349_, new_n28350_, new_n28352_,
    new_n28353_, new_n28354_, new_n28355_, new_n28356_, new_n28357_,
    new_n28358_, new_n28359_, new_n28360_, new_n28361_, new_n28362_,
    new_n28363_, new_n28364_, new_n28365_, new_n28366_, new_n28367_,
    new_n28368_, new_n28369_, new_n28370_, new_n28371_, new_n28372_,
    new_n28373_, new_n28374_, new_n28375_, new_n28376_, new_n28377_,
    new_n28378_, new_n28379_, new_n28380_, new_n28381_, new_n28382_,
    new_n28383_, new_n28384_, new_n28385_, new_n28386_, new_n28387_,
    new_n28388_, new_n28389_, new_n28390_, new_n28391_, new_n28392_,
    new_n28393_, new_n28394_, new_n28395_, new_n28396_, new_n28397_,
    new_n28398_, new_n28399_, new_n28400_, new_n28401_, new_n28402_,
    new_n28403_, new_n28404_, new_n28405_, new_n28406_, new_n28407_,
    new_n28408_, new_n28409_, new_n28410_, new_n28411_, new_n28412_,
    new_n28413_, new_n28414_, new_n28415_, new_n28416_, new_n28417_,
    new_n28418_, new_n28419_, new_n28420_, new_n28421_, new_n28422_,
    new_n28423_, new_n28424_, new_n28425_, new_n28426_, new_n28427_,
    new_n28428_, new_n28429_, new_n28430_, new_n28431_, new_n28432_,
    new_n28433_, new_n28434_, new_n28435_, new_n28436_, new_n28437_,
    new_n28438_, new_n28439_, new_n28440_, new_n28441_, new_n28442_,
    new_n28443_, new_n28444_, new_n28445_, new_n28446_, new_n28447_,
    new_n28448_, new_n28449_, new_n28450_, new_n28451_, new_n28452_,
    new_n28453_, new_n28454_, new_n28455_, new_n28456_, new_n28457_,
    new_n28458_, new_n28459_, new_n28460_, new_n28461_, new_n28462_,
    new_n28463_, new_n28464_, new_n28465_, new_n28466_, new_n28467_,
    new_n28468_, new_n28469_, new_n28470_, new_n28471_, new_n28472_,
    new_n28473_, new_n28474_, new_n28475_, new_n28476_, new_n28477_,
    new_n28478_, new_n28479_, new_n28480_, new_n28481_, new_n28482_,
    new_n28483_, new_n28484_, new_n28485_, new_n28486_, new_n28487_,
    new_n28488_, new_n28489_, new_n28490_, new_n28491_, new_n28492_,
    new_n28493_, new_n28494_, new_n28495_, new_n28496_, new_n28497_,
    new_n28498_, new_n28499_, new_n28500_, new_n28501_, new_n28502_,
    new_n28503_, new_n28504_, new_n28505_, new_n28506_, new_n28507_,
    new_n28508_, new_n28509_, new_n28510_, new_n28511_, new_n28512_,
    new_n28513_, new_n28514_, new_n28515_, new_n28516_, new_n28517_,
    new_n28518_, new_n28519_, new_n28520_, new_n28521_, new_n28522_,
    new_n28523_, new_n28524_, new_n28525_, new_n28526_, new_n28527_,
    new_n28528_, new_n28529_, new_n28530_, new_n28531_, new_n28532_,
    new_n28533_, new_n28534_, new_n28535_, new_n28536_, new_n28537_,
    new_n28538_, new_n28539_, new_n28540_, new_n28541_, new_n28542_,
    new_n28543_, new_n28544_, new_n28545_, new_n28546_, new_n28547_,
    new_n28548_, new_n28549_, new_n28550_, new_n28551_, new_n28552_,
    new_n28553_, new_n28554_, new_n28555_, new_n28556_, new_n28557_,
    new_n28558_, new_n28559_, new_n28560_, new_n28561_, new_n28562_,
    new_n28563_, new_n28564_, new_n28565_, new_n28566_, new_n28567_,
    new_n28568_, new_n28569_, new_n28570_, new_n28571_, new_n28572_,
    new_n28573_, new_n28574_, new_n28575_, new_n28576_, new_n28577_,
    new_n28578_, new_n28579_, new_n28580_, new_n28581_, new_n28582_,
    new_n28583_, new_n28584_, new_n28585_, new_n28586_, new_n28587_,
    new_n28588_, new_n28589_, new_n28590_, new_n28591_, new_n28592_,
    new_n28593_, new_n28594_, new_n28595_, new_n28596_, new_n28597_,
    new_n28598_, new_n28599_, new_n28600_, new_n28601_, new_n28602_,
    new_n28603_, new_n28604_, new_n28605_, new_n28606_, new_n28607_,
    new_n28608_, new_n28609_, new_n28610_, new_n28611_, new_n28612_,
    new_n28613_, new_n28614_, new_n28615_, new_n28616_, new_n28617_,
    new_n28618_, new_n28620_, new_n28621_, new_n28622_, new_n28623_,
    new_n28624_, new_n28625_, new_n28626_, new_n28627_, new_n28628_,
    new_n28629_, new_n28630_, new_n28631_, new_n28632_, new_n28633_,
    new_n28634_, new_n28635_, new_n28636_, new_n28637_, new_n28638_,
    new_n28639_, new_n28640_, new_n28641_, new_n28642_, new_n28643_,
    new_n28644_, new_n28645_, new_n28646_, new_n28647_, new_n28648_,
    new_n28649_, new_n28650_, new_n28651_, new_n28652_, new_n28653_,
    new_n28654_, new_n28655_, new_n28656_, new_n28657_, new_n28658_,
    new_n28659_, new_n28660_, new_n28661_, new_n28662_, new_n28663_,
    new_n28664_, new_n28665_, new_n28666_, new_n28667_, new_n28668_,
    new_n28669_, new_n28670_, new_n28671_, new_n28672_, new_n28673_,
    new_n28674_, new_n28675_, new_n28676_, new_n28677_, new_n28678_,
    new_n28679_, new_n28680_, new_n28681_, new_n28682_, new_n28683_,
    new_n28684_, new_n28685_, new_n28686_, new_n28687_, new_n28688_,
    new_n28689_, new_n28690_, new_n28691_, new_n28692_, new_n28693_,
    new_n28694_, new_n28695_, new_n28696_, new_n28697_, new_n28698_,
    new_n28699_, new_n28700_, new_n28701_, new_n28702_, new_n28703_,
    new_n28704_, new_n28705_, new_n28706_, new_n28707_, new_n28708_,
    new_n28709_, new_n28710_, new_n28711_, new_n28712_, new_n28713_,
    new_n28714_, new_n28715_, new_n28716_, new_n28717_, new_n28718_,
    new_n28719_, new_n28720_, new_n28721_, new_n28722_, new_n28723_,
    new_n28724_, new_n28725_, new_n28726_, new_n28727_, new_n28728_,
    new_n28729_, new_n28730_, new_n28731_, new_n28732_, new_n28733_,
    new_n28734_, new_n28735_, new_n28736_, new_n28737_, new_n28738_,
    new_n28739_, new_n28740_, new_n28741_, new_n28742_, new_n28743_,
    new_n28744_, new_n28745_, new_n28746_, new_n28747_, new_n28748_,
    new_n28749_, new_n28750_, new_n28751_, new_n28752_, new_n28753_,
    new_n28754_, new_n28755_, new_n28756_, new_n28757_, new_n28758_,
    new_n28759_, new_n28760_, new_n28761_, new_n28762_, new_n28763_,
    new_n28764_, new_n28765_, new_n28766_, new_n28767_, new_n28768_,
    new_n28769_, new_n28770_, new_n28772_, new_n28773_, new_n28774_,
    new_n28775_, new_n28776_, new_n28777_, new_n28778_, new_n28779_,
    new_n28780_, new_n28782_, new_n28783_, new_n28784_, new_n28785_,
    new_n28786_, new_n28787_, new_n28788_, new_n28789_, new_n28790_,
    new_n28791_, new_n28792_, new_n28793_, new_n28794_, new_n28795_,
    new_n28796_, new_n28797_, new_n28798_, new_n28799_, new_n28800_,
    new_n28801_, new_n28802_, new_n28803_, new_n28804_, new_n28805_,
    new_n28806_, new_n28807_, new_n28808_, new_n28809_, new_n28810_,
    new_n28811_, new_n28812_, new_n28813_, new_n28814_, new_n28815_,
    new_n28816_, new_n28817_, new_n28818_, new_n28819_, new_n28820_,
    new_n28821_, new_n28822_, new_n28823_, new_n28824_, new_n28825_,
    new_n28826_, new_n28827_, new_n28828_, new_n28829_, new_n28830_,
    new_n28831_, new_n28832_, new_n28833_, new_n28834_, new_n28835_,
    new_n28836_, new_n28837_, new_n28838_, new_n28839_, new_n28840_,
    new_n28841_, new_n28842_, new_n28843_, new_n28844_, new_n28845_,
    new_n28846_, new_n28847_, new_n28848_, new_n28849_, new_n28850_,
    new_n28851_, new_n28852_, new_n28853_, new_n28854_, new_n28855_,
    new_n28856_, new_n28857_, new_n28858_, new_n28859_, new_n28860_,
    new_n28861_, new_n28862_, new_n28863_, new_n28864_, new_n28865_,
    new_n28866_, new_n28867_, new_n28868_, new_n28869_, new_n28870_,
    new_n28871_, new_n28872_, new_n28873_, new_n28874_, new_n28875_,
    new_n28876_, new_n28877_, new_n28878_, new_n28879_, new_n28880_,
    new_n28881_, new_n28882_, new_n28883_, new_n28884_, new_n28885_,
    new_n28886_, new_n28887_, new_n28888_, new_n28889_, new_n28890_,
    new_n28891_, new_n28892_, new_n28893_, new_n28894_, new_n28895_,
    new_n28896_, new_n28897_, new_n28898_, new_n28899_, new_n28900_,
    new_n28901_, new_n28902_, new_n28903_, new_n28904_, new_n28905_,
    new_n28906_, new_n28907_, new_n28908_, new_n28909_, new_n28910_,
    new_n28911_, new_n28912_, new_n28913_, new_n28914_, new_n28915_,
    new_n28916_, new_n28917_, new_n28918_, new_n28919_, new_n28920_,
    new_n28921_, new_n28922_, new_n28923_, new_n28924_, new_n28925_,
    new_n28926_, new_n28927_, new_n28928_, new_n28929_, new_n28930_,
    new_n28931_, new_n28932_, new_n28933_, new_n28934_, new_n28935_,
    new_n28936_, new_n28937_, new_n28938_, new_n28939_, new_n28940_,
    new_n28941_, new_n28942_, new_n28943_, new_n28944_, new_n28945_,
    new_n28946_, new_n28947_, new_n28948_, new_n28949_, new_n28950_,
    new_n28951_, new_n28952_, new_n28953_, new_n28954_, new_n28955_,
    new_n28956_, new_n28957_, new_n28958_, new_n28959_, new_n28960_,
    new_n28961_, new_n28962_, new_n28963_, new_n28964_, new_n28965_,
    new_n28966_, new_n28967_, new_n28969_, new_n28970_, new_n28971_,
    new_n28972_, new_n28973_, new_n28974_, new_n28975_, new_n28976_,
    new_n28977_, new_n28978_, new_n28979_, new_n28980_, new_n28981_,
    new_n28982_, new_n28983_, new_n28984_, new_n28985_, new_n28986_,
    new_n28987_, new_n28988_, new_n28989_, new_n28990_, new_n28991_,
    new_n28992_, new_n28993_, new_n28994_, new_n28995_, new_n28996_,
    new_n28997_, new_n28998_, new_n28999_, new_n29000_, new_n29001_,
    new_n29002_, new_n29003_, new_n29004_, new_n29005_, new_n29006_,
    new_n29007_, new_n29008_, new_n29009_, new_n29010_, new_n29011_,
    new_n29012_, new_n29013_, new_n29014_, new_n29015_, new_n29016_,
    new_n29017_, new_n29018_, new_n29019_, new_n29020_, new_n29021_,
    new_n29022_, new_n29023_, new_n29024_, new_n29025_, new_n29026_,
    new_n29027_, new_n29028_, new_n29029_, new_n29030_, new_n29031_,
    new_n29032_, new_n29033_, new_n29034_, new_n29035_, new_n29036_,
    new_n29037_, new_n29038_, new_n29039_, new_n29040_, new_n29041_,
    new_n29042_, new_n29043_, new_n29044_, new_n29045_, new_n29046_,
    new_n29047_, new_n29048_, new_n29049_, new_n29050_, new_n29051_,
    new_n29052_, new_n29053_, new_n29054_, new_n29055_, new_n29056_,
    new_n29057_, new_n29058_, new_n29059_, new_n29060_, new_n29061_,
    new_n29062_, new_n29063_, new_n29064_, new_n29065_, new_n29066_,
    new_n29067_, new_n29068_, new_n29069_, new_n29070_, new_n29071_,
    new_n29072_, new_n29073_, new_n29074_, new_n29075_, new_n29076_,
    new_n29077_, new_n29078_, new_n29079_, new_n29080_, new_n29081_,
    new_n29082_, new_n29083_, new_n29084_, new_n29085_, new_n29086_,
    new_n29087_, new_n29088_, new_n29089_, new_n29090_, new_n29091_,
    new_n29092_, new_n29093_, new_n29094_, new_n29095_, new_n29096_,
    new_n29097_, new_n29098_, new_n29099_, new_n29100_, new_n29101_,
    new_n29102_, new_n29103_, new_n29104_, new_n29105_, new_n29106_,
    new_n29107_, new_n29108_, new_n29109_, new_n29110_, new_n29111_,
    new_n29112_, new_n29113_, new_n29114_, new_n29115_, new_n29116_,
    new_n29117_, new_n29118_, new_n29119_, new_n29120_, new_n29121_,
    new_n29122_, new_n29123_, new_n29124_, new_n29125_, new_n29126_,
    new_n29127_, new_n29128_, new_n29129_, new_n29130_, new_n29131_,
    new_n29132_, new_n29133_, new_n29134_, new_n29135_, new_n29136_,
    new_n29137_, new_n29138_, new_n29139_, new_n29140_, new_n29141_,
    new_n29142_, new_n29143_, new_n29144_, new_n29145_, new_n29146_,
    new_n29147_, new_n29148_, new_n29149_, new_n29150_, new_n29151_,
    new_n29152_, new_n29153_, new_n29154_, new_n29155_, new_n29156_,
    new_n29157_, new_n29158_, new_n29159_, new_n29160_, new_n29161_,
    new_n29162_, new_n29163_, new_n29164_, new_n29165_, new_n29166_,
    new_n29167_, new_n29168_, new_n29169_, new_n29170_, new_n29171_,
    new_n29172_, new_n29173_, new_n29174_, new_n29175_, new_n29176_,
    new_n29177_, new_n29178_, new_n29179_, new_n29180_, new_n29181_,
    new_n29182_, new_n29183_, new_n29184_, new_n29185_, new_n29186_,
    new_n29187_, new_n29188_, new_n29189_, new_n29190_, new_n29191_,
    new_n29192_, new_n29193_, new_n29194_, new_n29195_, new_n29196_,
    new_n29197_, new_n29198_, new_n29199_, new_n29200_, new_n29201_,
    new_n29202_, new_n29203_, new_n29204_, new_n29205_, new_n29206_,
    new_n29207_, new_n29208_, new_n29209_, new_n29210_, new_n29211_,
    new_n29212_, new_n29213_, new_n29214_, new_n29215_, new_n29216_,
    new_n29217_, new_n29218_, new_n29219_, new_n29220_, new_n29221_,
    new_n29222_, new_n29223_, new_n29224_, new_n29225_, new_n29226_,
    new_n29227_, new_n29228_, new_n29229_, new_n29231_, new_n29232_,
    new_n29233_, new_n29234_, new_n29235_, new_n29236_, new_n29237_,
    new_n29238_, new_n29239_, new_n29240_, new_n29241_, new_n29242_,
    new_n29243_, new_n29244_, new_n29245_, new_n29246_, new_n29247_,
    new_n29248_, new_n29249_, new_n29250_, new_n29251_, new_n29252_,
    new_n29253_, new_n29254_, new_n29255_, new_n29256_, new_n29257_,
    new_n29258_, new_n29259_, new_n29260_, new_n29261_, new_n29262_,
    new_n29263_, new_n29264_, new_n29265_, new_n29266_, new_n29267_,
    new_n29268_, new_n29269_, new_n29270_, new_n29271_, new_n29272_,
    new_n29273_, new_n29274_, new_n29275_, new_n29276_, new_n29277_,
    new_n29278_, new_n29279_, new_n29280_, new_n29281_, new_n29282_,
    new_n29283_, new_n29284_, new_n29285_, new_n29286_, new_n29287_,
    new_n29288_, new_n29289_, new_n29290_, new_n29291_, new_n29292_,
    new_n29293_, new_n29294_, new_n29296_, new_n29297_, new_n29298_,
    new_n29299_, new_n29300_, new_n29301_, new_n29302_, new_n29303_,
    new_n29304_, new_n29305_, new_n29306_, new_n29307_, new_n29308_,
    new_n29309_, new_n29310_, new_n29311_, new_n29312_, new_n29313_,
    new_n29314_, new_n29315_, new_n29316_, new_n29317_, new_n29318_,
    new_n29319_, new_n29320_, new_n29321_, new_n29322_, new_n29323_,
    new_n29324_, new_n29325_, new_n29326_, new_n29327_, new_n29328_,
    new_n29329_, new_n29330_, new_n29331_, new_n29332_, new_n29333_,
    new_n29334_, new_n29335_, new_n29336_, new_n29337_, new_n29338_,
    new_n29339_, new_n29340_, new_n29341_, new_n29342_, new_n29343_,
    new_n29344_, new_n29345_, new_n29346_, new_n29347_, new_n29348_,
    new_n29349_, new_n29350_, new_n29351_, new_n29352_, new_n29353_,
    new_n29354_, new_n29355_, new_n29356_, new_n29357_, new_n29358_,
    new_n29359_, new_n29360_, new_n29361_, new_n29362_, new_n29363_,
    new_n29364_, new_n29365_, new_n29366_, new_n29367_, new_n29368_,
    new_n29369_, new_n29370_, new_n29371_, new_n29372_, new_n29373_,
    new_n29374_, new_n29375_, new_n29376_, new_n29377_, new_n29378_,
    new_n29379_, new_n29380_, new_n29381_, new_n29382_, new_n29383_,
    new_n29384_, new_n29385_, new_n29386_, new_n29387_, new_n29388_,
    new_n29389_, new_n29390_, new_n29391_, new_n29392_, new_n29393_,
    new_n29394_, new_n29395_, new_n29396_, new_n29397_, new_n29398_,
    new_n29399_, new_n29400_, new_n29401_, new_n29402_, new_n29403_,
    new_n29404_, new_n29405_, new_n29406_, new_n29407_, new_n29408_,
    new_n29409_, new_n29410_, new_n29411_, new_n29412_, new_n29413_,
    new_n29414_, new_n29415_, new_n29416_, new_n29417_, new_n29418_,
    new_n29419_, new_n29420_, new_n29421_, new_n29422_, new_n29423_,
    new_n29424_, new_n29425_, new_n29426_, new_n29427_, new_n29428_,
    new_n29429_, new_n29430_, new_n29431_, new_n29432_, new_n29433_,
    new_n29434_, new_n29435_, new_n29436_, new_n29437_, new_n29438_,
    new_n29439_, new_n29440_, new_n29441_, new_n29442_, new_n29443_,
    new_n29444_, new_n29445_, new_n29446_, new_n29447_, new_n29448_,
    new_n29449_, new_n29450_, new_n29451_, new_n29452_, new_n29453_,
    new_n29454_, new_n29455_, new_n29456_, new_n29457_, new_n29458_,
    new_n29459_, new_n29460_, new_n29461_, new_n29462_, new_n29463_,
    new_n29464_, new_n29465_, new_n29466_, new_n29467_, new_n29468_,
    new_n29469_, new_n29470_, new_n29471_, new_n29472_, new_n29473_,
    new_n29474_, new_n29475_, new_n29476_, new_n29477_, new_n29478_,
    new_n29479_, new_n29480_, new_n29481_, new_n29482_, new_n29483_,
    new_n29484_, new_n29485_, new_n29486_, new_n29487_, new_n29488_,
    new_n29489_, new_n29490_, new_n29491_, new_n29492_, new_n29493_,
    new_n29494_, new_n29495_, new_n29496_, new_n29497_, new_n29498_,
    new_n29499_, new_n29500_, new_n29501_, new_n29502_, new_n29503_,
    new_n29504_, new_n29505_, new_n29506_, new_n29507_, new_n29508_,
    new_n29509_, new_n29510_, new_n29511_, new_n29512_, new_n29513_,
    new_n29514_, new_n29515_, new_n29516_, new_n29517_, new_n29518_,
    new_n29519_, new_n29520_, new_n29521_, new_n29522_, new_n29523_,
    new_n29524_, new_n29525_, new_n29526_, new_n29527_, new_n29528_,
    new_n29529_, new_n29530_, new_n29531_, new_n29532_, new_n29533_,
    new_n29534_, new_n29535_, new_n29536_, new_n29537_, new_n29538_,
    new_n29539_, new_n29540_, new_n29541_, new_n29542_, new_n29543_,
    new_n29544_, new_n29545_, new_n29546_, new_n29547_, new_n29548_,
    new_n29549_, new_n29550_, new_n29551_, new_n29552_, new_n29553_,
    new_n29554_, new_n29555_, new_n29556_, new_n29557_, new_n29558_,
    new_n29559_, new_n29560_, new_n29561_, new_n29562_, new_n29563_,
    new_n29564_, new_n29565_, new_n29566_, new_n29567_, new_n29568_,
    new_n29569_, new_n29570_, new_n29571_, new_n29572_, new_n29573_,
    new_n29574_, new_n29575_, new_n29576_, new_n29577_, new_n29578_,
    new_n29579_, new_n29580_, new_n29581_, new_n29582_, new_n29583_,
    new_n29584_, new_n29585_, new_n29586_, new_n29587_, new_n29588_,
    new_n29589_, new_n29590_, new_n29591_, new_n29592_, new_n29593_,
    new_n29594_, new_n29595_, new_n29596_, new_n29597_, new_n29598_,
    new_n29599_, new_n29600_, new_n29601_, new_n29602_, new_n29603_,
    new_n29604_, new_n29605_, new_n29606_, new_n29607_, new_n29608_,
    new_n29609_, new_n29610_, new_n29611_, new_n29612_, new_n29613_,
    new_n29614_, new_n29615_, new_n29616_, new_n29617_, new_n29618_,
    new_n29619_, new_n29620_, new_n29621_, new_n29622_, new_n29623_,
    new_n29624_, new_n29625_, new_n29626_, new_n29627_, new_n29628_,
    new_n29629_, new_n29630_, new_n29631_, new_n29632_, new_n29633_,
    new_n29634_, new_n29635_, new_n29636_, new_n29637_, new_n29638_,
    new_n29640_, new_n29641_, new_n29642_, new_n29643_, new_n29644_,
    new_n29645_, new_n29646_, new_n29647_, new_n29648_, new_n29649_,
    new_n29650_, new_n29651_, new_n29652_, new_n29653_, new_n29654_,
    new_n29655_, new_n29656_, new_n29657_, new_n29658_, new_n29659_,
    new_n29660_, new_n29661_, new_n29662_, new_n29663_, new_n29664_,
    new_n29665_, new_n29666_, new_n29667_, new_n29668_, new_n29669_,
    new_n29670_, new_n29671_, new_n29672_, new_n29673_, new_n29674_,
    new_n29675_, new_n29676_, new_n29677_, new_n29678_, new_n29679_,
    new_n29680_, new_n29681_, new_n29682_, new_n29683_, new_n29684_,
    new_n29685_, new_n29686_, new_n29687_, new_n29688_, new_n29689_,
    new_n29690_, new_n29691_, new_n29692_, new_n29693_, new_n29694_,
    new_n29695_, new_n29696_, new_n29697_, new_n29698_, new_n29699_,
    new_n29700_, new_n29701_, new_n29702_, new_n29703_, new_n29704_,
    new_n29705_, new_n29706_, new_n29707_, new_n29708_, new_n29709_,
    new_n29710_, new_n29711_, new_n29712_, new_n29713_, new_n29714_,
    new_n29715_, new_n29716_, new_n29717_, new_n29718_, new_n29719_,
    new_n29720_, new_n29721_, new_n29722_, new_n29723_, new_n29724_,
    new_n29725_, new_n29726_, new_n29727_, new_n29728_, new_n29729_,
    new_n29730_, new_n29731_, new_n29732_, new_n29733_, new_n29734_,
    new_n29735_, new_n29736_, new_n29737_, new_n29738_, new_n29739_,
    new_n29740_, new_n29741_, new_n29742_, new_n29743_, new_n29744_,
    new_n29745_, new_n29746_, new_n29747_, new_n29748_, new_n29749_,
    new_n29750_, new_n29751_, new_n29752_, new_n29753_, new_n29754_,
    new_n29755_, new_n29756_, new_n29757_, new_n29758_, new_n29759_,
    new_n29760_, new_n29761_, new_n29762_, new_n29763_, new_n29764_,
    new_n29765_, new_n29766_, new_n29767_, new_n29768_, new_n29769_,
    new_n29770_, new_n29771_, new_n29772_, new_n29773_, new_n29774_,
    new_n29775_, new_n29776_, new_n29777_, new_n29778_, new_n29779_,
    new_n29780_, new_n29781_, new_n29782_, new_n29783_, new_n29784_,
    new_n29785_, new_n29786_, new_n29787_, new_n29788_, new_n29789_,
    new_n29790_, new_n29791_, new_n29792_, new_n29793_, new_n29794_,
    new_n29795_, new_n29796_, new_n29797_, new_n29798_, new_n29799_,
    new_n29800_, new_n29801_, new_n29802_, new_n29803_, new_n29804_,
    new_n29805_, new_n29806_, new_n29807_, new_n29808_, new_n29809_,
    new_n29810_, new_n29811_, new_n29812_, new_n29813_, new_n29814_,
    new_n29815_, new_n29816_, new_n29817_, new_n29818_, new_n29819_,
    new_n29820_, new_n29821_, new_n29822_, new_n29823_, new_n29824_,
    new_n29825_, new_n29826_, new_n29827_, new_n29828_, new_n29829_,
    new_n29830_, new_n29831_, new_n29832_, new_n29833_, new_n29834_,
    new_n29835_, new_n29836_, new_n29837_, new_n29838_, new_n29839_,
    new_n29840_, new_n29841_, new_n29842_, new_n29843_, new_n29844_,
    new_n29845_, new_n29846_, new_n29847_, new_n29848_, new_n29849_,
    new_n29850_, new_n29851_, new_n29852_, new_n29853_, new_n29854_,
    new_n29855_, new_n29856_, new_n29858_, new_n29859_, new_n29860_,
    new_n29861_, new_n29862_, new_n29863_, new_n29864_, new_n29865_,
    new_n29866_, new_n29867_, new_n29868_, new_n29869_, new_n29870_,
    new_n29871_, new_n29872_, new_n29873_, new_n29874_, new_n29875_,
    new_n29876_, new_n29877_, new_n29878_, new_n29879_, new_n29880_,
    new_n29881_, new_n29882_, new_n29883_, new_n29884_, new_n29885_,
    new_n29886_, new_n29887_, new_n29888_, new_n29889_, new_n29890_,
    new_n29891_, new_n29892_, new_n29893_, new_n29894_, new_n29895_,
    new_n29896_, new_n29897_, new_n29898_, new_n29899_, new_n29900_,
    new_n29901_, new_n29902_, new_n29903_, new_n29904_, new_n29905_,
    new_n29906_, new_n29907_, new_n29908_, new_n29909_, new_n29910_,
    new_n29911_, new_n29912_, new_n29913_, new_n29914_, new_n29915_,
    new_n29916_, new_n29917_, new_n29919_, new_n29920_, new_n29921_,
    new_n29922_, new_n29923_, new_n29924_, new_n29925_, new_n29926_,
    new_n29927_, new_n29928_, new_n29929_, new_n29930_, new_n29931_,
    new_n29932_, new_n29933_, new_n29934_, new_n29935_, new_n29936_,
    new_n29937_, new_n29938_, new_n29939_, new_n29940_, new_n29941_,
    new_n29942_, new_n29943_, new_n29944_, new_n29945_, new_n29946_,
    new_n29947_, new_n29948_, new_n29949_, new_n29950_, new_n29951_,
    new_n29952_, new_n29953_, new_n29954_, new_n29955_, new_n29956_,
    new_n29957_, new_n29958_, new_n29959_, new_n29960_, new_n29961_,
    new_n29962_, new_n29963_, new_n29964_, new_n29965_, new_n29966_,
    new_n29967_, new_n29968_, new_n29969_, new_n29970_, new_n29971_,
    new_n29972_, new_n29973_, new_n29974_, new_n29975_, new_n29976_,
    new_n29977_, new_n29978_, new_n29979_, new_n29980_, new_n29981_,
    new_n29982_, new_n29983_, new_n29984_, new_n29985_, new_n29986_,
    new_n29987_, new_n29988_, new_n29989_, new_n29990_, new_n29991_,
    new_n29992_, new_n29993_, new_n29994_, new_n29995_, new_n29996_,
    new_n29997_, new_n29998_, new_n29999_, new_n30000_, new_n30001_,
    new_n30002_, new_n30003_, new_n30004_, new_n30005_, new_n30006_,
    new_n30007_, new_n30008_, new_n30009_, new_n30010_, new_n30011_,
    new_n30012_, new_n30013_, new_n30014_, new_n30015_, new_n30016_,
    new_n30017_, new_n30018_, new_n30019_, new_n30020_, new_n30021_,
    new_n30022_, new_n30023_, new_n30024_, new_n30025_, new_n30026_,
    new_n30027_, new_n30028_, new_n30029_, new_n30030_, new_n30031_,
    new_n30032_, new_n30033_, new_n30034_, new_n30035_, new_n30036_,
    new_n30037_, new_n30038_, new_n30039_, new_n30040_, new_n30041_,
    new_n30042_, new_n30043_, new_n30044_, new_n30045_, new_n30046_,
    new_n30047_, new_n30048_, new_n30049_, new_n30050_, new_n30051_,
    new_n30052_, new_n30053_, new_n30054_, new_n30055_, new_n30056_,
    new_n30057_, new_n30058_, new_n30059_, new_n30060_, new_n30061_,
    new_n30062_, new_n30063_, new_n30064_, new_n30065_, new_n30066_,
    new_n30067_, new_n30068_, new_n30069_, new_n30070_, new_n30071_,
    new_n30072_, new_n30073_, new_n30074_, new_n30075_, new_n30076_,
    new_n30077_, new_n30078_, new_n30079_, new_n30080_, new_n30081_,
    new_n30082_, new_n30083_, new_n30084_, new_n30085_, new_n30086_,
    new_n30087_, new_n30088_, new_n30089_, new_n30090_, new_n30091_,
    new_n30092_, new_n30093_, new_n30094_, new_n30095_, new_n30096_,
    new_n30097_, new_n30098_, new_n30099_, new_n30100_, new_n30101_,
    new_n30102_, new_n30103_, new_n30104_, new_n30105_, new_n30106_,
    new_n30107_, new_n30108_, new_n30109_, new_n30110_, new_n30111_,
    new_n30112_, new_n30113_, new_n30114_, new_n30115_, new_n30116_,
    new_n30117_, new_n30118_, new_n30119_, new_n30120_, new_n30121_,
    new_n30122_, new_n30123_, new_n30124_, new_n30125_, new_n30126_,
    new_n30127_, new_n30128_, new_n30129_, new_n30130_, new_n30131_,
    new_n30132_, new_n30133_, new_n30134_, new_n30135_, new_n30136_,
    new_n30137_, new_n30138_, new_n30139_, new_n30140_, new_n30141_,
    new_n30142_, new_n30143_, new_n30144_, new_n30145_, new_n30146_,
    new_n30147_, new_n30148_, new_n30149_, new_n30150_, new_n30151_,
    new_n30152_, new_n30153_, new_n30154_, new_n30155_, new_n30156_,
    new_n30157_, new_n30158_, new_n30159_, new_n30160_, new_n30161_,
    new_n30162_, new_n30163_, new_n30164_, new_n30165_, new_n30166_,
    new_n30167_, new_n30168_, new_n30169_, new_n30170_, new_n30171_,
    new_n30172_, new_n30173_, new_n30174_, new_n30175_, new_n30176_,
    new_n30177_, new_n30178_, new_n30179_, new_n30180_, new_n30181_,
    new_n30182_, new_n30183_, new_n30184_, new_n30185_, new_n30186_,
    new_n30187_, new_n30189_, new_n30190_, new_n30191_, new_n30192_,
    new_n30193_, new_n30194_, new_n30195_, new_n30196_, new_n30197_,
    new_n30198_, new_n30199_, new_n30200_, new_n30201_, new_n30202_,
    new_n30203_, new_n30204_, new_n30205_, new_n30206_, new_n30207_,
    new_n30208_, new_n30209_, new_n30210_, new_n30211_, new_n30212_,
    new_n30213_, new_n30214_, new_n30215_, new_n30216_, new_n30217_,
    new_n30218_, new_n30219_, new_n30220_, new_n30221_, new_n30222_,
    new_n30223_, new_n30224_, new_n30226_, new_n30227_, new_n30228_,
    new_n30229_, new_n30230_, new_n30231_, new_n30232_, new_n30233_,
    new_n30234_, new_n30235_, new_n30236_, new_n30237_, new_n30238_,
    new_n30239_, new_n30240_, new_n30241_, new_n30242_, new_n30243_,
    new_n30244_, new_n30245_, new_n30246_, new_n30247_, new_n30248_,
    new_n30249_, new_n30250_, new_n30251_, new_n30252_, new_n30253_,
    new_n30254_, new_n30255_, new_n30256_, new_n30257_, new_n30258_,
    new_n30259_, new_n30260_, new_n30261_, new_n30262_, new_n30263_,
    new_n30264_, new_n30265_, new_n30266_, new_n30267_, new_n30268_,
    new_n30269_, new_n30270_, new_n30271_, new_n30272_, new_n30273_,
    new_n30274_, new_n30275_, new_n30276_, new_n30277_, new_n30278_,
    new_n30279_, new_n30280_, new_n30281_, new_n30282_, new_n30283_,
    new_n30284_, new_n30285_, new_n30286_, new_n30287_, new_n30288_,
    new_n30289_, new_n30290_, new_n30291_, new_n30292_, new_n30293_,
    new_n30294_, new_n30295_, new_n30296_, new_n30297_, new_n30298_,
    new_n30299_, new_n30300_, new_n30301_, new_n30302_, new_n30303_,
    new_n30304_, new_n30305_, new_n30306_, new_n30307_, new_n30308_,
    new_n30309_, new_n30310_, new_n30311_, new_n30312_, new_n30313_,
    new_n30314_, new_n30315_, new_n30316_, new_n30317_, new_n30318_,
    new_n30319_, new_n30320_, new_n30321_, new_n30322_, new_n30323_,
    new_n30324_, new_n30325_, new_n30326_, new_n30327_, new_n30328_,
    new_n30329_, new_n30330_, new_n30331_, new_n30332_, new_n30333_,
    new_n30334_, new_n30335_, new_n30336_, new_n30337_, new_n30338_,
    new_n30339_, new_n30340_, new_n30341_, new_n30342_, new_n30343_,
    new_n30344_, new_n30345_, new_n30346_, new_n30347_, new_n30348_,
    new_n30349_, new_n30350_, new_n30351_, new_n30352_, new_n30353_,
    new_n30354_, new_n30355_, new_n30356_, new_n30357_, new_n30358_,
    new_n30359_, new_n30360_, new_n30361_, new_n30362_, new_n30363_,
    new_n30364_, new_n30365_, new_n30366_, new_n30367_, new_n30368_,
    new_n30369_, new_n30370_, new_n30371_, new_n30372_, new_n30373_,
    new_n30374_, new_n30375_, new_n30376_, new_n30377_, new_n30378_,
    new_n30379_, new_n30380_, new_n30381_, new_n30382_, new_n30383_,
    new_n30384_, new_n30385_, new_n30386_, new_n30387_, new_n30388_,
    new_n30389_, new_n30390_, new_n30391_, new_n30392_, new_n30393_,
    new_n30394_, new_n30395_, new_n30396_, new_n30397_, new_n30398_,
    new_n30399_, new_n30400_, new_n30401_, new_n30402_, new_n30403_,
    new_n30404_, new_n30405_, new_n30406_, new_n30407_, new_n30408_,
    new_n30409_, new_n30410_, new_n30411_, new_n30412_, new_n30413_,
    new_n30414_, new_n30416_, new_n30417_, new_n30418_, new_n30419_,
    new_n30420_, new_n30421_, new_n30422_, new_n30423_, new_n30424_,
    new_n30425_, new_n30426_, new_n30427_, new_n30428_, new_n30429_,
    new_n30430_, new_n30431_, new_n30432_, new_n30433_, new_n30434_,
    new_n30435_, new_n30436_, new_n30437_, new_n30438_, new_n30439_,
    new_n30440_, new_n30441_, new_n30442_, new_n30443_, new_n30444_,
    new_n30445_, new_n30446_, new_n30447_, new_n30448_, new_n30449_,
    new_n30450_, new_n30451_, new_n30452_, new_n30453_, new_n30454_,
    new_n30455_, new_n30456_, new_n30457_, new_n30458_, new_n30459_,
    new_n30460_, new_n30461_, new_n30462_, new_n30463_, new_n30464_,
    new_n30465_, new_n30466_, new_n30467_, new_n30468_, new_n30469_,
    new_n30470_, new_n30471_, new_n30472_, new_n30473_, new_n30474_,
    new_n30475_, new_n30476_, new_n30477_, new_n30478_, new_n30479_,
    new_n30480_, new_n30481_, new_n30482_, new_n30483_, new_n30484_,
    new_n30485_, new_n30486_, new_n30487_, new_n30488_, new_n30489_,
    new_n30490_, new_n30491_, new_n30492_, new_n30493_, new_n30494_,
    new_n30495_, new_n30496_, new_n30497_, new_n30498_, new_n30499_,
    new_n30500_, new_n30501_, new_n30502_, new_n30503_, new_n30504_,
    new_n30505_, new_n30506_, new_n30507_, new_n30508_, new_n30509_,
    new_n30510_, new_n30511_, new_n30512_, new_n30513_, new_n30514_,
    new_n30515_, new_n30516_, new_n30517_, new_n30518_, new_n30519_,
    new_n30520_, new_n30521_, new_n30522_, new_n30523_, new_n30524_,
    new_n30525_, new_n30526_, new_n30527_, new_n30528_, new_n30529_,
    new_n30530_, new_n30531_, new_n30532_, new_n30533_, new_n30534_,
    new_n30535_, new_n30536_, new_n30537_, new_n30538_, new_n30539_,
    new_n30540_, new_n30541_, new_n30542_, new_n30543_, new_n30544_,
    new_n30545_, new_n30546_, new_n30547_, new_n30548_, new_n30549_,
    new_n30550_, new_n30551_, new_n30552_, new_n30553_, new_n30554_,
    new_n30555_, new_n30556_, new_n30557_, new_n30558_, new_n30559_,
    new_n30560_, new_n30561_, new_n30562_, new_n30563_, new_n30564_,
    new_n30565_, new_n30566_, new_n30567_, new_n30568_, new_n30569_,
    new_n30570_, new_n30571_, new_n30572_, new_n30573_, new_n30574_,
    new_n30575_, new_n30576_, new_n30577_, new_n30578_, new_n30579_,
    new_n30580_, new_n30581_, new_n30582_, new_n30583_, new_n30584_,
    new_n30585_, new_n30586_, new_n30587_, new_n30588_, new_n30589_,
    new_n30590_, new_n30591_, new_n30592_, new_n30593_, new_n30594_,
    new_n30596_, new_n30597_, new_n30598_, new_n30599_, new_n30600_,
    new_n30601_, new_n30602_, new_n30603_, new_n30604_, new_n30605_,
    new_n30606_, new_n30607_, new_n30608_, new_n30609_, new_n30610_,
    new_n30611_, new_n30612_, new_n30613_, new_n30614_, new_n30615_,
    new_n30616_, new_n30617_, new_n30618_, new_n30619_, new_n30620_,
    new_n30621_, new_n30622_, new_n30623_, new_n30624_, new_n30625_,
    new_n30626_, new_n30627_, new_n30628_, new_n30629_, new_n30630_,
    new_n30631_, new_n30632_, new_n30633_, new_n30634_, new_n30635_,
    new_n30636_, new_n30637_, new_n30638_, new_n30639_, new_n30640_,
    new_n30641_, new_n30642_, new_n30643_, new_n30644_, new_n30645_,
    new_n30646_, new_n30647_, new_n30648_, new_n30649_, new_n30650_,
    new_n30651_, new_n30652_, new_n30653_, new_n30654_, new_n30655_,
    new_n30656_, new_n30657_, new_n30658_, new_n30659_, new_n30660_,
    new_n30661_, new_n30662_, new_n30663_, new_n30664_, new_n30665_,
    new_n30666_, new_n30667_, new_n30668_, new_n30669_, new_n30670_,
    new_n30671_, new_n30672_, new_n30673_, new_n30674_, new_n30675_,
    new_n30676_, new_n30677_, new_n30678_, new_n30679_, new_n30680_,
    new_n30681_, new_n30682_, new_n30683_, new_n30684_, new_n30685_,
    new_n30686_, new_n30687_, new_n30688_, new_n30689_, new_n30690_,
    new_n30691_, new_n30692_, new_n30693_, new_n30694_, new_n30695_,
    new_n30696_, new_n30697_, new_n30698_, new_n30699_, new_n30700_,
    new_n30701_, new_n30702_, new_n30703_, new_n30704_, new_n30705_,
    new_n30706_, new_n30707_, new_n30708_, new_n30709_, new_n30710_,
    new_n30711_, new_n30712_, new_n30713_, new_n30714_, new_n30715_,
    new_n30716_, new_n30717_, new_n30718_, new_n30719_, new_n30720_,
    new_n30721_, new_n30722_, new_n30723_, new_n30724_, new_n30725_,
    new_n30726_, new_n30727_, new_n30728_, new_n30729_, new_n30730_,
    new_n30731_, new_n30732_, new_n30733_, new_n30734_, new_n30735_,
    new_n30736_, new_n30737_, new_n30738_, new_n30739_, new_n30740_,
    new_n30741_, new_n30742_, new_n30743_, new_n30744_, new_n30745_,
    new_n30746_, new_n30747_, new_n30748_, new_n30749_, new_n30750_,
    new_n30751_, new_n30752_, new_n30753_, new_n30754_, new_n30755_,
    new_n30756_, new_n30757_, new_n30758_, new_n30760_, new_n30761_,
    new_n30762_, new_n30763_, new_n30764_, new_n30765_, new_n30766_,
    new_n30767_, new_n30768_, new_n30769_, new_n30770_, new_n30771_,
    new_n30772_, new_n30773_, new_n30774_, new_n30775_, new_n30776_,
    new_n30777_, new_n30778_, new_n30779_, new_n30780_, new_n30781_,
    new_n30782_, new_n30783_, new_n30784_, new_n30785_, new_n30786_,
    new_n30787_, new_n30788_, new_n30789_, new_n30790_, new_n30791_,
    new_n30792_, new_n30793_, new_n30794_, new_n30795_, new_n30796_,
    new_n30797_, new_n30798_, new_n30799_, new_n30800_, new_n30801_,
    new_n30802_, new_n30803_, new_n30804_, new_n30805_, new_n30806_,
    new_n30807_, new_n30808_, new_n30809_, new_n30810_, new_n30811_,
    new_n30812_, new_n30813_, new_n30814_, new_n30815_, new_n30816_,
    new_n30817_, new_n30818_, new_n30819_, new_n30820_, new_n30821_,
    new_n30822_, new_n30823_, new_n30824_, new_n30825_, new_n30826_,
    new_n30827_, new_n30828_, new_n30829_, new_n30830_, new_n30831_,
    new_n30832_, new_n30833_, new_n30834_, new_n30835_, new_n30836_,
    new_n30837_, new_n30838_, new_n30839_, new_n30840_, new_n30841_,
    new_n30842_, new_n30843_, new_n30844_, new_n30845_, new_n30846_,
    new_n30847_, new_n30848_, new_n30849_, new_n30850_, new_n30851_,
    new_n30852_, new_n30853_, new_n30854_, new_n30855_, new_n30856_,
    new_n30857_, new_n30858_, new_n30859_, new_n30860_, new_n30861_,
    new_n30862_, new_n30863_, new_n30864_, new_n30866_, new_n30867_,
    new_n30868_, new_n30869_, new_n30870_, new_n30871_, new_n30872_,
    new_n30873_, new_n30874_, new_n30875_, new_n30876_, new_n30877_,
    new_n30878_, new_n30879_, new_n30880_, new_n30881_, new_n30882_,
    new_n30883_, new_n30884_, new_n30885_, new_n30886_, new_n30887_,
    new_n30888_, new_n30889_, new_n30890_, new_n30891_, new_n30892_,
    new_n30893_, new_n30894_, new_n30895_, new_n30896_, new_n30897_,
    new_n30898_, new_n30899_, new_n30900_, new_n30901_, new_n30902_,
    new_n30903_, new_n30904_, new_n30905_, new_n30906_, new_n30907_,
    new_n30908_, new_n30909_, new_n30910_, new_n30911_, new_n30912_,
    new_n30913_, new_n30914_, new_n30915_, new_n30916_, new_n30917_,
    new_n30918_, new_n30919_, new_n30920_, new_n30921_, new_n30922_,
    new_n30923_, new_n30924_, new_n30925_, new_n30926_, new_n30927_,
    new_n30928_, new_n30929_, new_n30930_, new_n30931_, new_n30932_,
    new_n30933_, new_n30934_, new_n30935_, new_n30936_, new_n30937_,
    new_n30938_, new_n30939_, new_n30940_, new_n30941_, new_n30942_,
    new_n30943_, new_n30944_, new_n30945_, new_n30946_, new_n30947_,
    new_n30948_, new_n30949_, new_n30950_, new_n30951_, new_n30952_,
    new_n30953_, new_n30954_, new_n30955_, new_n30956_, new_n30957_,
    new_n30958_, new_n30959_, new_n30960_, new_n30961_, new_n30962_,
    new_n30963_, new_n30964_, new_n30965_, new_n30966_, new_n30967_,
    new_n30968_, new_n30969_, new_n30970_, new_n30971_, new_n30972_,
    new_n30973_, new_n30974_, new_n30975_, new_n30976_, new_n30977_,
    new_n30978_, new_n30979_, new_n30980_, new_n30981_, new_n30982_,
    new_n30983_, new_n30984_, new_n30985_, new_n30986_, new_n30987_,
    new_n30989_, new_n30990_, new_n30991_, new_n30993_, new_n30994_,
    new_n30995_, new_n30996_, new_n30997_, new_n30998_, new_n30999_,
    new_n31000_, new_n31002_, new_n31003_, new_n31004_, new_n31005_,
    new_n31006_, new_n31007_, new_n31008_, new_n31009_, new_n31010_,
    new_n31011_, new_n31012_, new_n31013_, new_n31014_, new_n31015_,
    new_n31016_, new_n31017_, new_n31018_, new_n31019_, new_n31020_,
    new_n31021_, new_n31022_, new_n31023_, new_n31024_, new_n31025_,
    new_n31026_, new_n31028_, new_n31029_, new_n31030_, new_n31031_,
    new_n31032_, new_n31033_, new_n31034_, new_n31035_, new_n31036_,
    new_n31037_, new_n31038_, new_n31039_, new_n31040_, new_n31041_,
    new_n31042_, new_n31043_, new_n31044_, new_n31045_, new_n31046_,
    new_n31047_, new_n31048_, new_n31049_, new_n31050_, new_n31051_,
    new_n31052_, new_n31053_, new_n31054_, new_n31055_, new_n31056_,
    new_n31057_, new_n31058_, new_n31059_, new_n31060_, new_n31061_,
    new_n31062_, new_n31063_, new_n31064_, new_n31065_, new_n31066_,
    new_n31067_, new_n31068_, new_n31069_, new_n31070_, new_n31071_,
    new_n31072_, new_n31073_, new_n31074_, new_n31075_, new_n31076_,
    new_n31077_, new_n31078_, new_n31079_, new_n31080_, new_n31081_,
    new_n31082_, new_n31083_, new_n31084_, new_n31085_, new_n31086_,
    new_n31087_, new_n31088_, new_n31089_, new_n31090_, new_n31091_,
    new_n31092_, new_n31093_, new_n31094_, new_n31095_, new_n31096_,
    new_n31097_, new_n31098_, new_n31099_, new_n31100_, new_n31101_,
    new_n31102_, new_n31103_, new_n31104_, new_n31105_, new_n31106_,
    new_n31107_, new_n31108_, new_n31109_, new_n31110_, new_n31111_,
    new_n31112_, new_n31113_, new_n31114_, new_n31115_, new_n31116_,
    new_n31117_, new_n31118_, new_n31119_, new_n31120_, new_n31121_,
    new_n31122_, new_n31123_, new_n31124_, new_n31125_, new_n31126_,
    new_n31127_, new_n31128_, new_n31129_, new_n31130_, new_n31131_,
    new_n31132_, new_n31133_, new_n31134_, new_n31135_, new_n31136_,
    new_n31137_, new_n31138_, new_n31139_, new_n31140_, new_n31141_,
    new_n31142_, new_n31143_, new_n31144_, new_n31145_, new_n31146_,
    new_n31147_, new_n31148_, new_n31149_, new_n31150_, new_n31151_,
    new_n31152_, new_n31153_, new_n31154_, new_n31155_, new_n31156_,
    new_n31157_, new_n31158_, new_n31159_, new_n31160_, new_n31161_,
    new_n31162_, new_n31163_, new_n31164_, new_n31165_, new_n31166_,
    new_n31167_, new_n31168_, new_n31169_, new_n31170_, new_n31171_,
    new_n31172_, new_n31173_, new_n31174_, new_n31175_, new_n31176_,
    new_n31177_, new_n31178_, new_n31179_, new_n31180_, new_n31181_,
    new_n31182_, new_n31183_, new_n31184_, new_n31185_, new_n31186_,
    new_n31187_, new_n31188_, new_n31189_, new_n31190_, new_n31191_,
    new_n31192_, new_n31193_, new_n31194_, new_n31195_, new_n31197_,
    new_n31198_, new_n31199_, new_n31200_, new_n31201_, new_n31202_,
    new_n31203_, new_n31204_, new_n31205_, new_n31206_, new_n31207_,
    new_n31208_, new_n31209_, new_n31210_, new_n31211_, new_n31212_,
    new_n31213_, new_n31214_, new_n31215_, new_n31216_, new_n31217_,
    new_n31218_, new_n31219_, new_n31220_, new_n31221_, new_n31222_,
    new_n31223_, new_n31224_, new_n31225_, new_n31226_, new_n31227_,
    new_n31228_, new_n31229_, new_n31230_, new_n31231_, new_n31232_,
    new_n31233_, new_n31234_, new_n31235_, new_n31236_, new_n31237_,
    new_n31238_, new_n31239_, new_n31240_, new_n31241_, new_n31242_,
    new_n31243_, new_n31244_, new_n31245_, new_n31246_, new_n31247_,
    new_n31248_, new_n31249_, new_n31250_, new_n31251_, new_n31252_,
    new_n31253_, new_n31254_, new_n31255_, new_n31256_, new_n31257_,
    new_n31258_, new_n31259_, new_n31260_, new_n31261_, new_n31262_,
    new_n31263_, new_n31264_, new_n31265_, new_n31266_, new_n31267_,
    new_n31268_, new_n31269_, new_n31270_, new_n31271_, new_n31272_,
    new_n31273_, new_n31274_, new_n31275_, new_n31276_, new_n31277_,
    new_n31278_, new_n31279_, new_n31280_, new_n31281_, new_n31282_,
    new_n31283_, new_n31284_, new_n31285_, new_n31286_, new_n31287_,
    new_n31288_, new_n31289_, new_n31290_, new_n31291_, new_n31292_,
    new_n31293_, new_n31294_, new_n31295_, new_n31296_, new_n31297_,
    new_n31298_, new_n31299_, new_n31300_, new_n31301_, new_n31302_,
    new_n31303_, new_n31304_, new_n31305_, new_n31306_, new_n31307_,
    new_n31308_, new_n31309_, new_n31310_, new_n31311_, new_n31312_,
    new_n31313_, new_n31314_, new_n31315_, new_n31316_, new_n31317_,
    new_n31318_, new_n31319_, new_n31320_, new_n31321_, new_n31322_,
    new_n31323_, new_n31324_, new_n31325_, new_n31326_, new_n31327_,
    new_n31328_, new_n31329_, new_n31330_, new_n31331_, new_n31332_,
    new_n31333_, new_n31334_, new_n31335_, new_n31337_, new_n31338_,
    new_n31339_, new_n31340_, new_n31341_, new_n31343_, new_n31344_,
    new_n31345_, new_n31346_, new_n31347_, new_n31349_, new_n31350_,
    new_n31351_, new_n31352_, new_n31353_, new_n31355_, new_n31356_,
    new_n31357_, new_n31358_, new_n31359_, new_n31361_, new_n31362_,
    new_n31363_, new_n31364_, new_n31365_, new_n31367_, new_n31368_,
    new_n31369_, new_n31370_, new_n31371_, new_n31373_, new_n31374_,
    new_n31375_, new_n31376_, new_n31377_, new_n31379_, new_n31380_,
    new_n31381_, new_n31382_, new_n31383_, new_n31384_, new_n31385_,
    new_n31386_, new_n31387_, new_n31388_, new_n31389_, new_n31390_,
    new_n31391_, new_n31392_, new_n31393_, new_n31394_, new_n31395_,
    new_n31396_, new_n31397_, new_n31398_, new_n31399_, new_n31400_,
    new_n31401_, new_n31403_, new_n31404_, new_n31405_, new_n31406_,
    new_n31407_, new_n31408_, new_n31409_, new_n31410_, new_n31411_,
    new_n31412_, new_n31413_, new_n31414_, new_n31415_, new_n31416_,
    new_n31417_, new_n31418_, new_n31419_, new_n31420_, new_n31421_,
    new_n31422_, new_n31423_, new_n31424_, new_n31425_, new_n31426_,
    new_n31427_, new_n31428_, new_n31429_, new_n31430_, new_n31431_,
    new_n31432_, new_n31433_, new_n31434_, new_n31435_, new_n31436_,
    new_n31437_, new_n31438_, new_n31439_, new_n31440_, new_n31441_,
    new_n31442_, new_n31443_, new_n31444_, new_n31445_, new_n31446_,
    new_n31447_, new_n31448_, new_n31449_, new_n31450_, new_n31451_,
    new_n31452_, new_n31453_, new_n31454_, new_n31455_, new_n31456_,
    new_n31457_, new_n31458_, new_n31459_, new_n31460_, new_n31461_,
    new_n31462_, new_n31463_, new_n31464_, new_n31465_, new_n31466_,
    new_n31467_, new_n31468_, new_n31469_, new_n31470_, new_n31471_,
    new_n31472_, new_n31473_, new_n31474_, new_n31475_, new_n31476_,
    new_n31477_, new_n31478_, new_n31479_, new_n31480_, new_n31481_,
    new_n31482_, new_n31483_, new_n31484_, new_n31485_, new_n31486_,
    new_n31487_, new_n31488_, new_n31489_, new_n31490_, new_n31491_,
    new_n31492_, new_n31493_, new_n31494_, new_n31495_, new_n31496_,
    new_n31497_, new_n31498_, new_n31499_, new_n31500_, new_n31501_,
    new_n31502_, new_n31503_, new_n31504_, new_n31505_, new_n31506_,
    new_n31507_, new_n31508_, new_n31509_, new_n31510_, new_n31511_,
    new_n31512_, new_n31513_, new_n31514_, new_n31515_, new_n31516_,
    new_n31517_, new_n31518_, new_n31519_, new_n31520_, new_n31521_,
    new_n31522_, new_n31523_, new_n31524_, new_n31525_, new_n31526_,
    new_n31527_, new_n31528_, new_n31529_, new_n31530_, new_n31531_,
    new_n31532_, new_n31533_, new_n31534_, new_n31535_, new_n31536_,
    new_n31537_, new_n31538_, new_n31539_, new_n31540_, new_n31541_,
    new_n31542_, new_n31543_, new_n31545_, new_n31546_, new_n31547_,
    new_n31548_, new_n31549_, new_n31550_, new_n31551_, new_n31552_,
    new_n31553_, new_n31554_, new_n31555_, new_n31556_, new_n31557_,
    new_n31558_, new_n31559_, new_n31560_, new_n31561_, new_n31562_,
    new_n31563_, new_n31564_, new_n31565_, new_n31566_, new_n31567_,
    new_n31568_, new_n31569_, new_n31570_, new_n31571_, new_n31572_,
    new_n31573_, new_n31574_, new_n31575_, new_n31576_, new_n31577_,
    new_n31579_, new_n31580_, new_n31581_, new_n31582_, new_n31583_,
    new_n31584_, new_n31585_, new_n31586_, new_n31587_, new_n31588_,
    new_n31589_, new_n31590_, new_n31591_, new_n31592_, new_n31593_,
    new_n31594_, new_n31595_, new_n31596_, new_n31597_, new_n31598_,
    new_n31599_, new_n31600_, new_n31601_, new_n31602_, new_n31603_,
    new_n31605_, new_n31606_, new_n31607_, new_n31608_, new_n31609_,
    new_n31610_, new_n31611_, new_n31612_, new_n31613_, new_n31614_,
    new_n31615_, new_n31616_, new_n31617_, new_n31618_, new_n31619_,
    new_n31620_, new_n31621_, new_n31622_, new_n31623_, new_n31624_,
    new_n31625_, new_n31626_, new_n31627_, new_n31628_, new_n31629_,
    new_n31630_, new_n31631_, new_n31632_, new_n31633_, new_n31634_,
    new_n31635_, new_n31636_, new_n31637_, new_n31638_, new_n31639_,
    new_n31640_, new_n31641_, new_n31642_, new_n31643_, new_n31644_,
    new_n31645_, new_n31646_, new_n31648_, new_n31649_, new_n31650_,
    new_n31651_, new_n31652_, new_n31653_, new_n31654_, new_n31655_,
    new_n31656_, new_n31657_, new_n31658_, new_n31659_, new_n31660_,
    new_n31661_, new_n31662_, new_n31663_, new_n31664_, new_n31665_,
    new_n31666_, new_n31667_, new_n31668_, new_n31669_, new_n31670_,
    new_n31671_, new_n31672_, new_n31673_, new_n31674_, new_n31675_,
    new_n31676_, new_n31677_, new_n31678_, new_n31679_, new_n31680_,
    new_n31681_, new_n31682_, new_n31683_, new_n31684_, new_n31685_,
    new_n31686_, new_n31687_, new_n31688_, new_n31689_, new_n31690_,
    new_n31691_, new_n31692_, new_n31693_, new_n31694_, new_n31695_,
    new_n31696_, new_n31697_, new_n31698_, new_n31699_, new_n31700_,
    new_n31701_, new_n31702_, new_n31703_, new_n31704_, new_n31705_,
    new_n31706_, new_n31707_, new_n31708_, new_n31709_, new_n31710_,
    new_n31711_, new_n31712_, new_n31713_, new_n31714_, new_n31715_,
    new_n31716_, new_n31717_, new_n31718_, new_n31719_, new_n31720_,
    new_n31721_, new_n31722_, new_n31723_, new_n31724_, new_n31725_,
    new_n31726_, new_n31727_, new_n31728_, new_n31729_, new_n31730_,
    new_n31731_, new_n31732_, new_n31733_, new_n31734_, new_n31735_,
    new_n31736_, new_n31737_, new_n31738_, new_n31739_, new_n31740_,
    new_n31741_, new_n31742_, new_n31743_, new_n31744_, new_n31745_,
    new_n31746_, new_n31747_, new_n31748_, new_n31749_, new_n31750_,
    new_n31751_, new_n31752_, new_n31753_, new_n31754_, new_n31755_,
    new_n31756_, new_n31757_, new_n31758_, new_n31759_, new_n31760_,
    new_n31761_, new_n31762_, new_n31763_, new_n31764_, new_n31765_,
    new_n31766_, new_n31767_, new_n31768_, new_n31769_, new_n31770_,
    new_n31771_, new_n31772_, new_n31773_, new_n31774_, new_n31775_,
    new_n31776_, new_n31777_, new_n31778_, new_n31780_, new_n31781_,
    new_n31782_, new_n31783_, new_n31784_, new_n31785_, new_n31786_,
    new_n31787_, new_n31788_, new_n31789_, new_n31790_, new_n31791_,
    new_n31792_, new_n31793_, new_n31794_, new_n31795_, new_n31796_,
    new_n31797_, new_n31798_, new_n31799_, new_n31800_, new_n31801_,
    new_n31802_, new_n31803_, new_n31804_, new_n31805_, new_n31806_,
    new_n31807_, new_n31808_, new_n31809_, new_n31810_, new_n31811_,
    new_n31812_, new_n31813_, new_n31814_, new_n31815_, new_n31816_,
    new_n31817_, new_n31818_, new_n31819_, new_n31820_, new_n31821_,
    new_n31822_, new_n31823_, new_n31824_, new_n31825_, new_n31826_,
    new_n31827_, new_n31828_, new_n31829_, new_n31830_, new_n31831_,
    new_n31832_, new_n31833_, new_n31834_, new_n31835_, new_n31836_,
    new_n31837_, new_n31838_, new_n31839_, new_n31840_, new_n31841_,
    new_n31842_, new_n31843_, new_n31844_, new_n31845_, new_n31846_,
    new_n31847_, new_n31848_, new_n31849_, new_n31850_, new_n31851_,
    new_n31852_, new_n31853_, new_n31854_, new_n31855_, new_n31856_,
    new_n31857_, new_n31858_, new_n31859_, new_n31860_, new_n31861_,
    new_n31862_, new_n31863_, new_n31864_, new_n31865_, new_n31866_,
    new_n31867_, new_n31868_, new_n31869_, new_n31870_, new_n31871_,
    new_n31872_, new_n31873_, new_n31874_, new_n31875_, new_n31876_,
    new_n31877_, new_n31878_, new_n31879_, new_n31880_, new_n31881_,
    new_n31882_, new_n31883_, new_n31884_, new_n31885_, new_n31886_,
    new_n31887_, new_n31888_, new_n31889_, new_n31890_, new_n31891_,
    new_n31892_, new_n31893_, new_n31894_, new_n31895_, new_n31896_,
    new_n31898_, new_n31899_, new_n31900_, new_n31901_, new_n31902_,
    new_n31903_, new_n31904_, new_n31905_, new_n31906_, new_n31907_,
    new_n31908_, new_n31909_, new_n31910_, new_n31911_, new_n31912_,
    new_n31913_, new_n31914_, new_n31915_, new_n31916_, new_n31917_,
    new_n31918_, new_n31919_, new_n31920_, new_n31921_, new_n31922_,
    new_n31923_, new_n31924_, new_n31925_, new_n31926_, new_n31927_,
    new_n31928_, new_n31930_, new_n31931_, new_n31932_, new_n31933_,
    new_n31934_, new_n31935_, new_n31936_, new_n31937_, new_n31938_,
    new_n31939_, new_n31940_, new_n31941_, new_n31942_, new_n31943_,
    new_n31944_, new_n31945_, new_n31946_, new_n31947_, new_n31948_,
    new_n31949_, new_n31950_, new_n31951_, new_n31952_, new_n31953_,
    new_n31954_, new_n31955_, new_n31957_, new_n31958_, new_n31959_,
    new_n31960_, new_n31961_, new_n31962_, new_n31963_, new_n31964_,
    new_n31965_, new_n31966_, new_n31967_, new_n31968_, new_n31969_,
    new_n31970_, new_n31971_, new_n31972_, new_n31973_, new_n31974_,
    new_n31975_, new_n31976_, new_n31977_, new_n31978_, new_n31979_,
    new_n31980_, new_n31981_, new_n31982_, new_n31983_, new_n31984_,
    new_n31985_, new_n31986_, new_n31987_, new_n31988_, new_n31989_,
    new_n31991_, new_n31992_, new_n31993_, new_n31994_, new_n31995_,
    new_n31996_, new_n31997_, new_n31998_, new_n31999_, new_n32000_,
    new_n32001_, new_n32002_, new_n32003_, new_n32004_, new_n32005_,
    new_n32006_, new_n32007_, new_n32008_, new_n32009_, new_n32010_,
    new_n32011_, new_n32012_, new_n32013_, new_n32014_, new_n32015_,
    new_n32016_, new_n32017_, new_n32018_, new_n32019_, new_n32020_,
    new_n32021_, new_n32022_, new_n32023_, new_n32024_, new_n32025_,
    new_n32026_, new_n32027_, new_n32028_, new_n32029_, new_n32030_,
    new_n32031_, new_n32032_, new_n32033_, new_n32034_, new_n32035_,
    new_n32036_, new_n32037_, new_n32038_, new_n32039_, new_n32040_,
    new_n32041_, new_n32042_, new_n32043_, new_n32044_, new_n32045_,
    new_n32046_, new_n32047_, new_n32048_, new_n32049_, new_n32050_,
    new_n32051_, new_n32052_, new_n32053_, new_n32054_, new_n32055_,
    new_n32056_, new_n32057_, new_n32058_, new_n32060_, new_n32061_,
    new_n32062_, new_n32063_, new_n32064_, new_n32065_, new_n32066_,
    new_n32067_, new_n32068_, new_n32069_, new_n32070_, new_n32071_,
    new_n32072_, new_n32073_, new_n32074_, new_n32075_, new_n32076_,
    new_n32077_, new_n32078_, new_n32079_, new_n32080_, new_n32081_,
    new_n32082_, new_n32083_, new_n32084_, new_n32085_, new_n32086_,
    new_n32087_, new_n32088_, new_n32089_, new_n32090_, new_n32091_,
    new_n32092_, new_n32093_, new_n32094_, new_n32095_, new_n32096_,
    new_n32097_, new_n32099_, new_n32100_, new_n32101_, new_n32102_,
    new_n32103_, new_n32104_, new_n32105_, new_n32106_, new_n32107_,
    new_n32108_, new_n32109_, new_n32110_, new_n32111_, new_n32112_,
    new_n32113_, new_n32114_, new_n32115_, new_n32116_, new_n32117_,
    new_n32118_, new_n32119_, new_n32120_, new_n32121_, new_n32122_,
    new_n32123_, new_n32125_, new_n32126_, new_n32127_, new_n32128_,
    new_n32129_, new_n32130_, new_n32131_, new_n32132_, new_n32133_,
    new_n32134_, new_n32135_, new_n32136_, new_n32137_, new_n32138_,
    new_n32139_, new_n32140_, new_n32141_, new_n32142_, new_n32143_,
    new_n32144_, new_n32145_, new_n32146_, new_n32147_, new_n32148_,
    new_n32149_, new_n32150_, new_n32151_, new_n32152_, new_n32153_,
    new_n32154_, new_n32155_, new_n32156_, new_n32157_, new_n32158_,
    new_n32159_, new_n32160_, new_n32161_, new_n32162_, new_n32163_,
    new_n32164_, new_n32165_, new_n32166_, new_n32167_, new_n32168_,
    new_n32169_, new_n32170_, new_n32172_, new_n32173_, new_n32174_,
    new_n32175_, new_n32176_, new_n32177_, new_n32178_, new_n32179_,
    new_n32180_, new_n32181_, new_n32182_, new_n32183_, new_n32184_,
    new_n32185_, new_n32186_, new_n32187_, new_n32188_, new_n32189_,
    new_n32190_, new_n32191_, new_n32193_, new_n32194_, new_n32195_,
    new_n32196_, new_n32197_, new_n32198_, new_n32199_, new_n32200_,
    new_n32201_, new_n32202_, new_n32203_, new_n32204_, new_n32205_,
    new_n32206_, new_n32207_, new_n32208_, new_n32209_, new_n32210_,
    new_n32211_, new_n32212_, new_n32213_, new_n32214_, new_n32215_,
    new_n32216_, new_n32217_, new_n32218_, new_n32219_, new_n32220_,
    new_n32221_, new_n32222_, new_n32223_, new_n32225_, new_n32226_,
    new_n32227_, new_n32228_, new_n32229_, new_n32230_, new_n32231_,
    new_n32232_, new_n32233_, new_n32234_, new_n32235_, new_n32236_,
    new_n32237_, new_n32238_, new_n32239_, new_n32240_, new_n32241_,
    new_n32242_, new_n32243_, new_n32244_, new_n32245_, new_n32246_,
    new_n32247_, new_n32248_, new_n32249_, new_n32250_, new_n32251_,
    new_n32252_, new_n32253_, new_n32254_, new_n32255_, new_n32256_,
    new_n32257_, new_n32258_, new_n32259_, new_n32260_, new_n32261_,
    new_n32262_, new_n32263_, new_n32264_, new_n32265_, new_n32266_,
    new_n32267_, new_n32268_, new_n32270_, new_n32271_, new_n32272_,
    new_n32273_, new_n32274_, new_n32275_, new_n32276_, new_n32277_,
    new_n32278_, new_n32279_, new_n32280_, new_n32281_, new_n32282_,
    new_n32283_, new_n32284_, new_n32285_, new_n32286_, new_n32287_,
    new_n32288_, new_n32289_, new_n32290_, new_n32291_, new_n32292_,
    new_n32293_, new_n32294_, new_n32295_, new_n32296_, new_n32297_,
    new_n32298_, new_n32299_, new_n32300_, new_n32301_, new_n32302_,
    new_n32303_, new_n32304_, new_n32305_, new_n32306_, new_n32308_,
    new_n32309_, new_n32310_, new_n32311_, new_n32312_, new_n32313_,
    new_n32314_, new_n32315_, new_n32316_, new_n32317_, new_n32318_,
    new_n32319_, new_n32320_, new_n32321_, new_n32322_, new_n32323_,
    new_n32324_, new_n32325_, new_n32326_, new_n32327_, new_n32328_,
    new_n32329_, new_n32330_, new_n32331_, new_n32332_, new_n32333_,
    new_n32334_, new_n32335_, new_n32336_, new_n32338_, new_n32339_,
    new_n32340_, new_n32341_, new_n32342_, new_n32343_, new_n32344_,
    new_n32345_, new_n32346_, new_n32347_, new_n32348_, new_n32349_,
    new_n32350_, new_n32351_, new_n32352_, new_n32353_, new_n32354_,
    new_n32355_, new_n32356_, new_n32357_, new_n32358_, new_n32359_,
    new_n32360_, new_n32361_, new_n32362_, new_n32364_, new_n32365_,
    new_n32366_, new_n32367_, new_n32368_, new_n32369_, new_n32370_,
    new_n32371_, new_n32372_, new_n32373_, new_n32374_, new_n32375_,
    new_n32376_, new_n32377_, new_n32378_, new_n32379_, new_n32380_,
    new_n32381_, new_n32382_, new_n32383_, new_n32384_, new_n32385_,
    new_n32386_, new_n32387_, new_n32388_, new_n32390_, new_n32391_,
    new_n32392_, new_n32393_, new_n32394_, new_n32395_, new_n32396_,
    new_n32397_, new_n32398_, new_n32399_, new_n32400_, new_n32401_,
    new_n32402_, new_n32403_, new_n32404_, new_n32405_, new_n32406_,
    new_n32407_, new_n32408_, new_n32409_, new_n32410_, new_n32411_,
    new_n32412_, new_n32413_, new_n32414_, new_n32415_, new_n32416_,
    new_n32417_, new_n32418_, new_n32419_, new_n32420_, new_n32421_,
    new_n32422_, new_n32423_, new_n32424_, new_n32425_, new_n32426_,
    new_n32427_, new_n32428_, new_n32430_, new_n32432_, new_n32433_,
    new_n32434_, new_n32435_, new_n32436_, new_n32437_, new_n32438_,
    new_n32439_, new_n32440_, new_n32441_, new_n32442_, new_n32443_,
    new_n32444_, new_n32445_, new_n32447_, new_n32448_, new_n32449_,
    new_n32450_, new_n32451_, new_n32452_, new_n32453_, new_n32454_,
    new_n32455_, new_n32456_, new_n32457_, new_n32461_, new_n32462_,
    new_n32464_, new_n32465_, new_n32466_, new_n32467_, new_n32468_,
    new_n32469_, new_n32470_, new_n32471_, new_n32472_, new_n32473_,
    new_n32475_, new_n32476_, new_n32478_, new_n32479_, new_n32481_,
    new_n32482_, new_n32484_, new_n32485_, new_n32487_, new_n32488_,
    new_n32490_, new_n32491_, new_n32493_, new_n32494_, new_n32496_,
    new_n32497_, new_n32499_, new_n32501_, new_n32502_, new_n32503_,
    new_n32504_, new_n32506_, new_n32507_, new_n32508_, new_n32509_,
    new_n32510_, new_n32511_, new_n32513_, new_n32514_, new_n32515_,
    new_n32516_, new_n32518_, new_n32519_, new_n32520_, new_n32521_,
    new_n32522_, new_n32523_, new_n32524_, new_n32525_, new_n32526_,
    new_n32527_, new_n32528_, new_n32529_, new_n32530_, new_n32531_,
    new_n32533_, new_n32535_, new_n32537_, new_n32539_, new_n32541_,
    new_n32543_, new_n32545_, new_n32547_, new_n32548_, new_n32549_,
    new_n32550_, new_n32551_, new_n32552_, new_n32553_, new_n32554_,
    new_n32555_, new_n32556_, new_n32557_, new_n32558_, new_n32559_,
    new_n32560_, new_n32561_, new_n32562_, new_n32564_, new_n32566_,
    new_n32568_, new_n32569_, new_n32570_, new_n32571_, new_n32573_,
    new_n32574_, new_n32575_, new_n32576_, new_n32577_, new_n32578_,
    new_n32580_, new_n32581_, new_n32582_, new_n32584_, new_n32585_,
    new_n32587_, new_n32588_, new_n32590_, new_n32591_, new_n32592_,
    new_n32593_, new_n32595_, new_n32597_, new_n32599_, new_n32600_,
    new_n32602_, new_n32604_, new_n32606_, new_n32608_, new_n32609_,
    new_n32611_, new_n32612_, new_n32614_, new_n32615_, new_n32616_,
    new_n32618_, new_n32619_, new_n32621_, new_n32622_, new_n32624_,
    new_n32625_, new_n32626_, new_n32628_, new_n32630_, new_n32631_,
    new_n32632_, new_n32633_, new_n32634_, new_n32635_, new_n32637_,
    new_n32639_, new_n32641_, new_n32643_, new_n32644_, new_n32646_,
    new_n32647_, new_n32649_, new_n32650_, new_n32652_, new_n32653_,
    new_n32655_, new_n32656_, new_n32657_, new_n32658_, new_n32660_,
    new_n32662_, new_n32664_, new_n32666_, new_n32668_, new_n32670_,
    new_n32672_, new_n32673_, new_n32675_, new_n32676_, new_n32678_,
    new_n32679_, new_n32681_, new_n32683_, new_n32685_, new_n32686_,
    new_n32688_, new_n32689_, new_n32691_, new_n32693_, new_n32695_,
    new_n32697_, new_n32698_, new_n32700_, new_n32701_, new_n32703_,
    new_n32705_, new_n32707_, new_n32708_, new_n32710_, new_n32712_,
    new_n32714_, new_n32716_, new_n32718_, new_n32720_, new_n32722_,
    new_n32723_, new_n32725_, new_n32727_, new_n32728_, new_n32730_,
    new_n32732_, new_n32734_, new_n32736_, new_n32738_, new_n32740_,
    new_n32741_, new_n32743_, new_n32745_, new_n32747_, new_n32748_,
    new_n32750_, new_n32751_, new_n32753_, new_n32754_, new_n32756_,
    new_n32758_, new_n32760_, new_n32762_, new_n32764_, new_n32766_,
    new_n32768_, new_n32770_, new_n32772_, new_n32773_, new_n32775_,
    new_n32777_, new_n32779_, new_n32781_, new_n32782_, new_n32784_,
    new_n32785_, new_n32787_, new_n32789_, new_n32791_, new_n32792_,
    new_n32794_, new_n32795_, new_n32797_, new_n32798_, new_n32800_,
    new_n32801_, new_n32803_, new_n32804_, new_n32806_, new_n32807_,
    new_n32809_, new_n32811_, new_n32812_, new_n32814_, new_n32815_,
    new_n32817_, new_n32818_, new_n32820_, new_n32822_, new_n32823_,
    new_n32825_, new_n32826_, new_n32828_, new_n32830_, new_n32832_,
    new_n32834_, new_n32835_, new_n32836_, new_n32838_, new_n32839_,
    new_n32841_, new_n32842_, new_n32844_, new_n32846_, new_n32848_,
    new_n32849_, new_n32851_, new_n32852_, new_n32854_, new_n32855_,
    new_n32857_, new_n32858_, new_n32860_, new_n32862_, new_n32863_,
    new_n32865_, new_n32866_, new_n32868_, new_n32869_, new_n32871_,
    new_n32872_, new_n32874_, new_n32876_, new_n32878_, new_n32880_,
    new_n32881_, new_n32883_, new_n32884_, new_n32886_, new_n32888_,
    new_n32890_, new_n32892_, new_n32894_, new_n32896_, new_n32898_,
    new_n32899_, new_n32901_, new_n32903_, new_n32905_, new_n32907_,
    new_n32909_, new_n32911_, new_n32913_, new_n32915_, new_n32917_,
    new_n32919_, new_n32921_, new_n32923_, new_n32925_, new_n32927_,
    new_n32928_, new_n32930_, new_n32931_, new_n32933_, new_n32935_,
    new_n32937_, new_n32938_, new_n32939_, new_n32940_, new_n32941_,
    new_n32942_, new_n32943_, new_n32944_, new_n32945_, new_n32946_,
    new_n32947_, new_n32948_, new_n32949_, new_n32950_, new_n32951_,
    new_n32952_, new_n32953_, new_n32954_, new_n32955_, new_n32956_,
    new_n32958_, new_n32960_, new_n32961_, new_n32963_, new_n32965_,
    new_n32967_, new_n32969_, new_n32971_, new_n32972_, new_n32974_,
    new_n32975_, new_n32976_, new_n32977_, new_n32978_, new_n32979_,
    new_n32980_, new_n32981_, new_n32982_, new_n32983_, new_n32984_,
    new_n32985_, new_n32986_, new_n32987_, new_n32988_, new_n32989_,
    new_n32990_, new_n32991_, new_n32992_, new_n32993_, new_n32994_,
    new_n32996_, new_n32997_, new_n32998_, new_n32999_, new_n33000_,
    new_n33001_, new_n33002_, new_n33003_, new_n33004_, new_n33005_,
    new_n33006_, new_n33007_, new_n33008_, new_n33010_, new_n33011_,
    new_n33012_, new_n33013_, new_n33014_, new_n33015_, new_n33016_,
    new_n33017_, new_n33018_, new_n33019_, new_n33020_, new_n33021_,
    new_n33022_, new_n33023_, new_n33024_, new_n33025_, new_n33026_,
    new_n33027_, new_n33028_, new_n33029_, new_n33030_, new_n33031_,
    new_n33032_, new_n33034_, new_n33036_, new_n33037_, new_n33038_,
    new_n33039_, new_n33040_, new_n33041_, new_n33042_, new_n33043_,
    new_n33044_, new_n33045_, new_n33046_, new_n33048_, new_n33049_,
    new_n33050_, new_n33051_, new_n33052_, new_n33053_, new_n33054_,
    new_n33055_, new_n33056_, new_n33057_, new_n33058_, new_n33060_,
    new_n33061_, new_n33062_, new_n33063_, new_n33064_, new_n33065_,
    new_n33066_, new_n33067_, new_n33068_, new_n33069_, new_n33070_,
    new_n33072_, new_n33073_, new_n33074_, new_n33075_, new_n33076_,
    new_n33077_, new_n33078_, new_n33079_, new_n33080_, new_n33081_,
    new_n33082_, new_n33084_, new_n33085_, new_n33086_, new_n33087_,
    new_n33088_, new_n33089_, new_n33090_, new_n33092_, new_n33093_,
    new_n33094_, new_n33095_, new_n33096_, new_n33097_, new_n33098_,
    new_n33100_, new_n33101_, new_n33102_, new_n33103_, new_n33104_,
    new_n33105_, new_n33106_, new_n33108_, new_n33109_, new_n33110_,
    new_n33111_, new_n33112_, new_n33113_, new_n33114_, new_n33118_,
    new_n33119_, new_n33121_, new_n33122_, new_n33124_, new_n33125_,
    new_n33127_, new_n33128_, new_n33130_, new_n33131_, new_n33133_,
    new_n33134_, new_n33136_, new_n33137_, new_n33139_, new_n33141_,
    new_n33142_, new_n33144_, new_n33146_, new_n33148_, new_n33149_,
    new_n33151_, new_n33152_, new_n33154_, new_n33156_, new_n33157_,
    new_n33159_, new_n33160_, new_n33162_, new_n33164_, new_n33166_,
    new_n33168_, new_n33170_, new_n33172_, new_n33173_, new_n33175_,
    new_n33176_, new_n33178_, new_n33179_, new_n33181_, new_n33182_,
    new_n33183_, new_n33184_, new_n33185_, new_n33186_, new_n33187_,
    new_n33188_, new_n33189_, new_n33191_, new_n33192_, new_n33194_,
    new_n33195_, new_n33197_, new_n33198_, new_n33200_, new_n33201_,
    new_n33203_, new_n33204_, new_n33206_, new_n33207_, new_n33208_,
    new_n33209_, new_n33211_, new_n33212_, new_n33214_, new_n33215_,
    new_n33217_, new_n33218_, new_n33220_, new_n33221_, new_n33223_,
    new_n33224_, new_n33226_, new_n33227_, new_n33229_, new_n33230_,
    new_n33231_, new_n33232_, new_n33234_, new_n33236_, new_n33237_,
    new_n33239_, new_n33240_, new_n33242_, new_n33243_, new_n33245_,
    new_n33246_, new_n33247_, new_n33248_, new_n33250_, new_n33252_,
    new_n33253_, new_n33255_, new_n33257_, new_n33258_, new_n33260_,
    new_n33262_, new_n33263_, new_n33265_, new_n33266_, new_n33268_,
    new_n33269_, new_n33271_, new_n33272_, new_n33274_, new_n33275_,
    new_n33277_, new_n33279_, new_n33280_, new_n33282_, new_n33283_,
    new_n33285_, new_n33286_, new_n33288_, new_n33289_, new_n33291_,
    new_n33292_, new_n33294_, new_n33295_, new_n33297_, new_n33298_,
    new_n33300_, new_n33301_, new_n33303_, new_n33305_, new_n33306_,
    new_n33307_, new_n33309_, new_n33310_, new_n33312_, new_n33314_,
    new_n33315_, new_n33317_, new_n33319_, new_n33320_, new_n33322_,
    new_n33324_, new_n33325_, new_n33327_, new_n33328_, new_n33330_,
    new_n33331_, new_n33333_, new_n33334_, new_n33336_, new_n33337_,
    new_n33339_, new_n33340_, new_n33342_, new_n33343_, new_n33344_,
    new_n33346_, new_n33347_, new_n33349_, new_n33350_, new_n33352_,
    new_n33353_, new_n33355_, new_n33356_, new_n33358_, new_n33360_,
    new_n33361_, new_n33363_, new_n33364_, new_n33366_, new_n33368_,
    new_n33369_, new_n33371_, new_n33372_, new_n33373_, new_n33374_,
    new_n33375_, new_n33376_, new_n33377_, new_n33378_, new_n33379_,
    new_n33380_, new_n33381_, new_n33382_, new_n33383_, new_n33384_,
    new_n33385_, new_n33386_, new_n33387_, new_n33388_, new_n33389_,
    new_n33390_, new_n33391_, new_n33392_, new_n33393_, new_n33394_,
    new_n33395_, new_n33396_, new_n33397_, new_n33398_, new_n33399_,
    new_n33400_, new_n33401_, new_n33402_, new_n33403_, new_n33404_,
    new_n33405_, new_n33406_, new_n33407_, new_n33408_, new_n33409_,
    new_n33410_, new_n33411_, new_n33412_, new_n33413_, new_n33414_,
    new_n33415_, new_n33416_, new_n33417_, new_n33418_, new_n33419_,
    new_n33420_, new_n33421_, new_n33422_, new_n33423_, new_n33424_,
    new_n33425_, new_n33426_, new_n33427_, new_n33428_, new_n33429_,
    new_n33430_, new_n33431_, new_n33432_, new_n33433_, new_n33434_,
    new_n33435_, new_n33436_, new_n33437_, new_n33438_, new_n33439_,
    new_n33440_, new_n33441_, new_n33443_, new_n33444_, new_n33446_,
    new_n33448_, new_n33449_, new_n33450_, new_n33452_, new_n33454_,
    new_n33455_, new_n33457_, new_n33458_, new_n33460_, new_n33461_,
    new_n33463_, new_n33464_, new_n33466_, new_n33468_, new_n33469_,
    new_n33471_, new_n33472_, new_n33474_, new_n33475_, new_n33477_,
    new_n33478_, new_n33480_, new_n33481_, new_n33483_, new_n33484_,
    new_n33486_, new_n33487_, new_n33489_, new_n33490_, new_n33492_,
    new_n33493_, new_n33495_, new_n33496_, new_n33498_, new_n33499_,
    new_n33500_, new_n33501_, new_n33503_, new_n33504_, new_n33505_,
    new_n33506_, new_n33507_, new_n33508_, new_n33509_, new_n33510_,
    new_n33511_, new_n33512_, new_n33513_, new_n33514_, new_n33515_,
    new_n33516_, new_n33518_, new_n33519_, new_n33521_, new_n33522_,
    new_n33524_, new_n33525_, new_n33527_, new_n33528_, new_n33529_,
    new_n33530_, new_n33531_, new_n33532_, new_n33533_, new_n33534_,
    new_n33535_, new_n33536_, new_n33537_, new_n33538_, new_n33539_,
    new_n33540_, new_n33541_, new_n33542_, new_n33543_, new_n33544_,
    new_n33545_, new_n33546_, new_n33547_, new_n33548_, new_n33549_,
    new_n33550_, new_n33551_, new_n33552_, new_n33553_, new_n33554_,
    new_n33555_, new_n33556_, new_n33557_, new_n33558_, new_n33559_,
    new_n33560_, new_n33561_, new_n33562_, new_n33563_, new_n33564_,
    new_n33565_, new_n33566_, new_n33567_, new_n33568_, new_n33569_,
    new_n33570_, new_n33571_, new_n33572_, new_n33573_, new_n33574_,
    new_n33575_, new_n33576_, new_n33577_, new_n33578_, new_n33579_,
    new_n33580_, new_n33581_, new_n33582_, new_n33583_, new_n33584_,
    new_n33585_, new_n33586_, new_n33587_, new_n33588_, new_n33589_,
    new_n33590_, new_n33591_, new_n33592_, new_n33593_, new_n33594_,
    new_n33595_, new_n33596_, new_n33597_, new_n33598_, new_n33599_,
    new_n33600_, new_n33601_, new_n33602_, new_n33603_, new_n33604_,
    new_n33605_, new_n33606_, new_n33607_, new_n33608_, new_n33609_,
    new_n33610_, new_n33611_, new_n33612_, new_n33613_, new_n33614_,
    new_n33615_, new_n33616_, new_n33617_, new_n33618_, new_n33619_,
    new_n33620_, new_n33621_, new_n33622_, new_n33623_, new_n33624_,
    new_n33625_, new_n33626_, new_n33627_, new_n33628_, new_n33629_,
    new_n33630_, new_n33631_, new_n33632_, new_n33633_, new_n33634_,
    new_n33635_, new_n33636_, new_n33637_, new_n33638_, new_n33639_,
    new_n33640_, new_n33641_, new_n33642_, new_n33643_, new_n33644_,
    new_n33645_, new_n33646_, new_n33647_, new_n33648_, new_n33649_,
    new_n33650_, new_n33651_, new_n33652_, new_n33653_, new_n33654_,
    new_n33655_, new_n33656_, new_n33657_, new_n33658_, new_n33659_,
    new_n33660_, new_n33661_, new_n33662_, new_n33663_, new_n33664_,
    new_n33665_, new_n33666_, new_n33667_, new_n33668_, new_n33669_,
    new_n33670_, new_n33671_, new_n33672_, new_n33673_, new_n33674_,
    new_n33675_, new_n33676_, new_n33677_, new_n33678_, new_n33679_,
    new_n33680_, new_n33681_, new_n33682_, new_n33683_, new_n33684_,
    new_n33685_, new_n33686_, new_n33687_, new_n33688_, new_n33689_,
    new_n33690_, new_n33691_, new_n33692_, new_n33693_, new_n33694_,
    new_n33695_, new_n33696_, new_n33697_, new_n33698_, new_n33699_,
    new_n33700_, new_n33701_, new_n33702_, new_n33703_, new_n33704_,
    new_n33705_, new_n33706_, new_n33707_, new_n33708_, new_n33709_,
    new_n33710_, new_n33711_, new_n33712_, new_n33713_, new_n33714_,
    new_n33715_, new_n33716_, new_n33717_, new_n33718_, new_n33719_,
    new_n33720_, new_n33721_, new_n33722_, new_n33723_, new_n33724_,
    new_n33725_, new_n33726_, new_n33727_, new_n33728_, new_n33729_,
    new_n33730_, new_n33731_, new_n33732_, new_n33733_, new_n33734_,
    new_n33735_, new_n33736_, new_n33737_, new_n33738_, new_n33739_,
    new_n33740_, new_n33741_, new_n33742_, new_n33743_, new_n33744_,
    new_n33745_, new_n33746_, new_n33747_, new_n33748_, new_n33749_,
    new_n33750_, new_n33751_, new_n33752_, new_n33753_, new_n33754_,
    new_n33755_, new_n33756_, new_n33757_, new_n33758_, new_n33759_,
    new_n33760_, new_n33761_, new_n33762_, new_n33763_, new_n33764_,
    new_n33765_, new_n33766_, new_n33767_, new_n33768_, new_n33769_,
    new_n33770_, new_n33771_, new_n33772_, new_n33773_, new_n33774_,
    new_n33775_, new_n33776_, new_n33777_, new_n33778_, new_n33779_,
    new_n33780_, new_n33781_, new_n33782_, new_n33783_, new_n33784_,
    new_n33785_, new_n33786_, new_n33787_, new_n33788_, new_n33789_,
    new_n33790_, new_n33791_, new_n33792_, new_n33793_, new_n33794_,
    new_n33795_, new_n33796_, new_n33797_, new_n33798_, new_n33799_,
    new_n33800_, new_n33801_, new_n33802_, new_n33803_, new_n33804_,
    new_n33805_, new_n33806_, new_n33807_, new_n33808_, new_n33809_,
    new_n33810_, new_n33811_, new_n33812_, new_n33813_, new_n33814_,
    new_n33815_, new_n33816_, new_n33817_, new_n33818_, new_n33819_,
    new_n33820_, new_n33821_, new_n33822_, new_n33823_, new_n33824_,
    new_n33825_, new_n33826_, new_n33827_, new_n33828_, new_n33829_,
    new_n33830_, new_n33831_, new_n33832_, new_n33833_, new_n33834_,
    new_n33835_, new_n33836_, new_n33837_, new_n33838_, new_n33839_,
    new_n33840_, new_n33841_, new_n33842_, new_n33843_, new_n33844_,
    new_n33845_, new_n33846_, new_n33847_, new_n33848_, new_n33849_,
    new_n33850_, new_n33851_, new_n33852_, new_n33853_, new_n33854_,
    new_n33855_, new_n33856_, new_n33857_, new_n33858_, new_n33859_,
    new_n33860_, new_n33861_, new_n33862_, new_n33863_, new_n33864_,
    new_n33865_, new_n33866_, new_n33867_, new_n33868_, new_n33869_,
    new_n33870_, new_n33871_, new_n33872_, new_n33873_, new_n33874_,
    new_n33875_, new_n33876_, new_n33877_, new_n33878_, new_n33879_,
    new_n33880_, new_n33881_, new_n33882_, new_n33883_, new_n33884_,
    new_n33885_, new_n33886_, new_n33887_, new_n33888_, new_n33889_,
    new_n33890_, new_n33891_, new_n33892_, new_n33893_, new_n33894_,
    new_n33895_, new_n33896_, new_n33897_, new_n33898_, new_n33899_,
    new_n33900_, new_n33901_, new_n33902_, new_n33903_, new_n33904_,
    new_n33905_, new_n33906_, new_n33907_, new_n33908_, new_n33909_,
    new_n33910_, new_n33911_, new_n33912_, new_n33913_, new_n33914_,
    new_n33915_, new_n33916_, new_n33917_, new_n33918_, new_n33919_,
    new_n33920_, new_n33921_, new_n33922_, new_n33923_, new_n33924_,
    new_n33925_, new_n33926_, new_n33927_, new_n33928_, new_n33929_,
    new_n33930_, new_n33931_, new_n33932_, new_n33933_, new_n33934_,
    new_n33935_, new_n33936_, new_n33937_, new_n33938_, new_n33939_,
    new_n33940_, new_n33941_, new_n33942_, new_n33943_, new_n33944_,
    new_n33945_, new_n33946_, new_n33947_, new_n33948_, new_n33949_,
    new_n33950_, new_n33951_, new_n33952_, new_n33953_, new_n33954_,
    new_n33955_, new_n33956_, new_n33957_, new_n33958_, new_n33959_,
    new_n33960_, new_n33961_, new_n33962_, new_n33963_, new_n33964_,
    new_n33965_, new_n33966_, new_n33967_, new_n33968_, new_n33969_,
    new_n33970_, new_n33971_, new_n33972_, new_n33973_, new_n33974_,
    new_n33975_, new_n33976_, new_n33977_, new_n33978_, new_n33979_,
    new_n33980_, new_n33981_, new_n33982_, new_n33983_, new_n33984_,
    new_n33985_, new_n33986_, new_n33987_, new_n33988_, new_n33989_,
    new_n33990_, new_n33991_, new_n33992_, new_n33993_, new_n33994_,
    new_n33995_, new_n33996_, new_n33997_, new_n33998_, new_n33999_,
    new_n34000_, new_n34001_, new_n34002_, new_n34003_, new_n34004_,
    new_n34005_, new_n34006_, new_n34007_, new_n34008_, new_n34009_,
    new_n34010_, new_n34011_, new_n34012_, new_n34013_, new_n34014_,
    new_n34015_, new_n34016_, new_n34017_, new_n34018_, new_n34019_,
    new_n34020_, new_n34021_, new_n34022_, new_n34023_, new_n34024_,
    new_n34025_, new_n34026_, new_n34027_, new_n34028_, new_n34029_,
    new_n34030_, new_n34031_, new_n34032_, new_n34033_, new_n34034_,
    new_n34035_, new_n34036_, new_n34037_, new_n34038_, new_n34039_,
    new_n34040_, new_n34041_, new_n34042_, new_n34043_, new_n34044_,
    new_n34045_, new_n34046_, new_n34047_, new_n34048_, new_n34049_,
    new_n34050_, new_n34051_, new_n34052_, new_n34053_, new_n34054_,
    new_n34055_, new_n34056_, new_n34057_, new_n34058_, new_n34059_,
    new_n34060_, new_n34061_, new_n34062_, new_n34063_, new_n34064_,
    new_n34065_, new_n34066_, new_n34067_, new_n34068_, new_n34069_,
    new_n34070_, new_n34071_, new_n34072_, new_n34073_, new_n34074_,
    new_n34075_, new_n34076_, new_n34077_, new_n34078_, new_n34079_,
    new_n34080_, new_n34081_, new_n34082_, new_n34083_, new_n34084_,
    new_n34085_, new_n34086_, new_n34087_, new_n34088_, new_n34089_,
    new_n34090_, new_n34091_, new_n34092_, new_n34093_, new_n34094_,
    new_n34095_, new_n34096_, new_n34097_, new_n34098_, new_n34099_,
    new_n34101_, new_n34102_, new_n34103_, new_n34104_, new_n34106_,
    new_n34107_, new_n34108_, new_n34110_, new_n34111_, new_n34112_,
    new_n34114_, new_n34115_, new_n34116_, new_n34118_, new_n34119_,
    new_n34120_, new_n34121_, new_n34123_, new_n34124_, new_n34126_,
    new_n34127_, new_n34128_, new_n34130_, new_n34131_, new_n34133_,
    new_n34134_, new_n34135_, new_n34136_, new_n34137_, new_n34139_,
    new_n34140_, new_n34141_, new_n34142_, new_n34143_, new_n34144_,
    new_n34145_, new_n34147_, new_n34148_, new_n34150_, new_n34151_,
    new_n34152_, new_n34153_, new_n34154_, new_n34156_, new_n34157_,
    new_n34159_, new_n34160_, new_n34161_, new_n34163_, new_n34164_,
    new_n34165_, new_n34167_, new_n34168_, new_n34170_, new_n34171_,
    new_n34173_, new_n34174_, new_n34176_, new_n34177_, new_n34179_,
    new_n34180_, new_n34182_, new_n34183_, new_n34185_, new_n34186_,
    new_n34187_, new_n34189_, new_n34190_, new_n34192_, new_n34193_,
    new_n34194_, new_n34196_, new_n34197_, new_n34198_, new_n34200_,
    new_n34201_, new_n34203_, new_n34204_, new_n34206_, new_n34207_,
    new_n34209_, new_n34210_, new_n34212_, new_n34213_, new_n34215_,
    new_n34216_, new_n34218_, new_n34219_, new_n34220_, new_n34221_,
    new_n34223_, new_n34224_, new_n34225_, new_n34226_, new_n34228_,
    new_n34229_, new_n34230_, new_n34232_, new_n34233_, new_n34235_,
    new_n34236_, new_n34238_, new_n34239_, new_n34241_, new_n34242_,
    new_n34244_, new_n34245_, new_n34247_, new_n34248_, new_n34250_,
    new_n34251_, new_n34253_, new_n34254_, new_n34256_, new_n34257_,
    new_n34259_, new_n34260_, new_n34262_, new_n34263_, new_n34265_,
    new_n34266_, new_n34268_, new_n34269_, new_n34271_, new_n34272_,
    new_n34274_, new_n34275_, new_n34277_, new_n34278_, new_n34280_,
    new_n34281_, new_n34283_, new_n34284_, new_n34286_, new_n34287_,
    new_n34289_, new_n34290_, new_n34292_, new_n34293_, new_n34295_,
    new_n34296_, new_n34298_, new_n34299_, new_n34301_, new_n34302_,
    new_n34304_, new_n34305_, new_n34307_, new_n34308_, new_n34310_,
    new_n34311_, new_n34313_, new_n34314_, new_n34316_, new_n34317_,
    new_n34319_, new_n34320_, new_n34322_, new_n34323_, new_n34325_,
    new_n34326_, new_n34328_, new_n34329_, new_n34331_, new_n34332_,
    new_n34333_, new_n34334_, new_n34335_, new_n34337_, new_n34338_,
    new_n34340_, new_n34341_, new_n34343_, new_n34344_, new_n34346_,
    new_n34347_, new_n34348_, new_n34349_, new_n34350_, new_n34351_,
    new_n34352_, new_n34353_, new_n34354_, new_n34355_, new_n34356_,
    new_n34357_, new_n34358_, new_n34359_, new_n34360_, new_n34361_,
    new_n34362_, new_n34363_, new_n34364_, new_n34365_, new_n34366_,
    new_n34367_, new_n34368_, new_n34369_, new_n34370_, new_n34371_,
    new_n34372_, new_n34373_, new_n34374_, new_n34375_, new_n34376_,
    new_n34377_, new_n34378_, new_n34379_, new_n34380_, new_n34381_,
    new_n34382_, new_n34383_, new_n34384_, new_n34386_, new_n34387_,
    new_n34388_, new_n34389_, new_n34390_, new_n34391_, new_n34392_,
    new_n34393_, new_n34394_, new_n34395_, new_n34396_, new_n34397_,
    new_n34398_, new_n34399_, new_n34400_, new_n34401_, new_n34402_,
    new_n34403_, new_n34404_, new_n34405_, new_n34406_, new_n34407_,
    new_n34408_, new_n34409_, new_n34410_, new_n34411_, new_n34412_,
    new_n34413_, new_n34414_, new_n34415_, new_n34417_, new_n34418_,
    new_n34420_, new_n34421_, new_n34422_, new_n34423_, new_n34424_,
    new_n34425_, new_n34426_, new_n34427_, new_n34428_, new_n34429_,
    new_n34430_, new_n34431_, new_n34432_, new_n34433_, new_n34434_,
    new_n34435_, new_n34436_, new_n34437_, new_n34438_, new_n34439_,
    new_n34440_, new_n34441_, new_n34443_, new_n34444_, new_n34445_,
    new_n34446_, new_n34447_, new_n34448_, new_n34449_, new_n34450_,
    new_n34451_, new_n34452_, new_n34453_, new_n34454_, new_n34455_,
    new_n34456_, new_n34457_, new_n34458_, new_n34459_, new_n34460_,
    new_n34461_, new_n34462_, new_n34463_, new_n34464_, new_n34465_,
    new_n34467_, new_n34468_, new_n34469_, new_n34470_, new_n34471_,
    new_n34472_, new_n34473_, new_n34474_, new_n34475_, new_n34476_,
    new_n34477_, new_n34478_, new_n34479_, new_n34480_, new_n34481_,
    new_n34482_, new_n34483_, new_n34484_, new_n34485_, new_n34486_,
    new_n34487_, new_n34488_, new_n34490_, new_n34491_, new_n34493_,
    new_n34494_, new_n34495_, new_n34496_, new_n34497_, new_n34498_,
    new_n34499_, new_n34500_, new_n34501_, new_n34502_, new_n34503_,
    new_n34504_, new_n34505_, new_n34506_, new_n34507_, new_n34508_,
    new_n34509_, new_n34511_, new_n34512_, new_n34513_, new_n34514_,
    new_n34515_, new_n34516_, new_n34517_, new_n34518_, new_n34519_,
    new_n34520_, new_n34521_, new_n34522_, new_n34523_, new_n34524_,
    new_n34525_, new_n34526_, new_n34528_, new_n34529_, new_n34530_,
    new_n34531_, new_n34532_, new_n34533_, new_n34534_, new_n34535_,
    new_n34536_, new_n34537_, new_n34538_, new_n34539_, new_n34540_,
    new_n34541_, new_n34542_, new_n34543_, new_n34544_, new_n34545_,
    new_n34546_, new_n34547_, new_n34548_, new_n34549_, new_n34551_,
    new_n34552_, new_n34553_, new_n34554_, new_n34555_, new_n34556_,
    new_n34557_, new_n34558_, new_n34559_, new_n34560_, new_n34561_,
    new_n34562_, new_n34563_, new_n34564_, new_n34565_, new_n34566_,
    new_n34567_, new_n34568_, new_n34569_, new_n34570_, new_n34571_,
    new_n34573_, new_n34574_, new_n34575_, new_n34576_, new_n34577_,
    new_n34578_, new_n34579_, new_n34580_, new_n34581_, new_n34582_,
    new_n34583_, new_n34584_, new_n34585_, new_n34586_, new_n34587_,
    new_n34588_, new_n34589_, new_n34590_, new_n34591_, new_n34592_,
    new_n34593_, new_n34594_, new_n34595_, new_n34596_, new_n34597_,
    new_n34599_, new_n34600_, new_n34601_, new_n34602_, new_n34603_,
    new_n34604_, new_n34605_, new_n34606_, new_n34607_, new_n34608_,
    new_n34609_, new_n34610_, new_n34611_, new_n34612_, new_n34613_,
    new_n34614_, new_n34615_, new_n34616_, new_n34617_, new_n34618_,
    new_n34619_, new_n34621_, new_n34622_, new_n34623_, new_n34624_,
    new_n34625_, new_n34626_, new_n34627_, new_n34628_, new_n34629_,
    new_n34630_, new_n34631_, new_n34632_, new_n34633_, new_n34634_,
    new_n34635_, new_n34636_, new_n34637_, new_n34638_, new_n34639_,
    new_n34640_, new_n34641_, new_n34643_, new_n34644_, new_n34645_,
    new_n34646_, new_n34647_, new_n34648_, new_n34649_, new_n34650_,
    new_n34651_, new_n34652_, new_n34653_, new_n34654_, new_n34655_,
    new_n34656_, new_n34657_, new_n34658_, new_n34660_, new_n34661_,
    new_n34662_, new_n34663_, new_n34664_, new_n34665_, new_n34666_,
    new_n34667_, new_n34668_, new_n34669_, new_n34670_, new_n34671_,
    new_n34672_, new_n34673_, new_n34674_, new_n34675_, new_n34677_,
    new_n34678_, new_n34679_, new_n34680_, new_n34681_, new_n34682_,
    new_n34683_, new_n34684_, new_n34685_, new_n34686_, new_n34687_,
    new_n34688_, new_n34689_, new_n34690_, new_n34691_, new_n34692_,
    new_n34693_, new_n34694_, new_n34695_, new_n34696_, new_n34697_,
    new_n34699_, new_n34700_, new_n34702_, new_n34703_, new_n34705_,
    new_n34706_, new_n34707_, new_n34708_, new_n34709_, new_n34710_,
    new_n34711_, new_n34712_, new_n34713_, new_n34714_, new_n34715_,
    new_n34716_, new_n34717_, new_n34718_, new_n34719_, new_n34720_,
    new_n34722_, new_n34723_, new_n34724_, new_n34726_, new_n34728_,
    new_n34729_, new_n34730_, new_n34731_, new_n34732_, new_n34733_,
    new_n34734_, new_n34735_, new_n34736_, new_n34737_, new_n34738_,
    new_n34739_, new_n34740_, new_n34741_, new_n34742_, new_n34743_,
    new_n34744_, new_n34745_, new_n34746_, new_n34747_, new_n34748_,
    new_n34749_, new_n34750_, new_n34751_, new_n34753_, new_n34754_,
    new_n34756_, new_n34757_, new_n34759_, new_n34760_, new_n34762_,
    new_n34763_, new_n34764_, new_n34765_, new_n34766_, new_n34767_,
    new_n34768_, new_n34769_, new_n34770_, new_n34771_, new_n34772_,
    new_n34773_, new_n34774_, new_n34775_, new_n34776_, new_n34777_,
    new_n34778_, new_n34779_, new_n34781_, new_n34782_, new_n34784_,
    new_n34785_, new_n34787_, new_n34788_, new_n34789_, new_n34790_,
    new_n34791_, new_n34792_, new_n34793_, new_n34794_, new_n34795_,
    new_n34796_, new_n34797_, new_n34798_, new_n34799_, new_n34800_,
    new_n34801_, new_n34802_, new_n34803_, new_n34805_, new_n34806_,
    new_n34808_, new_n34809_, new_n34810_, new_n34812_, new_n34813_,
    new_n34815_, new_n34816_, new_n34818_, new_n34819_, new_n34820_,
    new_n34822_, new_n34823_, new_n34825_, new_n34826_, new_n34828_,
    new_n34829_, new_n34831_, new_n34832_, new_n34834_, new_n34835_,
    new_n34837_, new_n34838_, new_n34840_, new_n34841_, new_n34843_,
    new_n34844_, new_n34846_, new_n34847_, new_n34849_, new_n34850_,
    new_n34851_, new_n34852_, new_n34853_, new_n34854_, new_n34855_,
    new_n34856_, new_n34857_, new_n34858_, new_n34859_, new_n34860_,
    new_n34861_, new_n34862_, new_n34863_, new_n34864_, new_n34865_,
    new_n34866_, new_n34867_, new_n34868_, new_n34869_, new_n34870_,
    new_n34872_, new_n34873_, new_n34874_, new_n34875_, new_n34876_,
    new_n34877_, new_n34878_, new_n34879_, new_n34880_, new_n34881_,
    new_n34882_, new_n34883_, new_n34884_, new_n34885_, new_n34886_,
    new_n34887_, new_n34888_, new_n34889_, new_n34890_, new_n34891_,
    new_n34892_, new_n34893_, new_n34894_, new_n34896_, new_n34897_,
    new_n34899_, new_n34900_, new_n34902_, new_n34903_, new_n34904_,
    new_n34905_, new_n34906_, new_n34907_, new_n34908_, new_n34909_,
    new_n34910_, new_n34911_, new_n34912_, new_n34913_, new_n34914_,
    new_n34915_, new_n34916_, new_n34917_, new_n34918_, new_n34919_,
    new_n34921_, new_n34922_, new_n34923_, new_n34924_, new_n34925_,
    new_n34926_, new_n34927_, new_n34928_, new_n34929_, new_n34930_,
    new_n34931_, new_n34932_, new_n34933_, new_n34934_, new_n34935_,
    new_n34936_, new_n34937_, new_n34939_, new_n34940_, new_n34941_,
    new_n34942_, new_n34943_, new_n34944_, new_n34945_, new_n34946_,
    new_n34947_, new_n34948_, new_n34949_, new_n34950_, new_n34951_,
    new_n34952_, new_n34953_, new_n34954_, new_n34955_, new_n34956_,
    new_n34957_, new_n34959_, new_n34960_, new_n34961_, new_n34962_,
    new_n34963_, new_n34964_, new_n34965_, new_n34966_, new_n34967_,
    new_n34968_, new_n34969_, new_n34970_, new_n34971_, new_n34972_,
    new_n34973_, new_n34974_, new_n34975_, new_n34976_, new_n34978_,
    new_n34979_, new_n34981_, new_n34982_, new_n34983_, new_n34984_,
    new_n34985_, new_n34986_, new_n34987_, new_n34988_, new_n34989_,
    new_n34990_, new_n34991_, new_n34992_, new_n34993_, new_n34994_,
    new_n34995_, new_n34996_, new_n34997_, new_n34998_, new_n34999_,
    new_n35000_, new_n35002_, new_n35003_, new_n35004_, new_n35005_,
    new_n35006_, new_n35007_, new_n35008_, new_n35009_, new_n35010_,
    new_n35011_, new_n35012_, new_n35013_, new_n35014_, new_n35015_,
    new_n35016_, new_n35017_, new_n35018_, new_n35020_, new_n35021_,
    new_n35022_, new_n35023_, new_n35024_, new_n35025_, new_n35026_,
    new_n35027_, new_n35028_, new_n35029_, new_n35030_, new_n35031_,
    new_n35032_, new_n35033_, new_n35034_, new_n35035_, new_n35036_,
    new_n35037_, new_n35038_, new_n35039_, new_n35041_, new_n35042_,
    new_n35043_, new_n35044_, new_n35045_, new_n35046_, new_n35047_,
    new_n35048_, new_n35049_, new_n35050_, new_n35051_, new_n35052_,
    new_n35053_, new_n35054_, new_n35055_, new_n35056_, new_n35057_,
    new_n35059_, new_n35060_, new_n35061_, new_n35062_, new_n35063_,
    new_n35064_, new_n35065_, new_n35066_, new_n35067_, new_n35068_,
    new_n35069_, new_n35070_, new_n35071_, new_n35072_, new_n35073_,
    new_n35074_, new_n35075_, new_n35076_, new_n35078_, new_n35079_,
    new_n35080_, new_n35081_, new_n35082_, new_n35083_, new_n35084_,
    new_n35085_, new_n35086_, new_n35087_, new_n35088_, new_n35089_,
    new_n35090_, new_n35091_, new_n35092_, new_n35093_, new_n35094_,
    new_n35095_, new_n35096_, new_n35097_, new_n35098_, new_n35099_,
    new_n35100_, new_n35101_, new_n35102_, new_n35103_, new_n35104_,
    new_n35105_, new_n35106_, new_n35107_, new_n35108_, new_n35109_,
    new_n35110_, new_n35111_, new_n35112_, new_n35113_, new_n35114_,
    new_n35115_, new_n35116_, new_n35117_, new_n35118_, new_n35119_,
    new_n35120_, new_n35121_, new_n35122_, new_n35123_, new_n35124_,
    new_n35125_, new_n35126_, new_n35127_, new_n35128_, new_n35129_,
    new_n35130_, new_n35131_, new_n35132_, new_n35134_, new_n35135_,
    new_n35136_, new_n35137_, new_n35138_, new_n35139_, new_n35140_,
    new_n35141_, new_n35142_, new_n35143_, new_n35144_, new_n35145_,
    new_n35146_, new_n35147_, new_n35148_, new_n35149_, new_n35150_,
    new_n35151_, new_n35152_, new_n35153_, new_n35154_, new_n35155_,
    new_n35156_, new_n35158_, new_n35159_, new_n35161_, new_n35162_,
    new_n35164_, new_n35165_, new_n35167_, new_n35168_, new_n35170_,
    new_n35171_, new_n35173_, new_n35174_, new_n35175_, new_n35177_,
    new_n35178_, new_n35180_, new_n35181_, new_n35183_, new_n35184_,
    new_n35185_, new_n35186_, new_n35187_, new_n35188_, new_n35189_,
    new_n35190_, new_n35191_, new_n35192_, new_n35193_, new_n35195_,
    new_n35196_, new_n35198_, new_n35199_, new_n35200_, new_n35201_,
    new_n35202_, new_n35203_, new_n35204_, new_n35205_, new_n35206_,
    new_n35207_, new_n35208_, new_n35209_, new_n35210_, new_n35211_,
    new_n35212_, new_n35213_, new_n35214_, new_n35215_, new_n35216_,
    new_n35217_, new_n35219_, new_n35220_, new_n35222_, new_n35223_,
    new_n35225_, new_n35226_, new_n35228_, new_n35229_, new_n35231_,
    new_n35232_, new_n35234_, new_n35235_, new_n35237_, new_n35238_,
    new_n35239_, new_n35241_, new_n35242_, new_n35244_, new_n35245_,
    new_n35247_, new_n35248_, new_n35250_, new_n35251_, new_n35252_,
    new_n35254_, new_n35255_, new_n35257_, new_n35258_, new_n35260_,
    new_n35261_, new_n35262_, new_n35263_, new_n35264_, new_n35265_,
    new_n35266_, new_n35268_, new_n35269_, new_n35271_, new_n35272_,
    new_n35274_, new_n35275_, new_n35276_, new_n35278_, new_n35279_,
    new_n35281_, new_n35282_, new_n35284_, new_n35285_, new_n35287_,
    new_n35288_, new_n35290_, new_n35291_, new_n35293_, new_n35294_,
    new_n35296_, new_n35297_, new_n35299_, new_n35300_, new_n35302_,
    new_n35303_, new_n35305_, new_n35306_, new_n35308_, new_n35309_,
    new_n35311_, new_n35312_, new_n35313_, new_n35315_, new_n35316_,
    new_n35318_, new_n35319_, new_n35321_, new_n35322_, new_n35323_,
    new_n35324_, new_n35325_, new_n35326_, new_n35327_, new_n35328_,
    new_n35329_, new_n35330_, new_n35331_, new_n35332_, new_n35333_,
    new_n35334_, new_n35335_, new_n35336_, new_n35337_, new_n35338_,
    new_n35340_, new_n35342_, new_n35343_, new_n35345_, new_n35346_,
    new_n35348_, new_n35349_, new_n35351_, new_n35352_, new_n35353_,
    new_n35354_, new_n35355_, new_n35356_, new_n35357_, new_n35358_,
    new_n35359_, new_n35361_, new_n35362_, new_n35364_, new_n35365_,
    new_n35366_, new_n35367_, new_n35368_, new_n35370_, new_n35372_,
    new_n35373_, new_n35375_, new_n35376_, new_n35377_, new_n35378_,
    new_n35380_, new_n35381_, new_n35383_, new_n35384_, new_n35385_,
    new_n35386_, new_n35387_, new_n35388_, new_n35389_, new_n35390_,
    new_n35391_, new_n35393_, new_n35394_, new_n35395_, new_n35397_,
    new_n35398_, new_n35400_, new_n35401_, new_n35402_, new_n35403_,
    new_n35407_, new_n35410_, new_n35412_, new_n35414_, new_n35416_,
    new_n35418_, new_n35420_, new_n35422_, new_n35424_, new_n35426_,
    new_n35428_, new_n35430_, new_n35431_, new_n35432_, new_n35434_,
    new_n35437_, new_n35438_, new_n35439_, new_n35441_, new_n35442_,
    new_n35444_, new_n35446_, new_n35448_, new_n35451_, new_n35453_,
    new_n35455_, new_n35457_, new_n35459_, new_n35461_, new_n35463_,
    new_n35465_, new_n35467_, new_n35469_, new_n35471_, new_n35473_,
    new_n35475_, new_n35480_, new_n35483_, new_n35486_, new_n35487_,
    new_n35488_, new_n35489_, new_n35490_, new_n35491_, new_n35492_,
    new_n35493_, new_n35494_, new_n35495_, new_n35496_, new_n35497_,
    new_n35498_, new_n35499_, new_n35502_, new_n35503_, new_n35504_,
    new_n35505_, new_n35506_, new_n35507_, new_n35508_, new_n35509_,
    new_n35510_, new_n35511_, new_n35512_, new_n35513_, new_n35516_,
    new_n35517_, new_n35518_, new_n35519_, new_n35520_, new_n35521_,
    new_n35522_, new_n35523_, new_n35524_, new_n35525_, new_n35526_,
    new_n35527_, new_n35530_, new_n35531_, new_n35532_, new_n35533_,
    new_n35534_, new_n35535_, new_n35536_, new_n35537_, new_n35538_,
    new_n35539_, new_n35540_, new_n35541_, new_n35543_, new_n35550_,
    new_n35553_, new_n35555_, new_n35559_, new_n35561_, new_n35564_,
    new_n35566_, new_n35569_, new_n35571_, new_n35573_, new_n35575_,
    new_n35578_, new_n35580_, new_n35582_, new_n35585_, new_n35587_,
    new_n35589_, new_n35591_, new_n35592_, new_n35593_, new_n35594_,
    new_n35595_, new_n35596_, new_n35598_, new_n35600_, new_n35602_,
    new_n35604_, new_n35606_, new_n35608_, new_n35610_, new_n35612_,
    new_n35613_, new_n35614_, new_n35615_, new_n35616_, new_n35617_,
    new_n35619_, new_n35621_, new_n35623_, new_n35625_, new_n35627_,
    new_n35629_, new_n35630_, new_n35631_, new_n35632_, new_n35634_,
    new_n35636_, new_n35637_, new_n35638_, new_n35639_, new_n35640_,
    new_n35641_, new_n35643_, new_n35644_, new_n35645_, new_n35646_,
    new_n35647_, new_n35648_, new_n35650_, new_n35651_, new_n35652_,
    new_n35653_, new_n35654_, new_n35655_, new_n35657_, new_n35659_,
    new_n35661_, new_n35663_, new_n35665_, new_n35667_, new_n35669_,
    new_n35671_, new_n35673_, new_n35675_, new_n35677_, new_n35679_,
    new_n35681_, new_n35683_, new_n35685_, new_n35687_, new_n35689_,
    new_n35691_, new_n35693_, new_n35695_, new_n35697_, new_n35699_,
    new_n35701_, new_n35703_, new_n35704_, new_n35705_, new_n35706_,
    new_n35707_, new_n35708_, new_n35709_, new_n35710_, new_n35711_,
    new_n35712_, new_n35713_, new_n35715_, new_n35717_, new_n35719_,
    new_n35721_, new_n35723_, new_n35725_, new_n35727_, new_n35728_,
    new_n35730_, new_n35732_, new_n35734_, new_n35736_, new_n35738_,
    new_n35740_, new_n35742_, new_n35744_, new_n35746_, new_n35748_,
    new_n35750_, new_n35752_, new_n35754_, new_n35757_, new_n35759_,
    new_n35761_, new_n35764_, new_n35766_, new_n35768_, new_n35770_,
    new_n35772_, new_n35774_, new_n35776_, new_n35778_, new_n35780_,
    new_n35782_, new_n35784_, new_n35786_, new_n35791_;
  INV_X1     g00000(.I(pi0215), .ZN(new_n2436_));
  NOR2_X1    g00001(.A1(pi0332), .A2(pi1144), .ZN(new_n2437_));
  INV_X1     g00002(.I(new_n2437_), .ZN(new_n2438_));
  NOR2_X1    g00003(.A1(new_n2438_), .A2(new_n2436_), .ZN(new_n2439_));
  INV_X1     g00004(.I(new_n2439_), .ZN(new_n2440_));
  INV_X1     g00005(.I(pi0221), .ZN(new_n2441_));
  INV_X1     g00006(.I(pi0929), .ZN(new_n2442_));
  INV_X1     g00007(.I(pi0833), .ZN(new_n2443_));
  NOR2_X1    g00008(.A1(new_n2443_), .A2(pi0216), .ZN(new_n2444_));
  NAND2_X1   g00009(.A1(new_n2444_), .A2(new_n2442_), .ZN(new_n2445_));
  INV_X1     g00010(.I(pi1144), .ZN(new_n2446_));
  INV_X1     g00011(.I(new_n2444_), .ZN(new_n2447_));
  NAND2_X1   g00012(.A1(new_n2447_), .A2(new_n2446_), .ZN(new_n2448_));
  AOI21_X1   g00013(.A1(new_n2448_), .A2(new_n2445_), .B(pi0332), .ZN(new_n2449_));
  INV_X1     g00014(.I(new_n2449_), .ZN(new_n2450_));
  NOR2_X1    g00015(.A1(new_n2450_), .A2(new_n2441_), .ZN(new_n2451_));
  INV_X1     g00016(.I(pi0265), .ZN(new_n2452_));
  OAI21_X1   g00017(.A1(new_n2452_), .A2(pi0332), .B(pi0216), .ZN(new_n2453_));
  NAND2_X1   g00018(.A1(new_n2453_), .A2(new_n2441_), .ZN(new_n2454_));
  INV_X1     g00019(.I(pi0153), .ZN(new_n2455_));
  NOR2_X1    g00020(.A1(new_n2455_), .A2(pi0332), .ZN(new_n2456_));
  INV_X1     g00021(.I(pi0105), .ZN(new_n2457_));
  INV_X1     g00022(.I(pi0228), .ZN(new_n2458_));
  NOR2_X1    g00023(.A1(new_n2457_), .A2(new_n2458_), .ZN(new_n2459_));
  INV_X1     g00024(.I(new_n2459_), .ZN(new_n2460_));
  AOI21_X1   g00025(.A1(new_n2460_), .A2(new_n2456_), .B(pi0216), .ZN(new_n2461_));
  INV_X1     g00026(.I(pi0095), .ZN(new_n2462_));
  NOR2_X1    g00027(.A1(new_n2462_), .A2(pi0479), .ZN(new_n2463_));
  AOI21_X1   g00028(.A1(new_n2463_), .A2(pi0234), .B(pi0332), .ZN(new_n2464_));
  NAND2_X1   g00029(.A1(new_n2464_), .A2(new_n2459_), .ZN(new_n2465_));
  AOI21_X1   g00030(.A1(new_n2465_), .A2(new_n2461_), .B(new_n2454_), .ZN(new_n2466_));
  OAI21_X1   g00031(.A1(new_n2451_), .A2(new_n2466_), .B(new_n2436_), .ZN(new_n2467_));
  NAND2_X1   g00032(.A1(new_n2467_), .A2(new_n2440_), .ZN(new_n2468_));
  INV_X1     g00033(.I(pi0059), .ZN(new_n2469_));
  NOR2_X1    g00034(.A1(pi0056), .A2(pi0062), .ZN(new_n2470_));
  INV_X1     g00035(.I(new_n2470_), .ZN(new_n2471_));
  INV_X1     g00036(.I(new_n2461_), .ZN(new_n2472_));
  INV_X1     g00037(.I(new_n2464_), .ZN(new_n2473_));
  NOR2_X1    g00038(.A1(pi0083), .A2(pi0103), .ZN(new_n2474_));
  INV_X1     g00039(.I(new_n2474_), .ZN(new_n2475_));
  NOR2_X1    g00040(.A1(pi0067), .A2(pi0069), .ZN(new_n2476_));
  INV_X1     g00041(.I(pi0048), .ZN(new_n2477_));
  INV_X1     g00042(.I(pi0049), .ZN(new_n2478_));
  INV_X1     g00043(.I(pi0089), .ZN(new_n2479_));
  NAND3_X1   g00044(.A1(new_n2477_), .A2(new_n2478_), .A3(new_n2479_), .ZN(new_n2480_));
  INV_X1     g00045(.I(pi0061), .ZN(new_n2481_));
  INV_X1     g00046(.I(pi0076), .ZN(new_n2482_));
  NOR2_X1    g00047(.A1(pi0085), .A2(pi0106), .ZN(new_n2483_));
  NAND3_X1   g00048(.A1(new_n2483_), .A2(new_n2481_), .A3(new_n2482_), .ZN(new_n2484_));
  NOR2_X1    g00049(.A1(pi0045), .A2(pi0104), .ZN(new_n2485_));
  INV_X1     g00050(.I(new_n2485_), .ZN(new_n2486_));
  NOR3_X1    g00051(.A1(new_n2484_), .A2(new_n2480_), .A3(new_n2486_), .ZN(new_n2487_));
  OR2_X2     g00052(.A1(pi0068), .A2(pi0084), .Z(new_n2488_));
  OR3_X2     g00053(.A1(pi0036), .A2(pi0082), .A3(pi0111), .Z(new_n2489_));
  NOR2_X1    g00054(.A1(new_n2489_), .A2(new_n2488_), .ZN(new_n2490_));
  NOR2_X1    g00055(.A1(pi0066), .A2(pi0073), .ZN(new_n2491_));
  NAND4_X1   g00056(.A1(new_n2487_), .A2(new_n2476_), .A3(new_n2490_), .A4(new_n2491_), .ZN(new_n2492_));
  NOR2_X1    g00057(.A1(pi0065), .A2(pi0071), .ZN(new_n2493_));
  INV_X1     g00058(.I(new_n2493_), .ZN(new_n2494_));
  INV_X1     g00059(.I(pi0064), .ZN(new_n2495_));
  NOR2_X1    g00060(.A1(pi0063), .A2(pi0107), .ZN(new_n2496_));
  NAND2_X1   g00061(.A1(new_n2496_), .A2(new_n2495_), .ZN(po1049));
  NOR2_X1    g00062(.A1(po1049), .A2(new_n2494_), .ZN(new_n2498_));
  INV_X1     g00063(.I(new_n2498_), .ZN(new_n2499_));
  INV_X1     g00064(.I(pi0081), .ZN(new_n2500_));
  INV_X1     g00065(.I(pi0102), .ZN(new_n2501_));
  INV_X1     g00066(.I(pi0077), .ZN(new_n2502_));
  NOR2_X1    g00067(.A1(pi0088), .A2(pi0098), .ZN(new_n2503_));
  NAND2_X1   g00068(.A1(new_n2503_), .A2(new_n2502_), .ZN(new_n2504_));
  NOR2_X1    g00069(.A1(new_n2504_), .A2(pi0050), .ZN(new_n2505_));
  NAND3_X1   g00070(.A1(new_n2505_), .A2(new_n2500_), .A3(new_n2501_), .ZN(new_n2506_));
  NOR4_X1    g00071(.A1(new_n2492_), .A2(new_n2475_), .A3(new_n2499_), .A4(new_n2506_), .ZN(new_n2507_));
  INV_X1     g00072(.I(pi0109), .ZN(new_n2508_));
  INV_X1     g00073(.I(pi0110), .ZN(new_n2509_));
  NAND2_X1   g00074(.A1(new_n2508_), .A2(new_n2509_), .ZN(new_n2510_));
  INV_X1     g00075(.I(pi0046), .ZN(new_n2511_));
  NOR2_X1    g00076(.A1(pi0097), .A2(pi0108), .ZN(new_n2512_));
  NAND2_X1   g00077(.A1(new_n2512_), .A2(new_n2511_), .ZN(new_n2513_));
  INV_X1     g00078(.I(pi0094), .ZN(new_n2514_));
  NOR3_X1    g00079(.A1(pi0053), .A2(pi0060), .A3(pi0086), .ZN(new_n2515_));
  NAND2_X1   g00080(.A1(new_n2515_), .A2(new_n2514_), .ZN(new_n2516_));
  NOR2_X1    g00081(.A1(pi0047), .A2(pi0091), .ZN(new_n2517_));
  INV_X1     g00082(.I(new_n2517_), .ZN(new_n2518_));
  NOR4_X1    g00083(.A1(new_n2516_), .A2(new_n2510_), .A3(new_n2513_), .A4(new_n2518_), .ZN(new_n2519_));
  NOR2_X1    g00084(.A1(pi0058), .A2(pi0090), .ZN(new_n2520_));
  NOR2_X1    g00085(.A1(pi0035), .A2(pi0093), .ZN(new_n2521_));
  NAND2_X1   g00086(.A1(new_n2520_), .A2(new_n2521_), .ZN(new_n2522_));
  NOR2_X1    g00087(.A1(new_n2522_), .A2(pi0070), .ZN(new_n2523_));
  NOR2_X1    g00088(.A1(pi0040), .A2(pi0072), .ZN(new_n2524_));
  NOR2_X1    g00089(.A1(pi0032), .A2(pi0095), .ZN(new_n2525_));
  NAND2_X1   g00090(.A1(new_n2524_), .A2(new_n2525_), .ZN(new_n2526_));
  NOR2_X1    g00091(.A1(pi0051), .A2(pi0096), .ZN(new_n2527_));
  INV_X1     g00092(.I(new_n2527_), .ZN(new_n2528_));
  NOR2_X1    g00093(.A1(new_n2526_), .A2(new_n2528_), .ZN(new_n2529_));
  NAND4_X1   g00094(.A1(new_n2507_), .A2(new_n2519_), .A3(new_n2523_), .A4(new_n2529_), .ZN(new_n2530_));
  INV_X1     g00095(.I(new_n2530_), .ZN(new_n2531_));
  NOR2_X1    g00096(.A1(new_n2531_), .A2(pi0234), .ZN(new_n2532_));
  NOR2_X1    g00097(.A1(pi0032), .A2(pi0040), .ZN(new_n2533_));
  INV_X1     g00098(.I(new_n2533_), .ZN(new_n2534_));
  NOR2_X1    g00099(.A1(new_n2534_), .A2(pi0095), .ZN(new_n2535_));
  INV_X1     g00100(.I(new_n2535_), .ZN(new_n2536_));
  INV_X1     g00101(.I(new_n2521_), .ZN(new_n2537_));
  NOR3_X1    g00102(.A1(pi0048), .A2(pi0049), .A3(pi0089), .ZN(new_n2538_));
  NOR4_X1    g00103(.A1(pi0061), .A2(pi0076), .A3(pi0085), .A4(pi0106), .ZN(new_n2539_));
  NAND3_X1   g00104(.A1(new_n2539_), .A2(new_n2538_), .A3(new_n2485_), .ZN(new_n2540_));
  NOR2_X1    g00105(.A1(pi0068), .A2(pi0084), .ZN(new_n2541_));
  NOR3_X1    g00106(.A1(pi0036), .A2(pi0082), .A3(pi0111), .ZN(new_n2542_));
  NAND2_X1   g00107(.A1(new_n2542_), .A2(new_n2541_), .ZN(new_n2543_));
  NOR2_X1    g00108(.A1(new_n2540_), .A2(new_n2543_), .ZN(new_n2544_));
  NAND4_X1   g00109(.A1(new_n2544_), .A2(new_n2474_), .A3(new_n2476_), .A4(new_n2491_), .ZN(new_n2545_));
  INV_X1     g00110(.I(new_n2519_), .ZN(new_n2546_));
  NOR4_X1    g00111(.A1(new_n2545_), .A2(new_n2499_), .A3(new_n2506_), .A4(new_n2546_), .ZN(new_n2547_));
  NAND2_X1   g00112(.A1(new_n2547_), .A2(new_n2520_), .ZN(new_n2548_));
  NOR2_X1    g00113(.A1(pi0072), .A2(pi0096), .ZN(new_n2549_));
  NOR2_X1    g00114(.A1(pi0051), .A2(pi0070), .ZN(new_n2550_));
  NAND2_X1   g00115(.A1(new_n2549_), .A2(new_n2550_), .ZN(new_n2551_));
  NOR3_X1    g00116(.A1(new_n2548_), .A2(new_n2537_), .A3(new_n2551_), .ZN(new_n2552_));
  INV_X1     g00117(.I(new_n2552_), .ZN(new_n2553_));
  NOR2_X1    g00118(.A1(new_n2553_), .A2(new_n2536_), .ZN(new_n2554_));
  NOR2_X1    g00119(.A1(new_n2554_), .A2(new_n2463_), .ZN(new_n2555_));
  AOI21_X1   g00120(.A1(new_n2555_), .A2(pi0234), .B(new_n2532_), .ZN(new_n2556_));
  AOI21_X1   g00121(.A1(new_n2556_), .A2(pi0137), .B(new_n2473_), .ZN(new_n2557_));
  NOR2_X1    g00122(.A1(pi0215), .A2(pi0221), .ZN(new_n2558_));
  INV_X1     g00123(.I(new_n2558_), .ZN(new_n2559_));
  NOR3_X1    g00124(.A1(new_n2557_), .A2(new_n2472_), .A3(new_n2559_), .ZN(new_n2560_));
  INV_X1     g00125(.I(new_n2560_), .ZN(new_n2561_));
  NOR2_X1    g00126(.A1(pi0054), .A2(pi0074), .ZN(new_n2562_));
  INV_X1     g00127(.I(new_n2562_), .ZN(new_n2563_));
  NOR2_X1    g00128(.A1(pi0075), .A2(pi0087), .ZN(new_n2564_));
  INV_X1     g00129(.I(new_n2564_), .ZN(new_n2565_));
  NOR2_X1    g00130(.A1(new_n2565_), .A2(pi0092), .ZN(new_n2566_));
  INV_X1     g00131(.I(new_n2566_), .ZN(new_n2567_));
  NOR2_X1    g00132(.A1(new_n2567_), .A2(new_n2563_), .ZN(new_n2568_));
  INV_X1     g00133(.I(new_n2568_), .ZN(new_n2569_));
  NOR2_X1    g00134(.A1(new_n2569_), .A2(pi0055), .ZN(new_n2570_));
  INV_X1     g00135(.I(new_n2570_), .ZN(new_n2571_));
  NOR2_X1    g00136(.A1(pi0038), .A2(pi0039), .ZN(new_n2572_));
  INV_X1     g00137(.I(new_n2572_), .ZN(new_n2573_));
  NOR2_X1    g00138(.A1(new_n2573_), .A2(pi0100), .ZN(new_n2574_));
  INV_X1     g00139(.I(new_n2574_), .ZN(new_n2575_));
  NOR2_X1    g00140(.A1(new_n2571_), .A2(new_n2575_), .ZN(new_n2576_));
  INV_X1     g00141(.I(new_n2576_), .ZN(new_n2577_));
  NOR3_X1    g00142(.A1(new_n2561_), .A2(new_n2471_), .A3(new_n2577_), .ZN(new_n2578_));
  NAND2_X1   g00143(.A1(new_n2578_), .A2(new_n2469_), .ZN(new_n2579_));
  NAND2_X1   g00144(.A1(new_n2579_), .A2(new_n2468_), .ZN(new_n2580_));
  NAND2_X1   g00145(.A1(new_n2580_), .A2(pi0057), .ZN(new_n2581_));
  INV_X1     g00146(.I(pi0057), .ZN(new_n2582_));
  NAND2_X1   g00147(.A1(new_n2468_), .A2(pi0059), .ZN(new_n2583_));
  OAI21_X1   g00148(.A1(new_n2578_), .A2(new_n2583_), .B(new_n2582_), .ZN(new_n2584_));
  NOR2_X1    g00149(.A1(new_n2449_), .A2(new_n2441_), .ZN(new_n2585_));
  INV_X1     g00150(.I(new_n2585_), .ZN(new_n2586_));
  INV_X1     g00151(.I(new_n2554_), .ZN(new_n2587_));
  NOR4_X1    g00152(.A1(new_n2587_), .A2(pi0137), .A3(pi0153), .A4(pi0332), .ZN(new_n2588_));
  INV_X1     g00153(.I(new_n2588_), .ZN(new_n2589_));
  NAND2_X1   g00154(.A1(new_n2531_), .A2(pi0137), .ZN(new_n2590_));
  AOI21_X1   g00155(.A1(new_n2590_), .A2(new_n2456_), .B(pi0228), .ZN(new_n2591_));
  NOR2_X1    g00156(.A1(new_n2456_), .A2(pi0105), .ZN(new_n2592_));
  INV_X1     g00157(.I(new_n2592_), .ZN(new_n2593_));
  OAI21_X1   g00158(.A1(new_n2557_), .A2(new_n2457_), .B(new_n2593_), .ZN(new_n2594_));
  AOI22_X1   g00159(.A1(new_n2594_), .A2(pi0228), .B1(new_n2589_), .B2(new_n2591_), .ZN(new_n2595_));
  OAI21_X1   g00160(.A1(new_n2595_), .A2(pi0216), .B(new_n2453_), .ZN(new_n2596_));
  AOI21_X1   g00161(.A1(new_n2596_), .A2(new_n2441_), .B(pi0215), .ZN(new_n2597_));
  AOI21_X1   g00162(.A1(new_n2597_), .A2(new_n2586_), .B(new_n2439_), .ZN(new_n2598_));
  NOR2_X1    g00163(.A1(new_n2468_), .A2(new_n2576_), .ZN(new_n2599_));
  AOI21_X1   g00164(.A1(new_n2598_), .A2(new_n2576_), .B(new_n2599_), .ZN(new_n2600_));
  AOI21_X1   g00165(.A1(new_n2600_), .A2(pi0056), .B(pi0062), .ZN(new_n2601_));
  INV_X1     g00166(.I(pi0055), .ZN(new_n2602_));
  NOR2_X1    g00167(.A1(pi0087), .A2(pi0100), .ZN(new_n2603_));
  INV_X1     g00168(.I(new_n2603_), .ZN(new_n2604_));
  NOR2_X1    g00169(.A1(pi0075), .A2(pi0092), .ZN(new_n2605_));
  INV_X1     g00170(.I(new_n2605_), .ZN(new_n2606_));
  NOR2_X1    g00171(.A1(new_n2563_), .A2(new_n2606_), .ZN(new_n2607_));
  INV_X1     g00172(.I(new_n2607_), .ZN(new_n2608_));
  NOR2_X1    g00173(.A1(new_n2608_), .A2(new_n2604_), .ZN(new_n2609_));
  INV_X1     g00174(.I(new_n2609_), .ZN(new_n2610_));
  NOR2_X1    g00175(.A1(new_n2610_), .A2(new_n2573_), .ZN(new_n2611_));
  INV_X1     g00176(.I(new_n2611_), .ZN(new_n2612_));
  AOI21_X1   g00177(.A1(new_n2468_), .A2(new_n2612_), .B(new_n2602_), .ZN(new_n2613_));
  INV_X1     g00178(.I(pi0216), .ZN(new_n2614_));
  NAND3_X1   g00179(.A1(new_n2530_), .A2(new_n2458_), .A3(new_n2456_), .ZN(new_n2615_));
  OAI21_X1   g00180(.A1(new_n2556_), .A2(pi0332), .B(pi0105), .ZN(new_n2616_));
  NAND3_X1   g00181(.A1(new_n2616_), .A2(pi0228), .A3(new_n2593_), .ZN(new_n2617_));
  NAND3_X1   g00182(.A1(new_n2617_), .A2(new_n2614_), .A3(new_n2615_), .ZN(new_n2618_));
  AOI21_X1   g00183(.A1(new_n2618_), .A2(new_n2453_), .B(pi0221), .ZN(new_n2619_));
  OAI21_X1   g00184(.A1(new_n2619_), .A2(new_n2585_), .B(new_n2436_), .ZN(new_n2620_));
  NOR2_X1    g00185(.A1(new_n2437_), .A2(new_n2436_), .ZN(new_n2621_));
  NOR2_X1    g00186(.A1(new_n2612_), .A2(new_n2621_), .ZN(new_n2622_));
  NAND2_X1   g00187(.A1(new_n2620_), .A2(new_n2622_), .ZN(new_n2623_));
  AOI21_X1   g00188(.A1(new_n2623_), .A2(new_n2613_), .B(pi0056), .ZN(new_n2624_));
  INV_X1     g00189(.I(pi0074), .ZN(new_n2625_));
  NOR2_X1    g00190(.A1(new_n2604_), .A2(pi0038), .ZN(new_n2626_));
  INV_X1     g00191(.I(pi0039), .ZN(new_n2627_));
  INV_X1     g00192(.I(pi0299), .ZN(new_n2628_));
  INV_X1     g00193(.I(pi0222), .ZN(new_n2629_));
  INV_X1     g00194(.I(pi0332), .ZN(new_n2630_));
  INV_X1     g00195(.I(pi0224), .ZN(new_n2631_));
  AOI21_X1   g00196(.A1(pi0265), .A2(new_n2630_), .B(new_n2631_), .ZN(new_n2632_));
  INV_X1     g00197(.I(new_n2632_), .ZN(new_n2633_));
  NOR2_X1    g00198(.A1(new_n2443_), .A2(pi0224), .ZN(new_n2634_));
  INV_X1     g00199(.I(new_n2634_), .ZN(new_n2635_));
  NOR2_X1    g00200(.A1(new_n2635_), .A2(pi0929), .ZN(new_n2636_));
  AOI22_X1   g00201(.A1(new_n2636_), .A2(new_n2630_), .B1(new_n2629_), .B2(new_n2633_), .ZN(new_n2637_));
  NOR2_X1    g00202(.A1(new_n2634_), .A2(new_n2629_), .ZN(new_n2638_));
  NOR2_X1    g00203(.A1(new_n2638_), .A2(pi0223), .ZN(new_n2639_));
  OAI22_X1   g00204(.A1(new_n2637_), .A2(pi0223), .B1(new_n2438_), .B2(new_n2639_), .ZN(new_n2640_));
  NOR2_X1    g00205(.A1(pi0222), .A2(pi0224), .ZN(new_n2641_));
  INV_X1     g00206(.I(new_n2641_), .ZN(new_n2642_));
  NOR2_X1    g00207(.A1(new_n2642_), .A2(pi0223), .ZN(new_n2643_));
  INV_X1     g00208(.I(new_n2643_), .ZN(new_n2644_));
  OAI21_X1   g00209(.A1(new_n2557_), .A2(new_n2644_), .B(new_n2640_), .ZN(new_n2645_));
  NAND2_X1   g00210(.A1(new_n2645_), .A2(new_n2628_), .ZN(new_n2646_));
  INV_X1     g00211(.I(new_n2646_), .ZN(new_n2647_));
  AOI21_X1   g00212(.A1(new_n2561_), .A2(new_n2468_), .B(new_n2628_), .ZN(new_n2648_));
  OAI21_X1   g00213(.A1(new_n2648_), .A2(new_n2647_), .B(new_n2627_), .ZN(new_n2649_));
  NOR2_X1    g00214(.A1(new_n2649_), .A2(new_n2606_), .ZN(new_n2650_));
  NAND2_X1   g00215(.A1(new_n2468_), .A2(pi0299), .ZN(new_n2651_));
  AOI21_X1   g00216(.A1(new_n2473_), .A2(new_n2643_), .B(pi0299), .ZN(new_n2652_));
  NAND2_X1   g00217(.A1(new_n2640_), .A2(new_n2652_), .ZN(new_n2653_));
  NAND2_X1   g00218(.A1(new_n2651_), .A2(new_n2653_), .ZN(new_n2654_));
  INV_X1     g00219(.I(new_n2654_), .ZN(new_n2655_));
  NOR2_X1    g00220(.A1(new_n2573_), .A2(pi0087), .ZN(new_n2656_));
  INV_X1     g00221(.I(new_n2656_), .ZN(new_n2657_));
  NOR2_X1    g00222(.A1(new_n2657_), .A2(pi0100), .ZN(new_n2658_));
  INV_X1     g00223(.I(new_n2658_), .ZN(new_n2659_));
  NOR2_X1    g00224(.A1(new_n2659_), .A2(new_n2606_), .ZN(new_n2660_));
  INV_X1     g00225(.I(new_n2660_), .ZN(new_n2661_));
  AOI22_X1   g00226(.A1(new_n2650_), .A2(new_n2626_), .B1(new_n2655_), .B2(new_n2661_), .ZN(new_n2662_));
  OR2_X2     g00227(.A1(new_n2662_), .A2(pi0054), .Z(new_n2663_));
  NAND2_X1   g00228(.A1(new_n2655_), .A2(pi0054), .ZN(new_n2664_));
  AOI21_X1   g00229(.A1(new_n2663_), .A2(new_n2664_), .B(new_n2625_), .ZN(new_n2665_));
  AOI21_X1   g00230(.A1(new_n2662_), .A2(pi0054), .B(pi0074), .ZN(new_n2666_));
  INV_X1     g00231(.I(new_n2640_), .ZN(new_n2667_));
  INV_X1     g00232(.I(pi0223), .ZN(new_n2668_));
  NOR3_X1    g00233(.A1(pi0144), .A2(pi0174), .A3(pi0189), .ZN(new_n2669_));
  INV_X1     g00234(.I(new_n2669_), .ZN(new_n2670_));
  INV_X1     g00235(.I(new_n2556_), .ZN(new_n2671_));
  INV_X1     g00236(.I(pi0198), .ZN(new_n2672_));
  AOI21_X1   g00237(.A1(new_n2672_), .A2(pi0142), .B(pi0137), .ZN(new_n2673_));
  OAI21_X1   g00238(.A1(new_n2671_), .A2(new_n2673_), .B(new_n2464_), .ZN(new_n2674_));
  NAND3_X1   g00239(.A1(new_n2674_), .A2(new_n2668_), .A3(new_n2670_), .ZN(new_n2675_));
  NAND2_X1   g00240(.A1(new_n2630_), .A2(pi0234), .ZN(new_n2676_));
  NOR3_X1    g00241(.A1(new_n2672_), .A2(pi0095), .A3(pi0137), .ZN(new_n2677_));
  NOR2_X1    g00242(.A1(new_n2555_), .A2(new_n2677_), .ZN(new_n2678_));
  NOR2_X1    g00243(.A1(new_n2670_), .A2(pi0223), .ZN(new_n2679_));
  INV_X1     g00244(.I(new_n2679_), .ZN(new_n2680_));
  NOR2_X1    g00245(.A1(pi0234), .A2(pi0332), .ZN(new_n2681_));
  OAI21_X1   g00246(.A1(pi0137), .A2(new_n2672_), .B(new_n2531_), .ZN(new_n2682_));
  AOI21_X1   g00247(.A1(new_n2682_), .A2(new_n2681_), .B(new_n2680_), .ZN(new_n2683_));
  OAI21_X1   g00248(.A1(new_n2678_), .A2(new_n2676_), .B(new_n2683_), .ZN(new_n2684_));
  AOI21_X1   g00249(.A1(new_n2675_), .A2(new_n2684_), .B(new_n2642_), .ZN(new_n2685_));
  OAI21_X1   g00250(.A1(new_n2685_), .A2(new_n2667_), .B(new_n2628_), .ZN(new_n2686_));
  AOI21_X1   g00251(.A1(pi0095), .A2(pi0234), .B(pi0137), .ZN(new_n2687_));
  NOR2_X1    g00252(.A1(pi0152), .A2(pi0161), .ZN(new_n2688_));
  INV_X1     g00253(.I(new_n2688_), .ZN(new_n2689_));
  NOR2_X1    g00254(.A1(new_n2689_), .A2(pi0166), .ZN(new_n2690_));
  NOR2_X1    g00255(.A1(new_n2690_), .A2(pi0146), .ZN(new_n2691_));
  OAI21_X1   g00256(.A1(new_n2691_), .A2(pi0210), .B(new_n2687_), .ZN(new_n2692_));
  NAND2_X1   g00257(.A1(new_n2556_), .A2(new_n2692_), .ZN(new_n2693_));
  AOI21_X1   g00258(.A1(new_n2693_), .A2(new_n2630_), .B(new_n2457_), .ZN(new_n2694_));
  NOR3_X1    g00259(.A1(new_n2694_), .A2(new_n2458_), .A3(new_n2592_), .ZN(new_n2695_));
  OAI21_X1   g00260(.A1(new_n2695_), .A2(new_n2472_), .B(new_n2453_), .ZN(new_n2696_));
  AOI21_X1   g00261(.A1(new_n2696_), .A2(new_n2441_), .B(pi0215), .ZN(new_n2697_));
  AOI21_X1   g00262(.A1(new_n2697_), .A2(new_n2586_), .B(new_n2439_), .ZN(new_n2698_));
  AOI21_X1   g00263(.A1(new_n2698_), .A2(pi0299), .B(new_n2659_), .ZN(new_n2699_));
  OAI21_X1   g00264(.A1(new_n2655_), .A2(new_n2658_), .B(pi0075), .ZN(new_n2700_));
  AOI21_X1   g00265(.A1(new_n2699_), .A2(new_n2686_), .B(new_n2700_), .ZN(new_n2701_));
  INV_X1     g00266(.I(pi0100), .ZN(new_n2702_));
  AOI21_X1   g00267(.A1(new_n2654_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n2703_));
  INV_X1     g00268(.I(pi0252), .ZN(new_n2704_));
  AOI21_X1   g00269(.A1(pi0210), .A2(new_n2704_), .B(new_n2691_), .ZN(new_n2705_));
  NOR2_X1    g00270(.A1(new_n2589_), .A2(new_n2705_), .ZN(new_n2706_));
  INV_X1     g00271(.I(new_n2691_), .ZN(new_n2707_));
  NOR2_X1    g00272(.A1(new_n2590_), .A2(new_n2707_), .ZN(new_n2708_));
  INV_X1     g00273(.I(pi0210), .ZN(new_n2709_));
  NOR2_X1    g00274(.A1(new_n2709_), .A2(pi0137), .ZN(new_n2710_));
  NOR4_X1    g00275(.A1(new_n2587_), .A2(pi0252), .A3(new_n2691_), .A4(new_n2710_), .ZN(new_n2711_));
  NOR4_X1    g00276(.A1(new_n2711_), .A2(new_n2455_), .A3(pi0332), .A4(new_n2708_), .ZN(new_n2712_));
  OAI21_X1   g00277(.A1(new_n2706_), .A2(new_n2712_), .B(new_n2458_), .ZN(new_n2713_));
  NAND2_X1   g00278(.A1(new_n2713_), .A2(new_n2614_), .ZN(new_n2714_));
  OAI21_X1   g00279(.A1(new_n2714_), .A2(new_n2695_), .B(new_n2453_), .ZN(new_n2715_));
  NAND2_X1   g00280(.A1(new_n2715_), .A2(new_n2441_), .ZN(new_n2716_));
  NAND3_X1   g00281(.A1(new_n2716_), .A2(new_n2436_), .A3(new_n2586_), .ZN(new_n2717_));
  NAND3_X1   g00282(.A1(new_n2717_), .A2(pi0299), .A3(new_n2440_), .ZN(new_n2718_));
  NAND3_X1   g00283(.A1(new_n2718_), .A2(new_n2572_), .A3(new_n2686_), .ZN(new_n2719_));
  AOI21_X1   g00284(.A1(new_n2719_), .A2(new_n2703_), .B(pi0087), .ZN(new_n2720_));
  NAND2_X1   g00285(.A1(new_n2655_), .A2(pi0039), .ZN(new_n2721_));
  NAND3_X1   g00286(.A1(new_n2649_), .A2(pi0038), .A3(new_n2721_), .ZN(new_n2722_));
  NAND2_X1   g00287(.A1(new_n2722_), .A2(new_n2702_), .ZN(new_n2723_));
  INV_X1     g00288(.I(pi0142), .ZN(new_n2724_));
  INV_X1     g00289(.I(pi0032), .ZN(new_n2725_));
  INV_X1     g00290(.I(new_n2524_), .ZN(new_n2726_));
  INV_X1     g00291(.I(new_n2507_), .ZN(new_n2727_));
  NOR2_X1    g00292(.A1(new_n2516_), .A2(new_n2513_), .ZN(new_n2728_));
  INV_X1     g00293(.I(new_n2728_), .ZN(new_n2729_));
  NOR2_X1    g00294(.A1(new_n2727_), .A2(new_n2729_), .ZN(new_n2730_));
  INV_X1     g00295(.I(new_n2730_), .ZN(new_n2731_));
  NOR2_X1    g00296(.A1(pi0058), .A2(pi0091), .ZN(new_n2732_));
  INV_X1     g00297(.I(new_n2732_), .ZN(new_n2733_));
  NOR3_X1    g00298(.A1(pi0047), .A2(pi0109), .A3(pi0110), .ZN(new_n2734_));
  INV_X1     g00299(.I(new_n2734_), .ZN(new_n2735_));
  NOR2_X1    g00300(.A1(new_n2735_), .A2(new_n2733_), .ZN(new_n2736_));
  INV_X1     g00301(.I(new_n2736_), .ZN(new_n2737_));
  NOR2_X1    g00302(.A1(new_n2731_), .A2(new_n2737_), .ZN(new_n2738_));
  INV_X1     g00303(.I(new_n2738_), .ZN(new_n2739_));
  NOR2_X1    g00304(.A1(pi0090), .A2(pi0093), .ZN(new_n2740_));
  INV_X1     g00305(.I(new_n2740_), .ZN(new_n2741_));
  INV_X1     g00306(.I(pi0096), .ZN(new_n2742_));
  INV_X1     g00307(.I(pi0035), .ZN(new_n2743_));
  INV_X1     g00308(.I(pi0051), .ZN(new_n2744_));
  NAND2_X1   g00309(.A1(new_n2743_), .A2(new_n2744_), .ZN(new_n2745_));
  NOR2_X1    g00310(.A1(new_n2745_), .A2(pi0070), .ZN(new_n2746_));
  NAND2_X1   g00311(.A1(new_n2746_), .A2(new_n2742_), .ZN(new_n2747_));
  NOR2_X1    g00312(.A1(new_n2747_), .A2(new_n2741_), .ZN(new_n2748_));
  INV_X1     g00313(.I(new_n2748_), .ZN(new_n2749_));
  NOR2_X1    g00314(.A1(new_n2739_), .A2(new_n2749_), .ZN(new_n2750_));
  INV_X1     g00315(.I(new_n2750_), .ZN(new_n2751_));
  NOR2_X1    g00316(.A1(new_n2751_), .A2(new_n2726_), .ZN(new_n2752_));
  AOI21_X1   g00317(.A1(new_n2752_), .A2(pi0225), .B(new_n2725_), .ZN(new_n2753_));
  INV_X1     g00318(.I(new_n2753_), .ZN(new_n2754_));
  NOR2_X1    g00319(.A1(new_n2729_), .A2(new_n2510_), .ZN(new_n2755_));
  INV_X1     g00320(.I(new_n2755_), .ZN(new_n2756_));
  NOR2_X1    g00321(.A1(new_n2756_), .A2(pi0047), .ZN(new_n2757_));
  INV_X1     g00322(.I(new_n2757_), .ZN(new_n2758_));
  NOR2_X1    g00323(.A1(new_n2758_), .A2(new_n2727_), .ZN(new_n2759_));
  INV_X1     g00324(.I(new_n2759_), .ZN(new_n2760_));
  INV_X1     g00325(.I(new_n2746_), .ZN(new_n2761_));
  INV_X1     g00326(.I(new_n2520_), .ZN(new_n2762_));
  NOR2_X1    g00327(.A1(new_n2762_), .A2(pi0093), .ZN(new_n2763_));
  INV_X1     g00328(.I(new_n2763_), .ZN(new_n2764_));
  NOR3_X1    g00329(.A1(new_n2764_), .A2(new_n2761_), .A3(pi0091), .ZN(new_n2765_));
  INV_X1     g00330(.I(new_n2765_), .ZN(new_n2766_));
  NOR2_X1    g00331(.A1(new_n2760_), .A2(new_n2766_), .ZN(new_n2767_));
  INV_X1     g00332(.I(new_n2767_), .ZN(new_n2768_));
  AOI21_X1   g00333(.A1(new_n2768_), .A2(pi0096), .B(new_n2726_), .ZN(new_n2769_));
  INV_X1     g00334(.I(pi0225), .ZN(new_n2770_));
  INV_X1     g00335(.I(pi0093), .ZN(new_n2771_));
  NAND3_X1   g00336(.A1(new_n2547_), .A2(new_n2771_), .A3(new_n2520_), .ZN(new_n2772_));
  NOR2_X1    g00337(.A1(new_n2772_), .A2(new_n2743_), .ZN(new_n2773_));
  AOI21_X1   g00338(.A1(new_n2773_), .A2(new_n2770_), .B(pi0070), .ZN(new_n2774_));
  INV_X1     g00339(.I(new_n2774_), .ZN(new_n2775_));
  NOR2_X1    g00340(.A1(new_n2775_), .A2(pi0051), .ZN(new_n2776_));
  INV_X1     g00341(.I(new_n2776_), .ZN(new_n2777_));
  INV_X1     g00342(.I(new_n2772_), .ZN(new_n2778_));
  NOR2_X1    g00343(.A1(new_n2778_), .A2(new_n2743_), .ZN(new_n2779_));
  NOR2_X1    g00344(.A1(new_n2777_), .A2(new_n2779_), .ZN(new_n2780_));
  INV_X1     g00345(.I(new_n2780_), .ZN(new_n2781_));
  NOR2_X1    g00346(.A1(pi0046), .A2(pi0109), .ZN(new_n2782_));
  NAND2_X1   g00347(.A1(new_n2782_), .A2(new_n2509_), .ZN(new_n2783_));
  INV_X1     g00348(.I(new_n2783_), .ZN(new_n2784_));
  NAND3_X1   g00349(.A1(new_n2784_), .A2(new_n2512_), .A3(new_n2517_), .ZN(new_n2785_));
  NOR2_X1    g00350(.A1(new_n2785_), .A2(pi0058), .ZN(new_n2786_));
  INV_X1     g00351(.I(new_n2786_), .ZN(new_n2787_));
  INV_X1     g00352(.I(pi0060), .ZN(new_n2788_));
  NOR2_X1    g00353(.A1(new_n2727_), .A2(new_n2788_), .ZN(new_n2789_));
  NOR2_X1    g00354(.A1(new_n2789_), .A2(pi0053), .ZN(new_n2790_));
  NOR2_X1    g00355(.A1(pi0086), .A2(pi0094), .ZN(new_n2791_));
  INV_X1     g00356(.I(new_n2791_), .ZN(new_n2792_));
  INV_X1     g00357(.I(pi0053), .ZN(new_n2793_));
  AOI21_X1   g00358(.A1(new_n2507_), .A2(new_n2788_), .B(new_n2793_), .ZN(new_n2794_));
  NOR2_X1    g00359(.A1(new_n2794_), .A2(new_n2792_), .ZN(new_n2795_));
  INV_X1     g00360(.I(new_n2795_), .ZN(new_n2796_));
  NOR2_X1    g00361(.A1(new_n2796_), .A2(new_n2790_), .ZN(new_n2797_));
  INV_X1     g00362(.I(new_n2797_), .ZN(new_n2798_));
  NOR2_X1    g00363(.A1(new_n2798_), .A2(new_n2787_), .ZN(new_n2799_));
  NAND2_X1   g00364(.A1(new_n2799_), .A2(new_n2740_), .ZN(new_n2800_));
  INV_X1     g00365(.I(new_n2800_), .ZN(new_n2801_));
  NOR2_X1    g00366(.A1(new_n2801_), .A2(pi0035), .ZN(new_n2802_));
  NOR2_X1    g00367(.A1(new_n2802_), .A2(new_n2781_), .ZN(new_n2803_));
  NOR2_X1    g00368(.A1(new_n2803_), .A2(pi0096), .ZN(new_n2804_));
  INV_X1     g00369(.I(new_n2804_), .ZN(new_n2805_));
  NAND2_X1   g00370(.A1(new_n2805_), .A2(new_n2769_), .ZN(new_n2806_));
  AOI21_X1   g00371(.A1(new_n2806_), .A2(new_n2725_), .B(pi0095), .ZN(new_n2807_));
  AOI21_X1   g00372(.A1(new_n2807_), .A2(new_n2754_), .B(new_n2463_), .ZN(new_n2808_));
  OR2_X2     g00373(.A1(new_n2808_), .A2(pi0137), .Z(new_n2809_));
  NOR2_X1    g00374(.A1(new_n2768_), .A2(new_n2742_), .ZN(new_n2810_));
  INV_X1     g00375(.I(new_n2810_), .ZN(new_n2811_));
  NOR2_X1    g00376(.A1(new_n2548_), .A2(new_n2537_), .ZN(new_n2812_));
  INV_X1     g00377(.I(new_n2812_), .ZN(new_n2813_));
  NOR2_X1    g00378(.A1(new_n2813_), .A2(pi0051), .ZN(new_n2814_));
  NAND2_X1   g00379(.A1(new_n2814_), .A2(new_n2524_), .ZN(new_n2815_));
  NOR2_X1    g00380(.A1(new_n2811_), .A2(new_n2815_), .ZN(new_n2816_));
  INV_X1     g00381(.I(new_n2816_), .ZN(new_n2817_));
  INV_X1     g00382(.I(pi0040), .ZN(new_n2818_));
  NOR2_X1    g00383(.A1(new_n2553_), .A2(new_n2818_), .ZN(new_n2819_));
  NOR2_X1    g00384(.A1(new_n2819_), .A2(pi0032), .ZN(new_n2820_));
  INV_X1     g00385(.I(pi0072), .ZN(new_n2821_));
  NOR2_X1    g00386(.A1(new_n2750_), .A2(new_n2821_), .ZN(new_n2822_));
  NOR2_X1    g00387(.A1(new_n2822_), .A2(pi0040), .ZN(new_n2823_));
  INV_X1     g00388(.I(new_n2476_), .ZN(new_n2824_));
  NAND4_X1   g00389(.A1(new_n2490_), .A2(new_n2538_), .A3(new_n2539_), .A4(new_n2485_), .ZN(new_n2825_));
  INV_X1     g00390(.I(new_n2491_), .ZN(new_n2826_));
  NOR4_X1    g00391(.A1(new_n2825_), .A2(new_n2475_), .A3(new_n2824_), .A4(new_n2826_), .ZN(new_n2827_));
  INV_X1     g00392(.I(new_n2506_), .ZN(new_n2828_));
  NAND4_X1   g00393(.A1(new_n2827_), .A2(new_n2498_), .A3(new_n2828_), .A4(new_n2519_), .ZN(new_n2829_));
  INV_X1     g00394(.I(new_n2523_), .ZN(new_n2830_));
  NOR2_X1    g00395(.A1(new_n2829_), .A2(new_n2830_), .ZN(new_n2831_));
  NOR2_X1    g00396(.A1(new_n2831_), .A2(new_n2744_), .ZN(new_n2832_));
  NOR2_X1    g00397(.A1(new_n2832_), .A2(pi0096), .ZN(new_n2833_));
  INV_X1     g00398(.I(new_n2833_), .ZN(new_n2834_));
  INV_X1     g00399(.I(pi0070), .ZN(new_n2835_));
  AOI21_X1   g00400(.A1(new_n2778_), .A2(pi0225), .B(new_n2743_), .ZN(new_n2836_));
  INV_X1     g00401(.I(new_n2836_), .ZN(new_n2837_));
  INV_X1     g00402(.I(pi0091), .ZN(new_n2838_));
  NOR2_X1    g00403(.A1(new_n2760_), .A2(new_n2838_), .ZN(new_n2839_));
  NOR2_X1    g00404(.A1(new_n2839_), .A2(new_n2762_), .ZN(new_n2840_));
  INV_X1     g00405(.I(new_n2840_), .ZN(new_n2841_));
  NOR2_X1    g00406(.A1(new_n2731_), .A2(pi0109), .ZN(new_n2842_));
  NOR2_X1    g00407(.A1(new_n2842_), .A2(new_n2509_), .ZN(new_n2843_));
  INV_X1     g00408(.I(pi0047), .ZN(new_n2844_));
  AOI21_X1   g00409(.A1(new_n2507_), .A2(new_n2755_), .B(new_n2844_), .ZN(new_n2845_));
  NOR3_X1    g00410(.A1(new_n2843_), .A2(pi0091), .A3(new_n2845_), .ZN(new_n2846_));
  NOR2_X1    g00411(.A1(pi0047), .A2(pi0110), .ZN(new_n2847_));
  NOR2_X1    g00412(.A1(new_n2730_), .A2(new_n2508_), .ZN(new_n2848_));
  INV_X1     g00413(.I(pi0108), .ZN(new_n2849_));
  INV_X1     g00414(.I(new_n2503_), .ZN(new_n2850_));
  NOR2_X1    g00415(.A1(pi0081), .A2(pi0102), .ZN(new_n2851_));
  INV_X1     g00416(.I(new_n2851_), .ZN(new_n2852_));
  NOR4_X1    g00417(.A1(new_n2545_), .A2(new_n2499_), .A3(new_n2850_), .A4(new_n2852_), .ZN(new_n2853_));
  INV_X1     g00418(.I(new_n2853_), .ZN(new_n2854_));
  NOR3_X1    g00419(.A1(pi0050), .A2(pi0053), .A3(pi0060), .ZN(new_n2855_));
  NAND2_X1   g00420(.A1(new_n2855_), .A2(new_n2502_), .ZN(new_n2856_));
  NOR2_X1    g00421(.A1(new_n2856_), .A2(new_n2792_), .ZN(new_n2857_));
  INV_X1     g00422(.I(new_n2857_), .ZN(new_n2858_));
  NOR2_X1    g00423(.A1(new_n2854_), .A2(new_n2858_), .ZN(new_n2859_));
  INV_X1     g00424(.I(new_n2859_), .ZN(new_n2860_));
  NOR2_X1    g00425(.A1(new_n2860_), .A2(pi0097), .ZN(new_n2861_));
  NOR2_X1    g00426(.A1(new_n2861_), .A2(new_n2849_), .ZN(new_n2862_));
  NOR2_X1    g00427(.A1(new_n2862_), .A2(pi0046), .ZN(new_n2863_));
  INV_X1     g00428(.I(pi0097), .ZN(new_n2864_));
  NOR2_X1    g00429(.A1(new_n2859_), .A2(new_n2864_), .ZN(new_n2865_));
  INV_X1     g00430(.I(new_n2855_), .ZN(new_n2866_));
  NOR2_X1    g00431(.A1(new_n2545_), .A2(new_n2499_), .ZN(new_n2867_));
  INV_X1     g00432(.I(new_n2867_), .ZN(new_n2868_));
  NOR2_X1    g00433(.A1(new_n2868_), .A2(new_n2852_), .ZN(new_n2869_));
  INV_X1     g00434(.I(new_n2869_), .ZN(new_n2870_));
  NOR2_X1    g00435(.A1(new_n2870_), .A2(new_n2504_), .ZN(new_n2871_));
  INV_X1     g00436(.I(new_n2871_), .ZN(new_n2872_));
  NOR2_X1    g00437(.A1(new_n2872_), .A2(new_n2866_), .ZN(new_n2873_));
  INV_X1     g00438(.I(new_n2873_), .ZN(new_n2874_));
  NOR3_X1    g00439(.A1(new_n2874_), .A2(pi0086), .A3(new_n2514_), .ZN(new_n2875_));
  NOR2_X1    g00440(.A1(new_n2875_), .A2(pi0097), .ZN(new_n2876_));
  INV_X1     g00441(.I(new_n2876_), .ZN(new_n2877_));
  AOI21_X1   g00442(.A1(new_n2874_), .A2(pi0086), .B(pi0094), .ZN(new_n2878_));
  INV_X1     g00443(.I(pi0086), .ZN(new_n2879_));
  INV_X1     g00444(.I(new_n2790_), .ZN(new_n2880_));
  AOI21_X1   g00445(.A1(new_n2872_), .A2(pi0050), .B(pi0060), .ZN(new_n2881_));
  NOR2_X1    g00446(.A1(new_n2854_), .A2(new_n2502_), .ZN(new_n2882_));
  NOR2_X1    g00447(.A1(new_n2882_), .A2(pi0050), .ZN(new_n2883_));
  INV_X1     g00448(.I(pi0088), .ZN(new_n2884_));
  NOR4_X1    g00449(.A1(new_n2545_), .A2(pi0098), .A3(new_n2499_), .A4(new_n2852_), .ZN(new_n2885_));
  NOR2_X1    g00450(.A1(new_n2885_), .A2(new_n2884_), .ZN(new_n2886_));
  INV_X1     g00451(.I(pi0098), .ZN(new_n2887_));
  NOR2_X1    g00452(.A1(new_n2869_), .A2(new_n2887_), .ZN(new_n2888_));
  NOR3_X1    g00453(.A1(new_n2888_), .A2(pi0077), .A3(new_n2886_), .ZN(new_n2889_));
  INV_X1     g00454(.I(new_n2889_), .ZN(new_n2890_));
  NOR2_X1    g00455(.A1(new_n2545_), .A2(new_n2494_), .ZN(new_n2891_));
  AOI21_X1   g00456(.A1(new_n2891_), .A2(new_n2496_), .B(new_n2495_), .ZN(new_n2892_));
  INV_X1     g00457(.I(new_n2892_), .ZN(new_n2893_));
  INV_X1     g00458(.I(pi0107), .ZN(new_n2894_));
  INV_X1     g00459(.I(pi0063), .ZN(new_n2895_));
  INV_X1     g00460(.I(new_n2891_), .ZN(new_n2896_));
  NOR2_X1    g00461(.A1(new_n2896_), .A2(new_n2895_), .ZN(new_n2897_));
  AOI21_X1   g00462(.A1(new_n2897_), .A2(new_n2894_), .B(pi0064), .ZN(new_n2898_));
  AOI21_X1   g00463(.A1(new_n2545_), .A2(pi0071), .B(pi0065), .ZN(new_n2899_));
  INV_X1     g00464(.I(new_n2899_), .ZN(new_n2900_));
  INV_X1     g00465(.I(pi0103), .ZN(new_n2901_));
  NOR2_X1    g00466(.A1(new_n2825_), .A2(new_n2826_), .ZN(new_n2902_));
  INV_X1     g00467(.I(new_n2902_), .ZN(new_n2903_));
  NOR2_X1    g00468(.A1(new_n2903_), .A2(pi0067), .ZN(new_n2904_));
  INV_X1     g00469(.I(new_n2904_), .ZN(new_n2905_));
  NOR4_X1    g00470(.A1(new_n2905_), .A2(pi0069), .A3(pi0083), .A4(new_n2901_), .ZN(new_n2906_));
  NOR2_X1    g00471(.A1(pi0069), .A2(pi0083), .ZN(new_n2907_));
  INV_X1     g00472(.I(pi0069), .ZN(new_n2908_));
  AOI21_X1   g00473(.A1(new_n2492_), .A2(pi0083), .B(pi0103), .ZN(new_n2909_));
  OAI21_X1   g00474(.A1(new_n2904_), .A2(new_n2908_), .B(new_n2909_), .ZN(new_n2910_));
  INV_X1     g00475(.I(pi0082), .ZN(new_n2911_));
  INV_X1     g00476(.I(pi0111), .ZN(new_n2912_));
  NAND2_X1   g00477(.A1(new_n2911_), .A2(new_n2912_), .ZN(new_n2913_));
  INV_X1     g00478(.I(new_n2913_), .ZN(new_n2914_));
  INV_X1     g00479(.I(pi0084), .ZN(new_n2915_));
  NOR2_X1    g00480(.A1(new_n2540_), .A2(new_n2826_), .ZN(new_n2916_));
  NAND2_X1   g00481(.A1(new_n2916_), .A2(new_n2915_), .ZN(new_n2917_));
  NOR2_X1    g00482(.A1(new_n2917_), .A2(pi0068), .ZN(new_n2918_));
  NAND2_X1   g00483(.A1(new_n2918_), .A2(new_n2914_), .ZN(new_n2919_));
  NAND2_X1   g00484(.A1(new_n2919_), .A2(pi0036), .ZN(new_n2920_));
  NAND2_X1   g00485(.A1(new_n2903_), .A2(pi0067), .ZN(new_n2921_));
  INV_X1     g00486(.I(pi0068), .ZN(new_n2922_));
  INV_X1     g00487(.I(new_n2917_), .ZN(new_n2923_));
  NAND4_X1   g00488(.A1(new_n2923_), .A2(new_n2922_), .A3(pi0082), .A4(new_n2912_), .ZN(new_n2924_));
  NOR2_X1    g00489(.A1(pi0036), .A2(pi0067), .ZN(new_n2925_));
  NAND2_X1   g00490(.A1(new_n2922_), .A2(new_n2912_), .ZN(new_n2926_));
  INV_X1     g00491(.I(pi0073), .ZN(new_n2927_));
  NOR2_X1    g00492(.A1(new_n2927_), .A2(pi0066), .ZN(new_n2928_));
  INV_X1     g00493(.I(pi0066), .ZN(new_n2929_));
  NOR2_X1    g00494(.A1(new_n2929_), .A2(pi0073), .ZN(new_n2930_));
  OAI21_X1   g00495(.A1(new_n2928_), .A2(new_n2930_), .B(new_n2487_), .ZN(new_n2931_));
  INV_X1     g00496(.I(new_n2931_), .ZN(new_n2932_));
  INV_X1     g00497(.I(pi0045), .ZN(new_n2933_));
  NOR3_X1    g00498(.A1(new_n2484_), .A2(new_n2480_), .A3(pi0104), .ZN(new_n2934_));
  NAND2_X1   g00499(.A1(new_n2483_), .A2(new_n2482_), .ZN(new_n2935_));
  AOI21_X1   g00500(.A1(pi0085), .A2(pi0106), .B(pi0076), .ZN(new_n2936_));
  OAI21_X1   g00501(.A1(new_n2936_), .A2(new_n2483_), .B(new_n2481_), .ZN(new_n2937_));
  AOI21_X1   g00502(.A1(new_n2937_), .A2(new_n2935_), .B(pi0048), .ZN(new_n2938_));
  OAI21_X1   g00503(.A1(new_n2938_), .A2(new_n2539_), .B(new_n2478_), .ZN(new_n2939_));
  NAND3_X1   g00504(.A1(new_n2539_), .A2(new_n2477_), .A3(new_n2479_), .ZN(new_n2940_));
  AOI21_X1   g00505(.A1(new_n2539_), .A2(new_n2477_), .B(new_n2479_), .ZN(new_n2941_));
  AOI21_X1   g00506(.A1(new_n2939_), .A2(new_n2940_), .B(new_n2941_), .ZN(new_n2942_));
  AOI21_X1   g00507(.A1(new_n2942_), .A2(new_n2933_), .B(new_n2934_), .ZN(new_n2943_));
  AOI21_X1   g00508(.A1(new_n2539_), .A2(new_n2538_), .B(new_n2485_), .ZN(new_n2944_));
  NOR3_X1    g00509(.A1(new_n2943_), .A2(new_n2487_), .A3(new_n2944_), .ZN(new_n2945_));
  AOI21_X1   g00510(.A1(new_n2945_), .A2(new_n2491_), .B(new_n2932_), .ZN(new_n2946_));
  NOR2_X1    g00511(.A1(new_n2916_), .A2(new_n2915_), .ZN(new_n2947_));
  AOI21_X1   g00512(.A1(new_n2946_), .A2(new_n2915_), .B(new_n2947_), .ZN(new_n2948_));
  OAI21_X1   g00513(.A1(new_n2918_), .A2(new_n2912_), .B(new_n2911_), .ZN(new_n2949_));
  AOI21_X1   g00514(.A1(pi0068), .A2(new_n2917_), .B(new_n2949_), .ZN(new_n2950_));
  OAI21_X1   g00515(.A1(new_n2948_), .A2(new_n2926_), .B(new_n2950_), .ZN(new_n2951_));
  NAND3_X1   g00516(.A1(new_n2951_), .A2(new_n2924_), .A3(new_n2925_), .ZN(new_n2952_));
  NAND3_X1   g00517(.A1(new_n2952_), .A2(new_n2920_), .A3(new_n2921_), .ZN(new_n2953_));
  AOI21_X1   g00518(.A1(new_n2953_), .A2(new_n2907_), .B(new_n2910_), .ZN(new_n2954_));
  NOR3_X1    g00519(.A1(new_n2954_), .A2(pi0071), .A3(new_n2906_), .ZN(new_n2955_));
  NOR2_X1    g00520(.A1(new_n2955_), .A2(new_n2900_), .ZN(new_n2956_));
  AOI21_X1   g00521(.A1(new_n2896_), .A2(pi0107), .B(pi0063), .ZN(new_n2957_));
  OAI21_X1   g00522(.A1(new_n2956_), .A2(pi0107), .B(new_n2957_), .ZN(new_n2958_));
  NAND2_X1   g00523(.A1(new_n2958_), .A2(new_n2898_), .ZN(new_n2959_));
  NAND2_X1   g00524(.A1(new_n2959_), .A2(new_n2893_), .ZN(new_n2960_));
  INV_X1     g00525(.I(new_n2957_), .ZN(new_n2961_));
  INV_X1     g00526(.I(pi0071), .ZN(new_n2962_));
  AND3_X2    g00527(.A1(new_n2827_), .A2(pi0065), .A3(new_n2962_), .Z(new_n2963_));
  NOR3_X1    g00528(.A1(new_n2956_), .A2(pi0107), .A3(new_n2963_), .ZN(new_n2964_));
  OAI21_X1   g00529(.A1(new_n2964_), .A2(new_n2961_), .B(new_n2495_), .ZN(new_n2965_));
  NAND2_X1   g00530(.A1(new_n2965_), .A2(new_n2893_), .ZN(new_n2966_));
  NAND3_X1   g00531(.A1(new_n2966_), .A2(new_n2960_), .A3(new_n2851_), .ZN(new_n2967_));
  NOR2_X1    g00532(.A1(new_n2867_), .A2(new_n2500_), .ZN(new_n2968_));
  NOR4_X1    g00533(.A1(new_n2540_), .A2(new_n2824_), .A3(new_n2543_), .A4(new_n2826_), .ZN(new_n2969_));
  NAND4_X1   g00534(.A1(new_n2969_), .A2(new_n2500_), .A3(new_n2474_), .A4(new_n2498_), .ZN(new_n2970_));
  AOI21_X1   g00535(.A1(pi0102), .A2(new_n2970_), .B(new_n2968_), .ZN(new_n2971_));
  AOI21_X1   g00536(.A1(new_n2967_), .A2(new_n2971_), .B(new_n2850_), .ZN(new_n2972_));
  OAI21_X1   g00537(.A1(new_n2972_), .A2(new_n2890_), .B(new_n2883_), .ZN(new_n2973_));
  AOI21_X1   g00538(.A1(new_n2973_), .A2(new_n2881_), .B(new_n2880_), .ZN(new_n2974_));
  OAI21_X1   g00539(.A1(new_n2974_), .A2(new_n2794_), .B(new_n2879_), .ZN(new_n2975_));
  AOI21_X1   g00540(.A1(new_n2975_), .A2(new_n2878_), .B(new_n2877_), .ZN(new_n2976_));
  OAI21_X1   g00541(.A1(new_n2976_), .A2(new_n2865_), .B(new_n2849_), .ZN(new_n2977_));
  INV_X1     g00542(.I(new_n2512_), .ZN(new_n2978_));
  NOR3_X1    g00543(.A1(new_n2860_), .A2(new_n2511_), .A3(new_n2978_), .ZN(new_n2979_));
  NOR2_X1    g00544(.A1(new_n2979_), .A2(pi0109), .ZN(new_n2980_));
  INV_X1     g00545(.I(new_n2980_), .ZN(new_n2981_));
  AOI21_X1   g00546(.A1(new_n2977_), .A2(new_n2863_), .B(new_n2981_), .ZN(new_n2982_));
  OAI21_X1   g00547(.A1(new_n2982_), .A2(new_n2848_), .B(new_n2847_), .ZN(new_n2983_));
  AOI21_X1   g00548(.A1(new_n2983_), .A2(new_n2846_), .B(new_n2841_), .ZN(new_n2984_));
  INV_X1     g00549(.I(pi0090), .ZN(new_n2985_));
  NOR2_X1    g00550(.A1(new_n2738_), .A2(new_n2985_), .ZN(new_n2986_));
  AOI21_X1   g00551(.A1(pi0058), .A2(new_n2829_), .B(new_n2986_), .ZN(new_n2987_));
  NAND2_X1   g00552(.A1(new_n2987_), .A2(new_n2771_), .ZN(new_n2988_));
  NOR2_X1    g00553(.A1(new_n2548_), .A2(new_n2771_), .ZN(new_n2989_));
  NOR2_X1    g00554(.A1(new_n2989_), .A2(pi0035), .ZN(new_n2990_));
  OAI21_X1   g00555(.A1(new_n2984_), .A2(new_n2988_), .B(new_n2990_), .ZN(new_n2991_));
  NAND3_X1   g00556(.A1(new_n2991_), .A2(new_n2835_), .A3(new_n2837_), .ZN(new_n2992_));
  AOI21_X1   g00557(.A1(new_n2992_), .A2(new_n2744_), .B(new_n2834_), .ZN(new_n2993_));
  OAI21_X1   g00558(.A1(new_n2993_), .A2(pi0072), .B(new_n2823_), .ZN(new_n2994_));
  NAND3_X1   g00559(.A1(new_n2994_), .A2(new_n2817_), .A3(new_n2820_), .ZN(new_n2995_));
  NAND2_X1   g00560(.A1(new_n2995_), .A2(new_n2754_), .ZN(new_n2996_));
  NAND2_X1   g00561(.A1(new_n2996_), .A2(new_n2462_), .ZN(new_n2997_));
  INV_X1     g00562(.I(pi0479), .ZN(new_n2998_));
  NOR2_X1    g00563(.A1(new_n2553_), .A2(new_n2534_), .ZN(new_n2999_));
  NOR2_X1    g00564(.A1(new_n2999_), .A2(new_n2462_), .ZN(new_n3000_));
  INV_X1     g00565(.I(new_n3000_), .ZN(new_n3001_));
  NOR2_X1    g00566(.A1(new_n3001_), .A2(new_n2998_), .ZN(new_n3002_));
  INV_X1     g00567(.I(new_n3002_), .ZN(new_n3003_));
  NAND3_X1   g00568(.A1(new_n2997_), .A2(pi0137), .A3(new_n3003_), .ZN(new_n3004_));
  AOI21_X1   g00569(.A1(new_n3004_), .A2(new_n2809_), .B(new_n2672_), .ZN(new_n3005_));
  NOR2_X1    g00570(.A1(pi0070), .A2(pi0096), .ZN(new_n3006_));
  INV_X1     g00571(.I(new_n3006_), .ZN(new_n3007_));
  NOR4_X1    g00572(.A1(new_n3007_), .A2(pi0035), .A3(pi0040), .A4(new_n2770_), .ZN(new_n3008_));
  NAND2_X1   g00573(.A1(new_n2778_), .A2(pi0841), .ZN(new_n3009_));
  NAND2_X1   g00574(.A1(new_n2744_), .A2(new_n2821_), .ZN(new_n3010_));
  NOR2_X1    g00575(.A1(new_n3009_), .A2(new_n3010_), .ZN(new_n3011_));
  AOI21_X1   g00576(.A1(new_n3011_), .A2(new_n3008_), .B(new_n2725_), .ZN(new_n3012_));
  INV_X1     g00577(.I(new_n3012_), .ZN(new_n3013_));
  AOI21_X1   g00578(.A1(new_n2995_), .A2(new_n3013_), .B(pi0095), .ZN(new_n3014_));
  OAI21_X1   g00579(.A1(new_n3014_), .A2(new_n3002_), .B(pi0137), .ZN(new_n3015_));
  INV_X1     g00580(.I(pi0137), .ZN(new_n3016_));
  AOI21_X1   g00581(.A1(new_n2807_), .A2(new_n3013_), .B(new_n2463_), .ZN(new_n3017_));
  NAND2_X1   g00582(.A1(new_n3017_), .A2(new_n3016_), .ZN(new_n3018_));
  NAND2_X1   g00583(.A1(new_n3015_), .A2(new_n3018_), .ZN(new_n3019_));
  NOR2_X1    g00584(.A1(new_n3019_), .A2(pi0198), .ZN(new_n3020_));
  OAI21_X1   g00585(.A1(new_n3020_), .A2(new_n3005_), .B(new_n2724_), .ZN(new_n3021_));
  INV_X1     g00586(.I(pi1091), .ZN(new_n3022_));
  INV_X1     g00587(.I(pi0957), .ZN(new_n3023_));
  NOR2_X1    g00588(.A1(new_n3023_), .A2(pi0833), .ZN(new_n3024_));
  NOR2_X1    g00589(.A1(new_n3024_), .A2(new_n3022_), .ZN(new_n3025_));
  INV_X1     g00590(.I(new_n3025_), .ZN(new_n3026_));
  NAND3_X1   g00591(.A1(new_n3015_), .A2(new_n3018_), .A3(new_n3026_), .ZN(new_n3027_));
  INV_X1     g00592(.I(new_n2463_), .ZN(new_n3028_));
  NAND2_X1   g00593(.A1(new_n2798_), .A2(new_n2864_), .ZN(new_n3029_));
  NAND2_X1   g00594(.A1(new_n2517_), .A2(new_n2782_), .ZN(new_n3030_));
  NOR3_X1    g00595(.A1(new_n2865_), .A2(pi0108), .A3(pi0110), .ZN(new_n3031_));
  INV_X1     g00596(.I(new_n3031_), .ZN(new_n3032_));
  NOR3_X1    g00597(.A1(new_n3032_), .A2(new_n2764_), .A3(new_n3030_), .ZN(new_n3033_));
  AOI21_X1   g00598(.A1(new_n3033_), .A2(new_n3029_), .B(pi0035), .ZN(new_n3034_));
  OAI21_X1   g00599(.A1(new_n2781_), .A2(new_n3034_), .B(new_n2742_), .ZN(new_n3035_));
  AOI21_X1   g00600(.A1(new_n3035_), .A2(new_n2769_), .B(pi0032), .ZN(new_n3036_));
  NOR2_X1    g00601(.A1(new_n3012_), .A2(pi0095), .ZN(new_n3037_));
  INV_X1     g00602(.I(new_n3037_), .ZN(new_n3038_));
  OAI21_X1   g00603(.A1(new_n3036_), .A2(new_n3038_), .B(new_n3028_), .ZN(new_n3039_));
  INV_X1     g00604(.I(pi1092), .ZN(new_n3040_));
  INV_X1     g00605(.I(pi1093), .ZN(new_n3041_));
  NOR2_X1    g00606(.A1(new_n3040_), .A2(new_n3041_), .ZN(new_n3042_));
  INV_X1     g00607(.I(new_n3042_), .ZN(new_n3043_));
  INV_X1     g00608(.I(pi0829), .ZN(new_n3044_));
  INV_X1     g00609(.I(pi0950), .ZN(new_n3045_));
  NOR2_X1    g00610(.A1(new_n3044_), .A2(new_n3045_), .ZN(new_n3046_));
  INV_X1     g00611(.I(new_n3046_), .ZN(new_n3047_));
  NOR2_X1    g00612(.A1(new_n3043_), .A2(new_n3047_), .ZN(new_n3048_));
  NAND2_X1   g00613(.A1(new_n3039_), .A2(new_n3048_), .ZN(new_n3049_));
  INV_X1     g00614(.I(new_n3017_), .ZN(new_n3050_));
  INV_X1     g00615(.I(new_n3048_), .ZN(new_n3051_));
  AOI21_X1   g00616(.A1(new_n3050_), .A2(new_n3051_), .B(pi0137), .ZN(new_n3052_));
  AOI21_X1   g00617(.A1(new_n3052_), .A2(new_n3049_), .B(new_n3026_), .ZN(new_n3053_));
  NAND2_X1   g00618(.A1(new_n3015_), .A2(new_n3053_), .ZN(new_n3054_));
  AOI21_X1   g00619(.A1(new_n3027_), .A2(new_n3054_), .B(pi0198), .ZN(new_n3055_));
  OAI21_X1   g00620(.A1(new_n3055_), .A2(new_n3005_), .B(pi0142), .ZN(new_n3056_));
  NAND4_X1   g00621(.A1(new_n3056_), .A2(new_n3021_), .A3(pi0234), .A4(new_n2630_), .ZN(new_n3057_));
  INV_X1     g00622(.I(new_n2549_), .ZN(new_n3058_));
  NOR2_X1    g00623(.A1(new_n3058_), .A2(pi0040), .ZN(new_n3059_));
  AOI21_X1   g00624(.A1(new_n2803_), .A2(new_n3059_), .B(pi0032), .ZN(new_n3060_));
  NOR2_X1    g00625(.A1(new_n3060_), .A2(pi0095), .ZN(new_n3061_));
  AOI21_X1   g00626(.A1(new_n3061_), .A2(new_n2754_), .B(pi0137), .ZN(new_n3062_));
  NOR2_X1    g00627(.A1(new_n3000_), .A2(new_n2463_), .ZN(new_n3063_));
  AOI21_X1   g00628(.A1(new_n2994_), .A2(new_n2820_), .B(new_n2753_), .ZN(new_n3064_));
  OAI21_X1   g00629(.A1(new_n3064_), .A2(pi0095), .B(new_n3063_), .ZN(new_n3065_));
  AOI21_X1   g00630(.A1(new_n3065_), .A2(pi0137), .B(new_n3062_), .ZN(new_n3066_));
  NAND2_X1   g00631(.A1(new_n3066_), .A2(pi0198), .ZN(new_n3067_));
  INV_X1     g00632(.I(new_n3060_), .ZN(new_n3068_));
  NAND2_X1   g00633(.A1(new_n3068_), .A2(new_n3037_), .ZN(new_n3069_));
  NAND2_X1   g00634(.A1(new_n3069_), .A2(new_n3016_), .ZN(new_n3070_));
  INV_X1     g00635(.I(new_n3063_), .ZN(new_n3071_));
  NAND2_X1   g00636(.A1(new_n2994_), .A2(new_n2820_), .ZN(new_n3072_));
  AOI21_X1   g00637(.A1(new_n3072_), .A2(new_n3013_), .B(pi0095), .ZN(new_n3073_));
  OAI21_X1   g00638(.A1(new_n3073_), .A2(new_n3071_), .B(pi0137), .ZN(new_n3074_));
  NAND2_X1   g00639(.A1(new_n3074_), .A2(new_n3070_), .ZN(new_n3075_));
  OAI21_X1   g00640(.A1(pi0198), .A2(new_n3075_), .B(new_n3067_), .ZN(new_n3076_));
  NAND2_X1   g00641(.A1(new_n3076_), .A2(new_n2724_), .ZN(new_n3077_));
  INV_X1     g00642(.I(new_n2681_), .ZN(new_n3078_));
  INV_X1     g00643(.I(new_n3059_), .ZN(new_n3079_));
  NOR2_X1    g00644(.A1(new_n3022_), .A2(new_n3041_), .ZN(new_n3080_));
  INV_X1     g00645(.I(new_n3080_), .ZN(new_n3081_));
  NAND2_X1   g00646(.A1(pi0950), .A2(pi1092), .ZN(new_n3082_));
  NOR2_X1    g00647(.A1(new_n3082_), .A2(new_n3044_), .ZN(new_n3083_));
  INV_X1     g00648(.I(new_n3083_), .ZN(new_n3084_));
  NOR4_X1    g00649(.A1(new_n3034_), .A2(new_n3024_), .A3(new_n3081_), .A4(new_n3084_), .ZN(new_n3085_));
  NOR2_X1    g00650(.A1(new_n3051_), .A2(new_n3026_), .ZN(new_n3086_));
  NOR2_X1    g00651(.A1(new_n2802_), .A2(new_n3086_), .ZN(new_n3087_));
  NOR2_X1    g00652(.A1(new_n3087_), .A2(new_n3085_), .ZN(new_n3088_));
  NOR3_X1    g00653(.A1(new_n3088_), .A2(new_n2781_), .A3(new_n3079_), .ZN(new_n3089_));
  OAI21_X1   g00654(.A1(new_n3089_), .A2(pi0032), .B(new_n3037_), .ZN(new_n3090_));
  NAND2_X1   g00655(.A1(new_n3090_), .A2(new_n3016_), .ZN(new_n3091_));
  NAND2_X1   g00656(.A1(new_n3074_), .A2(new_n3091_), .ZN(new_n3092_));
  OAI21_X1   g00657(.A1(pi0198), .A2(new_n3092_), .B(new_n3067_), .ZN(new_n3093_));
  AOI21_X1   g00658(.A1(new_n3093_), .A2(pi0142), .B(new_n3078_), .ZN(new_n3094_));
  NAND2_X1   g00659(.A1(new_n3094_), .A2(new_n3077_), .ZN(new_n3095_));
  NAND4_X1   g00660(.A1(new_n3057_), .A2(new_n3095_), .A3(new_n2668_), .A4(new_n2670_), .ZN(new_n3096_));
  INV_X1     g00661(.I(pi0234), .ZN(new_n3097_));
  NOR3_X1    g00662(.A1(new_n3055_), .A2(new_n3097_), .A3(new_n3005_), .ZN(new_n3098_));
  NOR2_X1    g00663(.A1(new_n3093_), .A2(pi0234), .ZN(new_n3099_));
  OAI21_X1   g00664(.A1(new_n3098_), .A2(new_n3099_), .B(new_n2630_), .ZN(new_n3100_));
  NAND2_X1   g00665(.A1(new_n3100_), .A2(new_n2679_), .ZN(new_n3101_));
  NAND2_X1   g00666(.A1(new_n3096_), .A2(new_n3101_), .ZN(new_n3102_));
  AOI21_X1   g00667(.A1(new_n3102_), .A2(new_n2641_), .B(pi0299), .ZN(new_n3103_));
  AOI21_X1   g00668(.A1(new_n3103_), .A2(new_n2640_), .B(pi0039), .ZN(new_n3104_));
  NOR2_X1    g00669(.A1(new_n2621_), .A2(new_n2628_), .ZN(new_n3105_));
  INV_X1     g00670(.I(new_n2451_), .ZN(new_n3106_));
  INV_X1     g00671(.I(pi0146), .ZN(new_n3107_));
  AOI21_X1   g00672(.A1(new_n3004_), .A2(new_n2809_), .B(new_n2709_), .ZN(new_n3108_));
  NOR2_X1    g00673(.A1(new_n3019_), .A2(pi0210), .ZN(new_n3109_));
  OAI21_X1   g00674(.A1(new_n3109_), .A2(new_n3108_), .B(new_n3107_), .ZN(new_n3110_));
  AOI21_X1   g00675(.A1(new_n3027_), .A2(new_n3054_), .B(pi0210), .ZN(new_n3111_));
  OAI21_X1   g00676(.A1(new_n3111_), .A2(new_n3108_), .B(pi0146), .ZN(new_n3112_));
  NAND4_X1   g00677(.A1(new_n3112_), .A2(new_n3110_), .A3(pi0234), .A4(new_n2630_), .ZN(new_n3113_));
  NAND2_X1   g00678(.A1(new_n3066_), .A2(pi0210), .ZN(new_n3114_));
  OAI21_X1   g00679(.A1(pi0210), .A2(new_n3075_), .B(new_n3114_), .ZN(new_n3115_));
  NAND2_X1   g00680(.A1(new_n3115_), .A2(new_n3107_), .ZN(new_n3116_));
  OAI21_X1   g00681(.A1(pi0210), .A2(new_n3092_), .B(new_n3114_), .ZN(new_n3117_));
  AOI21_X1   g00682(.A1(new_n3117_), .A2(pi0146), .B(new_n3078_), .ZN(new_n3118_));
  AOI21_X1   g00683(.A1(new_n3118_), .A2(new_n3116_), .B(new_n2690_), .ZN(new_n3119_));
  NAND2_X1   g00684(.A1(new_n3113_), .A2(new_n3119_), .ZN(new_n3120_));
  NOR3_X1    g00685(.A1(new_n3111_), .A2(new_n3097_), .A3(new_n3108_), .ZN(new_n3121_));
  NOR2_X1    g00686(.A1(new_n3117_), .A2(pi0234), .ZN(new_n3122_));
  OAI21_X1   g00687(.A1(new_n3121_), .A2(new_n3122_), .B(new_n2630_), .ZN(new_n3123_));
  NAND2_X1   g00688(.A1(new_n3123_), .A2(new_n2690_), .ZN(new_n3124_));
  AOI21_X1   g00689(.A1(new_n3120_), .A2(new_n3124_), .B(new_n2457_), .ZN(new_n3125_));
  OAI21_X1   g00690(.A1(new_n3125_), .A2(new_n2592_), .B(pi0228), .ZN(new_n3126_));
  INV_X1     g00691(.I(new_n2820_), .ZN(new_n3127_));
  INV_X1     g00692(.I(new_n2823_), .ZN(new_n3128_));
  INV_X1     g00693(.I(new_n2990_), .ZN(new_n3129_));
  INV_X1     g00694(.I(new_n2847_), .ZN(new_n3130_));
  NAND2_X1   g00695(.A1(new_n2977_), .A2(new_n2863_), .ZN(new_n3131_));
  AOI21_X1   g00696(.A1(new_n3131_), .A2(new_n2508_), .B(new_n2848_), .ZN(new_n3132_));
  OAI21_X1   g00697(.A1(new_n3132_), .A2(new_n3130_), .B(new_n2846_), .ZN(new_n3133_));
  AOI21_X1   g00698(.A1(new_n3133_), .A2(new_n2840_), .B(new_n2988_), .ZN(new_n3134_));
  NOR2_X1    g00699(.A1(new_n3134_), .A2(new_n3129_), .ZN(new_n3135_));
  NOR3_X1    g00700(.A1(new_n3135_), .A2(pi0070), .A3(new_n2836_), .ZN(new_n3136_));
  OAI21_X1   g00701(.A1(new_n3136_), .A2(pi0051), .B(new_n2833_), .ZN(new_n3137_));
  AOI21_X1   g00702(.A1(new_n3137_), .A2(new_n2821_), .B(new_n3128_), .ZN(new_n3138_));
  OR2_X2     g00703(.A1(new_n3138_), .A2(new_n3127_), .Z(new_n3139_));
  AOI21_X1   g00704(.A1(new_n3139_), .A2(new_n2754_), .B(pi0095), .ZN(new_n3140_));
  OAI21_X1   g00705(.A1(new_n3140_), .A2(new_n3071_), .B(pi0137), .ZN(new_n3141_));
  NAND2_X1   g00706(.A1(new_n3141_), .A2(pi0210), .ZN(new_n3142_));
  NAND2_X1   g00707(.A1(new_n3091_), .A2(new_n2707_), .ZN(new_n3143_));
  NAND2_X1   g00708(.A1(new_n3070_), .A2(new_n2691_), .ZN(new_n3144_));
  NAND2_X1   g00709(.A1(new_n3143_), .A2(new_n3144_), .ZN(new_n3145_));
  NAND3_X1   g00710(.A1(new_n3145_), .A2(new_n2709_), .A3(new_n3097_), .ZN(new_n3146_));
  NAND2_X1   g00711(.A1(new_n3139_), .A2(new_n3013_), .ZN(new_n3147_));
  NAND2_X1   g00712(.A1(new_n3147_), .A2(new_n2462_), .ZN(new_n3148_));
  AOI21_X1   g00713(.A1(new_n3148_), .A2(new_n3063_), .B(new_n3016_), .ZN(new_n3149_));
  OAI22_X1   g00714(.A1(new_n3142_), .A2(new_n3062_), .B1(new_n3149_), .B2(new_n3146_), .ZN(new_n3150_));
  NAND3_X1   g00715(.A1(new_n2707_), .A2(new_n3025_), .A3(new_n3048_), .ZN(new_n3151_));
  NAND3_X1   g00716(.A1(new_n3050_), .A2(new_n3001_), .A3(new_n3151_), .ZN(new_n3152_));
  NOR2_X1    g00717(.A1(new_n3049_), .A2(new_n3000_), .ZN(new_n3153_));
  NAND3_X1   g00718(.A1(new_n3153_), .A2(new_n2707_), .A3(new_n3025_), .ZN(new_n3154_));
  NAND3_X1   g00719(.A1(new_n3152_), .A2(new_n3016_), .A3(new_n3154_), .ZN(new_n3155_));
  OR3_X2     g00720(.A1(new_n3138_), .A2(new_n2816_), .A3(new_n3127_), .Z(new_n3156_));
  AOI21_X1   g00721(.A1(new_n3156_), .A2(new_n3013_), .B(pi0095), .ZN(new_n3157_));
  OAI21_X1   g00722(.A1(new_n3157_), .A2(new_n3000_), .B(pi0137), .ZN(new_n3158_));
  NAND2_X1   g00723(.A1(new_n3158_), .A2(new_n3155_), .ZN(new_n3159_));
  AOI21_X1   g00724(.A1(new_n3159_), .A2(new_n2709_), .B(new_n3097_), .ZN(new_n3160_));
  NOR2_X1    g00725(.A1(new_n3150_), .A2(new_n3160_), .ZN(new_n3161_));
  NOR2_X1    g00726(.A1(new_n3000_), .A2(new_n3016_), .ZN(new_n3162_));
  INV_X1     g00727(.I(new_n3162_), .ZN(new_n3163_));
  NAND2_X1   g00728(.A1(new_n3156_), .A2(new_n2754_), .ZN(new_n3164_));
  AOI21_X1   g00729(.A1(new_n3164_), .A2(new_n2462_), .B(new_n3163_), .ZN(new_n3165_));
  NOR3_X1    g00730(.A1(new_n2808_), .A2(pi0137), .A3(new_n3000_), .ZN(new_n3166_));
  NOR4_X1    g00731(.A1(new_n3165_), .A2(new_n2709_), .A3(new_n3097_), .A4(new_n3166_), .ZN(new_n3167_));
  OAI21_X1   g00732(.A1(new_n3161_), .A2(new_n3167_), .B(new_n2456_), .ZN(new_n3168_));
  INV_X1     g00733(.I(new_n2690_), .ZN(new_n3169_));
  NOR2_X1    g00734(.A1(new_n2812_), .A2(new_n2835_), .ZN(new_n3170_));
  NOR2_X1    g00735(.A1(new_n3170_), .A2(new_n2528_), .ZN(new_n3171_));
  INV_X1     g00736(.I(new_n3171_), .ZN(new_n3172_));
  NOR2_X1    g00737(.A1(new_n3172_), .A2(new_n2726_), .ZN(new_n3173_));
  AOI21_X1   g00738(.A1(new_n3173_), .A2(new_n2775_), .B(pi0032), .ZN(new_n3174_));
  INV_X1     g00739(.I(new_n3174_), .ZN(new_n3175_));
  NOR3_X1    g00740(.A1(new_n2811_), .A2(pi0032), .A3(new_n2726_), .ZN(new_n3176_));
  NOR2_X1    g00741(.A1(new_n3175_), .A2(new_n3176_), .ZN(new_n3177_));
  INV_X1     g00742(.I(new_n2752_), .ZN(new_n3178_));
  INV_X1     g00743(.I(pi0841), .ZN(new_n3179_));
  NOR2_X1    g00744(.A1(new_n2770_), .A2(new_n3179_), .ZN(new_n3180_));
  OAI21_X1   g00745(.A1(new_n3178_), .A2(new_n3180_), .B(pi0032), .ZN(new_n3181_));
  INV_X1     g00746(.I(new_n3181_), .ZN(new_n3182_));
  NOR3_X1    g00747(.A1(new_n3182_), .A2(pi0095), .A3(new_n3177_), .ZN(new_n3183_));
  NAND2_X1   g00748(.A1(new_n2999_), .A2(new_n2463_), .ZN(new_n3184_));
  INV_X1     g00749(.I(new_n3184_), .ZN(new_n3185_));
  NOR3_X1    g00750(.A1(new_n3183_), .A2(new_n3016_), .A3(new_n3185_), .ZN(new_n3186_));
  INV_X1     g00751(.I(new_n3186_), .ZN(new_n3187_));
  INV_X1     g00752(.I(new_n3086_), .ZN(new_n3188_));
  NOR2_X1    g00753(.A1(new_n3127_), .A2(new_n3188_), .ZN(new_n3189_));
  NOR2_X1    g00754(.A1(new_n2810_), .A2(pi0072), .ZN(new_n3190_));
  INV_X1     g00755(.I(new_n3190_), .ZN(new_n3191_));
  INV_X1     g00756(.I(new_n3170_), .ZN(new_n3192_));
  NAND3_X1   g00757(.A1(new_n2973_), .A2(new_n2793_), .A3(new_n2881_), .ZN(new_n3193_));
  NAND2_X1   g00758(.A1(new_n3193_), .A2(new_n2879_), .ZN(new_n3194_));
  AOI21_X1   g00759(.A1(new_n3194_), .A2(new_n2878_), .B(new_n2877_), .ZN(new_n3195_));
  OAI21_X1   g00760(.A1(new_n3195_), .A2(pi0097), .B(new_n2849_), .ZN(new_n3196_));
  NAND2_X1   g00761(.A1(new_n3196_), .A2(new_n2863_), .ZN(new_n3197_));
  AOI21_X1   g00762(.A1(new_n3197_), .A2(new_n2508_), .B(new_n2848_), .ZN(new_n3198_));
  OAI21_X1   g00763(.A1(new_n3198_), .A2(new_n3130_), .B(new_n2846_), .ZN(new_n3199_));
  AOI21_X1   g00764(.A1(new_n3199_), .A2(new_n2840_), .B(new_n2988_), .ZN(new_n3200_));
  OAI21_X1   g00765(.A1(new_n3200_), .A2(new_n2989_), .B(new_n2743_), .ZN(new_n3201_));
  NAND2_X1   g00766(.A1(new_n3201_), .A2(new_n2776_), .ZN(new_n3202_));
  AND3_X2    g00767(.A1(new_n3202_), .A2(new_n2833_), .A3(new_n3192_), .Z(new_n3203_));
  OAI21_X1   g00768(.A1(new_n3203_), .A2(new_n3191_), .B(new_n2823_), .ZN(new_n3204_));
  NAND2_X1   g00769(.A1(new_n3204_), .A2(new_n3189_), .ZN(new_n3205_));
  OAI21_X1   g00770(.A1(new_n3195_), .A2(new_n2865_), .B(new_n2849_), .ZN(new_n3206_));
  AOI21_X1   g00771(.A1(new_n3206_), .A2(new_n2863_), .B(pi0109), .ZN(new_n3207_));
  OAI21_X1   g00772(.A1(new_n3207_), .A2(new_n2848_), .B(new_n2847_), .ZN(new_n3208_));
  NAND2_X1   g00773(.A1(new_n3208_), .A2(new_n2846_), .ZN(new_n3209_));
  AOI21_X1   g00774(.A1(new_n3209_), .A2(new_n2840_), .B(new_n2988_), .ZN(new_n3210_));
  NOR2_X1    g00775(.A1(new_n3210_), .A2(new_n2989_), .ZN(new_n3211_));
  NOR2_X1    g00776(.A1(new_n3211_), .A2(pi0035), .ZN(new_n3212_));
  OAI21_X1   g00777(.A1(new_n3212_), .A2(new_n2777_), .B(new_n2833_), .ZN(new_n3213_));
  OAI21_X1   g00778(.A1(new_n3213_), .A2(new_n3170_), .B(new_n3190_), .ZN(new_n3214_));
  AOI21_X1   g00779(.A1(new_n3214_), .A2(new_n2823_), .B(new_n3127_), .ZN(new_n3215_));
  NAND2_X1   g00780(.A1(new_n3215_), .A2(new_n3188_), .ZN(new_n3216_));
  NAND3_X1   g00781(.A1(new_n3216_), .A2(new_n3205_), .A3(new_n3181_), .ZN(new_n3217_));
  AOI21_X1   g00782(.A1(new_n3217_), .A2(new_n2462_), .B(new_n3000_), .ZN(new_n3218_));
  OAI21_X1   g00783(.A1(new_n3218_), .A2(pi0137), .B(new_n3187_), .ZN(new_n3219_));
  NAND2_X1   g00784(.A1(new_n3219_), .A2(new_n2709_), .ZN(new_n3220_));
  AOI21_X1   g00785(.A1(new_n2752_), .A2(new_n2770_), .B(new_n2725_), .ZN(new_n3221_));
  OR2_X2     g00786(.A1(new_n3221_), .A2(pi0095), .Z(new_n3222_));
  OAI21_X1   g00787(.A1(new_n3222_), .A2(new_n3177_), .B(new_n3184_), .ZN(new_n3223_));
  NAND2_X1   g00788(.A1(new_n3223_), .A2(pi0137), .ZN(new_n3224_));
  NOR2_X1    g00789(.A1(new_n3000_), .A2(pi0137), .ZN(new_n3225_));
  OAI21_X1   g00790(.A1(new_n3215_), .A2(new_n3221_), .B(new_n2462_), .ZN(new_n3226_));
  AOI21_X1   g00791(.A1(new_n3226_), .A2(new_n3225_), .B(new_n2709_), .ZN(new_n3227_));
  AOI21_X1   g00792(.A1(new_n3227_), .A2(new_n3224_), .B(new_n3078_), .ZN(new_n3228_));
  AOI21_X1   g00793(.A1(new_n3220_), .A2(new_n3228_), .B(new_n3169_), .ZN(new_n3229_));
  NOR2_X1    g00794(.A1(new_n3182_), .A2(pi0095), .ZN(new_n3230_));
  AOI21_X1   g00795(.A1(new_n3230_), .A2(new_n3175_), .B(new_n3016_), .ZN(new_n3231_));
  OAI21_X1   g00796(.A1(new_n3203_), .A2(pi0072), .B(new_n2823_), .ZN(new_n3232_));
  NAND2_X1   g00797(.A1(new_n3232_), .A2(new_n3189_), .ZN(new_n3233_));
  OAI21_X1   g00798(.A1(new_n3213_), .A2(new_n3170_), .B(new_n2821_), .ZN(new_n3234_));
  AOI21_X1   g00799(.A1(new_n3234_), .A2(new_n2823_), .B(new_n3127_), .ZN(new_n3235_));
  NAND2_X1   g00800(.A1(new_n3235_), .A2(new_n3188_), .ZN(new_n3236_));
  NAND3_X1   g00801(.A1(new_n3236_), .A2(new_n3233_), .A3(new_n3181_), .ZN(new_n3237_));
  NAND2_X1   g00802(.A1(new_n3237_), .A2(new_n2462_), .ZN(new_n3238_));
  AOI21_X1   g00803(.A1(new_n3238_), .A2(new_n3063_), .B(pi0137), .ZN(new_n3239_));
  OAI21_X1   g00804(.A1(new_n3239_), .A2(new_n3231_), .B(new_n2709_), .ZN(new_n3240_));
  NOR2_X1    g00805(.A1(new_n3222_), .A2(new_n3016_), .ZN(new_n3241_));
  AOI21_X1   g00806(.A1(new_n3241_), .A2(new_n3175_), .B(new_n2709_), .ZN(new_n3242_));
  OAI21_X1   g00807(.A1(new_n3235_), .A2(new_n3221_), .B(new_n2462_), .ZN(new_n3243_));
  NAND3_X1   g00808(.A1(new_n3243_), .A2(new_n3016_), .A3(new_n3063_), .ZN(new_n3244_));
  AOI21_X1   g00809(.A1(new_n3244_), .A2(new_n3242_), .B(new_n2676_), .ZN(new_n3245_));
  NAND2_X1   g00810(.A1(new_n3240_), .A2(new_n3245_), .ZN(new_n3246_));
  AOI21_X1   g00811(.A1(new_n3229_), .A2(new_n3246_), .B(pi0153), .ZN(new_n3247_));
  NAND3_X1   g00812(.A1(new_n3219_), .A2(pi0146), .A3(new_n2709_), .ZN(new_n3248_));
  OAI21_X1   g00813(.A1(new_n3215_), .A2(new_n3182_), .B(new_n2462_), .ZN(new_n3249_));
  AOI21_X1   g00814(.A1(new_n3249_), .A2(new_n3001_), .B(pi0137), .ZN(new_n3250_));
  NOR2_X1    g00815(.A1(pi0146), .A2(pi0210), .ZN(new_n3251_));
  OAI21_X1   g00816(.A1(new_n3250_), .A2(new_n3186_), .B(new_n3251_), .ZN(new_n3252_));
  NAND3_X1   g00817(.A1(new_n3248_), .A2(new_n3228_), .A3(new_n3252_), .ZN(new_n3253_));
  OAI21_X1   g00818(.A1(new_n3235_), .A2(new_n3182_), .B(new_n2462_), .ZN(new_n3254_));
  AOI21_X1   g00819(.A1(new_n3254_), .A2(new_n3063_), .B(pi0137), .ZN(new_n3255_));
  OAI21_X1   g00820(.A1(new_n3255_), .A2(new_n3231_), .B(new_n3251_), .ZN(new_n3256_));
  AND2_X2    g00821(.A1(new_n3256_), .A2(new_n3245_), .Z(new_n3257_));
  OAI21_X1   g00822(.A1(new_n3240_), .A2(new_n3107_), .B(new_n3257_), .ZN(new_n3258_));
  NAND3_X1   g00823(.A1(new_n3253_), .A2(new_n3258_), .A3(new_n3169_), .ZN(new_n3259_));
  NAND2_X1   g00824(.A1(new_n3259_), .A2(new_n3247_), .ZN(new_n3260_));
  NAND3_X1   g00825(.A1(new_n3260_), .A2(new_n2458_), .A3(new_n3168_), .ZN(new_n3261_));
  AOI21_X1   g00826(.A1(new_n3126_), .A2(new_n3261_), .B(pi0216), .ZN(new_n3262_));
  OAI21_X1   g00827(.A1(new_n3262_), .A2(new_n2454_), .B(new_n3106_), .ZN(new_n3263_));
  OAI21_X1   g00828(.A1(new_n3263_), .A2(pi0215), .B(new_n3105_), .ZN(new_n3264_));
  INV_X1     g00829(.I(pi0038), .ZN(new_n3265_));
  AOI21_X1   g00830(.A1(new_n2598_), .A2(pi0299), .B(new_n2647_), .ZN(new_n3266_));
  OAI21_X1   g00831(.A1(new_n3266_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n3267_));
  AOI21_X1   g00832(.A1(new_n3264_), .A2(new_n3104_), .B(new_n3267_), .ZN(new_n3268_));
  OAI21_X1   g00833(.A1(new_n3268_), .A2(new_n2723_), .B(new_n2720_), .ZN(new_n3269_));
  NOR2_X1    g00834(.A1(pi0038), .A2(pi0100), .ZN(new_n3270_));
  INV_X1     g00835(.I(new_n3270_), .ZN(new_n3271_));
  NOR2_X1    g00836(.A1(new_n3271_), .A2(pi0039), .ZN(new_n3272_));
  INV_X1     g00837(.I(new_n3272_), .ZN(new_n3273_));
  NOR2_X1    g00838(.A1(new_n3266_), .A2(new_n3273_), .ZN(new_n3274_));
  AOI21_X1   g00839(.A1(new_n2655_), .A2(new_n3273_), .B(new_n3274_), .ZN(new_n3275_));
  AOI21_X1   g00840(.A1(new_n3275_), .A2(pi0087), .B(pi0075), .ZN(new_n3276_));
  AOI21_X1   g00841(.A1(new_n3269_), .A2(new_n3276_), .B(new_n2701_), .ZN(new_n3277_));
  NAND2_X1   g00842(.A1(new_n2655_), .A2(new_n2565_), .ZN(new_n3278_));
  OAI21_X1   g00843(.A1(new_n3275_), .A2(new_n2565_), .B(new_n3278_), .ZN(new_n3279_));
  AOI21_X1   g00844(.A1(new_n3279_), .A2(pi0092), .B(pi0054), .ZN(new_n3280_));
  OAI21_X1   g00845(.A1(new_n3277_), .A2(pi0092), .B(new_n3280_), .ZN(new_n3281_));
  AOI21_X1   g00846(.A1(new_n3281_), .A2(new_n2666_), .B(new_n2665_), .ZN(new_n3282_));
  OAI21_X1   g00847(.A1(new_n3282_), .A2(pi0055), .B(new_n2624_), .ZN(new_n3283_));
  INV_X1     g00848(.I(pi0056), .ZN(new_n3284_));
  NOR2_X1    g00849(.A1(new_n2468_), .A2(new_n3284_), .ZN(new_n3285_));
  NOR2_X1    g00850(.A1(new_n2600_), .A2(pi0056), .ZN(new_n3286_));
  OAI21_X1   g00851(.A1(new_n3286_), .A2(new_n3285_), .B(pi0062), .ZN(new_n3287_));
  NAND2_X1   g00852(.A1(new_n3287_), .A2(new_n2469_), .ZN(new_n3288_));
  AOI21_X1   g00853(.A1(new_n3283_), .A2(new_n2601_), .B(new_n3288_), .ZN(new_n3289_));
  OAI21_X1   g00854(.A1(new_n3289_), .A2(new_n2584_), .B(new_n2581_), .ZN(po0153));
  NOR2_X1    g00855(.A1(pi0057), .A2(pi0059), .ZN(new_n3291_));
  NOR2_X1    g00856(.A1(new_n2436_), .A2(pi1146), .ZN(new_n3292_));
  INV_X1     g00857(.I(pi0276), .ZN(new_n3293_));
  NOR2_X1    g00858(.A1(new_n2614_), .A2(new_n3293_), .ZN(new_n3294_));
  NAND2_X1   g00859(.A1(new_n2444_), .A2(pi0939), .ZN(new_n3295_));
  NAND2_X1   g00860(.A1(new_n2447_), .A2(pi1146), .ZN(new_n3296_));
  AOI21_X1   g00861(.A1(new_n3296_), .A2(new_n3295_), .B(new_n2441_), .ZN(new_n3297_));
  NOR2_X1    g00862(.A1(new_n3297_), .A2(pi0215), .ZN(new_n3298_));
  INV_X1     g00863(.I(new_n3298_), .ZN(new_n3299_));
  AOI21_X1   g00864(.A1(new_n2441_), .A2(new_n3294_), .B(new_n3299_), .ZN(new_n3300_));
  NOR2_X1    g00865(.A1(new_n3300_), .A2(new_n3292_), .ZN(new_n3301_));
  NOR2_X1    g00866(.A1(new_n2460_), .A2(new_n3028_), .ZN(new_n3302_));
  NOR2_X1    g00867(.A1(pi0216), .A2(pi0221), .ZN(new_n3303_));
  INV_X1     g00868(.I(new_n3303_), .ZN(new_n3304_));
  NOR2_X1    g00869(.A1(new_n3304_), .A2(pi0215), .ZN(new_n3305_));
  NAND2_X1   g00870(.A1(new_n3302_), .A2(new_n3305_), .ZN(new_n3306_));
  INV_X1     g00871(.I(new_n3306_), .ZN(new_n3307_));
  NOR2_X1    g00872(.A1(new_n3301_), .A2(new_n3307_), .ZN(new_n3308_));
  INV_X1     g00873(.I(new_n3308_), .ZN(new_n3309_));
  AOI21_X1   g00874(.A1(new_n2460_), .A2(new_n2614_), .B(new_n3294_), .ZN(new_n3310_));
  OAI21_X1   g00875(.A1(pi0221), .A2(new_n3310_), .B(new_n3298_), .ZN(new_n3311_));
  OAI21_X1   g00876(.A1(new_n2436_), .A2(pi1146), .B(new_n3311_), .ZN(new_n3312_));
  NOR2_X1    g00877(.A1(new_n3312_), .A2(pi0154), .ZN(new_n3313_));
  INV_X1     g00878(.I(new_n3312_), .ZN(new_n3314_));
  NOR2_X1    g00879(.A1(new_n3314_), .A2(pi0154), .ZN(new_n3315_));
  INV_X1     g00880(.I(new_n3315_), .ZN(new_n3316_));
  OAI22_X1   g00881(.A1(new_n3316_), .A2(new_n2436_), .B1(new_n3309_), .B2(new_n3313_), .ZN(new_n3317_));
  NOR2_X1    g00882(.A1(new_n2571_), .A2(pi0056), .ZN(new_n3318_));
  INV_X1     g00883(.I(new_n3318_), .ZN(new_n3319_));
  NOR2_X1    g00884(.A1(new_n3319_), .A2(new_n2575_), .ZN(new_n3320_));
  INV_X1     g00885(.I(pi0154), .ZN(new_n3321_));
  NOR2_X1    g00886(.A1(new_n2530_), .A2(pi0228), .ZN(new_n3322_));
  AOI21_X1   g00887(.A1(pi0215), .A2(pi1146), .B(new_n3297_), .ZN(new_n3323_));
  AND3_X2    g00888(.A1(new_n3322_), .A2(new_n2614_), .A3(new_n3323_), .Z(new_n3324_));
  OAI21_X1   g00889(.A1(new_n3321_), .A2(new_n3308_), .B(new_n3324_), .ZN(new_n3325_));
  INV_X1     g00890(.I(new_n3325_), .ZN(new_n3326_));
  NOR2_X1    g00891(.A1(new_n3326_), .A2(new_n3317_), .ZN(new_n3327_));
  NAND3_X1   g00892(.A1(new_n3327_), .A2(new_n2602_), .A3(new_n2611_), .ZN(new_n3328_));
  OAI22_X1   g00893(.A1(new_n3328_), .A2(pi0056), .B1(new_n3317_), .B2(new_n3320_), .ZN(new_n3329_));
  NAND2_X1   g00894(.A1(new_n3329_), .A2(pi0062), .ZN(new_n3330_));
  NAND2_X1   g00895(.A1(new_n3330_), .A2(new_n3291_), .ZN(new_n3331_));
  INV_X1     g00896(.I(new_n3317_), .ZN(new_n3332_));
  NAND2_X1   g00897(.A1(new_n3326_), .A2(new_n2611_), .ZN(new_n3333_));
  NAND3_X1   g00898(.A1(new_n3333_), .A2(new_n3332_), .A3(pi0055), .ZN(new_n3334_));
  NOR2_X1    g00899(.A1(pi0223), .A2(pi0299), .ZN(new_n3335_));
  INV_X1     g00900(.I(new_n3335_), .ZN(new_n3336_));
  NOR2_X1    g00901(.A1(new_n2642_), .A2(new_n3336_), .ZN(new_n3337_));
  INV_X1     g00902(.I(new_n3337_), .ZN(new_n3338_));
  NOR2_X1    g00903(.A1(new_n3338_), .A2(new_n3028_), .ZN(new_n3339_));
  INV_X1     g00904(.I(new_n3339_), .ZN(new_n3340_));
  INV_X1     g00905(.I(pi0939), .ZN(new_n3341_));
  NOR2_X1    g00906(.A1(new_n2635_), .A2(new_n3341_), .ZN(new_n3342_));
  INV_X1     g00907(.I(pi1146), .ZN(new_n3343_));
  NOR2_X1    g00908(.A1(new_n2634_), .A2(new_n3343_), .ZN(new_n3344_));
  OAI21_X1   g00909(.A1(new_n3342_), .A2(new_n3344_), .B(pi0222), .ZN(new_n3345_));
  NOR2_X1    g00910(.A1(new_n2631_), .A2(pi0222), .ZN(new_n3346_));
  INV_X1     g00911(.I(new_n3346_), .ZN(new_n3347_));
  OAI21_X1   g00912(.A1(new_n3293_), .A2(new_n3347_), .B(new_n3345_), .ZN(new_n3348_));
  NOR2_X1    g00913(.A1(new_n3348_), .A2(pi0223), .ZN(new_n3349_));
  NOR2_X1    g00914(.A1(new_n2668_), .A2(pi1146), .ZN(new_n3350_));
  NOR3_X1    g00915(.A1(new_n3349_), .A2(pi0299), .A3(new_n3350_), .ZN(new_n3351_));
  INV_X1     g00916(.I(new_n3351_), .ZN(new_n3352_));
  NAND2_X1   g00917(.A1(new_n3332_), .A2(pi0299), .ZN(new_n3353_));
  NAND3_X1   g00918(.A1(new_n3353_), .A2(new_n3340_), .A3(new_n3352_), .ZN(new_n3354_));
  INV_X1     g00919(.I(new_n3354_), .ZN(new_n3355_));
  AOI21_X1   g00920(.A1(new_n3355_), .A2(new_n2563_), .B(pi0055), .ZN(new_n3356_));
  NOR2_X1    g00921(.A1(new_n3327_), .A2(new_n2628_), .ZN(new_n3357_));
  INV_X1     g00922(.I(new_n3357_), .ZN(new_n3358_));
  OAI21_X1   g00923(.A1(new_n3358_), .A2(new_n3273_), .B(pi0087), .ZN(new_n3359_));
  INV_X1     g00924(.I(pi0161), .ZN(new_n3360_));
  INV_X1     g00925(.I(pi0166), .ZN(new_n3361_));
  NOR2_X1    g00926(.A1(new_n2530_), .A2(pi0252), .ZN(new_n3362_));
  INV_X1     g00927(.I(new_n3362_), .ZN(new_n3363_));
  NAND3_X1   g00928(.A1(new_n3363_), .A2(new_n3360_), .A3(new_n3361_), .ZN(new_n3364_));
  AOI21_X1   g00929(.A1(pi0146), .A2(pi0252), .B(new_n2530_), .ZN(new_n3365_));
  INV_X1     g00930(.I(new_n3365_), .ZN(new_n3366_));
  OAI21_X1   g00931(.A1(pi0161), .A2(pi0166), .B(new_n3366_), .ZN(new_n3367_));
  AOI21_X1   g00932(.A1(new_n3367_), .A2(new_n3364_), .B(pi0152), .ZN(new_n3368_));
  INV_X1     g00933(.I(pi0152), .ZN(new_n3369_));
  NOR2_X1    g00934(.A1(new_n3365_), .A2(new_n3369_), .ZN(new_n3370_));
  NOR2_X1    g00935(.A1(new_n3368_), .A2(new_n3370_), .ZN(new_n3371_));
  NAND3_X1   g00936(.A1(new_n3265_), .A2(new_n2614_), .A3(new_n2458_), .ZN(new_n3372_));
  NOR4_X1    g00937(.A1(new_n3372_), .A2(pi0039), .A3(pi0154), .A4(new_n2628_), .ZN(new_n3373_));
  NAND3_X1   g00938(.A1(new_n3371_), .A2(new_n3323_), .A3(new_n3373_), .ZN(new_n3374_));
  NAND2_X1   g00939(.A1(new_n3374_), .A2(pi0100), .ZN(new_n3375_));
  OAI21_X1   g00940(.A1(new_n3265_), .A2(pi0100), .B(new_n3375_), .ZN(new_n3376_));
  NAND2_X1   g00941(.A1(new_n3358_), .A2(new_n3354_), .ZN(new_n3377_));
  AOI21_X1   g00942(.A1(new_n3377_), .A2(pi0039), .B(new_n3271_), .ZN(new_n3378_));
  INV_X1     g00943(.I(new_n3350_), .ZN(new_n3379_));
  NOR2_X1    g00944(.A1(new_n2811_), .A2(new_n2526_), .ZN(new_n3380_));
  NOR2_X1    g00945(.A1(new_n3380_), .A2(new_n2463_), .ZN(new_n3381_));
  NOR2_X1    g00946(.A1(new_n3381_), .A2(pi0224), .ZN(new_n3382_));
  NOR2_X1    g00947(.A1(new_n2631_), .A2(new_n3293_), .ZN(new_n3383_));
  OAI21_X1   g00948(.A1(new_n3382_), .A2(new_n3383_), .B(new_n2629_), .ZN(new_n3384_));
  NAND3_X1   g00949(.A1(new_n3384_), .A2(new_n2668_), .A3(new_n3345_), .ZN(new_n3385_));
  AOI21_X1   g00950(.A1(new_n3385_), .A2(new_n3379_), .B(pi0299), .ZN(new_n3386_));
  NOR2_X1    g00951(.A1(new_n3381_), .A2(new_n3000_), .ZN(new_n3387_));
  NOR2_X1    g00952(.A1(new_n3381_), .A2(new_n2460_), .ZN(new_n3388_));
  AOI21_X1   g00953(.A1(new_n3387_), .A2(new_n2458_), .B(new_n3388_), .ZN(new_n3389_));
  INV_X1     g00954(.I(new_n3389_), .ZN(new_n3390_));
  NAND2_X1   g00955(.A1(new_n3390_), .A2(pi0154), .ZN(new_n3391_));
  INV_X1     g00956(.I(new_n3381_), .ZN(new_n3392_));
  INV_X1     g00957(.I(new_n2822_), .ZN(new_n3393_));
  NOR2_X1    g00958(.A1(new_n3170_), .A2(new_n2779_), .ZN(new_n3394_));
  NAND2_X1   g00959(.A1(new_n3135_), .A2(new_n2835_), .ZN(new_n3395_));
  NAND2_X1   g00960(.A1(new_n3395_), .A2(new_n3394_), .ZN(new_n3396_));
  AOI21_X1   g00961(.A1(new_n3396_), .A2(new_n2744_), .B(new_n2834_), .ZN(new_n3397_));
  OAI21_X1   g00962(.A1(new_n3397_), .A2(pi0072), .B(new_n3393_), .ZN(new_n3398_));
  NAND2_X1   g00963(.A1(new_n3398_), .A2(new_n2533_), .ZN(new_n3399_));
  NOR2_X1    g00964(.A1(new_n2552_), .A2(new_n2818_), .ZN(new_n3400_));
  AOI21_X1   g00965(.A1(new_n3178_), .A2(pi0032), .B(new_n3400_), .ZN(new_n3401_));
  AOI21_X1   g00966(.A1(new_n3399_), .A2(new_n3401_), .B(pi0095), .ZN(new_n3402_));
  NOR2_X1    g00967(.A1(new_n3402_), .A2(new_n3071_), .ZN(new_n3403_));
  INV_X1     g00968(.I(new_n3403_), .ZN(new_n3404_));
  OAI22_X1   g00969(.A1(new_n3404_), .A2(pi0228), .B1(new_n2460_), .B2(new_n3392_), .ZN(new_n3405_));
  OAI21_X1   g00970(.A1(new_n3405_), .A2(pi0154), .B(new_n3391_), .ZN(new_n3406_));
  INV_X1     g00971(.I(new_n3301_), .ZN(new_n3407_));
  NAND2_X1   g00972(.A1(new_n3407_), .A2(pi0299), .ZN(new_n3408_));
  AOI21_X1   g00973(.A1(new_n3406_), .A2(new_n3305_), .B(new_n3408_), .ZN(new_n3409_));
  OAI21_X1   g00974(.A1(new_n3409_), .A2(new_n3386_), .B(new_n2627_), .ZN(new_n3410_));
  AOI22_X1   g00975(.A1(new_n3410_), .A2(new_n3378_), .B1(new_n3354_), .B2(new_n3376_), .ZN(new_n3411_));
  OAI22_X1   g00976(.A1(new_n3411_), .A2(pi0087), .B1(new_n3355_), .B2(new_n3359_), .ZN(new_n3412_));
  AOI21_X1   g00977(.A1(new_n3355_), .A2(pi0075), .B(pi0092), .ZN(new_n3413_));
  OAI21_X1   g00978(.A1(new_n3412_), .A2(pi0075), .B(new_n3413_), .ZN(new_n3414_));
  NOR2_X1    g00979(.A1(new_n2575_), .A2(new_n2565_), .ZN(new_n3415_));
  NAND2_X1   g00980(.A1(new_n3357_), .A2(new_n3415_), .ZN(new_n3416_));
  NAND3_X1   g00981(.A1(new_n3416_), .A2(new_n3354_), .A3(pi0092), .ZN(new_n3417_));
  NAND3_X1   g00982(.A1(new_n3414_), .A2(new_n2562_), .A3(new_n3417_), .ZN(new_n3418_));
  NAND2_X1   g00983(.A1(new_n3418_), .A2(new_n3356_), .ZN(new_n3419_));
  NAND3_X1   g00984(.A1(new_n3419_), .A2(new_n3284_), .A3(new_n3334_), .ZN(new_n3420_));
  AOI21_X1   g00985(.A1(new_n3332_), .A2(new_n2577_), .B(new_n3284_), .ZN(new_n3421_));
  AOI21_X1   g00986(.A1(new_n3328_), .A2(new_n3421_), .B(pi0062), .ZN(new_n3422_));
  AOI21_X1   g00987(.A1(new_n3420_), .A2(new_n3422_), .B(new_n3331_), .ZN(new_n3423_));
  OAI21_X1   g00988(.A1(new_n3332_), .A2(new_n3291_), .B(pi0239), .ZN(new_n3424_));
  INV_X1     g00989(.I(new_n3291_), .ZN(new_n3425_));
  OAI21_X1   g00990(.A1(new_n3321_), .A2(new_n3407_), .B(new_n3324_), .ZN(new_n3426_));
  AOI21_X1   g00991(.A1(pi0154), .A2(new_n3407_), .B(new_n3315_), .ZN(new_n3427_));
  NAND4_X1   g00992(.A1(new_n3426_), .A2(new_n3427_), .A3(new_n2602_), .A4(new_n2611_), .ZN(new_n3428_));
  NAND2_X1   g00993(.A1(new_n3427_), .A2(new_n2577_), .ZN(new_n3429_));
  AND3_X2    g00994(.A1(new_n3428_), .A2(pi0056), .A3(new_n3429_), .Z(new_n3430_));
  INV_X1     g00995(.I(new_n3427_), .ZN(new_n3431_));
  OAI21_X1   g00996(.A1(new_n3426_), .A2(new_n2612_), .B(pi0055), .ZN(new_n3432_));
  OAI21_X1   g00997(.A1(new_n3432_), .A2(new_n3431_), .B(new_n3284_), .ZN(new_n3433_));
  AOI21_X1   g00998(.A1(new_n3427_), .A2(pi0299), .B(new_n3351_), .ZN(new_n3434_));
  AOI21_X1   g00999(.A1(new_n3434_), .A2(new_n2563_), .B(pi0055), .ZN(new_n3435_));
  INV_X1     g01000(.I(new_n3415_), .ZN(new_n3436_));
  NAND2_X1   g01001(.A1(new_n3434_), .A2(new_n3436_), .ZN(new_n3437_));
  NOR3_X1    g01002(.A1(new_n3324_), .A2(new_n2628_), .A3(new_n3312_), .ZN(new_n3438_));
  OAI21_X1   g01003(.A1(new_n3438_), .A2(new_n3351_), .B(new_n3321_), .ZN(new_n3439_));
  OAI21_X1   g01004(.A1(new_n3407_), .A2(new_n2628_), .B(new_n3352_), .ZN(new_n3440_));
  NAND2_X1   g01005(.A1(new_n3440_), .A2(pi0154), .ZN(new_n3441_));
  NAND4_X1   g01006(.A1(new_n3439_), .A2(new_n2564_), .A3(new_n3272_), .A4(new_n3441_), .ZN(new_n3442_));
  NAND3_X1   g01007(.A1(new_n3442_), .A2(new_n3437_), .A3(pi0092), .ZN(new_n3443_));
  INV_X1     g01008(.I(pi0092), .ZN(new_n3444_));
  AOI21_X1   g01009(.A1(new_n3434_), .A2(pi0038), .B(pi0100), .ZN(new_n3445_));
  NOR2_X1    g01010(.A1(new_n3312_), .A2(new_n2628_), .ZN(new_n3446_));
  NOR2_X1    g01011(.A1(new_n2530_), .A2(new_n2627_), .ZN(new_n3447_));
  OAI21_X1   g01012(.A1(new_n3397_), .A2(new_n3191_), .B(new_n3393_), .ZN(new_n3448_));
  NAND2_X1   g01013(.A1(new_n3448_), .A2(new_n2533_), .ZN(new_n3449_));
  AOI21_X1   g01014(.A1(new_n3449_), .A2(new_n3401_), .B(pi0095), .ZN(new_n3450_));
  NOR2_X1    g01015(.A1(new_n3450_), .A2(new_n3000_), .ZN(new_n3451_));
  AOI21_X1   g01016(.A1(new_n3451_), .A2(new_n2627_), .B(new_n3447_), .ZN(new_n3452_));
  INV_X1     g01017(.I(new_n3452_), .ZN(new_n3453_));
  NAND4_X1   g01018(.A1(new_n3453_), .A2(new_n2614_), .A3(new_n2458_), .A4(new_n3323_), .ZN(new_n3454_));
  AOI21_X1   g01019(.A1(new_n3454_), .A2(new_n3446_), .B(new_n3351_), .ZN(new_n3455_));
  AOI21_X1   g01020(.A1(new_n3440_), .A2(pi0154), .B(pi0038), .ZN(new_n3456_));
  OAI21_X1   g01021(.A1(new_n3455_), .A2(pi0154), .B(new_n3456_), .ZN(new_n3457_));
  INV_X1     g01022(.I(pi0087), .ZN(new_n3458_));
  OAI21_X1   g01023(.A1(new_n3375_), .A2(new_n3434_), .B(new_n3458_), .ZN(new_n3459_));
  AOI21_X1   g01024(.A1(new_n3457_), .A2(new_n3445_), .B(new_n3459_), .ZN(new_n3460_));
  NAND3_X1   g01025(.A1(new_n3439_), .A2(new_n3272_), .A3(new_n3441_), .ZN(new_n3461_));
  NAND2_X1   g01026(.A1(new_n3434_), .A2(new_n3273_), .ZN(new_n3462_));
  AOI21_X1   g01027(.A1(new_n3461_), .A2(new_n3462_), .B(new_n3458_), .ZN(new_n3463_));
  NOR3_X1    g01028(.A1(new_n3460_), .A2(pi0075), .A3(new_n3463_), .ZN(new_n3464_));
  INV_X1     g01029(.I(pi0075), .ZN(new_n3465_));
  NOR2_X1    g01030(.A1(new_n3434_), .A2(new_n3465_), .ZN(new_n3466_));
  OAI21_X1   g01031(.A1(new_n3464_), .A2(new_n3466_), .B(new_n3444_), .ZN(new_n3467_));
  NAND3_X1   g01032(.A1(new_n3467_), .A2(new_n2562_), .A3(new_n3443_), .ZN(new_n3468_));
  AOI21_X1   g01033(.A1(new_n3468_), .A2(new_n3435_), .B(new_n3433_), .ZN(new_n3469_));
  NOR3_X1    g01034(.A1(new_n3469_), .A2(pi0062), .A3(new_n3430_), .ZN(new_n3470_));
  INV_X1     g01035(.I(pi0062), .ZN(new_n3471_));
  INV_X1     g01036(.I(new_n3320_), .ZN(new_n3472_));
  NAND2_X1   g01037(.A1(new_n3427_), .A2(new_n3472_), .ZN(new_n3473_));
  AOI21_X1   g01038(.A1(new_n3428_), .A2(new_n3473_), .B(new_n3471_), .ZN(new_n3474_));
  NOR3_X1    g01039(.A1(new_n3470_), .A2(new_n3425_), .A3(new_n3474_), .ZN(new_n3475_));
  INV_X1     g01040(.I(pi0239), .ZN(new_n3476_));
  OAI21_X1   g01041(.A1(new_n3427_), .A2(new_n3291_), .B(new_n3476_), .ZN(new_n3477_));
  OAI22_X1   g01042(.A1(new_n3423_), .A2(new_n3424_), .B1(new_n3475_), .B2(new_n3477_), .ZN(po0154));
  INV_X1     g01043(.I(pi0235), .ZN(new_n3479_));
  NOR2_X1    g01044(.A1(new_n2436_), .A2(pi1145), .ZN(new_n3480_));
  NAND2_X1   g01045(.A1(new_n2444_), .A2(pi0927), .ZN(new_n3481_));
  NAND2_X1   g01046(.A1(new_n2447_), .A2(pi1145), .ZN(new_n3482_));
  AOI21_X1   g01047(.A1(new_n3482_), .A2(new_n3481_), .B(new_n2441_), .ZN(new_n3483_));
  NOR2_X1    g01048(.A1(new_n3483_), .A2(pi0215), .ZN(new_n3484_));
  INV_X1     g01049(.I(new_n3484_), .ZN(new_n3485_));
  AOI21_X1   g01050(.A1(pi0216), .A2(pi0274), .B(pi0221), .ZN(new_n3486_));
  INV_X1     g01051(.I(new_n3322_), .ZN(new_n3487_));
  NOR2_X1    g01052(.A1(new_n3487_), .A2(pi0151), .ZN(new_n3488_));
  NOR2_X1    g01053(.A1(new_n2459_), .A2(pi0151), .ZN(new_n3489_));
  NOR2_X1    g01054(.A1(new_n3302_), .A2(new_n3489_), .ZN(new_n3490_));
  OAI21_X1   g01055(.A1(new_n3488_), .A2(new_n3490_), .B(new_n2614_), .ZN(new_n3491_));
  AOI21_X1   g01056(.A1(new_n3491_), .A2(new_n3486_), .B(new_n3485_), .ZN(new_n3492_));
  NOR2_X1    g01057(.A1(new_n3492_), .A2(new_n3480_), .ZN(new_n3493_));
  NAND2_X1   g01058(.A1(new_n3493_), .A2(new_n3320_), .ZN(new_n3494_));
  INV_X1     g01059(.I(new_n3480_), .ZN(new_n3495_));
  OAI21_X1   g01060(.A1(new_n3489_), .A2(pi0216), .B(new_n3486_), .ZN(new_n3496_));
  NAND2_X1   g01061(.A1(new_n3484_), .A2(new_n3496_), .ZN(new_n3497_));
  NAND2_X1   g01062(.A1(new_n3497_), .A2(new_n3495_), .ZN(new_n3498_));
  INV_X1     g01063(.I(new_n3498_), .ZN(new_n3499_));
  INV_X1     g01064(.I(new_n3302_), .ZN(new_n3500_));
  NOR2_X1    g01065(.A1(new_n3500_), .A2(new_n2559_), .ZN(new_n3501_));
  INV_X1     g01066(.I(new_n3501_), .ZN(new_n3502_));
  AOI21_X1   g01067(.A1(pi0216), .A2(pi0274), .B(new_n3502_), .ZN(new_n3503_));
  NOR2_X1    g01068(.A1(new_n3499_), .A2(new_n3503_), .ZN(new_n3504_));
  INV_X1     g01069(.I(new_n3504_), .ZN(new_n3505_));
  NAND2_X1   g01070(.A1(new_n3472_), .A2(new_n3505_), .ZN(new_n3506_));
  AOI21_X1   g01071(.A1(new_n3494_), .A2(new_n3506_), .B(new_n3471_), .ZN(new_n3507_));
  NOR3_X1    g01072(.A1(new_n3507_), .A2(new_n3479_), .A3(new_n3425_), .ZN(new_n3508_));
  NOR3_X1    g01073(.A1(new_n3492_), .A2(new_n2612_), .A3(new_n3480_), .ZN(new_n3509_));
  NOR2_X1    g01074(.A1(new_n3504_), .A2(new_n2611_), .ZN(new_n3510_));
  OAI21_X1   g01075(.A1(new_n3509_), .A2(new_n3510_), .B(pi0055), .ZN(new_n3511_));
  INV_X1     g01076(.I(pi1145), .ZN(new_n3512_));
  NAND2_X1   g01077(.A1(new_n3512_), .A2(pi0223), .ZN(new_n3513_));
  INV_X1     g01078(.I(pi0927), .ZN(new_n3514_));
  NOR2_X1    g01079(.A1(new_n2635_), .A2(new_n3514_), .ZN(new_n3515_));
  NOR2_X1    g01080(.A1(new_n2634_), .A2(new_n3512_), .ZN(new_n3516_));
  OAI21_X1   g01081(.A1(new_n3515_), .A2(new_n3516_), .B(pi0222), .ZN(new_n3517_));
  NOR2_X1    g01082(.A1(new_n2631_), .A2(pi0274), .ZN(new_n3518_));
  NAND2_X1   g01083(.A1(new_n3518_), .A2(new_n2629_), .ZN(new_n3519_));
  NAND3_X1   g01084(.A1(new_n3517_), .A2(new_n2668_), .A3(new_n3519_), .ZN(new_n3520_));
  NAND3_X1   g01085(.A1(new_n3520_), .A2(new_n2628_), .A3(new_n3513_), .ZN(new_n3521_));
  INV_X1     g01086(.I(new_n3521_), .ZN(new_n3522_));
  NOR2_X1    g01087(.A1(new_n3522_), .A2(new_n3339_), .ZN(new_n3523_));
  INV_X1     g01088(.I(new_n3523_), .ZN(new_n3524_));
  AOI21_X1   g01089(.A1(new_n3505_), .A2(pi0299), .B(new_n3524_), .ZN(new_n3525_));
  AOI21_X1   g01090(.A1(new_n3525_), .A2(new_n2563_), .B(pi0055), .ZN(new_n3526_));
  AOI21_X1   g01091(.A1(new_n3493_), .A2(pi0299), .B(new_n3524_), .ZN(new_n3527_));
  OAI21_X1   g01092(.A1(new_n3527_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n3528_));
  OAI21_X1   g01093(.A1(new_n3382_), .A2(new_n3518_), .B(new_n2629_), .ZN(new_n3529_));
  NAND3_X1   g01094(.A1(new_n3529_), .A2(new_n2668_), .A3(new_n3517_), .ZN(new_n3530_));
  AOI21_X1   g01095(.A1(new_n3530_), .A2(new_n3513_), .B(pi0299), .ZN(new_n3531_));
  INV_X1     g01096(.I(new_n3486_), .ZN(new_n3532_));
  INV_X1     g01097(.I(pi0151), .ZN(new_n3533_));
  NAND2_X1   g01098(.A1(new_n3405_), .A2(new_n3533_), .ZN(new_n3534_));
  NAND2_X1   g01099(.A1(new_n3389_), .A2(pi0151), .ZN(new_n3535_));
  AOI21_X1   g01100(.A1(new_n3534_), .A2(new_n3535_), .B(pi0216), .ZN(new_n3536_));
  OAI21_X1   g01101(.A1(new_n3536_), .A2(new_n3532_), .B(new_n3484_), .ZN(new_n3537_));
  AOI21_X1   g01102(.A1(new_n3537_), .A2(new_n3495_), .B(new_n2628_), .ZN(new_n3538_));
  NOR3_X1    g01103(.A1(new_n3538_), .A2(pi0039), .A3(new_n3531_), .ZN(new_n3539_));
  AOI21_X1   g01104(.A1(new_n3525_), .A2(pi0038), .B(pi0100), .ZN(new_n3540_));
  OAI21_X1   g01105(.A1(new_n3539_), .A2(new_n3528_), .B(new_n3540_), .ZN(new_n3541_));
  AOI21_X1   g01106(.A1(new_n3525_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n3542_));
  NOR2_X1    g01107(.A1(new_n2460_), .A2(new_n2463_), .ZN(new_n3543_));
  INV_X1     g01108(.I(new_n3371_), .ZN(new_n3544_));
  NOR2_X1    g01109(.A1(new_n3544_), .A2(pi0228), .ZN(new_n3545_));
  NOR2_X1    g01110(.A1(new_n3545_), .A2(new_n3543_), .ZN(new_n3546_));
  AOI21_X1   g01111(.A1(new_n3546_), .A2(new_n3533_), .B(new_n3491_), .ZN(new_n3547_));
  OAI21_X1   g01112(.A1(new_n3547_), .A2(new_n3532_), .B(new_n3484_), .ZN(new_n3548_));
  NAND3_X1   g01113(.A1(new_n3548_), .A2(pi0299), .A3(new_n3495_), .ZN(new_n3549_));
  NAND3_X1   g01114(.A1(new_n3549_), .A2(new_n2572_), .A3(new_n3523_), .ZN(new_n3550_));
  NAND2_X1   g01115(.A1(new_n3550_), .A2(new_n3542_), .ZN(new_n3551_));
  NAND3_X1   g01116(.A1(new_n3541_), .A2(new_n3458_), .A3(new_n3551_), .ZN(new_n3552_));
  INV_X1     g01117(.I(new_n3525_), .ZN(new_n3553_));
  NOR2_X1    g01118(.A1(new_n3527_), .A2(new_n3273_), .ZN(new_n3554_));
  AOI21_X1   g01119(.A1(new_n3273_), .A2(new_n3553_), .B(new_n3554_), .ZN(new_n3555_));
  NAND2_X1   g01120(.A1(new_n3555_), .A2(pi0087), .ZN(new_n3556_));
  AOI21_X1   g01121(.A1(new_n3552_), .A2(new_n3556_), .B(pi0075), .ZN(new_n3557_));
  OAI21_X1   g01122(.A1(new_n3553_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n3558_));
  NOR2_X1    g01123(.A1(new_n3555_), .A2(new_n2565_), .ZN(new_n3559_));
  AOI21_X1   g01124(.A1(new_n2565_), .A2(new_n3553_), .B(new_n3559_), .ZN(new_n3560_));
  OAI22_X1   g01125(.A1(new_n3557_), .A2(new_n3558_), .B1(new_n3444_), .B2(new_n3560_), .ZN(new_n3561_));
  OAI21_X1   g01126(.A1(new_n3561_), .A2(new_n2563_), .B(new_n3526_), .ZN(new_n3562_));
  NAND3_X1   g01127(.A1(new_n3562_), .A2(new_n3284_), .A3(new_n3511_), .ZN(new_n3563_));
  NAND2_X1   g01128(.A1(new_n3504_), .A2(new_n2577_), .ZN(new_n3564_));
  OAI21_X1   g01129(.A1(new_n3493_), .A2(new_n2577_), .B(new_n3564_), .ZN(new_n3565_));
  AOI21_X1   g01130(.A1(new_n3565_), .A2(pi0056), .B(pi0062), .ZN(new_n3566_));
  NAND2_X1   g01131(.A1(new_n3563_), .A2(new_n3566_), .ZN(new_n3567_));
  NAND2_X1   g01132(.A1(new_n3503_), .A2(pi0235), .ZN(new_n3568_));
  NAND2_X1   g01133(.A1(new_n3568_), .A2(new_n3425_), .ZN(new_n3569_));
  AOI21_X1   g01134(.A1(pi0215), .A2(pi1145), .B(new_n3483_), .ZN(new_n3570_));
  NAND3_X1   g01135(.A1(new_n3322_), .A2(new_n2614_), .A3(new_n3570_), .ZN(new_n3571_));
  NOR2_X1    g01136(.A1(new_n3571_), .A2(new_n2577_), .ZN(new_n3572_));
  NAND2_X1   g01137(.A1(new_n3572_), .A2(new_n3284_), .ZN(new_n3573_));
  NAND3_X1   g01138(.A1(new_n3573_), .A2(pi0062), .A3(new_n3499_), .ZN(new_n3574_));
  NAND3_X1   g01139(.A1(new_n3574_), .A2(new_n3479_), .A3(new_n3291_), .ZN(new_n3575_));
  OAI21_X1   g01140(.A1(new_n3572_), .A2(new_n3498_), .B(pi0056), .ZN(new_n3576_));
  NAND2_X1   g01141(.A1(new_n3576_), .A2(new_n3471_), .ZN(new_n3577_));
  NOR2_X1    g01142(.A1(new_n3498_), .A2(new_n2628_), .ZN(new_n3578_));
  NOR2_X1    g01143(.A1(new_n3578_), .A2(new_n3522_), .ZN(new_n3579_));
  AOI21_X1   g01144(.A1(new_n3579_), .A2(new_n2563_), .B(pi0055), .ZN(new_n3580_));
  NAND2_X1   g01145(.A1(new_n3571_), .A2(new_n3578_), .ZN(new_n3581_));
  NAND3_X1   g01146(.A1(new_n3581_), .A2(new_n2574_), .A3(new_n3521_), .ZN(new_n3582_));
  OAI21_X1   g01147(.A1(new_n3582_), .A2(new_n2565_), .B(pi0092), .ZN(new_n3583_));
  AOI21_X1   g01148(.A1(new_n3436_), .A2(new_n3579_), .B(new_n3583_), .ZN(new_n3584_));
  NOR2_X1    g01149(.A1(new_n3544_), .A2(new_n2702_), .ZN(new_n3585_));
  AOI22_X1   g01150(.A1(new_n3453_), .A2(new_n2702_), .B1(new_n2627_), .B2(new_n3585_), .ZN(new_n3586_));
  NAND4_X1   g01151(.A1(new_n3570_), .A2(new_n3265_), .A3(new_n2614_), .A4(new_n2458_), .ZN(new_n3587_));
  OAI21_X1   g01152(.A1(new_n3586_), .A2(new_n3587_), .B(new_n3578_), .ZN(new_n3588_));
  NOR2_X1    g01153(.A1(new_n3522_), .A2(pi0087), .ZN(new_n3589_));
  NAND2_X1   g01154(.A1(new_n3579_), .A2(new_n3273_), .ZN(new_n3590_));
  NAND2_X1   g01155(.A1(new_n3582_), .A2(new_n3590_), .ZN(new_n3591_));
  AOI22_X1   g01156(.A1(new_n3588_), .A2(new_n3589_), .B1(pi0087), .B2(new_n3591_), .ZN(new_n3592_));
  NOR2_X1    g01157(.A1(new_n3579_), .A2(new_n3465_), .ZN(new_n3593_));
  AOI21_X1   g01158(.A1(new_n3592_), .A2(new_n3465_), .B(new_n3593_), .ZN(new_n3594_));
  OAI21_X1   g01159(.A1(new_n3594_), .A2(pi0092), .B(new_n2562_), .ZN(new_n3595_));
  OAI21_X1   g01160(.A1(new_n3595_), .A2(new_n3584_), .B(new_n3580_), .ZN(new_n3596_));
  NOR2_X1    g01161(.A1(new_n3571_), .A2(new_n2612_), .ZN(new_n3597_));
  NOR2_X1    g01162(.A1(new_n3597_), .A2(new_n2602_), .ZN(new_n3598_));
  AOI21_X1   g01163(.A1(new_n3598_), .A2(new_n3499_), .B(pi0056), .ZN(new_n3599_));
  AOI21_X1   g01164(.A1(new_n3596_), .A2(new_n3599_), .B(new_n3577_), .ZN(new_n3600_));
  OAI22_X1   g01165(.A1(new_n3600_), .A2(new_n3575_), .B1(new_n3499_), .B2(new_n3569_), .ZN(new_n3601_));
  AOI21_X1   g01166(.A1(new_n3567_), .A2(new_n3508_), .B(new_n3601_), .ZN(po0155));
  INV_X1     g01167(.I(pi0944), .ZN(new_n3603_));
  NOR2_X1    g01168(.A1(new_n2447_), .A2(new_n3603_), .ZN(new_n3604_));
  INV_X1     g01169(.I(pi1143), .ZN(new_n3605_));
  NOR2_X1    g01170(.A1(new_n2444_), .A2(new_n3605_), .ZN(new_n3606_));
  OAI21_X1   g01171(.A1(new_n3604_), .A2(new_n3606_), .B(pi0221), .ZN(new_n3607_));
  AOI21_X1   g01172(.A1(pi0216), .A2(pi0264), .B(pi0221), .ZN(new_n3608_));
  NAND2_X1   g01173(.A1(new_n2457_), .A2(new_n3107_), .ZN(new_n3609_));
  INV_X1     g01174(.I(pi0284), .ZN(new_n3610_));
  NOR2_X1    g01175(.A1(new_n2463_), .A2(new_n3610_), .ZN(new_n3611_));
  NAND2_X1   g01176(.A1(new_n3611_), .A2(pi0105), .ZN(new_n3612_));
  AOI21_X1   g01177(.A1(new_n3612_), .A2(new_n3609_), .B(new_n2458_), .ZN(new_n3613_));
  NOR2_X1    g01178(.A1(new_n3613_), .A2(new_n3302_), .ZN(new_n3614_));
  INV_X1     g01179(.I(new_n3614_), .ZN(new_n3615_));
  AOI21_X1   g01180(.A1(new_n3107_), .A2(new_n2458_), .B(new_n3615_), .ZN(new_n3616_));
  OAI21_X1   g01181(.A1(new_n3616_), .A2(pi0216), .B(new_n3608_), .ZN(new_n3617_));
  NAND3_X1   g01182(.A1(new_n3617_), .A2(new_n2436_), .A3(new_n3607_), .ZN(new_n3618_));
  NOR2_X1    g01183(.A1(new_n2436_), .A2(pi1143), .ZN(new_n3619_));
  INV_X1     g01184(.I(new_n3619_), .ZN(new_n3620_));
  NAND2_X1   g01185(.A1(new_n3618_), .A2(new_n3620_), .ZN(new_n3621_));
  AOI21_X1   g01186(.A1(pi0216), .A2(pi0264), .B(new_n3502_), .ZN(new_n3622_));
  NAND2_X1   g01187(.A1(new_n3622_), .A2(pi0238), .ZN(new_n3623_));
  AND3_X2    g01188(.A1(new_n3621_), .A2(new_n3425_), .A3(new_n3623_), .Z(new_n3624_));
  INV_X1     g01189(.I(pi0238), .ZN(new_n3625_));
  INV_X1     g01190(.I(new_n3607_), .ZN(new_n3626_));
  INV_X1     g01191(.I(new_n3608_), .ZN(new_n3627_));
  NOR2_X1    g01192(.A1(new_n2531_), .A2(pi0146), .ZN(new_n3628_));
  NOR2_X1    g01193(.A1(new_n2530_), .A2(new_n3610_), .ZN(new_n3629_));
  OAI21_X1   g01194(.A1(new_n3628_), .A2(new_n3629_), .B(new_n2458_), .ZN(new_n3630_));
  AOI21_X1   g01195(.A1(new_n3630_), .A2(new_n3614_), .B(pi0216), .ZN(new_n3631_));
  OAI21_X1   g01196(.A1(new_n3631_), .A2(new_n3627_), .B(new_n2436_), .ZN(new_n3632_));
  OAI21_X1   g01197(.A1(new_n3632_), .A2(new_n3626_), .B(new_n3620_), .ZN(new_n3633_));
  INV_X1     g01198(.I(new_n3621_), .ZN(new_n3634_));
  NAND2_X1   g01199(.A1(new_n3634_), .A2(new_n3472_), .ZN(new_n3635_));
  OAI21_X1   g01200(.A1(new_n3633_), .A2(new_n3472_), .B(new_n3635_), .ZN(new_n3636_));
  NAND2_X1   g01201(.A1(new_n3636_), .A2(pi0062), .ZN(new_n3637_));
  NAND3_X1   g01202(.A1(new_n3637_), .A2(new_n3625_), .A3(new_n3291_), .ZN(new_n3638_));
  NAND2_X1   g01203(.A1(new_n3634_), .A2(new_n2612_), .ZN(new_n3639_));
  OAI21_X1   g01204(.A1(new_n3633_), .A2(new_n2612_), .B(new_n3639_), .ZN(new_n3640_));
  NAND2_X1   g01205(.A1(new_n3640_), .A2(pi0055), .ZN(new_n3641_));
  NOR2_X1    g01206(.A1(new_n2635_), .A2(new_n3603_), .ZN(new_n3642_));
  NOR2_X1    g01207(.A1(new_n2634_), .A2(new_n3605_), .ZN(new_n3643_));
  OAI21_X1   g01208(.A1(new_n3642_), .A2(new_n3643_), .B(pi0222), .ZN(new_n3644_));
  AOI21_X1   g01209(.A1(pi0224), .A2(pi0264), .B(pi0222), .ZN(new_n3645_));
  NAND2_X1   g01210(.A1(new_n3611_), .A2(new_n2631_), .ZN(new_n3646_));
  NAND2_X1   g01211(.A1(new_n3646_), .A2(new_n3645_), .ZN(new_n3647_));
  NAND2_X1   g01212(.A1(new_n3644_), .A2(new_n3647_), .ZN(new_n3648_));
  NAND2_X1   g01213(.A1(new_n3648_), .A2(new_n2668_), .ZN(new_n3649_));
  NAND2_X1   g01214(.A1(pi0223), .A2(pi1143), .ZN(new_n3650_));
  AOI21_X1   g01215(.A1(new_n3649_), .A2(new_n3650_), .B(pi0299), .ZN(new_n3651_));
  INV_X1     g01216(.I(new_n3651_), .ZN(new_n3652_));
  NOR2_X1    g01217(.A1(new_n2644_), .A2(new_n3028_), .ZN(new_n3653_));
  NOR2_X1    g01218(.A1(new_n3652_), .A2(new_n3653_), .ZN(new_n3654_));
  AOI21_X1   g01219(.A1(new_n3634_), .A2(pi0299), .B(new_n3654_), .ZN(new_n3655_));
  AOI21_X1   g01220(.A1(new_n3655_), .A2(new_n2563_), .B(pi0055), .ZN(new_n3656_));
  INV_X1     g01221(.I(new_n3451_), .ZN(new_n3657_));
  NAND2_X1   g01222(.A1(new_n3657_), .A2(pi0146), .ZN(new_n3658_));
  NOR2_X1    g01223(.A1(new_n3107_), .A2(pi0284), .ZN(new_n3659_));
  AOI22_X1   g01224(.A1(new_n3658_), .A2(pi0284), .B1(new_n3387_), .B2(new_n3659_), .ZN(new_n3660_));
  NAND2_X1   g01225(.A1(new_n3404_), .A2(new_n3107_), .ZN(new_n3661_));
  AOI21_X1   g01226(.A1(new_n3660_), .A2(new_n3661_), .B(pi0228), .ZN(new_n3662_));
  NOR3_X1    g01227(.A1(new_n3662_), .A2(new_n3388_), .A3(new_n3613_), .ZN(new_n3663_));
  OAI21_X1   g01228(.A1(new_n3663_), .A2(pi0216), .B(new_n3608_), .ZN(new_n3664_));
  NAND3_X1   g01229(.A1(new_n3664_), .A2(new_n2436_), .A3(new_n3607_), .ZN(new_n3665_));
  AOI21_X1   g01230(.A1(new_n3665_), .A2(new_n3620_), .B(new_n2628_), .ZN(new_n3666_));
  NAND2_X1   g01231(.A1(new_n3650_), .A2(new_n2628_), .ZN(new_n3667_));
  INV_X1     g01232(.I(new_n3644_), .ZN(new_n3668_));
  OAI21_X1   g01233(.A1(new_n3392_), .A2(pi0284), .B(new_n2631_), .ZN(new_n3669_));
  AOI21_X1   g01234(.A1(new_n3669_), .A2(new_n3645_), .B(new_n3668_), .ZN(new_n3670_));
  INV_X1     g01235(.I(new_n3670_), .ZN(new_n3671_));
  INV_X1     g01236(.I(new_n3667_), .ZN(new_n3672_));
  AOI21_X1   g01237(.A1(new_n3392_), .A2(new_n3645_), .B(new_n3671_), .ZN(new_n3673_));
  OAI21_X1   g01238(.A1(new_n3673_), .A2(pi0223), .B(new_n3672_), .ZN(new_n3674_));
  NAND2_X1   g01239(.A1(new_n3674_), .A2(new_n2627_), .ZN(new_n3675_));
  INV_X1     g01240(.I(new_n3675_), .ZN(new_n3676_));
  OAI21_X1   g01241(.A1(new_n3667_), .A2(new_n3671_), .B(new_n3676_), .ZN(new_n3677_));
  OAI22_X1   g01242(.A1(new_n3633_), .A2(new_n2628_), .B1(new_n3652_), .B2(new_n3653_), .ZN(new_n3678_));
  NAND2_X1   g01243(.A1(new_n3678_), .A2(pi0039), .ZN(new_n3679_));
  OAI21_X1   g01244(.A1(new_n3666_), .A2(new_n3677_), .B(new_n3679_), .ZN(new_n3680_));
  AOI21_X1   g01245(.A1(new_n3655_), .A2(pi0038), .B(pi0100), .ZN(new_n3681_));
  OAI21_X1   g01246(.A1(new_n3680_), .A2(pi0038), .B(new_n3681_), .ZN(new_n3682_));
  AOI21_X1   g01247(.A1(new_n3655_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n3683_));
  NAND2_X1   g01248(.A1(new_n2690_), .A2(pi0252), .ZN(new_n3684_));
  NAND3_X1   g01249(.A1(new_n2531_), .A2(new_n3610_), .A3(new_n3684_), .ZN(new_n3685_));
  NAND2_X1   g01250(.A1(new_n3363_), .A2(pi0146), .ZN(new_n3686_));
  NAND3_X1   g01251(.A1(new_n3686_), .A2(new_n2458_), .A3(new_n3685_), .ZN(new_n3687_));
  AOI21_X1   g01252(.A1(new_n3687_), .A2(new_n3614_), .B(pi0216), .ZN(new_n3688_));
  OAI21_X1   g01253(.A1(new_n3688_), .A2(new_n3627_), .B(new_n2436_), .ZN(new_n3689_));
  OAI21_X1   g01254(.A1(new_n3689_), .A2(new_n3626_), .B(new_n3620_), .ZN(new_n3690_));
  OAI21_X1   g01255(.A1(new_n3690_), .A2(new_n2628_), .B(new_n2572_), .ZN(new_n3691_));
  OAI21_X1   g01256(.A1(new_n3691_), .A2(new_n3654_), .B(new_n3683_), .ZN(new_n3692_));
  NAND3_X1   g01257(.A1(new_n3682_), .A2(new_n3458_), .A3(new_n3692_), .ZN(new_n3693_));
  NOR2_X1    g01258(.A1(new_n3655_), .A2(new_n3272_), .ZN(new_n3694_));
  AOI21_X1   g01259(.A1(new_n3678_), .A2(new_n3272_), .B(new_n3694_), .ZN(new_n3695_));
  NAND2_X1   g01260(.A1(new_n3695_), .A2(pi0087), .ZN(new_n3696_));
  AOI21_X1   g01261(.A1(new_n3693_), .A2(new_n3696_), .B(pi0075), .ZN(new_n3697_));
  INV_X1     g01262(.I(new_n3655_), .ZN(new_n3698_));
  OAI21_X1   g01263(.A1(new_n3698_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n3699_));
  NOR2_X1    g01264(.A1(new_n3695_), .A2(new_n2565_), .ZN(new_n3700_));
  AOI21_X1   g01265(.A1(new_n2565_), .A2(new_n3698_), .B(new_n3700_), .ZN(new_n3701_));
  OAI22_X1   g01266(.A1(new_n3697_), .A2(new_n3699_), .B1(new_n3444_), .B2(new_n3701_), .ZN(new_n3702_));
  OAI21_X1   g01267(.A1(new_n3702_), .A2(new_n2563_), .B(new_n3656_), .ZN(new_n3703_));
  NAND3_X1   g01268(.A1(new_n3703_), .A2(new_n3284_), .A3(new_n3641_), .ZN(new_n3704_));
  NAND2_X1   g01269(.A1(new_n3633_), .A2(new_n2576_), .ZN(new_n3705_));
  OAI21_X1   g01270(.A1(new_n2576_), .A2(new_n3634_), .B(new_n3705_), .ZN(new_n3706_));
  AOI21_X1   g01271(.A1(new_n3706_), .A2(pi0056), .B(pi0062), .ZN(new_n3707_));
  AOI21_X1   g01272(.A1(new_n3704_), .A2(new_n3707_), .B(new_n3638_), .ZN(new_n3708_));
  INV_X1     g01273(.I(new_n3613_), .ZN(new_n3709_));
  AOI21_X1   g01274(.A1(new_n3630_), .A2(new_n3709_), .B(pi0216), .ZN(new_n3710_));
  OAI21_X1   g01275(.A1(new_n3710_), .A2(new_n3627_), .B(new_n2436_), .ZN(new_n3711_));
  OAI21_X1   g01276(.A1(new_n3711_), .A2(new_n3626_), .B(new_n3620_), .ZN(new_n3712_));
  NOR2_X1    g01277(.A1(new_n3712_), .A2(new_n3472_), .ZN(new_n3713_));
  NOR2_X1    g01278(.A1(new_n3634_), .A2(new_n3622_), .ZN(new_n3714_));
  NOR2_X1    g01279(.A1(new_n3714_), .A2(new_n3320_), .ZN(new_n3715_));
  OAI21_X1   g01280(.A1(new_n3713_), .A2(new_n3715_), .B(pi0062), .ZN(new_n3716_));
  NAND3_X1   g01281(.A1(new_n3716_), .A2(pi0238), .A3(new_n3291_), .ZN(new_n3717_));
  NOR2_X1    g01282(.A1(new_n3712_), .A2(new_n2612_), .ZN(new_n3718_));
  NOR2_X1    g01283(.A1(new_n3714_), .A2(new_n2611_), .ZN(new_n3719_));
  OAI21_X1   g01284(.A1(new_n3718_), .A2(new_n3719_), .B(pi0055), .ZN(new_n3720_));
  OAI21_X1   g01285(.A1(new_n3714_), .A2(new_n2628_), .B(new_n3652_), .ZN(new_n3721_));
  INV_X1     g01286(.I(new_n3721_), .ZN(new_n3722_));
  AOI21_X1   g01287(.A1(new_n3722_), .A2(new_n2563_), .B(pi0055), .ZN(new_n3723_));
  AOI21_X1   g01288(.A1(new_n3722_), .A2(pi0038), .B(pi0100), .ZN(new_n3724_));
  INV_X1     g01289(.I(new_n3712_), .ZN(new_n3725_));
  AOI21_X1   g01290(.A1(new_n3725_), .A2(pi0299), .B(new_n3651_), .ZN(new_n3726_));
  OAI21_X1   g01291(.A1(new_n3726_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n3727_));
  NOR2_X1    g01292(.A1(new_n3381_), .A2(new_n2457_), .ZN(new_n3728_));
  INV_X1     g01293(.I(new_n3728_), .ZN(new_n3729_));
  NAND2_X1   g01294(.A1(new_n3729_), .A2(new_n3613_), .ZN(new_n3730_));
  INV_X1     g01295(.I(new_n3387_), .ZN(new_n3731_));
  NAND2_X1   g01296(.A1(new_n3731_), .A2(new_n3107_), .ZN(new_n3732_));
  NAND2_X1   g01297(.A1(new_n3403_), .A2(pi0146), .ZN(new_n3733_));
  AOI21_X1   g01298(.A1(new_n3733_), .A2(new_n3732_), .B(new_n3610_), .ZN(new_n3734_));
  NOR3_X1    g01299(.A1(new_n3451_), .A2(pi0146), .A3(pi0284), .ZN(new_n3735_));
  OAI21_X1   g01300(.A1(new_n3734_), .A2(new_n3735_), .B(new_n2458_), .ZN(new_n3736_));
  AOI21_X1   g01301(.A1(new_n3736_), .A2(new_n3730_), .B(pi0216), .ZN(new_n3737_));
  OAI21_X1   g01302(.A1(new_n3737_), .A2(new_n3627_), .B(new_n3607_), .ZN(new_n3738_));
  OAI21_X1   g01303(.A1(new_n3738_), .A2(pi0215), .B(new_n3620_), .ZN(new_n3739_));
  AOI21_X1   g01304(.A1(new_n3739_), .A2(pi0299), .B(new_n3675_), .ZN(new_n3740_));
  OAI21_X1   g01305(.A1(new_n3740_), .A2(new_n3727_), .B(new_n3724_), .ZN(new_n3741_));
  AOI21_X1   g01306(.A1(new_n3722_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n3742_));
  AOI21_X1   g01307(.A1(new_n3687_), .A2(new_n3709_), .B(pi0216), .ZN(new_n3743_));
  OAI21_X1   g01308(.A1(new_n3743_), .A2(new_n3627_), .B(new_n2436_), .ZN(new_n3744_));
  OAI21_X1   g01309(.A1(new_n3744_), .A2(new_n3626_), .B(new_n3620_), .ZN(new_n3745_));
  OAI21_X1   g01310(.A1(new_n3745_), .A2(new_n2628_), .B(new_n2572_), .ZN(new_n3746_));
  OAI21_X1   g01311(.A1(new_n3746_), .A2(new_n3651_), .B(new_n3742_), .ZN(new_n3747_));
  NAND3_X1   g01312(.A1(new_n3741_), .A2(new_n3458_), .A3(new_n3747_), .ZN(new_n3748_));
  NOR2_X1    g01313(.A1(new_n3726_), .A2(new_n3273_), .ZN(new_n3749_));
  AOI21_X1   g01314(.A1(new_n3273_), .A2(new_n3721_), .B(new_n3749_), .ZN(new_n3750_));
  NAND2_X1   g01315(.A1(new_n3750_), .A2(pi0087), .ZN(new_n3751_));
  AOI21_X1   g01316(.A1(new_n3748_), .A2(new_n3751_), .B(pi0075), .ZN(new_n3752_));
  OAI21_X1   g01317(.A1(new_n3721_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n3753_));
  NOR2_X1    g01318(.A1(new_n3750_), .A2(new_n2565_), .ZN(new_n3754_));
  AOI21_X1   g01319(.A1(new_n2565_), .A2(new_n3721_), .B(new_n3754_), .ZN(new_n3755_));
  OAI22_X1   g01320(.A1(new_n3752_), .A2(new_n3753_), .B1(new_n3444_), .B2(new_n3755_), .ZN(new_n3756_));
  OAI21_X1   g01321(.A1(new_n3756_), .A2(new_n2563_), .B(new_n3723_), .ZN(new_n3757_));
  NAND3_X1   g01322(.A1(new_n3757_), .A2(new_n3284_), .A3(new_n3720_), .ZN(new_n3758_));
  NAND2_X1   g01323(.A1(new_n3714_), .A2(new_n2577_), .ZN(new_n3759_));
  OAI21_X1   g01324(.A1(new_n3725_), .A2(new_n2577_), .B(new_n3759_), .ZN(new_n3760_));
  AOI21_X1   g01325(.A1(new_n3760_), .A2(pi0056), .B(pi0062), .ZN(new_n3761_));
  AOI21_X1   g01326(.A1(new_n3758_), .A2(new_n3761_), .B(new_n3717_), .ZN(new_n3762_));
  NOR3_X1    g01327(.A1(new_n3708_), .A2(new_n3624_), .A3(new_n3762_), .ZN(po0156));
  NOR2_X1    g01328(.A1(new_n2436_), .A2(pi1142), .ZN(new_n3764_));
  INV_X1     g01329(.I(new_n3764_), .ZN(new_n3765_));
  INV_X1     g01330(.I(pi0932), .ZN(new_n3766_));
  NOR2_X1    g01331(.A1(new_n2447_), .A2(new_n3766_), .ZN(new_n3767_));
  INV_X1     g01332(.I(pi1142), .ZN(new_n3768_));
  NOR2_X1    g01333(.A1(new_n2444_), .A2(new_n3768_), .ZN(new_n3769_));
  OAI21_X1   g01334(.A1(new_n3767_), .A2(new_n3769_), .B(pi0221), .ZN(new_n3770_));
  INV_X1     g01335(.I(new_n3770_), .ZN(new_n3771_));
  AOI21_X1   g01336(.A1(pi0216), .A2(pi0277), .B(pi0221), .ZN(new_n3772_));
  INV_X1     g01337(.I(new_n3772_), .ZN(new_n3773_));
  INV_X1     g01338(.I(pi0262), .ZN(new_n3774_));
  NOR2_X1    g01339(.A1(new_n2463_), .A2(new_n3774_), .ZN(new_n3775_));
  INV_X1     g01340(.I(new_n3775_), .ZN(new_n3776_));
  NOR2_X1    g01341(.A1(new_n3776_), .A2(new_n2457_), .ZN(new_n3777_));
  INV_X1     g01342(.I(pi0172), .ZN(new_n3778_));
  NOR2_X1    g01343(.A1(new_n3778_), .A2(pi0105), .ZN(new_n3779_));
  OAI21_X1   g01344(.A1(new_n3777_), .A2(new_n3779_), .B(pi0228), .ZN(new_n3780_));
  NAND2_X1   g01345(.A1(new_n2531_), .A2(pi0262), .ZN(new_n3781_));
  NAND2_X1   g01346(.A1(new_n2530_), .A2(pi0172), .ZN(new_n3782_));
  AOI21_X1   g01347(.A1(new_n3781_), .A2(new_n3782_), .B(pi0228), .ZN(new_n3783_));
  INV_X1     g01348(.I(new_n3783_), .ZN(new_n3784_));
  AOI21_X1   g01349(.A1(new_n3784_), .A2(new_n3780_), .B(pi0216), .ZN(new_n3785_));
  OAI21_X1   g01350(.A1(new_n3785_), .A2(new_n3773_), .B(new_n2436_), .ZN(new_n3786_));
  OAI21_X1   g01351(.A1(new_n3786_), .A2(new_n3771_), .B(new_n3765_), .ZN(new_n3787_));
  INV_X1     g01352(.I(new_n3780_), .ZN(new_n3788_));
  AOI21_X1   g01353(.A1(pi0172), .A2(new_n2458_), .B(new_n3788_), .ZN(new_n3789_));
  OAI21_X1   g01354(.A1(new_n3789_), .A2(pi0216), .B(new_n3772_), .ZN(new_n3790_));
  NAND3_X1   g01355(.A1(new_n3790_), .A2(new_n2436_), .A3(new_n3770_), .ZN(new_n3791_));
  NAND2_X1   g01356(.A1(new_n3791_), .A2(new_n3765_), .ZN(new_n3792_));
  INV_X1     g01357(.I(new_n3792_), .ZN(new_n3793_));
  NAND2_X1   g01358(.A1(new_n3793_), .A2(new_n2612_), .ZN(new_n3794_));
  OAI21_X1   g01359(.A1(new_n3787_), .A2(new_n2612_), .B(new_n3794_), .ZN(new_n3795_));
  NAND2_X1   g01360(.A1(new_n3795_), .A2(pi0055), .ZN(new_n3796_));
  NOR2_X1    g01361(.A1(new_n2635_), .A2(new_n3766_), .ZN(new_n3797_));
  NOR2_X1    g01362(.A1(new_n2634_), .A2(new_n3768_), .ZN(new_n3798_));
  OAI21_X1   g01363(.A1(new_n3797_), .A2(new_n3798_), .B(pi0222), .ZN(new_n3799_));
  AOI21_X1   g01364(.A1(pi0224), .A2(pi0277), .B(pi0222), .ZN(new_n3800_));
  OAI21_X1   g01365(.A1(new_n3776_), .A2(pi0224), .B(new_n3800_), .ZN(new_n3801_));
  NAND2_X1   g01366(.A1(new_n3799_), .A2(new_n3801_), .ZN(new_n3802_));
  NAND2_X1   g01367(.A1(new_n3802_), .A2(new_n2668_), .ZN(new_n3803_));
  NAND2_X1   g01368(.A1(pi0223), .A2(pi1142), .ZN(new_n3804_));
  AOI21_X1   g01369(.A1(new_n3803_), .A2(new_n3804_), .B(pi0299), .ZN(new_n3805_));
  AOI21_X1   g01370(.A1(new_n3793_), .A2(pi0299), .B(new_n3805_), .ZN(new_n3806_));
  AOI21_X1   g01371(.A1(new_n3806_), .A2(new_n2563_), .B(pi0055), .ZN(new_n3807_));
  AOI21_X1   g01372(.A1(new_n3806_), .A2(pi0038), .B(pi0100), .ZN(new_n3808_));
  INV_X1     g01373(.I(new_n3787_), .ZN(new_n3809_));
  AOI21_X1   g01374(.A1(new_n3809_), .A2(pi0299), .B(new_n3805_), .ZN(new_n3810_));
  OAI21_X1   g01375(.A1(new_n3810_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n3811_));
  INV_X1     g01376(.I(new_n3380_), .ZN(new_n3812_));
  NOR2_X1    g01377(.A1(new_n3779_), .A2(new_n2458_), .ZN(new_n3813_));
  INV_X1     g01378(.I(new_n3813_), .ZN(new_n3814_));
  AOI21_X1   g01379(.A1(new_n3812_), .A2(new_n3777_), .B(new_n3814_), .ZN(new_n3815_));
  NOR2_X1    g01380(.A1(new_n3731_), .A2(new_n3774_), .ZN(new_n3816_));
  NOR2_X1    g01381(.A1(new_n3657_), .A2(pi0262), .ZN(new_n3817_));
  OAI21_X1   g01382(.A1(new_n3817_), .A2(new_n3816_), .B(pi0172), .ZN(new_n3818_));
  OAI21_X1   g01383(.A1(new_n3404_), .A2(new_n3774_), .B(new_n3778_), .ZN(new_n3819_));
  AOI21_X1   g01384(.A1(new_n3818_), .A2(new_n3819_), .B(pi0228), .ZN(new_n3820_));
  NOR3_X1    g01385(.A1(new_n3820_), .A2(pi0216), .A3(new_n3815_), .ZN(new_n3821_));
  OAI21_X1   g01386(.A1(new_n3821_), .A2(new_n3773_), .B(new_n3770_), .ZN(new_n3822_));
  OAI21_X1   g01387(.A1(new_n3822_), .A2(pi0215), .B(new_n3765_), .ZN(new_n3823_));
  NAND2_X1   g01388(.A1(new_n3804_), .A2(new_n2628_), .ZN(new_n3824_));
  INV_X1     g01389(.I(new_n3824_), .ZN(new_n3825_));
  INV_X1     g01390(.I(new_n3799_), .ZN(new_n3826_));
  OAI21_X1   g01391(.A1(new_n3392_), .A2(pi0262), .B(new_n2631_), .ZN(new_n3827_));
  AOI21_X1   g01392(.A1(new_n3827_), .A2(new_n3800_), .B(new_n3826_), .ZN(new_n3828_));
  INV_X1     g01393(.I(new_n3828_), .ZN(new_n3829_));
  AOI21_X1   g01394(.A1(new_n3392_), .A2(new_n3800_), .B(new_n3829_), .ZN(new_n3830_));
  OAI21_X1   g01395(.A1(new_n3830_), .A2(pi0223), .B(new_n3825_), .ZN(new_n3831_));
  NAND2_X1   g01396(.A1(new_n3831_), .A2(new_n2627_), .ZN(new_n3832_));
  AOI21_X1   g01397(.A1(new_n3823_), .A2(pi0299), .B(new_n3832_), .ZN(new_n3833_));
  OAI21_X1   g01398(.A1(new_n3833_), .A2(new_n3811_), .B(new_n3808_), .ZN(new_n3834_));
  AOI21_X1   g01399(.A1(new_n3806_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n3835_));
  NOR2_X1    g01400(.A1(new_n3544_), .A2(new_n3774_), .ZN(new_n3836_));
  NOR2_X1    g01401(.A1(new_n3371_), .A2(new_n3778_), .ZN(new_n3837_));
  OAI21_X1   g01402(.A1(new_n3836_), .A2(new_n3837_), .B(new_n2458_), .ZN(new_n3838_));
  AOI21_X1   g01403(.A1(new_n3838_), .A2(new_n3780_), .B(pi0216), .ZN(new_n3839_));
  OAI21_X1   g01404(.A1(new_n3839_), .A2(new_n3773_), .B(new_n2436_), .ZN(new_n3840_));
  OAI21_X1   g01405(.A1(new_n3840_), .A2(new_n3771_), .B(new_n3765_), .ZN(new_n3841_));
  OAI21_X1   g01406(.A1(new_n3841_), .A2(new_n2628_), .B(new_n2572_), .ZN(new_n3842_));
  OAI21_X1   g01407(.A1(new_n3842_), .A2(new_n3805_), .B(new_n3835_), .ZN(new_n3843_));
  NAND3_X1   g01408(.A1(new_n3834_), .A2(new_n3458_), .A3(new_n3843_), .ZN(new_n3844_));
  INV_X1     g01409(.I(new_n3806_), .ZN(new_n3845_));
  NOR2_X1    g01410(.A1(new_n3810_), .A2(new_n3273_), .ZN(new_n3846_));
  AOI21_X1   g01411(.A1(new_n3273_), .A2(new_n3845_), .B(new_n3846_), .ZN(new_n3847_));
  NAND2_X1   g01412(.A1(new_n3847_), .A2(pi0087), .ZN(new_n3848_));
  AOI21_X1   g01413(.A1(new_n3844_), .A2(new_n3848_), .B(pi0075), .ZN(new_n3849_));
  OAI21_X1   g01414(.A1(new_n3845_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n3850_));
  NOR2_X1    g01415(.A1(new_n3847_), .A2(new_n2565_), .ZN(new_n3851_));
  AOI21_X1   g01416(.A1(new_n2565_), .A2(new_n3845_), .B(new_n3851_), .ZN(new_n3852_));
  OAI22_X1   g01417(.A1(new_n3849_), .A2(new_n3850_), .B1(new_n3444_), .B2(new_n3852_), .ZN(new_n3853_));
  OAI21_X1   g01418(.A1(new_n3853_), .A2(new_n2563_), .B(new_n3807_), .ZN(new_n3854_));
  NAND3_X1   g01419(.A1(new_n3854_), .A2(new_n3284_), .A3(new_n3796_), .ZN(new_n3855_));
  NOR2_X1    g01420(.A1(new_n3809_), .A2(new_n2577_), .ZN(new_n3856_));
  NOR2_X1    g01421(.A1(new_n3793_), .A2(new_n2576_), .ZN(new_n3857_));
  OAI21_X1   g01422(.A1(new_n3856_), .A2(new_n3857_), .B(pi0056), .ZN(new_n3858_));
  NAND3_X1   g01423(.A1(new_n3855_), .A2(new_n3471_), .A3(new_n3858_), .ZN(new_n3859_));
  NAND2_X1   g01424(.A1(new_n3793_), .A2(new_n3472_), .ZN(new_n3860_));
  OAI21_X1   g01425(.A1(new_n3787_), .A2(new_n3472_), .B(new_n3860_), .ZN(new_n3861_));
  NAND2_X1   g01426(.A1(new_n3861_), .A2(pi0062), .ZN(new_n3862_));
  AND3_X2    g01427(.A1(new_n3859_), .A2(new_n3291_), .A3(new_n3862_), .Z(new_n3863_));
  OAI21_X1   g01428(.A1(new_n3793_), .A2(new_n3291_), .B(pi0249), .ZN(new_n3864_));
  INV_X1     g01429(.I(pi0249), .ZN(new_n3865_));
  NOR2_X1    g01430(.A1(new_n3788_), .A2(new_n3302_), .ZN(new_n3866_));
  AOI21_X1   g01431(.A1(new_n3784_), .A2(new_n3866_), .B(pi0216), .ZN(new_n3867_));
  OAI21_X1   g01432(.A1(new_n3867_), .A2(new_n3773_), .B(new_n2436_), .ZN(new_n3868_));
  OAI21_X1   g01433(.A1(new_n3868_), .A2(new_n3771_), .B(new_n3765_), .ZN(new_n3869_));
  NOR2_X1    g01434(.A1(new_n3792_), .A2(new_n3307_), .ZN(new_n3870_));
  NAND2_X1   g01435(.A1(new_n3870_), .A2(new_n2612_), .ZN(new_n3871_));
  OAI21_X1   g01436(.A1(new_n3869_), .A2(new_n2612_), .B(new_n3871_), .ZN(new_n3872_));
  NAND2_X1   g01437(.A1(new_n3872_), .A2(pi0055), .ZN(new_n3873_));
  INV_X1     g01438(.I(new_n3653_), .ZN(new_n3874_));
  NAND2_X1   g01439(.A1(new_n3805_), .A2(new_n3874_), .ZN(new_n3875_));
  INV_X1     g01440(.I(new_n3875_), .ZN(new_n3876_));
  AOI21_X1   g01441(.A1(new_n3870_), .A2(pi0299), .B(new_n3876_), .ZN(new_n3877_));
  AOI21_X1   g01442(.A1(new_n3877_), .A2(new_n2563_), .B(pi0055), .ZN(new_n3878_));
  NOR3_X1    g01443(.A1(new_n3731_), .A2(pi0172), .A3(pi0262), .ZN(new_n3879_));
  AOI21_X1   g01444(.A1(new_n3403_), .A2(new_n3774_), .B(new_n3778_), .ZN(new_n3880_));
  NOR2_X1    g01445(.A1(new_n3657_), .A2(new_n3774_), .ZN(new_n3881_));
  NOR4_X1    g01446(.A1(new_n3881_), .A2(pi0228), .A3(new_n3879_), .A4(new_n3880_), .ZN(new_n3882_));
  NAND2_X1   g01447(.A1(new_n3729_), .A2(new_n3815_), .ZN(new_n3883_));
  NAND2_X1   g01448(.A1(new_n3883_), .A2(new_n2614_), .ZN(new_n3884_));
  OAI21_X1   g01449(.A1(new_n3882_), .A2(new_n3884_), .B(new_n3772_), .ZN(new_n3885_));
  NAND3_X1   g01450(.A1(new_n3885_), .A2(new_n2436_), .A3(new_n3770_), .ZN(new_n3886_));
  AOI21_X1   g01451(.A1(new_n3886_), .A2(new_n3765_), .B(new_n2628_), .ZN(new_n3887_));
  INV_X1     g01452(.I(new_n3832_), .ZN(new_n3888_));
  OAI21_X1   g01453(.A1(new_n3824_), .A2(new_n3829_), .B(new_n3888_), .ZN(new_n3889_));
  OAI21_X1   g01454(.A1(new_n3869_), .A2(new_n2628_), .B(new_n3875_), .ZN(new_n3890_));
  NAND2_X1   g01455(.A1(new_n3890_), .A2(pi0039), .ZN(new_n3891_));
  OAI21_X1   g01456(.A1(new_n3887_), .A2(new_n3889_), .B(new_n3891_), .ZN(new_n3892_));
  AOI21_X1   g01457(.A1(new_n3877_), .A2(pi0038), .B(pi0100), .ZN(new_n3893_));
  OAI21_X1   g01458(.A1(new_n3892_), .A2(pi0038), .B(new_n3893_), .ZN(new_n3894_));
  AOI21_X1   g01459(.A1(new_n3877_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n3895_));
  AOI21_X1   g01460(.A1(new_n3838_), .A2(new_n3866_), .B(pi0216), .ZN(new_n3896_));
  OAI21_X1   g01461(.A1(new_n3896_), .A2(new_n3773_), .B(new_n2436_), .ZN(new_n3897_));
  OAI21_X1   g01462(.A1(new_n3897_), .A2(new_n3771_), .B(new_n3765_), .ZN(new_n3898_));
  OAI21_X1   g01463(.A1(new_n3898_), .A2(new_n2628_), .B(new_n2572_), .ZN(new_n3899_));
  OAI21_X1   g01464(.A1(new_n3899_), .A2(new_n3876_), .B(new_n3895_), .ZN(new_n3900_));
  NAND3_X1   g01465(.A1(new_n3894_), .A2(new_n3458_), .A3(new_n3900_), .ZN(new_n3901_));
  NOR2_X1    g01466(.A1(new_n3877_), .A2(new_n3272_), .ZN(new_n3902_));
  AOI21_X1   g01467(.A1(new_n3890_), .A2(new_n3272_), .B(new_n3902_), .ZN(new_n3903_));
  NAND2_X1   g01468(.A1(new_n3903_), .A2(pi0087), .ZN(new_n3904_));
  AOI21_X1   g01469(.A1(new_n3901_), .A2(new_n3904_), .B(pi0075), .ZN(new_n3905_));
  INV_X1     g01470(.I(new_n3877_), .ZN(new_n3906_));
  OAI21_X1   g01471(.A1(new_n3906_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n3907_));
  NOR2_X1    g01472(.A1(new_n3903_), .A2(new_n2565_), .ZN(new_n3908_));
  AOI21_X1   g01473(.A1(new_n2565_), .A2(new_n3906_), .B(new_n3908_), .ZN(new_n3909_));
  OAI22_X1   g01474(.A1(new_n3905_), .A2(new_n3907_), .B1(new_n3444_), .B2(new_n3909_), .ZN(new_n3910_));
  OAI21_X1   g01475(.A1(new_n3910_), .A2(new_n2563_), .B(new_n3878_), .ZN(new_n3911_));
  NAND3_X1   g01476(.A1(new_n3911_), .A2(new_n3284_), .A3(new_n3873_), .ZN(new_n3912_));
  NOR2_X1    g01477(.A1(new_n3870_), .A2(new_n2576_), .ZN(new_n3913_));
  AND2_X2    g01478(.A1(new_n3869_), .A2(new_n2576_), .Z(new_n3914_));
  OAI21_X1   g01479(.A1(new_n3914_), .A2(new_n3913_), .B(pi0056), .ZN(new_n3915_));
  NAND3_X1   g01480(.A1(new_n3912_), .A2(new_n3471_), .A3(new_n3915_), .ZN(new_n3916_));
  NAND2_X1   g01481(.A1(new_n3870_), .A2(new_n3472_), .ZN(new_n3917_));
  OAI21_X1   g01482(.A1(new_n3869_), .A2(new_n3472_), .B(new_n3917_), .ZN(new_n3918_));
  NAND2_X1   g01483(.A1(new_n3918_), .A2(pi0062), .ZN(new_n3919_));
  NAND3_X1   g01484(.A1(new_n3916_), .A2(new_n3291_), .A3(new_n3919_), .ZN(new_n3920_));
  OAI21_X1   g01485(.A1(new_n3792_), .A2(new_n3307_), .B(new_n3425_), .ZN(new_n3921_));
  NAND3_X1   g01486(.A1(new_n3920_), .A2(new_n3865_), .A3(new_n3921_), .ZN(new_n3922_));
  OAI21_X1   g01487(.A1(new_n3863_), .A2(new_n3864_), .B(new_n3922_), .ZN(po0157));
  INV_X1     g01488(.I(pi0935), .ZN(new_n3924_));
  NOR2_X1    g01489(.A1(new_n2447_), .A2(new_n3924_), .ZN(new_n3925_));
  INV_X1     g01490(.I(pi1141), .ZN(new_n3926_));
  NOR2_X1    g01491(.A1(new_n2444_), .A2(new_n3926_), .ZN(new_n3927_));
  OAI21_X1   g01492(.A1(new_n3925_), .A2(new_n3927_), .B(pi0221), .ZN(new_n3928_));
  INV_X1     g01493(.I(new_n3928_), .ZN(new_n3929_));
  AOI21_X1   g01494(.A1(pi0216), .A2(pi0270), .B(pi0221), .ZN(new_n3930_));
  INV_X1     g01495(.I(new_n3930_), .ZN(new_n3931_));
  INV_X1     g01496(.I(pi0171), .ZN(new_n3932_));
  NAND2_X1   g01497(.A1(new_n2457_), .A2(new_n3932_), .ZN(new_n3933_));
  INV_X1     g01498(.I(pi0861), .ZN(new_n3934_));
  NOR2_X1    g01499(.A1(new_n2463_), .A2(new_n3934_), .ZN(new_n3935_));
  NAND2_X1   g01500(.A1(new_n3935_), .A2(pi0105), .ZN(new_n3936_));
  AOI21_X1   g01501(.A1(new_n3936_), .A2(new_n3933_), .B(new_n2458_), .ZN(new_n3937_));
  NOR2_X1    g01502(.A1(new_n3937_), .A2(pi0216), .ZN(new_n3938_));
  NAND2_X1   g01503(.A1(new_n3932_), .A2(new_n2458_), .ZN(new_n3939_));
  AOI21_X1   g01504(.A1(new_n3938_), .A2(new_n3939_), .B(new_n3931_), .ZN(new_n3940_));
  NOR3_X1    g01505(.A1(new_n3940_), .A2(pi0215), .A3(new_n3929_), .ZN(new_n3941_));
  NOR2_X1    g01506(.A1(new_n2436_), .A2(pi1141), .ZN(new_n3942_));
  NOR2_X1    g01507(.A1(new_n3941_), .A2(new_n3942_), .ZN(new_n3943_));
  INV_X1     g01508(.I(new_n3943_), .ZN(new_n3944_));
  AOI21_X1   g01509(.A1(pi0216), .A2(pi0270), .B(new_n3502_), .ZN(new_n3945_));
  NAND2_X1   g01510(.A1(new_n3945_), .A2(pi0241), .ZN(new_n3946_));
  AND3_X2    g01511(.A1(new_n3944_), .A2(new_n3425_), .A3(new_n3946_), .Z(new_n3947_));
  INV_X1     g01512(.I(pi0241), .ZN(new_n3948_));
  INV_X1     g01513(.I(new_n3942_), .ZN(new_n3949_));
  INV_X1     g01514(.I(new_n3938_), .ZN(new_n3950_));
  NAND2_X1   g01515(.A1(new_n2530_), .A2(new_n3932_), .ZN(new_n3951_));
  OAI21_X1   g01516(.A1(new_n3934_), .A2(new_n2530_), .B(new_n3951_), .ZN(new_n3952_));
  AOI21_X1   g01517(.A1(new_n3952_), .A2(new_n2458_), .B(new_n3950_), .ZN(new_n3953_));
  OAI21_X1   g01518(.A1(new_n3953_), .A2(new_n3931_), .B(new_n3928_), .ZN(new_n3954_));
  OAI21_X1   g01519(.A1(new_n3954_), .A2(pi0215), .B(new_n3949_), .ZN(new_n3955_));
  NOR2_X1    g01520(.A1(new_n3955_), .A2(new_n3472_), .ZN(new_n3956_));
  NOR2_X1    g01521(.A1(new_n3944_), .A2(new_n3320_), .ZN(new_n3957_));
  OAI21_X1   g01522(.A1(new_n3956_), .A2(new_n3957_), .B(pi0062), .ZN(new_n3958_));
  NAND3_X1   g01523(.A1(new_n3958_), .A2(new_n3948_), .A3(new_n3291_), .ZN(new_n3959_));
  NOR2_X1    g01524(.A1(new_n3955_), .A2(new_n2612_), .ZN(new_n3960_));
  NOR2_X1    g01525(.A1(new_n3944_), .A2(new_n2611_), .ZN(new_n3961_));
  OAI21_X1   g01526(.A1(new_n3960_), .A2(new_n3961_), .B(pi0055), .ZN(new_n3962_));
  NOR2_X1    g01527(.A1(new_n2635_), .A2(new_n3924_), .ZN(new_n3963_));
  NOR2_X1    g01528(.A1(new_n2634_), .A2(new_n3926_), .ZN(new_n3964_));
  OAI21_X1   g01529(.A1(new_n3963_), .A2(new_n3964_), .B(pi0222), .ZN(new_n3965_));
  INV_X1     g01530(.I(new_n3965_), .ZN(new_n3966_));
  AOI21_X1   g01531(.A1(pi0224), .A2(pi0270), .B(pi0222), .ZN(new_n3967_));
  INV_X1     g01532(.I(new_n3967_), .ZN(new_n3968_));
  NOR2_X1    g01533(.A1(new_n3935_), .A2(pi0224), .ZN(new_n3969_));
  NOR2_X1    g01534(.A1(new_n3969_), .A2(new_n3968_), .ZN(new_n3970_));
  OAI21_X1   g01535(.A1(new_n3966_), .A2(new_n3970_), .B(new_n2668_), .ZN(new_n3971_));
  NAND2_X1   g01536(.A1(pi0223), .A2(pi1141), .ZN(new_n3972_));
  AOI21_X1   g01537(.A1(new_n3971_), .A2(new_n3972_), .B(pi0299), .ZN(new_n3973_));
  AOI21_X1   g01538(.A1(new_n3943_), .A2(pi0299), .B(new_n3973_), .ZN(new_n3974_));
  AOI21_X1   g01539(.A1(new_n3974_), .A2(new_n2563_), .B(pi0055), .ZN(new_n3975_));
  NAND2_X1   g01540(.A1(new_n3387_), .A2(pi0861), .ZN(new_n3976_));
  NAND3_X1   g01541(.A1(new_n3657_), .A2(new_n3932_), .A3(new_n3976_), .ZN(new_n3977_));
  NOR2_X1    g01542(.A1(new_n3387_), .A2(pi0171), .ZN(new_n3978_));
  NOR2_X1    g01543(.A1(new_n3404_), .A2(new_n3932_), .ZN(new_n3979_));
  OAI21_X1   g01544(.A1(new_n3979_), .A2(new_n3978_), .B(pi0861), .ZN(new_n3980_));
  AOI21_X1   g01545(.A1(new_n3980_), .A2(new_n3977_), .B(pi0228), .ZN(new_n3981_));
  NAND2_X1   g01546(.A1(new_n3729_), .A2(new_n3937_), .ZN(new_n3982_));
  NAND2_X1   g01547(.A1(new_n3982_), .A2(new_n2614_), .ZN(new_n3983_));
  OAI21_X1   g01548(.A1(new_n3981_), .A2(new_n3983_), .B(new_n3930_), .ZN(new_n3984_));
  NAND3_X1   g01549(.A1(new_n3984_), .A2(new_n2436_), .A3(new_n3928_), .ZN(new_n3985_));
  AOI21_X1   g01550(.A1(new_n3985_), .A2(new_n3949_), .B(new_n2628_), .ZN(new_n3986_));
  NAND2_X1   g01551(.A1(new_n3972_), .A2(new_n2628_), .ZN(new_n3987_));
  OAI21_X1   g01552(.A1(new_n3392_), .A2(new_n3934_), .B(new_n2631_), .ZN(new_n3988_));
  AOI21_X1   g01553(.A1(new_n3988_), .A2(new_n3967_), .B(new_n3966_), .ZN(new_n3989_));
  INV_X1     g01554(.I(new_n3989_), .ZN(new_n3990_));
  INV_X1     g01555(.I(new_n3987_), .ZN(new_n3991_));
  AOI21_X1   g01556(.A1(new_n3392_), .A2(new_n3967_), .B(new_n3990_), .ZN(new_n3992_));
  OAI21_X1   g01557(.A1(new_n3992_), .A2(pi0223), .B(new_n3991_), .ZN(new_n3993_));
  NAND2_X1   g01558(.A1(new_n3993_), .A2(new_n2627_), .ZN(new_n3994_));
  INV_X1     g01559(.I(new_n3994_), .ZN(new_n3995_));
  OAI21_X1   g01560(.A1(new_n3987_), .A2(new_n3990_), .B(new_n3995_), .ZN(new_n3996_));
  INV_X1     g01561(.I(new_n3955_), .ZN(new_n3997_));
  AOI21_X1   g01562(.A1(new_n3997_), .A2(pi0299), .B(new_n3973_), .ZN(new_n3998_));
  OAI22_X1   g01563(.A1(new_n3986_), .A2(new_n3996_), .B1(new_n2627_), .B2(new_n3998_), .ZN(new_n3999_));
  AOI21_X1   g01564(.A1(new_n3974_), .A2(pi0038), .B(pi0100), .ZN(new_n4000_));
  OAI21_X1   g01565(.A1(new_n3999_), .A2(pi0038), .B(new_n4000_), .ZN(new_n4001_));
  AOI21_X1   g01566(.A1(new_n3974_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n4002_));
  INV_X1     g01567(.I(new_n3973_), .ZN(new_n4003_));
  NOR2_X1    g01568(.A1(new_n3942_), .A2(new_n2628_), .ZN(new_n4004_));
  INV_X1     g01569(.I(new_n4004_), .ZN(new_n4005_));
  NOR2_X1    g01570(.A1(new_n3371_), .A2(pi0171), .ZN(new_n4006_));
  NOR2_X1    g01571(.A1(new_n3544_), .A2(new_n3934_), .ZN(new_n4007_));
  OAI21_X1   g01572(.A1(new_n4007_), .A2(new_n4006_), .B(new_n2458_), .ZN(new_n4008_));
  AOI21_X1   g01573(.A1(new_n4008_), .A2(new_n3938_), .B(new_n3931_), .ZN(new_n4009_));
  NOR3_X1    g01574(.A1(new_n4009_), .A2(pi0215), .A3(new_n3929_), .ZN(new_n4010_));
  OAI21_X1   g01575(.A1(new_n4010_), .A2(new_n4005_), .B(new_n4003_), .ZN(new_n4011_));
  OAI21_X1   g01576(.A1(new_n4011_), .A2(new_n2573_), .B(new_n4002_), .ZN(new_n4012_));
  NAND3_X1   g01577(.A1(new_n4001_), .A2(new_n3458_), .A3(new_n4012_), .ZN(new_n4013_));
  INV_X1     g01578(.I(new_n3974_), .ZN(new_n4014_));
  NOR2_X1    g01579(.A1(new_n3998_), .A2(new_n3273_), .ZN(new_n4015_));
  AOI21_X1   g01580(.A1(new_n3273_), .A2(new_n4014_), .B(new_n4015_), .ZN(new_n4016_));
  NAND2_X1   g01581(.A1(new_n4016_), .A2(pi0087), .ZN(new_n4017_));
  AOI21_X1   g01582(.A1(new_n4013_), .A2(new_n4017_), .B(pi0075), .ZN(new_n4018_));
  OAI21_X1   g01583(.A1(new_n4014_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4019_));
  NOR2_X1    g01584(.A1(new_n4016_), .A2(new_n2565_), .ZN(new_n4020_));
  AOI21_X1   g01585(.A1(new_n2565_), .A2(new_n4014_), .B(new_n4020_), .ZN(new_n4021_));
  OAI22_X1   g01586(.A1(new_n4018_), .A2(new_n4019_), .B1(new_n3444_), .B2(new_n4021_), .ZN(new_n4022_));
  OAI21_X1   g01587(.A1(new_n4022_), .A2(new_n2563_), .B(new_n3975_), .ZN(new_n4023_));
  NAND3_X1   g01588(.A1(new_n4023_), .A2(new_n3284_), .A3(new_n3962_), .ZN(new_n4024_));
  NAND2_X1   g01589(.A1(new_n3944_), .A2(new_n2577_), .ZN(new_n4025_));
  OAI21_X1   g01590(.A1(new_n3997_), .A2(new_n2577_), .B(new_n4025_), .ZN(new_n4026_));
  AOI21_X1   g01591(.A1(new_n4026_), .A2(pi0056), .B(pi0062), .ZN(new_n4027_));
  AOI21_X1   g01592(.A1(new_n4024_), .A2(new_n4027_), .B(new_n3959_), .ZN(new_n4028_));
  AOI21_X1   g01593(.A1(new_n3953_), .A2(new_n3500_), .B(new_n3931_), .ZN(new_n4029_));
  NOR3_X1    g01594(.A1(new_n4029_), .A2(pi0215), .A3(new_n3929_), .ZN(new_n4030_));
  NOR2_X1    g01595(.A1(new_n4030_), .A2(new_n3942_), .ZN(new_n4031_));
  INV_X1     g01596(.I(new_n4031_), .ZN(new_n4032_));
  NOR2_X1    g01597(.A1(new_n4032_), .A2(new_n3472_), .ZN(new_n4033_));
  NOR2_X1    g01598(.A1(new_n3943_), .A2(new_n3945_), .ZN(new_n4034_));
  NOR2_X1    g01599(.A1(new_n4034_), .A2(new_n3320_), .ZN(new_n4035_));
  OAI21_X1   g01600(.A1(new_n4033_), .A2(new_n4035_), .B(pi0062), .ZN(new_n4036_));
  NAND3_X1   g01601(.A1(new_n4036_), .A2(pi0241), .A3(new_n3291_), .ZN(new_n4037_));
  NOR2_X1    g01602(.A1(new_n4032_), .A2(new_n2612_), .ZN(new_n4038_));
  NOR2_X1    g01603(.A1(new_n4034_), .A2(new_n2611_), .ZN(new_n4039_));
  OAI21_X1   g01604(.A1(new_n4038_), .A2(new_n4039_), .B(pi0055), .ZN(new_n4040_));
  NOR2_X1    g01605(.A1(new_n3973_), .A2(new_n3339_), .ZN(new_n4041_));
  OAI21_X1   g01606(.A1(new_n4034_), .A2(new_n2628_), .B(new_n4041_), .ZN(new_n4042_));
  INV_X1     g01607(.I(new_n4042_), .ZN(new_n4043_));
  AOI21_X1   g01608(.A1(new_n4043_), .A2(new_n2563_), .B(pi0055), .ZN(new_n4044_));
  AOI21_X1   g01609(.A1(new_n4043_), .A2(pi0038), .B(pi0100), .ZN(new_n4045_));
  INV_X1     g01610(.I(new_n4041_), .ZN(new_n4046_));
  AOI21_X1   g01611(.A1(new_n4031_), .A2(pi0299), .B(new_n4046_), .ZN(new_n4047_));
  OAI21_X1   g01612(.A1(new_n4047_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n4048_));
  NOR2_X1    g01613(.A1(new_n3657_), .A2(new_n3934_), .ZN(new_n4049_));
  NOR2_X1    g01614(.A1(new_n3731_), .A2(pi0861), .ZN(new_n4050_));
  OAI21_X1   g01615(.A1(new_n4049_), .A2(new_n4050_), .B(pi0171), .ZN(new_n4051_));
  OAI21_X1   g01616(.A1(new_n3404_), .A2(pi0861), .B(new_n3932_), .ZN(new_n4052_));
  AOI21_X1   g01617(.A1(new_n4051_), .A2(new_n4052_), .B(pi0228), .ZN(new_n4053_));
  NOR3_X1    g01618(.A1(new_n4053_), .A2(new_n3388_), .A3(new_n3950_), .ZN(new_n4054_));
  OAI21_X1   g01619(.A1(new_n4054_), .A2(new_n3931_), .B(new_n3928_), .ZN(new_n4055_));
  OAI21_X1   g01620(.A1(new_n4055_), .A2(pi0215), .B(new_n3949_), .ZN(new_n4056_));
  AOI21_X1   g01621(.A1(new_n4056_), .A2(pi0299), .B(new_n3994_), .ZN(new_n4057_));
  OAI21_X1   g01622(.A1(new_n4057_), .A2(new_n4048_), .B(new_n4045_), .ZN(new_n4058_));
  AOI21_X1   g01623(.A1(new_n4043_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n4059_));
  AND3_X2    g01624(.A1(new_n4008_), .A2(new_n3500_), .A3(new_n3938_), .Z(new_n4060_));
  OAI21_X1   g01625(.A1(new_n4060_), .A2(new_n3931_), .B(new_n2436_), .ZN(new_n4061_));
  OAI21_X1   g01626(.A1(new_n4061_), .A2(new_n3929_), .B(new_n4004_), .ZN(new_n4062_));
  NAND3_X1   g01627(.A1(new_n4062_), .A2(new_n2572_), .A3(new_n4041_), .ZN(new_n4063_));
  NAND2_X1   g01628(.A1(new_n4063_), .A2(new_n4059_), .ZN(new_n4064_));
  NAND3_X1   g01629(.A1(new_n4058_), .A2(new_n3458_), .A3(new_n4064_), .ZN(new_n4065_));
  NOR2_X1    g01630(.A1(new_n4047_), .A2(new_n3273_), .ZN(new_n4066_));
  AOI21_X1   g01631(.A1(new_n3273_), .A2(new_n4042_), .B(new_n4066_), .ZN(new_n4067_));
  NAND2_X1   g01632(.A1(new_n4067_), .A2(pi0087), .ZN(new_n4068_));
  AOI21_X1   g01633(.A1(new_n4065_), .A2(new_n4068_), .B(pi0075), .ZN(new_n4069_));
  OAI21_X1   g01634(.A1(new_n4042_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4070_));
  NOR2_X1    g01635(.A1(new_n4067_), .A2(new_n2565_), .ZN(new_n4071_));
  AOI21_X1   g01636(.A1(new_n2565_), .A2(new_n4042_), .B(new_n4071_), .ZN(new_n4072_));
  OAI22_X1   g01637(.A1(new_n4069_), .A2(new_n4070_), .B1(new_n3444_), .B2(new_n4072_), .ZN(new_n4073_));
  OAI21_X1   g01638(.A1(new_n4073_), .A2(new_n2563_), .B(new_n4044_), .ZN(new_n4074_));
  NAND3_X1   g01639(.A1(new_n4074_), .A2(new_n3284_), .A3(new_n4040_), .ZN(new_n4075_));
  NAND2_X1   g01640(.A1(new_n4034_), .A2(new_n2577_), .ZN(new_n4076_));
  OAI21_X1   g01641(.A1(new_n4031_), .A2(new_n2577_), .B(new_n4076_), .ZN(new_n4077_));
  AOI21_X1   g01642(.A1(new_n4077_), .A2(pi0056), .B(pi0062), .ZN(new_n4078_));
  AOI21_X1   g01643(.A1(new_n4075_), .A2(new_n4078_), .B(new_n4037_), .ZN(new_n4079_));
  NOR3_X1    g01644(.A1(new_n4028_), .A2(new_n4079_), .A3(new_n3947_), .ZN(po0158));
  INV_X1     g01645(.I(pi0921), .ZN(new_n4081_));
  NOR2_X1    g01646(.A1(new_n2447_), .A2(new_n4081_), .ZN(new_n4082_));
  INV_X1     g01647(.I(pi1140), .ZN(new_n4083_));
  NOR2_X1    g01648(.A1(new_n2444_), .A2(new_n4083_), .ZN(new_n4084_));
  OAI21_X1   g01649(.A1(new_n4082_), .A2(new_n4084_), .B(pi0221), .ZN(new_n4085_));
  INV_X1     g01650(.I(new_n4085_), .ZN(new_n4086_));
  AOI21_X1   g01651(.A1(pi0216), .A2(pi0282), .B(pi0221), .ZN(new_n4087_));
  INV_X1     g01652(.I(new_n4087_), .ZN(new_n4088_));
  INV_X1     g01653(.I(pi0170), .ZN(new_n4089_));
  NAND2_X1   g01654(.A1(new_n2457_), .A2(new_n4089_), .ZN(new_n4090_));
  INV_X1     g01655(.I(pi0869), .ZN(new_n4091_));
  NOR2_X1    g01656(.A1(new_n2463_), .A2(new_n4091_), .ZN(new_n4092_));
  NAND2_X1   g01657(.A1(new_n4092_), .A2(pi0105), .ZN(new_n4093_));
  AOI21_X1   g01658(.A1(new_n4093_), .A2(new_n4090_), .B(new_n2458_), .ZN(new_n4094_));
  NOR2_X1    g01659(.A1(new_n4094_), .A2(pi0216), .ZN(new_n4095_));
  NAND2_X1   g01660(.A1(new_n4089_), .A2(new_n2458_), .ZN(new_n4096_));
  AOI21_X1   g01661(.A1(new_n4095_), .A2(new_n4096_), .B(new_n4088_), .ZN(new_n4097_));
  NOR3_X1    g01662(.A1(new_n4097_), .A2(pi0215), .A3(new_n4086_), .ZN(new_n4098_));
  NOR2_X1    g01663(.A1(new_n2436_), .A2(pi1140), .ZN(new_n4099_));
  NOR2_X1    g01664(.A1(new_n4098_), .A2(new_n4099_), .ZN(new_n4100_));
  INV_X1     g01665(.I(new_n4100_), .ZN(new_n4101_));
  AOI21_X1   g01666(.A1(pi0216), .A2(pi0282), .B(new_n3502_), .ZN(new_n4102_));
  NAND2_X1   g01667(.A1(new_n4102_), .A2(pi0248), .ZN(new_n4103_));
  AND3_X2    g01668(.A1(new_n4101_), .A2(new_n3425_), .A3(new_n4103_), .Z(new_n4104_));
  INV_X1     g01669(.I(pi0248), .ZN(new_n4105_));
  INV_X1     g01670(.I(new_n4099_), .ZN(new_n4106_));
  INV_X1     g01671(.I(new_n4095_), .ZN(new_n4107_));
  NAND2_X1   g01672(.A1(new_n2530_), .A2(new_n4089_), .ZN(new_n4108_));
  OAI21_X1   g01673(.A1(new_n4091_), .A2(new_n2530_), .B(new_n4108_), .ZN(new_n4109_));
  AOI21_X1   g01674(.A1(new_n4109_), .A2(new_n2458_), .B(new_n4107_), .ZN(new_n4110_));
  OAI21_X1   g01675(.A1(new_n4110_), .A2(new_n4088_), .B(new_n4085_), .ZN(new_n4111_));
  OAI21_X1   g01676(.A1(new_n4111_), .A2(pi0215), .B(new_n4106_), .ZN(new_n4112_));
  NOR2_X1    g01677(.A1(new_n4112_), .A2(new_n3472_), .ZN(new_n4113_));
  NOR2_X1    g01678(.A1(new_n4101_), .A2(new_n3320_), .ZN(new_n4114_));
  OAI21_X1   g01679(.A1(new_n4113_), .A2(new_n4114_), .B(pi0062), .ZN(new_n4115_));
  NAND3_X1   g01680(.A1(new_n4115_), .A2(new_n4105_), .A3(new_n3291_), .ZN(new_n4116_));
  NOR2_X1    g01681(.A1(new_n4112_), .A2(new_n2612_), .ZN(new_n4117_));
  NOR2_X1    g01682(.A1(new_n4101_), .A2(new_n2611_), .ZN(new_n4118_));
  OAI21_X1   g01683(.A1(new_n4117_), .A2(new_n4118_), .B(pi0055), .ZN(new_n4119_));
  NOR2_X1    g01684(.A1(new_n2635_), .A2(new_n4081_), .ZN(new_n4120_));
  NOR2_X1    g01685(.A1(new_n2634_), .A2(new_n4083_), .ZN(new_n4121_));
  OAI21_X1   g01686(.A1(new_n4120_), .A2(new_n4121_), .B(pi0222), .ZN(new_n4122_));
  INV_X1     g01687(.I(new_n4122_), .ZN(new_n4123_));
  AOI21_X1   g01688(.A1(pi0224), .A2(pi0282), .B(pi0222), .ZN(new_n4124_));
  INV_X1     g01689(.I(new_n4124_), .ZN(new_n4125_));
  NOR2_X1    g01690(.A1(new_n4092_), .A2(pi0224), .ZN(new_n4126_));
  NOR2_X1    g01691(.A1(new_n4126_), .A2(new_n4125_), .ZN(new_n4127_));
  OAI21_X1   g01692(.A1(new_n4123_), .A2(new_n4127_), .B(new_n2668_), .ZN(new_n4128_));
  NAND2_X1   g01693(.A1(pi0223), .A2(pi1140), .ZN(new_n4129_));
  AOI21_X1   g01694(.A1(new_n4128_), .A2(new_n4129_), .B(pi0299), .ZN(new_n4130_));
  AOI21_X1   g01695(.A1(new_n4100_), .A2(pi0299), .B(new_n4130_), .ZN(new_n4131_));
  AOI21_X1   g01696(.A1(new_n4131_), .A2(new_n2563_), .B(pi0055), .ZN(new_n4132_));
  NAND2_X1   g01697(.A1(new_n3387_), .A2(pi0869), .ZN(new_n4133_));
  NAND3_X1   g01698(.A1(new_n3657_), .A2(new_n4089_), .A3(new_n4133_), .ZN(new_n4134_));
  NOR2_X1    g01699(.A1(new_n3387_), .A2(pi0170), .ZN(new_n4135_));
  NOR2_X1    g01700(.A1(new_n3404_), .A2(new_n4089_), .ZN(new_n4136_));
  OAI21_X1   g01701(.A1(new_n4136_), .A2(new_n4135_), .B(pi0869), .ZN(new_n4137_));
  AOI21_X1   g01702(.A1(new_n4137_), .A2(new_n4134_), .B(pi0228), .ZN(new_n4138_));
  NAND2_X1   g01703(.A1(new_n3729_), .A2(new_n4094_), .ZN(new_n4139_));
  NAND2_X1   g01704(.A1(new_n4139_), .A2(new_n2614_), .ZN(new_n4140_));
  OAI21_X1   g01705(.A1(new_n4138_), .A2(new_n4140_), .B(new_n4087_), .ZN(new_n4141_));
  NAND3_X1   g01706(.A1(new_n4141_), .A2(new_n2436_), .A3(new_n4085_), .ZN(new_n4142_));
  AOI21_X1   g01707(.A1(new_n4142_), .A2(new_n4106_), .B(new_n2628_), .ZN(new_n4143_));
  NAND2_X1   g01708(.A1(new_n4129_), .A2(new_n2628_), .ZN(new_n4144_));
  OAI21_X1   g01709(.A1(new_n3392_), .A2(new_n4091_), .B(new_n2631_), .ZN(new_n4145_));
  AOI21_X1   g01710(.A1(new_n4145_), .A2(new_n4124_), .B(new_n4123_), .ZN(new_n4146_));
  INV_X1     g01711(.I(new_n4146_), .ZN(new_n4147_));
  INV_X1     g01712(.I(new_n4144_), .ZN(new_n4148_));
  AOI21_X1   g01713(.A1(new_n3392_), .A2(new_n4124_), .B(new_n4147_), .ZN(new_n4149_));
  OAI21_X1   g01714(.A1(new_n4149_), .A2(pi0223), .B(new_n4148_), .ZN(new_n4150_));
  NAND2_X1   g01715(.A1(new_n4150_), .A2(new_n2627_), .ZN(new_n4151_));
  INV_X1     g01716(.I(new_n4151_), .ZN(new_n4152_));
  OAI21_X1   g01717(.A1(new_n4144_), .A2(new_n4147_), .B(new_n4152_), .ZN(new_n4153_));
  INV_X1     g01718(.I(new_n4112_), .ZN(new_n4154_));
  AOI21_X1   g01719(.A1(new_n4154_), .A2(pi0299), .B(new_n4130_), .ZN(new_n4155_));
  OAI22_X1   g01720(.A1(new_n4143_), .A2(new_n4153_), .B1(new_n2627_), .B2(new_n4155_), .ZN(new_n4156_));
  AOI21_X1   g01721(.A1(new_n4131_), .A2(pi0038), .B(pi0100), .ZN(new_n4157_));
  OAI21_X1   g01722(.A1(new_n4156_), .A2(pi0038), .B(new_n4157_), .ZN(new_n4158_));
  AOI21_X1   g01723(.A1(new_n4131_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n4159_));
  INV_X1     g01724(.I(new_n4130_), .ZN(new_n4160_));
  NOR2_X1    g01725(.A1(new_n4099_), .A2(new_n2628_), .ZN(new_n4161_));
  INV_X1     g01726(.I(new_n4161_), .ZN(new_n4162_));
  NOR2_X1    g01727(.A1(new_n3371_), .A2(pi0170), .ZN(new_n4163_));
  NOR2_X1    g01728(.A1(new_n3544_), .A2(new_n4091_), .ZN(new_n4164_));
  OAI21_X1   g01729(.A1(new_n4164_), .A2(new_n4163_), .B(new_n2458_), .ZN(new_n4165_));
  AOI21_X1   g01730(.A1(new_n4165_), .A2(new_n4095_), .B(new_n4088_), .ZN(new_n4166_));
  NOR3_X1    g01731(.A1(new_n4166_), .A2(pi0215), .A3(new_n4086_), .ZN(new_n4167_));
  OAI21_X1   g01732(.A1(new_n4167_), .A2(new_n4162_), .B(new_n4160_), .ZN(new_n4168_));
  OAI21_X1   g01733(.A1(new_n4168_), .A2(new_n2573_), .B(new_n4159_), .ZN(new_n4169_));
  NAND3_X1   g01734(.A1(new_n4158_), .A2(new_n3458_), .A3(new_n4169_), .ZN(new_n4170_));
  INV_X1     g01735(.I(new_n4131_), .ZN(new_n4171_));
  NOR2_X1    g01736(.A1(new_n4155_), .A2(new_n3273_), .ZN(new_n4172_));
  AOI21_X1   g01737(.A1(new_n3273_), .A2(new_n4171_), .B(new_n4172_), .ZN(new_n4173_));
  NAND2_X1   g01738(.A1(new_n4173_), .A2(pi0087), .ZN(new_n4174_));
  AOI21_X1   g01739(.A1(new_n4170_), .A2(new_n4174_), .B(pi0075), .ZN(new_n4175_));
  OAI21_X1   g01740(.A1(new_n4171_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4176_));
  NOR2_X1    g01741(.A1(new_n4173_), .A2(new_n2565_), .ZN(new_n4177_));
  AOI21_X1   g01742(.A1(new_n2565_), .A2(new_n4171_), .B(new_n4177_), .ZN(new_n4178_));
  OAI22_X1   g01743(.A1(new_n4175_), .A2(new_n4176_), .B1(new_n3444_), .B2(new_n4178_), .ZN(new_n4179_));
  OAI21_X1   g01744(.A1(new_n4179_), .A2(new_n2563_), .B(new_n4132_), .ZN(new_n4180_));
  NAND3_X1   g01745(.A1(new_n4180_), .A2(new_n3284_), .A3(new_n4119_), .ZN(new_n4181_));
  NAND2_X1   g01746(.A1(new_n4101_), .A2(new_n2577_), .ZN(new_n4182_));
  OAI21_X1   g01747(.A1(new_n4154_), .A2(new_n2577_), .B(new_n4182_), .ZN(new_n4183_));
  AOI21_X1   g01748(.A1(new_n4183_), .A2(pi0056), .B(pi0062), .ZN(new_n4184_));
  AOI21_X1   g01749(.A1(new_n4181_), .A2(new_n4184_), .B(new_n4116_), .ZN(new_n4185_));
  AOI21_X1   g01750(.A1(new_n4110_), .A2(new_n3500_), .B(new_n4088_), .ZN(new_n4186_));
  NOR3_X1    g01751(.A1(new_n4186_), .A2(pi0215), .A3(new_n4086_), .ZN(new_n4187_));
  NOR2_X1    g01752(.A1(new_n4187_), .A2(new_n4099_), .ZN(new_n4188_));
  INV_X1     g01753(.I(new_n4188_), .ZN(new_n4189_));
  NOR2_X1    g01754(.A1(new_n4189_), .A2(new_n3472_), .ZN(new_n4190_));
  NOR2_X1    g01755(.A1(new_n4100_), .A2(new_n4102_), .ZN(new_n4191_));
  NOR2_X1    g01756(.A1(new_n4191_), .A2(new_n3320_), .ZN(new_n4192_));
  OAI21_X1   g01757(.A1(new_n4190_), .A2(new_n4192_), .B(pi0062), .ZN(new_n4193_));
  NAND3_X1   g01758(.A1(new_n4193_), .A2(pi0248), .A3(new_n3291_), .ZN(new_n4194_));
  NOR2_X1    g01759(.A1(new_n4189_), .A2(new_n2612_), .ZN(new_n4195_));
  NOR2_X1    g01760(.A1(new_n4191_), .A2(new_n2611_), .ZN(new_n4196_));
  OAI21_X1   g01761(.A1(new_n4195_), .A2(new_n4196_), .B(pi0055), .ZN(new_n4197_));
  NOR2_X1    g01762(.A1(new_n4130_), .A2(new_n3339_), .ZN(new_n4198_));
  OAI21_X1   g01763(.A1(new_n4191_), .A2(new_n2628_), .B(new_n4198_), .ZN(new_n4199_));
  INV_X1     g01764(.I(new_n4199_), .ZN(new_n4200_));
  AOI21_X1   g01765(.A1(new_n4200_), .A2(new_n2563_), .B(pi0055), .ZN(new_n4201_));
  AOI21_X1   g01766(.A1(new_n4200_), .A2(pi0038), .B(pi0100), .ZN(new_n4202_));
  INV_X1     g01767(.I(new_n4198_), .ZN(new_n4203_));
  AOI21_X1   g01768(.A1(new_n4188_), .A2(pi0299), .B(new_n4203_), .ZN(new_n4204_));
  OAI21_X1   g01769(.A1(new_n4204_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n4205_));
  NOR2_X1    g01770(.A1(new_n3657_), .A2(new_n4091_), .ZN(new_n4206_));
  NOR2_X1    g01771(.A1(new_n3731_), .A2(pi0869), .ZN(new_n4207_));
  OAI21_X1   g01772(.A1(new_n4206_), .A2(new_n4207_), .B(pi0170), .ZN(new_n4208_));
  OAI21_X1   g01773(.A1(new_n3404_), .A2(pi0869), .B(new_n4089_), .ZN(new_n4209_));
  AOI21_X1   g01774(.A1(new_n4208_), .A2(new_n4209_), .B(pi0228), .ZN(new_n4210_));
  NOR3_X1    g01775(.A1(new_n4210_), .A2(new_n3388_), .A3(new_n4107_), .ZN(new_n4211_));
  OAI21_X1   g01776(.A1(new_n4211_), .A2(new_n4088_), .B(new_n4085_), .ZN(new_n4212_));
  OAI21_X1   g01777(.A1(new_n4212_), .A2(pi0215), .B(new_n4106_), .ZN(new_n4213_));
  AOI21_X1   g01778(.A1(new_n4213_), .A2(pi0299), .B(new_n4151_), .ZN(new_n4214_));
  OAI21_X1   g01779(.A1(new_n4214_), .A2(new_n4205_), .B(new_n4202_), .ZN(new_n4215_));
  AOI21_X1   g01780(.A1(new_n4200_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n4216_));
  AND3_X2    g01781(.A1(new_n4165_), .A2(new_n3500_), .A3(new_n4095_), .Z(new_n4217_));
  OAI21_X1   g01782(.A1(new_n4217_), .A2(new_n4088_), .B(new_n2436_), .ZN(new_n4218_));
  OAI21_X1   g01783(.A1(new_n4218_), .A2(new_n4086_), .B(new_n4161_), .ZN(new_n4219_));
  NAND3_X1   g01784(.A1(new_n4219_), .A2(new_n2572_), .A3(new_n4198_), .ZN(new_n4220_));
  NAND2_X1   g01785(.A1(new_n4220_), .A2(new_n4216_), .ZN(new_n4221_));
  NAND3_X1   g01786(.A1(new_n4215_), .A2(new_n3458_), .A3(new_n4221_), .ZN(new_n4222_));
  NOR2_X1    g01787(.A1(new_n4204_), .A2(new_n3273_), .ZN(new_n4223_));
  AOI21_X1   g01788(.A1(new_n3273_), .A2(new_n4199_), .B(new_n4223_), .ZN(new_n4224_));
  NAND2_X1   g01789(.A1(new_n4224_), .A2(pi0087), .ZN(new_n4225_));
  AOI21_X1   g01790(.A1(new_n4222_), .A2(new_n4225_), .B(pi0075), .ZN(new_n4226_));
  OAI21_X1   g01791(.A1(new_n4199_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4227_));
  NOR2_X1    g01792(.A1(new_n4224_), .A2(new_n2565_), .ZN(new_n4228_));
  AOI21_X1   g01793(.A1(new_n2565_), .A2(new_n4199_), .B(new_n4228_), .ZN(new_n4229_));
  OAI22_X1   g01794(.A1(new_n4226_), .A2(new_n4227_), .B1(new_n3444_), .B2(new_n4229_), .ZN(new_n4230_));
  OAI21_X1   g01795(.A1(new_n4230_), .A2(new_n2563_), .B(new_n4201_), .ZN(new_n4231_));
  NAND3_X1   g01796(.A1(new_n4231_), .A2(new_n3284_), .A3(new_n4197_), .ZN(new_n4232_));
  NAND2_X1   g01797(.A1(new_n4191_), .A2(new_n2577_), .ZN(new_n4233_));
  OAI21_X1   g01798(.A1(new_n4188_), .A2(new_n2577_), .B(new_n4233_), .ZN(new_n4234_));
  AOI21_X1   g01799(.A1(new_n4234_), .A2(pi0056), .B(pi0062), .ZN(new_n4235_));
  AOI21_X1   g01800(.A1(new_n4232_), .A2(new_n4235_), .B(new_n4194_), .ZN(new_n4236_));
  NOR3_X1    g01801(.A1(new_n4185_), .A2(new_n4236_), .A3(new_n4104_), .ZN(po0159));
  INV_X1     g01802(.I(pi1139), .ZN(new_n4238_));
  INV_X1     g01803(.I(pi0920), .ZN(new_n4239_));
  NOR2_X1    g01804(.A1(pi0833), .A2(pi1139), .ZN(new_n4240_));
  AOI21_X1   g01805(.A1(pi0833), .A2(new_n4239_), .B(new_n4240_), .ZN(new_n4241_));
  OAI21_X1   g01806(.A1(new_n4241_), .A2(pi0216), .B(pi0221), .ZN(new_n4242_));
  AOI21_X1   g01807(.A1(pi0216), .A2(new_n4238_), .B(new_n4242_), .ZN(new_n4243_));
  AOI21_X1   g01808(.A1(pi0216), .A2(pi0281), .B(pi0221), .ZN(new_n4244_));
  NOR2_X1    g01809(.A1(new_n3322_), .A2(new_n3543_), .ZN(new_n4245_));
  INV_X1     g01810(.I(new_n4245_), .ZN(new_n4246_));
  NOR2_X1    g01811(.A1(pi0216), .A2(pi0862), .ZN(new_n4247_));
  NAND2_X1   g01812(.A1(new_n4246_), .A2(new_n4247_), .ZN(new_n4248_));
  AOI21_X1   g01813(.A1(new_n4248_), .A2(new_n4244_), .B(new_n4243_), .ZN(new_n4249_));
  INV_X1     g01814(.I(new_n4249_), .ZN(new_n4250_));
  NOR2_X1    g01815(.A1(new_n2436_), .A2(new_n4238_), .ZN(new_n4251_));
  INV_X1     g01816(.I(new_n4251_), .ZN(new_n4252_));
  INV_X1     g01817(.I(new_n4242_), .ZN(new_n4253_));
  NOR2_X1    g01818(.A1(new_n4253_), .A2(pi0216), .ZN(new_n4254_));
  INV_X1     g01819(.I(new_n4254_), .ZN(new_n4255_));
  NOR2_X1    g01820(.A1(new_n4246_), .A2(new_n4255_), .ZN(new_n4256_));
  INV_X1     g01821(.I(pi0148), .ZN(new_n4257_));
  NOR2_X1    g01822(.A1(new_n4257_), .A2(pi0215), .ZN(new_n4258_));
  NAND2_X1   g01823(.A1(new_n4250_), .A2(new_n4258_), .ZN(new_n4259_));
  OAI21_X1   g01824(.A1(new_n4259_), .A2(new_n4256_), .B(new_n4252_), .ZN(new_n4260_));
  NOR2_X1    g01825(.A1(new_n4255_), .A2(new_n4257_), .ZN(new_n4261_));
  AOI21_X1   g01826(.A1(new_n4261_), .A2(new_n2460_), .B(pi0215), .ZN(new_n4262_));
  AOI21_X1   g01827(.A1(new_n4250_), .A2(new_n4262_), .B(new_n4260_), .ZN(new_n4263_));
  INV_X1     g01828(.I(new_n4263_), .ZN(new_n4264_));
  NAND2_X1   g01829(.A1(new_n4264_), .A2(new_n2611_), .ZN(new_n4265_));
  INV_X1     g01830(.I(new_n4243_), .ZN(new_n4266_));
  INV_X1     g01831(.I(new_n4244_), .ZN(new_n4267_));
  NOR4_X1    g01832(.A1(new_n2460_), .A2(pi0216), .A3(pi0862), .A4(new_n2463_), .ZN(new_n4268_));
  OAI21_X1   g01833(.A1(new_n4267_), .A2(new_n4268_), .B(new_n4266_), .ZN(new_n4269_));
  NAND2_X1   g01834(.A1(new_n4262_), .A2(new_n4269_), .ZN(new_n4270_));
  NAND2_X1   g01835(.A1(new_n4270_), .A2(new_n4252_), .ZN(new_n4271_));
  NAND2_X1   g01836(.A1(new_n4271_), .A2(new_n2612_), .ZN(new_n4272_));
  AOI21_X1   g01837(.A1(new_n4265_), .A2(new_n4272_), .B(new_n2602_), .ZN(new_n4273_));
  NOR2_X1    g01838(.A1(new_n2668_), .A2(new_n4238_), .ZN(new_n4274_));
  NOR2_X1    g01839(.A1(new_n2635_), .A2(new_n4239_), .ZN(new_n4275_));
  NOR2_X1    g01840(.A1(new_n2634_), .A2(new_n4238_), .ZN(new_n4276_));
  OAI21_X1   g01841(.A1(new_n4275_), .A2(new_n4276_), .B(pi0222), .ZN(new_n4277_));
  INV_X1     g01842(.I(pi0281), .ZN(new_n4278_));
  NOR2_X1    g01843(.A1(new_n2631_), .A2(new_n4278_), .ZN(new_n4279_));
  OAI21_X1   g01844(.A1(pi0222), .A2(new_n4279_), .B(new_n4277_), .ZN(new_n4280_));
  AOI21_X1   g01845(.A1(new_n4280_), .A2(new_n2668_), .B(new_n4274_), .ZN(new_n4281_));
  NOR2_X1    g01846(.A1(new_n4281_), .A2(pi0299), .ZN(new_n4282_));
  INV_X1     g01847(.I(pi0862), .ZN(new_n4283_));
  INV_X1     g01848(.I(new_n4277_), .ZN(new_n4284_));
  NOR3_X1    g01849(.A1(new_n4284_), .A2(pi0224), .A3(new_n4274_), .ZN(new_n4285_));
  NAND2_X1   g01850(.A1(new_n4285_), .A2(new_n4283_), .ZN(new_n4286_));
  AOI21_X1   g01851(.A1(new_n4282_), .A2(new_n4286_), .B(new_n3339_), .ZN(new_n4287_));
  INV_X1     g01852(.I(new_n4287_), .ZN(new_n4288_));
  AOI21_X1   g01853(.A1(new_n4271_), .A2(pi0299), .B(new_n4288_), .ZN(new_n4289_));
  INV_X1     g01854(.I(new_n4289_), .ZN(new_n4290_));
  OAI21_X1   g01855(.A1(new_n4290_), .A2(new_n2562_), .B(new_n2602_), .ZN(new_n4291_));
  AOI21_X1   g01856(.A1(new_n4264_), .A2(pi0299), .B(new_n4288_), .ZN(new_n4292_));
  NAND2_X1   g01857(.A1(new_n4292_), .A2(pi0039), .ZN(new_n4293_));
  OAI21_X1   g01858(.A1(new_n3392_), .A2(new_n4286_), .B(new_n4282_), .ZN(new_n4294_));
  INV_X1     g01859(.I(new_n4258_), .ZN(new_n4295_));
  NOR2_X1    g01860(.A1(new_n3390_), .A2(pi0862), .ZN(new_n4296_));
  NOR2_X1    g01861(.A1(new_n2458_), .A2(pi0105), .ZN(new_n4297_));
  INV_X1     g01862(.I(new_n4297_), .ZN(new_n4298_));
  OAI21_X1   g01863(.A1(new_n3451_), .A2(pi0228), .B(new_n4298_), .ZN(new_n4299_));
  AOI21_X1   g01864(.A1(new_n4299_), .A2(pi0862), .B(new_n4296_), .ZN(new_n4300_));
  OAI21_X1   g01865(.A1(new_n4300_), .A2(pi0216), .B(new_n4244_), .ZN(new_n4301_));
  AOI21_X1   g01866(.A1(new_n4301_), .A2(new_n4266_), .B(new_n4295_), .ZN(new_n4302_));
  NOR2_X1    g01867(.A1(pi0148), .A2(pi0215), .ZN(new_n4303_));
  INV_X1     g01868(.I(new_n4303_), .ZN(new_n4304_));
  NAND2_X1   g01869(.A1(new_n3405_), .A2(new_n4247_), .ZN(new_n4305_));
  AOI21_X1   g01870(.A1(new_n4305_), .A2(new_n4244_), .B(new_n4243_), .ZN(new_n4306_));
  OAI21_X1   g01871(.A1(new_n4306_), .A2(new_n4304_), .B(new_n4252_), .ZN(new_n4307_));
  OAI21_X1   g01872(.A1(new_n4307_), .A2(new_n4302_), .B(pi0299), .ZN(new_n4308_));
  NAND3_X1   g01873(.A1(new_n4308_), .A2(new_n2627_), .A3(new_n4294_), .ZN(new_n4309_));
  AOI21_X1   g01874(.A1(new_n4309_), .A2(new_n4293_), .B(pi0038), .ZN(new_n4310_));
  OAI21_X1   g01875(.A1(new_n4290_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n4311_));
  OAI21_X1   g01876(.A1(new_n4290_), .A2(new_n2572_), .B(pi0100), .ZN(new_n4312_));
  NOR4_X1    g01877(.A1(new_n3545_), .A2(pi0216), .A3(new_n2459_), .A4(new_n4243_), .ZN(new_n4313_));
  OAI21_X1   g01878(.A1(new_n4313_), .A2(new_n4259_), .B(new_n4252_), .ZN(new_n4314_));
  AOI21_X1   g01879(.A1(new_n3546_), .A2(new_n4244_), .B(new_n4250_), .ZN(new_n4315_));
  NOR2_X1    g01880(.A1(new_n4315_), .A2(new_n4304_), .ZN(new_n4316_));
  OAI21_X1   g01881(.A1(new_n4316_), .A2(new_n4314_), .B(pi0299), .ZN(new_n4317_));
  AND3_X2    g01882(.A1(new_n4317_), .A2(new_n2572_), .A3(new_n4287_), .Z(new_n4318_));
  OAI22_X1   g01883(.A1(new_n4310_), .A2(new_n4311_), .B1(new_n4312_), .B2(new_n4318_), .ZN(new_n4319_));
  NOR2_X1    g01884(.A1(new_n4292_), .A2(new_n3273_), .ZN(new_n4320_));
  AOI21_X1   g01885(.A1(new_n3273_), .A2(new_n4290_), .B(new_n4320_), .ZN(new_n4321_));
  NAND2_X1   g01886(.A1(new_n4321_), .A2(pi0087), .ZN(new_n4322_));
  OAI21_X1   g01887(.A1(new_n4319_), .A2(pi0087), .B(new_n4322_), .ZN(new_n4323_));
  OAI21_X1   g01888(.A1(new_n4290_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4324_));
  AOI21_X1   g01889(.A1(new_n4323_), .A2(new_n3465_), .B(new_n4324_), .ZN(new_n4325_));
  NAND2_X1   g01890(.A1(new_n4290_), .A2(new_n2565_), .ZN(new_n4326_));
  OR2_X2     g01891(.A1(new_n4321_), .A2(new_n2565_), .Z(new_n4327_));
  AOI21_X1   g01892(.A1(new_n4327_), .A2(new_n4326_), .B(new_n3444_), .ZN(new_n4328_));
  NOR3_X1    g01893(.A1(new_n4325_), .A2(new_n2563_), .A3(new_n4328_), .ZN(new_n4329_));
  OAI21_X1   g01894(.A1(new_n4329_), .A2(new_n4291_), .B(new_n3284_), .ZN(new_n4330_));
  NOR2_X1    g01895(.A1(new_n4271_), .A2(new_n2576_), .ZN(new_n4331_));
  AOI21_X1   g01896(.A1(new_n4263_), .A2(new_n2576_), .B(new_n4331_), .ZN(new_n4332_));
  OAI22_X1   g01897(.A1(new_n4330_), .A2(new_n4273_), .B1(new_n3284_), .B2(new_n4332_), .ZN(new_n4333_));
  NOR2_X1    g01898(.A1(new_n4263_), .A2(new_n3472_), .ZN(new_n4334_));
  INV_X1     g01899(.I(new_n4271_), .ZN(new_n4335_));
  NOR2_X1    g01900(.A1(new_n4335_), .A2(new_n3320_), .ZN(new_n4336_));
  OAI21_X1   g01901(.A1(new_n4334_), .A2(new_n4336_), .B(pi0062), .ZN(new_n4337_));
  OAI21_X1   g01902(.A1(new_n4333_), .A2(pi0062), .B(new_n4337_), .ZN(new_n4338_));
  INV_X1     g01903(.I(pi0247), .ZN(new_n4339_));
  AOI21_X1   g01904(.A1(new_n4335_), .A2(new_n3425_), .B(new_n4339_), .ZN(new_n4340_));
  OAI21_X1   g01905(.A1(new_n4338_), .A2(new_n3425_), .B(new_n4340_), .ZN(new_n4341_));
  OAI21_X1   g01906(.A1(new_n3302_), .A2(new_n4283_), .B(new_n2614_), .ZN(new_n4342_));
  AOI21_X1   g01907(.A1(new_n3487_), .A2(new_n2460_), .B(new_n4342_), .ZN(new_n4343_));
  OAI21_X1   g01908(.A1(new_n4343_), .A2(new_n4267_), .B(new_n4266_), .ZN(new_n4344_));
  NAND2_X1   g01909(.A1(new_n4344_), .A2(new_n4303_), .ZN(new_n4345_));
  INV_X1     g01910(.I(new_n4345_), .ZN(new_n4346_));
  NOR2_X1    g01911(.A1(new_n4260_), .A2(new_n4346_), .ZN(new_n4347_));
  INV_X1     g01912(.I(new_n4347_), .ZN(new_n4348_));
  NAND2_X1   g01913(.A1(new_n4348_), .A2(new_n2611_), .ZN(new_n4349_));
  NOR2_X1    g01914(.A1(new_n4335_), .A2(new_n3307_), .ZN(new_n4350_));
  NAND2_X1   g01915(.A1(new_n4350_), .A2(new_n2612_), .ZN(new_n4351_));
  AOI21_X1   g01916(.A1(new_n4349_), .A2(new_n4351_), .B(new_n2602_), .ZN(new_n4352_));
  OAI21_X1   g01917(.A1(new_n4283_), .A2(new_n2463_), .B(new_n4285_), .ZN(new_n4353_));
  AND2_X2    g01918(.A1(new_n4282_), .A2(new_n4353_), .Z(new_n4354_));
  AOI21_X1   g01919(.A1(new_n4350_), .A2(pi0299), .B(new_n4354_), .ZN(new_n4355_));
  INV_X1     g01920(.I(new_n4355_), .ZN(new_n4356_));
  OAI21_X1   g01921(.A1(new_n4356_), .A2(new_n2562_), .B(new_n2602_), .ZN(new_n4357_));
  NOR2_X1    g01922(.A1(new_n4299_), .A2(pi0862), .ZN(new_n4358_));
  AOI21_X1   g01923(.A1(pi0862), .A2(new_n3390_), .B(new_n4358_), .ZN(new_n4359_));
  OAI21_X1   g01924(.A1(new_n4359_), .A2(pi0216), .B(new_n4244_), .ZN(new_n4360_));
  AOI21_X1   g01925(.A1(new_n4360_), .A2(new_n4266_), .B(new_n4304_), .ZN(new_n4361_));
  OAI21_X1   g01926(.A1(new_n3405_), .A2(new_n4255_), .B(new_n4258_), .ZN(new_n4362_));
  NOR2_X1    g01927(.A1(new_n4306_), .A2(new_n4362_), .ZN(new_n4363_));
  NOR4_X1    g01928(.A1(new_n4361_), .A2(new_n4363_), .A3(new_n2628_), .A4(new_n4251_), .ZN(new_n4364_));
  INV_X1     g01929(.I(new_n4281_), .ZN(new_n4365_));
  OAI21_X1   g01930(.A1(new_n3392_), .A2(new_n4283_), .B(new_n4285_), .ZN(new_n4366_));
  AOI21_X1   g01931(.A1(new_n4366_), .A2(new_n4365_), .B(pi0299), .ZN(new_n4367_));
  NOR3_X1    g01932(.A1(new_n4364_), .A2(pi0039), .A3(new_n4367_), .ZN(new_n4368_));
  AOI21_X1   g01933(.A1(new_n4348_), .A2(pi0299), .B(new_n4354_), .ZN(new_n4369_));
  NOR2_X1    g01934(.A1(new_n4369_), .A2(new_n2627_), .ZN(new_n4370_));
  NOR3_X1    g01935(.A1(new_n4368_), .A2(pi0038), .A3(new_n4370_), .ZN(new_n4371_));
  OAI21_X1   g01936(.A1(new_n4356_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n4372_));
  AOI21_X1   g01937(.A1(new_n4355_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n4373_));
  INV_X1     g01938(.I(new_n4315_), .ZN(new_n4374_));
  AOI21_X1   g01939(.A1(new_n3546_), .A2(new_n4254_), .B(new_n4295_), .ZN(new_n4375_));
  NOR3_X1    g01940(.A1(new_n3545_), .A2(new_n2459_), .A3(new_n4267_), .ZN(new_n4376_));
  OAI21_X1   g01941(.A1(new_n4376_), .A2(new_n4344_), .B(new_n4303_), .ZN(new_n4377_));
  NAND2_X1   g01942(.A1(new_n4377_), .A2(new_n4252_), .ZN(new_n4378_));
  AOI21_X1   g01943(.A1(new_n4375_), .A2(new_n4374_), .B(new_n4378_), .ZN(new_n4379_));
  OAI21_X1   g01944(.A1(new_n4379_), .A2(new_n2628_), .B(new_n2572_), .ZN(new_n4380_));
  OAI21_X1   g01945(.A1(new_n4380_), .A2(new_n4354_), .B(new_n4373_), .ZN(new_n4381_));
  OAI21_X1   g01946(.A1(new_n4371_), .A2(new_n4372_), .B(new_n4381_), .ZN(new_n4382_));
  NOR2_X1    g01947(.A1(new_n4369_), .A2(new_n3273_), .ZN(new_n4383_));
  AOI21_X1   g01948(.A1(new_n3273_), .A2(new_n4356_), .B(new_n4383_), .ZN(new_n4384_));
  NAND2_X1   g01949(.A1(new_n4384_), .A2(pi0087), .ZN(new_n4385_));
  OAI21_X1   g01950(.A1(new_n4382_), .A2(pi0087), .B(new_n4385_), .ZN(new_n4386_));
  OAI21_X1   g01951(.A1(new_n4356_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4387_));
  AOI21_X1   g01952(.A1(new_n4386_), .A2(new_n3465_), .B(new_n4387_), .ZN(new_n4388_));
  NAND2_X1   g01953(.A1(new_n4356_), .A2(new_n2565_), .ZN(new_n4389_));
  OR2_X2     g01954(.A1(new_n4384_), .A2(new_n2565_), .Z(new_n4390_));
  AOI21_X1   g01955(.A1(new_n4390_), .A2(new_n4389_), .B(new_n3444_), .ZN(new_n4391_));
  NOR3_X1    g01956(.A1(new_n4388_), .A2(new_n2563_), .A3(new_n4391_), .ZN(new_n4392_));
  OAI21_X1   g01957(.A1(new_n4392_), .A2(new_n4357_), .B(new_n3284_), .ZN(new_n4393_));
  NOR2_X1    g01958(.A1(new_n4350_), .A2(new_n2576_), .ZN(new_n4394_));
  NOR2_X1    g01959(.A1(new_n4348_), .A2(new_n2577_), .ZN(new_n4395_));
  OAI21_X1   g01960(.A1(new_n4395_), .A2(new_n4394_), .B(pi0056), .ZN(new_n4396_));
  OAI21_X1   g01961(.A1(new_n4393_), .A2(new_n4352_), .B(new_n4396_), .ZN(new_n4397_));
  NOR2_X1    g01962(.A1(new_n4347_), .A2(new_n3472_), .ZN(new_n4398_));
  INV_X1     g01963(.I(new_n4350_), .ZN(new_n4399_));
  NOR2_X1    g01964(.A1(new_n4399_), .A2(new_n3320_), .ZN(new_n4400_));
  OAI21_X1   g01965(.A1(new_n4398_), .A2(new_n4400_), .B(pi0062), .ZN(new_n4401_));
  OAI21_X1   g01966(.A1(new_n4397_), .A2(pi0062), .B(new_n4401_), .ZN(new_n4402_));
  AOI21_X1   g01967(.A1(new_n4399_), .A2(new_n3425_), .B(pi0247), .ZN(new_n4403_));
  OAI21_X1   g01968(.A1(new_n4402_), .A2(new_n3425_), .B(new_n4403_), .ZN(new_n4404_));
  NAND2_X1   g01969(.A1(new_n4404_), .A2(new_n4341_), .ZN(po0160));
  INV_X1     g01970(.I(pi0940), .ZN(new_n4406_));
  NOR2_X1    g01971(.A1(new_n2447_), .A2(new_n4406_), .ZN(new_n4407_));
  INV_X1     g01972(.I(pi1138), .ZN(new_n4408_));
  NOR2_X1    g01973(.A1(new_n2444_), .A2(new_n4408_), .ZN(new_n4409_));
  OAI21_X1   g01974(.A1(new_n4407_), .A2(new_n4409_), .B(pi0221), .ZN(new_n4410_));
  INV_X1     g01975(.I(new_n4410_), .ZN(new_n4411_));
  AOI21_X1   g01976(.A1(pi0216), .A2(pi0269), .B(pi0221), .ZN(new_n4412_));
  INV_X1     g01977(.I(new_n4412_), .ZN(new_n4413_));
  INV_X1     g01978(.I(pi0169), .ZN(new_n4414_));
  NAND2_X1   g01979(.A1(new_n2457_), .A2(new_n4414_), .ZN(new_n4415_));
  INV_X1     g01980(.I(pi0877), .ZN(new_n4416_));
  NOR2_X1    g01981(.A1(new_n2463_), .A2(new_n4416_), .ZN(new_n4417_));
  NAND2_X1   g01982(.A1(new_n4417_), .A2(pi0105), .ZN(new_n4418_));
  AOI21_X1   g01983(.A1(new_n4418_), .A2(new_n4415_), .B(new_n2458_), .ZN(new_n4419_));
  NOR2_X1    g01984(.A1(new_n4419_), .A2(pi0216), .ZN(new_n4420_));
  NAND2_X1   g01985(.A1(new_n4414_), .A2(new_n2458_), .ZN(new_n4421_));
  AOI21_X1   g01986(.A1(new_n4420_), .A2(new_n4421_), .B(new_n4413_), .ZN(new_n4422_));
  NOR3_X1    g01987(.A1(new_n4422_), .A2(pi0215), .A3(new_n4411_), .ZN(new_n4423_));
  NOR2_X1    g01988(.A1(new_n2436_), .A2(pi1138), .ZN(new_n4424_));
  NOR2_X1    g01989(.A1(new_n4423_), .A2(new_n4424_), .ZN(new_n4425_));
  INV_X1     g01990(.I(new_n4425_), .ZN(new_n4426_));
  AOI21_X1   g01991(.A1(pi0216), .A2(pi0269), .B(new_n3502_), .ZN(new_n4427_));
  NAND2_X1   g01992(.A1(new_n4427_), .A2(pi0246), .ZN(new_n4428_));
  AND3_X2    g01993(.A1(new_n4426_), .A2(new_n3425_), .A3(new_n4428_), .Z(new_n4429_));
  INV_X1     g01994(.I(pi0246), .ZN(new_n4430_));
  INV_X1     g01995(.I(new_n4424_), .ZN(new_n4431_));
  INV_X1     g01996(.I(new_n4420_), .ZN(new_n4432_));
  NAND2_X1   g01997(.A1(new_n2530_), .A2(new_n4414_), .ZN(new_n4433_));
  OAI21_X1   g01998(.A1(new_n4416_), .A2(new_n2530_), .B(new_n4433_), .ZN(new_n4434_));
  AOI21_X1   g01999(.A1(new_n4434_), .A2(new_n2458_), .B(new_n4432_), .ZN(new_n4435_));
  OAI21_X1   g02000(.A1(new_n4435_), .A2(new_n4413_), .B(new_n4410_), .ZN(new_n4436_));
  OAI21_X1   g02001(.A1(new_n4436_), .A2(pi0215), .B(new_n4431_), .ZN(new_n4437_));
  NOR2_X1    g02002(.A1(new_n4437_), .A2(new_n3472_), .ZN(new_n4438_));
  NOR2_X1    g02003(.A1(new_n4426_), .A2(new_n3320_), .ZN(new_n4439_));
  OAI21_X1   g02004(.A1(new_n4438_), .A2(new_n4439_), .B(pi0062), .ZN(new_n4440_));
  NAND3_X1   g02005(.A1(new_n4440_), .A2(new_n4430_), .A3(new_n3291_), .ZN(new_n4441_));
  NOR2_X1    g02006(.A1(new_n4437_), .A2(new_n2612_), .ZN(new_n4442_));
  NOR2_X1    g02007(.A1(new_n4426_), .A2(new_n2611_), .ZN(new_n4443_));
  OAI21_X1   g02008(.A1(new_n4442_), .A2(new_n4443_), .B(pi0055), .ZN(new_n4444_));
  NOR2_X1    g02009(.A1(new_n2635_), .A2(new_n4406_), .ZN(new_n4445_));
  NOR2_X1    g02010(.A1(new_n2634_), .A2(new_n4408_), .ZN(new_n4446_));
  OAI21_X1   g02011(.A1(new_n4445_), .A2(new_n4446_), .B(pi0222), .ZN(new_n4447_));
  INV_X1     g02012(.I(new_n4447_), .ZN(new_n4448_));
  AOI21_X1   g02013(.A1(pi0224), .A2(pi0269), .B(pi0222), .ZN(new_n4449_));
  INV_X1     g02014(.I(new_n4449_), .ZN(new_n4450_));
  NOR2_X1    g02015(.A1(new_n4417_), .A2(pi0224), .ZN(new_n4451_));
  NOR2_X1    g02016(.A1(new_n4451_), .A2(new_n4450_), .ZN(new_n4452_));
  OAI21_X1   g02017(.A1(new_n4448_), .A2(new_n4452_), .B(new_n2668_), .ZN(new_n4453_));
  NAND2_X1   g02018(.A1(pi0223), .A2(pi1138), .ZN(new_n4454_));
  AOI21_X1   g02019(.A1(new_n4453_), .A2(new_n4454_), .B(pi0299), .ZN(new_n4455_));
  AOI21_X1   g02020(.A1(new_n4425_), .A2(pi0299), .B(new_n4455_), .ZN(new_n4456_));
  AOI21_X1   g02021(.A1(new_n4456_), .A2(new_n2563_), .B(pi0055), .ZN(new_n4457_));
  NAND2_X1   g02022(.A1(new_n3387_), .A2(pi0877), .ZN(new_n4458_));
  NAND3_X1   g02023(.A1(new_n3657_), .A2(new_n4414_), .A3(new_n4458_), .ZN(new_n4459_));
  NOR2_X1    g02024(.A1(new_n3387_), .A2(pi0169), .ZN(new_n4460_));
  NOR2_X1    g02025(.A1(new_n3404_), .A2(new_n4414_), .ZN(new_n4461_));
  OAI21_X1   g02026(.A1(new_n4461_), .A2(new_n4460_), .B(pi0877), .ZN(new_n4462_));
  AOI21_X1   g02027(.A1(new_n4462_), .A2(new_n4459_), .B(pi0228), .ZN(new_n4463_));
  NAND2_X1   g02028(.A1(new_n3729_), .A2(new_n4419_), .ZN(new_n4464_));
  NAND2_X1   g02029(.A1(new_n4464_), .A2(new_n2614_), .ZN(new_n4465_));
  OAI21_X1   g02030(.A1(new_n4463_), .A2(new_n4465_), .B(new_n4412_), .ZN(new_n4466_));
  NAND3_X1   g02031(.A1(new_n4466_), .A2(new_n2436_), .A3(new_n4410_), .ZN(new_n4467_));
  AOI21_X1   g02032(.A1(new_n4467_), .A2(new_n4431_), .B(new_n2628_), .ZN(new_n4468_));
  NAND2_X1   g02033(.A1(new_n4454_), .A2(new_n2628_), .ZN(new_n4469_));
  OAI21_X1   g02034(.A1(new_n3392_), .A2(new_n4416_), .B(new_n2631_), .ZN(new_n4470_));
  AOI21_X1   g02035(.A1(new_n4470_), .A2(new_n4449_), .B(new_n4448_), .ZN(new_n4471_));
  INV_X1     g02036(.I(new_n4471_), .ZN(new_n4472_));
  INV_X1     g02037(.I(new_n4469_), .ZN(new_n4473_));
  AOI21_X1   g02038(.A1(new_n3392_), .A2(new_n4449_), .B(new_n4472_), .ZN(new_n4474_));
  OAI21_X1   g02039(.A1(new_n4474_), .A2(pi0223), .B(new_n4473_), .ZN(new_n4475_));
  NAND2_X1   g02040(.A1(new_n4475_), .A2(new_n2627_), .ZN(new_n4476_));
  INV_X1     g02041(.I(new_n4476_), .ZN(new_n4477_));
  OAI21_X1   g02042(.A1(new_n4469_), .A2(new_n4472_), .B(new_n4477_), .ZN(new_n4478_));
  INV_X1     g02043(.I(new_n4437_), .ZN(new_n4479_));
  AOI21_X1   g02044(.A1(new_n4479_), .A2(pi0299), .B(new_n4455_), .ZN(new_n4480_));
  OAI22_X1   g02045(.A1(new_n4468_), .A2(new_n4478_), .B1(new_n2627_), .B2(new_n4480_), .ZN(new_n4481_));
  AOI21_X1   g02046(.A1(new_n4456_), .A2(pi0038), .B(pi0100), .ZN(new_n4482_));
  OAI21_X1   g02047(.A1(new_n4481_), .A2(pi0038), .B(new_n4482_), .ZN(new_n4483_));
  AOI21_X1   g02048(.A1(new_n4456_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n4484_));
  INV_X1     g02049(.I(new_n4455_), .ZN(new_n4485_));
  NOR2_X1    g02050(.A1(new_n4424_), .A2(new_n2628_), .ZN(new_n4486_));
  INV_X1     g02051(.I(new_n4486_), .ZN(new_n4487_));
  NOR2_X1    g02052(.A1(new_n3371_), .A2(pi0169), .ZN(new_n4488_));
  NOR2_X1    g02053(.A1(new_n3544_), .A2(new_n4416_), .ZN(new_n4489_));
  OAI21_X1   g02054(.A1(new_n4489_), .A2(new_n4488_), .B(new_n2458_), .ZN(new_n4490_));
  AOI21_X1   g02055(.A1(new_n4490_), .A2(new_n4420_), .B(new_n4413_), .ZN(new_n4491_));
  NOR3_X1    g02056(.A1(new_n4491_), .A2(pi0215), .A3(new_n4411_), .ZN(new_n4492_));
  OAI21_X1   g02057(.A1(new_n4492_), .A2(new_n4487_), .B(new_n4485_), .ZN(new_n4493_));
  OAI21_X1   g02058(.A1(new_n4493_), .A2(new_n2573_), .B(new_n4484_), .ZN(new_n4494_));
  NAND3_X1   g02059(.A1(new_n4483_), .A2(new_n3458_), .A3(new_n4494_), .ZN(new_n4495_));
  INV_X1     g02060(.I(new_n4456_), .ZN(new_n4496_));
  NOR2_X1    g02061(.A1(new_n4480_), .A2(new_n3273_), .ZN(new_n4497_));
  AOI21_X1   g02062(.A1(new_n3273_), .A2(new_n4496_), .B(new_n4497_), .ZN(new_n4498_));
  NAND2_X1   g02063(.A1(new_n4498_), .A2(pi0087), .ZN(new_n4499_));
  AOI21_X1   g02064(.A1(new_n4495_), .A2(new_n4499_), .B(pi0075), .ZN(new_n4500_));
  OAI21_X1   g02065(.A1(new_n4496_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4501_));
  NOR2_X1    g02066(.A1(new_n4498_), .A2(new_n2565_), .ZN(new_n4502_));
  AOI21_X1   g02067(.A1(new_n2565_), .A2(new_n4496_), .B(new_n4502_), .ZN(new_n4503_));
  OAI22_X1   g02068(.A1(new_n4500_), .A2(new_n4501_), .B1(new_n3444_), .B2(new_n4503_), .ZN(new_n4504_));
  OAI21_X1   g02069(.A1(new_n4504_), .A2(new_n2563_), .B(new_n4457_), .ZN(new_n4505_));
  NAND3_X1   g02070(.A1(new_n4505_), .A2(new_n3284_), .A3(new_n4444_), .ZN(new_n4506_));
  NAND2_X1   g02071(.A1(new_n4426_), .A2(new_n2577_), .ZN(new_n4507_));
  OAI21_X1   g02072(.A1(new_n4479_), .A2(new_n2577_), .B(new_n4507_), .ZN(new_n4508_));
  AOI21_X1   g02073(.A1(new_n4508_), .A2(pi0056), .B(pi0062), .ZN(new_n4509_));
  AOI21_X1   g02074(.A1(new_n4506_), .A2(new_n4509_), .B(new_n4441_), .ZN(new_n4510_));
  AOI21_X1   g02075(.A1(new_n4435_), .A2(new_n3500_), .B(new_n4413_), .ZN(new_n4511_));
  NOR3_X1    g02076(.A1(new_n4511_), .A2(pi0215), .A3(new_n4411_), .ZN(new_n4512_));
  NOR2_X1    g02077(.A1(new_n4512_), .A2(new_n4424_), .ZN(new_n4513_));
  INV_X1     g02078(.I(new_n4513_), .ZN(new_n4514_));
  NOR2_X1    g02079(.A1(new_n4514_), .A2(new_n3472_), .ZN(new_n4515_));
  NOR2_X1    g02080(.A1(new_n4425_), .A2(new_n4427_), .ZN(new_n4516_));
  NOR2_X1    g02081(.A1(new_n4516_), .A2(new_n3320_), .ZN(new_n4517_));
  OAI21_X1   g02082(.A1(new_n4515_), .A2(new_n4517_), .B(pi0062), .ZN(new_n4518_));
  NAND3_X1   g02083(.A1(new_n4518_), .A2(pi0246), .A3(new_n3291_), .ZN(new_n4519_));
  NOR2_X1    g02084(.A1(new_n4514_), .A2(new_n2612_), .ZN(new_n4520_));
  NOR2_X1    g02085(.A1(new_n4516_), .A2(new_n2611_), .ZN(new_n4521_));
  OAI21_X1   g02086(.A1(new_n4520_), .A2(new_n4521_), .B(pi0055), .ZN(new_n4522_));
  NOR2_X1    g02087(.A1(new_n4455_), .A2(new_n3339_), .ZN(new_n4523_));
  OAI21_X1   g02088(.A1(new_n4516_), .A2(new_n2628_), .B(new_n4523_), .ZN(new_n4524_));
  INV_X1     g02089(.I(new_n4524_), .ZN(new_n4525_));
  AOI21_X1   g02090(.A1(new_n4525_), .A2(new_n2563_), .B(pi0055), .ZN(new_n4526_));
  AOI21_X1   g02091(.A1(new_n4525_), .A2(pi0038), .B(pi0100), .ZN(new_n4527_));
  INV_X1     g02092(.I(new_n4523_), .ZN(new_n4528_));
  AOI21_X1   g02093(.A1(new_n4513_), .A2(pi0299), .B(new_n4528_), .ZN(new_n4529_));
  OAI21_X1   g02094(.A1(new_n4529_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n4530_));
  NOR2_X1    g02095(.A1(new_n3657_), .A2(new_n4416_), .ZN(new_n4531_));
  NOR2_X1    g02096(.A1(new_n3731_), .A2(pi0877), .ZN(new_n4532_));
  OAI21_X1   g02097(.A1(new_n4531_), .A2(new_n4532_), .B(pi0169), .ZN(new_n4533_));
  OAI21_X1   g02098(.A1(new_n3404_), .A2(pi0877), .B(new_n4414_), .ZN(new_n4534_));
  AOI21_X1   g02099(.A1(new_n4533_), .A2(new_n4534_), .B(pi0228), .ZN(new_n4535_));
  NOR3_X1    g02100(.A1(new_n4535_), .A2(new_n3388_), .A3(new_n4432_), .ZN(new_n4536_));
  OAI21_X1   g02101(.A1(new_n4536_), .A2(new_n4413_), .B(new_n4410_), .ZN(new_n4537_));
  OAI21_X1   g02102(.A1(new_n4537_), .A2(pi0215), .B(new_n4431_), .ZN(new_n4538_));
  AOI21_X1   g02103(.A1(new_n4538_), .A2(pi0299), .B(new_n4476_), .ZN(new_n4539_));
  OAI21_X1   g02104(.A1(new_n4539_), .A2(new_n4530_), .B(new_n4527_), .ZN(new_n4540_));
  AOI21_X1   g02105(.A1(new_n4525_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n4541_));
  AND3_X2    g02106(.A1(new_n4490_), .A2(new_n3500_), .A3(new_n4420_), .Z(new_n4542_));
  OAI21_X1   g02107(.A1(new_n4542_), .A2(new_n4413_), .B(new_n2436_), .ZN(new_n4543_));
  OAI21_X1   g02108(.A1(new_n4543_), .A2(new_n4411_), .B(new_n4486_), .ZN(new_n4544_));
  NAND3_X1   g02109(.A1(new_n4544_), .A2(new_n2572_), .A3(new_n4523_), .ZN(new_n4545_));
  NAND2_X1   g02110(.A1(new_n4545_), .A2(new_n4541_), .ZN(new_n4546_));
  NAND3_X1   g02111(.A1(new_n4540_), .A2(new_n3458_), .A3(new_n4546_), .ZN(new_n4547_));
  NOR2_X1    g02112(.A1(new_n4529_), .A2(new_n3273_), .ZN(new_n4548_));
  AOI21_X1   g02113(.A1(new_n3273_), .A2(new_n4524_), .B(new_n4548_), .ZN(new_n4549_));
  NAND2_X1   g02114(.A1(new_n4549_), .A2(pi0087), .ZN(new_n4550_));
  AOI21_X1   g02115(.A1(new_n4547_), .A2(new_n4550_), .B(pi0075), .ZN(new_n4551_));
  OAI21_X1   g02116(.A1(new_n4524_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4552_));
  NOR2_X1    g02117(.A1(new_n4549_), .A2(new_n2565_), .ZN(new_n4553_));
  AOI21_X1   g02118(.A1(new_n2565_), .A2(new_n4524_), .B(new_n4553_), .ZN(new_n4554_));
  OAI22_X1   g02119(.A1(new_n4551_), .A2(new_n4552_), .B1(new_n3444_), .B2(new_n4554_), .ZN(new_n4555_));
  OAI21_X1   g02120(.A1(new_n4555_), .A2(new_n2563_), .B(new_n4526_), .ZN(new_n4556_));
  NAND3_X1   g02121(.A1(new_n4556_), .A2(new_n3284_), .A3(new_n4522_), .ZN(new_n4557_));
  NAND2_X1   g02122(.A1(new_n4516_), .A2(new_n2577_), .ZN(new_n4558_));
  OAI21_X1   g02123(.A1(new_n4513_), .A2(new_n2577_), .B(new_n4558_), .ZN(new_n4559_));
  AOI21_X1   g02124(.A1(new_n4559_), .A2(pi0056), .B(pi0062), .ZN(new_n4560_));
  AOI21_X1   g02125(.A1(new_n4557_), .A2(new_n4560_), .B(new_n4519_), .ZN(new_n4561_));
  NOR3_X1    g02126(.A1(new_n4510_), .A2(new_n4561_), .A3(new_n4429_), .ZN(po0161));
  INV_X1     g02127(.I(pi0933), .ZN(new_n4563_));
  NOR2_X1    g02128(.A1(new_n2447_), .A2(new_n4563_), .ZN(new_n4564_));
  INV_X1     g02129(.I(pi1137), .ZN(new_n4565_));
  NOR2_X1    g02130(.A1(new_n2444_), .A2(new_n4565_), .ZN(new_n4566_));
  OAI21_X1   g02131(.A1(new_n4564_), .A2(new_n4566_), .B(pi0221), .ZN(new_n4567_));
  INV_X1     g02132(.I(new_n4567_), .ZN(new_n4568_));
  AOI21_X1   g02133(.A1(pi0216), .A2(pi0280), .B(pi0221), .ZN(new_n4569_));
  INV_X1     g02134(.I(new_n4569_), .ZN(new_n4570_));
  INV_X1     g02135(.I(pi0168), .ZN(new_n4571_));
  NAND2_X1   g02136(.A1(new_n2457_), .A2(new_n4571_), .ZN(new_n4572_));
  INV_X1     g02137(.I(pi0878), .ZN(new_n4573_));
  NOR2_X1    g02138(.A1(new_n2463_), .A2(new_n4573_), .ZN(new_n4574_));
  NAND2_X1   g02139(.A1(new_n4574_), .A2(pi0105), .ZN(new_n4575_));
  AOI21_X1   g02140(.A1(new_n4575_), .A2(new_n4572_), .B(new_n2458_), .ZN(new_n4576_));
  NOR2_X1    g02141(.A1(new_n4576_), .A2(pi0216), .ZN(new_n4577_));
  NAND2_X1   g02142(.A1(new_n4571_), .A2(new_n2458_), .ZN(new_n4578_));
  AOI21_X1   g02143(.A1(new_n4577_), .A2(new_n4578_), .B(new_n4570_), .ZN(new_n4579_));
  NOR3_X1    g02144(.A1(new_n4579_), .A2(pi0215), .A3(new_n4568_), .ZN(new_n4580_));
  NOR2_X1    g02145(.A1(new_n2436_), .A2(pi1137), .ZN(new_n4581_));
  NOR2_X1    g02146(.A1(new_n4580_), .A2(new_n4581_), .ZN(new_n4582_));
  INV_X1     g02147(.I(new_n4582_), .ZN(new_n4583_));
  AOI21_X1   g02148(.A1(pi0216), .A2(pi0280), .B(new_n3502_), .ZN(new_n4584_));
  NAND2_X1   g02149(.A1(new_n4584_), .A2(pi0240), .ZN(new_n4585_));
  AND3_X2    g02150(.A1(new_n4583_), .A2(new_n3425_), .A3(new_n4585_), .Z(new_n4586_));
  INV_X1     g02151(.I(pi0240), .ZN(new_n4587_));
  INV_X1     g02152(.I(new_n4581_), .ZN(new_n4588_));
  INV_X1     g02153(.I(new_n4577_), .ZN(new_n4589_));
  NAND2_X1   g02154(.A1(new_n2530_), .A2(new_n4571_), .ZN(new_n4590_));
  OAI21_X1   g02155(.A1(new_n4573_), .A2(new_n2530_), .B(new_n4590_), .ZN(new_n4591_));
  AOI21_X1   g02156(.A1(new_n4591_), .A2(new_n2458_), .B(new_n4589_), .ZN(new_n4592_));
  OAI21_X1   g02157(.A1(new_n4592_), .A2(new_n4570_), .B(new_n4567_), .ZN(new_n4593_));
  OAI21_X1   g02158(.A1(new_n4593_), .A2(pi0215), .B(new_n4588_), .ZN(new_n4594_));
  NOR2_X1    g02159(.A1(new_n4594_), .A2(new_n3472_), .ZN(new_n4595_));
  NOR2_X1    g02160(.A1(new_n4583_), .A2(new_n3320_), .ZN(new_n4596_));
  OAI21_X1   g02161(.A1(new_n4595_), .A2(new_n4596_), .B(pi0062), .ZN(new_n4597_));
  NAND3_X1   g02162(.A1(new_n4597_), .A2(new_n4587_), .A3(new_n3291_), .ZN(new_n4598_));
  NOR2_X1    g02163(.A1(new_n4594_), .A2(new_n2612_), .ZN(new_n4599_));
  NOR2_X1    g02164(.A1(new_n4583_), .A2(new_n2611_), .ZN(new_n4600_));
  OAI21_X1   g02165(.A1(new_n4599_), .A2(new_n4600_), .B(pi0055), .ZN(new_n4601_));
  NOR2_X1    g02166(.A1(new_n2635_), .A2(new_n4563_), .ZN(new_n4602_));
  NOR2_X1    g02167(.A1(new_n2634_), .A2(new_n4565_), .ZN(new_n4603_));
  OAI21_X1   g02168(.A1(new_n4602_), .A2(new_n4603_), .B(pi0222), .ZN(new_n4604_));
  INV_X1     g02169(.I(new_n4604_), .ZN(new_n4605_));
  AOI21_X1   g02170(.A1(pi0224), .A2(pi0280), .B(pi0222), .ZN(new_n4606_));
  INV_X1     g02171(.I(new_n4606_), .ZN(new_n4607_));
  NOR2_X1    g02172(.A1(new_n4574_), .A2(pi0224), .ZN(new_n4608_));
  NOR2_X1    g02173(.A1(new_n4608_), .A2(new_n4607_), .ZN(new_n4609_));
  OAI21_X1   g02174(.A1(new_n4605_), .A2(new_n4609_), .B(new_n2668_), .ZN(new_n4610_));
  NAND2_X1   g02175(.A1(pi0223), .A2(pi1137), .ZN(new_n4611_));
  AOI21_X1   g02176(.A1(new_n4610_), .A2(new_n4611_), .B(pi0299), .ZN(new_n4612_));
  AOI21_X1   g02177(.A1(new_n4582_), .A2(pi0299), .B(new_n4612_), .ZN(new_n4613_));
  AOI21_X1   g02178(.A1(new_n4613_), .A2(new_n2563_), .B(pi0055), .ZN(new_n4614_));
  NAND2_X1   g02179(.A1(new_n3387_), .A2(pi0878), .ZN(new_n4615_));
  NAND3_X1   g02180(.A1(new_n3657_), .A2(new_n4571_), .A3(new_n4615_), .ZN(new_n4616_));
  NOR2_X1    g02181(.A1(new_n3387_), .A2(pi0168), .ZN(new_n4617_));
  NOR2_X1    g02182(.A1(new_n3404_), .A2(new_n4571_), .ZN(new_n4618_));
  OAI21_X1   g02183(.A1(new_n4618_), .A2(new_n4617_), .B(pi0878), .ZN(new_n4619_));
  AOI21_X1   g02184(.A1(new_n4619_), .A2(new_n4616_), .B(pi0228), .ZN(new_n4620_));
  NAND2_X1   g02185(.A1(new_n3729_), .A2(new_n4576_), .ZN(new_n4621_));
  NAND2_X1   g02186(.A1(new_n4621_), .A2(new_n2614_), .ZN(new_n4622_));
  OAI21_X1   g02187(.A1(new_n4620_), .A2(new_n4622_), .B(new_n4569_), .ZN(new_n4623_));
  NAND3_X1   g02188(.A1(new_n4623_), .A2(new_n2436_), .A3(new_n4567_), .ZN(new_n4624_));
  AOI21_X1   g02189(.A1(new_n4624_), .A2(new_n4588_), .B(new_n2628_), .ZN(new_n4625_));
  NAND2_X1   g02190(.A1(new_n4611_), .A2(new_n2628_), .ZN(new_n4626_));
  OAI21_X1   g02191(.A1(new_n3392_), .A2(new_n4573_), .B(new_n2631_), .ZN(new_n4627_));
  AOI21_X1   g02192(.A1(new_n4627_), .A2(new_n4606_), .B(new_n4605_), .ZN(new_n4628_));
  INV_X1     g02193(.I(new_n4628_), .ZN(new_n4629_));
  INV_X1     g02194(.I(new_n4626_), .ZN(new_n4630_));
  AOI21_X1   g02195(.A1(new_n3392_), .A2(new_n4606_), .B(new_n4629_), .ZN(new_n4631_));
  OAI21_X1   g02196(.A1(new_n4631_), .A2(pi0223), .B(new_n4630_), .ZN(new_n4632_));
  NAND2_X1   g02197(.A1(new_n4632_), .A2(new_n2627_), .ZN(new_n4633_));
  INV_X1     g02198(.I(new_n4633_), .ZN(new_n4634_));
  OAI21_X1   g02199(.A1(new_n4626_), .A2(new_n4629_), .B(new_n4634_), .ZN(new_n4635_));
  INV_X1     g02200(.I(new_n4594_), .ZN(new_n4636_));
  AOI21_X1   g02201(.A1(new_n4636_), .A2(pi0299), .B(new_n4612_), .ZN(new_n4637_));
  OAI22_X1   g02202(.A1(new_n4625_), .A2(new_n4635_), .B1(new_n2627_), .B2(new_n4637_), .ZN(new_n4638_));
  AOI21_X1   g02203(.A1(new_n4613_), .A2(pi0038), .B(pi0100), .ZN(new_n4639_));
  OAI21_X1   g02204(.A1(new_n4638_), .A2(pi0038), .B(new_n4639_), .ZN(new_n4640_));
  AOI21_X1   g02205(.A1(new_n4613_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n4641_));
  INV_X1     g02206(.I(new_n4612_), .ZN(new_n4642_));
  NOR2_X1    g02207(.A1(new_n4581_), .A2(new_n2628_), .ZN(new_n4643_));
  INV_X1     g02208(.I(new_n4643_), .ZN(new_n4644_));
  NOR2_X1    g02209(.A1(new_n3371_), .A2(pi0168), .ZN(new_n4645_));
  NOR2_X1    g02210(.A1(new_n3544_), .A2(new_n4573_), .ZN(new_n4646_));
  OAI21_X1   g02211(.A1(new_n4646_), .A2(new_n4645_), .B(new_n2458_), .ZN(new_n4647_));
  AOI21_X1   g02212(.A1(new_n4647_), .A2(new_n4577_), .B(new_n4570_), .ZN(new_n4648_));
  NOR3_X1    g02213(.A1(new_n4648_), .A2(pi0215), .A3(new_n4568_), .ZN(new_n4649_));
  OAI21_X1   g02214(.A1(new_n4649_), .A2(new_n4644_), .B(new_n4642_), .ZN(new_n4650_));
  OAI21_X1   g02215(.A1(new_n4650_), .A2(new_n2573_), .B(new_n4641_), .ZN(new_n4651_));
  NAND3_X1   g02216(.A1(new_n4640_), .A2(new_n3458_), .A3(new_n4651_), .ZN(new_n4652_));
  INV_X1     g02217(.I(new_n4613_), .ZN(new_n4653_));
  NOR2_X1    g02218(.A1(new_n4637_), .A2(new_n3273_), .ZN(new_n4654_));
  AOI21_X1   g02219(.A1(new_n3273_), .A2(new_n4653_), .B(new_n4654_), .ZN(new_n4655_));
  NAND2_X1   g02220(.A1(new_n4655_), .A2(pi0087), .ZN(new_n4656_));
  AOI21_X1   g02221(.A1(new_n4652_), .A2(new_n4656_), .B(pi0075), .ZN(new_n4657_));
  OAI21_X1   g02222(.A1(new_n4653_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4658_));
  NOR2_X1    g02223(.A1(new_n4655_), .A2(new_n2565_), .ZN(new_n4659_));
  AOI21_X1   g02224(.A1(new_n2565_), .A2(new_n4653_), .B(new_n4659_), .ZN(new_n4660_));
  OAI22_X1   g02225(.A1(new_n4657_), .A2(new_n4658_), .B1(new_n3444_), .B2(new_n4660_), .ZN(new_n4661_));
  OAI21_X1   g02226(.A1(new_n4661_), .A2(new_n2563_), .B(new_n4614_), .ZN(new_n4662_));
  NAND3_X1   g02227(.A1(new_n4662_), .A2(new_n3284_), .A3(new_n4601_), .ZN(new_n4663_));
  NAND2_X1   g02228(.A1(new_n4583_), .A2(new_n2577_), .ZN(new_n4664_));
  OAI21_X1   g02229(.A1(new_n4636_), .A2(new_n2577_), .B(new_n4664_), .ZN(new_n4665_));
  AOI21_X1   g02230(.A1(new_n4665_), .A2(pi0056), .B(pi0062), .ZN(new_n4666_));
  AOI21_X1   g02231(.A1(new_n4663_), .A2(new_n4666_), .B(new_n4598_), .ZN(new_n4667_));
  AOI21_X1   g02232(.A1(new_n4592_), .A2(new_n3500_), .B(new_n4570_), .ZN(new_n4668_));
  NOR3_X1    g02233(.A1(new_n4668_), .A2(pi0215), .A3(new_n4568_), .ZN(new_n4669_));
  NOR2_X1    g02234(.A1(new_n4669_), .A2(new_n4581_), .ZN(new_n4670_));
  INV_X1     g02235(.I(new_n4670_), .ZN(new_n4671_));
  NOR2_X1    g02236(.A1(new_n4671_), .A2(new_n3472_), .ZN(new_n4672_));
  NOR2_X1    g02237(.A1(new_n4582_), .A2(new_n4584_), .ZN(new_n4673_));
  NOR2_X1    g02238(.A1(new_n4673_), .A2(new_n3320_), .ZN(new_n4674_));
  OAI21_X1   g02239(.A1(new_n4672_), .A2(new_n4674_), .B(pi0062), .ZN(new_n4675_));
  NAND3_X1   g02240(.A1(new_n4675_), .A2(pi0240), .A3(new_n3291_), .ZN(new_n4676_));
  NOR2_X1    g02241(.A1(new_n4671_), .A2(new_n2612_), .ZN(new_n4677_));
  NOR2_X1    g02242(.A1(new_n4673_), .A2(new_n2611_), .ZN(new_n4678_));
  OAI21_X1   g02243(.A1(new_n4677_), .A2(new_n4678_), .B(pi0055), .ZN(new_n4679_));
  NOR2_X1    g02244(.A1(new_n4612_), .A2(new_n3339_), .ZN(new_n4680_));
  OAI21_X1   g02245(.A1(new_n4673_), .A2(new_n2628_), .B(new_n4680_), .ZN(new_n4681_));
  INV_X1     g02246(.I(new_n4681_), .ZN(new_n4682_));
  AOI21_X1   g02247(.A1(new_n4682_), .A2(new_n2563_), .B(pi0055), .ZN(new_n4683_));
  AOI21_X1   g02248(.A1(new_n4682_), .A2(pi0038), .B(pi0100), .ZN(new_n4684_));
  INV_X1     g02249(.I(new_n4680_), .ZN(new_n4685_));
  AOI21_X1   g02250(.A1(new_n4670_), .A2(pi0299), .B(new_n4685_), .ZN(new_n4686_));
  OAI21_X1   g02251(.A1(new_n4686_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n4687_));
  NOR2_X1    g02252(.A1(new_n3657_), .A2(new_n4573_), .ZN(new_n4688_));
  NOR2_X1    g02253(.A1(new_n3731_), .A2(pi0878), .ZN(new_n4689_));
  OAI21_X1   g02254(.A1(new_n4688_), .A2(new_n4689_), .B(pi0168), .ZN(new_n4690_));
  OAI21_X1   g02255(.A1(new_n3404_), .A2(pi0878), .B(new_n4571_), .ZN(new_n4691_));
  AOI21_X1   g02256(.A1(new_n4690_), .A2(new_n4691_), .B(pi0228), .ZN(new_n4692_));
  NOR3_X1    g02257(.A1(new_n4692_), .A2(new_n3388_), .A3(new_n4589_), .ZN(new_n4693_));
  OAI21_X1   g02258(.A1(new_n4693_), .A2(new_n4570_), .B(new_n4567_), .ZN(new_n4694_));
  OAI21_X1   g02259(.A1(new_n4694_), .A2(pi0215), .B(new_n4588_), .ZN(new_n4695_));
  AOI21_X1   g02260(.A1(new_n4695_), .A2(pi0299), .B(new_n4633_), .ZN(new_n4696_));
  OAI21_X1   g02261(.A1(new_n4696_), .A2(new_n4687_), .B(new_n4684_), .ZN(new_n4697_));
  AOI21_X1   g02262(.A1(new_n4682_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n4698_));
  AND3_X2    g02263(.A1(new_n4647_), .A2(new_n3500_), .A3(new_n4577_), .Z(new_n4699_));
  OAI21_X1   g02264(.A1(new_n4699_), .A2(new_n4570_), .B(new_n2436_), .ZN(new_n4700_));
  OAI21_X1   g02265(.A1(new_n4700_), .A2(new_n4568_), .B(new_n4643_), .ZN(new_n4701_));
  NAND3_X1   g02266(.A1(new_n4701_), .A2(new_n2572_), .A3(new_n4680_), .ZN(new_n4702_));
  NAND2_X1   g02267(.A1(new_n4702_), .A2(new_n4698_), .ZN(new_n4703_));
  NAND3_X1   g02268(.A1(new_n4697_), .A2(new_n3458_), .A3(new_n4703_), .ZN(new_n4704_));
  NOR2_X1    g02269(.A1(new_n4686_), .A2(new_n3273_), .ZN(new_n4705_));
  AOI21_X1   g02270(.A1(new_n3273_), .A2(new_n4681_), .B(new_n4705_), .ZN(new_n4706_));
  NAND2_X1   g02271(.A1(new_n4706_), .A2(pi0087), .ZN(new_n4707_));
  AOI21_X1   g02272(.A1(new_n4704_), .A2(new_n4707_), .B(pi0075), .ZN(new_n4708_));
  OAI21_X1   g02273(.A1(new_n4681_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4709_));
  NOR2_X1    g02274(.A1(new_n4706_), .A2(new_n2565_), .ZN(new_n4710_));
  AOI21_X1   g02275(.A1(new_n2565_), .A2(new_n4681_), .B(new_n4710_), .ZN(new_n4711_));
  OAI22_X1   g02276(.A1(new_n4708_), .A2(new_n4709_), .B1(new_n3444_), .B2(new_n4711_), .ZN(new_n4712_));
  OAI21_X1   g02277(.A1(new_n4712_), .A2(new_n2563_), .B(new_n4683_), .ZN(new_n4713_));
  NAND3_X1   g02278(.A1(new_n4713_), .A2(new_n3284_), .A3(new_n4679_), .ZN(new_n4714_));
  NAND2_X1   g02279(.A1(new_n4673_), .A2(new_n2577_), .ZN(new_n4715_));
  OAI21_X1   g02280(.A1(new_n4670_), .A2(new_n2577_), .B(new_n4715_), .ZN(new_n4716_));
  AOI21_X1   g02281(.A1(new_n4716_), .A2(pi0056), .B(pi0062), .ZN(new_n4717_));
  AOI21_X1   g02282(.A1(new_n4714_), .A2(new_n4717_), .B(new_n4676_), .ZN(new_n4718_));
  NOR3_X1    g02283(.A1(new_n4667_), .A2(new_n4718_), .A3(new_n4586_), .ZN(po0162));
  NOR2_X1    g02284(.A1(new_n2436_), .A2(pi1136), .ZN(new_n4720_));
  INV_X1     g02285(.I(new_n4720_), .ZN(new_n4721_));
  INV_X1     g02286(.I(pi0928), .ZN(new_n4722_));
  NOR2_X1    g02287(.A1(new_n2447_), .A2(new_n4722_), .ZN(new_n4723_));
  INV_X1     g02288(.I(pi1136), .ZN(new_n4724_));
  NOR2_X1    g02289(.A1(new_n2444_), .A2(new_n4724_), .ZN(new_n4725_));
  OAI21_X1   g02290(.A1(new_n4723_), .A2(new_n4725_), .B(pi0221), .ZN(new_n4726_));
  INV_X1     g02291(.I(pi0266), .ZN(new_n4727_));
  NOR2_X1    g02292(.A1(new_n2614_), .A2(new_n4727_), .ZN(new_n4728_));
  INV_X1     g02293(.I(pi0875), .ZN(new_n4729_));
  NAND2_X1   g02294(.A1(new_n2530_), .A2(pi0166), .ZN(new_n4730_));
  OAI21_X1   g02295(.A1(new_n4729_), .A2(new_n2530_), .B(new_n4730_), .ZN(new_n4731_));
  NOR2_X1    g02296(.A1(new_n3361_), .A2(pi0105), .ZN(new_n4732_));
  NOR2_X1    g02297(.A1(new_n2463_), .A2(new_n4729_), .ZN(new_n4733_));
  AOI21_X1   g02298(.A1(new_n4733_), .A2(pi0105), .B(new_n4732_), .ZN(new_n4734_));
  NOR2_X1    g02299(.A1(new_n4734_), .A2(new_n2458_), .ZN(new_n4735_));
  AOI21_X1   g02300(.A1(new_n4731_), .A2(new_n2458_), .B(new_n4735_), .ZN(new_n4736_));
  AOI21_X1   g02301(.A1(new_n4736_), .A2(new_n3500_), .B(pi0216), .ZN(new_n4737_));
  OAI21_X1   g02302(.A1(new_n4737_), .A2(new_n4728_), .B(new_n2441_), .ZN(new_n4738_));
  NAND3_X1   g02303(.A1(new_n4738_), .A2(new_n2436_), .A3(new_n4726_), .ZN(new_n4739_));
  NAND2_X1   g02304(.A1(new_n4739_), .A2(new_n4721_), .ZN(new_n4740_));
  INV_X1     g02305(.I(new_n4740_), .ZN(new_n4741_));
  NAND2_X1   g02306(.A1(new_n4741_), .A2(new_n2611_), .ZN(new_n4742_));
  INV_X1     g02307(.I(new_n4726_), .ZN(new_n4743_));
  INV_X1     g02308(.I(new_n4728_), .ZN(new_n4744_));
  NOR2_X1    g02309(.A1(new_n3361_), .A2(pi0228), .ZN(new_n4745_));
  OAI21_X1   g02310(.A1(new_n4735_), .A2(new_n4745_), .B(new_n2614_), .ZN(new_n4746_));
  AOI21_X1   g02311(.A1(new_n4746_), .A2(new_n4744_), .B(pi0221), .ZN(new_n4747_));
  NOR3_X1    g02312(.A1(new_n4747_), .A2(pi0215), .A3(new_n4743_), .ZN(new_n4748_));
  NOR2_X1    g02313(.A1(new_n4748_), .A2(new_n4720_), .ZN(new_n4749_));
  NOR2_X1    g02314(.A1(new_n4749_), .A2(new_n3307_), .ZN(new_n4750_));
  INV_X1     g02315(.I(new_n4750_), .ZN(new_n4751_));
  NAND2_X1   g02316(.A1(new_n4751_), .A2(new_n2612_), .ZN(new_n4752_));
  AOI21_X1   g02317(.A1(new_n4742_), .A2(new_n4752_), .B(new_n2602_), .ZN(new_n4753_));
  AOI21_X1   g02318(.A1(new_n4727_), .A2(pi0224), .B(pi0222), .ZN(new_n4754_));
  NAND3_X1   g02319(.A1(new_n3028_), .A2(new_n2631_), .A3(new_n4729_), .ZN(new_n4755_));
  AND2_X2    g02320(.A1(new_n4755_), .A2(new_n4754_), .Z(new_n4756_));
  NAND2_X1   g02321(.A1(new_n2634_), .A2(pi0928), .ZN(new_n4757_));
  NAND2_X1   g02322(.A1(new_n2635_), .A2(pi1136), .ZN(new_n4758_));
  AOI21_X1   g02323(.A1(new_n4758_), .A2(new_n4757_), .B(new_n2629_), .ZN(new_n4759_));
  OAI21_X1   g02324(.A1(new_n4756_), .A2(new_n4759_), .B(new_n2668_), .ZN(new_n4760_));
  NAND2_X1   g02325(.A1(pi0223), .A2(pi1136), .ZN(new_n4761_));
  AOI21_X1   g02326(.A1(new_n4760_), .A2(new_n4761_), .B(pi0299), .ZN(new_n4762_));
  AOI21_X1   g02327(.A1(new_n4751_), .A2(pi0299), .B(new_n4762_), .ZN(new_n4763_));
  INV_X1     g02328(.I(new_n4763_), .ZN(new_n4764_));
  OAI21_X1   g02329(.A1(new_n4764_), .A2(new_n2562_), .B(new_n2602_), .ZN(new_n4765_));
  OAI21_X1   g02330(.A1(new_n4764_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n4766_));
  AOI21_X1   g02331(.A1(new_n4741_), .A2(pi0299), .B(new_n4762_), .ZN(new_n4767_));
  OAI21_X1   g02332(.A1(new_n4767_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n4768_));
  NOR2_X1    g02333(.A1(new_n3728_), .A2(new_n2458_), .ZN(new_n4769_));
  AOI21_X1   g02334(.A1(new_n4769_), .A2(new_n4734_), .B(pi0216), .ZN(new_n4770_));
  NAND2_X1   g02335(.A1(new_n3404_), .A2(pi0166), .ZN(new_n4771_));
  NAND2_X1   g02336(.A1(new_n3387_), .A2(new_n3361_), .ZN(new_n4772_));
  AOI21_X1   g02337(.A1(new_n4771_), .A2(new_n4772_), .B(pi0875), .ZN(new_n4773_));
  OAI21_X1   g02338(.A1(new_n3451_), .A2(pi0166), .B(pi0875), .ZN(new_n4774_));
  NAND2_X1   g02339(.A1(new_n4774_), .A2(new_n2458_), .ZN(new_n4775_));
  OAI21_X1   g02340(.A1(new_n4773_), .A2(new_n4775_), .B(new_n4770_), .ZN(new_n4776_));
  AOI21_X1   g02341(.A1(new_n4776_), .A2(new_n4744_), .B(pi0221), .ZN(new_n4777_));
  NOR3_X1    g02342(.A1(new_n4777_), .A2(pi0215), .A3(new_n4743_), .ZN(new_n4778_));
  OAI21_X1   g02343(.A1(new_n4778_), .A2(new_n4720_), .B(pi0299), .ZN(new_n4779_));
  NAND2_X1   g02344(.A1(new_n4761_), .A2(new_n2628_), .ZN(new_n4780_));
  INV_X1     g02345(.I(new_n4780_), .ZN(new_n4781_));
  NOR2_X1    g02346(.A1(new_n3381_), .A2(new_n2642_), .ZN(new_n4782_));
  OR3_X2     g02347(.A1(new_n4782_), .A2(new_n4756_), .A3(new_n4759_), .Z(new_n4783_));
  NAND2_X1   g02348(.A1(new_n4783_), .A2(new_n2668_), .ZN(new_n4784_));
  AOI21_X1   g02349(.A1(new_n4784_), .A2(new_n4781_), .B(pi0039), .ZN(new_n4785_));
  AOI21_X1   g02350(.A1(new_n4779_), .A2(new_n4785_), .B(new_n4768_), .ZN(new_n4786_));
  OAI21_X1   g02351(.A1(new_n4764_), .A2(new_n2572_), .B(pi0100), .ZN(new_n4787_));
  NAND2_X1   g02352(.A1(new_n3362_), .A2(new_n2688_), .ZN(new_n4788_));
  NAND2_X1   g02353(.A1(new_n3365_), .A2(new_n2689_), .ZN(new_n4789_));
  NAND2_X1   g02354(.A1(new_n4789_), .A2(new_n4788_), .ZN(new_n4790_));
  NAND2_X1   g02355(.A1(new_n3365_), .A2(new_n4729_), .ZN(new_n4791_));
  AOI22_X1   g02356(.A1(new_n4790_), .A2(pi0875), .B1(pi0166), .B2(new_n4791_), .ZN(new_n4792_));
  NOR2_X1    g02357(.A1(new_n4792_), .A2(pi0228), .ZN(new_n4793_));
  NOR2_X1    g02358(.A1(new_n4793_), .A2(new_n4735_), .ZN(new_n4794_));
  NAND2_X1   g02359(.A1(new_n4794_), .A2(new_n3500_), .ZN(new_n4795_));
  AOI21_X1   g02360(.A1(new_n4795_), .A2(new_n2614_), .B(new_n4728_), .ZN(new_n4796_));
  OAI21_X1   g02361(.A1(new_n4796_), .A2(pi0221), .B(new_n2436_), .ZN(new_n4797_));
  OAI21_X1   g02362(.A1(new_n4797_), .A2(new_n4743_), .B(new_n4721_), .ZN(new_n4798_));
  OAI21_X1   g02363(.A1(new_n4798_), .A2(new_n2628_), .B(new_n2572_), .ZN(new_n4799_));
  NOR2_X1    g02364(.A1(new_n4799_), .A2(new_n4762_), .ZN(new_n4800_));
  OAI22_X1   g02365(.A1(new_n4786_), .A2(new_n4766_), .B1(new_n4787_), .B2(new_n4800_), .ZN(new_n4801_));
  NOR2_X1    g02366(.A1(new_n4767_), .A2(new_n3273_), .ZN(new_n4802_));
  AOI21_X1   g02367(.A1(new_n3273_), .A2(new_n4764_), .B(new_n4802_), .ZN(new_n4803_));
  NAND2_X1   g02368(.A1(new_n4803_), .A2(pi0087), .ZN(new_n4804_));
  OAI21_X1   g02369(.A1(new_n4801_), .A2(pi0087), .B(new_n4804_), .ZN(new_n4805_));
  OAI21_X1   g02370(.A1(new_n4764_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n4806_));
  AOI21_X1   g02371(.A1(new_n4805_), .A2(new_n3465_), .B(new_n4806_), .ZN(new_n4807_));
  NAND2_X1   g02372(.A1(new_n4764_), .A2(new_n2565_), .ZN(new_n4808_));
  OR2_X2     g02373(.A1(new_n4803_), .A2(new_n2565_), .Z(new_n4809_));
  AOI21_X1   g02374(.A1(new_n4809_), .A2(new_n4808_), .B(new_n3444_), .ZN(new_n4810_));
  NOR3_X1    g02375(.A1(new_n4807_), .A2(new_n2563_), .A3(new_n4810_), .ZN(new_n4811_));
  OAI21_X1   g02376(.A1(new_n4811_), .A2(new_n4765_), .B(new_n3284_), .ZN(new_n4812_));
  NOR2_X1    g02377(.A1(new_n4751_), .A2(new_n2576_), .ZN(new_n4813_));
  AOI21_X1   g02378(.A1(new_n4740_), .A2(new_n2576_), .B(new_n4813_), .ZN(new_n4814_));
  OAI22_X1   g02379(.A1(new_n4812_), .A2(new_n4753_), .B1(new_n3284_), .B2(new_n4814_), .ZN(new_n4815_));
  NAND2_X1   g02380(.A1(new_n4751_), .A2(new_n3472_), .ZN(new_n4816_));
  OAI21_X1   g02381(.A1(new_n4740_), .A2(new_n3472_), .B(new_n4816_), .ZN(new_n4817_));
  NAND2_X1   g02382(.A1(new_n4817_), .A2(pi0062), .ZN(new_n4818_));
  OAI21_X1   g02383(.A1(new_n4815_), .A2(pi0062), .B(new_n4818_), .ZN(new_n4819_));
  NOR2_X1    g02384(.A1(new_n4819_), .A2(new_n3425_), .ZN(new_n4820_));
  OAI21_X1   g02385(.A1(new_n4751_), .A2(new_n3291_), .B(pi0245), .ZN(new_n4821_));
  NAND2_X1   g02386(.A1(new_n4727_), .A2(pi0216), .ZN(new_n4822_));
  NAND2_X1   g02387(.A1(new_n4736_), .A2(new_n2614_), .ZN(new_n4823_));
  NAND3_X1   g02388(.A1(new_n4823_), .A2(new_n2441_), .A3(new_n4822_), .ZN(new_n4824_));
  NAND3_X1   g02389(.A1(new_n4824_), .A2(new_n2436_), .A3(new_n4726_), .ZN(new_n4825_));
  NAND2_X1   g02390(.A1(new_n4825_), .A2(new_n4721_), .ZN(new_n4826_));
  INV_X1     g02391(.I(new_n4826_), .ZN(new_n4827_));
  NAND2_X1   g02392(.A1(new_n4827_), .A2(new_n2611_), .ZN(new_n4828_));
  NAND2_X1   g02393(.A1(new_n4749_), .A2(new_n2612_), .ZN(new_n4829_));
  AOI21_X1   g02394(.A1(new_n4828_), .A2(new_n4829_), .B(new_n2602_), .ZN(new_n4830_));
  OAI21_X1   g02395(.A1(new_n2644_), .A2(new_n4733_), .B(new_n4762_), .ZN(new_n4831_));
  INV_X1     g02396(.I(new_n4831_), .ZN(new_n4832_));
  AOI21_X1   g02397(.A1(new_n4749_), .A2(pi0299), .B(new_n4832_), .ZN(new_n4833_));
  INV_X1     g02398(.I(new_n4833_), .ZN(new_n4834_));
  OAI21_X1   g02399(.A1(new_n4834_), .A2(new_n2562_), .B(new_n2602_), .ZN(new_n4835_));
  OAI21_X1   g02400(.A1(new_n4826_), .A2(new_n2628_), .B(new_n4831_), .ZN(new_n4836_));
  AOI21_X1   g02401(.A1(new_n4836_), .A2(pi0039), .B(pi0038), .ZN(new_n4837_));
  INV_X1     g02402(.I(new_n4770_), .ZN(new_n4838_));
  NOR2_X1    g02403(.A1(new_n3387_), .A2(new_n3361_), .ZN(new_n4839_));
  AOI21_X1   g02404(.A1(new_n3403_), .A2(new_n3361_), .B(new_n4839_), .ZN(new_n4840_));
  NAND2_X1   g02405(.A1(new_n4729_), .A2(pi0166), .ZN(new_n4841_));
  OAI22_X1   g02406(.A1(new_n4840_), .A2(new_n4729_), .B1(new_n3451_), .B2(new_n4841_), .ZN(new_n4842_));
  AOI21_X1   g02407(.A1(new_n4842_), .A2(new_n2458_), .B(new_n4769_), .ZN(new_n4843_));
  OAI21_X1   g02408(.A1(new_n4843_), .A2(new_n4838_), .B(new_n4744_), .ZN(new_n4844_));
  AOI21_X1   g02409(.A1(new_n4844_), .A2(new_n2441_), .B(new_n4743_), .ZN(new_n4845_));
  AOI21_X1   g02410(.A1(new_n4845_), .A2(new_n2436_), .B(new_n4720_), .ZN(new_n4846_));
  INV_X1     g02411(.I(new_n4759_), .ZN(new_n4847_));
  INV_X1     g02412(.I(new_n4785_), .ZN(new_n4848_));
  INV_X1     g02413(.I(new_n4782_), .ZN(new_n4849_));
  AOI21_X1   g02414(.A1(new_n4849_), .A2(new_n4756_), .B(new_n4780_), .ZN(new_n4850_));
  AOI21_X1   g02415(.A1(new_n4847_), .A2(new_n4850_), .B(new_n4848_), .ZN(new_n4851_));
  OAI21_X1   g02416(.A1(new_n4846_), .A2(new_n2628_), .B(new_n4851_), .ZN(new_n4852_));
  OAI21_X1   g02417(.A1(new_n4834_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n4853_));
  AOI21_X1   g02418(.A1(new_n4852_), .A2(new_n4837_), .B(new_n4853_), .ZN(new_n4854_));
  OAI21_X1   g02419(.A1(new_n4834_), .A2(new_n2572_), .B(pi0100), .ZN(new_n4855_));
  NOR2_X1    g02420(.A1(new_n4720_), .A2(new_n2628_), .ZN(new_n4856_));
  NAND2_X1   g02421(.A1(new_n4794_), .A2(new_n2614_), .ZN(new_n4857_));
  NAND3_X1   g02422(.A1(new_n4857_), .A2(new_n2441_), .A3(new_n4822_), .ZN(new_n4858_));
  NAND3_X1   g02423(.A1(new_n4858_), .A2(new_n2436_), .A3(new_n4726_), .ZN(new_n4859_));
  AOI21_X1   g02424(.A1(new_n4859_), .A2(new_n4856_), .B(new_n4832_), .ZN(new_n4860_));
  AOI21_X1   g02425(.A1(new_n4860_), .A2(new_n2572_), .B(new_n4855_), .ZN(new_n4861_));
  NOR3_X1    g02426(.A1(new_n4854_), .A2(pi0087), .A3(new_n4861_), .ZN(new_n4862_));
  NAND2_X1   g02427(.A1(new_n4836_), .A2(new_n3272_), .ZN(new_n4863_));
  OAI21_X1   g02428(.A1(new_n3272_), .A2(new_n4833_), .B(new_n4863_), .ZN(new_n4864_));
  NOR2_X1    g02429(.A1(new_n4864_), .A2(new_n3458_), .ZN(new_n4865_));
  OAI21_X1   g02430(.A1(new_n4862_), .A2(new_n4865_), .B(new_n3465_), .ZN(new_n4866_));
  AOI21_X1   g02431(.A1(new_n4833_), .A2(pi0075), .B(pi0092), .ZN(new_n4867_));
  NAND2_X1   g02432(.A1(new_n4864_), .A2(new_n2564_), .ZN(new_n4868_));
  OAI21_X1   g02433(.A1(new_n2564_), .A2(new_n4833_), .B(new_n4868_), .ZN(new_n4869_));
  AOI22_X1   g02434(.A1(new_n4866_), .A2(new_n4867_), .B1(pi0092), .B2(new_n4869_), .ZN(new_n4870_));
  AOI21_X1   g02435(.A1(new_n4870_), .A2(new_n2562_), .B(new_n4835_), .ZN(new_n4871_));
  NOR3_X1    g02436(.A1(new_n4871_), .A2(pi0056), .A3(new_n4830_), .ZN(new_n4872_));
  NAND2_X1   g02437(.A1(new_n4826_), .A2(new_n2576_), .ZN(new_n4873_));
  OAI21_X1   g02438(.A1(new_n4720_), .A2(new_n4748_), .B(new_n2577_), .ZN(new_n4874_));
  AOI21_X1   g02439(.A1(new_n4873_), .A2(new_n4874_), .B(new_n3284_), .ZN(new_n4875_));
  NOR3_X1    g02440(.A1(new_n4872_), .A2(pi0062), .A3(new_n4875_), .ZN(new_n4876_));
  NAND2_X1   g02441(.A1(new_n4827_), .A2(new_n3320_), .ZN(new_n4877_));
  NAND2_X1   g02442(.A1(new_n3472_), .A2(new_n4749_), .ZN(new_n4878_));
  AOI21_X1   g02443(.A1(new_n4877_), .A2(new_n4878_), .B(new_n3471_), .ZN(new_n4879_));
  NOR3_X1    g02444(.A1(new_n4876_), .A2(new_n3425_), .A3(new_n4879_), .ZN(new_n4880_));
  INV_X1     g02445(.I(pi0245), .ZN(new_n4881_));
  OAI21_X1   g02446(.A1(new_n4749_), .A2(new_n3291_), .B(new_n4881_), .ZN(new_n4882_));
  OAI22_X1   g02447(.A1(new_n4820_), .A2(new_n4821_), .B1(new_n4880_), .B2(new_n4882_), .ZN(po0163));
  NOR2_X1    g02448(.A1(new_n2436_), .A2(pi1135), .ZN(new_n4884_));
  INV_X1     g02449(.I(new_n4884_), .ZN(new_n4885_));
  INV_X1     g02450(.I(pi0938), .ZN(new_n4886_));
  NOR2_X1    g02451(.A1(new_n2447_), .A2(new_n4886_), .ZN(new_n4887_));
  INV_X1     g02452(.I(pi1135), .ZN(new_n4888_));
  NOR2_X1    g02453(.A1(new_n2444_), .A2(new_n4888_), .ZN(new_n4889_));
  OAI21_X1   g02454(.A1(new_n4887_), .A2(new_n4889_), .B(pi0221), .ZN(new_n4890_));
  INV_X1     g02455(.I(pi0279), .ZN(new_n4891_));
  NOR2_X1    g02456(.A1(new_n2614_), .A2(new_n4891_), .ZN(new_n4892_));
  INV_X1     g02457(.I(pi0879), .ZN(new_n4893_));
  NAND2_X1   g02458(.A1(new_n2530_), .A2(pi0161), .ZN(new_n4894_));
  OAI21_X1   g02459(.A1(new_n4893_), .A2(new_n2530_), .B(new_n4894_), .ZN(new_n4895_));
  NOR2_X1    g02460(.A1(new_n3360_), .A2(pi0105), .ZN(new_n4896_));
  NOR2_X1    g02461(.A1(new_n2463_), .A2(new_n4893_), .ZN(new_n4897_));
  AOI21_X1   g02462(.A1(new_n4897_), .A2(pi0105), .B(new_n4896_), .ZN(new_n4898_));
  NOR2_X1    g02463(.A1(new_n4898_), .A2(new_n2458_), .ZN(new_n4899_));
  AOI21_X1   g02464(.A1(new_n4895_), .A2(new_n2458_), .B(new_n4899_), .ZN(new_n4900_));
  AOI21_X1   g02465(.A1(new_n4900_), .A2(new_n3500_), .B(pi0216), .ZN(new_n4901_));
  OAI21_X1   g02466(.A1(new_n4901_), .A2(new_n4892_), .B(new_n2441_), .ZN(new_n4902_));
  NAND3_X1   g02467(.A1(new_n4902_), .A2(new_n2436_), .A3(new_n4890_), .ZN(new_n4903_));
  NAND2_X1   g02468(.A1(new_n4903_), .A2(new_n4885_), .ZN(new_n4904_));
  INV_X1     g02469(.I(new_n4904_), .ZN(new_n4905_));
  NAND2_X1   g02470(.A1(new_n4905_), .A2(new_n2611_), .ZN(new_n4906_));
  INV_X1     g02471(.I(new_n4890_), .ZN(new_n4907_));
  INV_X1     g02472(.I(new_n4892_), .ZN(new_n4908_));
  NOR2_X1    g02473(.A1(new_n3360_), .A2(pi0228), .ZN(new_n4909_));
  OAI21_X1   g02474(.A1(new_n4899_), .A2(new_n4909_), .B(new_n2614_), .ZN(new_n4910_));
  AOI21_X1   g02475(.A1(new_n4910_), .A2(new_n4908_), .B(pi0221), .ZN(new_n4911_));
  NOR3_X1    g02476(.A1(new_n4911_), .A2(pi0215), .A3(new_n4907_), .ZN(new_n4912_));
  NOR2_X1    g02477(.A1(new_n4912_), .A2(new_n4884_), .ZN(new_n4913_));
  NOR2_X1    g02478(.A1(new_n4913_), .A2(new_n3307_), .ZN(new_n4914_));
  INV_X1     g02479(.I(new_n4914_), .ZN(new_n4915_));
  NAND2_X1   g02480(.A1(new_n4915_), .A2(new_n2612_), .ZN(new_n4916_));
  AOI21_X1   g02481(.A1(new_n4906_), .A2(new_n4916_), .B(new_n2602_), .ZN(new_n4917_));
  NOR2_X1    g02482(.A1(new_n2635_), .A2(new_n4886_), .ZN(new_n4918_));
  NOR2_X1    g02483(.A1(new_n2634_), .A2(new_n4888_), .ZN(new_n4919_));
  OAI21_X1   g02484(.A1(new_n4918_), .A2(new_n4919_), .B(pi0222), .ZN(new_n4920_));
  AOI21_X1   g02485(.A1(new_n4891_), .A2(pi0224), .B(pi0222), .ZN(new_n4921_));
  NAND3_X1   g02486(.A1(new_n3028_), .A2(new_n2631_), .A3(new_n4893_), .ZN(new_n4922_));
  AND2_X2    g02487(.A1(new_n4922_), .A2(new_n4921_), .Z(new_n4923_));
  INV_X1     g02488(.I(new_n4923_), .ZN(new_n4924_));
  NAND2_X1   g02489(.A1(new_n4924_), .A2(new_n4920_), .ZN(new_n4925_));
  NAND2_X1   g02490(.A1(new_n4925_), .A2(new_n2668_), .ZN(new_n4926_));
  NAND2_X1   g02491(.A1(pi0223), .A2(pi1135), .ZN(new_n4927_));
  AOI21_X1   g02492(.A1(new_n4926_), .A2(new_n4927_), .B(pi0299), .ZN(new_n4928_));
  AOI21_X1   g02493(.A1(new_n4915_), .A2(pi0299), .B(new_n4928_), .ZN(new_n4929_));
  INV_X1     g02494(.I(new_n4929_), .ZN(new_n4930_));
  OAI21_X1   g02495(.A1(new_n4930_), .A2(new_n2562_), .B(new_n2602_), .ZN(new_n4931_));
  AOI21_X1   g02496(.A1(new_n4769_), .A2(new_n4898_), .B(pi0216), .ZN(new_n4932_));
  NAND2_X1   g02497(.A1(new_n3404_), .A2(pi0161), .ZN(new_n4933_));
  NAND2_X1   g02498(.A1(new_n3387_), .A2(new_n3360_), .ZN(new_n4934_));
  AOI21_X1   g02499(.A1(new_n4933_), .A2(new_n4934_), .B(pi0879), .ZN(new_n4935_));
  OAI21_X1   g02500(.A1(new_n3451_), .A2(pi0161), .B(pi0879), .ZN(new_n4936_));
  NAND2_X1   g02501(.A1(new_n4936_), .A2(new_n2458_), .ZN(new_n4937_));
  OAI21_X1   g02502(.A1(new_n4935_), .A2(new_n4937_), .B(new_n4932_), .ZN(new_n4938_));
  AOI21_X1   g02503(.A1(new_n4938_), .A2(new_n4908_), .B(pi0221), .ZN(new_n4939_));
  NOR3_X1    g02504(.A1(new_n4939_), .A2(pi0215), .A3(new_n4907_), .ZN(new_n4940_));
  OAI21_X1   g02505(.A1(new_n4940_), .A2(new_n4884_), .B(pi0299), .ZN(new_n4941_));
  NAND2_X1   g02506(.A1(new_n4927_), .A2(new_n2628_), .ZN(new_n4942_));
  INV_X1     g02507(.I(new_n4942_), .ZN(new_n4943_));
  OAI21_X1   g02508(.A1(new_n4782_), .A2(new_n4925_), .B(new_n2668_), .ZN(new_n4944_));
  AOI21_X1   g02509(.A1(new_n4944_), .A2(new_n4943_), .B(pi0039), .ZN(new_n4945_));
  AOI21_X1   g02510(.A1(new_n4905_), .A2(pi0299), .B(new_n4928_), .ZN(new_n4946_));
  INV_X1     g02511(.I(new_n4946_), .ZN(new_n4947_));
  AOI22_X1   g02512(.A1(new_n4941_), .A2(new_n4945_), .B1(pi0039), .B2(new_n4947_), .ZN(new_n4948_));
  OAI21_X1   g02513(.A1(new_n4930_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n4949_));
  AOI21_X1   g02514(.A1(new_n4948_), .A2(new_n3265_), .B(new_n4949_), .ZN(new_n4950_));
  INV_X1     g02515(.I(new_n4928_), .ZN(new_n4951_));
  OAI21_X1   g02516(.A1(new_n4930_), .A2(new_n2572_), .B(pi0100), .ZN(new_n4952_));
  NOR3_X1    g02517(.A1(new_n3363_), .A2(pi0152), .A3(pi0166), .ZN(new_n4953_));
  AOI21_X1   g02518(.A1(new_n3369_), .A2(new_n3361_), .B(new_n3366_), .ZN(new_n4954_));
  OAI21_X1   g02519(.A1(new_n4954_), .A2(new_n4953_), .B(pi0879), .ZN(new_n4955_));
  OAI21_X1   g02520(.A1(new_n3366_), .A2(pi0879), .B(pi0161), .ZN(new_n4956_));
  AOI21_X1   g02521(.A1(new_n4955_), .A2(new_n4956_), .B(pi0228), .ZN(new_n4957_));
  OR2_X2     g02522(.A1(new_n4957_), .A2(new_n4899_), .Z(new_n4958_));
  OAI21_X1   g02523(.A1(new_n4958_), .A2(new_n3302_), .B(new_n2614_), .ZN(new_n4959_));
  NAND2_X1   g02524(.A1(new_n4959_), .A2(new_n4908_), .ZN(new_n4960_));
  AOI21_X1   g02525(.A1(new_n4960_), .A2(new_n2441_), .B(pi0215), .ZN(new_n4961_));
  AOI21_X1   g02526(.A1(new_n4961_), .A2(new_n4890_), .B(new_n4884_), .ZN(new_n4962_));
  AOI21_X1   g02527(.A1(new_n4962_), .A2(pi0299), .B(new_n2573_), .ZN(new_n4963_));
  AOI21_X1   g02528(.A1(new_n4963_), .A2(new_n4951_), .B(new_n4952_), .ZN(new_n4964_));
  NOR3_X1    g02529(.A1(new_n4950_), .A2(pi0087), .A3(new_n4964_), .ZN(new_n4965_));
  NAND2_X1   g02530(.A1(new_n4930_), .A2(new_n3273_), .ZN(new_n4966_));
  OAI21_X1   g02531(.A1(new_n4946_), .A2(new_n3273_), .B(new_n4966_), .ZN(new_n4967_));
  NOR2_X1    g02532(.A1(new_n4967_), .A2(new_n3458_), .ZN(new_n4968_));
  OAI21_X1   g02533(.A1(new_n4965_), .A2(new_n4968_), .B(new_n3465_), .ZN(new_n4969_));
  AOI21_X1   g02534(.A1(new_n4929_), .A2(pi0075), .B(pi0092), .ZN(new_n4970_));
  NAND2_X1   g02535(.A1(new_n4967_), .A2(new_n2564_), .ZN(new_n4971_));
  OAI21_X1   g02536(.A1(new_n2564_), .A2(new_n4929_), .B(new_n4971_), .ZN(new_n4972_));
  AOI22_X1   g02537(.A1(new_n4969_), .A2(new_n4970_), .B1(pi0092), .B2(new_n4972_), .ZN(new_n4973_));
  AOI21_X1   g02538(.A1(new_n4973_), .A2(new_n2562_), .B(new_n4931_), .ZN(new_n4974_));
  NOR3_X1    g02539(.A1(new_n4974_), .A2(pi0056), .A3(new_n4917_), .ZN(new_n4975_));
  NAND2_X1   g02540(.A1(new_n4904_), .A2(new_n2576_), .ZN(new_n4976_));
  NAND2_X1   g02541(.A1(new_n4914_), .A2(new_n2577_), .ZN(new_n4977_));
  AOI21_X1   g02542(.A1(new_n4976_), .A2(new_n4977_), .B(new_n3284_), .ZN(new_n4978_));
  NOR3_X1    g02543(.A1(new_n4975_), .A2(pi0062), .A3(new_n4978_), .ZN(new_n4979_));
  NAND2_X1   g02544(.A1(new_n4905_), .A2(new_n3320_), .ZN(new_n4980_));
  NAND2_X1   g02545(.A1(new_n4915_), .A2(new_n3472_), .ZN(new_n4981_));
  AOI21_X1   g02546(.A1(new_n4980_), .A2(new_n4981_), .B(new_n3471_), .ZN(new_n4982_));
  NOR3_X1    g02547(.A1(new_n4979_), .A2(new_n3425_), .A3(new_n4982_), .ZN(new_n4983_));
  OAI21_X1   g02548(.A1(new_n4915_), .A2(new_n3291_), .B(pi0244), .ZN(new_n4984_));
  NOR2_X1    g02549(.A1(new_n2614_), .A2(pi0279), .ZN(new_n4985_));
  AOI21_X1   g02550(.A1(new_n4900_), .A2(new_n2614_), .B(new_n4985_), .ZN(new_n4986_));
  NAND2_X1   g02551(.A1(new_n4986_), .A2(new_n2441_), .ZN(new_n4987_));
  AND3_X2    g02552(.A1(new_n4987_), .A2(new_n2436_), .A3(new_n4890_), .Z(new_n4988_));
  NOR2_X1    g02553(.A1(new_n4988_), .A2(new_n4884_), .ZN(new_n4989_));
  INV_X1     g02554(.I(new_n4913_), .ZN(new_n4990_));
  NOR2_X1    g02555(.A1(new_n4990_), .A2(new_n3320_), .ZN(new_n4991_));
  AOI21_X1   g02556(.A1(new_n4989_), .A2(new_n3320_), .B(new_n4991_), .ZN(new_n4992_));
  OAI21_X1   g02557(.A1(new_n4992_), .A2(new_n3471_), .B(new_n3291_), .ZN(new_n4993_));
  NOR3_X1    g02558(.A1(new_n4988_), .A2(new_n2612_), .A3(new_n4884_), .ZN(new_n4994_));
  NOR2_X1    g02559(.A1(new_n4990_), .A2(new_n2611_), .ZN(new_n4995_));
  OAI21_X1   g02560(.A1(new_n4994_), .A2(new_n4995_), .B(pi0055), .ZN(new_n4996_));
  OAI21_X1   g02561(.A1(new_n2644_), .A2(new_n4897_), .B(new_n4928_), .ZN(new_n4997_));
  INV_X1     g02562(.I(new_n4997_), .ZN(new_n4998_));
  AOI21_X1   g02563(.A1(pi0299), .A2(new_n4913_), .B(new_n4998_), .ZN(new_n4999_));
  AOI21_X1   g02564(.A1(new_n4999_), .A2(new_n2563_), .B(pi0055), .ZN(new_n5000_));
  INV_X1     g02565(.I(new_n4769_), .ZN(new_n5001_));
  INV_X1     g02566(.I(new_n4932_), .ZN(new_n5002_));
  NAND2_X1   g02567(.A1(new_n3731_), .A2(pi0161), .ZN(new_n5003_));
  NAND2_X1   g02568(.A1(new_n3403_), .A2(new_n3360_), .ZN(new_n5004_));
  AOI21_X1   g02569(.A1(new_n5004_), .A2(new_n5003_), .B(new_n4893_), .ZN(new_n5005_));
  NOR3_X1    g02570(.A1(new_n3451_), .A2(new_n3360_), .A3(pi0879), .ZN(new_n5006_));
  OAI21_X1   g02571(.A1(new_n5005_), .A2(new_n5006_), .B(new_n2458_), .ZN(new_n5007_));
  AOI21_X1   g02572(.A1(new_n5007_), .A2(new_n5001_), .B(new_n5002_), .ZN(new_n5008_));
  OAI21_X1   g02573(.A1(new_n5008_), .A2(new_n4892_), .B(new_n2441_), .ZN(new_n5009_));
  NAND3_X1   g02574(.A1(new_n5009_), .A2(new_n2436_), .A3(new_n4890_), .ZN(new_n5010_));
  AOI21_X1   g02575(.A1(new_n5010_), .A2(new_n4885_), .B(new_n2628_), .ZN(new_n5011_));
  NAND2_X1   g02576(.A1(new_n4849_), .A2(new_n4923_), .ZN(new_n5012_));
  AOI21_X1   g02577(.A1(new_n5012_), .A2(new_n4920_), .B(pi0223), .ZN(new_n5013_));
  OAI21_X1   g02578(.A1(new_n5013_), .A2(new_n4942_), .B(new_n2627_), .ZN(new_n5014_));
  AOI21_X1   g02579(.A1(new_n4989_), .A2(pi0299), .B(new_n4998_), .ZN(new_n5015_));
  OAI22_X1   g02580(.A1(new_n5011_), .A2(new_n5014_), .B1(new_n2627_), .B2(new_n5015_), .ZN(new_n5016_));
  AOI21_X1   g02581(.A1(new_n4999_), .A2(pi0038), .B(pi0100), .ZN(new_n5017_));
  OAI21_X1   g02582(.A1(new_n5016_), .A2(pi0038), .B(new_n5017_), .ZN(new_n5018_));
  AOI21_X1   g02583(.A1(new_n4999_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n5019_));
  NAND2_X1   g02584(.A1(new_n4885_), .A2(pi0299), .ZN(new_n5020_));
  NOR2_X1    g02585(.A1(new_n4958_), .A2(pi0216), .ZN(new_n5021_));
  NOR3_X1    g02586(.A1(new_n5021_), .A2(pi0221), .A3(new_n4985_), .ZN(new_n5022_));
  NOR3_X1    g02587(.A1(new_n5022_), .A2(pi0215), .A3(new_n4907_), .ZN(new_n5023_));
  OAI21_X1   g02588(.A1(new_n5023_), .A2(new_n5020_), .B(new_n4997_), .ZN(new_n5024_));
  OAI21_X1   g02589(.A1(new_n5024_), .A2(new_n2573_), .B(new_n5019_), .ZN(new_n5025_));
  NAND3_X1   g02590(.A1(new_n5018_), .A2(new_n3458_), .A3(new_n5025_), .ZN(new_n5026_));
  INV_X1     g02591(.I(new_n4999_), .ZN(new_n5027_));
  NOR2_X1    g02592(.A1(new_n5015_), .A2(new_n3273_), .ZN(new_n5028_));
  AOI21_X1   g02593(.A1(new_n3273_), .A2(new_n5027_), .B(new_n5028_), .ZN(new_n5029_));
  NAND2_X1   g02594(.A1(new_n5029_), .A2(pi0087), .ZN(new_n5030_));
  AOI21_X1   g02595(.A1(new_n5026_), .A2(new_n5030_), .B(pi0075), .ZN(new_n5031_));
  OAI21_X1   g02596(.A1(new_n5027_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n5032_));
  NOR2_X1    g02597(.A1(new_n5029_), .A2(new_n2565_), .ZN(new_n5033_));
  AOI21_X1   g02598(.A1(new_n2565_), .A2(new_n5027_), .B(new_n5033_), .ZN(new_n5034_));
  OAI22_X1   g02599(.A1(new_n5031_), .A2(new_n5032_), .B1(new_n3444_), .B2(new_n5034_), .ZN(new_n5035_));
  OAI21_X1   g02600(.A1(new_n5035_), .A2(new_n2563_), .B(new_n5000_), .ZN(new_n5036_));
  NAND3_X1   g02601(.A1(new_n5036_), .A2(new_n3284_), .A3(new_n4996_), .ZN(new_n5037_));
  NAND2_X1   g02602(.A1(new_n4990_), .A2(new_n2577_), .ZN(new_n5038_));
  OAI21_X1   g02603(.A1(new_n4989_), .A2(new_n2577_), .B(new_n5038_), .ZN(new_n5039_));
  AOI21_X1   g02604(.A1(new_n5039_), .A2(pi0056), .B(pi0062), .ZN(new_n5040_));
  AOI21_X1   g02605(.A1(new_n5037_), .A2(new_n5040_), .B(new_n4993_), .ZN(new_n5041_));
  INV_X1     g02606(.I(pi0244), .ZN(new_n5042_));
  OAI21_X1   g02607(.A1(new_n4913_), .A2(new_n3291_), .B(new_n5042_), .ZN(new_n5043_));
  OAI22_X1   g02608(.A1(new_n4983_), .A2(new_n4984_), .B1(new_n5041_), .B2(new_n5043_), .ZN(po0164));
  INV_X1     g02609(.I(pi1134), .ZN(new_n5045_));
  AOI21_X1   g02610(.A1(pi0216), .A2(pi0278), .B(pi0221), .ZN(new_n5046_));
  INV_X1     g02611(.I(pi0846), .ZN(new_n5047_));
  NOR2_X1    g02612(.A1(new_n2463_), .A2(new_n5047_), .ZN(new_n5048_));
  NOR2_X1    g02613(.A1(new_n3369_), .A2(pi0105), .ZN(new_n5049_));
  AOI21_X1   g02614(.A1(new_n5048_), .A2(pi0105), .B(new_n5049_), .ZN(new_n5050_));
  NOR2_X1    g02615(.A1(new_n5050_), .A2(new_n2458_), .ZN(new_n5051_));
  NOR2_X1    g02616(.A1(new_n3369_), .A2(pi0228), .ZN(new_n5052_));
  OAI21_X1   g02617(.A1(new_n5051_), .A2(new_n5052_), .B(new_n2614_), .ZN(new_n5053_));
  NAND2_X1   g02618(.A1(new_n5053_), .A2(new_n5046_), .ZN(new_n5054_));
  INV_X1     g02619(.I(pi0930), .ZN(new_n5055_));
  NOR2_X1    g02620(.A1(new_n2441_), .A2(pi0216), .ZN(new_n5056_));
  NAND3_X1   g02621(.A1(new_n5056_), .A2(pi0833), .A3(new_n5055_), .ZN(new_n5057_));
  AOI21_X1   g02622(.A1(new_n5054_), .A2(new_n5057_), .B(pi0215), .ZN(new_n5058_));
  AOI21_X1   g02623(.A1(new_n5058_), .A2(new_n3425_), .B(pi0242), .ZN(new_n5059_));
  INV_X1     g02624(.I(new_n5057_), .ZN(new_n5060_));
  INV_X1     g02625(.I(new_n5046_), .ZN(new_n5061_));
  NAND2_X1   g02626(.A1(new_n2531_), .A2(pi0846), .ZN(new_n5062_));
  NAND2_X1   g02627(.A1(new_n2530_), .A2(pi0152), .ZN(new_n5063_));
  AOI21_X1   g02628(.A1(new_n5062_), .A2(new_n5063_), .B(pi0228), .ZN(new_n5064_));
  NOR2_X1    g02629(.A1(new_n5064_), .A2(new_n5051_), .ZN(new_n5065_));
  NOR2_X1    g02630(.A1(new_n5065_), .A2(pi0216), .ZN(new_n5066_));
  NOR2_X1    g02631(.A1(new_n5066_), .A2(new_n5061_), .ZN(new_n5067_));
  OAI21_X1   g02632(.A1(new_n5067_), .A2(new_n5060_), .B(new_n2436_), .ZN(new_n5068_));
  NAND2_X1   g02633(.A1(new_n5068_), .A2(new_n3320_), .ZN(new_n5069_));
  INV_X1     g02634(.I(new_n5058_), .ZN(new_n5070_));
  NAND2_X1   g02635(.A1(new_n3472_), .A2(new_n5070_), .ZN(new_n5071_));
  AOI21_X1   g02636(.A1(new_n5069_), .A2(new_n5071_), .B(new_n3471_), .ZN(new_n5072_));
  NAND2_X1   g02637(.A1(new_n5068_), .A2(new_n2611_), .ZN(new_n5073_));
  NAND2_X1   g02638(.A1(new_n5070_), .A2(new_n2612_), .ZN(new_n5074_));
  AOI21_X1   g02639(.A1(new_n5073_), .A2(new_n5074_), .B(new_n2602_), .ZN(new_n5075_));
  AOI21_X1   g02640(.A1(pi0224), .A2(pi0278), .B(pi0222), .ZN(new_n5076_));
  INV_X1     g02641(.I(new_n5076_), .ZN(new_n5077_));
  NAND2_X1   g02642(.A1(new_n5048_), .A2(new_n2631_), .ZN(new_n5078_));
  INV_X1     g02643(.I(new_n5078_), .ZN(new_n5079_));
  NOR2_X1    g02644(.A1(new_n5079_), .A2(new_n5077_), .ZN(new_n5080_));
  NOR2_X1    g02645(.A1(new_n2629_), .A2(pi0224), .ZN(new_n5081_));
  INV_X1     g02646(.I(new_n5081_), .ZN(new_n5082_));
  NOR3_X1    g02647(.A1(new_n5082_), .A2(new_n2443_), .A3(pi0930), .ZN(new_n5083_));
  INV_X1     g02648(.I(new_n5083_), .ZN(new_n5084_));
  INV_X1     g02649(.I(new_n5080_), .ZN(new_n5085_));
  NAND3_X1   g02650(.A1(new_n5085_), .A2(new_n2639_), .A3(new_n5084_), .ZN(new_n5086_));
  NAND2_X1   g02651(.A1(new_n5086_), .A2(new_n2628_), .ZN(new_n5087_));
  NOR2_X1    g02652(.A1(new_n5087_), .A2(new_n3653_), .ZN(new_n5088_));
  AOI21_X1   g02653(.A1(new_n5088_), .A2(new_n2639_), .B(pi0299), .ZN(new_n5089_));
  INV_X1     g02654(.I(new_n5089_), .ZN(new_n5090_));
  AOI21_X1   g02655(.A1(new_n2668_), .A2(new_n5080_), .B(new_n5090_), .ZN(new_n5091_));
  AOI21_X1   g02656(.A1(pi0299), .A2(new_n5070_), .B(new_n5091_), .ZN(new_n5092_));
  INV_X1     g02657(.I(new_n5092_), .ZN(new_n5093_));
  OAI21_X1   g02658(.A1(new_n5093_), .A2(new_n2562_), .B(new_n2602_), .ZN(new_n5094_));
  AOI21_X1   g02659(.A1(new_n5068_), .A2(pi0299), .B(new_n5091_), .ZN(new_n5095_));
  OAI21_X1   g02660(.A1(new_n5095_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n5096_));
  OAI21_X1   g02661(.A1(new_n3392_), .A2(pi0846), .B(new_n2631_), .ZN(new_n5097_));
  AOI21_X1   g02662(.A1(new_n5097_), .A2(new_n5076_), .B(new_n5083_), .ZN(new_n5098_));
  OAI21_X1   g02663(.A1(new_n5098_), .A2(new_n3336_), .B(new_n2627_), .ZN(new_n5099_));
  AOI21_X1   g02664(.A1(new_n3812_), .A2(new_n5079_), .B(new_n5077_), .ZN(new_n5100_));
  AOI21_X1   g02665(.A1(new_n3335_), .A2(new_n5100_), .B(new_n5099_), .ZN(new_n5101_));
  OAI21_X1   g02666(.A1(new_n3369_), .A2(pi0105), .B(pi0228), .ZN(new_n5102_));
  NOR2_X1    g02667(.A1(new_n3381_), .A2(new_n5102_), .ZN(new_n5103_));
  AOI21_X1   g02668(.A1(new_n3381_), .A2(new_n5047_), .B(new_n2457_), .ZN(new_n5104_));
  OAI21_X1   g02669(.A1(new_n5104_), .A2(new_n5102_), .B(new_n2614_), .ZN(new_n5105_));
  NAND2_X1   g02670(.A1(new_n5047_), .A2(pi0152), .ZN(new_n5106_));
  OAI21_X1   g02671(.A1(new_n3451_), .A2(new_n5106_), .B(new_n2458_), .ZN(new_n5107_));
  NAND2_X1   g02672(.A1(new_n3731_), .A2(pi0152), .ZN(new_n5108_));
  OAI21_X1   g02673(.A1(new_n3404_), .A2(pi0152), .B(new_n5108_), .ZN(new_n5109_));
  AOI21_X1   g02674(.A1(new_n5109_), .A2(pi0846), .B(new_n5107_), .ZN(new_n5110_));
  NOR3_X1    g02675(.A1(new_n5110_), .A2(new_n5103_), .A3(new_n5105_), .ZN(new_n5111_));
  OAI21_X1   g02676(.A1(new_n5111_), .A2(new_n5061_), .B(new_n5057_), .ZN(new_n5112_));
  NOR2_X1    g02677(.A1(new_n2628_), .A2(pi0215), .ZN(new_n5113_));
  NAND2_X1   g02678(.A1(new_n5112_), .A2(new_n5113_), .ZN(new_n5114_));
  AOI21_X1   g02679(.A1(new_n5114_), .A2(new_n5101_), .B(new_n5096_), .ZN(new_n5115_));
  OAI21_X1   g02680(.A1(new_n5093_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n5116_));
  OAI21_X1   g02681(.A1(new_n5093_), .A2(new_n2572_), .B(pi0100), .ZN(new_n5117_));
  OAI22_X1   g02682(.A1(new_n3368_), .A2(new_n5047_), .B1(new_n3369_), .B2(new_n3365_), .ZN(new_n5118_));
  NAND2_X1   g02683(.A1(new_n5118_), .A2(new_n2458_), .ZN(new_n5119_));
  INV_X1     g02684(.I(new_n5119_), .ZN(new_n5120_));
  OAI21_X1   g02685(.A1(new_n5120_), .A2(new_n5051_), .B(new_n2614_), .ZN(new_n5121_));
  NAND2_X1   g02686(.A1(new_n5121_), .A2(new_n5046_), .ZN(new_n5122_));
  AOI21_X1   g02687(.A1(new_n5122_), .A2(new_n5057_), .B(pi0215), .ZN(new_n5123_));
  NOR2_X1    g02688(.A1(new_n5123_), .A2(new_n2628_), .ZN(new_n5124_));
  NOR3_X1    g02689(.A1(new_n5124_), .A2(new_n2573_), .A3(new_n5091_), .ZN(new_n5125_));
  OAI22_X1   g02690(.A1(new_n5115_), .A2(new_n5116_), .B1(new_n5117_), .B2(new_n5125_), .ZN(new_n5126_));
  NOR2_X1    g02691(.A1(new_n5095_), .A2(new_n3273_), .ZN(new_n5127_));
  AOI21_X1   g02692(.A1(new_n3273_), .A2(new_n5093_), .B(new_n5127_), .ZN(new_n5128_));
  NAND2_X1   g02693(.A1(new_n5128_), .A2(pi0087), .ZN(new_n5129_));
  OAI21_X1   g02694(.A1(new_n5126_), .A2(pi0087), .B(new_n5129_), .ZN(new_n5130_));
  OAI21_X1   g02695(.A1(new_n5093_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n5131_));
  AOI21_X1   g02696(.A1(new_n5130_), .A2(new_n3465_), .B(new_n5131_), .ZN(new_n5132_));
  NAND2_X1   g02697(.A1(new_n5093_), .A2(new_n2565_), .ZN(new_n5133_));
  OR2_X2     g02698(.A1(new_n5128_), .A2(new_n2565_), .Z(new_n5134_));
  AOI21_X1   g02699(.A1(new_n5134_), .A2(new_n5133_), .B(new_n3444_), .ZN(new_n5135_));
  NOR3_X1    g02700(.A1(new_n5132_), .A2(new_n2563_), .A3(new_n5135_), .ZN(new_n5136_));
  OAI21_X1   g02701(.A1(new_n5136_), .A2(new_n5094_), .B(new_n3284_), .ZN(new_n5137_));
  NOR2_X1    g02702(.A1(new_n5068_), .A2(new_n2577_), .ZN(new_n5138_));
  AOI21_X1   g02703(.A1(new_n2577_), .A2(new_n5058_), .B(new_n5138_), .ZN(new_n5139_));
  OAI22_X1   g02704(.A1(new_n5137_), .A2(new_n5075_), .B1(new_n3284_), .B2(new_n5139_), .ZN(new_n5140_));
  OAI21_X1   g02705(.A1(new_n5140_), .A2(pi0062), .B(new_n3291_), .ZN(new_n5141_));
  OAI21_X1   g02706(.A1(new_n5141_), .A2(new_n5072_), .B(new_n5059_), .ZN(new_n5142_));
  INV_X1     g02707(.I(pi0242), .ZN(new_n5143_));
  NOR2_X1    g02708(.A1(new_n5070_), .A2(new_n3307_), .ZN(new_n5144_));
  AOI21_X1   g02709(.A1(new_n5144_), .A2(new_n3425_), .B(new_n5143_), .ZN(new_n5145_));
  INV_X1     g02710(.I(new_n5064_), .ZN(new_n5146_));
  NOR2_X1    g02711(.A1(new_n5051_), .A2(new_n3302_), .ZN(new_n5147_));
  AOI21_X1   g02712(.A1(new_n5146_), .A2(new_n5147_), .B(pi0216), .ZN(new_n5148_));
  NOR2_X1    g02713(.A1(new_n5148_), .A2(new_n5061_), .ZN(new_n5149_));
  INV_X1     g02714(.I(new_n5149_), .ZN(new_n5150_));
  AOI21_X1   g02715(.A1(new_n5150_), .A2(new_n5057_), .B(pi0215), .ZN(new_n5151_));
  NOR2_X1    g02716(.A1(new_n5151_), .A2(new_n2612_), .ZN(new_n5152_));
  NOR2_X1    g02717(.A1(new_n5144_), .A2(new_n2611_), .ZN(new_n5153_));
  OAI21_X1   g02718(.A1(new_n5152_), .A2(new_n5153_), .B(pi0055), .ZN(new_n5154_));
  INV_X1     g02719(.I(new_n5144_), .ZN(new_n5155_));
  AOI21_X1   g02720(.A1(new_n5155_), .A2(pi0299), .B(new_n5089_), .ZN(new_n5156_));
  AOI21_X1   g02721(.A1(new_n5156_), .A2(new_n2563_), .B(pi0055), .ZN(new_n5157_));
  INV_X1     g02722(.I(new_n5151_), .ZN(new_n5158_));
  AOI21_X1   g02723(.A1(new_n5158_), .A2(pi0299), .B(new_n5089_), .ZN(new_n5159_));
  OAI21_X1   g02724(.A1(new_n5159_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n5160_));
  NOR2_X1    g02725(.A1(new_n3387_), .A2(pi0152), .ZN(new_n5161_));
  NOR2_X1    g02726(.A1(new_n3404_), .A2(new_n3369_), .ZN(new_n5162_));
  OAI21_X1   g02727(.A1(new_n5162_), .A2(new_n5161_), .B(new_n5047_), .ZN(new_n5163_));
  NAND3_X1   g02728(.A1(new_n3657_), .A2(new_n3369_), .A3(pi0846), .ZN(new_n5164_));
  AOI21_X1   g02729(.A1(new_n5163_), .A2(new_n5164_), .B(pi0228), .ZN(new_n5165_));
  OAI21_X1   g02730(.A1(new_n5165_), .A2(new_n5105_), .B(new_n5046_), .ZN(new_n5166_));
  NAND2_X1   g02731(.A1(new_n5166_), .A2(new_n5057_), .ZN(new_n5167_));
  AOI21_X1   g02732(.A1(new_n5167_), .A2(new_n5113_), .B(new_n5099_), .ZN(new_n5168_));
  AOI21_X1   g02733(.A1(new_n5156_), .A2(pi0038), .B(pi0100), .ZN(new_n5169_));
  OAI21_X1   g02734(.A1(new_n5168_), .A2(new_n5160_), .B(new_n5169_), .ZN(new_n5170_));
  AOI21_X1   g02735(.A1(new_n5156_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n5171_));
  NAND2_X1   g02736(.A1(new_n5119_), .A2(new_n5147_), .ZN(new_n5172_));
  AOI21_X1   g02737(.A1(new_n5172_), .A2(new_n2614_), .B(new_n5061_), .ZN(new_n5173_));
  NOR2_X1    g02738(.A1(new_n5173_), .A2(new_n5060_), .ZN(new_n5174_));
  OAI21_X1   g02739(.A1(new_n5174_), .A2(pi0215), .B(pi0299), .ZN(new_n5175_));
  NAND3_X1   g02740(.A1(new_n5175_), .A2(new_n2572_), .A3(new_n5090_), .ZN(new_n5176_));
  NAND2_X1   g02741(.A1(new_n5176_), .A2(new_n5171_), .ZN(new_n5177_));
  NAND3_X1   g02742(.A1(new_n5170_), .A2(new_n3458_), .A3(new_n5177_), .ZN(new_n5178_));
  INV_X1     g02743(.I(new_n5156_), .ZN(new_n5179_));
  NOR2_X1    g02744(.A1(new_n5159_), .A2(new_n3273_), .ZN(new_n5180_));
  AOI21_X1   g02745(.A1(new_n3273_), .A2(new_n5179_), .B(new_n5180_), .ZN(new_n5181_));
  NAND2_X1   g02746(.A1(new_n5181_), .A2(pi0087), .ZN(new_n5182_));
  AOI21_X1   g02747(.A1(new_n5178_), .A2(new_n5182_), .B(pi0075), .ZN(new_n5183_));
  OAI21_X1   g02748(.A1(new_n5179_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n5184_));
  NOR2_X1    g02749(.A1(new_n5181_), .A2(new_n2565_), .ZN(new_n5185_));
  AOI21_X1   g02750(.A1(new_n2565_), .A2(new_n5179_), .B(new_n5185_), .ZN(new_n5186_));
  OAI22_X1   g02751(.A1(new_n5183_), .A2(new_n5184_), .B1(new_n3444_), .B2(new_n5186_), .ZN(new_n5187_));
  OAI21_X1   g02752(.A1(new_n5187_), .A2(new_n2563_), .B(new_n5157_), .ZN(new_n5188_));
  NAND3_X1   g02753(.A1(new_n5188_), .A2(new_n3284_), .A3(new_n5154_), .ZN(new_n5189_));
  NOR2_X1    g02754(.A1(new_n5158_), .A2(new_n2577_), .ZN(new_n5190_));
  NOR2_X1    g02755(.A1(new_n5155_), .A2(new_n2576_), .ZN(new_n5191_));
  OAI21_X1   g02756(.A1(new_n5190_), .A2(new_n5191_), .B(pi0056), .ZN(new_n5192_));
  NAND3_X1   g02757(.A1(new_n5189_), .A2(new_n3471_), .A3(new_n5192_), .ZN(new_n5193_));
  NOR2_X1    g02758(.A1(new_n5151_), .A2(new_n3472_), .ZN(new_n5194_));
  NOR2_X1    g02759(.A1(new_n3320_), .A2(new_n5144_), .ZN(new_n5195_));
  OAI21_X1   g02760(.A1(new_n5194_), .A2(new_n5195_), .B(pi0062), .ZN(new_n5196_));
  NAND3_X1   g02761(.A1(new_n5193_), .A2(new_n3291_), .A3(new_n5196_), .ZN(new_n5197_));
  AOI21_X1   g02762(.A1(new_n5197_), .A2(new_n5145_), .B(new_n5045_), .ZN(new_n5198_));
  NAND2_X1   g02763(.A1(new_n2447_), .A2(pi0221), .ZN(new_n5199_));
  NAND2_X1   g02764(.A1(new_n5199_), .A2(new_n2436_), .ZN(new_n5200_));
  NOR2_X1    g02765(.A1(new_n5200_), .A2(new_n5060_), .ZN(new_n5201_));
  INV_X1     g02766(.I(new_n5201_), .ZN(new_n5202_));
  NOR2_X1    g02767(.A1(new_n5067_), .A2(new_n5202_), .ZN(new_n5203_));
  INV_X1     g02768(.I(new_n5203_), .ZN(new_n5204_));
  NAND2_X1   g02769(.A1(new_n5204_), .A2(new_n2611_), .ZN(new_n5205_));
  NAND2_X1   g02770(.A1(new_n5054_), .A2(new_n5201_), .ZN(new_n5206_));
  NAND2_X1   g02771(.A1(new_n5206_), .A2(new_n2612_), .ZN(new_n5207_));
  AOI21_X1   g02772(.A1(new_n5205_), .A2(new_n5207_), .B(new_n2602_), .ZN(new_n5208_));
  INV_X1     g02773(.I(new_n5087_), .ZN(new_n5209_));
  AOI21_X1   g02774(.A1(new_n5206_), .A2(pi0299), .B(new_n5209_), .ZN(new_n5210_));
  INV_X1     g02775(.I(new_n5210_), .ZN(new_n5211_));
  OAI21_X1   g02776(.A1(new_n5211_), .A2(new_n2562_), .B(new_n2602_), .ZN(new_n5212_));
  AOI21_X1   g02777(.A1(new_n5204_), .A2(pi0299), .B(new_n5209_), .ZN(new_n5213_));
  NOR2_X1    g02778(.A1(new_n5213_), .A2(new_n2627_), .ZN(new_n5214_));
  NOR2_X1    g02779(.A1(new_n5214_), .A2(pi0038), .ZN(new_n5215_));
  NOR2_X1    g02780(.A1(new_n2638_), .A2(new_n3336_), .ZN(new_n5216_));
  INV_X1     g02781(.I(new_n5216_), .ZN(new_n5217_));
  NOR2_X1    g02782(.A1(new_n5100_), .A2(new_n5217_), .ZN(new_n5218_));
  AOI21_X1   g02783(.A1(new_n5218_), .A2(new_n5084_), .B(pi0039), .ZN(new_n5219_));
  NAND2_X1   g02784(.A1(new_n5199_), .A2(new_n5113_), .ZN(new_n5220_));
  OAI21_X1   g02785(.A1(new_n5112_), .A2(new_n5220_), .B(new_n5219_), .ZN(new_n5221_));
  OAI21_X1   g02786(.A1(new_n5211_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n5222_));
  AOI21_X1   g02787(.A1(new_n5221_), .A2(new_n5215_), .B(new_n5222_), .ZN(new_n5223_));
  OAI21_X1   g02788(.A1(new_n5211_), .A2(new_n2572_), .B(pi0100), .ZN(new_n5224_));
  NAND2_X1   g02789(.A1(new_n5122_), .A2(new_n5201_), .ZN(new_n5225_));
  AOI21_X1   g02790(.A1(new_n5225_), .A2(pi0299), .B(new_n5209_), .ZN(new_n5226_));
  AOI21_X1   g02791(.A1(new_n5226_), .A2(new_n2572_), .B(new_n5224_), .ZN(new_n5227_));
  NOR3_X1    g02792(.A1(new_n5223_), .A2(pi0087), .A3(new_n5227_), .ZN(new_n5228_));
  NAND2_X1   g02793(.A1(new_n5211_), .A2(new_n3273_), .ZN(new_n5229_));
  OAI21_X1   g02794(.A1(new_n5213_), .A2(new_n3273_), .B(new_n5229_), .ZN(new_n5230_));
  NOR2_X1    g02795(.A1(new_n5230_), .A2(new_n3458_), .ZN(new_n5231_));
  OAI21_X1   g02796(.A1(new_n5228_), .A2(new_n5231_), .B(new_n3465_), .ZN(new_n5232_));
  AOI21_X1   g02797(.A1(new_n5210_), .A2(pi0075), .B(pi0092), .ZN(new_n5233_));
  NAND2_X1   g02798(.A1(new_n5230_), .A2(new_n2564_), .ZN(new_n5234_));
  OAI21_X1   g02799(.A1(new_n2564_), .A2(new_n5210_), .B(new_n5234_), .ZN(new_n5235_));
  AOI22_X1   g02800(.A1(new_n5232_), .A2(new_n5233_), .B1(pi0092), .B2(new_n5235_), .ZN(new_n5236_));
  AOI21_X1   g02801(.A1(new_n5236_), .A2(new_n2562_), .B(new_n5212_), .ZN(new_n5237_));
  NOR3_X1    g02802(.A1(new_n5237_), .A2(pi0056), .A3(new_n5208_), .ZN(new_n5238_));
  NAND2_X1   g02803(.A1(new_n5203_), .A2(new_n2576_), .ZN(new_n5239_));
  INV_X1     g02804(.I(new_n5206_), .ZN(new_n5240_));
  NAND2_X1   g02805(.A1(new_n2577_), .A2(new_n5240_), .ZN(new_n5241_));
  AOI21_X1   g02806(.A1(new_n5239_), .A2(new_n5241_), .B(new_n3284_), .ZN(new_n5242_));
  NOR3_X1    g02807(.A1(new_n5238_), .A2(pi0062), .A3(new_n5242_), .ZN(new_n5243_));
  NAND2_X1   g02808(.A1(new_n5204_), .A2(new_n3320_), .ZN(new_n5244_));
  NAND2_X1   g02809(.A1(new_n3472_), .A2(new_n5206_), .ZN(new_n5245_));
  AOI21_X1   g02810(.A1(new_n5244_), .A2(new_n5245_), .B(new_n3471_), .ZN(new_n5246_));
  NOR3_X1    g02811(.A1(new_n5243_), .A2(new_n3425_), .A3(new_n5246_), .ZN(new_n5247_));
  OAI21_X1   g02812(.A1(new_n5206_), .A2(new_n3291_), .B(new_n5143_), .ZN(new_n5248_));
  NOR2_X1    g02813(.A1(new_n5240_), .A2(new_n3307_), .ZN(new_n5249_));
  INV_X1     g02814(.I(new_n5249_), .ZN(new_n5250_));
  NAND2_X1   g02815(.A1(new_n5250_), .A2(new_n2577_), .ZN(new_n5251_));
  NOR2_X1    g02816(.A1(new_n5149_), .A2(new_n5202_), .ZN(new_n5252_));
  INV_X1     g02817(.I(new_n5252_), .ZN(new_n5253_));
  OAI21_X1   g02818(.A1(new_n5253_), .A2(new_n2577_), .B(new_n5251_), .ZN(new_n5254_));
  NAND2_X1   g02819(.A1(new_n5254_), .A2(pi0056), .ZN(new_n5255_));
  NAND2_X1   g02820(.A1(new_n5249_), .A2(new_n2612_), .ZN(new_n5256_));
  OAI21_X1   g02821(.A1(new_n5252_), .A2(new_n2612_), .B(new_n5256_), .ZN(new_n5257_));
  AOI21_X1   g02822(.A1(new_n5257_), .A2(pi0055), .B(pi0056), .ZN(new_n5258_));
  AOI21_X1   g02823(.A1(new_n5249_), .A2(pi0299), .B(new_n5088_), .ZN(new_n5259_));
  INV_X1     g02824(.I(new_n5259_), .ZN(new_n5260_));
  OAI21_X1   g02825(.A1(new_n5260_), .A2(new_n2562_), .B(new_n2602_), .ZN(new_n5261_));
  NAND2_X1   g02826(.A1(new_n5260_), .A2(new_n2565_), .ZN(new_n5262_));
  AOI21_X1   g02827(.A1(new_n5253_), .A2(pi0299), .B(new_n5088_), .ZN(new_n5263_));
  NAND2_X1   g02828(.A1(new_n5260_), .A2(new_n3273_), .ZN(new_n5264_));
  OAI21_X1   g02829(.A1(new_n5263_), .A2(new_n3273_), .B(new_n5264_), .ZN(new_n5265_));
  NAND2_X1   g02830(.A1(new_n5265_), .A2(new_n2564_), .ZN(new_n5266_));
  AOI21_X1   g02831(.A1(new_n5266_), .A2(new_n5262_), .B(new_n3444_), .ZN(new_n5267_));
  OAI21_X1   g02832(.A1(new_n5263_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n5268_));
  AOI21_X1   g02833(.A1(new_n5098_), .A2(new_n5216_), .B(pi0039), .ZN(new_n5269_));
  INV_X1     g02834(.I(new_n5220_), .ZN(new_n5270_));
  NAND3_X1   g02835(.A1(new_n5166_), .A2(new_n5057_), .A3(new_n5270_), .ZN(new_n5271_));
  AOI21_X1   g02836(.A1(new_n5271_), .A2(new_n5269_), .B(new_n5268_), .ZN(new_n5272_));
  OAI21_X1   g02837(.A1(new_n5260_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n5273_));
  OAI21_X1   g02838(.A1(new_n5260_), .A2(new_n2572_), .B(pi0100), .ZN(new_n5274_));
  NOR2_X1    g02839(.A1(new_n5173_), .A2(new_n5202_), .ZN(new_n5275_));
  NOR2_X1    g02840(.A1(new_n5275_), .A2(new_n2628_), .ZN(new_n5276_));
  NOR3_X1    g02841(.A1(new_n5276_), .A2(new_n2573_), .A3(new_n5088_), .ZN(new_n5277_));
  OAI22_X1   g02842(.A1(new_n5272_), .A2(new_n5273_), .B1(new_n5274_), .B2(new_n5277_), .ZN(new_n5278_));
  OR2_X2     g02843(.A1(new_n5265_), .A2(new_n3458_), .Z(new_n5279_));
  OAI21_X1   g02844(.A1(new_n5278_), .A2(pi0087), .B(new_n5279_), .ZN(new_n5280_));
  OAI21_X1   g02845(.A1(new_n5260_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n5281_));
  AOI21_X1   g02846(.A1(new_n5280_), .A2(new_n3465_), .B(new_n5281_), .ZN(new_n5282_));
  NOR3_X1    g02847(.A1(new_n5282_), .A2(new_n2563_), .A3(new_n5267_), .ZN(new_n5283_));
  OAI21_X1   g02848(.A1(new_n5283_), .A2(new_n5261_), .B(new_n5258_), .ZN(new_n5284_));
  NAND3_X1   g02849(.A1(new_n5284_), .A2(new_n3471_), .A3(new_n5255_), .ZN(new_n5285_));
  NOR2_X1    g02850(.A1(new_n5252_), .A2(new_n3472_), .ZN(new_n5286_));
  NOR2_X1    g02851(.A1(new_n5250_), .A2(new_n3320_), .ZN(new_n5287_));
  OAI21_X1   g02852(.A1(new_n5286_), .A2(new_n5287_), .B(pi0062), .ZN(new_n5288_));
  AND3_X2    g02853(.A1(new_n5285_), .A2(new_n3291_), .A3(new_n5288_), .Z(new_n5289_));
  OAI21_X1   g02854(.A1(new_n5249_), .A2(new_n3291_), .B(pi0242), .ZN(new_n5290_));
  OAI22_X1   g02855(.A1(new_n5289_), .A2(new_n5290_), .B1(new_n5247_), .B2(new_n5248_), .ZN(new_n5291_));
  AOI22_X1   g02856(.A1(new_n5045_), .A2(new_n5291_), .B1(new_n5198_), .B2(new_n5142_), .ZN(po0165));
  NOR3_X1    g02857(.A1(new_n2577_), .A2(new_n2471_), .A3(new_n2530_), .ZN(new_n5294_));
  NAND2_X1   g02858(.A1(pi0057), .A2(pi0059), .ZN(new_n5295_));
  AOI21_X1   g02859(.A1(new_n5294_), .A2(new_n5295_), .B(new_n3291_), .ZN(new_n5296_));
  NOR2_X1    g02860(.A1(new_n2587_), .A2(new_n3273_), .ZN(new_n5297_));
  AOI21_X1   g02861(.A1(new_n5297_), .A2(new_n2570_), .B(new_n3284_), .ZN(new_n5298_));
  NOR2_X1    g02862(.A1(new_n2567_), .A2(pi0054), .ZN(new_n5299_));
  AOI21_X1   g02863(.A1(new_n5297_), .A2(new_n5299_), .B(new_n2625_), .ZN(new_n5300_));
  INV_X1     g02864(.I(new_n5300_), .ZN(new_n5301_));
  NOR2_X1    g02865(.A1(new_n5297_), .A2(new_n3458_), .ZN(new_n5302_));
  NOR2_X1    g02866(.A1(new_n5302_), .A2(pi0075), .ZN(new_n5303_));
  INV_X1     g02867(.I(new_n5303_), .ZN(new_n5304_));
  NOR2_X1    g02868(.A1(pi0054), .A2(pi0092), .ZN(new_n5305_));
  NOR2_X1    g02869(.A1(new_n2669_), .A2(pi0142), .ZN(new_n5306_));
  NOR2_X1    g02870(.A1(new_n5306_), .A2(pi0299), .ZN(new_n5307_));
  AOI21_X1   g02871(.A1(new_n2707_), .A2(pi0299), .B(new_n5307_), .ZN(new_n5308_));
  INV_X1     g02872(.I(new_n5308_), .ZN(new_n5309_));
  NOR2_X1    g02873(.A1(pi0041), .A2(pi0099), .ZN(new_n5310_));
  INV_X1     g02874(.I(new_n5310_), .ZN(new_n5311_));
  NOR2_X1    g02875(.A1(new_n5311_), .A2(pi0101), .ZN(new_n5312_));
  INV_X1     g02876(.I(new_n5312_), .ZN(new_n5313_));
  NOR3_X1    g02877(.A1(pi0042), .A2(pi0043), .A3(pi0052), .ZN(new_n5314_));
  NOR2_X1    g02878(.A1(pi0113), .A2(pi0116), .ZN(new_n5315_));
  INV_X1     g02879(.I(new_n5315_), .ZN(new_n5316_));
  NOR2_X1    g02880(.A1(pi0114), .A2(pi0115), .ZN(new_n5317_));
  INV_X1     g02881(.I(new_n5317_), .ZN(new_n5318_));
  NOR2_X1    g02882(.A1(new_n5316_), .A2(new_n5318_), .ZN(new_n5319_));
  NAND2_X1   g02883(.A1(new_n5319_), .A2(new_n5314_), .ZN(new_n5320_));
  NOR2_X1    g02884(.A1(new_n5320_), .A2(new_n5313_), .ZN(new_n5321_));
  INV_X1     g02885(.I(new_n5321_), .ZN(new_n5322_));
  NOR2_X1    g02886(.A1(new_n5322_), .A2(pi0044), .ZN(new_n5323_));
  NOR2_X1    g02887(.A1(new_n5323_), .A2(new_n5309_), .ZN(new_n5324_));
  INV_X1     g02888(.I(pi0683), .ZN(new_n5325_));
  INV_X1     g02889(.I(new_n5323_), .ZN(po1057));
  INV_X1     g02890(.I(pi0250), .ZN(new_n5327_));
  NOR2_X1    g02891(.A1(new_n5327_), .A2(pi0129), .ZN(new_n5328_));
  NOR2_X1    g02892(.A1(pi0824), .A2(pi0829), .ZN(new_n5329_));
  NOR2_X1    g02893(.A1(new_n5329_), .A2(new_n3082_), .ZN(new_n5330_));
  INV_X1     g02894(.I(new_n5330_), .ZN(new_n5331_));
  NOR2_X1    g02895(.A1(new_n5331_), .A2(pi1093), .ZN(po0740));
  AOI21_X1   g02896(.A1(po0740), .A2(new_n5327_), .B(new_n5328_), .ZN(new_n5333_));
  INV_X1     g02897(.I(new_n5333_), .ZN(new_n5334_));
  AOI21_X1   g02898(.A1(po1057), .A2(new_n5325_), .B(new_n5334_), .ZN(new_n5335_));
  NOR2_X1    g02899(.A1(new_n2530_), .A2(pi0039), .ZN(new_n5336_));
  INV_X1     g02900(.I(new_n5336_), .ZN(new_n5337_));
  NOR3_X1    g02901(.A1(new_n5337_), .A2(pi0038), .A3(new_n2702_), .ZN(new_n5338_));
  INV_X1     g02902(.I(new_n5338_), .ZN(new_n5339_));
  AOI21_X1   g02903(.A1(new_n5324_), .A2(new_n5335_), .B(new_n5339_), .ZN(new_n5340_));
  NOR2_X1    g02904(.A1(new_n3362_), .A2(new_n5308_), .ZN(new_n5341_));
  INV_X1     g02905(.I(new_n5341_), .ZN(new_n5342_));
  AOI21_X1   g02906(.A1(new_n5340_), .A2(new_n5342_), .B(pi0087), .ZN(new_n5343_));
  INV_X1     g02907(.I(new_n5343_), .ZN(new_n5344_));
  NOR2_X1    g02908(.A1(new_n2587_), .A2(pi0039), .ZN(new_n5345_));
  INV_X1     g02909(.I(new_n5345_), .ZN(new_n5346_));
  NOR2_X1    g02910(.A1(new_n5346_), .A2(new_n3265_), .ZN(new_n5347_));
  INV_X1     g02911(.I(new_n5347_), .ZN(new_n5348_));
  NOR2_X1    g02912(.A1(new_n2672_), .A2(pi0299), .ZN(new_n5349_));
  AOI21_X1   g02913(.A1(pi0210), .A2(pi0299), .B(new_n5349_), .ZN(new_n5350_));
  INV_X1     g02914(.I(new_n5350_), .ZN(new_n5351_));
  NAND2_X1   g02915(.A1(new_n3178_), .A2(new_n5351_), .ZN(new_n5352_));
  NOR2_X1    g02916(.A1(new_n2551_), .A2(pi0035), .ZN(new_n5353_));
  INV_X1     g02917(.I(new_n5353_), .ZN(new_n5354_));
  NOR3_X1    g02918(.A1(new_n3009_), .A2(pi0040), .A3(new_n5354_), .ZN(new_n5355_));
  INV_X1     g02919(.I(new_n5355_), .ZN(new_n5356_));
  NAND2_X1   g02920(.A1(new_n5356_), .A2(new_n5350_), .ZN(new_n5357_));
  AOI21_X1   g02921(.A1(new_n5352_), .A2(new_n5357_), .B(new_n2725_), .ZN(new_n5358_));
  INV_X1     g02922(.I(pi0058), .ZN(new_n5359_));
  NOR2_X1    g02923(.A1(new_n2829_), .A2(new_n5359_), .ZN(new_n5360_));
  NOR2_X1    g02924(.A1(new_n5360_), .A2(pi0090), .ZN(new_n5361_));
  INV_X1     g02925(.I(new_n5361_), .ZN(new_n5362_));
  INV_X1     g02926(.I(new_n2845_), .ZN(new_n5363_));
  NAND2_X1   g02927(.A1(new_n5363_), .A2(new_n2732_), .ZN(new_n5364_));
  INV_X1     g02928(.I(new_n2843_), .ZN(new_n5365_));
  INV_X1     g02929(.I(new_n2848_), .ZN(new_n5366_));
  INV_X1     g02930(.I(new_n2972_), .ZN(new_n5367_));
  NAND4_X1   g02931(.A1(new_n5367_), .A2(new_n2791_), .A3(new_n2855_), .A4(new_n2889_), .ZN(new_n5368_));
  AOI21_X1   g02932(.A1(new_n5368_), .A2(new_n2876_), .B(new_n2865_), .ZN(new_n5369_));
  OAI21_X1   g02933(.A1(new_n5369_), .A2(pi0108), .B(new_n2863_), .ZN(new_n5370_));
  NAND3_X1   g02934(.A1(new_n5370_), .A2(new_n2509_), .A3(new_n2980_), .ZN(new_n5371_));
  NAND3_X1   g02935(.A1(new_n5371_), .A2(new_n5365_), .A3(new_n5366_), .ZN(new_n5372_));
  AOI21_X1   g02936(.A1(new_n5372_), .A2(new_n2844_), .B(new_n5364_), .ZN(new_n5373_));
  OAI22_X1   g02937(.A1(new_n5373_), .A2(new_n5362_), .B1(new_n2985_), .B2(new_n2738_), .ZN(new_n5374_));
  INV_X1     g02938(.I(new_n2548_), .ZN(new_n5375_));
  AOI21_X1   g02939(.A1(new_n5375_), .A2(new_n3179_), .B(new_n2771_), .ZN(new_n5376_));
  NOR2_X1    g02940(.A1(new_n5376_), .A2(pi0035), .ZN(new_n5377_));
  INV_X1     g02941(.I(new_n5377_), .ZN(new_n5378_));
  AOI21_X1   g02942(.A1(new_n5374_), .A2(new_n2771_), .B(new_n5378_), .ZN(new_n5379_));
  OAI21_X1   g02943(.A1(new_n5379_), .A2(new_n2773_), .B(new_n2835_), .ZN(new_n5380_));
  AOI21_X1   g02944(.A1(new_n5380_), .A2(new_n2744_), .B(new_n2834_), .ZN(new_n5381_));
  OAI21_X1   g02945(.A1(new_n5381_), .A2(new_n3191_), .B(new_n2823_), .ZN(new_n5382_));
  AOI21_X1   g02946(.A1(new_n5382_), .A2(new_n2820_), .B(new_n5358_), .ZN(new_n5383_));
  OAI21_X1   g02947(.A1(new_n5383_), .A2(pi0095), .B(new_n3001_), .ZN(new_n5384_));
  NAND2_X1   g02948(.A1(new_n5384_), .A2(new_n2627_), .ZN(new_n5385_));
  INV_X1     g02949(.I(pi0835), .ZN(new_n5386_));
  INV_X1     g02950(.I(pi0984), .ZN(new_n5387_));
  NOR2_X1    g02951(.A1(new_n5386_), .A2(new_n5387_), .ZN(new_n5388_));
  INV_X1     g02952(.I(pi0979), .ZN(new_n5389_));
  OAI21_X1   g02953(.A1(pi0252), .A2(pi1001), .B(new_n5389_), .ZN(new_n5390_));
  NOR2_X1    g02954(.A1(new_n5390_), .A2(new_n5388_), .ZN(new_n5391_));
  INV_X1     g02955(.I(new_n5391_), .ZN(new_n5392_));
  NOR2_X1    g02956(.A1(new_n5392_), .A2(pi0287), .ZN(new_n5393_));
  NAND2_X1   g02957(.A1(new_n5393_), .A2(pi0835), .ZN(new_n5394_));
  INV_X1     g02958(.I(new_n5394_), .ZN(new_n5395_));
  NAND2_X1   g02959(.A1(new_n5395_), .A2(pi0950), .ZN(new_n5396_));
  NOR2_X1    g02960(.A1(new_n5396_), .A2(new_n3188_), .ZN(new_n5397_));
  NOR2_X1    g02961(.A1(pi0332), .A2(pi0468), .ZN(new_n5398_));
  INV_X1     g02962(.I(pi0681), .ZN(new_n5399_));
  INV_X1     g02963(.I(pi0662), .ZN(new_n5400_));
  NAND2_X1   g02964(.A1(new_n5400_), .A2(pi0680), .ZN(new_n5401_));
  NOR2_X1    g02965(.A1(new_n5401_), .A2(pi0661), .ZN(new_n5402_));
  NAND2_X1   g02966(.A1(new_n5402_), .A2(new_n5399_), .ZN(new_n5403_));
  INV_X1     g02967(.I(new_n5403_), .ZN(new_n5404_));
  INV_X1     g02968(.I(pi0614), .ZN(new_n5405_));
  INV_X1     g02969(.I(pi0642), .ZN(new_n5406_));
  NAND2_X1   g02970(.A1(new_n5405_), .A2(new_n5406_), .ZN(new_n5407_));
  NOR2_X1    g02971(.A1(new_n5407_), .A2(pi0616), .ZN(new_n5408_));
  NAND2_X1   g02972(.A1(new_n5408_), .A2(pi0603), .ZN(new_n5409_));
  INV_X1     g02973(.I(new_n5409_), .ZN(new_n5410_));
  NOR2_X1    g02974(.A1(new_n5410_), .A2(new_n5404_), .ZN(new_n5411_));
  INV_X1     g02975(.I(new_n5411_), .ZN(po1101));
  NOR2_X1    g02976(.A1(po1101), .A2(new_n5398_), .ZN(new_n5413_));
  INV_X1     g02977(.I(pi0970), .ZN(new_n5414_));
  INV_X1     g02978(.I(pi0972), .ZN(new_n5415_));
  INV_X1     g02979(.I(pi0975), .ZN(new_n5416_));
  NAND3_X1   g02980(.A1(new_n5414_), .A2(new_n5415_), .A3(new_n5416_), .ZN(new_n5417_));
  NOR4_X1    g02981(.A1(new_n5417_), .A2(pi0960), .A3(pi0963), .A4(pi0978), .ZN(new_n5418_));
  INV_X1     g02982(.I(new_n5418_), .ZN(new_n5419_));
  NOR2_X1    g02983(.A1(pi0907), .A2(pi0947), .ZN(new_n5420_));
  INV_X1     g02984(.I(new_n5420_), .ZN(new_n5421_));
  NOR2_X1    g02985(.A1(new_n5419_), .A2(new_n5421_), .ZN(new_n5422_));
  AOI21_X1   g02986(.A1(new_n5398_), .A2(new_n5422_), .B(new_n5413_), .ZN(new_n5423_));
  NAND4_X1   g02987(.A1(new_n5423_), .A2(new_n5397_), .A3(pi0216), .A4(pi0221), .ZN(new_n5424_));
  NAND2_X1   g02988(.A1(new_n5424_), .A2(new_n2531_), .ZN(new_n5425_));
  AOI21_X1   g02989(.A1(new_n5425_), .A2(new_n2436_), .B(new_n2628_), .ZN(new_n5426_));
  INV_X1     g02990(.I(new_n5413_), .ZN(new_n5427_));
  INV_X1     g02991(.I(pi0824), .ZN(new_n5428_));
  NOR2_X1    g02992(.A1(new_n3025_), .A2(new_n3041_), .ZN(new_n5429_));
  OAI22_X1   g02993(.A1(new_n5429_), .A2(new_n5329_), .B1(new_n5428_), .B2(pi1091), .ZN(new_n5430_));
  INV_X1     g02994(.I(new_n5430_), .ZN(new_n5431_));
  NOR2_X1    g02995(.A1(new_n5431_), .A2(new_n3082_), .ZN(new_n5432_));
  INV_X1     g02996(.I(new_n5432_), .ZN(po0950));
  NOR2_X1    g02997(.A1(po0950), .A2(new_n5394_), .ZN(new_n5434_));
  AOI21_X1   g02998(.A1(new_n5434_), .A2(new_n5427_), .B(new_n2530_), .ZN(new_n5435_));
  NOR2_X1    g02999(.A1(new_n5435_), .A2(new_n5422_), .ZN(new_n5436_));
  INV_X1     g03000(.I(new_n5398_), .ZN(new_n5437_));
  NOR2_X1    g03001(.A1(new_n2587_), .A2(new_n5437_), .ZN(new_n5438_));
  OAI21_X1   g03002(.A1(new_n5434_), .A2(new_n5398_), .B(po1101), .ZN(new_n5439_));
  AOI22_X1   g03003(.A1(new_n5438_), .A2(po1101), .B1(new_n2531_), .B2(new_n5439_), .ZN(new_n5440_));
  AOI21_X1   g03004(.A1(new_n5440_), .A2(new_n5422_), .B(new_n5436_), .ZN(new_n5441_));
  OAI21_X1   g03005(.A1(new_n5441_), .A2(new_n2436_), .B(new_n5426_), .ZN(new_n5442_));
  NOR4_X1    g03006(.A1(pi0969), .A2(pi0971), .A3(pi0974), .A4(pi0977), .ZN(new_n5443_));
  NOR4_X1    g03007(.A1(pi0587), .A2(pi0602), .A3(pi0961), .A4(pi0967), .ZN(new_n5444_));
  NAND2_X1   g03008(.A1(new_n5443_), .A2(new_n5444_), .ZN(new_n5445_));
  INV_X1     g03009(.I(new_n5445_), .ZN(new_n5446_));
  NOR2_X1    g03010(.A1(new_n5435_), .A2(new_n5446_), .ZN(new_n5447_));
  AOI21_X1   g03011(.A1(new_n5440_), .A2(new_n5446_), .B(new_n5447_), .ZN(new_n5448_));
  NOR2_X1    g03012(.A1(new_n5411_), .A2(new_n5398_), .ZN(new_n5449_));
  NOR2_X1    g03013(.A1(new_n5446_), .A2(new_n5437_), .ZN(new_n5450_));
  NOR2_X1    g03014(.A1(new_n5449_), .A2(new_n5450_), .ZN(new_n5451_));
  INV_X1     g03015(.I(new_n5451_), .ZN(new_n5452_));
  NAND4_X1   g03016(.A1(new_n5397_), .A2(pi0222), .A3(new_n5452_), .A4(pi0224), .ZN(new_n5453_));
  NAND2_X1   g03017(.A1(new_n5453_), .A2(new_n2531_), .ZN(new_n5454_));
  AOI21_X1   g03018(.A1(new_n5454_), .A2(new_n2668_), .B(pi0299), .ZN(new_n5455_));
  OAI21_X1   g03019(.A1(new_n5448_), .A2(new_n2668_), .B(new_n5455_), .ZN(new_n5456_));
  NAND3_X1   g03020(.A1(new_n5442_), .A2(new_n5456_), .A3(pi0039), .ZN(new_n5457_));
  NAND3_X1   g03021(.A1(new_n5385_), .A2(new_n3265_), .A3(new_n5457_), .ZN(new_n5458_));
  AOI21_X1   g03022(.A1(new_n5458_), .A2(new_n5348_), .B(pi0100), .ZN(new_n5459_));
  OAI21_X1   g03023(.A1(new_n5459_), .A2(new_n5344_), .B(new_n5305_), .ZN(new_n5460_));
  OAI21_X1   g03024(.A1(new_n5460_), .A2(new_n5304_), .B(new_n2625_), .ZN(new_n5461_));
  NAND3_X1   g03025(.A1(new_n5461_), .A2(new_n2602_), .A3(new_n5301_), .ZN(new_n5462_));
  AOI21_X1   g03026(.A1(new_n5462_), .A2(new_n3284_), .B(new_n5298_), .ZN(new_n5463_));
  AOI21_X1   g03027(.A1(new_n5297_), .A2(new_n3318_), .B(new_n3471_), .ZN(new_n5464_));
  INV_X1     g03028(.I(new_n5464_), .ZN(new_n5465_));
  OAI21_X1   g03029(.A1(new_n5463_), .A2(pi0062), .B(new_n5465_), .ZN(new_n5466_));
  OAI22_X1   g03030(.A1(new_n5466_), .A2(new_n3425_), .B1(new_n2582_), .B2(new_n5296_), .ZN(po0167));
  INV_X1     g03031(.I(pi1090), .ZN(po0170));
  INV_X1     g03032(.I(pi0030), .ZN(new_n5469_));
  NOR2_X1    g03033(.A1(new_n5469_), .A2(new_n2458_), .ZN(new_n5470_));
  AOI21_X1   g03034(.A1(new_n3322_), .A2(new_n2611_), .B(new_n5470_), .ZN(new_n5471_));
  NAND2_X1   g03035(.A1(new_n5403_), .A2(new_n5437_), .ZN(new_n5472_));
  INV_X1     g03036(.I(pi0907), .ZN(new_n5473_));
  NAND2_X1   g03037(.A1(new_n5398_), .A2(new_n5473_), .ZN(new_n5474_));
  NAND2_X1   g03038(.A1(new_n5472_), .A2(new_n5474_), .ZN(new_n5475_));
  NAND2_X1   g03039(.A1(new_n2470_), .A2(new_n2602_), .ZN(new_n5476_));
  NOR2_X1    g03040(.A1(new_n5476_), .A2(pi0059), .ZN(new_n5477_));
  NOR2_X1    g03041(.A1(new_n5477_), .A2(pi0228), .ZN(new_n5478_));
  NOR4_X1    g03042(.A1(new_n5471_), .A2(new_n2582_), .A3(new_n5475_), .A4(new_n5478_), .ZN(new_n5479_));
  NOR2_X1    g03043(.A1(new_n5471_), .A2(new_n5475_), .ZN(new_n5480_));
  NAND2_X1   g03044(.A1(new_n5476_), .A2(new_n2458_), .ZN(new_n5481_));
  NAND2_X1   g03045(.A1(new_n5480_), .A2(new_n5481_), .ZN(new_n5482_));
  AOI21_X1   g03046(.A1(new_n5482_), .A2(pi0059), .B(pi0057), .ZN(new_n5483_));
  INV_X1     g03047(.I(new_n5470_), .ZN(new_n5484_));
  NOR2_X1    g03048(.A1(new_n5475_), .A2(new_n2628_), .ZN(new_n5485_));
  INV_X1     g03049(.I(pi0602), .ZN(new_n5486_));
  NAND2_X1   g03050(.A1(new_n5398_), .A2(new_n5486_), .ZN(new_n5487_));
  NAND2_X1   g03051(.A1(new_n5472_), .A2(new_n5487_), .ZN(new_n5488_));
  INV_X1     g03052(.I(new_n5488_), .ZN(new_n5489_));
  AOI21_X1   g03053(.A1(new_n2628_), .A2(new_n5489_), .B(new_n5485_), .ZN(new_n5490_));
  NOR2_X1    g03054(.A1(new_n5490_), .A2(new_n5484_), .ZN(new_n5491_));
  NOR2_X1    g03055(.A1(new_n2606_), .A2(pi0054), .ZN(new_n5492_));
  OAI21_X1   g03056(.A1(new_n3322_), .A2(new_n5470_), .B(new_n2627_), .ZN(new_n5493_));
  NOR2_X1    g03057(.A1(new_n5493_), .A2(new_n5490_), .ZN(new_n5494_));
  AOI22_X1   g03058(.A1(new_n5494_), .A2(new_n2626_), .B1(new_n2659_), .B2(new_n5491_), .ZN(new_n5495_));
  AOI21_X1   g03059(.A1(new_n5495_), .A2(new_n5492_), .B(new_n2625_), .ZN(new_n5496_));
  OAI21_X1   g03060(.A1(new_n5491_), .A2(new_n5492_), .B(new_n5496_), .ZN(new_n5497_));
  NAND2_X1   g03061(.A1(new_n5497_), .A2(new_n2602_), .ZN(new_n5498_));
  INV_X1     g03062(.I(pi0054), .ZN(new_n5499_));
  NOR4_X1    g03063(.A1(new_n2530_), .A2(new_n5325_), .A3(new_n5323_), .A4(new_n5334_), .ZN(new_n5500_));
  INV_X1     g03064(.I(new_n5500_), .ZN(new_n5501_));
  AOI21_X1   g03065(.A1(new_n5437_), .A2(new_n5403_), .B(new_n5501_), .ZN(new_n5502_));
  NAND2_X1   g03066(.A1(new_n5502_), .A2(new_n5306_), .ZN(new_n5503_));
  INV_X1     g03067(.I(new_n5306_), .ZN(new_n5504_));
  INV_X1     g03068(.I(new_n5438_), .ZN(new_n5505_));
  NAND2_X1   g03069(.A1(new_n2531_), .A2(new_n5404_), .ZN(new_n5506_));
  OAI21_X1   g03070(.A1(new_n5505_), .A2(new_n5404_), .B(new_n5506_), .ZN(new_n5507_));
  NAND3_X1   g03071(.A1(new_n5507_), .A2(pi0252), .A3(new_n5504_), .ZN(new_n5508_));
  AOI22_X1   g03072(.A1(new_n5508_), .A2(new_n5503_), .B1(new_n5486_), .B2(new_n5398_), .ZN(new_n5509_));
  OAI21_X1   g03073(.A1(new_n5488_), .A2(new_n5484_), .B(new_n2628_), .ZN(new_n5510_));
  AOI21_X1   g03074(.A1(new_n5509_), .A2(new_n2458_), .B(new_n5510_), .ZN(new_n5511_));
  NOR2_X1    g03075(.A1(new_n5475_), .A2(new_n5484_), .ZN(new_n5512_));
  NOR2_X1    g03076(.A1(new_n5512_), .A2(new_n2628_), .ZN(new_n5513_));
  INV_X1     g03077(.I(new_n5513_), .ZN(new_n5514_));
  NAND2_X1   g03078(.A1(new_n5474_), .A2(new_n2458_), .ZN(new_n5515_));
  NAND3_X1   g03079(.A1(new_n5507_), .A2(pi0252), .A3(new_n2707_), .ZN(new_n5516_));
  NAND2_X1   g03080(.A1(new_n5502_), .A2(new_n2691_), .ZN(new_n5517_));
  AOI21_X1   g03081(.A1(new_n5516_), .A2(new_n5517_), .B(new_n5515_), .ZN(new_n5518_));
  OAI21_X1   g03082(.A1(new_n5518_), .A2(new_n5514_), .B(new_n2572_), .ZN(new_n5519_));
  NOR2_X1    g03083(.A1(new_n5511_), .A2(new_n5519_), .ZN(new_n5520_));
  INV_X1     g03084(.I(new_n5491_), .ZN(new_n5521_));
  OAI21_X1   g03085(.A1(new_n5521_), .A2(new_n2572_), .B(pi0100), .ZN(new_n5522_));
  NOR2_X1    g03086(.A1(new_n2458_), .A2(pi0030), .ZN(new_n5523_));
  NOR2_X1    g03087(.A1(new_n2629_), .A2(pi0223), .ZN(new_n5524_));
  INV_X1     g03088(.I(new_n5524_), .ZN(new_n5525_));
  NOR2_X1    g03089(.A1(new_n2530_), .A2(new_n5394_), .ZN(new_n5526_));
  INV_X1     g03090(.I(new_n5526_), .ZN(new_n5527_));
  NOR2_X1    g03091(.A1(new_n5428_), .A2(new_n3041_), .ZN(new_n5528_));
  INV_X1     g03092(.I(new_n5528_), .ZN(new_n5529_));
  NOR2_X1    g03093(.A1(new_n5529_), .A2(new_n3082_), .ZN(new_n5530_));
  INV_X1     g03094(.I(new_n5530_), .ZN(new_n5531_));
  INV_X1     g03095(.I(new_n3024_), .ZN(new_n5532_));
  NOR2_X1    g03096(.A1(new_n5532_), .A2(new_n3022_), .ZN(new_n5533_));
  NOR2_X1    g03097(.A1(new_n5531_), .A2(new_n5533_), .ZN(new_n5534_));
  AOI21_X1   g03098(.A1(new_n3086_), .A2(pi1091), .B(new_n5534_), .ZN(new_n5535_));
  NOR2_X1    g03099(.A1(new_n5527_), .A2(new_n5535_), .ZN(new_n5536_));
  NAND2_X1   g03100(.A1(new_n5536_), .A2(pi0224), .ZN(new_n5537_));
  NOR2_X1    g03101(.A1(new_n3024_), .A2(pi0829), .ZN(new_n5538_));
  NOR2_X1    g03102(.A1(new_n5538_), .A2(new_n3022_), .ZN(new_n5539_));
  NOR2_X1    g03103(.A1(new_n5531_), .A2(new_n5539_), .ZN(new_n5540_));
  NAND2_X1   g03104(.A1(new_n5526_), .A2(new_n5540_), .ZN(new_n5541_));
  INV_X1     g03105(.I(new_n5541_), .ZN(new_n5542_));
  NAND2_X1   g03106(.A1(new_n5542_), .A2(new_n2631_), .ZN(new_n5543_));
  AOI21_X1   g03107(.A1(new_n5537_), .A2(new_n5543_), .B(new_n5525_), .ZN(new_n5544_));
  INV_X1     g03108(.I(new_n5544_), .ZN(new_n5545_));
  AOI21_X1   g03109(.A1(new_n5545_), .A2(new_n2458_), .B(new_n5523_), .ZN(new_n5546_));
  AOI21_X1   g03110(.A1(new_n5546_), .A2(new_n5489_), .B(pi0299), .ZN(new_n5547_));
  INV_X1     g03111(.I(new_n5475_), .ZN(new_n5548_));
  NOR2_X1    g03112(.A1(new_n2441_), .A2(pi0215), .ZN(new_n5549_));
  INV_X1     g03113(.I(new_n5549_), .ZN(new_n5550_));
  INV_X1     g03114(.I(new_n5536_), .ZN(new_n5551_));
  NOR2_X1    g03115(.A1(new_n5542_), .A2(pi0216), .ZN(new_n5552_));
  AOI21_X1   g03116(.A1(pi0216), .A2(new_n5551_), .B(new_n5552_), .ZN(new_n5553_));
  NAND2_X1   g03117(.A1(new_n5553_), .A2(new_n2458_), .ZN(new_n5554_));
  OAI21_X1   g03118(.A1(new_n5554_), .A2(new_n5550_), .B(new_n5484_), .ZN(new_n5555_));
  AOI21_X1   g03119(.A1(new_n5555_), .A2(new_n5548_), .B(new_n2628_), .ZN(new_n5556_));
  NOR3_X1    g03120(.A1(new_n5556_), .A2(new_n5547_), .A3(new_n2627_), .ZN(new_n5557_));
  NOR2_X1    g03121(.A1(new_n2822_), .A2(new_n2536_), .ZN(new_n5558_));
  INV_X1     g03122(.I(new_n5558_), .ZN(new_n5559_));
  AOI21_X1   g03123(.A1(new_n2760_), .A2(pi0091), .B(pi0058), .ZN(new_n5560_));
  INV_X1     g03124(.I(new_n5560_), .ZN(new_n5561_));
  NOR2_X1    g03125(.A1(new_n2848_), .A2(new_n3130_), .ZN(new_n5562_));
  INV_X1     g03126(.I(new_n2878_), .ZN(new_n5563_));
  NOR2_X1    g03127(.A1(new_n5563_), .A2(new_n2513_), .ZN(new_n5564_));
  INV_X1     g03128(.I(new_n5564_), .ZN(new_n5565_));
  INV_X1     g03129(.I(new_n2794_), .ZN(new_n5566_));
  NOR2_X1    g03130(.A1(new_n2900_), .A2(po1049), .ZN(new_n5567_));
  INV_X1     g03131(.I(new_n2925_), .ZN(new_n5568_));
  NAND3_X1   g03132(.A1(new_n2945_), .A2(pi0085), .A3(new_n2491_), .ZN(new_n5569_));
  NAND2_X1   g03133(.A1(new_n5569_), .A2(new_n2931_), .ZN(new_n5570_));
  NAND2_X1   g03134(.A1(new_n5570_), .A2(new_n2541_), .ZN(new_n5571_));
  NAND2_X1   g03135(.A1(pi0068), .A2(pi0084), .ZN(new_n5572_));
  NAND3_X1   g03136(.A1(new_n2916_), .A2(new_n2488_), .A3(new_n5572_), .ZN(new_n5573_));
  NAND2_X1   g03137(.A1(new_n5571_), .A2(new_n5573_), .ZN(new_n5574_));
  NAND2_X1   g03138(.A1(new_n5574_), .A2(new_n2914_), .ZN(new_n5575_));
  AOI21_X1   g03139(.A1(new_n5575_), .A2(new_n2924_), .B(new_n5568_), .ZN(new_n5576_));
  INV_X1     g03140(.I(pi0067), .ZN(new_n5577_));
  OAI21_X1   g03141(.A1(new_n2903_), .A2(new_n5577_), .B(new_n2907_), .ZN(new_n5578_));
  NOR2_X1    g03142(.A1(new_n5576_), .A2(new_n5578_), .ZN(new_n5579_));
  OAI21_X1   g03143(.A1(new_n5579_), .A2(new_n2910_), .B(new_n2962_), .ZN(new_n5580_));
  AOI21_X1   g03144(.A1(new_n5580_), .A2(new_n5567_), .B(pi0081), .ZN(new_n5581_));
  NOR3_X1    g03145(.A1(new_n2968_), .A2(pi0102), .A3(new_n2504_), .ZN(new_n5582_));
  INV_X1     g03146(.I(new_n5582_), .ZN(new_n5583_));
  OAI21_X1   g03147(.A1(new_n5581_), .A2(new_n5583_), .B(new_n2883_), .ZN(new_n5584_));
  NAND2_X1   g03148(.A1(new_n5584_), .A2(new_n2881_), .ZN(new_n5585_));
  NAND2_X1   g03149(.A1(new_n5585_), .A2(new_n2790_), .ZN(new_n5586_));
  AOI21_X1   g03150(.A1(new_n5586_), .A2(new_n5566_), .B(pi0086), .ZN(new_n5587_));
  NOR2_X1    g03151(.A1(new_n5587_), .A2(new_n5565_), .ZN(new_n5588_));
  OAI21_X1   g03152(.A1(new_n5588_), .A2(new_n2981_), .B(new_n5562_), .ZN(new_n5589_));
  INV_X1     g03153(.I(pi0314), .ZN(new_n5590_));
  NOR2_X1    g03154(.A1(new_n5590_), .A2(pi0091), .ZN(new_n5591_));
  AOI21_X1   g03155(.A1(new_n5589_), .A2(new_n5591_), .B(new_n5561_), .ZN(new_n5592_));
  INV_X1     g03156(.I(new_n2881_), .ZN(new_n5593_));
  NAND2_X1   g03157(.A1(new_n2906_), .A2(new_n5567_), .ZN(new_n5594_));
  AOI21_X1   g03158(.A1(new_n5581_), .A2(new_n5594_), .B(new_n5583_), .ZN(new_n5595_));
  NOR3_X1    g03159(.A1(new_n5595_), .A2(pi0050), .A3(new_n2882_), .ZN(new_n5596_));
  OAI21_X1   g03160(.A1(new_n5596_), .A2(new_n5593_), .B(new_n2790_), .ZN(new_n5597_));
  NAND2_X1   g03161(.A1(new_n5597_), .A2(new_n5566_), .ZN(new_n5598_));
  AOI21_X1   g03162(.A1(new_n5598_), .A2(new_n2879_), .B(new_n5565_), .ZN(new_n5599_));
  OAI21_X1   g03163(.A1(new_n5599_), .A2(new_n2981_), .B(new_n5562_), .ZN(new_n5600_));
  NOR2_X1    g03164(.A1(pi0091), .A2(pi0314), .ZN(new_n5601_));
  NAND2_X1   g03165(.A1(new_n5600_), .A2(new_n5601_), .ZN(new_n5602_));
  NAND2_X1   g03166(.A1(new_n5602_), .A2(new_n5592_), .ZN(new_n5603_));
  AOI21_X1   g03167(.A1(new_n5603_), .A2(new_n2985_), .B(new_n2986_), .ZN(new_n5604_));
  NAND2_X1   g03168(.A1(new_n5375_), .A2(pi0841), .ZN(new_n5605_));
  AOI21_X1   g03169(.A1(new_n5605_), .A2(pi0093), .B(pi0035), .ZN(new_n5606_));
  OAI21_X1   g03170(.A1(new_n5604_), .A2(pi0093), .B(new_n5606_), .ZN(new_n5607_));
  NAND2_X1   g03171(.A1(new_n5607_), .A2(new_n2835_), .ZN(new_n5608_));
  AOI21_X1   g03172(.A1(new_n5608_), .A2(new_n3171_), .B(pi0072), .ZN(new_n5609_));
  OAI21_X1   g03173(.A1(new_n5609_), .A2(new_n5559_), .B(new_n3184_), .ZN(new_n5610_));
  NOR2_X1    g03174(.A1(new_n2772_), .A2(pi0841), .ZN(new_n5611_));
  NAND3_X1   g03175(.A1(new_n5611_), .A2(new_n2746_), .A3(new_n3059_), .ZN(new_n5612_));
  NOR2_X1    g03176(.A1(new_n5612_), .A2(new_n2725_), .ZN(new_n5613_));
  INV_X1     g03177(.I(new_n5613_), .ZN(new_n5614_));
  NOR2_X1    g03178(.A1(new_n5614_), .A2(pi0095), .ZN(new_n5615_));
  INV_X1     g03179(.I(new_n5615_), .ZN(new_n5616_));
  NOR2_X1    g03180(.A1(new_n5616_), .A2(pi0210), .ZN(new_n5617_));
  OAI21_X1   g03181(.A1(new_n5610_), .A2(new_n5617_), .B(new_n5437_), .ZN(new_n5618_));
  OAI21_X1   g03182(.A1(new_n5599_), .A2(new_n2979_), .B(new_n2734_), .ZN(new_n5619_));
  AOI21_X1   g03183(.A1(new_n5619_), .A2(new_n5601_), .B(new_n5561_), .ZN(new_n5620_));
  OAI21_X1   g03184(.A1(new_n5588_), .A2(new_n2979_), .B(new_n2734_), .ZN(new_n5621_));
  NAND2_X1   g03185(.A1(new_n5621_), .A2(new_n5591_), .ZN(new_n5622_));
  AOI21_X1   g03186(.A1(new_n5620_), .A2(new_n5622_), .B(pi0090), .ZN(new_n5623_));
  OAI21_X1   g03187(.A1(new_n5623_), .A2(new_n2986_), .B(new_n2771_), .ZN(new_n5624_));
  AOI21_X1   g03188(.A1(new_n5624_), .A2(new_n5606_), .B(pi0070), .ZN(new_n5625_));
  OAI21_X1   g03189(.A1(new_n5625_), .A2(new_n3172_), .B(new_n2821_), .ZN(new_n5626_));
  AOI21_X1   g03190(.A1(new_n5626_), .A2(new_n5558_), .B(new_n3185_), .ZN(new_n5627_));
  OAI21_X1   g03191(.A1(pi0210), .A2(new_n5616_), .B(new_n5627_), .ZN(new_n5628_));
  NAND2_X1   g03192(.A1(new_n5628_), .A2(new_n5398_), .ZN(new_n5629_));
  NAND2_X1   g03193(.A1(new_n5629_), .A2(new_n5618_), .ZN(new_n5630_));
  INV_X1     g03194(.I(pi0158), .ZN(new_n5631_));
  INV_X1     g03195(.I(pi0159), .ZN(new_n5632_));
  NOR2_X1    g03196(.A1(new_n5631_), .A2(new_n5632_), .ZN(new_n5633_));
  INV_X1     g03197(.I(new_n5633_), .ZN(new_n5634_));
  INV_X1     g03198(.I(pi0160), .ZN(new_n5635_));
  INV_X1     g03199(.I(pi0197), .ZN(new_n5636_));
  NOR2_X1    g03200(.A1(new_n5635_), .A2(new_n5636_), .ZN(new_n5637_));
  INV_X1     g03201(.I(new_n5637_), .ZN(new_n5638_));
  NOR2_X1    g03202(.A1(new_n5634_), .A2(new_n5638_), .ZN(new_n5639_));
  NAND3_X1   g03203(.A1(new_n5630_), .A2(new_n5548_), .A3(new_n5639_), .ZN(new_n5640_));
  INV_X1     g03204(.I(new_n5639_), .ZN(new_n5641_));
  NOR2_X1    g03205(.A1(new_n5610_), .A2(new_n5617_), .ZN(new_n5642_));
  NOR2_X1    g03206(.A1(new_n5642_), .A2(new_n5475_), .ZN(new_n5643_));
  NAND2_X1   g03207(.A1(new_n5643_), .A2(new_n5641_), .ZN(new_n5644_));
  AOI21_X1   g03208(.A1(new_n5640_), .A2(new_n5644_), .B(pi0228), .ZN(new_n5645_));
  OAI21_X1   g03209(.A1(new_n5645_), .A2(new_n5514_), .B(pi0232), .ZN(new_n5646_));
  NOR2_X1    g03210(.A1(new_n5616_), .A2(pi0198), .ZN(new_n5647_));
  INV_X1     g03211(.I(new_n5647_), .ZN(new_n5648_));
  AOI21_X1   g03212(.A1(new_n5627_), .A2(new_n5648_), .B(new_n5437_), .ZN(new_n5649_));
  NOR2_X1    g03213(.A1(new_n5610_), .A2(new_n5647_), .ZN(new_n5650_));
  NOR2_X1    g03214(.A1(new_n5650_), .A2(new_n5398_), .ZN(new_n5651_));
  NOR2_X1    g03215(.A1(new_n5651_), .A2(new_n5649_), .ZN(new_n5652_));
  NOR2_X1    g03216(.A1(new_n5652_), .A2(pi0228), .ZN(new_n5653_));
  NOR2_X1    g03217(.A1(new_n5653_), .A2(new_n5470_), .ZN(new_n5654_));
  NOR2_X1    g03218(.A1(new_n5654_), .A2(new_n5488_), .ZN(new_n5655_));
  INV_X1     g03219(.I(pi0145), .ZN(new_n5656_));
  INV_X1     g03220(.I(pi0180), .ZN(new_n5657_));
  INV_X1     g03221(.I(pi0181), .ZN(new_n5658_));
  INV_X1     g03222(.I(pi0182), .ZN(new_n5659_));
  NOR4_X1    g03223(.A1(new_n5656_), .A2(new_n5657_), .A3(new_n5658_), .A4(new_n5659_), .ZN(new_n5660_));
  AOI21_X1   g03224(.A1(new_n5650_), .A2(new_n2458_), .B(new_n5523_), .ZN(new_n5661_));
  INV_X1     g03225(.I(new_n5661_), .ZN(new_n5662_));
  OAI21_X1   g03226(.A1(new_n5662_), .A2(new_n5488_), .B(new_n2628_), .ZN(new_n5663_));
  NAND2_X1   g03227(.A1(new_n5660_), .A2(new_n2628_), .ZN(new_n5664_));
  AOI22_X1   g03228(.A1(new_n5655_), .A2(new_n5660_), .B1(new_n5663_), .B2(new_n5664_), .ZN(new_n5665_));
  INV_X1     g03229(.I(pi0232), .ZN(new_n5666_));
  NAND2_X1   g03230(.A1(new_n5643_), .A2(new_n2458_), .ZN(new_n5667_));
  NAND2_X1   g03231(.A1(new_n5667_), .A2(new_n5513_), .ZN(new_n5668_));
  NAND3_X1   g03232(.A1(new_n5663_), .A2(new_n5668_), .A3(new_n5666_), .ZN(new_n5669_));
  OAI21_X1   g03233(.A1(new_n5665_), .A2(new_n5646_), .B(new_n5669_), .ZN(new_n5670_));
  AOI21_X1   g03234(.A1(new_n5670_), .A2(new_n2627_), .B(new_n5557_), .ZN(new_n5671_));
  NOR3_X1    g03235(.A1(new_n5494_), .A2(new_n3265_), .A3(new_n5491_), .ZN(new_n5672_));
  AOI21_X1   g03236(.A1(new_n5671_), .A2(new_n3265_), .B(new_n5672_), .ZN(new_n5673_));
  OAI22_X1   g03237(.A1(new_n5673_), .A2(pi0100), .B1(new_n5520_), .B2(new_n5522_), .ZN(new_n5674_));
  NAND2_X1   g03238(.A1(new_n5491_), .A2(pi0087), .ZN(new_n5675_));
  OAI21_X1   g03239(.A1(new_n5674_), .A2(pi0087), .B(new_n5675_), .ZN(new_n5676_));
  AOI21_X1   g03240(.A1(new_n5495_), .A2(pi0075), .B(pi0092), .ZN(new_n5677_));
  OAI21_X1   g03241(.A1(new_n5676_), .A2(pi0075), .B(new_n5677_), .ZN(new_n5678_));
  NOR2_X1    g03242(.A1(new_n5495_), .A2(pi0075), .ZN(new_n5679_));
  NOR2_X1    g03243(.A1(new_n5521_), .A2(new_n3465_), .ZN(new_n5680_));
  OAI21_X1   g03244(.A1(new_n5679_), .A2(new_n5680_), .B(pi0092), .ZN(new_n5681_));
  NAND3_X1   g03245(.A1(new_n5678_), .A2(new_n5499_), .A3(new_n5681_), .ZN(new_n5682_));
  NAND2_X1   g03246(.A1(new_n5495_), .A2(new_n2605_), .ZN(new_n5683_));
  OAI21_X1   g03247(.A1(new_n2605_), .A2(new_n5491_), .B(new_n5683_), .ZN(new_n5684_));
  AOI21_X1   g03248(.A1(new_n5684_), .A2(pi0054), .B(pi0074), .ZN(new_n5685_));
  AOI21_X1   g03249(.A1(new_n5682_), .A2(new_n5685_), .B(new_n5498_), .ZN(new_n5686_));
  OAI21_X1   g03250(.A1(new_n5480_), .A2(new_n2602_), .B(new_n2470_), .ZN(new_n5687_));
  AOI21_X1   g03251(.A1(new_n5512_), .A2(new_n2471_), .B(pi0059), .ZN(new_n5688_));
  OAI21_X1   g03252(.A1(new_n5686_), .A2(new_n5687_), .B(new_n5688_), .ZN(new_n5689_));
  AOI21_X1   g03253(.A1(new_n5689_), .A2(new_n5483_), .B(new_n5479_), .ZN(po0171));
  NAND2_X1   g03254(.A1(new_n5409_), .A2(new_n5437_), .ZN(new_n5691_));
  INV_X1     g03255(.I(pi0947), .ZN(new_n5692_));
  NAND2_X1   g03256(.A1(new_n5398_), .A2(new_n5692_), .ZN(new_n5693_));
  NAND2_X1   g03257(.A1(new_n5691_), .A2(new_n5693_), .ZN(new_n5694_));
  NOR4_X1    g03258(.A1(new_n5471_), .A2(new_n2582_), .A3(new_n5478_), .A4(new_n5694_), .ZN(new_n5695_));
  NOR2_X1    g03259(.A1(new_n5471_), .A2(new_n5694_), .ZN(new_n5696_));
  NAND2_X1   g03260(.A1(new_n5696_), .A2(new_n5481_), .ZN(new_n5697_));
  AOI21_X1   g03261(.A1(new_n5697_), .A2(pi0059), .B(pi0057), .ZN(new_n5698_));
  INV_X1     g03262(.I(new_n5694_), .ZN(new_n5699_));
  INV_X1     g03263(.I(pi0587), .ZN(new_n5700_));
  NAND2_X1   g03264(.A1(new_n5398_), .A2(new_n5700_), .ZN(new_n5701_));
  NAND2_X1   g03265(.A1(new_n5691_), .A2(new_n5701_), .ZN(new_n5702_));
  NOR2_X1    g03266(.A1(new_n5702_), .A2(pi0299), .ZN(new_n5703_));
  AOI21_X1   g03267(.A1(pi0299), .A2(new_n5699_), .B(new_n5703_), .ZN(new_n5704_));
  NOR2_X1    g03268(.A1(new_n5704_), .A2(new_n5484_), .ZN(new_n5705_));
  NOR2_X1    g03269(.A1(new_n5493_), .A2(new_n5704_), .ZN(new_n5706_));
  AOI22_X1   g03270(.A1(new_n5706_), .A2(new_n2626_), .B1(new_n2659_), .B2(new_n5705_), .ZN(new_n5707_));
  AOI21_X1   g03271(.A1(new_n5707_), .A2(new_n5492_), .B(new_n2625_), .ZN(new_n5708_));
  OAI21_X1   g03272(.A1(new_n5492_), .A2(new_n5705_), .B(new_n5708_), .ZN(new_n5709_));
  NAND2_X1   g03273(.A1(new_n5709_), .A2(new_n2602_), .ZN(new_n5710_));
  NOR2_X1    g03274(.A1(new_n5694_), .A2(new_n5484_), .ZN(new_n5711_));
  NOR2_X1    g03275(.A1(new_n5711_), .A2(new_n2628_), .ZN(new_n5712_));
  INV_X1     g03276(.I(new_n5712_), .ZN(new_n5713_));
  NAND2_X1   g03277(.A1(new_n2531_), .A2(new_n5410_), .ZN(new_n5714_));
  NAND2_X1   g03278(.A1(new_n5438_), .A2(new_n5409_), .ZN(new_n5715_));
  AOI21_X1   g03279(.A1(new_n5715_), .A2(new_n5714_), .B(new_n2704_), .ZN(new_n5716_));
  OAI21_X1   g03280(.A1(new_n5409_), .A2(new_n5398_), .B(new_n5692_), .ZN(new_n5717_));
  NAND3_X1   g03281(.A1(new_n5716_), .A2(new_n2707_), .A3(new_n5717_), .ZN(new_n5718_));
  NAND4_X1   g03282(.A1(new_n5500_), .A2(new_n2691_), .A3(new_n5691_), .A4(new_n5693_), .ZN(new_n5719_));
  AOI21_X1   g03283(.A1(new_n5718_), .A2(new_n5719_), .B(pi0228), .ZN(new_n5720_));
  OAI21_X1   g03284(.A1(new_n5720_), .A2(new_n5713_), .B(new_n2572_), .ZN(new_n5721_));
  OAI21_X1   g03285(.A1(new_n5409_), .A2(new_n5398_), .B(new_n5700_), .ZN(new_n5722_));
  NAND2_X1   g03286(.A1(new_n5722_), .A2(new_n2458_), .ZN(new_n5723_));
  INV_X1     g03287(.I(new_n5691_), .ZN(new_n5724_));
  NOR3_X1    g03288(.A1(new_n5501_), .A2(pi0142), .A3(new_n5724_), .ZN(new_n5725_));
  AOI21_X1   g03289(.A1(new_n5716_), .A2(pi0142), .B(new_n5725_), .ZN(new_n5726_));
  INV_X1     g03290(.I(new_n5702_), .ZN(new_n5727_));
  NOR2_X1    g03291(.A1(new_n2670_), .A2(pi0228), .ZN(new_n5728_));
  AOI21_X1   g03292(.A1(new_n5727_), .A2(new_n5470_), .B(new_n5728_), .ZN(new_n5729_));
  OAI21_X1   g03293(.A1(new_n5726_), .A2(new_n5723_), .B(new_n5729_), .ZN(new_n5730_));
  NAND2_X1   g03294(.A1(new_n5716_), .A2(new_n5701_), .ZN(new_n5731_));
  NAND2_X1   g03295(.A1(new_n5731_), .A2(new_n5728_), .ZN(new_n5732_));
  AOI21_X1   g03296(.A1(new_n5730_), .A2(new_n5732_), .B(pi0299), .ZN(new_n5733_));
  AOI21_X1   g03297(.A1(new_n5705_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n5734_));
  OAI21_X1   g03298(.A1(new_n5733_), .A2(new_n5721_), .B(new_n5734_), .ZN(new_n5735_));
  INV_X1     g03299(.I(new_n5660_), .ZN(new_n5736_));
  NAND2_X1   g03300(.A1(new_n5661_), .A2(new_n5727_), .ZN(new_n5737_));
  NAND2_X1   g03301(.A1(new_n5737_), .A2(new_n5736_), .ZN(new_n5738_));
  OAI21_X1   g03302(.A1(new_n5654_), .A2(new_n5702_), .B(new_n5660_), .ZN(new_n5739_));
  AOI21_X1   g03303(.A1(new_n5739_), .A2(new_n5738_), .B(pi0299), .ZN(new_n5740_));
  NAND3_X1   g03304(.A1(new_n5630_), .A2(new_n5639_), .A3(new_n5699_), .ZN(new_n5741_));
  NOR2_X1    g03305(.A1(new_n5642_), .A2(new_n5694_), .ZN(new_n5742_));
  NAND2_X1   g03306(.A1(new_n5742_), .A2(new_n5641_), .ZN(new_n5743_));
  AOI21_X1   g03307(.A1(new_n5741_), .A2(new_n5743_), .B(pi0228), .ZN(new_n5744_));
  OAI21_X1   g03308(.A1(new_n5744_), .A2(new_n5713_), .B(pi0232), .ZN(new_n5745_));
  NAND2_X1   g03309(.A1(new_n5737_), .A2(new_n2628_), .ZN(new_n5746_));
  NAND2_X1   g03310(.A1(new_n5742_), .A2(new_n2458_), .ZN(new_n5747_));
  NAND2_X1   g03311(.A1(new_n5747_), .A2(new_n5712_), .ZN(new_n5748_));
  NAND3_X1   g03312(.A1(new_n5746_), .A2(new_n5748_), .A3(new_n5666_), .ZN(new_n5749_));
  OAI21_X1   g03313(.A1(new_n5740_), .A2(new_n5745_), .B(new_n5749_), .ZN(new_n5750_));
  NAND2_X1   g03314(.A1(new_n5546_), .A2(new_n5727_), .ZN(new_n5751_));
  NAND2_X1   g03315(.A1(new_n5751_), .A2(new_n2628_), .ZN(new_n5752_));
  NAND2_X1   g03316(.A1(new_n5752_), .A2(pi0039), .ZN(new_n5753_));
  AOI21_X1   g03317(.A1(new_n5554_), .A2(new_n5484_), .B(new_n5550_), .ZN(new_n5754_));
  NOR2_X1    g03318(.A1(new_n5550_), .A2(new_n2628_), .ZN(new_n5755_));
  INV_X1     g03319(.I(new_n5755_), .ZN(new_n5756_));
  AOI22_X1   g03320(.A1(new_n5754_), .A2(new_n5699_), .B1(new_n5713_), .B2(new_n5756_), .ZN(new_n5757_));
  OAI21_X1   g03321(.A1(new_n5753_), .A2(new_n5757_), .B(new_n3265_), .ZN(new_n5758_));
  AOI21_X1   g03322(.A1(new_n5750_), .A2(new_n2627_), .B(new_n5758_), .ZN(new_n5759_));
  NOR3_X1    g03323(.A1(new_n5706_), .A2(new_n3265_), .A3(new_n5705_), .ZN(new_n5760_));
  OAI21_X1   g03324(.A1(new_n5759_), .A2(new_n5760_), .B(new_n2702_), .ZN(new_n5761_));
  NAND3_X1   g03325(.A1(new_n5761_), .A2(new_n3458_), .A3(new_n5735_), .ZN(new_n5762_));
  NAND2_X1   g03326(.A1(new_n5705_), .A2(pi0087), .ZN(new_n5763_));
  NAND3_X1   g03327(.A1(new_n5762_), .A2(new_n3465_), .A3(new_n5763_), .ZN(new_n5764_));
  AOI21_X1   g03328(.A1(new_n5707_), .A2(pi0075), .B(pi0092), .ZN(new_n5765_));
  NAND2_X1   g03329(.A1(new_n5764_), .A2(new_n5765_), .ZN(new_n5766_));
  NOR2_X1    g03330(.A1(new_n5707_), .A2(pi0075), .ZN(new_n5767_));
  NOR3_X1    g03331(.A1(new_n5704_), .A2(new_n3465_), .A3(new_n5484_), .ZN(new_n5768_));
  OAI21_X1   g03332(.A1(new_n5767_), .A2(new_n5768_), .B(pi0092), .ZN(new_n5769_));
  NAND3_X1   g03333(.A1(new_n5766_), .A2(new_n5499_), .A3(new_n5769_), .ZN(new_n5770_));
  NAND2_X1   g03334(.A1(new_n5707_), .A2(new_n2605_), .ZN(new_n5771_));
  OAI21_X1   g03335(.A1(new_n2605_), .A2(new_n5705_), .B(new_n5771_), .ZN(new_n5772_));
  AOI21_X1   g03336(.A1(new_n5772_), .A2(pi0054), .B(pi0074), .ZN(new_n5773_));
  AOI21_X1   g03337(.A1(new_n5770_), .A2(new_n5773_), .B(new_n5710_), .ZN(new_n5774_));
  OAI21_X1   g03338(.A1(new_n5696_), .A2(new_n2602_), .B(new_n2470_), .ZN(new_n5775_));
  AOI21_X1   g03339(.A1(new_n5711_), .A2(new_n2471_), .B(pi0059), .ZN(new_n5776_));
  OAI21_X1   g03340(.A1(new_n5774_), .A2(new_n5775_), .B(new_n5776_), .ZN(new_n5777_));
  AOI21_X1   g03341(.A1(new_n5777_), .A2(new_n5698_), .B(new_n5695_), .ZN(po0172));
  NOR3_X1    g03342(.A1(new_n5437_), .A2(new_n5469_), .A3(new_n2458_), .ZN(new_n5779_));
  INV_X1     g03343(.I(new_n5779_), .ZN(new_n5780_));
  NOR2_X1    g03344(.A1(new_n5780_), .A2(new_n5414_), .ZN(new_n5781_));
  NOR2_X1    g03345(.A1(new_n5505_), .A2(pi0228), .ZN(new_n5782_));
  NAND2_X1   g03346(.A1(new_n5782_), .A2(pi0970), .ZN(new_n5783_));
  OAI21_X1   g03347(.A1(new_n5783_), .A2(new_n2612_), .B(pi0055), .ZN(new_n5784_));
  OAI21_X1   g03348(.A1(new_n5784_), .A2(new_n5781_), .B(new_n2470_), .ZN(new_n5785_));
  INV_X1     g03349(.I(pi0967), .ZN(new_n5786_));
  NAND2_X1   g03350(.A1(pi0299), .A2(pi0970), .ZN(new_n5787_));
  OAI21_X1   g03351(.A1(pi0299), .A2(new_n5786_), .B(new_n5787_), .ZN(new_n5788_));
  NAND2_X1   g03352(.A1(new_n5779_), .A2(new_n5788_), .ZN(new_n5789_));
  INV_X1     g03353(.I(new_n5789_), .ZN(new_n5790_));
  OAI21_X1   g03354(.A1(new_n5790_), .A2(new_n5492_), .B(pi0074), .ZN(new_n5791_));
  INV_X1     g03355(.I(new_n2626_), .ZN(new_n5792_));
  NAND2_X1   g03356(.A1(new_n2554_), .A2(new_n2458_), .ZN(new_n5793_));
  AOI21_X1   g03357(.A1(new_n5793_), .A2(new_n5484_), .B(new_n5437_), .ZN(new_n5794_));
  INV_X1     g03358(.I(new_n5794_), .ZN(new_n5795_));
  OAI21_X1   g03359(.A1(new_n5795_), .A2(new_n5786_), .B(new_n2628_), .ZN(new_n5796_));
  NOR2_X1    g03360(.A1(new_n5781_), .A2(new_n2628_), .ZN(new_n5797_));
  NAND2_X1   g03361(.A1(new_n5783_), .A2(new_n5797_), .ZN(new_n5798_));
  NAND3_X1   g03362(.A1(new_n5798_), .A2(new_n2627_), .A3(new_n5796_), .ZN(new_n5799_));
  OAI22_X1   g03363(.A1(new_n5799_), .A2(new_n5792_), .B1(new_n2658_), .B2(new_n5789_), .ZN(new_n5800_));
  INV_X1     g03364(.I(new_n5800_), .ZN(new_n5801_));
  AOI21_X1   g03365(.A1(new_n5801_), .A2(new_n5492_), .B(new_n5791_), .ZN(new_n5802_));
  NAND2_X1   g03366(.A1(new_n5800_), .A2(new_n2605_), .ZN(new_n5803_));
  NAND2_X1   g03367(.A1(new_n5790_), .A2(new_n2606_), .ZN(new_n5804_));
  NAND3_X1   g03368(.A1(new_n5803_), .A2(pi0054), .A3(new_n5804_), .ZN(new_n5805_));
  NAND2_X1   g03369(.A1(new_n5805_), .A2(new_n2625_), .ZN(new_n5806_));
  NAND2_X1   g03370(.A1(new_n5500_), .A2(new_n5398_), .ZN(new_n5807_));
  NOR2_X1    g03371(.A1(new_n5807_), .A2(new_n2707_), .ZN(new_n5808_));
  NOR3_X1    g03372(.A1(new_n5505_), .A2(new_n2704_), .A3(new_n2691_), .ZN(new_n5809_));
  OAI21_X1   g03373(.A1(new_n5809_), .A2(new_n5808_), .B(new_n2458_), .ZN(new_n5810_));
  OAI21_X1   g03374(.A1(new_n5810_), .A2(new_n5414_), .B(new_n5797_), .ZN(new_n5811_));
  NAND2_X1   g03375(.A1(new_n5811_), .A2(new_n2572_), .ZN(new_n5812_));
  AOI21_X1   g03376(.A1(new_n5398_), .A2(pi0030), .B(new_n2458_), .ZN(new_n5813_));
  OAI21_X1   g03377(.A1(new_n5505_), .A2(new_n2704_), .B(new_n5504_), .ZN(new_n5814_));
  NAND2_X1   g03378(.A1(new_n5807_), .A2(new_n5306_), .ZN(new_n5815_));
  NAND2_X1   g03379(.A1(new_n5814_), .A2(new_n5815_), .ZN(new_n5816_));
  AOI21_X1   g03380(.A1(new_n5816_), .A2(new_n2458_), .B(new_n5813_), .ZN(new_n5817_));
  AOI21_X1   g03381(.A1(new_n5817_), .A2(pi0967), .B(pi0299), .ZN(new_n5818_));
  NOR2_X1    g03382(.A1(new_n5812_), .A2(new_n5818_), .ZN(new_n5819_));
  OAI21_X1   g03383(.A1(new_n5789_), .A2(new_n2572_), .B(pi0100), .ZN(new_n5820_));
  AOI21_X1   g03384(.A1(new_n5790_), .A2(pi0039), .B(new_n3265_), .ZN(new_n5821_));
  NOR2_X1    g03385(.A1(new_n5813_), .A2(new_n2627_), .ZN(new_n5822_));
  OAI21_X1   g03386(.A1(new_n5545_), .A2(new_n5437_), .B(new_n2458_), .ZN(new_n5823_));
  NAND2_X1   g03387(.A1(new_n5823_), .A2(new_n2628_), .ZN(new_n5824_));
  NAND3_X1   g03388(.A1(new_n5553_), .A2(new_n5398_), .A3(new_n5549_), .ZN(new_n5825_));
  NAND2_X1   g03389(.A1(new_n5825_), .A2(new_n2458_), .ZN(new_n5826_));
  NAND2_X1   g03390(.A1(new_n5826_), .A2(pi0299), .ZN(new_n5827_));
  OAI22_X1   g03391(.A1(new_n5827_), .A2(new_n5414_), .B1(new_n5824_), .B2(new_n5786_), .ZN(new_n5828_));
  AOI21_X1   g03392(.A1(new_n5828_), .A2(new_n5822_), .B(pi0038), .ZN(new_n5829_));
  NOR2_X1    g03393(.A1(new_n5642_), .A2(new_n5437_), .ZN(new_n5830_));
  NAND3_X1   g03394(.A1(new_n5830_), .A2(new_n2458_), .A3(pi0970), .ZN(new_n5831_));
  AND2_X2    g03395(.A1(new_n5831_), .A2(new_n5797_), .Z(new_n5832_));
  NOR2_X1    g03396(.A1(new_n5662_), .A2(new_n5437_), .ZN(new_n5833_));
  AOI21_X1   g03397(.A1(new_n5833_), .A2(pi0967), .B(pi0299), .ZN(new_n5834_));
  NOR3_X1    g03398(.A1(new_n5834_), .A2(pi0232), .A3(new_n5832_), .ZN(new_n5835_));
  OAI21_X1   g03399(.A1(new_n5650_), .A2(new_n5660_), .B(new_n5780_), .ZN(new_n5836_));
  AND2_X2    g03400(.A1(new_n5649_), .A2(new_n2458_), .Z(new_n5837_));
  OAI22_X1   g03401(.A1(new_n5833_), .A2(new_n5660_), .B1(new_n5836_), .B2(new_n5837_), .ZN(new_n5838_));
  OAI21_X1   g03402(.A1(new_n5838_), .A2(new_n5786_), .B(new_n2628_), .ZN(new_n5839_));
  NAND2_X1   g03403(.A1(new_n5839_), .A2(pi0232), .ZN(new_n5840_));
  NOR2_X1    g03404(.A1(new_n5642_), .A2(new_n5637_), .ZN(new_n5841_));
  NOR2_X1    g03405(.A1(new_n5629_), .A2(new_n5638_), .ZN(new_n5842_));
  OAI21_X1   g03406(.A1(new_n5842_), .A2(new_n5841_), .B(new_n5398_), .ZN(new_n5843_));
  OAI21_X1   g03407(.A1(new_n5843_), .A2(pi0228), .B(new_n5780_), .ZN(new_n5844_));
  NAND3_X1   g03408(.A1(new_n5844_), .A2(pi0970), .A3(new_n5633_), .ZN(new_n5845_));
  NOR2_X1    g03409(.A1(new_n5634_), .A2(new_n2628_), .ZN(new_n5846_));
  OR2_X2     g03410(.A1(new_n5832_), .A2(new_n5846_), .Z(new_n5847_));
  AOI21_X1   g03411(.A1(new_n5847_), .A2(new_n5845_), .B(new_n5840_), .ZN(new_n5848_));
  OAI21_X1   g03412(.A1(new_n5848_), .A2(new_n5835_), .B(new_n2627_), .ZN(new_n5849_));
  AOI22_X1   g03413(.A1(new_n5849_), .A2(new_n5829_), .B1(new_n5799_), .B2(new_n5821_), .ZN(new_n5850_));
  OAI22_X1   g03414(.A1(new_n5850_), .A2(pi0100), .B1(new_n5819_), .B2(new_n5820_), .ZN(new_n5851_));
  NAND2_X1   g03415(.A1(new_n5790_), .A2(pi0087), .ZN(new_n5852_));
  OAI21_X1   g03416(.A1(new_n5851_), .A2(pi0087), .B(new_n5852_), .ZN(new_n5853_));
  AOI21_X1   g03417(.A1(new_n5801_), .A2(pi0075), .B(pi0092), .ZN(new_n5854_));
  OAI21_X1   g03418(.A1(new_n5853_), .A2(pi0075), .B(new_n5854_), .ZN(new_n5855_));
  NAND2_X1   g03419(.A1(new_n5790_), .A2(pi0075), .ZN(new_n5856_));
  OAI21_X1   g03420(.A1(new_n5801_), .A2(pi0075), .B(new_n5856_), .ZN(new_n5857_));
  AOI21_X1   g03421(.A1(new_n5857_), .A2(pi0092), .B(pi0054), .ZN(new_n5858_));
  AOI21_X1   g03422(.A1(new_n5855_), .A2(new_n5858_), .B(new_n5806_), .ZN(new_n5859_));
  NOR3_X1    g03423(.A1(new_n5859_), .A2(pi0055), .A3(new_n5802_), .ZN(new_n5860_));
  AOI21_X1   g03424(.A1(new_n5781_), .A2(new_n2471_), .B(pi0059), .ZN(new_n5861_));
  OAI21_X1   g03425(.A1(new_n5860_), .A2(new_n5785_), .B(new_n5861_), .ZN(new_n5862_));
  INV_X1     g03426(.I(new_n5781_), .ZN(new_n5863_));
  INV_X1     g03427(.I(new_n5476_), .ZN(new_n5864_));
  NOR2_X1    g03428(.A1(new_n5783_), .A2(new_n2612_), .ZN(new_n5865_));
  AOI21_X1   g03429(.A1(new_n5865_), .A2(new_n5864_), .B(new_n2469_), .ZN(new_n5866_));
  AOI21_X1   g03430(.A1(new_n5866_), .A2(new_n5863_), .B(pi0057), .ZN(new_n5867_));
  NAND2_X1   g03431(.A1(new_n5865_), .A2(new_n5477_), .ZN(new_n5868_));
  NAND2_X1   g03432(.A1(new_n5868_), .A2(new_n5863_), .ZN(new_n5869_));
  AOI22_X1   g03433(.A1(new_n5862_), .A2(new_n5867_), .B1(pi0057), .B2(new_n5869_), .ZN(po0173));
  NOR2_X1    g03434(.A1(new_n5780_), .A2(new_n5415_), .ZN(new_n5871_));
  NAND2_X1   g03435(.A1(new_n5782_), .A2(pi0972), .ZN(new_n5872_));
  OAI21_X1   g03436(.A1(new_n5872_), .A2(new_n2612_), .B(pi0055), .ZN(new_n5873_));
  OAI21_X1   g03437(.A1(new_n5873_), .A2(new_n5871_), .B(new_n2470_), .ZN(new_n5874_));
  INV_X1     g03438(.I(pi0961), .ZN(new_n5875_));
  NAND2_X1   g03439(.A1(pi0299), .A2(pi0972), .ZN(new_n5876_));
  OAI21_X1   g03440(.A1(pi0299), .A2(new_n5875_), .B(new_n5876_), .ZN(new_n5877_));
  NAND2_X1   g03441(.A1(new_n5779_), .A2(new_n5877_), .ZN(new_n5878_));
  INV_X1     g03442(.I(new_n5878_), .ZN(new_n5879_));
  OAI21_X1   g03443(.A1(new_n5879_), .A2(new_n5492_), .B(pi0074), .ZN(new_n5880_));
  OAI21_X1   g03444(.A1(new_n5795_), .A2(new_n5875_), .B(new_n2628_), .ZN(new_n5881_));
  NOR2_X1    g03445(.A1(new_n5871_), .A2(new_n2628_), .ZN(new_n5882_));
  NAND2_X1   g03446(.A1(new_n5872_), .A2(new_n5882_), .ZN(new_n5883_));
  NAND3_X1   g03447(.A1(new_n5883_), .A2(new_n2627_), .A3(new_n5881_), .ZN(new_n5884_));
  OAI22_X1   g03448(.A1(new_n5884_), .A2(new_n5792_), .B1(new_n2658_), .B2(new_n5878_), .ZN(new_n5885_));
  INV_X1     g03449(.I(new_n5885_), .ZN(new_n5886_));
  AOI21_X1   g03450(.A1(new_n5886_), .A2(new_n5492_), .B(new_n5880_), .ZN(new_n5887_));
  NAND2_X1   g03451(.A1(new_n5885_), .A2(new_n2605_), .ZN(new_n5888_));
  NAND2_X1   g03452(.A1(new_n5879_), .A2(new_n2606_), .ZN(new_n5889_));
  NAND3_X1   g03453(.A1(new_n5888_), .A2(pi0054), .A3(new_n5889_), .ZN(new_n5890_));
  NAND2_X1   g03454(.A1(new_n5890_), .A2(new_n2625_), .ZN(new_n5891_));
  OAI21_X1   g03455(.A1(new_n5810_), .A2(new_n5415_), .B(new_n5882_), .ZN(new_n5892_));
  NAND2_X1   g03456(.A1(new_n5892_), .A2(new_n2572_), .ZN(new_n5893_));
  AOI21_X1   g03457(.A1(new_n5817_), .A2(pi0961), .B(pi0299), .ZN(new_n5894_));
  NOR2_X1    g03458(.A1(new_n5893_), .A2(new_n5894_), .ZN(new_n5895_));
  OAI21_X1   g03459(.A1(new_n5878_), .A2(new_n2572_), .B(pi0100), .ZN(new_n5896_));
  AOI21_X1   g03460(.A1(new_n5879_), .A2(pi0039), .B(new_n3265_), .ZN(new_n5897_));
  OAI22_X1   g03461(.A1(new_n5827_), .A2(new_n5415_), .B1(new_n5824_), .B2(new_n5875_), .ZN(new_n5898_));
  AOI21_X1   g03462(.A1(new_n5898_), .A2(new_n5822_), .B(pi0038), .ZN(new_n5899_));
  NAND3_X1   g03463(.A1(new_n5830_), .A2(new_n2458_), .A3(pi0972), .ZN(new_n5900_));
  AND2_X2    g03464(.A1(new_n5900_), .A2(new_n5882_), .Z(new_n5901_));
  AOI21_X1   g03465(.A1(new_n5833_), .A2(pi0961), .B(pi0299), .ZN(new_n5902_));
  NOR3_X1    g03466(.A1(new_n5902_), .A2(pi0232), .A3(new_n5901_), .ZN(new_n5903_));
  OAI21_X1   g03467(.A1(new_n5838_), .A2(new_n5875_), .B(new_n2628_), .ZN(new_n5904_));
  NAND2_X1   g03468(.A1(new_n5904_), .A2(pi0232), .ZN(new_n5905_));
  NAND3_X1   g03469(.A1(new_n5844_), .A2(pi0972), .A3(new_n5633_), .ZN(new_n5906_));
  OR2_X2     g03470(.A1(new_n5901_), .A2(new_n5846_), .Z(new_n5907_));
  AOI21_X1   g03471(.A1(new_n5907_), .A2(new_n5906_), .B(new_n5905_), .ZN(new_n5908_));
  OAI21_X1   g03472(.A1(new_n5908_), .A2(new_n5903_), .B(new_n2627_), .ZN(new_n5909_));
  AOI22_X1   g03473(.A1(new_n5909_), .A2(new_n5899_), .B1(new_n5884_), .B2(new_n5897_), .ZN(new_n5910_));
  OAI22_X1   g03474(.A1(new_n5910_), .A2(pi0100), .B1(new_n5895_), .B2(new_n5896_), .ZN(new_n5911_));
  NAND2_X1   g03475(.A1(new_n5879_), .A2(pi0087), .ZN(new_n5912_));
  OAI21_X1   g03476(.A1(new_n5911_), .A2(pi0087), .B(new_n5912_), .ZN(new_n5913_));
  AOI21_X1   g03477(.A1(new_n5886_), .A2(pi0075), .B(pi0092), .ZN(new_n5914_));
  OAI21_X1   g03478(.A1(new_n5913_), .A2(pi0075), .B(new_n5914_), .ZN(new_n5915_));
  NAND2_X1   g03479(.A1(new_n5879_), .A2(pi0075), .ZN(new_n5916_));
  OAI21_X1   g03480(.A1(new_n5886_), .A2(pi0075), .B(new_n5916_), .ZN(new_n5917_));
  AOI21_X1   g03481(.A1(new_n5917_), .A2(pi0092), .B(pi0054), .ZN(new_n5918_));
  AOI21_X1   g03482(.A1(new_n5915_), .A2(new_n5918_), .B(new_n5891_), .ZN(new_n5919_));
  NOR3_X1    g03483(.A1(new_n5919_), .A2(pi0055), .A3(new_n5887_), .ZN(new_n5920_));
  AOI21_X1   g03484(.A1(new_n5871_), .A2(new_n2471_), .B(pi0059), .ZN(new_n5921_));
  OAI21_X1   g03485(.A1(new_n5920_), .A2(new_n5874_), .B(new_n5921_), .ZN(new_n5922_));
  INV_X1     g03486(.I(new_n5871_), .ZN(new_n5923_));
  NOR2_X1    g03487(.A1(new_n5872_), .A2(new_n2612_), .ZN(new_n5924_));
  AOI21_X1   g03488(.A1(new_n5924_), .A2(new_n5864_), .B(new_n2469_), .ZN(new_n5925_));
  AOI21_X1   g03489(.A1(new_n5925_), .A2(new_n5923_), .B(pi0057), .ZN(new_n5926_));
  NAND2_X1   g03490(.A1(new_n5924_), .A2(new_n5477_), .ZN(new_n5927_));
  NAND2_X1   g03491(.A1(new_n5927_), .A2(new_n5923_), .ZN(new_n5928_));
  AOI22_X1   g03492(.A1(new_n5922_), .A2(new_n5926_), .B1(pi0057), .B2(new_n5928_), .ZN(po0174));
  INV_X1     g03493(.I(pi0960), .ZN(new_n5930_));
  NOR2_X1    g03494(.A1(new_n5780_), .A2(new_n5930_), .ZN(new_n5931_));
  NAND2_X1   g03495(.A1(new_n5782_), .A2(pi0960), .ZN(new_n5932_));
  OAI21_X1   g03496(.A1(new_n5932_), .A2(new_n2612_), .B(pi0055), .ZN(new_n5933_));
  OAI21_X1   g03497(.A1(new_n5933_), .A2(new_n5931_), .B(new_n2470_), .ZN(new_n5934_));
  INV_X1     g03498(.I(pi0977), .ZN(new_n5935_));
  NAND2_X1   g03499(.A1(pi0299), .A2(pi0960), .ZN(new_n5936_));
  OAI21_X1   g03500(.A1(pi0299), .A2(new_n5935_), .B(new_n5936_), .ZN(new_n5937_));
  NAND2_X1   g03501(.A1(new_n5779_), .A2(new_n5937_), .ZN(new_n5938_));
  INV_X1     g03502(.I(new_n5938_), .ZN(new_n5939_));
  OAI21_X1   g03503(.A1(new_n5939_), .A2(new_n5492_), .B(pi0074), .ZN(new_n5940_));
  OAI21_X1   g03504(.A1(new_n5795_), .A2(new_n5935_), .B(new_n2628_), .ZN(new_n5941_));
  NOR2_X1    g03505(.A1(new_n5931_), .A2(new_n2628_), .ZN(new_n5942_));
  NAND2_X1   g03506(.A1(new_n5932_), .A2(new_n5942_), .ZN(new_n5943_));
  NAND3_X1   g03507(.A1(new_n5943_), .A2(new_n2627_), .A3(new_n5941_), .ZN(new_n5944_));
  OAI22_X1   g03508(.A1(new_n5944_), .A2(new_n5792_), .B1(new_n2658_), .B2(new_n5938_), .ZN(new_n5945_));
  INV_X1     g03509(.I(new_n5945_), .ZN(new_n5946_));
  AOI21_X1   g03510(.A1(new_n5946_), .A2(new_n5492_), .B(new_n5940_), .ZN(new_n5947_));
  NAND2_X1   g03511(.A1(new_n5945_), .A2(new_n2605_), .ZN(new_n5948_));
  NAND2_X1   g03512(.A1(new_n5939_), .A2(new_n2606_), .ZN(new_n5949_));
  NAND3_X1   g03513(.A1(new_n5948_), .A2(pi0054), .A3(new_n5949_), .ZN(new_n5950_));
  NAND2_X1   g03514(.A1(new_n5950_), .A2(new_n2625_), .ZN(new_n5951_));
  OAI21_X1   g03515(.A1(new_n5810_), .A2(new_n5930_), .B(new_n5942_), .ZN(new_n5952_));
  NAND2_X1   g03516(.A1(new_n5952_), .A2(new_n2572_), .ZN(new_n5953_));
  AOI21_X1   g03517(.A1(new_n5817_), .A2(pi0977), .B(pi0299), .ZN(new_n5954_));
  NOR2_X1    g03518(.A1(new_n5953_), .A2(new_n5954_), .ZN(new_n5955_));
  OAI21_X1   g03519(.A1(new_n5938_), .A2(new_n2572_), .B(pi0100), .ZN(new_n5956_));
  AOI21_X1   g03520(.A1(new_n5939_), .A2(pi0039), .B(new_n3265_), .ZN(new_n5957_));
  OAI22_X1   g03521(.A1(new_n5827_), .A2(new_n5930_), .B1(new_n5824_), .B2(new_n5935_), .ZN(new_n5958_));
  AOI21_X1   g03522(.A1(new_n5958_), .A2(new_n5822_), .B(pi0038), .ZN(new_n5959_));
  NAND3_X1   g03523(.A1(new_n5830_), .A2(new_n2458_), .A3(pi0960), .ZN(new_n5960_));
  AND2_X2    g03524(.A1(new_n5960_), .A2(new_n5942_), .Z(new_n5961_));
  AOI21_X1   g03525(.A1(new_n5833_), .A2(pi0977), .B(pi0299), .ZN(new_n5962_));
  NOR3_X1    g03526(.A1(new_n5962_), .A2(pi0232), .A3(new_n5961_), .ZN(new_n5963_));
  OAI21_X1   g03527(.A1(new_n5838_), .A2(new_n5935_), .B(new_n2628_), .ZN(new_n5964_));
  NAND2_X1   g03528(.A1(new_n5964_), .A2(pi0232), .ZN(new_n5965_));
  NAND3_X1   g03529(.A1(new_n5844_), .A2(pi0960), .A3(new_n5633_), .ZN(new_n5966_));
  OR2_X2     g03530(.A1(new_n5961_), .A2(new_n5846_), .Z(new_n5967_));
  AOI21_X1   g03531(.A1(new_n5967_), .A2(new_n5966_), .B(new_n5965_), .ZN(new_n5968_));
  OAI21_X1   g03532(.A1(new_n5968_), .A2(new_n5963_), .B(new_n2627_), .ZN(new_n5969_));
  AOI22_X1   g03533(.A1(new_n5969_), .A2(new_n5959_), .B1(new_n5944_), .B2(new_n5957_), .ZN(new_n5970_));
  OAI22_X1   g03534(.A1(new_n5970_), .A2(pi0100), .B1(new_n5955_), .B2(new_n5956_), .ZN(new_n5971_));
  NAND2_X1   g03535(.A1(new_n5939_), .A2(pi0087), .ZN(new_n5972_));
  OAI21_X1   g03536(.A1(new_n5971_), .A2(pi0087), .B(new_n5972_), .ZN(new_n5973_));
  AOI21_X1   g03537(.A1(new_n5946_), .A2(pi0075), .B(pi0092), .ZN(new_n5974_));
  OAI21_X1   g03538(.A1(new_n5973_), .A2(pi0075), .B(new_n5974_), .ZN(new_n5975_));
  NAND2_X1   g03539(.A1(new_n5939_), .A2(pi0075), .ZN(new_n5976_));
  OAI21_X1   g03540(.A1(new_n5946_), .A2(pi0075), .B(new_n5976_), .ZN(new_n5977_));
  AOI21_X1   g03541(.A1(new_n5977_), .A2(pi0092), .B(pi0054), .ZN(new_n5978_));
  AOI21_X1   g03542(.A1(new_n5975_), .A2(new_n5978_), .B(new_n5951_), .ZN(new_n5979_));
  NOR3_X1    g03543(.A1(new_n5979_), .A2(pi0055), .A3(new_n5947_), .ZN(new_n5980_));
  AOI21_X1   g03544(.A1(new_n5931_), .A2(new_n2471_), .B(pi0059), .ZN(new_n5981_));
  OAI21_X1   g03545(.A1(new_n5980_), .A2(new_n5934_), .B(new_n5981_), .ZN(new_n5982_));
  INV_X1     g03546(.I(new_n5931_), .ZN(new_n5983_));
  NOR2_X1    g03547(.A1(new_n5932_), .A2(new_n2612_), .ZN(new_n5984_));
  AOI21_X1   g03548(.A1(new_n5984_), .A2(new_n5864_), .B(new_n2469_), .ZN(new_n5985_));
  AOI21_X1   g03549(.A1(new_n5985_), .A2(new_n5983_), .B(pi0057), .ZN(new_n5986_));
  NAND2_X1   g03550(.A1(new_n5984_), .A2(new_n5477_), .ZN(new_n5987_));
  NAND2_X1   g03551(.A1(new_n5987_), .A2(new_n5983_), .ZN(new_n5988_));
  AOI22_X1   g03552(.A1(new_n5982_), .A2(new_n5986_), .B1(pi0057), .B2(new_n5988_), .ZN(po0175));
  INV_X1     g03553(.I(pi0963), .ZN(new_n5990_));
  NOR2_X1    g03554(.A1(new_n5780_), .A2(new_n5990_), .ZN(new_n5991_));
  NAND2_X1   g03555(.A1(new_n5782_), .A2(pi0963), .ZN(new_n5992_));
  OAI21_X1   g03556(.A1(new_n5992_), .A2(new_n2612_), .B(pi0055), .ZN(new_n5993_));
  OAI21_X1   g03557(.A1(new_n5993_), .A2(new_n5991_), .B(new_n2470_), .ZN(new_n5994_));
  INV_X1     g03558(.I(pi0969), .ZN(new_n5995_));
  NAND2_X1   g03559(.A1(pi0299), .A2(pi0963), .ZN(new_n5996_));
  OAI21_X1   g03560(.A1(pi0299), .A2(new_n5995_), .B(new_n5996_), .ZN(new_n5997_));
  NAND2_X1   g03561(.A1(new_n5779_), .A2(new_n5997_), .ZN(new_n5998_));
  INV_X1     g03562(.I(new_n5998_), .ZN(new_n5999_));
  OAI21_X1   g03563(.A1(new_n5999_), .A2(new_n5492_), .B(pi0074), .ZN(new_n6000_));
  OAI21_X1   g03564(.A1(new_n5795_), .A2(new_n5995_), .B(new_n2628_), .ZN(new_n6001_));
  NOR2_X1    g03565(.A1(new_n5991_), .A2(new_n2628_), .ZN(new_n6002_));
  NAND2_X1   g03566(.A1(new_n5992_), .A2(new_n6002_), .ZN(new_n6003_));
  NAND3_X1   g03567(.A1(new_n6003_), .A2(new_n2627_), .A3(new_n6001_), .ZN(new_n6004_));
  OAI22_X1   g03568(.A1(new_n6004_), .A2(new_n5792_), .B1(new_n2658_), .B2(new_n5998_), .ZN(new_n6005_));
  INV_X1     g03569(.I(new_n6005_), .ZN(new_n6006_));
  AOI21_X1   g03570(.A1(new_n6006_), .A2(new_n5492_), .B(new_n6000_), .ZN(new_n6007_));
  NAND2_X1   g03571(.A1(new_n6005_), .A2(new_n2605_), .ZN(new_n6008_));
  NAND2_X1   g03572(.A1(new_n5999_), .A2(new_n2606_), .ZN(new_n6009_));
  NAND3_X1   g03573(.A1(new_n6008_), .A2(pi0054), .A3(new_n6009_), .ZN(new_n6010_));
  NAND2_X1   g03574(.A1(new_n6010_), .A2(new_n2625_), .ZN(new_n6011_));
  OAI21_X1   g03575(.A1(new_n5810_), .A2(new_n5990_), .B(new_n6002_), .ZN(new_n6012_));
  NAND2_X1   g03576(.A1(new_n6012_), .A2(new_n2572_), .ZN(new_n6013_));
  AOI21_X1   g03577(.A1(new_n5817_), .A2(pi0969), .B(pi0299), .ZN(new_n6014_));
  NOR2_X1    g03578(.A1(new_n6013_), .A2(new_n6014_), .ZN(new_n6015_));
  OAI21_X1   g03579(.A1(new_n5998_), .A2(new_n2572_), .B(pi0100), .ZN(new_n6016_));
  AOI21_X1   g03580(.A1(new_n5999_), .A2(pi0039), .B(new_n3265_), .ZN(new_n6017_));
  OAI22_X1   g03581(.A1(new_n5827_), .A2(new_n5990_), .B1(new_n5824_), .B2(new_n5995_), .ZN(new_n6018_));
  AOI21_X1   g03582(.A1(new_n6018_), .A2(new_n5822_), .B(pi0038), .ZN(new_n6019_));
  NAND3_X1   g03583(.A1(new_n5830_), .A2(new_n2458_), .A3(pi0963), .ZN(new_n6020_));
  AND2_X2    g03584(.A1(new_n6020_), .A2(new_n6002_), .Z(new_n6021_));
  AOI21_X1   g03585(.A1(new_n5833_), .A2(pi0969), .B(pi0299), .ZN(new_n6022_));
  NOR3_X1    g03586(.A1(new_n6022_), .A2(pi0232), .A3(new_n6021_), .ZN(new_n6023_));
  OAI21_X1   g03587(.A1(new_n5838_), .A2(new_n5995_), .B(new_n2628_), .ZN(new_n6024_));
  NAND2_X1   g03588(.A1(new_n6024_), .A2(pi0232), .ZN(new_n6025_));
  NAND3_X1   g03589(.A1(new_n5844_), .A2(pi0963), .A3(new_n5633_), .ZN(new_n6026_));
  OR2_X2     g03590(.A1(new_n6021_), .A2(new_n5846_), .Z(new_n6027_));
  AOI21_X1   g03591(.A1(new_n6027_), .A2(new_n6026_), .B(new_n6025_), .ZN(new_n6028_));
  OAI21_X1   g03592(.A1(new_n6028_), .A2(new_n6023_), .B(new_n2627_), .ZN(new_n6029_));
  AOI22_X1   g03593(.A1(new_n6029_), .A2(new_n6019_), .B1(new_n6004_), .B2(new_n6017_), .ZN(new_n6030_));
  OAI22_X1   g03594(.A1(new_n6030_), .A2(pi0100), .B1(new_n6015_), .B2(new_n6016_), .ZN(new_n6031_));
  NAND2_X1   g03595(.A1(new_n5999_), .A2(pi0087), .ZN(new_n6032_));
  OAI21_X1   g03596(.A1(new_n6031_), .A2(pi0087), .B(new_n6032_), .ZN(new_n6033_));
  AOI21_X1   g03597(.A1(new_n6006_), .A2(pi0075), .B(pi0092), .ZN(new_n6034_));
  OAI21_X1   g03598(.A1(new_n6033_), .A2(pi0075), .B(new_n6034_), .ZN(new_n6035_));
  NAND2_X1   g03599(.A1(new_n5999_), .A2(pi0075), .ZN(new_n6036_));
  OAI21_X1   g03600(.A1(new_n6006_), .A2(pi0075), .B(new_n6036_), .ZN(new_n6037_));
  AOI21_X1   g03601(.A1(new_n6037_), .A2(pi0092), .B(pi0054), .ZN(new_n6038_));
  AOI21_X1   g03602(.A1(new_n6035_), .A2(new_n6038_), .B(new_n6011_), .ZN(new_n6039_));
  NOR3_X1    g03603(.A1(new_n6039_), .A2(pi0055), .A3(new_n6007_), .ZN(new_n6040_));
  AOI21_X1   g03604(.A1(new_n5991_), .A2(new_n2471_), .B(pi0059), .ZN(new_n6041_));
  OAI21_X1   g03605(.A1(new_n6040_), .A2(new_n5994_), .B(new_n6041_), .ZN(new_n6042_));
  INV_X1     g03606(.I(new_n5991_), .ZN(new_n6043_));
  NOR2_X1    g03607(.A1(new_n5992_), .A2(new_n2612_), .ZN(new_n6044_));
  AOI21_X1   g03608(.A1(new_n6044_), .A2(new_n5864_), .B(new_n2469_), .ZN(new_n6045_));
  AOI21_X1   g03609(.A1(new_n6045_), .A2(new_n6043_), .B(pi0057), .ZN(new_n6046_));
  NAND2_X1   g03610(.A1(new_n6044_), .A2(new_n5477_), .ZN(new_n6047_));
  NAND2_X1   g03611(.A1(new_n6047_), .A2(new_n6043_), .ZN(new_n6048_));
  AOI22_X1   g03612(.A1(new_n6042_), .A2(new_n6046_), .B1(pi0057), .B2(new_n6048_), .ZN(po0176));
  NOR2_X1    g03613(.A1(new_n5780_), .A2(new_n5416_), .ZN(new_n6050_));
  NAND2_X1   g03614(.A1(new_n5782_), .A2(pi0975), .ZN(new_n6051_));
  OAI21_X1   g03615(.A1(new_n6051_), .A2(new_n2612_), .B(pi0055), .ZN(new_n6052_));
  OAI21_X1   g03616(.A1(new_n6052_), .A2(new_n6050_), .B(new_n2470_), .ZN(new_n6053_));
  INV_X1     g03617(.I(pi0971), .ZN(new_n6054_));
  NAND2_X1   g03618(.A1(pi0299), .A2(pi0975), .ZN(new_n6055_));
  OAI21_X1   g03619(.A1(pi0299), .A2(new_n6054_), .B(new_n6055_), .ZN(new_n6056_));
  NAND2_X1   g03620(.A1(new_n5779_), .A2(new_n6056_), .ZN(new_n6057_));
  INV_X1     g03621(.I(new_n6057_), .ZN(new_n6058_));
  OAI21_X1   g03622(.A1(new_n6058_), .A2(new_n5492_), .B(pi0074), .ZN(new_n6059_));
  OAI21_X1   g03623(.A1(new_n5795_), .A2(new_n6054_), .B(new_n2628_), .ZN(new_n6060_));
  NOR2_X1    g03624(.A1(new_n6050_), .A2(new_n2628_), .ZN(new_n6061_));
  NAND2_X1   g03625(.A1(new_n6051_), .A2(new_n6061_), .ZN(new_n6062_));
  NAND3_X1   g03626(.A1(new_n6062_), .A2(new_n2627_), .A3(new_n6060_), .ZN(new_n6063_));
  OAI22_X1   g03627(.A1(new_n6063_), .A2(new_n5792_), .B1(new_n2658_), .B2(new_n6057_), .ZN(new_n6064_));
  INV_X1     g03628(.I(new_n6064_), .ZN(new_n6065_));
  AOI21_X1   g03629(.A1(new_n6065_), .A2(new_n5492_), .B(new_n6059_), .ZN(new_n6066_));
  NAND2_X1   g03630(.A1(new_n6064_), .A2(new_n2605_), .ZN(new_n6067_));
  NAND2_X1   g03631(.A1(new_n6058_), .A2(new_n2606_), .ZN(new_n6068_));
  NAND3_X1   g03632(.A1(new_n6067_), .A2(pi0054), .A3(new_n6068_), .ZN(new_n6069_));
  NAND2_X1   g03633(.A1(new_n6069_), .A2(new_n2625_), .ZN(new_n6070_));
  OAI21_X1   g03634(.A1(new_n5810_), .A2(new_n5416_), .B(new_n6061_), .ZN(new_n6071_));
  NAND2_X1   g03635(.A1(new_n6071_), .A2(new_n2572_), .ZN(new_n6072_));
  AOI21_X1   g03636(.A1(new_n5817_), .A2(pi0971), .B(pi0299), .ZN(new_n6073_));
  NOR2_X1    g03637(.A1(new_n6072_), .A2(new_n6073_), .ZN(new_n6074_));
  OAI21_X1   g03638(.A1(new_n6057_), .A2(new_n2572_), .B(pi0100), .ZN(new_n6075_));
  AOI21_X1   g03639(.A1(new_n6058_), .A2(pi0039), .B(new_n3265_), .ZN(new_n6076_));
  OAI22_X1   g03640(.A1(new_n5827_), .A2(new_n5416_), .B1(new_n5824_), .B2(new_n6054_), .ZN(new_n6077_));
  AOI21_X1   g03641(.A1(new_n6077_), .A2(new_n5822_), .B(pi0038), .ZN(new_n6078_));
  NAND3_X1   g03642(.A1(new_n5830_), .A2(new_n2458_), .A3(pi0975), .ZN(new_n6079_));
  AND2_X2    g03643(.A1(new_n6079_), .A2(new_n6061_), .Z(new_n6080_));
  AOI21_X1   g03644(.A1(new_n5833_), .A2(pi0971), .B(pi0299), .ZN(new_n6081_));
  NOR3_X1    g03645(.A1(new_n6081_), .A2(pi0232), .A3(new_n6080_), .ZN(new_n6082_));
  OAI21_X1   g03646(.A1(new_n5838_), .A2(new_n6054_), .B(new_n2628_), .ZN(new_n6083_));
  NAND2_X1   g03647(.A1(new_n6083_), .A2(pi0232), .ZN(new_n6084_));
  NAND3_X1   g03648(.A1(new_n5844_), .A2(pi0975), .A3(new_n5633_), .ZN(new_n6085_));
  OR2_X2     g03649(.A1(new_n6080_), .A2(new_n5846_), .Z(new_n6086_));
  AOI21_X1   g03650(.A1(new_n6086_), .A2(new_n6085_), .B(new_n6084_), .ZN(new_n6087_));
  OAI21_X1   g03651(.A1(new_n6087_), .A2(new_n6082_), .B(new_n2627_), .ZN(new_n6088_));
  AOI22_X1   g03652(.A1(new_n6088_), .A2(new_n6078_), .B1(new_n6063_), .B2(new_n6076_), .ZN(new_n6089_));
  OAI22_X1   g03653(.A1(new_n6089_), .A2(pi0100), .B1(new_n6074_), .B2(new_n6075_), .ZN(new_n6090_));
  NAND2_X1   g03654(.A1(new_n6058_), .A2(pi0087), .ZN(new_n6091_));
  OAI21_X1   g03655(.A1(new_n6090_), .A2(pi0087), .B(new_n6091_), .ZN(new_n6092_));
  AOI21_X1   g03656(.A1(new_n6065_), .A2(pi0075), .B(pi0092), .ZN(new_n6093_));
  OAI21_X1   g03657(.A1(new_n6092_), .A2(pi0075), .B(new_n6093_), .ZN(new_n6094_));
  NAND2_X1   g03658(.A1(new_n6058_), .A2(pi0075), .ZN(new_n6095_));
  OAI21_X1   g03659(.A1(new_n6065_), .A2(pi0075), .B(new_n6095_), .ZN(new_n6096_));
  AOI21_X1   g03660(.A1(new_n6096_), .A2(pi0092), .B(pi0054), .ZN(new_n6097_));
  AOI21_X1   g03661(.A1(new_n6094_), .A2(new_n6097_), .B(new_n6070_), .ZN(new_n6098_));
  NOR3_X1    g03662(.A1(new_n6098_), .A2(pi0055), .A3(new_n6066_), .ZN(new_n6099_));
  AOI21_X1   g03663(.A1(new_n6050_), .A2(new_n2471_), .B(pi0059), .ZN(new_n6100_));
  OAI21_X1   g03664(.A1(new_n6099_), .A2(new_n6053_), .B(new_n6100_), .ZN(new_n6101_));
  INV_X1     g03665(.I(new_n6050_), .ZN(new_n6102_));
  NOR2_X1    g03666(.A1(new_n6051_), .A2(new_n2612_), .ZN(new_n6103_));
  AOI21_X1   g03667(.A1(new_n6103_), .A2(new_n5864_), .B(new_n2469_), .ZN(new_n6104_));
  AOI21_X1   g03668(.A1(new_n6104_), .A2(new_n6102_), .B(pi0057), .ZN(new_n6105_));
  NAND2_X1   g03669(.A1(new_n6103_), .A2(new_n5477_), .ZN(new_n6106_));
  NAND2_X1   g03670(.A1(new_n6106_), .A2(new_n6102_), .ZN(new_n6107_));
  AOI22_X1   g03671(.A1(new_n6101_), .A2(new_n6105_), .B1(pi0057), .B2(new_n6107_), .ZN(po0177));
  INV_X1     g03672(.I(pi0978), .ZN(new_n6109_));
  NOR2_X1    g03673(.A1(new_n5780_), .A2(new_n6109_), .ZN(new_n6110_));
  INV_X1     g03674(.I(new_n6110_), .ZN(new_n6111_));
  NAND3_X1   g03675(.A1(new_n5782_), .A2(pi0978), .A3(new_n2611_), .ZN(new_n6112_));
  NAND3_X1   g03676(.A1(new_n6112_), .A2(pi0055), .A3(new_n6111_), .ZN(new_n6113_));
  NAND2_X1   g03677(.A1(new_n6113_), .A2(new_n2470_), .ZN(new_n6114_));
  INV_X1     g03678(.I(pi0974), .ZN(new_n6115_));
  NOR2_X1    g03679(.A1(new_n6115_), .A2(pi0299), .ZN(new_n6116_));
  AOI21_X1   g03680(.A1(pi0299), .A2(pi0978), .B(new_n6116_), .ZN(new_n6117_));
  NOR2_X1    g03681(.A1(new_n5780_), .A2(new_n6117_), .ZN(new_n6118_));
  OAI21_X1   g03682(.A1(new_n6118_), .A2(new_n5492_), .B(pi0074), .ZN(new_n6119_));
  NOR2_X1    g03683(.A1(new_n5795_), .A2(new_n6117_), .ZN(new_n6120_));
  INV_X1     g03684(.I(new_n6120_), .ZN(new_n6121_));
  AOI21_X1   g03685(.A1(new_n2458_), .A2(new_n2659_), .B(new_n6121_), .ZN(new_n6122_));
  INV_X1     g03686(.I(new_n6122_), .ZN(new_n6123_));
  AOI21_X1   g03687(.A1(new_n6123_), .A2(new_n5492_), .B(new_n6119_), .ZN(new_n6124_));
  NAND2_X1   g03688(.A1(new_n6122_), .A2(new_n2605_), .ZN(new_n6125_));
  NAND2_X1   g03689(.A1(new_n6118_), .A2(new_n2606_), .ZN(new_n6126_));
  NAND3_X1   g03690(.A1(new_n6125_), .A2(pi0054), .A3(new_n6126_), .ZN(new_n6127_));
  NAND2_X1   g03691(.A1(new_n6127_), .A2(new_n2625_), .ZN(new_n6128_));
  NOR2_X1    g03692(.A1(new_n6110_), .A2(new_n2628_), .ZN(new_n6129_));
  OAI21_X1   g03693(.A1(new_n5810_), .A2(new_n6109_), .B(new_n6129_), .ZN(new_n6130_));
  NAND2_X1   g03694(.A1(new_n6130_), .A2(new_n2572_), .ZN(new_n6131_));
  AOI21_X1   g03695(.A1(new_n5817_), .A2(pi0974), .B(pi0299), .ZN(new_n6132_));
  AOI21_X1   g03696(.A1(new_n6118_), .A2(new_n2573_), .B(new_n2702_), .ZN(new_n6133_));
  OAI21_X1   g03697(.A1(new_n6131_), .A2(new_n6132_), .B(new_n6133_), .ZN(new_n6134_));
  NAND2_X1   g03698(.A1(new_n6121_), .A2(new_n2627_), .ZN(new_n6135_));
  OAI21_X1   g03699(.A1(new_n2627_), .A2(new_n6118_), .B(new_n6135_), .ZN(new_n6136_));
  OAI22_X1   g03700(.A1(new_n5827_), .A2(new_n6109_), .B1(new_n5824_), .B2(new_n6115_), .ZN(new_n6137_));
  AOI21_X1   g03701(.A1(new_n6137_), .A2(new_n5822_), .B(pi0038), .ZN(new_n6138_));
  NAND3_X1   g03702(.A1(new_n5830_), .A2(new_n2458_), .A3(pi0978), .ZN(new_n6139_));
  AND2_X2    g03703(.A1(new_n6139_), .A2(new_n6129_), .Z(new_n6140_));
  AOI21_X1   g03704(.A1(new_n5833_), .A2(pi0974), .B(pi0299), .ZN(new_n6141_));
  NOR3_X1    g03705(.A1(new_n6141_), .A2(pi0232), .A3(new_n6140_), .ZN(new_n6142_));
  OAI21_X1   g03706(.A1(new_n5838_), .A2(new_n6115_), .B(new_n2628_), .ZN(new_n6143_));
  NAND2_X1   g03707(.A1(new_n6143_), .A2(pi0232), .ZN(new_n6144_));
  NAND3_X1   g03708(.A1(new_n5844_), .A2(pi0978), .A3(new_n5633_), .ZN(new_n6145_));
  OR2_X2     g03709(.A1(new_n6140_), .A2(new_n5846_), .Z(new_n6146_));
  AOI21_X1   g03710(.A1(new_n6146_), .A2(new_n6145_), .B(new_n6144_), .ZN(new_n6147_));
  OAI21_X1   g03711(.A1(new_n6147_), .A2(new_n6142_), .B(new_n2627_), .ZN(new_n6148_));
  AOI22_X1   g03712(.A1(new_n6148_), .A2(new_n6138_), .B1(pi0038), .B2(new_n6136_), .ZN(new_n6149_));
  OAI21_X1   g03713(.A1(new_n6149_), .A2(pi0100), .B(new_n6134_), .ZN(new_n6150_));
  NAND2_X1   g03714(.A1(new_n6118_), .A2(pi0087), .ZN(new_n6151_));
  OAI21_X1   g03715(.A1(new_n6150_), .A2(pi0087), .B(new_n6151_), .ZN(new_n6152_));
  AOI21_X1   g03716(.A1(new_n6123_), .A2(pi0075), .B(pi0092), .ZN(new_n6153_));
  OAI21_X1   g03717(.A1(new_n6152_), .A2(pi0075), .B(new_n6153_), .ZN(new_n6154_));
  NAND2_X1   g03718(.A1(new_n6118_), .A2(pi0075), .ZN(new_n6155_));
  OAI21_X1   g03719(.A1(new_n6123_), .A2(pi0075), .B(new_n6155_), .ZN(new_n6156_));
  AOI21_X1   g03720(.A1(new_n6156_), .A2(pi0092), .B(pi0054), .ZN(new_n6157_));
  AOI21_X1   g03721(.A1(new_n6154_), .A2(new_n6157_), .B(new_n6128_), .ZN(new_n6158_));
  NOR3_X1    g03722(.A1(new_n6158_), .A2(pi0055), .A3(new_n6124_), .ZN(new_n6159_));
  AOI21_X1   g03723(.A1(new_n6110_), .A2(new_n2471_), .B(pi0059), .ZN(new_n6160_));
  OAI21_X1   g03724(.A1(new_n6159_), .A2(new_n6114_), .B(new_n6160_), .ZN(new_n6161_));
  INV_X1     g03725(.I(new_n6112_), .ZN(new_n6162_));
  AOI21_X1   g03726(.A1(new_n6162_), .A2(new_n5864_), .B(new_n2469_), .ZN(new_n6163_));
  AOI21_X1   g03727(.A1(new_n6163_), .A2(new_n6111_), .B(pi0057), .ZN(new_n6164_));
  INV_X1     g03728(.I(new_n5477_), .ZN(new_n6165_));
  OAI21_X1   g03729(.A1(new_n6112_), .A2(new_n6165_), .B(new_n6111_), .ZN(new_n6166_));
  AOI22_X1   g03730(.A1(new_n6161_), .A2(new_n6164_), .B1(pi0057), .B2(new_n6166_), .ZN(po0178));
  INV_X1     g03731(.I(pi0954), .ZN(po1110));
  NOR3_X1    g03732(.A1(new_n2587_), .A2(new_n2569_), .A3(new_n3273_), .ZN(new_n6169_));
  NOR2_X1    g03733(.A1(new_n6169_), .A2(new_n2602_), .ZN(new_n6170_));
  NOR2_X1    g03734(.A1(new_n6170_), .A2(pi0056), .ZN(new_n6171_));
  NOR2_X1    g03735(.A1(new_n2530_), .A2(new_n3273_), .ZN(new_n6172_));
  INV_X1     g03736(.I(new_n6172_), .ZN(new_n6173_));
  NOR3_X1    g03737(.A1(new_n6173_), .A2(pi0092), .A3(new_n2565_), .ZN(new_n6174_));
  NOR2_X1    g03738(.A1(new_n6174_), .A2(new_n5499_), .ZN(new_n6175_));
  INV_X1     g03739(.I(new_n6175_), .ZN(new_n6176_));
  NOR2_X1    g03740(.A1(new_n5337_), .A2(new_n5792_), .ZN(new_n6177_));
  NOR2_X1    g03741(.A1(new_n6177_), .A2(new_n3465_), .ZN(new_n6178_));
  AOI21_X1   g03742(.A1(new_n6172_), .A2(new_n2564_), .B(new_n3444_), .ZN(new_n6179_));
  NOR2_X1    g03743(.A1(new_n6178_), .A2(new_n6179_), .ZN(new_n6180_));
  INV_X1     g03744(.I(new_n6180_), .ZN(new_n6181_));
  NAND3_X1   g03745(.A1(new_n5544_), .A2(new_n2628_), .A3(new_n5452_), .ZN(new_n6182_));
  NAND4_X1   g03746(.A1(new_n5553_), .A2(pi0299), .A3(new_n5423_), .A4(new_n5549_), .ZN(new_n6183_));
  NAND3_X1   g03747(.A1(new_n6183_), .A2(pi0039), .A3(new_n6182_), .ZN(new_n6184_));
  NOR2_X1    g03748(.A1(new_n5642_), .A2(new_n2628_), .ZN(new_n6185_));
  NOR2_X1    g03749(.A1(new_n5650_), .A2(pi0299), .ZN(new_n6186_));
  OAI21_X1   g03750(.A1(new_n6185_), .A2(new_n6186_), .B(new_n5666_), .ZN(new_n6187_));
  NAND3_X1   g03751(.A1(new_n5642_), .A2(pi0299), .A3(new_n5634_), .ZN(new_n6188_));
  NOR2_X1    g03752(.A1(new_n5842_), .A2(new_n5841_), .ZN(new_n6189_));
  NAND3_X1   g03753(.A1(new_n6189_), .A2(new_n5618_), .A3(new_n5846_), .ZN(new_n6190_));
  OAI22_X1   g03754(.A1(new_n5610_), .A2(new_n5647_), .B1(new_n5437_), .B2(new_n5736_), .ZN(new_n6191_));
  NAND2_X1   g03755(.A1(new_n5649_), .A2(new_n5660_), .ZN(new_n6192_));
  NAND3_X1   g03756(.A1(new_n6192_), .A2(new_n6191_), .A3(new_n2628_), .ZN(new_n6193_));
  NAND4_X1   g03757(.A1(new_n6190_), .A2(pi0232), .A3(new_n6188_), .A4(new_n6193_), .ZN(new_n6194_));
  NAND3_X1   g03758(.A1(new_n6194_), .A2(new_n2627_), .A3(new_n6187_), .ZN(new_n6195_));
  AND3_X2    g03759(.A1(new_n6195_), .A2(new_n3265_), .A3(new_n6184_), .Z(new_n6196_));
  NOR2_X1    g03760(.A1(new_n6196_), .A2(new_n5347_), .ZN(new_n6197_));
  OAI21_X1   g03761(.A1(new_n6197_), .A2(pi0100), .B(new_n5339_), .ZN(new_n6198_));
  AOI21_X1   g03762(.A1(new_n6198_), .A2(new_n5343_), .B(new_n2606_), .ZN(new_n6199_));
  OAI21_X1   g03763(.A1(new_n6199_), .A2(new_n6181_), .B(new_n5499_), .ZN(new_n6200_));
  AOI21_X1   g03764(.A1(new_n6200_), .A2(new_n6176_), .B(pi0074), .ZN(new_n6201_));
  OAI21_X1   g03765(.A1(new_n6201_), .A2(new_n5300_), .B(new_n2602_), .ZN(new_n6202_));
  NAND3_X1   g03766(.A1(new_n6202_), .A2(new_n3471_), .A3(new_n6171_), .ZN(new_n6203_));
  AOI21_X1   g03767(.A1(new_n6203_), .A2(new_n3291_), .B(new_n5296_), .ZN(po0195));
  NAND2_X1   g03768(.A1(po0195), .A2(po1110), .ZN(new_n6205_));
  OAI21_X1   g03769(.A1(pi0024), .A2(po1110), .B(new_n6205_), .ZN(po0182));
  NOR2_X1    g03770(.A1(new_n3487_), .A2(new_n3436_), .ZN(new_n6207_));
  OAI21_X1   g03771(.A1(new_n6207_), .A2(new_n2459_), .B(pi0092), .ZN(new_n6208_));
  NAND2_X1   g03772(.A1(new_n6208_), .A2(new_n2562_), .ZN(new_n6209_));
  AOI21_X1   g03773(.A1(new_n2460_), .A2(pi0075), .B(pi0092), .ZN(new_n6210_));
  NAND2_X1   g03774(.A1(new_n3371_), .A2(pi0299), .ZN(new_n6211_));
  NAND2_X1   g03775(.A1(new_n5504_), .A2(pi0252), .ZN(new_n6212_));
  NAND3_X1   g03776(.A1(new_n2531_), .A2(new_n2628_), .A3(new_n6212_), .ZN(new_n6213_));
  AOI21_X1   g03777(.A1(new_n6211_), .A2(new_n6213_), .B(new_n2702_), .ZN(new_n6214_));
  AOI21_X1   g03778(.A1(new_n6214_), .A2(new_n3322_), .B(pi0039), .ZN(new_n6215_));
  NAND3_X1   g03779(.A1(new_n3451_), .A2(new_n2702_), .A3(new_n2458_), .ZN(new_n6216_));
  OAI21_X1   g03780(.A1(new_n3487_), .A2(pi0100), .B(pi0039), .ZN(new_n6217_));
  NAND2_X1   g03781(.A1(new_n6217_), .A2(new_n3265_), .ZN(new_n6218_));
  AOI21_X1   g03782(.A1(new_n6216_), .A2(new_n6215_), .B(new_n6218_), .ZN(new_n6219_));
  OAI21_X1   g03783(.A1(new_n6219_), .A2(new_n2459_), .B(new_n3458_), .ZN(new_n6220_));
  OAI21_X1   g03784(.A1(new_n3487_), .A2(new_n2575_), .B(new_n2460_), .ZN(new_n6221_));
  AOI21_X1   g03785(.A1(new_n6221_), .A2(pi0087), .B(pi0075), .ZN(new_n6222_));
  NAND2_X1   g03786(.A1(new_n6220_), .A2(new_n6222_), .ZN(new_n6223_));
  AOI21_X1   g03787(.A1(new_n6223_), .A2(new_n6210_), .B(new_n6209_), .ZN(new_n6224_));
  OAI21_X1   g03788(.A1(new_n2459_), .A2(new_n2562_), .B(new_n2602_), .ZN(new_n6225_));
  INV_X1     g03789(.I(new_n5299_), .ZN(new_n6226_));
  NOR2_X1    g03790(.A1(new_n6226_), .A2(new_n2575_), .ZN(new_n6227_));
  NAND2_X1   g03791(.A1(new_n3322_), .A2(new_n6227_), .ZN(new_n6228_));
  OAI21_X1   g03792(.A1(new_n6228_), .A2(pi0074), .B(new_n2460_), .ZN(new_n6229_));
  AOI21_X1   g03793(.A1(new_n6229_), .A2(pi0055), .B(pi0056), .ZN(new_n6230_));
  OAI21_X1   g03794(.A1(new_n6224_), .A2(new_n6225_), .B(new_n6230_), .ZN(new_n6231_));
  AOI21_X1   g03795(.A1(new_n3322_), .A2(new_n2576_), .B(new_n3284_), .ZN(new_n6232_));
  AOI21_X1   g03796(.A1(new_n6232_), .A2(new_n2460_), .B(pi0062), .ZN(new_n6233_));
  NOR2_X1    g03797(.A1(new_n3487_), .A2(new_n2575_), .ZN(new_n6234_));
  NAND2_X1   g03798(.A1(new_n6234_), .A2(new_n3318_), .ZN(new_n6235_));
  NAND2_X1   g03799(.A1(new_n6235_), .A2(new_n2460_), .ZN(new_n6236_));
  AOI22_X1   g03800(.A1(new_n6231_), .A2(new_n6233_), .B1(pi0062), .B2(new_n6236_), .ZN(new_n6237_));
  NAND2_X1   g03801(.A1(new_n2459_), .A2(new_n3425_), .ZN(new_n6238_));
  OAI21_X1   g03802(.A1(new_n6237_), .A2(new_n3425_), .B(new_n6238_), .ZN(po0183));
  INV_X1     g03803(.I(pi0119), .ZN(new_n6240_));
  NAND2_X1   g03804(.A1(new_n2458_), .A2(pi0252), .ZN(new_n6241_));
  AOI21_X1   g03805(.A1(new_n6241_), .A2(new_n6240_), .B(pi0468), .ZN(new_n6242_));
  NAND2_X1   g03806(.A1(pi0119), .A2(pi1056), .ZN(new_n6243_));
  NAND2_X1   g03807(.A1(new_n6242_), .A2(new_n6243_), .ZN(po0184));
  NAND2_X1   g03808(.A1(pi0119), .A2(pi1077), .ZN(new_n6245_));
  NAND2_X1   g03809(.A1(new_n6242_), .A2(new_n6245_), .ZN(po0185));
  NAND2_X1   g03810(.A1(pi0119), .A2(pi1073), .ZN(new_n6247_));
  NAND2_X1   g03811(.A1(new_n6242_), .A2(new_n6247_), .ZN(po0186));
  NAND2_X1   g03812(.A1(pi0119), .A2(pi1041), .ZN(new_n6249_));
  NAND2_X1   g03813(.A1(new_n6242_), .A2(new_n6249_), .ZN(po0187));
  INV_X1     g03814(.I(pi0588), .ZN(new_n6251_));
  NAND2_X1   g03815(.A1(new_n5477_), .A2(new_n2582_), .ZN(po1038));
  NOR2_X1    g03816(.A1(pi0590), .A2(pi0591), .ZN(new_n6253_));
  INV_X1     g03817(.I(new_n6253_), .ZN(new_n6254_));
  INV_X1     g03818(.I(pi0567), .ZN(new_n6255_));
  NOR2_X1    g03819(.A1(new_n3041_), .A2(pi0122), .ZN(new_n6256_));
  INV_X1     g03820(.I(new_n6256_), .ZN(new_n6257_));
  NOR2_X1    g03821(.A1(new_n3082_), .A2(new_n5428_), .ZN(new_n6258_));
  INV_X1     g03822(.I(new_n6258_), .ZN(new_n6259_));
  NOR2_X1    g03823(.A1(new_n6259_), .A2(pi0098), .ZN(new_n6260_));
  INV_X1     g03824(.I(new_n6260_), .ZN(new_n6261_));
  NOR2_X1    g03825(.A1(new_n6261_), .A2(new_n6257_), .ZN(new_n6262_));
  INV_X1     g03826(.I(new_n6262_), .ZN(new_n6263_));
  NOR2_X1    g03827(.A1(new_n6263_), .A2(pi1091), .ZN(new_n6264_));
  INV_X1     g03828(.I(new_n6264_), .ZN(new_n6265_));
  NOR2_X1    g03829(.A1(new_n6265_), .A2(new_n6255_), .ZN(new_n6266_));
  AOI21_X1   g03830(.A1(new_n6266_), .A2(new_n6254_), .B(new_n6251_), .ZN(new_n6267_));
  INV_X1     g03831(.I(pi0592), .ZN(new_n6268_));
  INV_X1     g03832(.I(new_n6266_), .ZN(new_n6269_));
  NOR2_X1    g03833(.A1(new_n6269_), .A2(new_n6268_), .ZN(new_n6270_));
  NOR2_X1    g03834(.A1(new_n6269_), .A2(pi0592), .ZN(new_n6271_));
  INV_X1     g03835(.I(new_n6271_), .ZN(new_n6272_));
  INV_X1     g03836(.I(pi1197), .ZN(new_n6273_));
  INV_X1     g03837(.I(pi1198), .ZN(new_n6274_));
  XNOR2_X1   g03838(.A1(pi0421), .A2(pi0459), .ZN(new_n6275_));
  XOR2_X1    g03839(.A1(pi0432), .A2(pi0454), .Z(new_n6276_));
  XOR2_X1    g03840(.A1(new_n6275_), .A2(new_n6276_), .Z(new_n6277_));
  INV_X1     g03841(.I(pi0423), .ZN(new_n6278_));
  XOR2_X1    g03842(.A1(pi0419), .A2(pi0420), .Z(new_n6279_));
  XOR2_X1    g03843(.A1(new_n6279_), .A2(new_n6278_), .Z(new_n6280_));
  XNOR2_X1   g03844(.A1(pi0424), .A2(pi0425), .ZN(new_n6281_));
  XOR2_X1    g03845(.A1(new_n6280_), .A2(new_n6281_), .Z(new_n6282_));
  XOR2_X1    g03846(.A1(new_n6282_), .A2(new_n6277_), .Z(new_n6283_));
  NOR2_X1    g03847(.A1(pi0418), .A2(pi0437), .ZN(new_n6284_));
  INV_X1     g03848(.I(pi0418), .ZN(new_n6285_));
  INV_X1     g03849(.I(pi0437), .ZN(new_n6286_));
  NOR2_X1    g03850(.A1(new_n6285_), .A2(new_n6286_), .ZN(new_n6287_));
  OAI21_X1   g03851(.A1(new_n6287_), .A2(new_n6284_), .B(pi0417), .ZN(new_n6288_));
  INV_X1     g03852(.I(pi0417), .ZN(new_n6289_));
  NOR2_X1    g03853(.A1(new_n6286_), .A2(pi0418), .ZN(new_n6290_));
  NOR2_X1    g03854(.A1(new_n6285_), .A2(pi0437), .ZN(new_n6291_));
  OAI21_X1   g03855(.A1(new_n6290_), .A2(new_n6291_), .B(new_n6289_), .ZN(new_n6292_));
  NAND2_X1   g03856(.A1(new_n6288_), .A2(new_n6292_), .ZN(new_n6293_));
  XOR2_X1    g03857(.A1(pi0453), .A2(pi0464), .Z(new_n6294_));
  XOR2_X1    g03858(.A1(new_n6293_), .A2(new_n6294_), .Z(new_n6295_));
  XOR2_X1    g03859(.A1(new_n6295_), .A2(pi0431), .Z(new_n6296_));
  INV_X1     g03860(.I(pi0438), .ZN(new_n6297_));
  XOR2_X1    g03861(.A1(pi0415), .A2(pi0416), .Z(new_n6298_));
  XOR2_X1    g03862(.A1(new_n6298_), .A2(new_n6297_), .Z(new_n6299_));
  XOR2_X1    g03863(.A1(new_n6296_), .A2(new_n6299_), .Z(new_n6300_));
  OAI22_X1   g03864(.A1(new_n6300_), .A2(new_n6273_), .B1(new_n6274_), .B2(new_n6283_), .ZN(new_n6301_));
  INV_X1     g03865(.I(pi1196), .ZN(new_n6302_));
  NOR2_X1    g03866(.A1(new_n6302_), .A2(pi0592), .ZN(new_n6303_));
  INV_X1     g03867(.I(new_n6303_), .ZN(new_n6304_));
  XOR2_X1    g03868(.A1(pi0443), .A2(pi0444), .Z(new_n6305_));
  INV_X1     g03869(.I(pi0436), .ZN(new_n6306_));
  XNOR2_X1   g03870(.A1(pi0429), .A2(pi0435), .ZN(new_n6307_));
  XOR2_X1    g03871(.A1(pi0414), .A2(pi0422), .Z(new_n6308_));
  INV_X1     g03872(.I(pi0434), .ZN(new_n6309_));
  NAND2_X1   g03873(.A1(new_n6309_), .A2(pi0446), .ZN(new_n6310_));
  INV_X1     g03874(.I(pi0446), .ZN(new_n6311_));
  NAND2_X1   g03875(.A1(new_n6311_), .A2(pi0434), .ZN(new_n6312_));
  AOI21_X1   g03876(.A1(new_n6310_), .A2(new_n6312_), .B(new_n6308_), .ZN(new_n6313_));
  XNOR2_X1   g03877(.A1(pi0434), .A2(pi0446), .ZN(new_n6314_));
  AOI21_X1   g03878(.A1(new_n6308_), .A2(new_n6314_), .B(new_n6313_), .ZN(new_n6315_));
  XOR2_X1    g03879(.A1(new_n6315_), .A2(new_n6307_), .Z(new_n6316_));
  XOR2_X1    g03880(.A1(new_n6316_), .A2(new_n6306_), .Z(new_n6317_));
  XOR2_X1    g03881(.A1(new_n6317_), .A2(new_n6305_), .Z(new_n6318_));
  NOR2_X1    g03882(.A1(new_n6318_), .A2(new_n6304_), .ZN(new_n6319_));
  OR2_X2     g03883(.A1(new_n6319_), .A2(new_n6301_), .Z(new_n6320_));
  NOR2_X1    g03884(.A1(new_n6320_), .A2(new_n6272_), .ZN(new_n6321_));
  INV_X1     g03885(.I(pi0451), .ZN(new_n6322_));
  NOR2_X1    g03886(.A1(new_n6322_), .A2(pi0449), .ZN(new_n6323_));
  INV_X1     g03887(.I(pi0449), .ZN(new_n6324_));
  NOR2_X1    g03888(.A1(new_n6324_), .A2(pi0451), .ZN(new_n6325_));
  OAI21_X1   g03889(.A1(new_n6323_), .A2(new_n6325_), .B(pi0433), .ZN(new_n6326_));
  INV_X1     g03890(.I(pi0433), .ZN(new_n6327_));
  NOR2_X1    g03891(.A1(pi0449), .A2(pi0451), .ZN(new_n6328_));
  NOR2_X1    g03892(.A1(new_n6324_), .A2(new_n6322_), .ZN(new_n6329_));
  OAI21_X1   g03893(.A1(new_n6329_), .A2(new_n6328_), .B(new_n6327_), .ZN(new_n6330_));
  NAND2_X1   g03894(.A1(new_n6330_), .A2(new_n6326_), .ZN(new_n6331_));
  XOR2_X1    g03895(.A1(pi0426), .A2(pi0427), .Z(new_n6332_));
  INV_X1     g03896(.I(pi0428), .ZN(new_n6333_));
  NAND2_X1   g03897(.A1(new_n6333_), .A2(pi0430), .ZN(new_n6334_));
  INV_X1     g03898(.I(pi0430), .ZN(new_n6335_));
  NAND2_X1   g03899(.A1(new_n6335_), .A2(pi0428), .ZN(new_n6336_));
  AOI21_X1   g03900(.A1(new_n6334_), .A2(new_n6336_), .B(new_n6332_), .ZN(new_n6337_));
  XNOR2_X1   g03901(.A1(pi0428), .A2(pi0430), .ZN(new_n6338_));
  AOI21_X1   g03902(.A1(new_n6332_), .A2(new_n6338_), .B(new_n6337_), .ZN(new_n6339_));
  XOR2_X1    g03903(.A1(new_n6339_), .A2(pi0445), .Z(new_n6340_));
  XOR2_X1    g03904(.A1(new_n6340_), .A2(pi0448), .Z(new_n6341_));
  XOR2_X1    g03905(.A1(new_n6341_), .A2(new_n6331_), .Z(new_n6342_));
  NAND2_X1   g03906(.A1(new_n6342_), .A2(pi1199), .ZN(new_n6343_));
  AOI21_X1   g03907(.A1(new_n6321_), .A2(new_n6343_), .B(new_n6270_), .ZN(new_n6344_));
  OAI21_X1   g03908(.A1(new_n6344_), .A2(new_n6254_), .B(new_n6267_), .ZN(new_n6345_));
  INV_X1     g03909(.I(pi0285), .ZN(new_n6346_));
  INV_X1     g03910(.I(pi0289), .ZN(new_n6347_));
  NAND2_X1   g03911(.A1(new_n6346_), .A2(new_n6347_), .ZN(new_n6348_));
  NOR3_X1    g03912(.A1(new_n6348_), .A2(pi0286), .A3(pi0288), .ZN(new_n6349_));
  INV_X1     g03913(.I(new_n6349_), .ZN(new_n6350_));
  NAND3_X1   g03914(.A1(new_n6345_), .A2(po1038), .A3(new_n6350_), .ZN(new_n6351_));
  INV_X1     g03915(.I(pi0590), .ZN(new_n6352_));
  NOR2_X1    g03916(.A1(new_n6266_), .A2(new_n6352_), .ZN(new_n6353_));
  XOR2_X1    g03917(.A1(pi0335), .A2(pi0407), .Z(new_n6354_));
  INV_X1     g03918(.I(new_n6354_), .ZN(new_n6355_));
  INV_X1     g03919(.I(pi0463), .ZN(new_n6356_));
  NOR2_X1    g03920(.A1(new_n6356_), .A2(pi0413), .ZN(new_n6357_));
  INV_X1     g03921(.I(pi0413), .ZN(new_n6358_));
  NOR2_X1    g03922(.A1(new_n6358_), .A2(pi0463), .ZN(new_n6359_));
  OAI21_X1   g03923(.A1(new_n6357_), .A2(new_n6359_), .B(new_n6355_), .ZN(new_n6360_));
  XOR2_X1    g03924(.A1(pi0413), .A2(pi0463), .Z(new_n6361_));
  OAI21_X1   g03925(.A1(new_n6355_), .A2(new_n6361_), .B(new_n6360_), .ZN(new_n6362_));
  XOR2_X1    g03926(.A1(new_n6362_), .A2(pi0334), .Z(new_n6363_));
  XOR2_X1    g03927(.A1(new_n6363_), .A2(pi0393), .Z(new_n6364_));
  XNOR2_X1   g03928(.A1(pi0391), .A2(pi0392), .ZN(new_n6365_));
  INV_X1     g03929(.I(new_n6365_), .ZN(new_n6366_));
  XOR2_X1    g03930(.A1(pi0328), .A2(pi0394), .Z(new_n6367_));
  INV_X1     g03931(.I(pi0396), .ZN(new_n6368_));
  NAND2_X1   g03932(.A1(new_n6368_), .A2(pi0408), .ZN(new_n6369_));
  INV_X1     g03933(.I(pi0408), .ZN(new_n6370_));
  NAND2_X1   g03934(.A1(new_n6370_), .A2(pi0396), .ZN(new_n6371_));
  AOI21_X1   g03935(.A1(new_n6369_), .A2(new_n6371_), .B(new_n6367_), .ZN(new_n6372_));
  XNOR2_X1   g03936(.A1(pi0396), .A2(pi0408), .ZN(new_n6373_));
  AOI21_X1   g03937(.A1(new_n6367_), .A2(new_n6373_), .B(new_n6372_), .ZN(new_n6374_));
  XOR2_X1    g03938(.A1(pi0329), .A2(pi0395), .Z(new_n6375_));
  XOR2_X1    g03939(.A1(new_n6375_), .A2(pi0398), .Z(new_n6376_));
  XNOR2_X1   g03940(.A1(pi0399), .A2(pi0400), .ZN(new_n6377_));
  XOR2_X1    g03941(.A1(new_n6376_), .A2(new_n6377_), .Z(new_n6378_));
  XOR2_X1    g03942(.A1(new_n6378_), .A2(new_n6374_), .Z(new_n6379_));
  INV_X1     g03943(.I(pi1199), .ZN(new_n6380_));
  INV_X1     g03944(.I(new_n6270_), .ZN(new_n6381_));
  INV_X1     g03945(.I(pi0411), .ZN(new_n6382_));
  XNOR2_X1   g03946(.A1(pi0404), .A2(pi0412), .ZN(new_n6383_));
  NOR2_X1    g03947(.A1(pi0324), .A2(pi0456), .ZN(new_n6384_));
  INV_X1     g03948(.I(pi0324), .ZN(new_n6385_));
  INV_X1     g03949(.I(pi0456), .ZN(new_n6386_));
  NOR2_X1    g03950(.A1(new_n6385_), .A2(new_n6386_), .ZN(new_n6387_));
  OAI21_X1   g03951(.A1(new_n6387_), .A2(new_n6384_), .B(pi0319), .ZN(new_n6388_));
  INV_X1     g03952(.I(pi0319), .ZN(new_n6389_));
  NOR2_X1    g03953(.A1(new_n6386_), .A2(pi0324), .ZN(new_n6390_));
  NOR2_X1    g03954(.A1(new_n6385_), .A2(pi0456), .ZN(new_n6391_));
  OAI21_X1   g03955(.A1(new_n6390_), .A2(new_n6391_), .B(new_n6389_), .ZN(new_n6392_));
  NAND2_X1   g03956(.A1(new_n6388_), .A2(new_n6392_), .ZN(new_n6393_));
  XOR2_X1    g03957(.A1(new_n6393_), .A2(pi0397), .Z(new_n6394_));
  XOR2_X1    g03958(.A1(new_n6394_), .A2(new_n6383_), .Z(new_n6395_));
  XNOR2_X1   g03959(.A1(pi0390), .A2(pi0410), .ZN(new_n6396_));
  NOR2_X1    g03960(.A1(new_n6395_), .A2(new_n6396_), .ZN(new_n6397_));
  XOR2_X1    g03961(.A1(pi0390), .A2(pi0410), .Z(new_n6398_));
  INV_X1     g03962(.I(new_n6398_), .ZN(new_n6399_));
  AOI21_X1   g03963(.A1(new_n6395_), .A2(new_n6399_), .B(new_n6397_), .ZN(new_n6400_));
  OR2_X2     g03964(.A1(new_n6400_), .A2(new_n6382_), .Z(new_n6401_));
  NAND2_X1   g03965(.A1(new_n6400_), .A2(new_n6382_), .ZN(new_n6402_));
  NAND2_X1   g03966(.A1(new_n6401_), .A2(new_n6402_), .ZN(new_n6403_));
  INV_X1     g03967(.I(new_n6403_), .ZN(new_n6404_));
  OAI21_X1   g03968(.A1(new_n6404_), .A2(new_n6304_), .B(new_n6266_), .ZN(new_n6405_));
  NAND2_X1   g03969(.A1(new_n6403_), .A2(pi1196), .ZN(new_n6406_));
  XNOR2_X1   g03970(.A1(pi0318), .A2(pi0409), .ZN(new_n6407_));
  XNOR2_X1   g03971(.A1(pi0402), .A2(pi0406), .ZN(new_n6408_));
  XOR2_X1    g03972(.A1(pi0325), .A2(pi0405), .Z(new_n6409_));
  XOR2_X1    g03973(.A1(pi0326), .A2(pi0403), .Z(new_n6410_));
  XOR2_X1    g03974(.A1(new_n6409_), .A2(new_n6410_), .Z(new_n6411_));
  XOR2_X1    g03975(.A1(new_n6411_), .A2(pi0401), .Z(new_n6412_));
  XOR2_X1    g03976(.A1(new_n6412_), .A2(new_n6408_), .Z(new_n6413_));
  AND2_X2    g03977(.A1(new_n6413_), .A2(new_n6407_), .Z(new_n6414_));
  NOR2_X1    g03978(.A1(new_n6413_), .A2(new_n6407_), .ZN(new_n6415_));
  NOR2_X1    g03979(.A1(new_n6414_), .A2(new_n6415_), .ZN(new_n6416_));
  NOR2_X1    g03980(.A1(new_n6416_), .A2(new_n6265_), .ZN(new_n6417_));
  NAND4_X1   g03981(.A1(new_n6406_), .A2(pi0567), .A3(new_n6268_), .A4(new_n6417_), .ZN(new_n6418_));
  AND2_X2    g03982(.A1(new_n6418_), .A2(pi1199), .Z(new_n6419_));
  AOI22_X1   g03983(.A1(new_n6419_), .A2(new_n6381_), .B1(new_n6380_), .B2(new_n6405_), .ZN(new_n6420_));
  OAI21_X1   g03984(.A1(new_n6274_), .A2(new_n6270_), .B(new_n6420_), .ZN(new_n6421_));
  INV_X1     g03985(.I(pi0333), .ZN(new_n6422_));
  NOR2_X1    g03986(.A1(new_n6381_), .A2(new_n6273_), .ZN(new_n6423_));
  AOI21_X1   g03987(.A1(new_n6420_), .A2(new_n6273_), .B(new_n6423_), .ZN(new_n6424_));
  NOR2_X1    g03988(.A1(new_n6424_), .A2(new_n6422_), .ZN(new_n6425_));
  AOI21_X1   g03989(.A1(new_n6422_), .A2(new_n6420_), .B(new_n6425_), .ZN(new_n6426_));
  AOI21_X1   g03990(.A1(new_n6379_), .A2(new_n6421_), .B(new_n6426_), .ZN(new_n6427_));
  XOR2_X1    g03991(.A1(pi0391), .A2(pi0392), .Z(new_n6428_));
  INV_X1     g03992(.I(new_n6428_), .ZN(new_n6429_));
  NAND2_X1   g03993(.A1(new_n6424_), .A2(new_n6422_), .ZN(new_n6430_));
  NAND2_X1   g03994(.A1(new_n6430_), .A2(new_n6420_), .ZN(new_n6431_));
  AOI21_X1   g03995(.A1(new_n6379_), .A2(new_n6421_), .B(new_n6431_), .ZN(new_n6432_));
  AOI22_X1   g03996(.A1(new_n6427_), .A2(new_n6366_), .B1(new_n6429_), .B2(new_n6432_), .ZN(new_n6433_));
  NAND2_X1   g03997(.A1(new_n6433_), .A2(new_n6364_), .ZN(new_n6434_));
  INV_X1     g03998(.I(new_n6364_), .ZN(new_n6435_));
  AOI22_X1   g03999(.A1(new_n6427_), .A2(new_n6429_), .B1(new_n6366_), .B2(new_n6432_), .ZN(new_n6436_));
  NAND2_X1   g04000(.A1(new_n6436_), .A2(new_n6435_), .ZN(new_n6437_));
  AOI21_X1   g04001(.A1(new_n6434_), .A2(new_n6437_), .B(pi0590), .ZN(new_n6438_));
  OAI21_X1   g04002(.A1(new_n6438_), .A2(new_n6353_), .B(pi0591), .ZN(new_n6439_));
  INV_X1     g04003(.I(pi0591), .ZN(new_n6440_));
  XNOR2_X1   g04004(.A1(pi0357), .A2(pi0461), .ZN(new_n6441_));
  INV_X1     g04005(.I(new_n6441_), .ZN(new_n6442_));
  INV_X1     g04006(.I(pi0351), .ZN(new_n6443_));
  NOR2_X1    g04007(.A1(new_n6443_), .A2(new_n6380_), .ZN(new_n6444_));
  NAND2_X1   g04008(.A1(new_n6270_), .A2(new_n6444_), .ZN(new_n6445_));
  NOR2_X1    g04009(.A1(pi0345), .A2(pi0346), .ZN(new_n6446_));
  INV_X1     g04010(.I(pi0345), .ZN(new_n6447_));
  INV_X1     g04011(.I(pi0346), .ZN(new_n6448_));
  NOR2_X1    g04012(.A1(new_n6447_), .A2(new_n6448_), .ZN(new_n6449_));
  OAI21_X1   g04013(.A1(new_n6449_), .A2(new_n6446_), .B(pi0323), .ZN(new_n6450_));
  INV_X1     g04014(.I(pi0323), .ZN(new_n6451_));
  NOR2_X1    g04015(.A1(new_n6448_), .A2(pi0345), .ZN(new_n6452_));
  NOR2_X1    g04016(.A1(new_n6447_), .A2(pi0346), .ZN(new_n6453_));
  OAI21_X1   g04017(.A1(new_n6452_), .A2(new_n6453_), .B(new_n6451_), .ZN(new_n6454_));
  NAND2_X1   g04018(.A1(new_n6450_), .A2(new_n6454_), .ZN(new_n6455_));
  XNOR2_X1   g04019(.A1(pi0358), .A2(pi0450), .ZN(new_n6456_));
  XNOR2_X1   g04020(.A1(new_n6455_), .A2(new_n6456_), .ZN(new_n6457_));
  XOR2_X1    g04021(.A1(pi0327), .A2(pi0343), .Z(new_n6458_));
  INV_X1     g04022(.I(pi0344), .ZN(new_n6459_));
  NAND2_X1   g04023(.A1(new_n6459_), .A2(pi0362), .ZN(new_n6460_));
  INV_X1     g04024(.I(pi0362), .ZN(new_n6461_));
  NAND2_X1   g04025(.A1(new_n6461_), .A2(pi0344), .ZN(new_n6462_));
  AOI21_X1   g04026(.A1(new_n6460_), .A2(new_n6462_), .B(new_n6458_), .ZN(new_n6463_));
  XNOR2_X1   g04027(.A1(pi0344), .A2(pi0362), .ZN(new_n6464_));
  AOI21_X1   g04028(.A1(new_n6458_), .A2(new_n6464_), .B(new_n6463_), .ZN(new_n6465_));
  XOR2_X1    g04029(.A1(new_n6457_), .A2(new_n6465_), .Z(new_n6466_));
  NOR2_X1    g04030(.A1(new_n6466_), .A2(new_n6273_), .ZN(new_n6467_));
  NOR2_X1    g04031(.A1(pi0342), .A2(pi0460), .ZN(new_n6468_));
  INV_X1     g04032(.I(pi0342), .ZN(new_n6469_));
  INV_X1     g04033(.I(pi0460), .ZN(new_n6470_));
  NOR2_X1    g04034(.A1(new_n6469_), .A2(new_n6470_), .ZN(new_n6471_));
  OAI21_X1   g04035(.A1(new_n6471_), .A2(new_n6468_), .B(pi0320), .ZN(new_n6472_));
  INV_X1     g04036(.I(pi0320), .ZN(new_n6473_));
  NOR2_X1    g04037(.A1(new_n6470_), .A2(pi0342), .ZN(new_n6474_));
  NOR2_X1    g04038(.A1(new_n6469_), .A2(pi0460), .ZN(new_n6475_));
  OAI21_X1   g04039(.A1(new_n6474_), .A2(new_n6475_), .B(new_n6473_), .ZN(new_n6476_));
  NAND2_X1   g04040(.A1(new_n6472_), .A2(new_n6476_), .ZN(new_n6477_));
  INV_X1     g04041(.I(new_n6477_), .ZN(new_n6478_));
  XNOR2_X1   g04042(.A1(pi0361), .A2(pi0441), .ZN(new_n6479_));
  NOR2_X1    g04043(.A1(new_n6478_), .A2(new_n6479_), .ZN(new_n6480_));
  NAND2_X1   g04044(.A1(new_n6478_), .A2(new_n6479_), .ZN(new_n6481_));
  INV_X1     g04045(.I(new_n6481_), .ZN(new_n6482_));
  NOR2_X1    g04046(.A1(new_n6482_), .A2(new_n6480_), .ZN(new_n6483_));
  XOR2_X1    g04047(.A1(new_n6483_), .A2(pi0458), .Z(new_n6484_));
  INV_X1     g04048(.I(pi0355), .ZN(new_n6485_));
  NOR2_X1    g04049(.A1(pi0452), .A2(pi0455), .ZN(new_n6486_));
  INV_X1     g04050(.I(pi0452), .ZN(new_n6487_));
  INV_X1     g04051(.I(pi0455), .ZN(new_n6488_));
  NOR2_X1    g04052(.A1(new_n6487_), .A2(new_n6488_), .ZN(new_n6489_));
  NOR2_X1    g04053(.A1(new_n6489_), .A2(new_n6486_), .ZN(new_n6490_));
  XOR2_X1    g04054(.A1(new_n6490_), .A2(new_n6485_), .Z(new_n6491_));
  XOR2_X1    g04055(.A1(new_n6490_), .A2(pi0355), .Z(new_n6492_));
  INV_X1     g04056(.I(new_n6492_), .ZN(new_n6493_));
  NAND2_X1   g04057(.A1(new_n6484_), .A2(new_n6493_), .ZN(new_n6494_));
  OAI21_X1   g04058(.A1(new_n6484_), .A2(new_n6491_), .B(new_n6494_), .ZN(new_n6495_));
  INV_X1     g04059(.I(new_n6495_), .ZN(new_n6496_));
  NOR2_X1    g04060(.A1(new_n6496_), .A2(new_n6302_), .ZN(new_n6497_));
  INV_X1     g04061(.I(new_n6497_), .ZN(new_n6498_));
  XNOR2_X1   g04062(.A1(pi0321), .A2(pi0347), .ZN(new_n6499_));
  XNOR2_X1   g04063(.A1(pi0348), .A2(pi0349), .ZN(new_n6500_));
  INV_X1     g04064(.I(pi0359), .ZN(new_n6501_));
  NOR2_X1    g04065(.A1(new_n6501_), .A2(pi0322), .ZN(new_n6502_));
  INV_X1     g04066(.I(pi0322), .ZN(new_n6503_));
  NOR2_X1    g04067(.A1(new_n6503_), .A2(pi0359), .ZN(new_n6504_));
  OAI21_X1   g04068(.A1(new_n6502_), .A2(new_n6504_), .B(pi0315), .ZN(new_n6505_));
  INV_X1     g04069(.I(pi0315), .ZN(new_n6506_));
  NOR2_X1    g04070(.A1(pi0322), .A2(pi0359), .ZN(new_n6507_));
  NOR2_X1    g04071(.A1(new_n6503_), .A2(new_n6501_), .ZN(new_n6508_));
  OAI21_X1   g04072(.A1(new_n6508_), .A2(new_n6507_), .B(new_n6506_), .ZN(new_n6509_));
  NAND2_X1   g04073(.A1(new_n6509_), .A2(new_n6505_), .ZN(new_n6510_));
  XOR2_X1    g04074(.A1(new_n6510_), .A2(pi0316), .Z(new_n6511_));
  XOR2_X1    g04075(.A1(new_n6511_), .A2(new_n6500_), .Z(new_n6512_));
  XOR2_X1    g04076(.A1(new_n6512_), .A2(new_n6499_), .Z(new_n6513_));
  XOR2_X1    g04077(.A1(new_n6513_), .A2(pi0350), .Z(new_n6514_));
  NAND2_X1   g04078(.A1(new_n6498_), .A2(new_n6514_), .ZN(new_n6515_));
  INV_X1     g04079(.I(new_n6515_), .ZN(new_n6516_));
  NAND3_X1   g04080(.A1(new_n6516_), .A2(pi1198), .A3(new_n6271_), .ZN(new_n6517_));
  INV_X1     g04081(.I(pi0441), .ZN(new_n6518_));
  XOR2_X1    g04082(.A1(pi0361), .A2(pi0458), .Z(new_n6519_));
  NOR2_X1    g04083(.A1(new_n6491_), .A2(new_n6519_), .ZN(new_n6520_));
  AOI21_X1   g04084(.A1(new_n6493_), .A2(new_n6519_), .B(new_n6520_), .ZN(new_n6521_));
  XOR2_X1    g04085(.A1(new_n6521_), .A2(new_n6518_), .Z(new_n6522_));
  OAI21_X1   g04086(.A1(new_n6522_), .A2(pi0592), .B(new_n6266_), .ZN(new_n6523_));
  NOR2_X1    g04087(.A1(new_n6523_), .A2(new_n6478_), .ZN(new_n6524_));
  NOR2_X1    g04088(.A1(new_n6496_), .A2(pi0592), .ZN(new_n6525_));
  NAND2_X1   g04089(.A1(new_n6266_), .A2(new_n6478_), .ZN(new_n6526_));
  OAI21_X1   g04090(.A1(new_n6525_), .A2(new_n6526_), .B(pi1196), .ZN(new_n6527_));
  OAI21_X1   g04091(.A1(new_n6527_), .A2(new_n6524_), .B(new_n6274_), .ZN(new_n6528_));
  AOI21_X1   g04092(.A1(new_n6517_), .A2(new_n6528_), .B(new_n6467_), .ZN(new_n6529_));
  OAI21_X1   g04093(.A1(new_n6529_), .A2(pi0592), .B(new_n6266_), .ZN(new_n6530_));
  OAI21_X1   g04094(.A1(new_n6530_), .A2(new_n6444_), .B(new_n6445_), .ZN(new_n6531_));
  XOR2_X1    g04095(.A1(pi0357), .A2(pi0461), .Z(new_n6532_));
  INV_X1     g04096(.I(new_n6532_), .ZN(new_n6533_));
  NOR2_X1    g04097(.A1(new_n6380_), .A2(pi0351), .ZN(new_n6534_));
  NAND2_X1   g04098(.A1(new_n6270_), .A2(new_n6534_), .ZN(new_n6535_));
  OAI21_X1   g04099(.A1(new_n6530_), .A2(new_n6534_), .B(new_n6535_), .ZN(new_n6536_));
  AOI22_X1   g04100(.A1(new_n6442_), .A2(new_n6531_), .B1(new_n6536_), .B2(new_n6533_), .ZN(new_n6537_));
  XOR2_X1    g04101(.A1(pi0352), .A2(pi0353), .Z(new_n6538_));
  INV_X1     g04102(.I(new_n6538_), .ZN(new_n6539_));
  INV_X1     g04103(.I(pi0462), .ZN(new_n6540_));
  NOR2_X1    g04104(.A1(new_n6540_), .A2(pi0360), .ZN(new_n6541_));
  INV_X1     g04105(.I(pi0360), .ZN(new_n6542_));
  NOR2_X1    g04106(.A1(new_n6542_), .A2(pi0462), .ZN(new_n6543_));
  OAI21_X1   g04107(.A1(new_n6541_), .A2(new_n6543_), .B(new_n6539_), .ZN(new_n6544_));
  XOR2_X1    g04108(.A1(pi0360), .A2(pi0462), .Z(new_n6545_));
  OAI21_X1   g04109(.A1(new_n6539_), .A2(new_n6545_), .B(new_n6544_), .ZN(new_n6546_));
  XOR2_X1    g04110(.A1(new_n6546_), .A2(pi0354), .Z(new_n6547_));
  XOR2_X1    g04111(.A1(new_n6547_), .A2(pi0356), .Z(new_n6548_));
  NAND2_X1   g04112(.A1(new_n6537_), .A2(new_n6548_), .ZN(new_n6549_));
  INV_X1     g04113(.I(new_n6548_), .ZN(new_n6550_));
  AOI22_X1   g04114(.A1(new_n6442_), .A2(new_n6536_), .B1(new_n6531_), .B2(new_n6533_), .ZN(new_n6551_));
  NAND2_X1   g04115(.A1(new_n6551_), .A2(new_n6550_), .ZN(new_n6552_));
  AOI21_X1   g04116(.A1(new_n6549_), .A2(new_n6552_), .B(new_n6352_), .ZN(new_n6553_));
  XNOR2_X1   g04117(.A1(pi0338), .A2(pi0388), .ZN(new_n6554_));
  XOR2_X1    g04118(.A1(pi0337), .A2(pi0339), .Z(new_n6555_));
  XOR2_X1    g04119(.A1(new_n6555_), .A2(pi0380), .Z(new_n6556_));
  INV_X1     g04120(.I(pi0386), .ZN(new_n6557_));
  NOR2_X1    g04121(.A1(new_n6557_), .A2(pi0372), .ZN(new_n6558_));
  INV_X1     g04122(.I(pi0372), .ZN(new_n6559_));
  NOR2_X1    g04123(.A1(new_n6559_), .A2(pi0386), .ZN(new_n6560_));
  OAI21_X1   g04124(.A1(new_n6558_), .A2(new_n6560_), .B(pi0363), .ZN(new_n6561_));
  INV_X1     g04125(.I(pi0363), .ZN(new_n6562_));
  NOR2_X1    g04126(.A1(pi0372), .A2(pi0386), .ZN(new_n6563_));
  NOR2_X1    g04127(.A1(new_n6559_), .A2(new_n6557_), .ZN(new_n6564_));
  OAI21_X1   g04128(.A1(new_n6564_), .A2(new_n6563_), .B(new_n6562_), .ZN(new_n6565_));
  NAND2_X1   g04129(.A1(new_n6565_), .A2(new_n6561_), .ZN(new_n6566_));
  XOR2_X1    g04130(.A1(new_n6566_), .A2(pi0387), .Z(new_n6567_));
  XOR2_X1    g04131(.A1(new_n6567_), .A2(new_n6556_), .Z(new_n6568_));
  XOR2_X1    g04132(.A1(new_n6568_), .A2(new_n6554_), .Z(new_n6569_));
  INV_X1     g04133(.I(new_n6569_), .ZN(new_n6570_));
  NOR2_X1    g04134(.A1(new_n6570_), .A2(new_n6302_), .ZN(new_n6571_));
  XOR2_X1    g04135(.A1(pi0365), .A2(pi0447), .Z(new_n6572_));
  XOR2_X1    g04136(.A1(pi0336), .A2(pi0364), .Z(new_n6573_));
  INV_X1     g04137(.I(new_n6573_), .ZN(new_n6574_));
  INV_X1     g04138(.I(pi0383), .ZN(new_n6575_));
  NOR2_X1    g04139(.A1(new_n6575_), .A2(pi0366), .ZN(new_n6576_));
  INV_X1     g04140(.I(pi0366), .ZN(new_n6577_));
  NOR2_X1    g04141(.A1(new_n6577_), .A2(pi0383), .ZN(new_n6578_));
  OAI21_X1   g04142(.A1(new_n6576_), .A2(new_n6578_), .B(new_n6574_), .ZN(new_n6579_));
  XOR2_X1    g04143(.A1(pi0366), .A2(pi0383), .Z(new_n6580_));
  OAI21_X1   g04144(.A1(new_n6574_), .A2(new_n6580_), .B(new_n6579_), .ZN(new_n6581_));
  XOR2_X1    g04145(.A1(new_n6581_), .A2(new_n6572_), .Z(new_n6582_));
  INV_X1     g04146(.I(pi0367), .ZN(new_n6583_));
  XOR2_X1    g04147(.A1(pi0368), .A2(pi0389), .Z(new_n6584_));
  XOR2_X1    g04148(.A1(new_n6584_), .A2(new_n6583_), .Z(new_n6585_));
  XOR2_X1    g04149(.A1(new_n6584_), .A2(pi0367), .Z(new_n6586_));
  INV_X1     g04150(.I(new_n6586_), .ZN(new_n6587_));
  NAND2_X1   g04151(.A1(new_n6582_), .A2(new_n6587_), .ZN(new_n6588_));
  OAI21_X1   g04152(.A1(new_n6582_), .A2(new_n6585_), .B(new_n6588_), .ZN(new_n6589_));
  NAND2_X1   g04153(.A1(new_n6589_), .A2(pi1197), .ZN(new_n6590_));
  INV_X1     g04154(.I(new_n6590_), .ZN(new_n6591_));
  NOR2_X1    g04155(.A1(new_n6571_), .A2(new_n6591_), .ZN(new_n6592_));
  INV_X1     g04156(.I(new_n6592_), .ZN(new_n6593_));
  INV_X1     g04157(.I(pi0377), .ZN(new_n6594_));
  XNOR2_X1   g04158(.A1(pi0379), .A2(pi0382), .ZN(new_n6595_));
  XNOR2_X1   g04159(.A1(pi0381), .A2(pi0439), .ZN(new_n6596_));
  INV_X1     g04160(.I(pi0385), .ZN(new_n6597_));
  NOR2_X1    g04161(.A1(new_n6597_), .A2(pi0378), .ZN(new_n6598_));
  INV_X1     g04162(.I(pi0378), .ZN(new_n6599_));
  NOR2_X1    g04163(.A1(new_n6599_), .A2(pi0385), .ZN(new_n6600_));
  OAI21_X1   g04164(.A1(new_n6598_), .A2(new_n6600_), .B(pi0317), .ZN(new_n6601_));
  INV_X1     g04165(.I(pi0317), .ZN(new_n6602_));
  NOR2_X1    g04166(.A1(pi0378), .A2(pi0385), .ZN(new_n6603_));
  NOR2_X1    g04167(.A1(new_n6599_), .A2(new_n6597_), .ZN(new_n6604_));
  OAI21_X1   g04168(.A1(new_n6604_), .A2(new_n6603_), .B(new_n6602_), .ZN(new_n6605_));
  NAND2_X1   g04169(.A1(new_n6605_), .A2(new_n6601_), .ZN(new_n6606_));
  XOR2_X1    g04170(.A1(new_n6606_), .A2(pi0376), .Z(new_n6607_));
  XOR2_X1    g04171(.A1(new_n6607_), .A2(new_n6596_), .Z(new_n6608_));
  XOR2_X1    g04172(.A1(new_n6608_), .A2(new_n6595_), .Z(new_n6609_));
  XOR2_X1    g04173(.A1(new_n6609_), .A2(new_n6594_), .Z(new_n6610_));
  NOR2_X1    g04174(.A1(new_n6593_), .A2(new_n6610_), .ZN(new_n6611_));
  OAI21_X1   g04175(.A1(new_n6611_), .A2(new_n6268_), .B(new_n6266_), .ZN(new_n6612_));
  NAND2_X1   g04176(.A1(new_n6612_), .A2(pi1199), .ZN(new_n6613_));
  OAI21_X1   g04177(.A1(new_n6268_), .A2(new_n6592_), .B(new_n6613_), .ZN(new_n6614_));
  NOR2_X1    g04178(.A1(new_n6614_), .A2(new_n6381_), .ZN(new_n6615_));
  XNOR2_X1   g04179(.A1(pi0369), .A2(pi0370), .ZN(new_n6616_));
  XOR2_X1    g04180(.A1(pi0371), .A2(pi0374), .Z(new_n6617_));
  XNOR2_X1   g04181(.A1(pi0369), .A2(pi0370), .ZN(new_n6618_));
  NOR2_X1    g04182(.A1(new_n6618_), .A2(new_n6617_), .ZN(new_n6619_));
  AOI21_X1   g04183(.A1(new_n6616_), .A2(new_n6617_), .B(new_n6619_), .ZN(new_n6620_));
  NOR2_X1    g04184(.A1(pi0440), .A2(pi0442), .ZN(new_n6621_));
  INV_X1     g04185(.I(pi0440), .ZN(new_n6622_));
  INV_X1     g04186(.I(pi0442), .ZN(new_n6623_));
  NOR2_X1    g04187(.A1(new_n6622_), .A2(new_n6623_), .ZN(new_n6624_));
  OAI21_X1   g04188(.A1(new_n6624_), .A2(new_n6621_), .B(pi0384), .ZN(new_n6625_));
  INV_X1     g04189(.I(pi0384), .ZN(new_n6626_));
  NOR2_X1    g04190(.A1(new_n6623_), .A2(pi0440), .ZN(new_n6627_));
  NOR2_X1    g04191(.A1(new_n6622_), .A2(pi0442), .ZN(new_n6628_));
  OAI21_X1   g04192(.A1(new_n6627_), .A2(new_n6628_), .B(new_n6626_), .ZN(new_n6629_));
  NAND2_X1   g04193(.A1(new_n6625_), .A2(new_n6629_), .ZN(new_n6630_));
  INV_X1     g04194(.I(new_n6630_), .ZN(new_n6631_));
  XNOR2_X1   g04195(.A1(pi0373), .A2(pi0375), .ZN(new_n6632_));
  NOR2_X1    g04196(.A1(new_n6631_), .A2(new_n6632_), .ZN(new_n6633_));
  INV_X1     g04197(.I(new_n6633_), .ZN(new_n6634_));
  NAND2_X1   g04198(.A1(new_n6631_), .A2(new_n6632_), .ZN(new_n6635_));
  NAND2_X1   g04199(.A1(new_n6634_), .A2(new_n6635_), .ZN(new_n6636_));
  XNOR2_X1   g04200(.A1(new_n6636_), .A2(new_n6620_), .ZN(new_n6637_));
  OAI21_X1   g04201(.A1(new_n6274_), .A2(new_n6637_), .B(new_n6615_), .ZN(new_n6638_));
  AND3_X2    g04202(.A1(new_n6638_), .A2(new_n6352_), .A3(new_n6272_), .Z(new_n6639_));
  OAI21_X1   g04203(.A1(new_n6553_), .A2(new_n6639_), .B(new_n6440_), .ZN(new_n6640_));
  NAND2_X1   g04204(.A1(new_n6439_), .A2(new_n6640_), .ZN(new_n6641_));
  AOI21_X1   g04205(.A1(new_n6641_), .A2(new_n6251_), .B(new_n6351_), .ZN(new_n6642_));
  INV_X1     g04206(.I(po1038), .ZN(new_n6643_));
  INV_X1     g04207(.I(new_n5305_), .ZN(new_n6644_));
  NOR2_X1    g04208(.A1(new_n6644_), .A2(pi0074), .ZN(new_n6645_));
  NOR2_X1    g04209(.A1(new_n6269_), .A2(new_n6645_), .ZN(new_n6646_));
  INV_X1     g04210(.I(new_n6646_), .ZN(new_n6647_));
  INV_X1     g04211(.I(new_n6645_), .ZN(new_n6648_));
  NOR2_X1    g04212(.A1(new_n2575_), .A2(pi0075), .ZN(new_n6649_));
  INV_X1     g04213(.I(new_n6649_), .ZN(new_n6650_));
  NAND2_X1   g04214(.A1(new_n2531_), .A2(po0740), .ZN(new_n6651_));
  AOI21_X1   g04215(.A1(new_n6651_), .A2(pi0087), .B(new_n6650_), .ZN(new_n6652_));
  NOR2_X1    g04216(.A1(new_n3044_), .A2(pi0122), .ZN(new_n6653_));
  INV_X1     g04217(.I(new_n6653_), .ZN(new_n6654_));
  NOR2_X1    g04218(.A1(new_n6654_), .A2(new_n3082_), .ZN(new_n6655_));
  INV_X1     g04219(.I(new_n6655_), .ZN(new_n6656_));
  NAND2_X1   g04220(.A1(new_n5611_), .A2(new_n2746_), .ZN(new_n6657_));
  NAND2_X1   g04221(.A1(new_n6657_), .A2(pi0096), .ZN(new_n6658_));
  INV_X1     g04222(.I(new_n6658_), .ZN(new_n6659_));
  NOR2_X1    g04223(.A1(new_n6659_), .A2(new_n2526_), .ZN(new_n6660_));
  INV_X1     g04224(.I(new_n6660_), .ZN(new_n6661_));
  NOR2_X1    g04225(.A1(new_n2739_), .A2(pi0841), .ZN(new_n6662_));
  AOI21_X1   g04226(.A1(new_n6662_), .A2(pi0090), .B(pi0093), .ZN(new_n6663_));
  INV_X1     g04227(.I(new_n6663_), .ZN(new_n6664_));
  NOR2_X1    g04228(.A1(new_n5378_), .A2(pi0070), .ZN(new_n6665_));
  AOI21_X1   g04229(.A1(new_n6664_), .A2(new_n6665_), .B(pi0051), .ZN(new_n6666_));
  NOR2_X1    g04230(.A1(pi0050), .A2(pi0077), .ZN(new_n6667_));
  INV_X1     g04231(.I(new_n6667_), .ZN(new_n6668_));
  NOR2_X1    g04232(.A1(new_n6668_), .A2(pi0094), .ZN(new_n6669_));
  INV_X1     g04233(.I(new_n6669_), .ZN(new_n6670_));
  INV_X1     g04234(.I(new_n2515_), .ZN(new_n6671_));
  NOR2_X1    g04235(.A1(new_n6671_), .A2(pi0088), .ZN(new_n6672_));
  INV_X1     g04236(.I(new_n6672_), .ZN(new_n6673_));
  NOR4_X1    g04237(.A1(new_n2870_), .A2(new_n2887_), .A3(new_n6670_), .A4(new_n6673_), .ZN(new_n6674_));
  OAI21_X1   g04238(.A1(new_n6674_), .A2(pi0097), .B(new_n2786_), .ZN(new_n6675_));
  NOR2_X1    g04239(.A1(new_n2741_), .A2(pi0035), .ZN(new_n6676_));
  INV_X1     g04240(.I(new_n6676_), .ZN(new_n6677_));
  NOR2_X1    g04241(.A1(new_n6677_), .A2(pi0070), .ZN(new_n6678_));
  INV_X1     g04242(.I(new_n6678_), .ZN(new_n6679_));
  OAI21_X1   g04243(.A1(new_n6675_), .A2(new_n6679_), .B(new_n6666_), .ZN(new_n6680_));
  OAI21_X1   g04244(.A1(new_n2744_), .A2(new_n2831_), .B(new_n6680_), .ZN(new_n6681_));
  AND2_X2    g04245(.A1(new_n6681_), .A2(new_n2742_), .Z(new_n6682_));
  NOR3_X1    g04246(.A1(new_n6682_), .A2(new_n6656_), .A3(new_n6661_), .ZN(new_n6683_));
  NOR2_X1    g04247(.A1(new_n2526_), .A2(pi0096), .ZN(new_n6684_));
  INV_X1     g04248(.I(new_n6684_), .ZN(new_n6685_));
  NOR2_X1    g04249(.A1(new_n6681_), .A2(new_n6685_), .ZN(new_n6686_));
  INV_X1     g04250(.I(new_n6686_), .ZN(new_n6687_));
  NOR2_X1    g04251(.A1(new_n6687_), .A2(new_n5331_), .ZN(new_n6688_));
  AOI21_X1   g04252(.A1(new_n6654_), .A2(new_n6688_), .B(new_n6683_), .ZN(new_n6689_));
  NOR2_X1    g04253(.A1(new_n6689_), .A2(pi1093), .ZN(new_n6690_));
  OAI21_X1   g04254(.A1(new_n6690_), .A2(pi0087), .B(new_n6652_), .ZN(new_n6691_));
  AOI21_X1   g04255(.A1(new_n6691_), .A2(new_n6255_), .B(new_n6648_), .ZN(new_n6692_));
  NOR2_X1    g04256(.A1(new_n2690_), .A2(new_n2628_), .ZN(new_n6693_));
  NOR2_X1    g04257(.A1(new_n2669_), .A2(pi0299), .ZN(new_n6694_));
  NOR2_X1    g04258(.A1(new_n6693_), .A2(new_n6694_), .ZN(new_n6695_));
  INV_X1     g04259(.I(new_n6695_), .ZN(new_n6696_));
  NOR2_X1    g04260(.A1(new_n5437_), .A2(new_n5666_), .ZN(new_n6697_));
  INV_X1     g04261(.I(new_n6697_), .ZN(new_n6698_));
  NOR2_X1    g04262(.A1(new_n6696_), .A2(new_n6698_), .ZN(new_n6699_));
  NOR2_X1    g04263(.A1(new_n6699_), .A2(new_n2659_), .ZN(new_n6700_));
  INV_X1     g04264(.I(new_n6700_), .ZN(new_n6701_));
  AOI21_X1   g04265(.A1(new_n6701_), .A2(new_n6264_), .B(new_n3465_), .ZN(new_n6702_));
  NOR2_X1    g04266(.A1(new_n6656_), .A2(new_n3041_), .ZN(new_n6703_));
  NOR2_X1    g04267(.A1(new_n5323_), .A2(new_n3024_), .ZN(new_n6704_));
  INV_X1     g04268(.I(new_n6704_), .ZN(new_n6705_));
  NOR3_X1    g04269(.A1(new_n2530_), .A2(pi0024), .A3(new_n2704_), .ZN(new_n6706_));
  INV_X1     g04270(.I(new_n6706_), .ZN(new_n6707_));
  NOR2_X1    g04271(.A1(new_n6707_), .A2(new_n6705_), .ZN(new_n6708_));
  AOI21_X1   g04272(.A1(new_n6708_), .A2(new_n6703_), .B(new_n3022_), .ZN(new_n6709_));
  NOR2_X1    g04273(.A1(new_n6709_), .A2(new_n6701_), .ZN(new_n6710_));
  OAI21_X1   g04274(.A1(pi1091), .A2(new_n6262_), .B(new_n6710_), .ZN(new_n6711_));
  NOR2_X1    g04275(.A1(new_n3024_), .A2(new_n3041_), .ZN(new_n6712_));
  INV_X1     g04276(.I(new_n6712_), .ZN(new_n6713_));
  INV_X1     g04277(.I(pi0122), .ZN(new_n6714_));
  NOR2_X1    g04278(.A1(new_n2834_), .A2(new_n2526_), .ZN(new_n6715_));
  INV_X1     g04279(.I(new_n6715_), .ZN(new_n6716_));
  NOR2_X1    g04280(.A1(new_n6666_), .A2(new_n6716_), .ZN(new_n6717_));
  INV_X1     g04281(.I(new_n2839_), .ZN(new_n6718_));
  NOR2_X1    g04282(.A1(new_n6718_), .A2(pi0024), .ZN(new_n6719_));
  INV_X1     g04283(.I(new_n6719_), .ZN(new_n6720_));
  NAND4_X1   g04284(.A1(new_n2734_), .A2(new_n2511_), .A3(pi0097), .A4(new_n2849_), .ZN(new_n6721_));
  NOR2_X1    g04285(.A1(new_n2860_), .A2(new_n6721_), .ZN(new_n6722_));
  INV_X1     g04286(.I(new_n6722_), .ZN(new_n6723_));
  OAI21_X1   g04287(.A1(new_n6723_), .A2(pi0091), .B(new_n6720_), .ZN(new_n6724_));
  NAND3_X1   g04288(.A1(new_n6724_), .A2(new_n2520_), .A3(new_n6665_), .ZN(new_n6725_));
  AOI21_X1   g04289(.A1(new_n6725_), .A2(new_n6666_), .B(new_n2832_), .ZN(new_n6726_));
  NOR2_X1    g04290(.A1(new_n6726_), .A2(pi0096), .ZN(new_n6727_));
  NOR2_X1    g04291(.A1(new_n6661_), .A2(new_n3084_), .ZN(new_n6728_));
  INV_X1     g04292(.I(new_n6728_), .ZN(new_n6729_));
  INV_X1     g04293(.I(new_n6717_), .ZN(new_n6730_));
  NOR2_X1    g04294(.A1(new_n6730_), .A2(new_n6259_), .ZN(new_n6731_));
  INV_X1     g04295(.I(new_n6731_), .ZN(new_n6732_));
  OAI22_X1   g04296(.A1(new_n6732_), .A2(pi0829), .B1(new_n6727_), .B2(new_n6729_), .ZN(new_n6733_));
  NOR2_X1    g04297(.A1(new_n5331_), .A2(new_n6714_), .ZN(new_n6734_));
  AOI22_X1   g04298(.A1(new_n6733_), .A2(new_n6714_), .B1(new_n6717_), .B2(new_n6734_), .ZN(new_n6735_));
  NOR2_X1    g04299(.A1(new_n6735_), .A2(new_n6713_), .ZN(new_n6736_));
  OR3_X2     g04300(.A1(new_n6690_), .A2(new_n3022_), .A3(new_n6736_), .Z(new_n6737_));
  NAND2_X1   g04301(.A1(new_n6737_), .A2(new_n2627_), .ZN(new_n6738_));
  NOR2_X1    g04302(.A1(new_n6690_), .A2(pi1091), .ZN(new_n6739_));
  NOR2_X1    g04303(.A1(new_n6261_), .A2(pi0122), .ZN(new_n6740_));
  NOR2_X1    g04304(.A1(new_n6732_), .A2(new_n6714_), .ZN(new_n6741_));
  OAI21_X1   g04305(.A1(new_n6741_), .A2(new_n6740_), .B(pi1093), .ZN(new_n6742_));
  AOI21_X1   g04306(.A1(new_n6739_), .A2(new_n6742_), .B(new_n6738_), .ZN(new_n6743_));
  NOR2_X1    g04307(.A1(new_n5082_), .A2(pi0223), .ZN(new_n6744_));
  INV_X1     g04308(.I(new_n5449_), .ZN(new_n6745_));
  NOR2_X1    g04309(.A1(new_n3043_), .A2(new_n3022_), .ZN(new_n6746_));
  INV_X1     g04310(.I(new_n6746_), .ZN(new_n6747_));
  NOR3_X1    g04311(.A1(new_n5527_), .A2(new_n3024_), .A3(new_n3047_), .ZN(new_n6748_));
  INV_X1     g04312(.I(new_n6748_), .ZN(new_n6749_));
  NOR2_X1    g04313(.A1(new_n6749_), .A2(new_n6747_), .ZN(new_n6750_));
  INV_X1     g04314(.I(new_n6750_), .ZN(new_n6751_));
  NOR2_X1    g04315(.A1(new_n6751_), .A2(new_n6745_), .ZN(new_n6752_));
  INV_X1     g04316(.I(new_n6752_), .ZN(new_n6753_));
  AOI21_X1   g04317(.A1(new_n6753_), .A2(new_n6265_), .B(new_n5445_), .ZN(new_n6754_));
  NOR2_X1    g04318(.A1(new_n6751_), .A2(new_n5413_), .ZN(new_n6755_));
  INV_X1     g04319(.I(new_n6755_), .ZN(new_n6756_));
  AOI21_X1   g04320(.A1(new_n6756_), .A2(new_n6265_), .B(new_n5446_), .ZN(new_n6757_));
  OAI21_X1   g04321(.A1(new_n6754_), .A2(new_n6757_), .B(new_n6744_), .ZN(new_n6758_));
  INV_X1     g04322(.I(new_n6744_), .ZN(new_n6759_));
  AOI21_X1   g04323(.A1(new_n6264_), .A2(new_n6759_), .B(pi0299), .ZN(new_n6760_));
  NOR2_X1    g04324(.A1(new_n5550_), .A2(pi0216), .ZN(new_n6761_));
  INV_X1     g04325(.I(new_n6761_), .ZN(new_n6762_));
  OAI21_X1   g04326(.A1(new_n6752_), .A2(new_n6264_), .B(new_n5422_), .ZN(new_n6763_));
  INV_X1     g04327(.I(new_n5422_), .ZN(new_n6764_));
  OAI21_X1   g04328(.A1(new_n6755_), .A2(new_n6264_), .B(new_n6764_), .ZN(new_n6765_));
  AOI21_X1   g04329(.A1(new_n6763_), .A2(new_n6765_), .B(new_n6762_), .ZN(new_n6766_));
  OAI21_X1   g04330(.A1(new_n6265_), .A2(new_n6761_), .B(pi0299), .ZN(new_n6767_));
  OAI21_X1   g04331(.A1(new_n6766_), .A2(new_n6767_), .B(pi0039), .ZN(new_n6768_));
  AOI21_X1   g04332(.A1(new_n6758_), .A2(new_n6760_), .B(new_n6768_), .ZN(new_n6769_));
  NOR3_X1    g04333(.A1(new_n6743_), .A2(pi0038), .A3(new_n6769_), .ZN(new_n6770_));
  NOR2_X1    g04334(.A1(new_n6264_), .A2(new_n3265_), .ZN(new_n6771_));
  OAI21_X1   g04335(.A1(new_n6770_), .A2(new_n6771_), .B(new_n2702_), .ZN(new_n6772_));
  NOR2_X1    g04336(.A1(new_n6264_), .A2(new_n2702_), .ZN(new_n6773_));
  NOR2_X1    g04337(.A1(new_n6699_), .A2(new_n2458_), .ZN(new_n6774_));
  NOR3_X1    g04338(.A1(new_n6705_), .A2(new_n2530_), .A3(new_n6656_), .ZN(new_n6775_));
  NAND2_X1   g04339(.A1(new_n6775_), .A2(new_n3080_), .ZN(new_n6776_));
  INV_X1     g04340(.I(new_n6776_), .ZN(new_n6777_));
  NAND3_X1   g04341(.A1(new_n6777_), .A2(new_n2572_), .A3(new_n6774_), .ZN(new_n6778_));
  AOI21_X1   g04342(.A1(new_n6778_), .A2(new_n6773_), .B(pi0087), .ZN(new_n6779_));
  NAND2_X1   g04343(.A1(new_n6772_), .A2(new_n6779_), .ZN(new_n6780_));
  NOR2_X1    g04344(.A1(new_n5532_), .A2(new_n3041_), .ZN(new_n6781_));
  NOR3_X1    g04345(.A1(new_n2530_), .A2(new_n5331_), .A3(new_n6781_), .ZN(new_n6782_));
  OR2_X2     g04346(.A1(new_n6782_), .A2(new_n3022_), .Z(new_n6783_));
  NAND2_X1   g04347(.A1(new_n6651_), .A2(new_n3022_), .ZN(new_n6784_));
  INV_X1     g04348(.I(new_n6784_), .ZN(new_n6785_));
  NOR2_X1    g04349(.A1(new_n2530_), .A2(new_n6259_), .ZN(new_n6786_));
  AOI21_X1   g04350(.A1(new_n6786_), .A2(pi0122), .B(new_n6740_), .ZN(new_n6787_));
  OAI21_X1   g04351(.A1(new_n6787_), .A2(new_n3041_), .B(new_n6785_), .ZN(new_n6788_));
  NAND3_X1   g04352(.A1(new_n6788_), .A2(new_n3272_), .A3(new_n6783_), .ZN(new_n6789_));
  NAND2_X1   g04353(.A1(new_n6789_), .A2(new_n6265_), .ZN(new_n6790_));
  AOI21_X1   g04354(.A1(new_n6790_), .A2(pi0087), .B(pi0075), .ZN(new_n6791_));
  AOI22_X1   g04355(.A1(new_n6780_), .A2(new_n6791_), .B1(new_n6702_), .B2(new_n6711_), .ZN(new_n6792_));
  OAI21_X1   g04356(.A1(new_n6792_), .A2(new_n6255_), .B(new_n6692_), .ZN(new_n6793_));
  NAND2_X1   g04357(.A1(new_n6793_), .A2(new_n6647_), .ZN(new_n6794_));
  AOI21_X1   g04358(.A1(new_n6794_), .A2(new_n6254_), .B(new_n6349_), .ZN(new_n6795_));
  NOR2_X1    g04359(.A1(new_n6794_), .A2(new_n6268_), .ZN(new_n6796_));
  NAND3_X1   g04360(.A1(new_n6708_), .A2(pi1091), .A3(new_n6655_), .ZN(new_n6797_));
  NOR2_X1    g04361(.A1(new_n6797_), .A2(new_n3041_), .ZN(new_n6798_));
  AOI21_X1   g04362(.A1(new_n6798_), .A2(new_n6700_), .B(new_n3465_), .ZN(new_n6799_));
  NOR2_X1    g04363(.A1(new_n3458_), .A2(pi0100), .ZN(new_n6800_));
  INV_X1     g04364(.I(new_n6800_), .ZN(new_n6801_));
  NOR2_X1    g04365(.A1(new_n6801_), .A2(new_n2573_), .ZN(new_n6802_));
  NAND3_X1   g04366(.A1(new_n6783_), .A2(new_n6784_), .A3(new_n6802_), .ZN(new_n6803_));
  NAND2_X1   g04367(.A1(new_n6803_), .A2(new_n3465_), .ZN(new_n6804_));
  NOR2_X1    g04368(.A1(new_n6751_), .A2(new_n5451_), .ZN(new_n6805_));
  NOR2_X1    g04369(.A1(new_n5525_), .A2(pi0299), .ZN(new_n6806_));
  NAND2_X1   g04370(.A1(new_n6805_), .A2(new_n6806_), .ZN(new_n6807_));
  OAI21_X1   g04371(.A1(new_n6807_), .A2(pi0224), .B(pi0039), .ZN(new_n6808_));
  INV_X1     g04372(.I(new_n5423_), .ZN(new_n6809_));
  NOR2_X1    g04373(.A1(new_n6762_), .A2(new_n2628_), .ZN(new_n6810_));
  INV_X1     g04374(.I(new_n6810_), .ZN(new_n6811_));
  NOR3_X1    g04375(.A1(new_n6751_), .A2(new_n6809_), .A3(new_n6811_), .ZN(new_n6812_));
  OAI21_X1   g04376(.A1(new_n6808_), .A2(new_n6812_), .B(new_n3265_), .ZN(new_n6813_));
  INV_X1     g04377(.I(new_n6739_), .ZN(new_n6814_));
  NAND2_X1   g04378(.A1(new_n6737_), .A2(new_n6814_), .ZN(new_n6815_));
  AOI21_X1   g04379(.A1(new_n6815_), .A2(new_n2627_), .B(new_n6813_), .ZN(new_n6816_));
  NOR2_X1    g04380(.A1(new_n6816_), .A2(pi0100), .ZN(new_n6817_));
  INV_X1     g04381(.I(new_n6817_), .ZN(new_n6818_));
  INV_X1     g04382(.I(new_n6774_), .ZN(new_n6819_));
  NOR2_X1    g04383(.A1(new_n6819_), .A2(new_n2573_), .ZN(new_n6820_));
  AOI21_X1   g04384(.A1(new_n6777_), .A2(new_n6820_), .B(new_n2702_), .ZN(new_n6821_));
  NOR2_X1    g04385(.A1(new_n6821_), .A2(pi0087), .ZN(new_n6822_));
  AOI21_X1   g04386(.A1(new_n6818_), .A2(new_n6822_), .B(new_n6804_), .ZN(new_n6823_));
  OAI21_X1   g04387(.A1(new_n6823_), .A2(new_n6799_), .B(pi0567), .ZN(new_n6824_));
  NAND2_X1   g04388(.A1(new_n6824_), .A2(new_n6692_), .ZN(new_n6825_));
  INV_X1     g04389(.I(new_n6825_), .ZN(new_n6826_));
  NOR2_X1    g04390(.A1(new_n6826_), .A2(pi0592), .ZN(new_n6827_));
  NOR2_X1    g04391(.A1(new_n6796_), .A2(new_n6827_), .ZN(new_n6828_));
  XOR2_X1    g04392(.A1(pi0436), .A2(pi0444), .Z(new_n6829_));
  INV_X1     g04393(.I(new_n6829_), .ZN(new_n6830_));
  XOR2_X1    g04394(.A1(new_n6316_), .A2(new_n6830_), .Z(new_n6831_));
  INV_X1     g04395(.I(new_n6831_), .ZN(new_n6832_));
  NAND2_X1   g04396(.A1(new_n6268_), .A2(pi0443), .ZN(new_n6833_));
  NOR2_X1    g04397(.A1(new_n6825_), .A2(new_n6833_), .ZN(new_n6834_));
  AOI21_X1   g04398(.A1(new_n6794_), .A2(new_n6833_), .B(new_n6834_), .ZN(new_n6835_));
  OAI21_X1   g04399(.A1(new_n6835_), .A2(new_n6832_), .B(pi1196), .ZN(new_n6836_));
  NOR2_X1    g04400(.A1(pi0443), .A2(pi0592), .ZN(new_n6837_));
  INV_X1     g04401(.I(new_n6837_), .ZN(new_n6838_));
  NOR2_X1    g04402(.A1(new_n6825_), .A2(new_n6838_), .ZN(new_n6839_));
  AOI21_X1   g04403(.A1(new_n6794_), .A2(new_n6838_), .B(new_n6839_), .ZN(new_n6840_));
  NOR2_X1    g04404(.A1(new_n6840_), .A2(new_n6831_), .ZN(new_n6841_));
  NOR2_X1    g04405(.A1(new_n6836_), .A2(new_n6841_), .ZN(new_n6842_));
  NOR2_X1    g04406(.A1(new_n6794_), .A2(pi1196), .ZN(new_n6843_));
  NOR3_X1    g04407(.A1(new_n6842_), .A2(new_n6301_), .A3(new_n6843_), .ZN(new_n6844_));
  AOI21_X1   g04408(.A1(new_n6301_), .A2(new_n6828_), .B(new_n6844_), .ZN(new_n6845_));
  AOI21_X1   g04409(.A1(new_n6845_), .A2(new_n6380_), .B(new_n6254_), .ZN(new_n6846_));
  INV_X1     g04410(.I(new_n6828_), .ZN(new_n6847_));
  XOR2_X1    g04411(.A1(pi0427), .A2(pi0428), .Z(new_n6848_));
  INV_X1     g04412(.I(new_n6848_), .ZN(new_n6849_));
  XNOR2_X1   g04413(.A1(pi0427), .A2(pi0428), .ZN(new_n6850_));
  INV_X1     g04414(.I(new_n6850_), .ZN(new_n6851_));
  AOI22_X1   g04415(.A1(new_n6845_), .A2(new_n6851_), .B1(new_n6847_), .B2(new_n6849_), .ZN(new_n6852_));
  XOR2_X1    g04416(.A1(pi0426), .A2(pi0430), .Z(new_n6853_));
  INV_X1     g04417(.I(new_n6853_), .ZN(new_n6854_));
  OAI22_X1   g04418(.A1(new_n6845_), .A2(new_n6848_), .B1(new_n6847_), .B2(new_n6850_), .ZN(new_n6855_));
  XNOR2_X1   g04419(.A1(pi0426), .A2(pi0430), .ZN(new_n6856_));
  INV_X1     g04420(.I(new_n6856_), .ZN(new_n6857_));
  AOI22_X1   g04421(.A1(new_n6852_), .A2(new_n6854_), .B1(new_n6855_), .B2(new_n6857_), .ZN(new_n6858_));
  INV_X1     g04422(.I(pi0445), .ZN(new_n6859_));
  XOR2_X1    g04423(.A1(new_n6331_), .A2(pi0448), .Z(new_n6860_));
  XOR2_X1    g04424(.A1(new_n6860_), .A2(new_n6859_), .Z(new_n6861_));
  AND2_X2    g04425(.A1(new_n6858_), .A2(new_n6861_), .Z(new_n6862_));
  NAND2_X1   g04426(.A1(new_n6855_), .A2(new_n6854_), .ZN(new_n6863_));
  NAND2_X1   g04427(.A1(new_n6852_), .A2(new_n6857_), .ZN(new_n6864_));
  NAND2_X1   g04428(.A1(new_n6864_), .A2(new_n6863_), .ZN(new_n6865_));
  NOR2_X1    g04429(.A1(new_n6865_), .A2(new_n6861_), .ZN(new_n6866_));
  OAI21_X1   g04430(.A1(new_n6862_), .A2(new_n6866_), .B(pi1199), .ZN(new_n6867_));
  NAND2_X1   g04431(.A1(new_n6867_), .A2(new_n6846_), .ZN(new_n6868_));
  INV_X1     g04432(.I(new_n6799_), .ZN(new_n6869_));
  NOR2_X1    g04433(.A1(new_n3041_), .A2(pi1091), .ZN(new_n6870_));
  INV_X1     g04434(.I(new_n6870_), .ZN(new_n6871_));
  NOR2_X1    g04435(.A1(new_n6782_), .A2(new_n6870_), .ZN(new_n6872_));
  INV_X1     g04436(.I(new_n6872_), .ZN(new_n6873_));
  OAI21_X1   g04437(.A1(new_n6786_), .A2(new_n6871_), .B(new_n6873_), .ZN(new_n6874_));
  OAI21_X1   g04438(.A1(new_n6874_), .A2(new_n3273_), .B(pi0087), .ZN(new_n6875_));
  INV_X1     g04439(.I(new_n6813_), .ZN(new_n6876_));
  OAI21_X1   g04440(.A1(new_n6736_), .A2(new_n3022_), .B(new_n6876_), .ZN(new_n6877_));
  NOR3_X1    g04441(.A1(new_n6877_), .A2(new_n5531_), .A3(new_n6730_), .ZN(new_n6878_));
  INV_X1     g04442(.I(new_n6878_), .ZN(new_n6879_));
  AOI21_X1   g04443(.A1(new_n6817_), .A2(new_n6879_), .B(new_n6821_), .ZN(new_n6880_));
  OAI21_X1   g04444(.A1(new_n6880_), .A2(pi0087), .B(new_n6875_), .ZN(new_n6881_));
  NAND2_X1   g04445(.A1(new_n6881_), .A2(new_n3465_), .ZN(new_n6882_));
  NAND2_X1   g04446(.A1(new_n6882_), .A2(new_n6869_), .ZN(new_n6883_));
  NAND2_X1   g04447(.A1(new_n6883_), .A2(pi0567), .ZN(new_n6884_));
  NAND2_X1   g04448(.A1(new_n6884_), .A2(new_n6692_), .ZN(new_n6885_));
  INV_X1     g04449(.I(new_n6885_), .ZN(new_n6886_));
  NOR2_X1    g04450(.A1(new_n6886_), .A2(new_n6268_), .ZN(new_n6887_));
  NOR2_X1    g04451(.A1(new_n6887_), .A2(new_n6827_), .ZN(new_n6888_));
  NAND2_X1   g04452(.A1(new_n6888_), .A2(new_n6301_), .ZN(new_n6889_));
  INV_X1     g04453(.I(new_n6317_), .ZN(new_n6890_));
  INV_X1     g04454(.I(pi0444), .ZN(new_n6891_));
  AOI21_X1   g04455(.A1(new_n6886_), .A2(new_n6838_), .B(new_n6839_), .ZN(new_n6892_));
  NOR2_X1    g04456(.A1(new_n6892_), .A2(new_n6891_), .ZN(new_n6893_));
  AOI21_X1   g04457(.A1(new_n6886_), .A2(new_n6833_), .B(new_n6834_), .ZN(new_n6894_));
  NOR2_X1    g04458(.A1(new_n6894_), .A2(pi0444), .ZN(new_n6895_));
  NOR3_X1    g04459(.A1(new_n6893_), .A2(new_n6895_), .A3(new_n6890_), .ZN(new_n6896_));
  NOR2_X1    g04460(.A1(new_n6894_), .A2(new_n6891_), .ZN(new_n6897_));
  NOR2_X1    g04461(.A1(new_n6892_), .A2(pi0444), .ZN(new_n6898_));
  NOR3_X1    g04462(.A1(new_n6897_), .A2(new_n6898_), .A3(new_n6317_), .ZN(new_n6899_));
  OAI21_X1   g04463(.A1(new_n6896_), .A2(new_n6899_), .B(pi1196), .ZN(new_n6900_));
  NOR2_X1    g04464(.A1(new_n6886_), .A2(pi1196), .ZN(new_n6901_));
  NOR2_X1    g04465(.A1(new_n6901_), .A2(new_n6301_), .ZN(new_n6902_));
  NAND2_X1   g04466(.A1(new_n6900_), .A2(new_n6902_), .ZN(new_n6903_));
  NAND2_X1   g04467(.A1(new_n6903_), .A2(new_n6889_), .ZN(new_n6904_));
  NOR2_X1    g04468(.A1(new_n6904_), .A2(pi1199), .ZN(new_n6905_));
  NOR2_X1    g04469(.A1(new_n6905_), .A2(new_n6254_), .ZN(new_n6906_));
  OAI22_X1   g04470(.A1(new_n6904_), .A2(new_n6848_), .B1(new_n6850_), .B2(new_n6888_), .ZN(new_n6907_));
  OAI22_X1   g04471(.A1(new_n6904_), .A2(new_n6850_), .B1(new_n6848_), .B2(new_n6888_), .ZN(new_n6908_));
  AOI22_X1   g04472(.A1(new_n6854_), .A2(new_n6908_), .B1(new_n6907_), .B2(new_n6857_), .ZN(new_n6909_));
  NAND2_X1   g04473(.A1(new_n6909_), .A2(new_n6859_), .ZN(new_n6910_));
  AOI22_X1   g04474(.A1(new_n6854_), .A2(new_n6907_), .B1(new_n6908_), .B2(new_n6857_), .ZN(new_n6911_));
  NAND2_X1   g04475(.A1(new_n6911_), .A2(pi0445), .ZN(new_n6912_));
  AOI21_X1   g04476(.A1(new_n6910_), .A2(new_n6912_), .B(new_n6860_), .ZN(new_n6913_));
  AND2_X2    g04477(.A1(new_n6909_), .A2(pi0445), .Z(new_n6914_));
  AND2_X2    g04478(.A1(new_n6911_), .A2(new_n6859_), .Z(new_n6915_));
  OAI21_X1   g04479(.A1(new_n6914_), .A2(new_n6915_), .B(new_n6860_), .ZN(new_n6916_));
  NAND2_X1   g04480(.A1(new_n6916_), .A2(pi1199), .ZN(new_n6917_));
  OAI21_X1   g04481(.A1(new_n6917_), .A2(new_n6913_), .B(new_n6906_), .ZN(new_n6918_));
  AOI21_X1   g04482(.A1(new_n6886_), .A2(new_n6254_), .B(new_n6350_), .ZN(new_n6919_));
  AOI22_X1   g04483(.A1(new_n6918_), .A2(new_n6919_), .B1(new_n6795_), .B2(new_n6868_), .ZN(new_n6920_));
  OAI21_X1   g04484(.A1(new_n6920_), .A2(new_n6251_), .B(new_n6643_), .ZN(new_n6921_));
  NOR2_X1    g04485(.A1(new_n6273_), .A2(pi0333), .ZN(new_n6922_));
  NAND2_X1   g04486(.A1(new_n6828_), .A2(new_n6922_), .ZN(new_n6923_));
  NAND2_X1   g04487(.A1(new_n6379_), .A2(pi1198), .ZN(new_n6924_));
  NOR2_X1    g04488(.A1(new_n6403_), .A2(new_n6265_), .ZN(new_n6925_));
  INV_X1     g04489(.I(new_n6925_), .ZN(new_n6926_));
  NOR3_X1    g04490(.A1(new_n6926_), .A2(new_n6255_), .A3(new_n6645_), .ZN(new_n6927_));
  OR2_X2     g04491(.A1(new_n6927_), .A2(new_n6304_), .Z(new_n6928_));
  OAI21_X1   g04492(.A1(new_n6403_), .A2(new_n6263_), .B(new_n3022_), .ZN(new_n6929_));
  OAI21_X1   g04493(.A1(new_n6926_), .A2(new_n6700_), .B(pi0075), .ZN(new_n6930_));
  AOI21_X1   g04494(.A1(new_n6710_), .A2(new_n6929_), .B(new_n6930_), .ZN(new_n6931_));
  AOI21_X1   g04495(.A1(new_n6925_), .A2(new_n3273_), .B(new_n3458_), .ZN(new_n6932_));
  NOR2_X1    g04496(.A1(new_n6404_), .A2(new_n6784_), .ZN(new_n6933_));
  OAI21_X1   g04497(.A1(new_n6789_), .A2(new_n6933_), .B(new_n6932_), .ZN(new_n6934_));
  OAI21_X1   g04498(.A1(new_n6404_), .A2(new_n6814_), .B(new_n6743_), .ZN(new_n6935_));
  AOI21_X1   g04499(.A1(new_n6925_), .A2(new_n6762_), .B(new_n2628_), .ZN(new_n6936_));
  AOI21_X1   g04500(.A1(new_n6926_), .A2(new_n6756_), .B(new_n5422_), .ZN(new_n6937_));
  AOI21_X1   g04501(.A1(new_n6926_), .A2(new_n6753_), .B(new_n6764_), .ZN(new_n6938_));
  OAI21_X1   g04502(.A1(new_n6937_), .A2(new_n6938_), .B(new_n6761_), .ZN(new_n6939_));
  NAND2_X1   g04503(.A1(new_n6939_), .A2(new_n6936_), .ZN(new_n6940_));
  AOI21_X1   g04504(.A1(new_n6926_), .A2(new_n6756_), .B(new_n5446_), .ZN(new_n6941_));
  AOI21_X1   g04505(.A1(new_n6926_), .A2(new_n6753_), .B(new_n5445_), .ZN(new_n6942_));
  OAI21_X1   g04506(.A1(new_n6941_), .A2(new_n6942_), .B(new_n6744_), .ZN(new_n6943_));
  AOI21_X1   g04507(.A1(new_n6925_), .A2(new_n6759_), .B(pi0299), .ZN(new_n6944_));
  AOI21_X1   g04508(.A1(new_n6943_), .A2(new_n6944_), .B(new_n2627_), .ZN(new_n6945_));
  NAND2_X1   g04509(.A1(new_n6945_), .A2(new_n6940_), .ZN(new_n6946_));
  NAND3_X1   g04510(.A1(new_n6935_), .A2(new_n3265_), .A3(new_n6946_), .ZN(new_n6947_));
  NAND2_X1   g04511(.A1(new_n6926_), .A2(pi0038), .ZN(new_n6948_));
  AOI21_X1   g04512(.A1(new_n6947_), .A2(new_n6948_), .B(pi0100), .ZN(new_n6949_));
  INV_X1     g04513(.I(new_n6821_), .ZN(new_n6950_));
  NOR2_X1    g04514(.A1(new_n6925_), .A2(new_n6950_), .ZN(new_n6951_));
  OAI21_X1   g04515(.A1(new_n6949_), .A2(new_n6951_), .B(new_n3458_), .ZN(new_n6952_));
  AOI21_X1   g04516(.A1(new_n6952_), .A2(new_n6934_), .B(pi0075), .ZN(new_n6953_));
  OAI21_X1   g04517(.A1(new_n6953_), .A2(new_n6931_), .B(pi0567), .ZN(new_n6954_));
  AOI21_X1   g04518(.A1(new_n6954_), .A2(new_n6692_), .B(new_n6928_), .ZN(new_n6955_));
  OAI21_X1   g04519(.A1(new_n6794_), .A2(pi1196), .B(new_n6380_), .ZN(new_n6956_));
  OAI21_X1   g04520(.A1(new_n6955_), .A2(new_n6956_), .B(new_n6924_), .ZN(new_n6957_));
  NOR2_X1    g04521(.A1(new_n6416_), .A2(new_n6261_), .ZN(new_n6958_));
  AOI21_X1   g04522(.A1(new_n6927_), .A2(new_n6958_), .B(new_n6304_), .ZN(new_n6959_));
  INV_X1     g04523(.I(new_n6416_), .ZN(new_n6960_));
  NAND2_X1   g04524(.A1(new_n6268_), .A2(new_n6302_), .ZN(new_n6961_));
  AOI21_X1   g04525(.A1(new_n6960_), .A2(new_n6646_), .B(new_n6961_), .ZN(new_n6962_));
  NOR2_X1    g04526(.A1(new_n6959_), .A2(new_n6962_), .ZN(new_n6963_));
  OAI21_X1   g04527(.A1(new_n6692_), .A2(new_n6963_), .B(pi1199), .ZN(new_n6964_));
  NOR2_X1    g04528(.A1(new_n6926_), .A2(new_n6416_), .ZN(new_n6965_));
  INV_X1     g04529(.I(new_n6965_), .ZN(new_n6966_));
  OAI21_X1   g04530(.A1(new_n6966_), .A2(new_n6700_), .B(pi0075), .ZN(new_n6967_));
  NAND2_X1   g04531(.A1(new_n6966_), .A2(new_n3022_), .ZN(new_n6968_));
  AOI21_X1   g04532(.A1(new_n6710_), .A2(new_n6968_), .B(new_n6967_), .ZN(new_n6969_));
  AOI21_X1   g04533(.A1(new_n6777_), .A2(pi0228), .B(pi0232), .ZN(new_n6970_));
  NAND2_X1   g04534(.A1(new_n6966_), .A2(new_n6970_), .ZN(new_n6971_));
  INV_X1     g04535(.I(new_n6693_), .ZN(new_n6972_));
  AOI21_X1   g04536(.A1(new_n6972_), .A2(new_n5398_), .B(new_n6694_), .ZN(new_n6973_));
  NAND2_X1   g04537(.A1(new_n6973_), .A2(pi0228), .ZN(new_n6974_));
  AOI21_X1   g04538(.A1(new_n6965_), .A2(new_n6974_), .B(new_n5666_), .ZN(new_n6975_));
  INV_X1     g04539(.I(new_n6973_), .ZN(new_n6976_));
  AOI21_X1   g04540(.A1(new_n6966_), .A2(new_n6776_), .B(new_n6976_), .ZN(new_n6977_));
  INV_X1     g04541(.I(new_n6694_), .ZN(new_n6978_));
  NOR2_X1    g04542(.A1(new_n6776_), .A2(new_n6978_), .ZN(new_n6979_));
  OAI21_X1   g04543(.A1(new_n6977_), .A2(new_n6979_), .B(pi0228), .ZN(new_n6980_));
  AOI21_X1   g04544(.A1(new_n6980_), .A2(new_n6975_), .B(new_n2573_), .ZN(new_n6981_));
  OAI21_X1   g04545(.A1(new_n6966_), .A2(new_n2572_), .B(pi0100), .ZN(new_n6982_));
  AOI21_X1   g04546(.A1(new_n6981_), .A2(new_n6971_), .B(new_n6982_), .ZN(new_n6983_));
  AOI21_X1   g04547(.A1(new_n6965_), .A2(new_n6759_), .B(pi0299), .ZN(new_n6984_));
  AOI21_X1   g04548(.A1(new_n6966_), .A2(new_n6753_), .B(new_n5445_), .ZN(new_n6985_));
  AOI21_X1   g04549(.A1(new_n6966_), .A2(new_n6756_), .B(new_n5446_), .ZN(new_n6986_));
  OAI21_X1   g04550(.A1(new_n6985_), .A2(new_n6986_), .B(new_n6744_), .ZN(new_n6987_));
  AOI21_X1   g04551(.A1(new_n6987_), .A2(new_n6984_), .B(new_n2627_), .ZN(new_n6988_));
  AOI21_X1   g04552(.A1(new_n6966_), .A2(new_n6753_), .B(new_n6764_), .ZN(new_n6989_));
  AOI21_X1   g04553(.A1(new_n6966_), .A2(new_n6756_), .B(new_n5422_), .ZN(new_n6990_));
  NOR2_X1    g04554(.A1(new_n6989_), .A2(new_n6990_), .ZN(new_n6991_));
  AOI21_X1   g04555(.A1(new_n6417_), .A2(new_n6762_), .B(new_n2628_), .ZN(new_n6992_));
  OAI22_X1   g04556(.A1(new_n6991_), .A2(new_n6762_), .B1(new_n6936_), .B2(new_n6992_), .ZN(new_n6993_));
  NAND2_X1   g04557(.A1(new_n6993_), .A2(new_n6988_), .ZN(new_n6994_));
  AOI21_X1   g04558(.A1(new_n6731_), .A2(new_n6960_), .B(new_n6714_), .ZN(new_n6995_));
  OAI21_X1   g04559(.A1(new_n6958_), .A2(pi0122), .B(pi1093), .ZN(new_n6996_));
  OAI21_X1   g04560(.A1(new_n6995_), .A2(new_n6996_), .B(new_n6739_), .ZN(new_n6997_));
  INV_X1     g04561(.I(new_n6997_), .ZN(new_n6998_));
  OAI21_X1   g04562(.A1(new_n6935_), .A2(new_n6998_), .B(new_n6994_), .ZN(new_n6999_));
  OAI21_X1   g04563(.A1(new_n6966_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n7000_));
  AOI21_X1   g04564(.A1(new_n6999_), .A2(new_n3265_), .B(new_n7000_), .ZN(new_n7001_));
  OAI21_X1   g04565(.A1(new_n7001_), .A2(new_n6983_), .B(new_n3458_), .ZN(new_n7002_));
  AOI21_X1   g04566(.A1(new_n6965_), .A2(new_n3273_), .B(new_n3458_), .ZN(new_n7003_));
  INV_X1     g04567(.I(new_n6789_), .ZN(new_n7004_));
  OAI21_X1   g04568(.A1(new_n6960_), .A2(new_n6784_), .B(new_n7004_), .ZN(new_n7005_));
  OAI21_X1   g04569(.A1(new_n6933_), .A2(new_n7005_), .B(new_n7003_), .ZN(new_n7006_));
  AOI21_X1   g04570(.A1(new_n7002_), .A2(new_n7006_), .B(pi0075), .ZN(new_n7007_));
  OAI21_X1   g04571(.A1(new_n7007_), .A2(new_n6969_), .B(new_n6959_), .ZN(new_n7008_));
  AOI21_X1   g04572(.A1(new_n6417_), .A2(new_n3273_), .B(new_n3458_), .ZN(new_n7009_));
  NAND2_X1   g04573(.A1(new_n7005_), .A2(new_n7009_), .ZN(new_n7010_));
  INV_X1     g04574(.I(new_n6417_), .ZN(new_n7011_));
  AOI21_X1   g04575(.A1(new_n6756_), .A2(new_n7011_), .B(new_n5446_), .ZN(new_n7012_));
  AOI21_X1   g04576(.A1(new_n6753_), .A2(new_n7011_), .B(new_n5445_), .ZN(new_n7013_));
  OAI21_X1   g04577(.A1(new_n7012_), .A2(new_n7013_), .B(new_n6744_), .ZN(new_n7014_));
  AOI21_X1   g04578(.A1(new_n6417_), .A2(new_n6759_), .B(pi0299), .ZN(new_n7015_));
  NAND2_X1   g04579(.A1(new_n7014_), .A2(new_n7015_), .ZN(new_n7016_));
  AOI21_X1   g04580(.A1(new_n6756_), .A2(new_n7011_), .B(new_n5422_), .ZN(new_n7017_));
  AOI21_X1   g04581(.A1(new_n6753_), .A2(new_n7011_), .B(new_n6764_), .ZN(new_n7018_));
  OAI21_X1   g04582(.A1(new_n7017_), .A2(new_n7018_), .B(new_n6761_), .ZN(new_n7019_));
  AOI21_X1   g04583(.A1(new_n7019_), .A2(new_n6992_), .B(new_n2627_), .ZN(new_n7020_));
  NAND2_X1   g04584(.A1(new_n7020_), .A2(new_n7016_), .ZN(new_n7021_));
  NAND3_X1   g04585(.A1(new_n6997_), .A2(new_n2627_), .A3(new_n6737_), .ZN(new_n7022_));
  NAND3_X1   g04586(.A1(new_n7022_), .A2(new_n3265_), .A3(new_n7021_), .ZN(new_n7023_));
  NAND2_X1   g04587(.A1(new_n7011_), .A2(pi0038), .ZN(new_n7024_));
  AOI21_X1   g04588(.A1(new_n7023_), .A2(new_n7024_), .B(pi0100), .ZN(new_n7025_));
  NOR2_X1    g04589(.A1(new_n6417_), .A2(new_n6950_), .ZN(new_n7026_));
  OAI21_X1   g04590(.A1(new_n7025_), .A2(new_n7026_), .B(new_n3458_), .ZN(new_n7027_));
  AOI21_X1   g04591(.A1(new_n7027_), .A2(new_n7010_), .B(pi0075), .ZN(new_n7028_));
  OAI21_X1   g04592(.A1(new_n6416_), .A2(new_n6263_), .B(new_n3022_), .ZN(new_n7029_));
  OAI21_X1   g04593(.A1(new_n7011_), .A2(new_n6700_), .B(pi0075), .ZN(new_n7030_));
  AOI21_X1   g04594(.A1(new_n6710_), .A2(new_n7029_), .B(new_n7030_), .ZN(new_n7031_));
  OAI21_X1   g04595(.A1(new_n7028_), .A2(new_n7031_), .B(new_n6962_), .ZN(new_n7032_));
  NAND2_X1   g04596(.A1(new_n7008_), .A2(new_n7032_), .ZN(new_n7033_));
  AOI21_X1   g04597(.A1(new_n7033_), .A2(pi0567), .B(new_n6964_), .ZN(new_n7034_));
  INV_X1     g04598(.I(new_n6924_), .ZN(new_n7035_));
  AOI21_X1   g04599(.A1(new_n6827_), .A2(new_n7035_), .B(new_n6796_), .ZN(new_n7036_));
  OAI21_X1   g04600(.A1(new_n6957_), .A2(new_n7034_), .B(new_n7036_), .ZN(new_n7037_));
  OAI21_X1   g04601(.A1(new_n7037_), .A2(new_n6922_), .B(new_n6923_), .ZN(new_n7038_));
  NOR2_X1    g04602(.A1(new_n6422_), .A2(new_n6273_), .ZN(new_n7039_));
  NAND2_X1   g04603(.A1(new_n6828_), .A2(new_n7039_), .ZN(new_n7040_));
  OAI21_X1   g04604(.A1(new_n7037_), .A2(new_n7039_), .B(new_n7040_), .ZN(new_n7041_));
  AOI22_X1   g04605(.A1(new_n6366_), .A2(new_n7038_), .B1(new_n7041_), .B2(new_n6429_), .ZN(new_n7042_));
  AOI21_X1   g04606(.A1(new_n7042_), .A2(new_n6435_), .B(new_n6440_), .ZN(new_n7043_));
  AOI22_X1   g04607(.A1(new_n6366_), .A2(new_n7041_), .B1(new_n7038_), .B2(new_n6429_), .ZN(new_n7044_));
  NAND2_X1   g04608(.A1(new_n7044_), .A2(new_n6364_), .ZN(new_n7045_));
  AOI21_X1   g04609(.A1(new_n7043_), .A2(new_n7045_), .B(pi0590), .ZN(new_n7046_));
  XOR2_X1    g04610(.A1(pi0373), .A2(pi0375), .Z(new_n7047_));
  OAI21_X1   g04611(.A1(new_n6630_), .A2(new_n7047_), .B(new_n6634_), .ZN(new_n7048_));
  INV_X1     g04612(.I(pi0371), .ZN(new_n7049_));
  INV_X1     g04613(.I(new_n6618_), .ZN(new_n7050_));
  INV_X1     g04614(.I(pi0374), .ZN(new_n7051_));
  NOR2_X1    g04615(.A1(new_n7051_), .A2(new_n6274_), .ZN(new_n7052_));
  NOR2_X1    g04616(.A1(new_n6825_), .A2(new_n6268_), .ZN(new_n7053_));
  AOI21_X1   g04617(.A1(new_n6794_), .A2(new_n6268_), .B(new_n7053_), .ZN(new_n7054_));
  INV_X1     g04618(.I(new_n7054_), .ZN(new_n7055_));
  NAND2_X1   g04619(.A1(new_n7055_), .A2(new_n7052_), .ZN(new_n7056_));
  INV_X1     g04620(.I(new_n6794_), .ZN(new_n7057_));
  AOI21_X1   g04621(.A1(new_n7057_), .A2(new_n6380_), .B(new_n6593_), .ZN(new_n7058_));
  INV_X1     g04622(.I(new_n6609_), .ZN(new_n7059_));
  NOR2_X1    g04623(.A1(new_n6594_), .A2(new_n6268_), .ZN(new_n7060_));
  AOI21_X1   g04624(.A1(new_n6825_), .A2(new_n7060_), .B(new_n7059_), .ZN(new_n7061_));
  INV_X1     g04625(.I(new_n7060_), .ZN(new_n7062_));
  NAND2_X1   g04626(.A1(new_n7057_), .A2(new_n7062_), .ZN(new_n7063_));
  NOR2_X1    g04627(.A1(new_n6268_), .A2(pi0377), .ZN(new_n7064_));
  AOI21_X1   g04628(.A1(new_n6825_), .A2(new_n7064_), .B(new_n6609_), .ZN(new_n7065_));
  OAI21_X1   g04629(.A1(pi0377), .A2(new_n6268_), .B(new_n7057_), .ZN(new_n7066_));
  AOI22_X1   g04630(.A1(new_n7066_), .A2(new_n7065_), .B1(new_n7061_), .B2(new_n7063_), .ZN(new_n7067_));
  NAND2_X1   g04631(.A1(new_n7067_), .A2(pi1199), .ZN(new_n7068_));
  AOI22_X1   g04632(.A1(new_n7068_), .A2(new_n7058_), .B1(new_n6593_), .B2(new_n7055_), .ZN(new_n7069_));
  OAI21_X1   g04633(.A1(new_n7069_), .A2(new_n7052_), .B(new_n7056_), .ZN(new_n7070_));
  NOR2_X1    g04634(.A1(new_n6274_), .A2(pi0374), .ZN(new_n7071_));
  NAND2_X1   g04635(.A1(new_n7055_), .A2(new_n7071_), .ZN(new_n7072_));
  OAI21_X1   g04636(.A1(new_n7069_), .A2(new_n7071_), .B(new_n7072_), .ZN(new_n7073_));
  AOI22_X1   g04637(.A1(new_n6616_), .A2(new_n7073_), .B1(new_n7070_), .B2(new_n7050_), .ZN(new_n7074_));
  NAND2_X1   g04638(.A1(new_n7074_), .A2(new_n7049_), .ZN(new_n7075_));
  AOI22_X1   g04639(.A1(new_n6616_), .A2(new_n7070_), .B1(new_n7073_), .B2(new_n7050_), .ZN(new_n7076_));
  NAND2_X1   g04640(.A1(new_n7076_), .A2(pi0371), .ZN(new_n7077_));
  AOI21_X1   g04641(.A1(new_n7075_), .A2(new_n7077_), .B(new_n7048_), .ZN(new_n7078_));
  AND2_X2    g04642(.A1(new_n7074_), .A2(pi0371), .Z(new_n7079_));
  AND2_X2    g04643(.A1(new_n7076_), .A2(new_n7049_), .Z(new_n7080_));
  OAI21_X1   g04644(.A1(new_n7079_), .A2(new_n7080_), .B(new_n7048_), .ZN(new_n7081_));
  NAND2_X1   g04645(.A1(new_n7081_), .A2(new_n6440_), .ZN(new_n7082_));
  OAI21_X1   g04646(.A1(new_n7082_), .A2(new_n7078_), .B(new_n7046_), .ZN(new_n7083_));
  NAND2_X1   g04647(.A1(new_n6828_), .A2(new_n6534_), .ZN(new_n7084_));
  INV_X1     g04648(.I(new_n6467_), .ZN(new_n7085_));
  INV_X1     g04649(.I(pi0350), .ZN(new_n7086_));
  NAND2_X1   g04650(.A1(new_n7086_), .A2(new_n6268_), .ZN(new_n7087_));
  INV_X1     g04651(.I(new_n6513_), .ZN(new_n7088_));
  OAI21_X1   g04652(.A1(new_n6826_), .A2(new_n7087_), .B(new_n7088_), .ZN(new_n7089_));
  AOI21_X1   g04653(.A1(new_n7057_), .A2(new_n7087_), .B(new_n7089_), .ZN(new_n7090_));
  NOR2_X1    g04654(.A1(new_n7086_), .A2(pi0592), .ZN(new_n7091_));
  INV_X1     g04655(.I(new_n7091_), .ZN(new_n7092_));
  OAI21_X1   g04656(.A1(new_n6826_), .A2(new_n7092_), .B(new_n6513_), .ZN(new_n7093_));
  AOI21_X1   g04657(.A1(new_n7057_), .A2(new_n7092_), .B(new_n7093_), .ZN(new_n7094_));
  NOR3_X1    g04658(.A1(new_n7090_), .A2(new_n7094_), .A3(new_n6497_), .ZN(new_n7095_));
  OAI21_X1   g04659(.A1(new_n6828_), .A2(new_n6498_), .B(pi1198), .ZN(new_n7096_));
  NOR2_X1    g04660(.A1(new_n7095_), .A2(new_n7096_), .ZN(new_n7097_));
  XOR2_X1    g04661(.A1(new_n6484_), .A2(pi0355), .Z(new_n7098_));
  NAND2_X1   g04662(.A1(new_n6794_), .A2(pi0455), .ZN(new_n7099_));
  OAI21_X1   g04663(.A1(new_n6847_), .A2(pi0455), .B(new_n7099_), .ZN(new_n7100_));
  NAND2_X1   g04664(.A1(new_n7100_), .A2(pi0452), .ZN(new_n7101_));
  NAND2_X1   g04665(.A1(new_n6794_), .A2(new_n6488_), .ZN(new_n7102_));
  OAI21_X1   g04666(.A1(new_n6847_), .A2(new_n6488_), .B(new_n7102_), .ZN(new_n7103_));
  NAND2_X1   g04667(.A1(new_n7103_), .A2(new_n6487_), .ZN(new_n7104_));
  AOI21_X1   g04668(.A1(new_n7101_), .A2(new_n7104_), .B(new_n7098_), .ZN(new_n7105_));
  OAI21_X1   g04669(.A1(new_n7103_), .A2(new_n6487_), .B(new_n7098_), .ZN(new_n7106_));
  NOR2_X1    g04670(.A1(new_n7100_), .A2(pi0452), .ZN(new_n7107_));
  OAI21_X1   g04671(.A1(new_n7106_), .A2(new_n7107_), .B(pi1196), .ZN(new_n7108_));
  OAI21_X1   g04672(.A1(new_n7108_), .A2(new_n7105_), .B(new_n6274_), .ZN(new_n7109_));
  OAI21_X1   g04673(.A1(new_n7109_), .A2(new_n6843_), .B(new_n7085_), .ZN(new_n7110_));
  OAI22_X1   g04674(.A1(new_n7110_), .A2(new_n7097_), .B1(new_n7085_), .B2(new_n6828_), .ZN(new_n7111_));
  OAI21_X1   g04675(.A1(new_n7111_), .A2(new_n6534_), .B(new_n7084_), .ZN(new_n7112_));
  NAND2_X1   g04676(.A1(new_n6828_), .A2(new_n6444_), .ZN(new_n7113_));
  OAI21_X1   g04677(.A1(new_n7111_), .A2(new_n6444_), .B(new_n7113_), .ZN(new_n7114_));
  AOI22_X1   g04678(.A1(new_n6442_), .A2(new_n7112_), .B1(new_n7114_), .B2(new_n6533_), .ZN(new_n7115_));
  NAND2_X1   g04679(.A1(new_n7115_), .A2(new_n6550_), .ZN(new_n7116_));
  AOI22_X1   g04680(.A1(new_n6442_), .A2(new_n7114_), .B1(new_n7112_), .B2(new_n6533_), .ZN(new_n7117_));
  NAND2_X1   g04681(.A1(new_n7117_), .A2(new_n6548_), .ZN(new_n7118_));
  NAND3_X1   g04682(.A1(new_n7116_), .A2(new_n7118_), .A3(new_n6440_), .ZN(new_n7119_));
  AOI21_X1   g04683(.A1(new_n6794_), .A2(pi0591), .B(new_n6352_), .ZN(new_n7120_));
  AOI21_X1   g04684(.A1(new_n7119_), .A2(new_n7120_), .B(new_n6349_), .ZN(new_n7121_));
  AOI21_X1   g04685(.A1(new_n7121_), .A2(new_n7083_), .B(pi0588), .ZN(new_n7122_));
  NAND2_X1   g04686(.A1(new_n6888_), .A2(new_n6534_), .ZN(new_n7123_));
  NOR2_X1    g04687(.A1(new_n6886_), .A2(new_n7091_), .ZN(new_n7124_));
  OAI21_X1   g04688(.A1(new_n7124_), .A2(new_n7093_), .B(new_n6498_), .ZN(new_n7125_));
  AOI21_X1   g04689(.A1(new_n6885_), .A2(new_n7087_), .B(new_n7089_), .ZN(new_n7126_));
  NOR2_X1    g04690(.A1(new_n7125_), .A2(new_n7126_), .ZN(new_n7127_));
  OAI21_X1   g04691(.A1(new_n6888_), .A2(new_n6498_), .B(pi1198), .ZN(new_n7128_));
  NOR2_X1    g04692(.A1(new_n7127_), .A2(new_n7128_), .ZN(new_n7129_));
  INV_X1     g04693(.I(new_n6888_), .ZN(new_n7130_));
  XNOR2_X1   g04694(.A1(pi0452), .A2(pi0455), .ZN(new_n7131_));
  OAI22_X1   g04695(.A1(new_n7130_), .A2(new_n6490_), .B1(new_n6885_), .B2(new_n7131_), .ZN(new_n7132_));
  NAND2_X1   g04696(.A1(new_n7132_), .A2(pi0355), .ZN(new_n7133_));
  OAI22_X1   g04697(.A1(new_n7130_), .A2(new_n7131_), .B1(new_n6490_), .B2(new_n6885_), .ZN(new_n7134_));
  NAND2_X1   g04698(.A1(new_n7134_), .A2(new_n6485_), .ZN(new_n7135_));
  INV_X1     g04699(.I(pi0458), .ZN(new_n7136_));
  XOR2_X1    g04700(.A1(new_n6483_), .A2(new_n7136_), .Z(new_n7137_));
  NAND3_X1   g04701(.A1(new_n7133_), .A2(new_n7135_), .A3(new_n7137_), .ZN(new_n7138_));
  INV_X1     g04702(.I(new_n7137_), .ZN(new_n7139_));
  NAND2_X1   g04703(.A1(new_n7134_), .A2(pi0355), .ZN(new_n7140_));
  NAND2_X1   g04704(.A1(new_n7132_), .A2(new_n6485_), .ZN(new_n7141_));
  NAND3_X1   g04705(.A1(new_n7140_), .A2(new_n7141_), .A3(new_n7139_), .ZN(new_n7142_));
  AOI21_X1   g04706(.A1(new_n7138_), .A2(new_n7142_), .B(new_n6302_), .ZN(new_n7143_));
  OR3_X2     g04707(.A1(new_n7143_), .A2(pi1198), .A3(new_n6901_), .Z(new_n7144_));
  NAND2_X1   g04708(.A1(new_n7144_), .A2(new_n7085_), .ZN(new_n7145_));
  OAI22_X1   g04709(.A1(new_n7145_), .A2(new_n7129_), .B1(new_n7085_), .B2(new_n6888_), .ZN(new_n7146_));
  OAI21_X1   g04710(.A1(new_n7146_), .A2(new_n6534_), .B(new_n7123_), .ZN(new_n7147_));
  NAND2_X1   g04711(.A1(new_n6888_), .A2(new_n6444_), .ZN(new_n7148_));
  OAI21_X1   g04712(.A1(new_n7146_), .A2(new_n6444_), .B(new_n7148_), .ZN(new_n7149_));
  AOI22_X1   g04713(.A1(new_n6442_), .A2(new_n7147_), .B1(new_n7149_), .B2(new_n6533_), .ZN(new_n7150_));
  NAND2_X1   g04714(.A1(new_n7150_), .A2(new_n6550_), .ZN(new_n7151_));
  AOI22_X1   g04715(.A1(new_n6442_), .A2(new_n7149_), .B1(new_n7147_), .B2(new_n6533_), .ZN(new_n7152_));
  NAND2_X1   g04716(.A1(new_n7152_), .A2(new_n6548_), .ZN(new_n7153_));
  NAND3_X1   g04717(.A1(new_n7151_), .A2(new_n7153_), .A3(new_n6440_), .ZN(new_n7154_));
  AOI21_X1   g04718(.A1(new_n6886_), .A2(pi0591), .B(new_n6352_), .ZN(new_n7155_));
  NAND2_X1   g04719(.A1(new_n7154_), .A2(new_n7155_), .ZN(new_n7156_));
  INV_X1     g04720(.I(new_n6362_), .ZN(new_n7157_));
  INV_X1     g04721(.I(pi0393), .ZN(new_n7158_));
  OAI21_X1   g04722(.A1(new_n6406_), .A2(pi0075), .B(new_n6960_), .ZN(new_n7159_));
  NOR2_X1    g04723(.A1(new_n6879_), .A2(new_n7159_), .ZN(new_n7160_));
  OAI21_X1   g04724(.A1(new_n6818_), .A2(new_n7160_), .B(new_n6822_), .ZN(new_n7161_));
  NOR2_X1    g04725(.A1(pi0075), .A2(pi0592), .ZN(new_n7162_));
  NAND2_X1   g04726(.A1(new_n6873_), .A2(new_n6802_), .ZN(new_n7163_));
  NAND2_X1   g04727(.A1(new_n6960_), .A2(new_n6786_), .ZN(new_n7164_));
  AOI21_X1   g04728(.A1(new_n7164_), .A2(new_n6870_), .B(new_n7163_), .ZN(new_n7165_));
  AOI21_X1   g04729(.A1(new_n6404_), .A2(new_n6786_), .B(new_n6871_), .ZN(new_n7166_));
  NAND2_X1   g04730(.A1(new_n7166_), .A2(pi1196), .ZN(new_n7167_));
  NAND2_X1   g04731(.A1(new_n7167_), .A2(new_n7165_), .ZN(new_n7168_));
  NAND4_X1   g04732(.A1(new_n7161_), .A2(pi1199), .A3(new_n7162_), .A4(new_n7168_), .ZN(new_n7169_));
  INV_X1     g04733(.I(new_n7162_), .ZN(new_n7170_));
  NAND2_X1   g04734(.A1(new_n6883_), .A2(new_n7170_), .ZN(new_n7171_));
  AOI21_X1   g04735(.A1(new_n6404_), .A2(new_n6878_), .B(new_n6818_), .ZN(new_n7172_));
  NOR3_X1    g04736(.A1(new_n7172_), .A2(pi0087), .A3(new_n6821_), .ZN(new_n7173_));
  NOR2_X1    g04737(.A1(new_n7166_), .A2(new_n7163_), .ZN(new_n7174_));
  NOR4_X1    g04738(.A1(new_n7173_), .A2(new_n6302_), .A3(new_n7170_), .A4(new_n7174_), .ZN(new_n7175_));
  NOR2_X1    g04739(.A1(new_n6882_), .A2(pi1196), .ZN(new_n7176_));
  OAI21_X1   g04740(.A1(new_n7175_), .A2(new_n7176_), .B(new_n6380_), .ZN(new_n7177_));
  NAND3_X1   g04741(.A1(new_n7177_), .A2(new_n7169_), .A3(new_n7171_), .ZN(new_n7178_));
  NAND2_X1   g04742(.A1(new_n6692_), .A2(new_n6924_), .ZN(new_n7179_));
  AOI21_X1   g04743(.A1(new_n7178_), .A2(pi0567), .B(new_n7179_), .ZN(new_n7180_));
  AOI21_X1   g04744(.A1(new_n6888_), .A2(new_n7035_), .B(new_n7180_), .ZN(new_n7181_));
  NOR2_X1    g04745(.A1(new_n7181_), .A2(new_n7039_), .ZN(new_n7182_));
  AOI21_X1   g04746(.A1(new_n6888_), .A2(new_n7039_), .B(new_n7182_), .ZN(new_n7183_));
  INV_X1     g04747(.I(new_n7183_), .ZN(new_n7184_));
  MUX2_X1    g04748(.I0(new_n7181_), .I1(new_n7130_), .S(new_n6922_), .Z(new_n7185_));
  INV_X1     g04749(.I(new_n7185_), .ZN(new_n7186_));
  AOI22_X1   g04750(.A1(new_n7184_), .A2(new_n6429_), .B1(new_n6366_), .B2(new_n7186_), .ZN(new_n7187_));
  NOR2_X1    g04751(.A1(new_n7187_), .A2(new_n7158_), .ZN(new_n7188_));
  AOI22_X1   g04752(.A1(new_n7184_), .A2(new_n6366_), .B1(new_n6429_), .B2(new_n7186_), .ZN(new_n7189_));
  INV_X1     g04753(.I(new_n7189_), .ZN(new_n7190_));
  AOI21_X1   g04754(.A1(new_n7158_), .A2(new_n7190_), .B(new_n7188_), .ZN(new_n7191_));
  AND2_X2    g04755(.A1(new_n7191_), .A2(pi0334), .Z(new_n7192_));
  NAND2_X1   g04756(.A1(new_n7190_), .A2(pi0393), .ZN(new_n7193_));
  OAI21_X1   g04757(.A1(pi0393), .A2(new_n7187_), .B(new_n7193_), .ZN(new_n7194_));
  NOR2_X1    g04758(.A1(new_n7194_), .A2(pi0334), .ZN(new_n7195_));
  OAI21_X1   g04759(.A1(new_n7195_), .A2(new_n7192_), .B(new_n7157_), .ZN(new_n7196_));
  INV_X1     g04760(.I(pi0334), .ZN(new_n7197_));
  NAND2_X1   g04761(.A1(new_n7191_), .A2(new_n7197_), .ZN(new_n7198_));
  OAI21_X1   g04762(.A1(new_n7197_), .A2(new_n7194_), .B(new_n7198_), .ZN(new_n7199_));
  AOI21_X1   g04763(.A1(new_n7199_), .A2(new_n6362_), .B(new_n6440_), .ZN(new_n7200_));
  AOI21_X1   g04764(.A1(new_n7200_), .A2(new_n7196_), .B(pi0590), .ZN(new_n7201_));
  NOR2_X1    g04765(.A1(new_n6885_), .A2(pi0592), .ZN(new_n7202_));
  NOR2_X1    g04766(.A1(new_n7202_), .A2(new_n7053_), .ZN(new_n7203_));
  INV_X1     g04767(.I(new_n7203_), .ZN(new_n7204_));
  NOR2_X1    g04768(.A1(new_n7204_), .A2(new_n6590_), .ZN(new_n7205_));
  NOR2_X1    g04769(.A1(new_n6886_), .A2(new_n6591_), .ZN(new_n7206_));
  OAI21_X1   g04770(.A1(new_n7205_), .A2(new_n7206_), .B(new_n6570_), .ZN(new_n7207_));
  AOI21_X1   g04771(.A1(new_n6302_), .A2(new_n6590_), .B(new_n7204_), .ZN(new_n7208_));
  NOR3_X1    g04772(.A1(new_n6886_), .A2(pi1196), .A3(new_n6591_), .ZN(new_n7209_));
  OAI21_X1   g04773(.A1(new_n7208_), .A2(new_n7209_), .B(new_n6569_), .ZN(new_n7210_));
  AOI21_X1   g04774(.A1(new_n7210_), .A2(new_n7207_), .B(pi1199), .ZN(new_n7211_));
  INV_X1     g04775(.I(new_n7211_), .ZN(new_n7212_));
  OAI21_X1   g04776(.A1(new_n6886_), .A2(new_n7064_), .B(new_n7065_), .ZN(new_n7213_));
  NAND2_X1   g04777(.A1(new_n6885_), .A2(new_n7062_), .ZN(new_n7214_));
  AOI21_X1   g04778(.A1(new_n7214_), .A2(new_n7061_), .B(new_n6593_), .ZN(new_n7215_));
  AOI22_X1   g04779(.A1(new_n7215_), .A2(new_n7213_), .B1(new_n7203_), .B2(new_n6593_), .ZN(new_n7216_));
  OAI21_X1   g04780(.A1(new_n6380_), .A2(new_n7216_), .B(new_n7212_), .ZN(new_n7217_));
  XNOR2_X1   g04781(.A1(pi0369), .A2(pi0374), .ZN(new_n7218_));
  NAND2_X1   g04782(.A1(new_n6274_), .A2(pi1199), .ZN(new_n7219_));
  OAI22_X1   g04783(.A1(new_n7216_), .A2(new_n7219_), .B1(new_n6274_), .B2(new_n7204_), .ZN(new_n7220_));
  NOR2_X1    g04784(.A1(new_n7212_), .A2(pi1198), .ZN(new_n7221_));
  NOR2_X1    g04785(.A1(new_n7221_), .A2(new_n7220_), .ZN(new_n7222_));
  INV_X1     g04786(.I(new_n7222_), .ZN(new_n7223_));
  XOR2_X1    g04787(.A1(pi0369), .A2(pi0374), .Z(new_n7224_));
  OAI22_X1   g04788(.A1(new_n7223_), .A2(new_n7224_), .B1(new_n7217_), .B2(new_n7218_), .ZN(new_n7225_));
  INV_X1     g04789(.I(new_n7225_), .ZN(new_n7226_));
  XNOR2_X1   g04790(.A1(pi0370), .A2(pi0371), .ZN(new_n7227_));
  NOR2_X1    g04791(.A1(new_n7223_), .A2(new_n7218_), .ZN(new_n7228_));
  NOR2_X1    g04792(.A1(new_n7217_), .A2(new_n7224_), .ZN(new_n7229_));
  NOR2_X1    g04793(.A1(new_n7228_), .A2(new_n7229_), .ZN(new_n7230_));
  XOR2_X1    g04794(.A1(pi0370), .A2(pi0371), .Z(new_n7231_));
  OAI22_X1   g04795(.A1(new_n7226_), .A2(new_n7227_), .B1(new_n7230_), .B2(new_n7231_), .ZN(new_n7232_));
  NAND2_X1   g04796(.A1(new_n7232_), .A2(pi0373), .ZN(new_n7233_));
  INV_X1     g04797(.I(pi0373), .ZN(new_n7234_));
  INV_X1     g04798(.I(new_n7231_), .ZN(new_n7235_));
  NAND2_X1   g04799(.A1(new_n7225_), .A2(new_n7235_), .ZN(new_n7236_));
  OAI21_X1   g04800(.A1(new_n7227_), .A2(new_n7230_), .B(new_n7236_), .ZN(new_n7237_));
  NAND2_X1   g04801(.A1(new_n7237_), .A2(new_n7234_), .ZN(new_n7238_));
  NAND3_X1   g04802(.A1(new_n7238_), .A2(new_n7233_), .A3(pi0375), .ZN(new_n7239_));
  INV_X1     g04803(.I(pi0375), .ZN(new_n7240_));
  NAND2_X1   g04804(.A1(new_n7237_), .A2(pi0373), .ZN(new_n7241_));
  NAND2_X1   g04805(.A1(new_n7232_), .A2(new_n7234_), .ZN(new_n7242_));
  NAND3_X1   g04806(.A1(new_n7241_), .A2(new_n7242_), .A3(new_n7240_), .ZN(new_n7243_));
  AOI21_X1   g04807(.A1(new_n7239_), .A2(new_n7243_), .B(new_n6630_), .ZN(new_n7244_));
  AND3_X2    g04808(.A1(new_n7238_), .A2(new_n7240_), .A3(new_n7233_), .Z(new_n7245_));
  AND3_X2    g04809(.A1(new_n7241_), .A2(new_n7242_), .A3(pi0375), .Z(new_n7246_));
  OAI21_X1   g04810(.A1(new_n7245_), .A2(new_n7246_), .B(new_n6630_), .ZN(new_n7247_));
  NAND2_X1   g04811(.A1(new_n7247_), .A2(new_n6440_), .ZN(new_n7248_));
  OAI21_X1   g04812(.A1(new_n7248_), .A2(new_n7244_), .B(new_n7201_), .ZN(new_n7249_));
  NAND3_X1   g04813(.A1(new_n7249_), .A2(new_n6349_), .A3(new_n7156_), .ZN(new_n7250_));
  AOI21_X1   g04814(.A1(new_n7250_), .A2(new_n7122_), .B(new_n6921_), .ZN(new_n7251_));
  NOR3_X1    g04815(.A1(new_n7251_), .A2(pi0217), .A3(new_n6642_), .ZN(new_n7252_));
  NOR3_X1    g04816(.A1(pi1161), .A2(pi1162), .A3(pi1163), .ZN(new_n7253_));
  NAND3_X1   g04817(.A1(new_n6266_), .A2(po1038), .A3(new_n6350_), .ZN(new_n7254_));
  NAND2_X1   g04818(.A1(new_n7254_), .A2(pi0217), .ZN(new_n7255_));
  NAND2_X1   g04819(.A1(new_n6794_), .A2(new_n6350_), .ZN(new_n7256_));
  NAND2_X1   g04820(.A1(new_n6886_), .A2(new_n6349_), .ZN(new_n7257_));
  AOI21_X1   g04821(.A1(new_n7257_), .A2(new_n7256_), .B(po1038), .ZN(new_n7258_));
  OAI21_X1   g04822(.A1(new_n7258_), .A2(new_n7255_), .B(new_n7253_), .ZN(new_n7259_));
  INV_X1     g04823(.I(pi1163), .ZN(new_n7260_));
  NAND4_X1   g04824(.A1(new_n3042_), .A2(pi1161), .A3(pi1162), .A4(new_n7260_), .ZN(new_n7261_));
  OAI22_X1   g04825(.A1(new_n7252_), .A2(new_n7259_), .B1(pi0031), .B2(new_n7261_), .ZN(po0189));
  NOR2_X1    g04826(.A1(pi0055), .A2(pi0074), .ZN(new_n7263_));
  INV_X1     g04827(.I(new_n7263_), .ZN(new_n7264_));
  NOR3_X1    g04828(.A1(new_n3425_), .A2(new_n7264_), .A3(new_n2471_), .ZN(new_n7265_));
  INV_X1     g04829(.I(new_n7265_), .ZN(new_n7266_));
  NOR2_X1    g04830(.A1(new_n7266_), .A2(new_n6644_), .ZN(new_n7267_));
  INV_X1     g04831(.I(new_n7267_), .ZN(new_n7268_));
  NAND2_X1   g04832(.A1(new_n5355_), .A2(pi0032), .ZN(new_n7269_));
  NOR3_X1    g04833(.A1(new_n2783_), .A2(new_n2978_), .A3(pi0094), .ZN(new_n7270_));
  INV_X1     g04834(.I(new_n7270_), .ZN(new_n7271_));
  NOR2_X1    g04835(.A1(new_n2733_), .A2(pi0047), .ZN(new_n7272_));
  INV_X1     g04836(.I(new_n7272_), .ZN(new_n7273_));
  NOR2_X1    g04837(.A1(new_n7271_), .A2(new_n7273_), .ZN(new_n7274_));
  INV_X1     g04838(.I(pi0050), .ZN(new_n7275_));
  NOR3_X1    g04839(.A1(new_n2872_), .A2(new_n7275_), .A3(new_n6671_), .ZN(new_n7276_));
  NAND3_X1   g04840(.A1(new_n7276_), .A2(new_n2771_), .A3(new_n7274_), .ZN(new_n7277_));
  INV_X1     g04841(.I(pi0024), .ZN(new_n7278_));
  NAND2_X1   g04842(.A1(new_n7278_), .A2(new_n2985_), .ZN(new_n7279_));
  NOR3_X1    g04843(.A1(new_n5354_), .A2(pi0040), .A3(new_n7279_), .ZN(new_n7280_));
  INV_X1     g04844(.I(new_n7280_), .ZN(new_n7281_));
  NOR2_X1    g04845(.A1(new_n7277_), .A2(new_n7281_), .ZN(new_n7282_));
  NAND2_X1   g04846(.A1(new_n7282_), .A2(new_n2725_), .ZN(new_n7283_));
  AOI21_X1   g04847(.A1(new_n7283_), .A2(new_n7269_), .B(new_n5350_), .ZN(new_n7284_));
  NAND2_X1   g04848(.A1(new_n7278_), .A2(new_n3179_), .ZN(new_n7285_));
  NAND3_X1   g04849(.A1(new_n2752_), .A2(pi0032), .A3(new_n7285_), .ZN(new_n7286_));
  NOR3_X1    g04850(.A1(new_n3082_), .A2(new_n3044_), .A3(pi1093), .ZN(new_n7287_));
  NOR2_X1    g04851(.A1(new_n3086_), .A2(new_n7287_), .ZN(new_n7288_));
  INV_X1     g04852(.I(new_n7288_), .ZN(po0840));
  OAI21_X1   g04853(.A1(po0840), .A2(new_n6349_), .B(new_n3016_), .ZN(new_n7290_));
  NAND2_X1   g04854(.A1(new_n3059_), .A2(new_n2550_), .ZN(new_n7291_));
  NOR3_X1    g04855(.A1(new_n7290_), .A2(new_n6677_), .A3(new_n7291_), .ZN(new_n7292_));
  INV_X1     g04856(.I(new_n7274_), .ZN(new_n7293_));
  NOR3_X1    g04857(.A1(new_n2826_), .A2(pi0049), .A3(pi0068), .ZN(new_n7294_));
  NAND4_X1   g04858(.A1(new_n7294_), .A2(pi0076), .A3(new_n2915_), .A4(new_n2914_), .ZN(new_n7295_));
  NOR2_X1    g04859(.A1(pi0089), .A2(pi0102), .ZN(new_n7296_));
  NOR2_X1    g04860(.A1(pi0064), .A2(pi0081), .ZN(new_n7297_));
  NAND4_X1   g04861(.A1(new_n2496_), .A2(new_n6667_), .A3(new_n7296_), .A4(new_n7297_), .ZN(new_n7298_));
  NOR2_X1    g04862(.A1(pi0045), .A2(pi0048), .ZN(new_n7299_));
  INV_X1     g04863(.I(new_n7299_), .ZN(new_n7300_));
  NAND2_X1   g04864(.A1(new_n2493_), .A2(new_n2907_), .ZN(new_n7301_));
  NOR4_X1    g04865(.A1(new_n7301_), .A2(pi0061), .A3(new_n7300_), .A4(pi0104), .ZN(new_n7302_));
  INV_X1     g04866(.I(new_n7302_), .ZN(new_n7303_));
  NAND2_X1   g04867(.A1(new_n2503_), .A2(new_n2925_), .ZN(new_n7304_));
  NOR4_X1    g04868(.A1(new_n7304_), .A2(pi0085), .A3(pi0103), .A4(pi0106), .ZN(new_n7305_));
  INV_X1     g04869(.I(new_n7305_), .ZN(new_n7306_));
  NOR4_X1    g04870(.A1(new_n7303_), .A2(new_n7306_), .A3(new_n7295_), .A4(new_n7298_), .ZN(new_n7307_));
  NAND2_X1   g04871(.A1(new_n7307_), .A2(new_n2515_), .ZN(new_n7308_));
  NOR2_X1    g04872(.A1(new_n7308_), .A2(new_n7293_), .ZN(new_n7309_));
  NAND2_X1   g04873(.A1(new_n7309_), .A2(pi0024), .ZN(new_n7310_));
  NOR2_X1    g04874(.A1(new_n2872_), .A2(new_n7275_), .ZN(new_n7311_));
  NAND2_X1   g04875(.A1(new_n2728_), .A2(new_n2736_), .ZN(new_n7312_));
  INV_X1     g04876(.I(new_n7312_), .ZN(new_n7313_));
  OAI21_X1   g04877(.A1(new_n7311_), .A2(new_n7307_), .B(new_n7313_), .ZN(new_n7314_));
  OAI21_X1   g04878(.A1(new_n7314_), .A2(pi0024), .B(new_n7310_), .ZN(new_n7315_));
  AOI22_X1   g04879(.A1(new_n7292_), .A2(new_n7315_), .B1(new_n7282_), .B2(new_n7290_), .ZN(new_n7316_));
  OAI21_X1   g04880(.A1(new_n7316_), .A2(pi0032), .B(new_n7286_), .ZN(new_n7317_));
  AOI21_X1   g04881(.A1(new_n7317_), .A2(new_n5350_), .B(new_n7284_), .ZN(new_n7318_));
  NOR3_X1    g04882(.A1(new_n7318_), .A2(pi0095), .A3(new_n2575_), .ZN(new_n7319_));
  NOR4_X1    g04883(.A1(po1057), .A2(new_n2530_), .A3(new_n5309_), .A4(new_n5334_), .ZN(new_n7320_));
  NAND2_X1   g04884(.A1(new_n7320_), .A2(new_n3016_), .ZN(new_n7321_));
  INV_X1     g04885(.I(pi0129), .ZN(new_n7322_));
  NOR2_X1    g04886(.A1(new_n2530_), .A2(new_n7322_), .ZN(new_n7323_));
  NOR2_X1    g04887(.A1(new_n5323_), .A2(new_n6699_), .ZN(new_n7324_));
  NOR2_X1    g04888(.A1(new_n7324_), .A2(new_n2704_), .ZN(new_n7325_));
  NAND4_X1   g04889(.A1(new_n7325_), .A2(new_n3016_), .A3(new_n7323_), .A4(new_n5309_), .ZN(new_n7326_));
  NOR2_X1    g04890(.A1(new_n2573_), .A2(new_n2702_), .ZN(new_n7327_));
  INV_X1     g04891(.I(new_n7327_), .ZN(new_n7328_));
  AOI21_X1   g04892(.A1(new_n7326_), .A2(new_n7321_), .B(new_n7328_), .ZN(new_n7329_));
  OAI21_X1   g04893(.A1(new_n7319_), .A2(new_n7329_), .B(new_n2564_), .ZN(new_n7330_));
  NOR2_X1    g04894(.A1(new_n2526_), .A2(new_n3007_), .ZN(new_n7331_));
  INV_X1     g04895(.I(new_n7331_), .ZN(new_n7332_));
  NAND2_X1   g04896(.A1(new_n2812_), .A2(new_n7278_), .ZN(new_n7333_));
  NOR3_X1    g04897(.A1(new_n7333_), .A2(pi0051), .A3(new_n7332_), .ZN(new_n7334_));
  INV_X1     g04898(.I(new_n7334_), .ZN(new_n7335_));
  NOR2_X1    g04899(.A1(new_n2659_), .A2(new_n3465_), .ZN(new_n7336_));
  INV_X1     g04900(.I(new_n7336_), .ZN(new_n7337_));
  NOR2_X1    g04901(.A1(new_n7335_), .A2(new_n7337_), .ZN(new_n7338_));
  NOR4_X1    g04902(.A1(new_n7325_), .A2(pi0137), .A3(new_n5324_), .A4(po0840), .ZN(new_n7339_));
  NAND2_X1   g04903(.A1(new_n7338_), .A2(new_n7339_), .ZN(new_n7340_));
  AOI21_X1   g04904(.A1(new_n7330_), .A2(new_n7340_), .B(new_n7268_), .ZN(po0190));
  NOR2_X1    g04905(.A1(pi0075), .A2(pi0100), .ZN(new_n7342_));
  XNOR2_X1   g04906(.A1(pi0149), .A2(pi0157), .ZN(new_n7343_));
  NOR2_X1    g04907(.A1(new_n7343_), .A2(new_n5437_), .ZN(new_n7344_));
  INV_X1     g04908(.I(new_n7344_), .ZN(new_n7345_));
  NOR2_X1    g04909(.A1(new_n7345_), .A2(new_n5666_), .ZN(new_n7346_));
  NOR2_X1    g04910(.A1(new_n7346_), .A2(new_n7342_), .ZN(new_n7347_));
  INV_X1     g04911(.I(new_n7342_), .ZN(new_n7348_));
  NOR2_X1    g04912(.A1(new_n6698_), .A2(new_n7348_), .ZN(new_n7349_));
  INV_X1     g04913(.I(new_n7349_), .ZN(new_n7350_));
  NOR2_X1    g04914(.A1(new_n7350_), .A2(new_n4414_), .ZN(new_n7351_));
  OAI21_X1   g04915(.A1(new_n7347_), .A2(new_n7351_), .B(pi0074), .ZN(new_n7352_));
  INV_X1     g04916(.I(new_n7352_), .ZN(new_n7353_));
  AOI21_X1   g04917(.A1(pi0164), .A2(new_n7349_), .B(new_n7347_), .ZN(new_n7354_));
  NOR2_X1    g04918(.A1(new_n7354_), .A2(pi0074), .ZN(new_n7355_));
  NOR3_X1    g04919(.A1(new_n7355_), .A2(new_n3291_), .A3(new_n7353_), .ZN(new_n7356_));
  NOR2_X1    g04920(.A1(new_n7354_), .A2(new_n5499_), .ZN(new_n7357_));
  INV_X1     g04921(.I(new_n7357_), .ZN(new_n7358_));
  INV_X1     g04922(.I(pi0164), .ZN(new_n7359_));
  NOR2_X1    g04923(.A1(new_n6698_), .A2(new_n7359_), .ZN(new_n7360_));
  INV_X1     g04924(.I(new_n7360_), .ZN(new_n7361_));
  NOR2_X1    g04925(.A1(new_n7361_), .A2(new_n3265_), .ZN(new_n7362_));
  AOI21_X1   g04926(.A1(new_n7342_), .A2(new_n7362_), .B(new_n7347_), .ZN(new_n7363_));
  NAND2_X1   g04927(.A1(new_n7358_), .A2(new_n7363_), .ZN(new_n7364_));
  AOI21_X1   g04928(.A1(new_n7364_), .A2(new_n2625_), .B(new_n7353_), .ZN(new_n7365_));
  OAI21_X1   g04929(.A1(new_n7365_), .A2(new_n2470_), .B(new_n3291_), .ZN(new_n7366_));
  XOR2_X1    g04930(.A1(pi0178), .A2(pi0183), .Z(new_n7367_));
  NAND3_X1   g04931(.A1(new_n7367_), .A2(new_n2628_), .A3(new_n5398_), .ZN(new_n7368_));
  OAI21_X1   g04932(.A1(new_n7345_), .A2(new_n2628_), .B(new_n7368_), .ZN(new_n7369_));
  NAND2_X1   g04933(.A1(new_n7369_), .A2(pi0232), .ZN(new_n7370_));
  NAND2_X1   g04934(.A1(new_n7370_), .A2(pi0100), .ZN(new_n7371_));
  INV_X1     g04935(.I(new_n7371_), .ZN(new_n7372_));
  NAND2_X1   g04936(.A1(new_n7370_), .A2(pi0075), .ZN(new_n7373_));
  INV_X1     g04937(.I(new_n7373_), .ZN(new_n7374_));
  NOR2_X1    g04938(.A1(new_n7372_), .A2(new_n7374_), .ZN(new_n7375_));
  NOR2_X1    g04939(.A1(pi0191), .A2(pi0299), .ZN(new_n7376_));
  AOI21_X1   g04940(.A1(new_n4414_), .A2(pi0299), .B(new_n7376_), .ZN(new_n7377_));
  INV_X1     g04941(.I(new_n7377_), .ZN(new_n7378_));
  OAI21_X1   g04942(.A1(new_n7350_), .A2(new_n7378_), .B(new_n7375_), .ZN(new_n7379_));
  AOI21_X1   g04943(.A1(new_n7379_), .A2(pi0074), .B(pi0055), .ZN(new_n7380_));
  INV_X1     g04944(.I(pi0186), .ZN(new_n7381_));
  NOR2_X1    g04945(.A1(new_n7381_), .A2(pi0299), .ZN(new_n7382_));
  AOI21_X1   g04946(.A1(pi0164), .A2(pi0299), .B(new_n7382_), .ZN(new_n7383_));
  NOR2_X1    g04947(.A1(new_n6698_), .A2(new_n7383_), .ZN(new_n7384_));
  NAND2_X1   g04948(.A1(new_n7384_), .A2(new_n7342_), .ZN(new_n7385_));
  AOI21_X1   g04949(.A1(new_n7375_), .A2(new_n7385_), .B(new_n5499_), .ZN(new_n7386_));
  NOR2_X1    g04950(.A1(new_n3444_), .A2(pi0075), .ZN(new_n7387_));
  NOR2_X1    g04951(.A1(new_n3265_), .A2(pi0100), .ZN(new_n7388_));
  AOI21_X1   g04952(.A1(new_n7388_), .A2(new_n7384_), .B(new_n7372_), .ZN(new_n7389_));
  INV_X1     g04953(.I(new_n7389_), .ZN(new_n7390_));
  AOI21_X1   g04954(.A1(new_n3321_), .A2(pi0299), .B(new_n5666_), .ZN(new_n7391_));
  INV_X1     g04955(.I(new_n7391_), .ZN(new_n7392_));
  NOR2_X1    g04956(.A1(pi0176), .A2(pi0299), .ZN(new_n7393_));
  NOR3_X1    g04957(.A1(new_n7392_), .A2(new_n5437_), .A3(new_n7393_), .ZN(new_n7394_));
  AND3_X2    g04958(.A1(new_n5345_), .A2(new_n2626_), .A3(new_n7394_), .Z(new_n7395_));
  OAI21_X1   g04959(.A1(new_n7395_), .A2(new_n7390_), .B(new_n7387_), .ZN(new_n7396_));
  NOR2_X1    g04960(.A1(new_n5336_), .A2(new_n6698_), .ZN(new_n7397_));
  INV_X1     g04961(.I(new_n7397_), .ZN(new_n7398_));
  NOR2_X1    g04962(.A1(new_n7398_), .A2(new_n7381_), .ZN(new_n7399_));
  NOR2_X1    g04963(.A1(new_n5345_), .A2(new_n6698_), .ZN(new_n7400_));
  NAND2_X1   g04964(.A1(new_n7400_), .A2(pi0299), .ZN(new_n7401_));
  NOR2_X1    g04965(.A1(new_n7401_), .A2(pi0186), .ZN(new_n7402_));
  OAI21_X1   g04966(.A1(new_n7402_), .A2(new_n7399_), .B(pi0164), .ZN(new_n7403_));
  INV_X1     g04967(.I(new_n7403_), .ZN(new_n7404_));
  NAND2_X1   g04968(.A1(new_n7400_), .A2(new_n2628_), .ZN(new_n7405_));
  NOR3_X1    g04969(.A1(new_n7405_), .A2(pi0164), .A3(new_n7381_), .ZN(new_n7406_));
  NOR3_X1    g04970(.A1(new_n7404_), .A2(new_n7406_), .A3(new_n3265_), .ZN(new_n7407_));
  INV_X1     g04971(.I(new_n7407_), .ZN(new_n7408_));
  INV_X1     g04972(.I(new_n2496_), .ZN(new_n7409_));
  NOR3_X1    g04973(.A1(new_n2796_), .A2(new_n2522_), .A3(new_n2785_), .ZN(new_n7410_));
  INV_X1     g04974(.I(new_n7410_), .ZN(new_n7411_));
  NAND2_X1   g04975(.A1(new_n2793_), .A2(new_n2788_), .ZN(new_n7412_));
  NAND2_X1   g04976(.A1(new_n2505_), .A2(new_n2501_), .ZN(new_n7413_));
  INV_X1     g04977(.I(new_n7413_), .ZN(new_n7414_));
  NAND3_X1   g04978(.A1(new_n7414_), .A2(new_n2493_), .A3(new_n7297_), .ZN(new_n7415_));
  INV_X1     g04979(.I(pi0036), .ZN(new_n7416_));
  NOR2_X1    g04980(.A1(new_n2824_), .A2(pi0068), .ZN(new_n7417_));
  NOR2_X1    g04981(.A1(new_n2475_), .A2(pi0111), .ZN(new_n7418_));
  NAND3_X1   g04982(.A1(new_n7417_), .A2(new_n7418_), .A3(new_n7416_), .ZN(new_n7419_));
  NOR3_X1    g04983(.A1(new_n7415_), .A2(new_n2540_), .A3(new_n7419_), .ZN(new_n7420_));
  NAND4_X1   g04984(.A1(new_n7420_), .A2(new_n2911_), .A3(new_n2915_), .A4(new_n2928_), .ZN(new_n7421_));
  OAI21_X1   g04985(.A1(new_n7421_), .A2(new_n7412_), .B(new_n2496_), .ZN(new_n7422_));
  AOI21_X1   g04986(.A1(new_n7311_), .A2(new_n2788_), .B(new_n2880_), .ZN(new_n7423_));
  NOR2_X1    g04987(.A1(new_n7415_), .A2(new_n2545_), .ZN(new_n7424_));
  INV_X1     g04988(.I(new_n7424_), .ZN(new_n7425_));
  NOR2_X1    g04989(.A1(new_n7425_), .A2(pi0060), .ZN(new_n7426_));
  INV_X1     g04990(.I(new_n7426_), .ZN(new_n7427_));
  AOI21_X1   g04991(.A1(pi0053), .A2(new_n7427_), .B(new_n7423_), .ZN(new_n7428_));
  OAI21_X1   g04992(.A1(new_n7428_), .A2(new_n7422_), .B(new_n2791_), .ZN(new_n7429_));
  OR3_X2     g04993(.A1(new_n7429_), .A2(new_n7409_), .A3(new_n7411_), .Z(new_n7430_));
  NAND2_X1   g04994(.A1(new_n7430_), .A2(new_n2835_), .ZN(new_n7431_));
  INV_X1     g04995(.I(new_n7431_), .ZN(new_n7432_));
  NOR2_X1    g04996(.A1(new_n3172_), .A2(new_n2526_), .ZN(new_n7433_));
  INV_X1     g04997(.I(new_n7433_), .ZN(new_n7434_));
  NOR2_X1    g04998(.A1(new_n7432_), .A2(new_n7434_), .ZN(new_n7435_));
  NOR2_X1    g04999(.A1(new_n7435_), .A2(new_n5617_), .ZN(new_n7436_));
  NOR2_X1    g05000(.A1(new_n6662_), .A2(new_n2985_), .ZN(new_n7437_));
  NOR3_X1    g05001(.A1(new_n7437_), .A2(new_n2537_), .A3(new_n5361_), .ZN(new_n7438_));
  INV_X1     g05002(.I(new_n7438_), .ZN(new_n7439_));
  NAND2_X1   g05003(.A1(new_n7432_), .A2(new_n7439_), .ZN(new_n7440_));
  NAND2_X1   g05004(.A1(new_n7440_), .A2(new_n7433_), .ZN(new_n7441_));
  INV_X1     g05005(.I(new_n7441_), .ZN(new_n7442_));
  NAND2_X1   g05006(.A1(new_n7442_), .A2(pi0172), .ZN(new_n7443_));
  NAND3_X1   g05007(.A1(new_n7443_), .A2(new_n3369_), .A3(new_n7436_), .ZN(new_n7444_));
  OAI21_X1   g05008(.A1(new_n7423_), .A2(new_n7411_), .B(new_n2835_), .ZN(new_n7445_));
  INV_X1     g05009(.I(new_n7445_), .ZN(new_n7446_));
  NOR2_X1    g05010(.A1(new_n7446_), .A2(new_n7434_), .ZN(new_n7447_));
  NOR2_X1    g05011(.A1(new_n7447_), .A2(new_n5617_), .ZN(new_n7448_));
  AOI21_X1   g05012(.A1(new_n7446_), .A2(new_n7439_), .B(new_n7434_), .ZN(new_n7449_));
  NAND2_X1   g05013(.A1(new_n7449_), .A2(pi0172), .ZN(new_n7450_));
  NAND3_X1   g05014(.A1(new_n7450_), .A2(new_n7448_), .A3(pi0152), .ZN(new_n7451_));
  NAND4_X1   g05015(.A1(new_n7444_), .A2(pi0149), .A3(new_n5398_), .A4(new_n7451_), .ZN(new_n7452_));
  NOR2_X1    g05016(.A1(new_n3184_), .A2(new_n5437_), .ZN(new_n7453_));
  AOI21_X1   g05017(.A1(new_n7453_), .A2(pi0158), .B(new_n2628_), .ZN(new_n7454_));
  INV_X1     g05018(.I(pi0149), .ZN(new_n7455_));
  INV_X1     g05019(.I(new_n2525_), .ZN(new_n7456_));
  NOR3_X1    g05020(.A1(new_n7456_), .A2(new_n5437_), .A3(pi0040), .ZN(new_n7457_));
  NOR2_X1    g05021(.A1(new_n7437_), .A2(new_n2747_), .ZN(new_n7458_));
  NAND3_X1   g05022(.A1(new_n7458_), .A2(new_n2821_), .A3(new_n2771_), .ZN(new_n7459_));
  NOR2_X1    g05023(.A1(new_n7459_), .A2(new_n5361_), .ZN(new_n7460_));
  NAND2_X1   g05024(.A1(new_n7460_), .A2(new_n7457_), .ZN(new_n7461_));
  INV_X1     g05025(.I(new_n7461_), .ZN(new_n7462_));
  NOR2_X1    g05026(.A1(new_n7421_), .A2(new_n7312_), .ZN(new_n7463_));
  NAND2_X1   g05027(.A1(new_n7463_), .A2(new_n2496_), .ZN(new_n7464_));
  AOI21_X1   g05028(.A1(new_n5361_), .A2(new_n7464_), .B(new_n7459_), .ZN(new_n7465_));
  NAND2_X1   g05029(.A1(new_n7465_), .A2(new_n7457_), .ZN(new_n7466_));
  INV_X1     g05030(.I(new_n7466_), .ZN(new_n7467_));
  AOI21_X1   g05031(.A1(new_n7467_), .A2(new_n3369_), .B(new_n7462_), .ZN(new_n7468_));
  NAND2_X1   g05032(.A1(new_n2748_), .A2(new_n2821_), .ZN(new_n7469_));
  NOR2_X1    g05033(.A1(new_n7464_), .A2(new_n7469_), .ZN(new_n7470_));
  INV_X1     g05034(.I(new_n7470_), .ZN(new_n7471_));
  NOR2_X1    g05035(.A1(new_n7471_), .A2(new_n7456_), .ZN(new_n7472_));
  INV_X1     g05036(.I(new_n7472_), .ZN(new_n7473_));
  NOR3_X1    g05037(.A1(new_n7473_), .A2(pi0040), .A3(new_n5437_), .ZN(new_n7474_));
  NAND2_X1   g05038(.A1(new_n7474_), .A2(new_n3778_), .ZN(new_n7475_));
  OAI22_X1   g05039(.A1(new_n7468_), .A2(new_n3778_), .B1(pi0152), .B2(new_n7475_), .ZN(new_n7476_));
  NAND2_X1   g05040(.A1(new_n7476_), .A2(new_n7455_), .ZN(new_n7477_));
  AND3_X2    g05041(.A1(new_n7452_), .A2(new_n7454_), .A3(new_n7477_), .Z(new_n7478_));
  INV_X1     g05042(.I(pi0183), .ZN(new_n7479_));
  NOR2_X1    g05043(.A1(new_n5437_), .A2(new_n7479_), .ZN(new_n7480_));
  NOR2_X1    g05044(.A1(new_n7435_), .A2(new_n5647_), .ZN(new_n7481_));
  OAI21_X1   g05045(.A1(new_n7434_), .A2(new_n7446_), .B(new_n5648_), .ZN(new_n7482_));
  NAND2_X1   g05046(.A1(new_n7482_), .A2(pi0174), .ZN(new_n7483_));
  OAI21_X1   g05047(.A1(new_n7481_), .A2(pi0174), .B(new_n7483_), .ZN(new_n7484_));
  NAND2_X1   g05048(.A1(new_n7484_), .A2(new_n7480_), .ZN(new_n7485_));
  NOR2_X1    g05049(.A1(pi0174), .A2(pi0183), .ZN(new_n7486_));
  AOI21_X1   g05050(.A1(new_n7474_), .A2(new_n7486_), .B(pi0193), .ZN(new_n7487_));
  INV_X1     g05051(.I(pi0174), .ZN(new_n7488_));
  NOR2_X1    g05052(.A1(new_n7449_), .A2(new_n5647_), .ZN(new_n7489_));
  NOR2_X1    g05053(.A1(new_n7489_), .A2(new_n5437_), .ZN(new_n7490_));
  INV_X1     g05054(.I(new_n7490_), .ZN(new_n7491_));
  NOR2_X1    g05055(.A1(new_n7462_), .A2(pi0183), .ZN(new_n7492_));
  AOI21_X1   g05056(.A1(new_n7491_), .A2(pi0183), .B(new_n7492_), .ZN(new_n7493_));
  OAI21_X1   g05057(.A1(new_n7466_), .A2(pi0183), .B(new_n7488_), .ZN(new_n7494_));
  INV_X1     g05058(.I(new_n7480_), .ZN(new_n7495_));
  NOR2_X1    g05059(.A1(new_n7435_), .A2(new_n5615_), .ZN(new_n7496_));
  NOR2_X1    g05060(.A1(new_n7496_), .A2(pi0198), .ZN(new_n7497_));
  NOR2_X1    g05061(.A1(new_n7497_), .A2(new_n7442_), .ZN(new_n7498_));
  NOR2_X1    g05062(.A1(new_n7498_), .A2(new_n7495_), .ZN(new_n7499_));
  OAI22_X1   g05063(.A1(new_n7499_), .A2(new_n7494_), .B1(new_n7488_), .B2(new_n7493_), .ZN(new_n7500_));
  AOI22_X1   g05064(.A1(new_n7500_), .A2(pi0193), .B1(new_n7485_), .B2(new_n7487_), .ZN(new_n7501_));
  NAND2_X1   g05065(.A1(new_n7453_), .A2(pi0180), .ZN(new_n7502_));
  NAND2_X1   g05066(.A1(new_n7502_), .A2(new_n2628_), .ZN(new_n7503_));
  NOR2_X1    g05067(.A1(new_n5666_), .A2(pi0039), .ZN(new_n7504_));
  OAI21_X1   g05068(.A1(new_n7501_), .A2(new_n7503_), .B(new_n7504_), .ZN(new_n7505_));
  NOR2_X1    g05069(.A1(new_n2627_), .A2(new_n5666_), .ZN(new_n7506_));
  INV_X1     g05070(.I(new_n7506_), .ZN(new_n7507_));
  NOR2_X1    g05071(.A1(new_n5550_), .A2(new_n2614_), .ZN(new_n7508_));
  NOR3_X1    g05072(.A1(new_n5551_), .A2(new_n5437_), .A3(new_n5422_), .ZN(new_n7509_));
  NAND2_X1   g05073(.A1(new_n7509_), .A2(pi0154), .ZN(new_n7510_));
  NOR3_X1    g05074(.A1(new_n5541_), .A2(new_n5437_), .A3(new_n5422_), .ZN(new_n7511_));
  NAND2_X1   g05075(.A1(new_n7511_), .A2(new_n3321_), .ZN(new_n7512_));
  AOI21_X1   g05076(.A1(new_n7510_), .A2(new_n7512_), .B(pi0152), .ZN(new_n7513_));
  NOR3_X1    g05077(.A1(new_n6751_), .A2(new_n5437_), .A3(new_n5422_), .ZN(new_n7514_));
  AND3_X2    g05078(.A1(new_n7514_), .A2(pi0152), .A3(pi0154), .Z(new_n7515_));
  OAI21_X1   g05079(.A1(new_n7515_), .A2(new_n7513_), .B(new_n7508_), .ZN(new_n7516_));
  NAND2_X1   g05080(.A1(new_n7516_), .A2(pi0299), .ZN(new_n7517_));
  INV_X1     g05081(.I(pi0176), .ZN(new_n7518_));
  NOR2_X1    g05082(.A1(new_n5525_), .A2(new_n2631_), .ZN(new_n7519_));
  INV_X1     g05083(.I(new_n5450_), .ZN(new_n7520_));
  NOR2_X1    g05084(.A1(new_n5541_), .A2(new_n7520_), .ZN(new_n7521_));
  NAND2_X1   g05085(.A1(new_n7521_), .A2(new_n7519_), .ZN(new_n7522_));
  NOR2_X1    g05086(.A1(new_n7522_), .A2(pi0174), .ZN(new_n7523_));
  AOI21_X1   g05087(.A1(new_n7523_), .A2(new_n7518_), .B(pi0299), .ZN(new_n7524_));
  INV_X1     g05088(.I(new_n7519_), .ZN(new_n7525_));
  NOR3_X1    g05089(.A1(new_n6751_), .A2(new_n7520_), .A3(new_n7525_), .ZN(new_n7526_));
  NOR3_X1    g05090(.A1(new_n5551_), .A2(new_n7520_), .A3(new_n7525_), .ZN(new_n7527_));
  OR2_X2     g05091(.A1(new_n7527_), .A2(pi0174), .Z(new_n7528_));
  OAI21_X1   g05092(.A1(new_n7526_), .A2(new_n7488_), .B(new_n7528_), .ZN(new_n7529_));
  OAI21_X1   g05093(.A1(new_n7529_), .A2(new_n7518_), .B(new_n7524_), .ZN(new_n7530_));
  NAND2_X1   g05094(.A1(new_n7517_), .A2(new_n7530_), .ZN(new_n7531_));
  OAI22_X1   g05095(.A1(new_n7505_), .A2(new_n7478_), .B1(new_n7507_), .B2(new_n7531_), .ZN(new_n7532_));
  OAI21_X1   g05096(.A1(new_n7532_), .A2(pi0038), .B(new_n7408_), .ZN(new_n7533_));
  AOI21_X1   g05097(.A1(new_n7384_), .A2(pi0038), .B(new_n3458_), .ZN(new_n7534_));
  OR2_X2     g05098(.A1(new_n7534_), .A2(pi0100), .Z(new_n7535_));
  AOI21_X1   g05099(.A1(new_n7533_), .A2(new_n3458_), .B(new_n7535_), .ZN(new_n7536_));
  OAI21_X1   g05100(.A1(new_n7536_), .A2(new_n7372_), .B(new_n2605_), .ZN(new_n7537_));
  NAND3_X1   g05101(.A1(new_n7537_), .A2(new_n7373_), .A3(new_n7396_), .ZN(new_n7538_));
  AOI21_X1   g05102(.A1(new_n7538_), .A2(new_n5499_), .B(new_n7386_), .ZN(new_n7539_));
  OAI21_X1   g05103(.A1(new_n7539_), .A2(pi0074), .B(new_n7380_), .ZN(new_n7540_));
  INV_X1     g05104(.I(new_n7346_), .ZN(new_n7541_));
  NOR2_X1    g05105(.A1(new_n7541_), .A2(new_n3465_), .ZN(new_n7542_));
  INV_X1     g05106(.I(new_n7362_), .ZN(new_n7543_));
  OAI22_X1   g05107(.A1(new_n7543_), .A2(new_n6801_), .B1(new_n2702_), .B2(new_n7346_), .ZN(new_n7544_));
  AOI21_X1   g05108(.A1(new_n7361_), .A2(pi0038), .B(new_n2604_), .ZN(new_n7545_));
  NOR2_X1    g05109(.A1(new_n6698_), .A2(new_n7455_), .ZN(new_n7546_));
  INV_X1     g05110(.I(new_n7546_), .ZN(new_n7547_));
  OAI21_X1   g05111(.A1(new_n5346_), .A2(new_n7547_), .B(new_n3265_), .ZN(new_n7548_));
  AOI21_X1   g05112(.A1(new_n7548_), .A2(new_n7545_), .B(new_n7544_), .ZN(new_n7549_));
  AOI21_X1   g05113(.A1(new_n7549_), .A2(new_n3465_), .B(new_n7542_), .ZN(new_n7550_));
  NAND2_X1   g05114(.A1(new_n7363_), .A2(pi0092), .ZN(new_n7551_));
  OAI21_X1   g05115(.A1(new_n7550_), .A2(pi0092), .B(new_n7551_), .ZN(new_n7552_));
  OAI21_X1   g05116(.A1(new_n7552_), .A2(pi0054), .B(new_n7358_), .ZN(new_n7553_));
  AOI21_X1   g05117(.A1(new_n7553_), .A2(new_n2625_), .B(new_n2602_), .ZN(new_n7554_));
  AOI21_X1   g05118(.A1(new_n7554_), .A2(new_n7352_), .B(new_n2471_), .ZN(new_n7555_));
  AOI21_X1   g05119(.A1(new_n7540_), .A2(new_n7555_), .B(new_n7366_), .ZN(new_n7556_));
  OR2_X2     g05120(.A1(new_n7556_), .A2(new_n7356_), .Z(new_n7557_));
  INV_X1     g05121(.I(pi0033), .ZN(new_n7558_));
  INV_X1     g05122(.I(pi0034), .ZN(new_n7559_));
  INV_X1     g05123(.I(pi0079), .ZN(new_n7560_));
  NOR4_X1    g05124(.A1(pi0138), .A2(pi0139), .A3(pi0195), .A4(pi0196), .ZN(new_n7561_));
  INV_X1     g05125(.I(new_n7561_), .ZN(new_n7562_));
  NOR2_X1    g05126(.A1(new_n7562_), .A2(pi0118), .ZN(new_n7563_));
  NAND3_X1   g05127(.A1(new_n7563_), .A2(new_n7559_), .A3(new_n7560_), .ZN(new_n7564_));
  NAND2_X1   g05128(.A1(new_n7564_), .A2(new_n7558_), .ZN(new_n7565_));
  INV_X1     g05129(.I(new_n7542_), .ZN(new_n7566_));
  INV_X1     g05130(.I(new_n7545_), .ZN(new_n7567_));
  NOR2_X1    g05131(.A1(new_n7409_), .A2(pi0040), .ZN(new_n7568_));
  INV_X1     g05132(.I(new_n2551_), .ZN(new_n7569_));
  NOR2_X1    g05133(.A1(new_n2785_), .A2(new_n2792_), .ZN(new_n7570_));
  INV_X1     g05134(.I(new_n7570_), .ZN(new_n7571_));
  NOR2_X1    g05135(.A1(new_n7571_), .A2(pi0053), .ZN(new_n7572_));
  INV_X1     g05136(.I(new_n7572_), .ZN(new_n7573_));
  NOR2_X1    g05137(.A1(new_n7427_), .A2(new_n7573_), .ZN(new_n7574_));
  INV_X1     g05138(.I(new_n7574_), .ZN(new_n7575_));
  NOR2_X1    g05139(.A1(new_n7575_), .A2(pi0058), .ZN(new_n7576_));
  INV_X1     g05140(.I(new_n7576_), .ZN(new_n7577_));
  NOR2_X1    g05141(.A1(new_n7577_), .A2(new_n6677_), .ZN(new_n7578_));
  NAND3_X1   g05142(.A1(new_n7578_), .A2(new_n2725_), .A3(new_n7569_), .ZN(new_n7579_));
  NOR2_X1    g05143(.A1(new_n7579_), .A2(pi0095), .ZN(new_n7580_));
  NAND3_X1   g05144(.A1(new_n7580_), .A2(new_n2627_), .A3(new_n7547_), .ZN(new_n7581_));
  AOI21_X1   g05145(.A1(new_n7581_), .A2(new_n7568_), .B(pi0038), .ZN(new_n7582_));
  INV_X1     g05146(.I(new_n7568_), .ZN(new_n7583_));
  NOR2_X1    g05147(.A1(new_n7583_), .A2(pi0038), .ZN(new_n7584_));
  INV_X1     g05148(.I(new_n7584_), .ZN(new_n7585_));
  AOI21_X1   g05149(.A1(new_n7543_), .A2(new_n7585_), .B(pi0100), .ZN(new_n7586_));
  AOI22_X1   g05150(.A1(new_n7586_), .A2(pi0087), .B1(pi0100), .B2(new_n7541_), .ZN(new_n7587_));
  OAI21_X1   g05151(.A1(new_n7582_), .A2(new_n7567_), .B(new_n7587_), .ZN(new_n7588_));
  OAI21_X1   g05152(.A1(new_n7588_), .A2(pi0075), .B(new_n7566_), .ZN(new_n7589_));
  NAND2_X1   g05153(.A1(new_n7586_), .A2(new_n3465_), .ZN(new_n7590_));
  NAND2_X1   g05154(.A1(new_n7590_), .A2(pi0092), .ZN(new_n7591_));
  OAI21_X1   g05155(.A1(new_n7591_), .A2(new_n7347_), .B(new_n5499_), .ZN(new_n7592_));
  AOI21_X1   g05156(.A1(new_n7589_), .A2(new_n3444_), .B(new_n7592_), .ZN(new_n7593_));
  OAI21_X1   g05157(.A1(new_n7593_), .A2(new_n7357_), .B(new_n2625_), .ZN(new_n7594_));
  NAND3_X1   g05158(.A1(new_n7594_), .A2(pi0055), .A3(new_n7352_), .ZN(new_n7595_));
  NOR2_X1    g05159(.A1(new_n7583_), .A2(new_n3271_), .ZN(new_n7596_));
  INV_X1     g05160(.I(new_n7580_), .ZN(new_n7597_));
  NOR2_X1    g05161(.A1(pi0039), .A2(pi0087), .ZN(new_n7598_));
  INV_X1     g05162(.I(new_n7598_), .ZN(new_n7599_));
  NOR2_X1    g05163(.A1(new_n7597_), .A2(new_n7599_), .ZN(new_n7600_));
  INV_X1     g05164(.I(new_n7600_), .ZN(new_n7601_));
  OAI21_X1   g05165(.A1(new_n7601_), .A2(new_n7394_), .B(new_n7596_), .ZN(new_n7602_));
  NAND2_X1   g05166(.A1(new_n7602_), .A2(new_n7389_), .ZN(new_n7603_));
  AOI21_X1   g05167(.A1(new_n7603_), .A2(new_n7387_), .B(new_n7374_), .ZN(new_n7604_));
  INV_X1     g05168(.I(new_n5397_), .ZN(new_n7605_));
  NOR4_X1    g05169(.A1(new_n5396_), .A2(new_n3040_), .A3(new_n5529_), .A4(new_n5539_), .ZN(new_n7606_));
  INV_X1     g05170(.I(new_n7606_), .ZN(new_n7607_));
  AOI21_X1   g05171(.A1(new_n7605_), .A2(new_n7607_), .B(new_n7597_), .ZN(new_n7608_));
  AOI21_X1   g05172(.A1(new_n7608_), .A2(new_n5449_), .B(new_n7583_), .ZN(new_n7609_));
  NOR2_X1    g05173(.A1(new_n7583_), .A2(new_n7519_), .ZN(new_n7610_));
  NOR2_X1    g05174(.A1(new_n7609_), .A2(new_n7610_), .ZN(new_n7611_));
  INV_X1     g05175(.I(new_n7611_), .ZN(new_n7612_));
  INV_X1     g05176(.I(new_n7610_), .ZN(new_n7613_));
  NOR2_X1    g05177(.A1(new_n7597_), .A2(new_n7607_), .ZN(new_n7614_));
  AOI21_X1   g05178(.A1(new_n7614_), .A2(new_n5398_), .B(new_n7583_), .ZN(new_n7615_));
  NOR2_X1    g05179(.A1(new_n7615_), .A2(new_n5446_), .ZN(new_n7616_));
  NAND3_X1   g05180(.A1(new_n7616_), .A2(pi0174), .A3(new_n7613_), .ZN(new_n7617_));
  NAND2_X1   g05181(.A1(new_n7612_), .A2(new_n7617_), .ZN(new_n7618_));
  NOR2_X1    g05182(.A1(new_n7583_), .A2(new_n7508_), .ZN(new_n7619_));
  NOR2_X1    g05183(.A1(new_n7619_), .A2(new_n2628_), .ZN(new_n7620_));
  INV_X1     g05184(.I(new_n7609_), .ZN(new_n7621_));
  OAI21_X1   g05185(.A1(new_n7597_), .A2(new_n7607_), .B(new_n7568_), .ZN(new_n7622_));
  NAND3_X1   g05186(.A1(new_n7622_), .A2(new_n5398_), .A3(new_n6764_), .ZN(new_n7623_));
  NOR2_X1    g05187(.A1(new_n7623_), .A2(new_n3369_), .ZN(new_n7624_));
  OAI21_X1   g05188(.A1(new_n7621_), .A2(new_n7624_), .B(pi0154), .ZN(new_n7625_));
  NOR2_X1    g05189(.A1(new_n7597_), .A2(new_n7605_), .ZN(new_n7626_));
  AOI21_X1   g05190(.A1(new_n7626_), .A2(new_n5427_), .B(new_n7583_), .ZN(new_n7627_));
  INV_X1     g05191(.I(new_n7627_), .ZN(new_n7628_));
  NOR3_X1    g05192(.A1(new_n7628_), .A2(pi0152), .A3(new_n5437_), .ZN(new_n7629_));
  AOI21_X1   g05193(.A1(new_n7608_), .A2(new_n5398_), .B(new_n7583_), .ZN(new_n7630_));
  NOR2_X1    g05194(.A1(new_n7630_), .A2(new_n5422_), .ZN(new_n7631_));
  NOR2_X1    g05195(.A1(new_n7631_), .A2(new_n7621_), .ZN(new_n7632_));
  OR3_X2     g05196(.A1(new_n7632_), .A2(pi0154), .A3(new_n7629_), .Z(new_n7633_));
  NAND3_X1   g05197(.A1(new_n7633_), .A2(new_n7508_), .A3(new_n7625_), .ZN(new_n7634_));
  AOI22_X1   g05198(.A1(new_n7634_), .A2(new_n7620_), .B1(new_n2628_), .B2(new_n7618_), .ZN(new_n7635_));
  NOR3_X1    g05199(.A1(new_n7635_), .A2(new_n7518_), .A3(new_n5666_), .ZN(new_n7636_));
  INV_X1     g05200(.I(new_n7620_), .ZN(new_n7637_));
  NOR2_X1    g05201(.A1(new_n7630_), .A2(new_n5446_), .ZN(new_n7638_));
  INV_X1     g05202(.I(new_n7638_), .ZN(new_n7639_));
  AOI21_X1   g05203(.A1(new_n7639_), .A2(new_n7609_), .B(new_n7610_), .ZN(new_n7640_));
  INV_X1     g05204(.I(new_n7640_), .ZN(new_n7641_));
  OAI22_X1   g05205(.A1(new_n7641_), .A2(pi0299), .B1(new_n7632_), .B2(new_n7637_), .ZN(new_n7642_));
  NAND2_X1   g05206(.A1(new_n7642_), .A2(new_n5666_), .ZN(new_n7643_));
  INV_X1     g05207(.I(new_n7643_), .ZN(new_n7644_));
  NAND2_X1   g05208(.A1(new_n7626_), .A2(new_n5450_), .ZN(new_n7645_));
  INV_X1     g05209(.I(new_n7645_), .ZN(new_n7646_));
  AOI21_X1   g05210(.A1(new_n7646_), .A2(new_n7519_), .B(new_n7583_), .ZN(new_n7647_));
  OR2_X2     g05211(.A1(new_n7647_), .A2(pi0299), .Z(new_n7648_));
  NAND2_X1   g05212(.A1(new_n7518_), .A2(pi0232), .ZN(new_n7649_));
  AOI21_X1   g05213(.A1(new_n7635_), .A2(new_n7648_), .B(new_n7649_), .ZN(new_n7650_));
  NOR4_X1    g05214(.A1(new_n7636_), .A2(new_n7650_), .A3(new_n2627_), .A4(new_n7644_), .ZN(new_n7651_));
  OAI21_X1   g05215(.A1(new_n7578_), .A2(new_n7409_), .B(pi0070), .ZN(new_n7652_));
  AOI21_X1   g05216(.A1(new_n2537_), .A2(new_n2496_), .B(pi0070), .ZN(new_n7653_));
  NOR2_X1    g05217(.A1(new_n7577_), .A2(pi0841), .ZN(new_n7654_));
  INV_X1     g05218(.I(new_n7654_), .ZN(new_n7655_));
  NAND2_X1   g05219(.A1(new_n7655_), .A2(new_n2496_), .ZN(new_n7656_));
  AOI21_X1   g05220(.A1(new_n7656_), .A2(pi0090), .B(new_n2537_), .ZN(new_n7657_));
  INV_X1     g05221(.I(new_n7657_), .ZN(new_n7658_));
  AOI21_X1   g05222(.A1(new_n7575_), .A2(new_n2496_), .B(new_n5359_), .ZN(new_n7659_));
  INV_X1     g05223(.I(new_n7659_), .ZN(new_n7660_));
  AOI21_X1   g05224(.A1(new_n7409_), .A2(new_n2792_), .B(new_n2785_), .ZN(new_n7661_));
  NAND2_X1   g05225(.A1(new_n7429_), .A2(new_n7661_), .ZN(new_n7662_));
  AOI21_X1   g05226(.A1(new_n2785_), .A2(new_n2496_), .B(pi0058), .ZN(new_n7663_));
  NAND2_X1   g05227(.A1(new_n7662_), .A2(new_n7663_), .ZN(new_n7664_));
  AOI21_X1   g05228(.A1(new_n7664_), .A2(new_n7660_), .B(pi0090), .ZN(new_n7665_));
  OAI21_X1   g05229(.A1(new_n7665_), .A2(new_n7658_), .B(new_n7653_), .ZN(new_n7666_));
  NAND2_X1   g05230(.A1(new_n7666_), .A2(new_n7652_), .ZN(new_n7667_));
  NOR2_X1    g05231(.A1(new_n3058_), .A2(pi0051), .ZN(new_n7668_));
  NOR2_X1    g05232(.A1(new_n7668_), .A2(new_n2496_), .ZN(new_n7669_));
  AOI21_X1   g05233(.A1(new_n7667_), .A2(new_n7668_), .B(new_n7669_), .ZN(new_n7670_));
  AOI21_X1   g05234(.A1(new_n7670_), .A2(new_n2818_), .B(pi0032), .ZN(new_n7671_));
  NOR2_X1    g05235(.A1(new_n7568_), .A2(new_n2725_), .ZN(new_n7672_));
  OAI21_X1   g05236(.A1(new_n7671_), .A2(new_n7672_), .B(new_n2462_), .ZN(new_n7673_));
  NOR2_X1    g05237(.A1(new_n7568_), .A2(new_n2462_), .ZN(new_n7674_));
  INV_X1     g05238(.I(new_n7674_), .ZN(new_n7675_));
  NAND2_X1   g05239(.A1(new_n7579_), .A2(new_n2496_), .ZN(new_n7676_));
  INV_X1     g05240(.I(new_n7676_), .ZN(new_n7677_));
  NOR2_X1    g05241(.A1(pi0040), .A2(pi0479), .ZN(new_n7678_));
  AOI22_X1   g05242(.A1(new_n7677_), .A2(new_n7678_), .B1(new_n3028_), .B2(new_n7675_), .ZN(new_n7679_));
  INV_X1     g05243(.I(new_n7679_), .ZN(new_n7680_));
  NAND2_X1   g05244(.A1(new_n7673_), .A2(new_n7680_), .ZN(new_n7681_));
  INV_X1     g05245(.I(new_n7469_), .ZN(new_n7682_));
  AOI21_X1   g05246(.A1(new_n7654_), .A2(new_n7682_), .B(new_n7583_), .ZN(new_n7683_));
  NOR2_X1    g05247(.A1(new_n7683_), .A2(new_n2725_), .ZN(new_n7684_));
  OAI21_X1   g05248(.A1(new_n7671_), .A2(new_n7684_), .B(new_n2462_), .ZN(new_n7685_));
  NOR2_X1    g05249(.A1(new_n7685_), .A2(new_n5351_), .ZN(new_n7686_));
  OAI21_X1   g05250(.A1(new_n7686_), .A2(new_n7681_), .B(new_n5666_), .ZN(new_n7687_));
  INV_X1     g05251(.I(new_n7687_), .ZN(new_n7688_));
  NOR2_X1    g05252(.A1(new_n2628_), .A2(pi0158), .ZN(new_n7689_));
  NOR2_X1    g05253(.A1(new_n7685_), .A2(pi0210), .ZN(new_n7690_));
  NOR2_X1    g05254(.A1(new_n7690_), .A2(new_n7681_), .ZN(new_n7691_));
  NOR2_X1    g05255(.A1(new_n7691_), .A2(new_n5398_), .ZN(new_n7692_));
  AOI21_X1   g05256(.A1(new_n5354_), .A2(new_n2496_), .B(pi0032), .ZN(new_n7693_));
  AOI21_X1   g05257(.A1(pi0093), .A2(new_n7409_), .B(new_n5354_), .ZN(new_n7694_));
  NAND2_X1   g05258(.A1(new_n7655_), .A2(pi0090), .ZN(new_n7695_));
  NAND2_X1   g05259(.A1(new_n7660_), .A2(new_n2985_), .ZN(new_n7696_));
  AOI21_X1   g05260(.A1(new_n7695_), .A2(new_n7696_), .B(new_n7409_), .ZN(new_n7697_));
  OAI21_X1   g05261(.A1(new_n7697_), .A2(pi0093), .B(new_n7694_), .ZN(new_n7698_));
  AOI21_X1   g05262(.A1(new_n7409_), .A2(pi0032), .B(pi0040), .ZN(new_n7699_));
  INV_X1     g05263(.I(new_n7699_), .ZN(new_n7700_));
  AOI21_X1   g05264(.A1(new_n7698_), .A2(new_n7693_), .B(new_n7700_), .ZN(new_n7701_));
  NOR2_X1    g05265(.A1(new_n7701_), .A2(pi0095), .ZN(new_n7702_));
  NOR2_X1    g05266(.A1(new_n7702_), .A2(new_n7679_), .ZN(new_n7703_));
  NOR2_X1    g05267(.A1(new_n7703_), .A2(new_n5437_), .ZN(new_n7704_));
  OAI21_X1   g05268(.A1(new_n7692_), .A2(new_n7704_), .B(new_n3369_), .ZN(new_n7705_));
  NAND2_X1   g05269(.A1(new_n7463_), .A2(new_n2985_), .ZN(new_n7706_));
  NAND2_X1   g05270(.A1(new_n7697_), .A2(new_n7706_), .ZN(new_n7707_));
  NAND2_X1   g05271(.A1(new_n7707_), .A2(new_n2771_), .ZN(new_n7708_));
  NAND2_X1   g05272(.A1(new_n7708_), .A2(new_n7694_), .ZN(new_n7709_));
  AOI21_X1   g05273(.A1(new_n7709_), .A2(new_n7693_), .B(new_n7700_), .ZN(new_n7710_));
  NOR2_X1    g05274(.A1(new_n7710_), .A2(pi0095), .ZN(new_n7711_));
  NOR2_X1    g05275(.A1(new_n7711_), .A2(new_n7679_), .ZN(new_n7712_));
  NOR2_X1    g05276(.A1(new_n7712_), .A2(new_n5437_), .ZN(new_n7713_));
  OAI21_X1   g05277(.A1(new_n7692_), .A2(new_n7713_), .B(pi0152), .ZN(new_n7714_));
  AOI21_X1   g05278(.A1(new_n7705_), .A2(new_n7714_), .B(pi0172), .ZN(new_n7715_));
  NOR3_X1    g05279(.A1(new_n7312_), .A2(new_n2741_), .A3(new_n5354_), .ZN(new_n7716_));
  INV_X1     g05280(.I(new_n7716_), .ZN(new_n7717_));
  OR3_X2     g05281(.A1(new_n7421_), .A2(pi0032), .A3(new_n7717_), .Z(new_n7718_));
  NAND2_X1   g05282(.A1(new_n7718_), .A2(new_n7568_), .ZN(new_n7719_));
  AOI21_X1   g05283(.A1(new_n7719_), .A2(new_n2462_), .B(new_n5437_), .ZN(new_n7720_));
  NAND2_X1   g05284(.A1(new_n7680_), .A2(new_n7720_), .ZN(new_n7721_));
  INV_X1     g05285(.I(new_n7691_), .ZN(new_n7722_));
  NOR2_X1    g05286(.A1(new_n7722_), .A2(new_n5398_), .ZN(new_n7723_));
  INV_X1     g05287(.I(new_n7723_), .ZN(new_n7724_));
  NAND3_X1   g05288(.A1(new_n7724_), .A2(pi0152), .A3(new_n7721_), .ZN(new_n7725_));
  AOI21_X1   g05289(.A1(new_n2462_), .A2(new_n7583_), .B(new_n7679_), .ZN(new_n7726_));
  NOR2_X1    g05290(.A1(new_n7726_), .A2(new_n5437_), .ZN(new_n7727_));
  OAI21_X1   g05291(.A1(new_n7692_), .A2(new_n7727_), .B(new_n3369_), .ZN(new_n7728_));
  AOI21_X1   g05292(.A1(new_n7725_), .A2(new_n7728_), .B(new_n3778_), .ZN(new_n7729_));
  OAI21_X1   g05293(.A1(new_n7729_), .A2(new_n7715_), .B(new_n7689_), .ZN(new_n7730_));
  NOR2_X1    g05294(.A1(new_n5631_), .A2(new_n2628_), .ZN(new_n7731_));
  NOR3_X1    g05295(.A1(new_n7711_), .A2(new_n5437_), .A3(new_n7674_), .ZN(new_n7732_));
  NOR2_X1    g05296(.A1(new_n7723_), .A2(new_n7732_), .ZN(new_n7733_));
  NAND2_X1   g05297(.A1(new_n7733_), .A2(pi0152), .ZN(new_n7734_));
  NOR3_X1    g05298(.A1(new_n7702_), .A2(new_n5437_), .A3(new_n7674_), .ZN(new_n7735_));
  NOR2_X1    g05299(.A1(new_n7723_), .A2(new_n7735_), .ZN(new_n7736_));
  NAND2_X1   g05300(.A1(new_n7736_), .A2(new_n3369_), .ZN(new_n7737_));
  AOI21_X1   g05301(.A1(new_n7734_), .A2(new_n7737_), .B(pi0172), .ZN(new_n7738_));
  NAND2_X1   g05302(.A1(new_n7568_), .A2(new_n5398_), .ZN(new_n7739_));
  NAND3_X1   g05303(.A1(new_n7724_), .A2(new_n3369_), .A3(new_n7739_), .ZN(new_n7740_));
  NAND2_X1   g05304(.A1(new_n7720_), .A2(new_n7675_), .ZN(new_n7741_));
  NAND3_X1   g05305(.A1(new_n7724_), .A2(pi0152), .A3(new_n7741_), .ZN(new_n7742_));
  AOI21_X1   g05306(.A1(new_n7740_), .A2(new_n7742_), .B(new_n3778_), .ZN(new_n7743_));
  OAI21_X1   g05307(.A1(new_n7738_), .A2(new_n7743_), .B(new_n7731_), .ZN(new_n7744_));
  NAND3_X1   g05308(.A1(new_n7744_), .A2(pi0149), .A3(new_n7730_), .ZN(new_n7745_));
  NOR2_X1    g05309(.A1(new_n3059_), .A2(new_n7568_), .ZN(new_n7746_));
  NAND2_X1   g05310(.A1(new_n3058_), .A2(new_n2496_), .ZN(new_n7747_));
  AOI21_X1   g05311(.A1(pi0051), .A2(new_n7409_), .B(new_n3058_), .ZN(new_n7748_));
  INV_X1     g05312(.I(new_n7652_), .ZN(new_n7749_));
  INV_X1     g05313(.I(new_n2522_), .ZN(new_n7750_));
  OAI22_X1   g05314(.A1(new_n7664_), .A2(new_n6677_), .B1(new_n2496_), .B2(new_n7750_), .ZN(new_n7751_));
  AOI21_X1   g05315(.A1(new_n7751_), .A2(new_n2835_), .B(new_n7749_), .ZN(new_n7752_));
  OAI21_X1   g05316(.A1(new_n7752_), .A2(pi0051), .B(new_n7748_), .ZN(new_n7753_));
  NAND3_X1   g05317(.A1(new_n7753_), .A2(new_n2818_), .A3(new_n7747_), .ZN(new_n7754_));
  NAND2_X1   g05318(.A1(new_n7754_), .A2(new_n2725_), .ZN(new_n7755_));
  NOR2_X1    g05319(.A1(new_n2496_), .A2(pi0040), .ZN(new_n7756_));
  NOR2_X1    g05320(.A1(new_n7756_), .A2(new_n2725_), .ZN(new_n7757_));
  INV_X1     g05321(.I(new_n7757_), .ZN(new_n7758_));
  NAND2_X1   g05322(.A1(new_n7755_), .A2(new_n7758_), .ZN(new_n7759_));
  INV_X1     g05323(.I(new_n7759_), .ZN(new_n7760_));
  OAI21_X1   g05324(.A1(new_n7760_), .A2(new_n7746_), .B(new_n2462_), .ZN(new_n7761_));
  AND2_X2    g05325(.A1(new_n7761_), .A2(new_n7675_), .Z(new_n7762_));
  OAI21_X1   g05326(.A1(new_n7683_), .A2(pi0040), .B(pi0032), .ZN(new_n7763_));
  AOI21_X1   g05327(.A1(new_n7755_), .A2(new_n7763_), .B(pi0095), .ZN(new_n7764_));
  NOR2_X1    g05328(.A1(new_n7756_), .A2(new_n2462_), .ZN(new_n7765_));
  OR2_X2     g05329(.A1(new_n7764_), .A2(new_n7765_), .Z(new_n7766_));
  NAND2_X1   g05330(.A1(new_n7762_), .A2(new_n7766_), .ZN(new_n7767_));
  AOI21_X1   g05331(.A1(new_n7767_), .A2(new_n2709_), .B(new_n5437_), .ZN(new_n7768_));
  AOI21_X1   g05332(.A1(new_n7768_), .A2(new_n7762_), .B(new_n7723_), .ZN(new_n7769_));
  NAND2_X1   g05333(.A1(new_n7769_), .A2(pi0152), .ZN(new_n7770_));
  INV_X1     g05334(.I(new_n7672_), .ZN(new_n7771_));
  INV_X1     g05335(.I(new_n7669_), .ZN(new_n7772_));
  AOI21_X1   g05336(.A1(new_n7428_), .A2(new_n7570_), .B(new_n7409_), .ZN(new_n7773_));
  NOR2_X1    g05337(.A1(new_n7773_), .A2(pi0058), .ZN(new_n7774_));
  AOI22_X1   g05338(.A1(new_n7774_), .A2(new_n6676_), .B1(new_n7409_), .B2(new_n2522_), .ZN(new_n7775_));
  OAI21_X1   g05339(.A1(new_n7775_), .A2(pi0070), .B(new_n7652_), .ZN(new_n7776_));
  NAND2_X1   g05340(.A1(new_n7776_), .A2(new_n7668_), .ZN(new_n7777_));
  NAND2_X1   g05341(.A1(new_n7777_), .A2(new_n7772_), .ZN(new_n7778_));
  NOR2_X1    g05342(.A1(new_n7778_), .A2(pi0040), .ZN(new_n7779_));
  NOR2_X1    g05343(.A1(new_n7779_), .A2(pi0032), .ZN(new_n7780_));
  INV_X1     g05344(.I(new_n7780_), .ZN(new_n7781_));
  AOI21_X1   g05345(.A1(new_n7781_), .A2(new_n7771_), .B(pi0095), .ZN(new_n7782_));
  INV_X1     g05346(.I(new_n7684_), .ZN(new_n7783_));
  AOI21_X1   g05347(.A1(new_n7781_), .A2(new_n7783_), .B(pi0095), .ZN(new_n7784_));
  OAI21_X1   g05348(.A1(new_n7784_), .A2(new_n7674_), .B(new_n2709_), .ZN(new_n7785_));
  NAND2_X1   g05349(.A1(new_n7785_), .A2(new_n5398_), .ZN(new_n7786_));
  OR3_X2     g05350(.A1(new_n7786_), .A2(new_n7674_), .A3(new_n7782_), .Z(new_n7787_));
  NAND3_X1   g05351(.A1(new_n7787_), .A2(new_n7724_), .A3(new_n3369_), .ZN(new_n7788_));
  AOI21_X1   g05352(.A1(new_n7770_), .A2(new_n7788_), .B(new_n3778_), .ZN(new_n7789_));
  INV_X1     g05353(.I(new_n7653_), .ZN(new_n7790_));
  OAI21_X1   g05354(.A1(new_n7773_), .A2(pi0058), .B(new_n7660_), .ZN(new_n7791_));
  AOI21_X1   g05355(.A1(new_n7791_), .A2(new_n2985_), .B(new_n7658_), .ZN(new_n7792_));
  OAI21_X1   g05356(.A1(new_n7792_), .A2(new_n7790_), .B(new_n7652_), .ZN(new_n7793_));
  AOI21_X1   g05357(.A1(new_n7793_), .A2(new_n7668_), .B(new_n7669_), .ZN(new_n7794_));
  INV_X1     g05358(.I(new_n7794_), .ZN(new_n7795_));
  OAI21_X1   g05359(.A1(new_n7795_), .A2(pi0040), .B(new_n2725_), .ZN(new_n7796_));
  AOI21_X1   g05360(.A1(new_n7796_), .A2(new_n7771_), .B(pi0095), .ZN(new_n7797_));
  NOR3_X1    g05361(.A1(new_n7797_), .A2(new_n5437_), .A3(new_n7674_), .ZN(new_n7798_));
  AOI21_X1   g05362(.A1(new_n7796_), .A2(new_n7783_), .B(pi0095), .ZN(new_n7799_));
  INV_X1     g05363(.I(new_n7799_), .ZN(new_n7800_));
  NOR2_X1    g05364(.A1(new_n7800_), .A2(pi0210), .ZN(new_n7801_));
  INV_X1     g05365(.I(new_n7801_), .ZN(new_n7802_));
  AOI21_X1   g05366(.A1(new_n7798_), .A2(new_n7802_), .B(new_n7723_), .ZN(new_n7803_));
  NAND2_X1   g05367(.A1(new_n7803_), .A2(new_n3369_), .ZN(new_n7804_));
  NAND2_X1   g05368(.A1(new_n7673_), .A2(new_n7675_), .ZN(new_n7805_));
  NOR2_X1    g05369(.A1(new_n7690_), .A2(new_n7805_), .ZN(new_n7806_));
  AOI21_X1   g05370(.A1(new_n5398_), .A2(new_n7806_), .B(new_n7723_), .ZN(new_n7807_));
  NAND2_X1   g05371(.A1(new_n7807_), .A2(pi0152), .ZN(new_n7808_));
  AOI21_X1   g05372(.A1(new_n7804_), .A2(new_n7808_), .B(pi0172), .ZN(new_n7809_));
  OAI21_X1   g05373(.A1(new_n7789_), .A2(new_n7809_), .B(new_n7731_), .ZN(new_n7810_));
  NOR2_X1    g05374(.A1(new_n7722_), .A2(new_n3369_), .ZN(new_n7811_));
  NOR2_X1    g05375(.A1(new_n7797_), .A2(new_n7679_), .ZN(new_n7812_));
  INV_X1     g05376(.I(new_n7812_), .ZN(new_n7813_));
  NOR2_X1    g05377(.A1(new_n7801_), .A2(new_n7813_), .ZN(new_n7814_));
  INV_X1     g05378(.I(new_n7814_), .ZN(new_n7815_));
  NOR3_X1    g05379(.A1(new_n7815_), .A2(pi0152), .A3(new_n5437_), .ZN(new_n7816_));
  OAI21_X1   g05380(.A1(new_n7816_), .A2(new_n7811_), .B(new_n3778_), .ZN(new_n7817_));
  NAND2_X1   g05381(.A1(new_n7761_), .A2(new_n7680_), .ZN(new_n7818_));
  INV_X1     g05382(.I(new_n7818_), .ZN(new_n7819_));
  NOR2_X1    g05383(.A1(new_n7568_), .A2(new_n5437_), .ZN(new_n7820_));
  OAI21_X1   g05384(.A1(new_n7768_), .A2(new_n7820_), .B(new_n7819_), .ZN(new_n7821_));
  NOR2_X1    g05385(.A1(new_n7821_), .A2(new_n3369_), .ZN(new_n7822_));
  INV_X1     g05386(.I(new_n7820_), .ZN(new_n7823_));
  NOR2_X1    g05387(.A1(new_n7782_), .A2(new_n7679_), .ZN(new_n7824_));
  INV_X1     g05388(.I(new_n7824_), .ZN(new_n7825_));
  AOI21_X1   g05389(.A1(new_n7786_), .A2(new_n7823_), .B(new_n7825_), .ZN(new_n7826_));
  INV_X1     g05390(.I(new_n7826_), .ZN(new_n7827_));
  NOR2_X1    g05391(.A1(new_n7827_), .A2(pi0152), .ZN(new_n7828_));
  OAI21_X1   g05392(.A1(new_n7822_), .A2(new_n7828_), .B(pi0172), .ZN(new_n7829_));
  NAND4_X1   g05393(.A1(new_n7829_), .A2(new_n7689_), .A3(new_n7724_), .A4(new_n7817_), .ZN(new_n7830_));
  NAND3_X1   g05394(.A1(new_n7830_), .A2(new_n7810_), .A3(new_n7455_), .ZN(new_n7831_));
  NAND2_X1   g05395(.A1(new_n7831_), .A2(new_n7745_), .ZN(new_n7832_));
  NOR2_X1    g05396(.A1(new_n7685_), .A2(pi0198), .ZN(new_n7833_));
  NOR2_X1    g05397(.A1(new_n7833_), .A2(new_n7681_), .ZN(new_n7834_));
  INV_X1     g05398(.I(new_n7834_), .ZN(new_n7835_));
  NOR2_X1    g05399(.A1(new_n7835_), .A2(new_n5398_), .ZN(new_n7836_));
  NOR2_X1    g05400(.A1(new_n7836_), .A2(new_n7732_), .ZN(new_n7837_));
  NAND2_X1   g05401(.A1(new_n7837_), .A2(pi0183), .ZN(new_n7838_));
  NOR2_X1    g05402(.A1(new_n5437_), .A2(pi0040), .ZN(new_n7839_));
  NOR2_X1    g05403(.A1(new_n7833_), .A2(new_n7805_), .ZN(new_n7840_));
  AOI21_X1   g05404(.A1(new_n7839_), .A2(new_n7840_), .B(new_n7836_), .ZN(new_n7841_));
  NAND2_X1   g05405(.A1(new_n7841_), .A2(new_n7479_), .ZN(new_n7842_));
  AOI21_X1   g05406(.A1(new_n7842_), .A2(new_n7838_), .B(new_n7488_), .ZN(new_n7843_));
  OR2_X2     g05407(.A1(new_n7836_), .A2(new_n7735_), .Z(new_n7844_));
  NOR2_X1    g05408(.A1(new_n7844_), .A2(new_n7479_), .ZN(new_n7845_));
  NOR2_X1    g05409(.A1(new_n7800_), .A2(pi0198), .ZN(new_n7846_));
  INV_X1     g05410(.I(new_n7846_), .ZN(new_n7847_));
  AOI21_X1   g05411(.A1(new_n7798_), .A2(new_n7847_), .B(new_n7836_), .ZN(new_n7848_));
  AOI21_X1   g05412(.A1(new_n7479_), .A2(new_n7848_), .B(new_n7845_), .ZN(new_n7849_));
  NOR2_X1    g05413(.A1(new_n7849_), .A2(pi0174), .ZN(new_n7850_));
  OAI21_X1   g05414(.A1(new_n7850_), .A2(new_n7843_), .B(pi0180), .ZN(new_n7851_));
  OAI21_X1   g05415(.A1(new_n7849_), .A2(pi0095), .B(new_n7488_), .ZN(new_n7852_));
  AOI21_X1   g05416(.A1(new_n7713_), .A2(pi0183), .B(new_n7488_), .ZN(new_n7853_));
  NAND2_X1   g05417(.A1(new_n7835_), .A2(new_n7495_), .ZN(new_n7854_));
  AOI21_X1   g05418(.A1(new_n7854_), .A2(new_n7853_), .B(pi0180), .ZN(new_n7855_));
  OAI21_X1   g05419(.A1(new_n7852_), .A2(new_n7679_), .B(new_n7855_), .ZN(new_n7856_));
  AOI21_X1   g05420(.A1(new_n7856_), .A2(new_n7851_), .B(pi0193), .ZN(new_n7857_));
  INV_X1     g05421(.I(pi0193), .ZN(new_n7858_));
  AOI21_X1   g05422(.A1(new_n7778_), .A2(new_n2818_), .B(pi0032), .ZN(new_n7859_));
  INV_X1     g05423(.I(new_n7859_), .ZN(new_n7860_));
  AOI21_X1   g05424(.A1(new_n7860_), .A2(new_n7758_), .B(pi0095), .ZN(new_n7861_));
  NOR2_X1    g05425(.A1(new_n7861_), .A2(new_n7765_), .ZN(new_n7862_));
  AOI21_X1   g05426(.A1(new_n7860_), .A2(new_n7763_), .B(pi0095), .ZN(new_n7863_));
  NOR3_X1    g05427(.A1(new_n7863_), .A2(pi0198), .A3(new_n7765_), .ZN(new_n7864_));
  AOI21_X1   g05428(.A1(pi0198), .A2(new_n7862_), .B(new_n7864_), .ZN(new_n7865_));
  AOI21_X1   g05429(.A1(new_n7865_), .A2(new_n7839_), .B(new_n7836_), .ZN(new_n7866_));
  NAND2_X1   g05430(.A1(new_n7866_), .A2(new_n7479_), .ZN(new_n7867_));
  INV_X1     g05431(.I(new_n7836_), .ZN(new_n7868_));
  NAND3_X1   g05432(.A1(new_n7868_), .A2(pi0183), .A3(new_n7739_), .ZN(new_n7869_));
  AOI21_X1   g05433(.A1(new_n7867_), .A2(new_n7869_), .B(pi0174), .ZN(new_n7870_));
  NAND3_X1   g05434(.A1(new_n7868_), .A2(pi0183), .A3(new_n7741_), .ZN(new_n7871_));
  AOI21_X1   g05435(.A1(new_n7767_), .A2(new_n2672_), .B(new_n5437_), .ZN(new_n7872_));
  AOI21_X1   g05436(.A1(new_n7872_), .A2(new_n7762_), .B(new_n7836_), .ZN(new_n7873_));
  NAND2_X1   g05437(.A1(new_n7873_), .A2(new_n7479_), .ZN(new_n7874_));
  AOI21_X1   g05438(.A1(new_n7874_), .A2(new_n7871_), .B(new_n7488_), .ZN(new_n7875_));
  NOR3_X1    g05439(.A1(new_n7875_), .A2(new_n5657_), .A3(new_n7870_), .ZN(new_n7876_));
  INV_X1     g05440(.I(new_n7721_), .ZN(new_n7877_));
  NOR2_X1    g05441(.A1(new_n7836_), .A2(new_n7877_), .ZN(new_n7878_));
  NAND2_X1   g05442(.A1(new_n7878_), .A2(pi0183), .ZN(new_n7879_));
  OAI21_X1   g05443(.A1(new_n7872_), .A2(new_n7820_), .B(new_n7819_), .ZN(new_n7880_));
  NAND3_X1   g05444(.A1(new_n7880_), .A2(new_n7479_), .A3(new_n7868_), .ZN(new_n7881_));
  AOI21_X1   g05445(.A1(new_n7881_), .A2(new_n7879_), .B(new_n7488_), .ZN(new_n7882_));
  AOI21_X1   g05446(.A1(new_n2672_), .A2(new_n7784_), .B(new_n7825_), .ZN(new_n7883_));
  AOI21_X1   g05447(.A1(new_n5398_), .A2(new_n7883_), .B(new_n7836_), .ZN(new_n7884_));
  AND2_X2    g05448(.A1(new_n7884_), .A2(new_n7479_), .Z(new_n7885_));
  AOI21_X1   g05449(.A1(new_n7835_), .A2(new_n5437_), .B(new_n7727_), .ZN(new_n7886_));
  NOR2_X1    g05450(.A1(new_n7886_), .A2(new_n7479_), .ZN(new_n7887_));
  OAI21_X1   g05451(.A1(new_n7885_), .A2(new_n7887_), .B(new_n7488_), .ZN(new_n7888_));
  NAND2_X1   g05452(.A1(new_n7888_), .A2(new_n5657_), .ZN(new_n7889_));
  NOR2_X1    g05453(.A1(new_n7882_), .A2(new_n7889_), .ZN(new_n7890_));
  NOR3_X1    g05454(.A1(new_n7890_), .A2(new_n7876_), .A3(new_n7858_), .ZN(new_n7891_));
  OAI21_X1   g05455(.A1(new_n7857_), .A2(new_n7891_), .B(new_n2628_), .ZN(new_n7892_));
  AOI21_X1   g05456(.A1(new_n7892_), .A2(new_n7832_), .B(new_n5666_), .ZN(new_n7893_));
  NOR3_X1    g05457(.A1(new_n7893_), .A2(pi0039), .A3(new_n7688_), .ZN(new_n7894_));
  NOR3_X1    g05458(.A1(new_n7894_), .A2(pi0038), .A3(new_n7651_), .ZN(new_n7895_));
  NOR3_X1    g05459(.A1(new_n7895_), .A2(pi0100), .A3(new_n7407_), .ZN(new_n7896_));
  NOR3_X1    g05460(.A1(new_n7896_), .A2(pi0087), .A3(new_n7372_), .ZN(new_n7897_));
  OAI21_X1   g05461(.A1(new_n7583_), .A2(new_n3271_), .B(pi0087), .ZN(new_n7898_));
  OAI21_X1   g05462(.A1(new_n7390_), .A2(new_n7898_), .B(new_n2605_), .ZN(new_n7899_));
  OAI21_X1   g05463(.A1(new_n7897_), .A2(new_n7899_), .B(new_n7604_), .ZN(new_n7900_));
  AOI21_X1   g05464(.A1(new_n7900_), .A2(new_n5499_), .B(new_n7386_), .ZN(new_n7901_));
  OAI21_X1   g05465(.A1(new_n7901_), .A2(pi0074), .B(new_n7380_), .ZN(new_n7902_));
  NAND3_X1   g05466(.A1(new_n7902_), .A2(new_n2470_), .A3(new_n7595_), .ZN(new_n7903_));
  NOR3_X1    g05467(.A1(new_n7585_), .A2(new_n2563_), .A3(new_n7348_), .ZN(new_n7904_));
  INV_X1     g05468(.I(new_n7904_), .ZN(new_n7905_));
  NOR2_X1    g05469(.A1(new_n7905_), .A2(new_n2470_), .ZN(new_n7906_));
  NOR2_X1    g05470(.A1(new_n7366_), .A2(new_n7906_), .ZN(new_n7907_));
  AOI21_X1   g05471(.A1(new_n7903_), .A2(new_n7907_), .B(new_n7356_), .ZN(new_n7908_));
  NAND2_X1   g05472(.A1(new_n7908_), .A2(new_n7565_), .ZN(new_n7909_));
  OAI21_X1   g05473(.A1(new_n7557_), .A2(new_n7565_), .B(new_n7909_), .ZN(new_n7910_));
  NOR2_X1    g05474(.A1(new_n7557_), .A2(new_n7558_), .ZN(new_n7911_));
  AOI21_X1   g05475(.A1(new_n7908_), .A2(new_n7558_), .B(new_n7911_), .ZN(new_n7912_));
  NOR2_X1    g05476(.A1(new_n7912_), .A2(po1110), .ZN(new_n7913_));
  AOI21_X1   g05477(.A1(new_n7910_), .A2(po1110), .B(new_n7913_), .ZN(po0191));
  NOR2_X1    g05478(.A1(pi0033), .A2(pi0954), .ZN(new_n7915_));
  NOR2_X1    g05479(.A1(pi0149), .A2(pi0157), .ZN(new_n7916_));
  XNOR2_X1   g05480(.A1(pi0162), .A2(pi0197), .ZN(new_n7917_));
  NAND2_X1   g05481(.A1(new_n7917_), .A2(new_n7916_), .ZN(new_n7918_));
  OR2_X2     g05482(.A1(new_n7917_), .A2(new_n7916_), .Z(new_n7919_));
  NAND4_X1   g05483(.A1(new_n7919_), .A2(pi0232), .A3(new_n5398_), .A4(new_n7918_), .ZN(new_n7920_));
  NOR2_X1    g05484(.A1(new_n7920_), .A2(new_n7342_), .ZN(new_n7921_));
  INV_X1     g05485(.I(new_n7921_), .ZN(new_n7922_));
  AOI21_X1   g05486(.A1(new_n7349_), .A2(pi0148), .B(new_n2625_), .ZN(new_n7923_));
  NAND2_X1   g05487(.A1(new_n7922_), .A2(new_n7923_), .ZN(new_n7924_));
  INV_X1     g05488(.I(pi0167), .ZN(new_n7925_));
  NOR2_X1    g05489(.A1(new_n7350_), .A2(new_n7925_), .ZN(new_n7926_));
  NOR2_X1    g05490(.A1(new_n7921_), .A2(new_n7926_), .ZN(new_n7927_));
  NAND2_X1   g05491(.A1(new_n7927_), .A2(new_n2625_), .ZN(new_n7928_));
  NAND2_X1   g05492(.A1(new_n7928_), .A2(new_n7924_), .ZN(new_n7929_));
  INV_X1     g05493(.I(new_n7929_), .ZN(new_n7930_));
  NAND2_X1   g05494(.A1(new_n7930_), .A2(new_n3425_), .ZN(new_n7931_));
  NOR2_X1    g05495(.A1(pi0178), .A2(pi0183), .ZN(new_n7932_));
  NOR2_X1    g05496(.A1(new_n5437_), .A2(new_n7932_), .ZN(new_n7933_));
  INV_X1     g05497(.I(pi0140), .ZN(new_n7934_));
  NOR2_X1    g05498(.A1(new_n7934_), .A2(new_n5656_), .ZN(new_n7935_));
  INV_X1     g05499(.I(new_n7935_), .ZN(new_n7936_));
  NAND2_X1   g05500(.A1(new_n7934_), .A2(new_n5656_), .ZN(new_n7937_));
  NAND2_X1   g05501(.A1(new_n7936_), .A2(new_n7937_), .ZN(new_n7938_));
  NAND2_X1   g05502(.A1(new_n7938_), .A2(new_n7933_), .ZN(new_n7939_));
  NAND2_X1   g05503(.A1(new_n7936_), .A2(new_n7932_), .ZN(new_n7940_));
  INV_X1     g05504(.I(new_n7940_), .ZN(new_n7941_));
  NAND3_X1   g05505(.A1(new_n7941_), .A2(new_n5398_), .A3(new_n7937_), .ZN(new_n7942_));
  NAND3_X1   g05506(.A1(new_n7942_), .A2(new_n2628_), .A3(new_n7939_), .ZN(new_n7943_));
  NAND3_X1   g05507(.A1(new_n7919_), .A2(new_n5398_), .A3(new_n7918_), .ZN(new_n7944_));
  AOI21_X1   g05508(.A1(new_n7944_), .A2(pi0299), .B(new_n5666_), .ZN(new_n7945_));
  NAND2_X1   g05509(.A1(new_n7945_), .A2(new_n7943_), .ZN(new_n7946_));
  NAND2_X1   g05510(.A1(new_n7946_), .A2(pi0100), .ZN(new_n7947_));
  INV_X1     g05511(.I(new_n7947_), .ZN(new_n7948_));
  NAND2_X1   g05512(.A1(new_n7946_), .A2(pi0075), .ZN(new_n7949_));
  INV_X1     g05513(.I(new_n7949_), .ZN(new_n7950_));
  NOR2_X1    g05514(.A1(new_n7948_), .A2(new_n7950_), .ZN(new_n7951_));
  NOR2_X1    g05515(.A1(pi0141), .A2(pi0299), .ZN(new_n7952_));
  AOI21_X1   g05516(.A1(new_n4257_), .A2(pi0299), .B(new_n7952_), .ZN(new_n7953_));
  INV_X1     g05517(.I(new_n7953_), .ZN(new_n7954_));
  NOR2_X1    g05518(.A1(new_n6698_), .A2(new_n7954_), .ZN(new_n7955_));
  OAI21_X1   g05519(.A1(new_n7348_), .A2(new_n7955_), .B(new_n7951_), .ZN(new_n7956_));
  AOI21_X1   g05520(.A1(new_n7956_), .A2(pi0074), .B(pi0055), .ZN(new_n7957_));
  INV_X1     g05521(.I(pi0188), .ZN(new_n7958_));
  NOR2_X1    g05522(.A1(new_n7958_), .A2(pi0299), .ZN(new_n7959_));
  AOI21_X1   g05523(.A1(pi0167), .A2(pi0299), .B(new_n7959_), .ZN(new_n7960_));
  NOR2_X1    g05524(.A1(new_n6698_), .A2(new_n7960_), .ZN(new_n7961_));
  NOR2_X1    g05525(.A1(new_n7961_), .A2(pi0100), .ZN(new_n7962_));
  INV_X1     g05526(.I(new_n7962_), .ZN(new_n7963_));
  NOR2_X1    g05527(.A1(new_n7963_), .A2(pi0075), .ZN(new_n7964_));
  INV_X1     g05528(.I(new_n7964_), .ZN(new_n7965_));
  AOI21_X1   g05529(.A1(new_n7951_), .A2(new_n7965_), .B(new_n5499_), .ZN(new_n7966_));
  AOI21_X1   g05530(.A1(new_n7961_), .A2(pi0038), .B(new_n7584_), .ZN(new_n7967_));
  INV_X1     g05531(.I(pi0155), .ZN(new_n7968_));
  NOR2_X1    g05532(.A1(pi0177), .A2(pi0299), .ZN(new_n7969_));
  AOI21_X1   g05533(.A1(new_n7968_), .A2(pi0299), .B(new_n7969_), .ZN(new_n7970_));
  OAI21_X1   g05534(.A1(pi0038), .A2(new_n7970_), .B(new_n6697_), .ZN(new_n7971_));
  AOI21_X1   g05535(.A1(new_n7600_), .A2(new_n7971_), .B(new_n7967_), .ZN(new_n7972_));
  OAI21_X1   g05536(.A1(new_n7972_), .A2(pi0100), .B(new_n7947_), .ZN(new_n7973_));
  NAND2_X1   g05537(.A1(new_n7973_), .A2(new_n7387_), .ZN(new_n7974_));
  NOR2_X1    g05538(.A1(new_n7925_), .A2(new_n7958_), .ZN(new_n7975_));
  AOI22_X1   g05539(.A1(new_n7401_), .A2(new_n7958_), .B1(new_n7398_), .B2(new_n7975_), .ZN(new_n7976_));
  NOR2_X1    g05540(.A1(new_n7405_), .A2(new_n7958_), .ZN(new_n7977_));
  NOR2_X1    g05541(.A1(new_n7977_), .A2(pi0167), .ZN(new_n7978_));
  INV_X1     g05542(.I(new_n7978_), .ZN(new_n7979_));
  AOI21_X1   g05543(.A1(new_n7979_), .A2(new_n7976_), .B(new_n3265_), .ZN(new_n7980_));
  NAND2_X1   g05544(.A1(pi0159), .A2(pi0299), .ZN(new_n7981_));
  NOR3_X1    g05545(.A1(new_n7723_), .A2(new_n3107_), .A3(new_n7732_), .ZN(new_n7982_));
  AND3_X2    g05546(.A1(new_n7724_), .A2(new_n3107_), .A3(new_n7741_), .Z(new_n7983_));
  OAI21_X1   g05547(.A1(new_n7983_), .A2(new_n7982_), .B(pi0161), .ZN(new_n7984_));
  INV_X1     g05548(.I(pi0162), .ZN(new_n7985_));
  NAND3_X1   g05549(.A1(new_n7724_), .A2(new_n3107_), .A3(new_n7739_), .ZN(new_n7986_));
  NAND2_X1   g05550(.A1(new_n7736_), .A2(pi0146), .ZN(new_n7987_));
  NAND2_X1   g05551(.A1(new_n7987_), .A2(new_n7986_), .ZN(new_n7988_));
  AOI21_X1   g05552(.A1(new_n7988_), .A2(new_n3360_), .B(new_n7985_), .ZN(new_n7989_));
  AOI21_X1   g05553(.A1(new_n7989_), .A2(new_n7984_), .B(new_n7981_), .ZN(new_n7990_));
  AND2_X2    g05554(.A1(new_n7807_), .A2(pi0146), .Z(new_n7991_));
  AOI21_X1   g05555(.A1(new_n7769_), .A2(new_n3107_), .B(new_n7991_), .ZN(new_n7992_));
  NAND2_X1   g05556(.A1(new_n7803_), .A2(pi0146), .ZN(new_n7993_));
  NAND3_X1   g05557(.A1(new_n7787_), .A2(new_n7724_), .A3(new_n3107_), .ZN(new_n7994_));
  NAND2_X1   g05558(.A1(new_n7993_), .A2(new_n7994_), .ZN(new_n7995_));
  AOI21_X1   g05559(.A1(new_n7995_), .A2(new_n3360_), .B(pi0162), .ZN(new_n7996_));
  OAI21_X1   g05560(.A1(new_n3360_), .A2(new_n7992_), .B(new_n7996_), .ZN(new_n7997_));
  NAND2_X1   g05561(.A1(new_n7997_), .A2(new_n7990_), .ZN(new_n7998_));
  NOR2_X1    g05562(.A1(new_n7884_), .A2(pi0142), .ZN(new_n7999_));
  OAI21_X1   g05563(.A1(new_n7834_), .A2(new_n5398_), .B(pi0142), .ZN(new_n8000_));
  NOR2_X1    g05564(.A1(new_n7846_), .A2(new_n7813_), .ZN(new_n8001_));
  INV_X1     g05565(.I(new_n8001_), .ZN(new_n8002_));
  AOI21_X1   g05566(.A1(new_n8002_), .A2(new_n5398_), .B(new_n8000_), .ZN(new_n8003_));
  NOR3_X1    g05567(.A1(new_n7999_), .A2(new_n8003_), .A3(pi0140), .ZN(new_n8004_));
  OAI21_X1   g05568(.A1(new_n8000_), .A2(new_n7704_), .B(pi0140), .ZN(new_n8005_));
  AOI21_X1   g05569(.A1(new_n2724_), .A2(new_n7886_), .B(new_n8005_), .ZN(new_n8006_));
  OAI21_X1   g05570(.A1(new_n8004_), .A2(new_n8006_), .B(new_n5658_), .ZN(new_n8007_));
  AND3_X2    g05571(.A1(new_n7868_), .A2(new_n2724_), .A3(new_n7739_), .Z(new_n8008_));
  NOR2_X1    g05572(.A1(new_n7844_), .A2(new_n2724_), .ZN(new_n8009_));
  OAI21_X1   g05573(.A1(new_n8009_), .A2(new_n8008_), .B(pi0140), .ZN(new_n8010_));
  AND2_X2    g05574(.A1(new_n7848_), .A2(pi0142), .Z(new_n8011_));
  AND2_X2    g05575(.A1(new_n7866_), .A2(new_n2724_), .Z(new_n8012_));
  OAI21_X1   g05576(.A1(new_n8012_), .A2(new_n8011_), .B(new_n7934_), .ZN(new_n8013_));
  NAND2_X1   g05577(.A1(new_n8013_), .A2(new_n8010_), .ZN(new_n8014_));
  AOI21_X1   g05578(.A1(new_n8014_), .A2(pi0181), .B(pi0144), .ZN(new_n8015_));
  AOI21_X1   g05579(.A1(new_n8015_), .A2(new_n8007_), .B(pi0299), .ZN(new_n8016_));
  NAND2_X1   g05580(.A1(new_n7837_), .A2(pi0142), .ZN(new_n8017_));
  NAND3_X1   g05581(.A1(new_n7868_), .A2(new_n2724_), .A3(new_n7741_), .ZN(new_n8018_));
  AOI21_X1   g05582(.A1(new_n8017_), .A2(new_n8018_), .B(new_n7934_), .ZN(new_n8019_));
  NAND2_X1   g05583(.A1(new_n7841_), .A2(pi0142), .ZN(new_n8020_));
  NAND2_X1   g05584(.A1(new_n7873_), .A2(new_n2724_), .ZN(new_n8021_));
  AOI21_X1   g05585(.A1(new_n8021_), .A2(new_n8020_), .B(pi0140), .ZN(new_n8022_));
  OAI21_X1   g05586(.A1(new_n8022_), .A2(new_n8019_), .B(pi0181), .ZN(new_n8023_));
  NAND3_X1   g05587(.A1(new_n7880_), .A2(new_n2724_), .A3(new_n7868_), .ZN(new_n8024_));
  NAND2_X1   g05588(.A1(new_n7835_), .A2(pi0142), .ZN(new_n8025_));
  AOI21_X1   g05589(.A1(new_n8024_), .A2(new_n8025_), .B(pi0140), .ZN(new_n8026_));
  OAI21_X1   g05590(.A1(new_n8000_), .A2(new_n7713_), .B(pi0140), .ZN(new_n8027_));
  NOR2_X1    g05591(.A1(new_n7878_), .A2(pi0142), .ZN(new_n8028_));
  NOR2_X1    g05592(.A1(new_n8028_), .A2(new_n8027_), .ZN(new_n8029_));
  OAI21_X1   g05593(.A1(new_n8026_), .A2(new_n8029_), .B(new_n5658_), .ZN(new_n8030_));
  NAND3_X1   g05594(.A1(new_n8030_), .A2(new_n8023_), .A3(pi0144), .ZN(new_n8031_));
  NAND2_X1   g05595(.A1(new_n8016_), .A2(new_n8031_), .ZN(new_n8032_));
  NOR2_X1    g05596(.A1(new_n2628_), .A2(pi0159), .ZN(new_n8033_));
  NAND2_X1   g05597(.A1(new_n7691_), .A2(pi0161), .ZN(new_n8034_));
  NOR2_X1    g05598(.A1(new_n7815_), .A2(new_n5437_), .ZN(new_n8035_));
  NAND2_X1   g05599(.A1(new_n8035_), .A2(new_n3360_), .ZN(new_n8036_));
  AOI21_X1   g05600(.A1(new_n8036_), .A2(new_n8034_), .B(new_n3107_), .ZN(new_n8037_));
  OR2_X2     g05601(.A1(new_n7821_), .A2(new_n3360_), .Z(new_n8038_));
  NAND2_X1   g05602(.A1(new_n7826_), .A2(new_n3360_), .ZN(new_n8039_));
  AOI21_X1   g05603(.A1(new_n8038_), .A2(new_n8039_), .B(pi0146), .ZN(new_n8040_));
  NOR4_X1    g05604(.A1(new_n8040_), .A2(pi0162), .A3(new_n7723_), .A4(new_n8037_), .ZN(new_n8041_));
  NOR2_X1    g05605(.A1(new_n7692_), .A2(new_n7704_), .ZN(new_n8042_));
  NOR2_X1    g05606(.A1(new_n8042_), .A2(new_n3107_), .ZN(new_n8043_));
  NOR2_X1    g05607(.A1(new_n7692_), .A2(new_n7727_), .ZN(new_n8044_));
  NOR2_X1    g05608(.A1(new_n8044_), .A2(pi0146), .ZN(new_n8045_));
  OAI21_X1   g05609(.A1(new_n8043_), .A2(new_n8045_), .B(new_n3360_), .ZN(new_n8046_));
  NOR2_X1    g05610(.A1(new_n7692_), .A2(new_n7713_), .ZN(new_n8047_));
  NOR2_X1    g05611(.A1(new_n8047_), .A2(new_n3107_), .ZN(new_n8048_));
  NOR3_X1    g05612(.A1(new_n7723_), .A2(pi0146), .A3(new_n7877_), .ZN(new_n8049_));
  OAI21_X1   g05613(.A1(new_n8048_), .A2(new_n8049_), .B(pi0161), .ZN(new_n8050_));
  AOI21_X1   g05614(.A1(new_n8046_), .A2(new_n8050_), .B(new_n7985_), .ZN(new_n8051_));
  OAI21_X1   g05615(.A1(new_n8041_), .A2(new_n8051_), .B(new_n8033_), .ZN(new_n8052_));
  NAND3_X1   g05616(.A1(new_n8032_), .A2(new_n7998_), .A3(new_n8052_), .ZN(new_n8053_));
  NAND2_X1   g05617(.A1(new_n8053_), .A2(pi0232), .ZN(new_n8054_));
  AOI21_X1   g05618(.A1(new_n8054_), .A2(new_n7687_), .B(new_n2573_), .ZN(new_n8055_));
  INV_X1     g05619(.I(pi0177), .ZN(new_n8056_));
  NOR2_X1    g05620(.A1(new_n8056_), .A2(pi0299), .ZN(new_n8057_));
  INV_X1     g05621(.I(pi0144), .ZN(new_n8058_));
  NOR4_X1    g05622(.A1(new_n7615_), .A2(new_n8058_), .A3(new_n5446_), .A4(new_n7610_), .ZN(new_n8059_));
  OAI21_X1   g05623(.A1(new_n7611_), .A2(new_n8059_), .B(new_n8057_), .ZN(new_n8060_));
  NAND2_X1   g05624(.A1(new_n7641_), .A2(pi0144), .ZN(new_n8061_));
  NAND3_X1   g05625(.A1(new_n7612_), .A2(new_n8058_), .A3(new_n7647_), .ZN(new_n8062_));
  NAND3_X1   g05626(.A1(new_n8061_), .A2(new_n7969_), .A3(new_n8062_), .ZN(new_n8063_));
  AOI21_X1   g05627(.A1(new_n8063_), .A2(new_n8060_), .B(new_n5666_), .ZN(new_n8064_));
  OAI21_X1   g05628(.A1(new_n8064_), .A2(new_n7644_), .B(new_n3265_), .ZN(new_n8065_));
  NOR2_X1    g05629(.A1(pi0038), .A2(pi0155), .ZN(new_n8066_));
  NOR3_X1    g05630(.A1(new_n7628_), .A2(pi0161), .A3(new_n5437_), .ZN(new_n8067_));
  OAI21_X1   g05631(.A1(new_n7632_), .A2(new_n8067_), .B(new_n7508_), .ZN(new_n8068_));
  NAND2_X1   g05632(.A1(new_n8068_), .A2(new_n8066_), .ZN(new_n8069_));
  INV_X1     g05633(.I(new_n7508_), .ZN(new_n8070_));
  NOR2_X1    g05634(.A1(new_n7623_), .A2(new_n3360_), .ZN(new_n8071_));
  NOR3_X1    g05635(.A1(new_n7621_), .A2(new_n8071_), .A3(new_n8070_), .ZN(new_n8072_));
  NAND2_X1   g05636(.A1(new_n3265_), .A2(pi0155), .ZN(new_n8073_));
  OAI21_X1   g05637(.A1(new_n8072_), .A2(new_n8073_), .B(new_n8069_), .ZN(new_n8074_));
  NAND3_X1   g05638(.A1(new_n8074_), .A2(pi0232), .A3(new_n7620_), .ZN(new_n8075_));
  AOI21_X1   g05639(.A1(new_n8065_), .A2(new_n8075_), .B(new_n2627_), .ZN(new_n8076_));
  NOR4_X1    g05640(.A1(new_n8055_), .A2(pi0087), .A3(new_n7980_), .A4(new_n8076_), .ZN(new_n8077_));
  OAI21_X1   g05641(.A1(new_n7967_), .A2(new_n3458_), .B(new_n2702_), .ZN(new_n8078_));
  OAI21_X1   g05642(.A1(new_n8077_), .A2(new_n8078_), .B(new_n7947_), .ZN(new_n8079_));
  AOI21_X1   g05643(.A1(new_n8079_), .A2(new_n2605_), .B(new_n7950_), .ZN(new_n8080_));
  AOI21_X1   g05644(.A1(new_n8080_), .A2(new_n7974_), .B(pi0054), .ZN(new_n8081_));
  OAI21_X1   g05645(.A1(new_n8081_), .A2(new_n7966_), .B(new_n2625_), .ZN(new_n8082_));
  NAND2_X1   g05646(.A1(new_n7924_), .A2(pi0055), .ZN(new_n8083_));
  NAND2_X1   g05647(.A1(new_n7920_), .A2(new_n7348_), .ZN(new_n8084_));
  NOR2_X1    g05648(.A1(new_n7601_), .A2(pi0232), .ZN(new_n8085_));
  NAND2_X1   g05649(.A1(new_n5398_), .A2(pi0162), .ZN(new_n8086_));
  NAND2_X1   g05650(.A1(new_n7600_), .A2(new_n8086_), .ZN(new_n8087_));
  AOI21_X1   g05651(.A1(new_n8087_), .A2(new_n7584_), .B(pi0100), .ZN(new_n8088_));
  NAND2_X1   g05652(.A1(new_n6697_), .A2(pi0167), .ZN(new_n8089_));
  OAI22_X1   g05653(.A1(new_n8088_), .A2(new_n8085_), .B1(new_n3265_), .B2(new_n8089_), .ZN(new_n8090_));
  OAI21_X1   g05654(.A1(new_n8090_), .A2(pi0075), .B(new_n8084_), .ZN(new_n8091_));
  NOR2_X1    g05655(.A1(new_n7585_), .A2(new_n7348_), .ZN(new_n8092_));
  AOI21_X1   g05656(.A1(new_n7926_), .A2(pi0038), .B(pi0054), .ZN(new_n8093_));
  NAND2_X1   g05657(.A1(new_n8093_), .A2(new_n7922_), .ZN(new_n8094_));
  NOR2_X1    g05658(.A1(new_n8094_), .A2(new_n8092_), .ZN(new_n8095_));
  OAI22_X1   g05659(.A1(new_n8091_), .A2(pi0092), .B1(new_n5305_), .B2(new_n8095_), .ZN(new_n8096_));
  NAND2_X1   g05660(.A1(new_n7927_), .A2(pi0054), .ZN(new_n8097_));
  AOI21_X1   g05661(.A1(new_n8096_), .A2(new_n8097_), .B(pi0074), .ZN(new_n8098_));
  OAI21_X1   g05662(.A1(new_n8098_), .A2(new_n8083_), .B(new_n2470_), .ZN(new_n8099_));
  AOI21_X1   g05663(.A1(new_n8082_), .A2(new_n7957_), .B(new_n8099_), .ZN(new_n8100_));
  OAI21_X1   g05664(.A1(pi0074), .A2(new_n8094_), .B(new_n7930_), .ZN(new_n8101_));
  AOI21_X1   g05665(.A1(new_n8101_), .A2(new_n2471_), .B(new_n3425_), .ZN(new_n8102_));
  AOI21_X1   g05666(.A1(new_n7905_), .A2(new_n2471_), .B(new_n3425_), .ZN(new_n8103_));
  NOR2_X1    g05667(.A1(new_n8102_), .A2(new_n8103_), .ZN(new_n8104_));
  OAI21_X1   g05668(.A1(new_n8100_), .A2(new_n8104_), .B(new_n7931_), .ZN(new_n8105_));
  INV_X1     g05669(.I(new_n7957_), .ZN(new_n8106_));
  INV_X1     g05670(.I(new_n7966_), .ZN(new_n8107_));
  INV_X1     g05671(.I(new_n7387_), .ZN(new_n8108_));
  NOR2_X1    g05672(.A1(new_n7948_), .A2(new_n3270_), .ZN(new_n8109_));
  AOI21_X1   g05673(.A1(new_n8109_), .A2(new_n7963_), .B(new_n3458_), .ZN(new_n8110_));
  OR2_X2     g05674(.A1(new_n7960_), .A2(new_n3265_), .Z(new_n8111_));
  NAND3_X1   g05675(.A1(new_n2554_), .A2(new_n2572_), .A3(new_n7970_), .ZN(new_n8112_));
  AOI21_X1   g05676(.A1(new_n8112_), .A2(new_n8111_), .B(new_n6698_), .ZN(new_n8113_));
  OAI21_X1   g05677(.A1(new_n8113_), .A2(pi0100), .B(new_n7947_), .ZN(new_n8114_));
  AOI21_X1   g05678(.A1(new_n8114_), .A2(new_n3458_), .B(new_n8110_), .ZN(new_n8115_));
  OAI21_X1   g05679(.A1(new_n8115_), .A2(new_n8108_), .B(new_n7949_), .ZN(new_n8116_));
  INV_X1     g05680(.I(new_n8110_), .ZN(new_n8117_));
  NAND3_X1   g05681(.A1(new_n7453_), .A2(pi0159), .A3(new_n7985_), .ZN(new_n8118_));
  NAND3_X1   g05682(.A1(new_n8118_), .A2(pi0299), .A3(new_n8086_), .ZN(new_n8119_));
  NAND2_X1   g05683(.A1(new_n7442_), .A2(new_n3107_), .ZN(new_n8120_));
  AOI21_X1   g05684(.A1(new_n8120_), .A2(new_n7436_), .B(pi0161), .ZN(new_n8121_));
  INV_X1     g05685(.I(new_n7448_), .ZN(new_n8122_));
  INV_X1     g05686(.I(new_n7449_), .ZN(new_n8123_));
  NOR2_X1    g05687(.A1(new_n8123_), .A2(pi0146), .ZN(new_n8124_));
  OAI21_X1   g05688(.A1(new_n8124_), .A2(new_n8122_), .B(pi0161), .ZN(new_n8125_));
  AOI21_X1   g05689(.A1(new_n3185_), .A2(pi0159), .B(new_n2628_), .ZN(new_n8126_));
  NAND2_X1   g05690(.A1(new_n8125_), .A2(new_n8126_), .ZN(new_n8127_));
  OAI21_X1   g05691(.A1(new_n8121_), .A2(new_n8127_), .B(new_n8119_), .ZN(new_n8128_));
  NAND2_X1   g05692(.A1(new_n7474_), .A2(pi0146), .ZN(new_n8129_));
  NAND2_X1   g05693(.A1(new_n7467_), .A2(new_n3107_), .ZN(new_n8130_));
  AOI21_X1   g05694(.A1(new_n8130_), .A2(new_n8129_), .B(pi0161), .ZN(new_n8131_));
  NOR3_X1    g05695(.A1(new_n7461_), .A2(pi0146), .A3(new_n3360_), .ZN(new_n8132_));
  OAI21_X1   g05696(.A1(new_n8131_), .A2(new_n8132_), .B(new_n7985_), .ZN(new_n8133_));
  NAND2_X1   g05697(.A1(new_n8128_), .A2(new_n8133_), .ZN(new_n8134_));
  NOR2_X1    g05698(.A1(new_n8123_), .A2(pi0142), .ZN(new_n8135_));
  NOR3_X1    g05699(.A1(new_n8135_), .A2(new_n7934_), .A3(new_n7482_), .ZN(new_n8136_));
  AOI21_X1   g05700(.A1(new_n7462_), .A2(new_n2724_), .B(pi0140), .ZN(new_n8137_));
  NOR2_X1    g05701(.A1(new_n8136_), .A2(new_n8137_), .ZN(new_n8138_));
  OAI22_X1   g05702(.A1(new_n8138_), .A2(new_n8058_), .B1(new_n7934_), .B2(new_n5398_), .ZN(new_n8139_));
  NAND2_X1   g05703(.A1(new_n7442_), .A2(new_n2724_), .ZN(new_n8140_));
  NAND3_X1   g05704(.A1(new_n8140_), .A2(pi0140), .A3(new_n7481_), .ZN(new_n8141_));
  NOR2_X1    g05705(.A1(new_n7467_), .A2(pi0142), .ZN(new_n8142_));
  NOR2_X1    g05706(.A1(new_n7474_), .A2(new_n2724_), .ZN(new_n8143_));
  OAI21_X1   g05707(.A1(new_n8142_), .A2(new_n8143_), .B(new_n7934_), .ZN(new_n8144_));
  AOI21_X1   g05708(.A1(new_n8141_), .A2(new_n8144_), .B(pi0144), .ZN(new_n8145_));
  AOI21_X1   g05709(.A1(new_n7453_), .A2(pi0181), .B(pi0299), .ZN(new_n8146_));
  OAI21_X1   g05710(.A1(new_n8145_), .A2(new_n8139_), .B(new_n8146_), .ZN(new_n8147_));
  NAND3_X1   g05711(.A1(new_n8147_), .A2(new_n8134_), .A3(pi0232), .ZN(new_n8148_));
  AOI21_X1   g05712(.A1(new_n8148_), .A2(new_n2572_), .B(new_n7980_), .ZN(new_n8149_));
  NOR2_X1    g05713(.A1(new_n2627_), .A2(pi0038), .ZN(new_n8150_));
  NOR2_X1    g05714(.A1(new_n7526_), .A2(new_n8058_), .ZN(new_n8151_));
  NOR2_X1    g05715(.A1(new_n7527_), .A2(pi0144), .ZN(new_n8152_));
  OAI21_X1   g05716(.A1(new_n8151_), .A2(new_n8152_), .B(new_n8057_), .ZN(new_n8153_));
  OAI21_X1   g05717(.A1(new_n7522_), .A2(pi0144), .B(new_n7969_), .ZN(new_n8154_));
  NAND3_X1   g05718(.A1(new_n8153_), .A2(pi0232), .A3(new_n8154_), .ZN(new_n8155_));
  NOR4_X1    g05719(.A1(new_n5551_), .A2(pi0161), .A3(new_n5437_), .A4(new_n5422_), .ZN(new_n8156_));
  AOI21_X1   g05720(.A1(new_n7514_), .A2(pi0161), .B(new_n8156_), .ZN(new_n8157_));
  OAI21_X1   g05721(.A1(new_n8157_), .A2(new_n8070_), .B(pi0155), .ZN(new_n8158_));
  INV_X1     g05722(.I(new_n7511_), .ZN(new_n8159_));
  NAND2_X1   g05723(.A1(new_n7508_), .A2(new_n3360_), .ZN(new_n8160_));
  OAI21_X1   g05724(.A1(new_n8159_), .A2(new_n8160_), .B(new_n7968_), .ZN(new_n8161_));
  AOI21_X1   g05725(.A1(new_n8158_), .A2(new_n8161_), .B(new_n2628_), .ZN(new_n8162_));
  OAI21_X1   g05726(.A1(new_n8162_), .A2(new_n8155_), .B(new_n8150_), .ZN(new_n8163_));
  NAND2_X1   g05727(.A1(new_n8149_), .A2(new_n8163_), .ZN(new_n8164_));
  AOI21_X1   g05728(.A1(new_n8164_), .A2(new_n2702_), .B(new_n7948_), .ZN(new_n8165_));
  OAI21_X1   g05729(.A1(new_n8165_), .A2(pi0087), .B(new_n8117_), .ZN(new_n8166_));
  AOI21_X1   g05730(.A1(new_n8166_), .A2(new_n2605_), .B(new_n8116_), .ZN(new_n8167_));
  OAI21_X1   g05731(.A1(new_n8167_), .A2(pi0054), .B(new_n8107_), .ZN(new_n8168_));
  AOI21_X1   g05732(.A1(new_n8168_), .A2(new_n2625_), .B(new_n8106_), .ZN(new_n8169_));
  NOR2_X1    g05733(.A1(pi0038), .A2(pi0087), .ZN(new_n8170_));
  NAND4_X1   g05734(.A1(new_n7504_), .A2(new_n3444_), .A3(pi0162), .A4(new_n8170_), .ZN(new_n8171_));
  OAI22_X1   g05735(.A1(new_n5505_), .A2(new_n8171_), .B1(new_n3265_), .B2(new_n8089_), .ZN(new_n8172_));
  NAND2_X1   g05736(.A1(new_n8172_), .A2(new_n7342_), .ZN(new_n8173_));
  NOR2_X1    g05737(.A1(new_n7926_), .A2(new_n5499_), .ZN(new_n8174_));
  AOI21_X1   g05738(.A1(new_n8173_), .A2(new_n5499_), .B(new_n8174_), .ZN(new_n8175_));
  NOR3_X1    g05739(.A1(new_n8175_), .A2(pi0074), .A3(new_n7921_), .ZN(new_n8176_));
  OAI21_X1   g05740(.A1(new_n8176_), .A2(new_n8083_), .B(new_n2470_), .ZN(new_n8177_));
  OAI21_X1   g05741(.A1(new_n8169_), .A2(new_n8177_), .B(new_n8102_), .ZN(new_n8178_));
  AND2_X2    g05742(.A1(new_n8178_), .A2(new_n7931_), .Z(new_n8179_));
  NOR2_X1    g05743(.A1(new_n8179_), .A2(new_n7559_), .ZN(new_n8180_));
  AOI21_X1   g05744(.A1(new_n8105_), .A2(new_n7559_), .B(new_n8180_), .ZN(new_n8181_));
  NOR2_X1    g05745(.A1(new_n8181_), .A2(new_n7915_), .ZN(new_n8182_));
  NAND2_X1   g05746(.A1(new_n7563_), .A2(new_n7560_), .ZN(new_n8183_));
  NAND2_X1   g05747(.A1(new_n8183_), .A2(new_n7559_), .ZN(new_n8184_));
  NAND2_X1   g05748(.A1(new_n8105_), .A2(new_n8184_), .ZN(new_n8185_));
  OAI21_X1   g05749(.A1(new_n8179_), .A2(new_n8184_), .B(new_n8185_), .ZN(new_n8186_));
  AOI21_X1   g05750(.A1(new_n8186_), .A2(new_n7915_), .B(new_n8182_), .ZN(po0192));
  NOR3_X1    g05751(.A1(new_n7335_), .A2(new_n2471_), .A3(new_n2612_), .ZN(new_n8188_));
  INV_X1     g05752(.I(new_n8188_), .ZN(new_n8189_));
  NOR2_X1    g05753(.A1(new_n8189_), .A2(pi0055), .ZN(new_n8190_));
  NAND2_X1   g05754(.A1(new_n8190_), .A2(pi0059), .ZN(new_n8191_));
  AOI21_X1   g05755(.A1(new_n5360_), .A2(new_n2985_), .B(pi0093), .ZN(new_n8192_));
  OAI21_X1   g05756(.A1(new_n5376_), .A2(new_n8192_), .B(new_n2743_), .ZN(new_n8193_));
  AOI21_X1   g05757(.A1(new_n3009_), .A2(pi0035), .B(new_n7291_), .ZN(new_n8194_));
  AND2_X2    g05758(.A1(new_n8193_), .A2(new_n8194_), .Z(new_n8195_));
  OAI21_X1   g05759(.A1(new_n8195_), .A2(new_n2819_), .B(pi1082), .ZN(new_n8196_));
  NOR2_X1    g05760(.A1(new_n8196_), .A2(new_n7456_), .ZN(new_n8197_));
  NOR2_X1    g05761(.A1(new_n5351_), .A2(pi0137), .ZN(new_n8198_));
  NOR4_X1    g05762(.A1(new_n8198_), .A2(pi0122), .A3(po0740), .A4(new_n6350_), .ZN(new_n8199_));
  INV_X1     g05763(.I(new_n6703_), .ZN(new_n8200_));
  NOR4_X1    g05764(.A1(new_n8200_), .A2(new_n8198_), .A3(new_n3026_), .A4(new_n6349_), .ZN(new_n8201_));
  INV_X1     g05765(.I(new_n8193_), .ZN(new_n8202_));
  NOR2_X1    g05766(.A1(new_n8202_), .A2(new_n5350_), .ZN(new_n8203_));
  NOR3_X1    g05767(.A1(new_n8203_), .A2(new_n8199_), .A3(new_n8201_), .ZN(new_n8204_));
  NAND2_X1   g05768(.A1(new_n7309_), .A2(new_n2740_), .ZN(new_n8205_));
  NAND2_X1   g05769(.A1(new_n8202_), .A2(new_n8205_), .ZN(new_n8206_));
  NAND3_X1   g05770(.A1(new_n8206_), .A2(new_n2525_), .A3(new_n8194_), .ZN(new_n8207_));
  NOR2_X1    g05771(.A1(new_n8204_), .A2(new_n8207_), .ZN(new_n8208_));
  NAND4_X1   g05772(.A1(new_n6662_), .A2(pi0032), .A3(new_n2771_), .A4(new_n7280_), .ZN(new_n8209_));
  NAND2_X1   g05773(.A1(new_n8195_), .A2(new_n2725_), .ZN(new_n8210_));
  NAND2_X1   g05774(.A1(new_n5350_), .A2(new_n2462_), .ZN(new_n8211_));
  AOI21_X1   g05775(.A1(new_n8210_), .A2(new_n8209_), .B(new_n8211_), .ZN(new_n8212_));
  NOR4_X1    g05776(.A1(new_n8208_), .A2(new_n8197_), .A3(new_n8212_), .A4(pi0038), .ZN(new_n8213_));
  NAND2_X1   g05777(.A1(new_n7335_), .A2(pi0038), .ZN(new_n8214_));
  NAND3_X1   g05778(.A1(new_n8214_), .A2(new_n2627_), .A3(new_n2702_), .ZN(new_n8215_));
  INV_X1     g05779(.I(new_n7323_), .ZN(new_n8216_));
  INV_X1     g05780(.I(new_n7324_), .ZN(new_n8217_));
  NOR2_X1    g05781(.A1(new_n3081_), .A2(new_n5532_), .ZN(new_n8218_));
  NOR2_X1    g05782(.A1(new_n8218_), .A2(new_n6259_), .ZN(new_n8219_));
  INV_X1     g05783(.I(new_n8219_), .ZN(new_n8220_));
  NOR2_X1    g05784(.A1(new_n8220_), .A2(new_n5325_), .ZN(new_n8221_));
  NOR3_X1    g05785(.A1(new_n5323_), .A2(new_n2704_), .A3(new_n8221_), .ZN(new_n8222_));
  NOR2_X1    g05786(.A1(new_n8217_), .A2(new_n8222_), .ZN(new_n8223_));
  INV_X1     g05787(.I(new_n6699_), .ZN(new_n8224_));
  AOI22_X1   g05788(.A1(new_n6693_), .A2(pi0146), .B1(pi0142), .B2(new_n6694_), .ZN(new_n8225_));
  AOI22_X1   g05789(.A1(new_n8222_), .A2(new_n8224_), .B1(new_n6696_), .B2(new_n8225_), .ZN(new_n8226_));
  NAND2_X1   g05790(.A1(new_n3016_), .A2(pi0252), .ZN(new_n8227_));
  AOI22_X1   g05791(.A1(new_n8223_), .A2(new_n5309_), .B1(new_n8226_), .B2(new_n8227_), .ZN(new_n8228_));
  NOR2_X1    g05792(.A1(new_n8228_), .A2(new_n8216_), .ZN(new_n8229_));
  AOI21_X1   g05793(.A1(pi0137), .A2(new_n7320_), .B(new_n8229_), .ZN(new_n8230_));
  OAI22_X1   g05794(.A1(new_n8213_), .A2(new_n8215_), .B1(new_n7328_), .B2(new_n8230_), .ZN(new_n8231_));
  NOR3_X1    g05795(.A1(new_n5324_), .A2(new_n3016_), .A3(po0840), .ZN(new_n8232_));
  OR2_X2     g05796(.A1(new_n8232_), .A2(new_n7325_), .Z(new_n8233_));
  AOI22_X1   g05797(.A1(new_n8231_), .A2(new_n2564_), .B1(new_n7338_), .B2(new_n8233_), .ZN(new_n8234_));
  OAI21_X1   g05798(.A1(new_n8234_), .A2(pi0092), .B(new_n5499_), .ZN(new_n8235_));
  NAND2_X1   g05799(.A1(new_n6174_), .A2(new_n7278_), .ZN(new_n8236_));
  NAND2_X1   g05800(.A1(new_n8236_), .A2(pi0054), .ZN(new_n8237_));
  NOR2_X1    g05801(.A1(new_n5476_), .A2(pi0074), .ZN(new_n8238_));
  NAND4_X1   g05802(.A1(new_n8235_), .A2(new_n2469_), .A3(new_n8237_), .A4(new_n8238_), .ZN(new_n8239_));
  AOI21_X1   g05803(.A1(new_n8239_), .A2(new_n8191_), .B(pi0057), .ZN(po0193));
  INV_X1     g05804(.I(po0740), .ZN(new_n8241_));
  INV_X1     g05805(.I(new_n7297_), .ZN(new_n8242_));
  NOR2_X1    g05806(.A1(new_n8242_), .A2(pi0102), .ZN(new_n8243_));
  INV_X1     g05807(.I(new_n8243_), .ZN(new_n8244_));
  NOR4_X1    g05808(.A1(new_n8244_), .A2(new_n7409_), .A3(new_n2850_), .A4(pi0065), .ZN(new_n8245_));
  INV_X1     g05809(.I(new_n8245_), .ZN(new_n8246_));
  NOR2_X1    g05810(.A1(new_n8246_), .A2(pi0069), .ZN(new_n8247_));
  NOR2_X1    g05811(.A1(pi0067), .A2(pi0103), .ZN(new_n8248_));
  NAND4_X1   g05812(.A1(new_n8247_), .A2(pi0036), .A3(new_n2962_), .A4(new_n8248_), .ZN(new_n8249_));
  NOR3_X1    g05813(.A1(new_n8249_), .A2(pi0083), .A3(new_n2919_), .ZN(new_n8250_));
  NOR2_X1    g05814(.A1(new_n2787_), .A2(new_n2858_), .ZN(new_n8251_));
  AOI22_X1   g05815(.A1(new_n6719_), .A2(new_n5359_), .B1(new_n8250_), .B2(new_n8251_), .ZN(new_n8252_));
  NOR3_X1    g05816(.A1(new_n5354_), .A2(new_n2536_), .A3(new_n2741_), .ZN(new_n8253_));
  INV_X1     g05817(.I(new_n8253_), .ZN(new_n8254_));
  NOR2_X1    g05818(.A1(po1038), .A2(new_n2563_), .ZN(new_n8255_));
  INV_X1     g05819(.I(new_n8255_), .ZN(new_n8256_));
  NOR2_X1    g05820(.A1(new_n8256_), .A2(new_n3436_), .ZN(new_n8257_));
  INV_X1     g05821(.I(new_n8257_), .ZN(new_n8258_));
  NOR2_X1    g05822(.A1(new_n8258_), .A2(pi0092), .ZN(new_n8259_));
  INV_X1     g05823(.I(new_n8259_), .ZN(new_n8260_));
  NOR2_X1    g05824(.A1(new_n8260_), .A2(new_n8254_), .ZN(new_n8261_));
  INV_X1     g05825(.I(new_n8261_), .ZN(new_n8262_));
  NOR3_X1    g05826(.A1(new_n8252_), .A2(new_n8241_), .A3(new_n8262_), .ZN(po0194));
  NOR2_X1    g05827(.A1(new_n2610_), .A2(po1038), .ZN(new_n8264_));
  INV_X1     g05828(.I(new_n8264_), .ZN(new_n8265_));
  NOR4_X1    g05829(.A1(new_n2751_), .A2(new_n7278_), .A3(pi0039), .A4(new_n2526_), .ZN(new_n8266_));
  NAND2_X1   g05830(.A1(new_n8266_), .A2(pi0038), .ZN(new_n8267_));
  NOR4_X1    g05831(.A1(new_n2546_), .A2(new_n2522_), .A3(new_n2536_), .A4(new_n2551_), .ZN(new_n8268_));
  AND4_X2    g05832(.A1(new_n2627_), .A2(new_n8268_), .A3(new_n3179_), .A4(new_n7414_), .Z(new_n8269_));
  INV_X1     g05833(.I(new_n7419_), .ZN(new_n8270_));
  NAND3_X1   g05834(.A1(new_n2911_), .A2(new_n2915_), .A3(pi0089), .ZN(new_n8271_));
  NAND4_X1   g05835(.A1(new_n2933_), .A2(new_n2478_), .A3(new_n2929_), .A4(new_n2927_), .ZN(new_n8272_));
  NOR4_X1    g05836(.A1(new_n8272_), .A2(pi0048), .A3(pi0065), .A4(new_n8271_), .ZN(new_n8273_));
  NOR4_X1    g05837(.A1(new_n2484_), .A2(pi0071), .A3(new_n7409_), .A4(pi0104), .ZN(new_n8274_));
  NAND3_X1   g05838(.A1(new_n8270_), .A2(new_n8273_), .A3(new_n8274_), .ZN(new_n8275_));
  OAI21_X1   g05839(.A1(new_n8275_), .A2(new_n2630_), .B(new_n2495_), .ZN(new_n8276_));
  NOR2_X1    g05840(.A1(new_n2892_), .A2(pi0081), .ZN(new_n8277_));
  NAND4_X1   g05841(.A1(new_n8277_), .A2(new_n8269_), .A3(new_n3265_), .A4(new_n8276_), .ZN(new_n8278_));
  AOI21_X1   g05842(.A1(new_n8267_), .A2(new_n8278_), .B(new_n8265_), .ZN(po0196));
  NOR2_X1    g05843(.A1(new_n8265_), .A2(pi0038), .ZN(new_n8280_));
  INV_X1     g05844(.I(new_n8280_), .ZN(new_n8281_));
  INV_X1     g05845(.I(pi0287), .ZN(new_n8282_));
  NAND4_X1   g05846(.A1(new_n2547_), .A2(new_n8282_), .A3(new_n2523_), .A4(new_n2529_), .ZN(new_n8283_));
  AOI21_X1   g05847(.A1(new_n3082_), .A2(new_n5387_), .B(new_n5386_), .ZN(new_n8284_));
  OR2_X2     g05848(.A1(new_n8284_), .A2(new_n5390_), .Z(new_n8285_));
  NAND2_X1   g05849(.A1(new_n5430_), .A2(new_n8285_), .ZN(new_n8286_));
  OAI21_X1   g05850(.A1(new_n6745_), .A2(new_n8286_), .B(new_n5391_), .ZN(new_n8287_));
  NOR2_X1    g05851(.A1(new_n8287_), .A2(new_n8283_), .ZN(new_n8288_));
  NOR2_X1    g05852(.A1(new_n8288_), .A2(new_n5445_), .ZN(new_n8289_));
  OAI21_X1   g05853(.A1(new_n5413_), .A2(new_n8286_), .B(new_n5391_), .ZN(new_n8290_));
  NOR2_X1    g05854(.A1(new_n8290_), .A2(new_n8283_), .ZN(new_n8291_));
  NOR2_X1    g05855(.A1(new_n8291_), .A2(new_n5446_), .ZN(new_n8292_));
  OAI21_X1   g05856(.A1(new_n8289_), .A2(new_n8292_), .B(new_n2628_), .ZN(new_n8293_));
  NOR2_X1    g05857(.A1(new_n8286_), .A2(new_n3041_), .ZN(new_n8294_));
  NOR4_X1    g05858(.A1(new_n8283_), .A2(pi0223), .A3(new_n5392_), .A4(new_n8294_), .ZN(new_n8295_));
  NOR2_X1    g05859(.A1(new_n8293_), .A2(new_n8295_), .ZN(new_n8296_));
  INV_X1     g05860(.I(pi0786), .ZN(new_n8297_));
  NOR2_X1    g05861(.A1(new_n8288_), .A2(new_n6764_), .ZN(new_n8298_));
  NOR2_X1    g05862(.A1(new_n8291_), .A2(new_n5422_), .ZN(new_n8299_));
  OAI21_X1   g05863(.A1(new_n8298_), .A2(new_n8299_), .B(pi0299), .ZN(new_n8300_));
  NOR4_X1    g05864(.A1(new_n8283_), .A2(pi0215), .A3(new_n5392_), .A4(new_n8294_), .ZN(new_n8301_));
  OAI22_X1   g05865(.A1(new_n8300_), .A2(new_n8301_), .B1(new_n8297_), .B2(pi1082), .ZN(new_n8302_));
  NOR2_X1    g05866(.A1(new_n8297_), .A2(pi1082), .ZN(new_n8303_));
  INV_X1     g05867(.I(new_n5113_), .ZN(new_n8304_));
  OAI22_X1   g05868(.A1(new_n6809_), .A2(new_n8304_), .B1(new_n3336_), .B2(new_n5451_), .ZN(new_n8305_));
  NAND4_X1   g05869(.A1(new_n8305_), .A2(po0740), .A3(new_n5526_), .A4(new_n8303_), .ZN(new_n8306_));
  OAI21_X1   g05870(.A1(new_n8302_), .A2(new_n8296_), .B(new_n8306_), .ZN(new_n8307_));
  NAND2_X1   g05871(.A1(new_n8307_), .A2(pi0039), .ZN(new_n8308_));
  OAI21_X1   g05872(.A1(new_n2772_), .A2(pi0841), .B(pi0035), .ZN(new_n8309_));
  NAND3_X1   g05873(.A1(new_n8309_), .A2(new_n2533_), .A3(new_n7569_), .ZN(new_n8310_));
  OAI21_X1   g05874(.A1(po0740), .A2(pi0986), .B(pi0252), .ZN(new_n8311_));
  INV_X1     g05875(.I(new_n8311_), .ZN(new_n8312_));
  NOR2_X1    g05876(.A1(new_n2727_), .A2(new_n2844_), .ZN(new_n8313_));
  NAND4_X1   g05877(.A1(new_n2478_), .A2(new_n2922_), .A3(new_n2911_), .A4(pi0048), .ZN(new_n8314_));
  NOR2_X1    g05878(.A1(pi0066), .A2(pi0084), .ZN(new_n8315_));
  NAND2_X1   g05879(.A1(new_n7297_), .A2(new_n8315_), .ZN(new_n8316_));
  NOR3_X1    g05880(.A1(new_n8316_), .A2(pi0065), .A3(pi0069), .ZN(new_n8317_));
  INV_X1     g05881(.I(new_n8317_), .ZN(new_n8318_));
  NOR4_X1    g05882(.A1(new_n8318_), .A2(pi0045), .A3(new_n8314_), .A4(pi0073), .ZN(new_n8319_));
  INV_X1     g05883(.I(new_n7296_), .ZN(new_n8320_));
  NOR3_X1    g05884(.A1(new_n7304_), .A2(new_n6668_), .A3(new_n8320_), .ZN(new_n8321_));
  NAND4_X1   g05885(.A1(new_n8319_), .A2(new_n7418_), .A3(new_n8274_), .A4(new_n8321_), .ZN(new_n8322_));
  NOR3_X1    g05886(.A1(new_n8322_), .A2(pi0047), .A3(pi0841), .ZN(new_n8323_));
  OAI22_X1   g05887(.A1(new_n8323_), .A2(new_n8313_), .B1(new_n5590_), .B2(new_n8312_), .ZN(new_n8324_));
  NOR3_X1    g05888(.A1(new_n8324_), .A2(new_n2756_), .A3(new_n2733_), .ZN(new_n8325_));
  NAND4_X1   g05889(.A1(new_n5363_), .A2(pi0314), .A3(new_n2732_), .A4(new_n8311_), .ZN(new_n8326_));
  OAI21_X1   g05890(.A1(new_n2861_), .A2(new_n2849_), .B(new_n2784_), .ZN(new_n8327_));
  NAND3_X1   g05891(.A1(new_n2515_), .A2(new_n2514_), .A3(new_n3179_), .ZN(new_n8328_));
  OR4_X2     g05892(.A1(pi0097), .A2(new_n8327_), .A3(new_n8322_), .A4(new_n8328_), .Z(new_n8329_));
  NOR2_X1    g05893(.A1(new_n2783_), .A2(new_n2849_), .ZN(new_n8330_));
  AOI21_X1   g05894(.A1(new_n2861_), .A2(new_n8330_), .B(pi0047), .ZN(new_n8331_));
  AOI21_X1   g05895(.A1(new_n8329_), .A2(new_n8331_), .B(new_n8326_), .ZN(new_n8332_));
  OAI21_X1   g05896(.A1(new_n8332_), .A2(new_n8325_), .B(new_n2740_), .ZN(new_n8333_));
  AOI21_X1   g05897(.A1(new_n8333_), .A2(new_n2743_), .B(new_n8310_), .ZN(new_n8334_));
  NOR2_X1    g05898(.A1(new_n5614_), .A2(new_n5350_), .ZN(new_n8335_));
  NOR2_X1    g05899(.A1(pi0039), .A2(pi0095), .ZN(new_n8336_));
  OAI21_X1   g05900(.A1(new_n8334_), .A2(new_n8335_), .B(new_n8336_), .ZN(new_n8337_));
  AOI21_X1   g05901(.A1(new_n8337_), .A2(new_n8308_), .B(new_n8281_), .ZN(po0197));
  NAND3_X1   g05902(.A1(new_n2505_), .A2(new_n2763_), .A3(pi0102), .ZN(new_n8339_));
  NOR4_X1    g05903(.A1(new_n2970_), .A2(new_n2546_), .A3(new_n5354_), .A4(new_n8339_), .ZN(new_n8340_));
  NAND3_X1   g05904(.A1(new_n8340_), .A2(pi1082), .A3(new_n2535_), .ZN(new_n8341_));
  OAI21_X1   g05905(.A1(new_n2552_), .A2(new_n2818_), .B(new_n2525_), .ZN(new_n8342_));
  NOR2_X1    g05906(.A1(new_n8340_), .A2(pi0040), .ZN(new_n8343_));
  OR3_X2     g05907(.A1(new_n8342_), .A2(pi1082), .A3(new_n8343_), .Z(new_n8344_));
  AOI21_X1   g05908(.A1(new_n8344_), .A2(new_n8341_), .B(new_n8260_), .ZN(po0198));
  INV_X1     g05909(.I(pi0041), .ZN(new_n8346_));
  NOR2_X1    g05910(.A1(new_n8346_), .A2(pi0039), .ZN(new_n8347_));
  NOR2_X1    g05911(.A1(new_n5437_), .A2(pi0166), .ZN(new_n8348_));
  INV_X1     g05912(.I(new_n8348_), .ZN(new_n8349_));
  NOR3_X1    g05913(.A1(new_n8349_), .A2(pi0152), .A3(new_n3360_), .ZN(new_n8350_));
  INV_X1     g05914(.I(new_n8350_), .ZN(new_n8351_));
  NOR2_X1    g05915(.A1(new_n8351_), .A2(new_n7507_), .ZN(new_n8352_));
  NOR4_X1    g05916(.A1(new_n8352_), .A2(pi0072), .A3(new_n6643_), .A4(new_n8347_), .ZN(new_n8353_));
  NOR2_X1    g05917(.A1(new_n5437_), .A2(pi0189), .ZN(new_n8354_));
  INV_X1     g05918(.I(new_n8354_), .ZN(new_n8355_));
  NOR2_X1    g05919(.A1(new_n8355_), .A2(new_n8058_), .ZN(new_n8356_));
  AOI21_X1   g05920(.A1(new_n8356_), .A2(new_n7488_), .B(pi0299), .ZN(new_n8357_));
  INV_X1     g05921(.I(new_n8357_), .ZN(new_n8358_));
  AOI21_X1   g05922(.A1(new_n8351_), .A2(new_n6978_), .B(new_n5666_), .ZN(new_n8359_));
  AND2_X2    g05923(.A1(new_n8359_), .A2(new_n8358_), .Z(new_n8360_));
  INV_X1     g05924(.I(new_n8360_), .ZN(new_n8361_));
  AOI21_X1   g05925(.A1(new_n8361_), .A2(new_n2821_), .B(new_n2627_), .ZN(new_n8362_));
  NOR2_X1    g05926(.A1(pi0041), .A2(pi0072), .ZN(new_n8363_));
  NOR2_X1    g05927(.A1(new_n8363_), .A2(pi0039), .ZN(new_n8364_));
  NOR2_X1    g05928(.A1(new_n8362_), .A2(new_n8364_), .ZN(new_n8365_));
  INV_X1     g05929(.I(new_n8365_), .ZN(new_n8366_));
  AOI21_X1   g05930(.A1(new_n8366_), .A2(new_n6648_), .B(po1038), .ZN(new_n8367_));
  INV_X1     g05931(.I(new_n8362_), .ZN(new_n8368_));
  NOR2_X1    g05932(.A1(new_n6819_), .A2(new_n3026_), .ZN(new_n8369_));
  INV_X1     g05933(.I(new_n8369_), .ZN(new_n8370_));
  NOR2_X1    g05934(.A1(new_n2821_), .A2(pi0041), .ZN(new_n8371_));
  NOR2_X1    g05935(.A1(new_n5320_), .A2(pi0099), .ZN(new_n8372_));
  INV_X1     g05936(.I(pi0101), .ZN(new_n8373_));
  NOR2_X1    g05937(.A1(new_n8373_), .A2(pi0072), .ZN(new_n8374_));
  NOR2_X1    g05938(.A1(new_n8374_), .A2(pi0041), .ZN(new_n8375_));
  INV_X1     g05939(.I(new_n8375_), .ZN(new_n8376_));
  INV_X1     g05940(.I(pi0044), .ZN(new_n8377_));
  NOR2_X1    g05941(.A1(new_n2751_), .A2(new_n2536_), .ZN(new_n8378_));
  INV_X1     g05942(.I(new_n8378_), .ZN(new_n8379_));
  NOR2_X1    g05943(.A1(new_n8379_), .A2(new_n8200_), .ZN(new_n8380_));
  INV_X1     g05944(.I(new_n8380_), .ZN(new_n8381_));
  NOR3_X1    g05945(.A1(new_n8381_), .A2(pi0024), .A3(new_n2704_), .ZN(new_n8382_));
  NAND2_X1   g05946(.A1(new_n8382_), .A2(new_n8377_), .ZN(new_n8383_));
  NOR3_X1    g05947(.A1(new_n8383_), .A2(new_n8372_), .A3(new_n8376_), .ZN(new_n8384_));
  NOR2_X1    g05948(.A1(new_n2530_), .A2(pi0044), .ZN(new_n8385_));
  INV_X1     g05949(.I(new_n8385_), .ZN(new_n8386_));
  NOR2_X1    g05950(.A1(new_n8386_), .A2(pi0101), .ZN(new_n8387_));
  INV_X1     g05951(.I(new_n8387_), .ZN(new_n8388_));
  NOR2_X1    g05952(.A1(new_n8388_), .A2(new_n8200_), .ZN(new_n8389_));
  INV_X1     g05953(.I(new_n8389_), .ZN(new_n8390_));
  NOR2_X1    g05954(.A1(new_n8390_), .A2(new_n6707_), .ZN(new_n8391_));
  NOR2_X1    g05955(.A1(new_n8391_), .A2(new_n8346_), .ZN(new_n8392_));
  NOR4_X1    g05956(.A1(new_n8384_), .A2(new_n3026_), .A3(new_n8371_), .A4(new_n8392_), .ZN(new_n8393_));
  AOI22_X1   g05957(.A1(new_n8393_), .A2(new_n6774_), .B1(new_n8363_), .B2(new_n8370_), .ZN(new_n8394_));
  AOI21_X1   g05958(.A1(new_n8394_), .A2(new_n2627_), .B(new_n5792_), .ZN(new_n8395_));
  OAI21_X1   g05959(.A1(new_n8366_), .A2(new_n2626_), .B(pi0075), .ZN(new_n8396_));
  AOI21_X1   g05960(.A1(new_n8395_), .A2(new_n8368_), .B(new_n8396_), .ZN(new_n8397_));
  AOI21_X1   g05961(.A1(new_n2458_), .A2(new_n8363_), .B(new_n3273_), .ZN(new_n8398_));
  NOR2_X1    g05962(.A1(new_n8387_), .A2(new_n8346_), .ZN(new_n8399_));
  NOR3_X1    g05963(.A1(new_n8379_), .A2(pi0044), .A3(new_n8376_), .ZN(new_n8400_));
  NOR2_X1    g05964(.A1(new_n8400_), .A2(new_n8371_), .ZN(new_n8401_));
  NAND2_X1   g05965(.A1(new_n8401_), .A2(pi0228), .ZN(new_n8402_));
  OAI21_X1   g05966(.A1(new_n8402_), .A2(new_n8399_), .B(new_n8398_), .ZN(new_n8403_));
  NAND2_X1   g05967(.A1(new_n8364_), .A2(new_n3271_), .ZN(new_n8404_));
  NAND4_X1   g05968(.A1(new_n8403_), .A2(pi0087), .A3(new_n8368_), .A4(new_n8404_), .ZN(new_n8405_));
  NAND2_X1   g05969(.A1(new_n8405_), .A2(new_n3465_), .ZN(new_n8406_));
  NOR2_X1    g05970(.A1(new_n2530_), .A2(new_n8282_), .ZN(new_n8407_));
  NAND2_X1   g05971(.A1(new_n8360_), .A2(new_n8407_), .ZN(new_n8408_));
  OAI21_X1   g05972(.A1(pi0072), .A2(new_n8360_), .B(new_n8408_), .ZN(new_n8409_));
  AOI21_X1   g05973(.A1(new_n8409_), .A2(pi0039), .B(new_n3271_), .ZN(new_n8410_));
  INV_X1     g05974(.I(pi0949), .ZN(new_n8411_));
  NAND2_X1   g05975(.A1(new_n2842_), .A2(new_n7272_), .ZN(new_n8412_));
  NOR2_X1    g05976(.A1(new_n8412_), .A2(new_n2509_), .ZN(new_n8413_));
  INV_X1     g05977(.I(new_n8413_), .ZN(new_n8414_));
  NOR4_X1    g05978(.A1(new_n8414_), .A2(pi0480), .A3(new_n8411_), .A4(new_n2749_), .ZN(new_n8415_));
  INV_X1     g05979(.I(pi0901), .ZN(new_n8416_));
  NOR2_X1    g05980(.A1(new_n8416_), .A2(pi0959), .ZN(new_n8417_));
  NOR2_X1    g05981(.A1(new_n8415_), .A2(new_n8417_), .ZN(new_n8418_));
  NOR2_X1    g05982(.A1(new_n2704_), .A2(pi0250), .ZN(new_n8419_));
  INV_X1     g05983(.I(new_n8419_), .ZN(new_n8420_));
  NOR3_X1    g05984(.A1(new_n8418_), .A2(new_n2536_), .A3(new_n8420_), .ZN(new_n8421_));
  NOR4_X1    g05985(.A1(new_n2749_), .A2(pi0047), .A3(pi0480), .A4(new_n8411_), .ZN(new_n8422_));
  NAND2_X1   g05986(.A1(new_n2512_), .A2(new_n2782_), .ZN(new_n8423_));
  INV_X1     g05987(.I(new_n8423_), .ZN(new_n8424_));
  AOI21_X1   g05988(.A1(new_n2875_), .A2(new_n8424_), .B(pi0110), .ZN(new_n8425_));
  NOR3_X1    g05989(.A1(new_n8425_), .A2(new_n2733_), .A3(new_n2843_), .ZN(new_n8426_));
  INV_X1     g05990(.I(pi0480), .ZN(new_n8427_));
  NAND2_X1   g05991(.A1(new_n8427_), .A2(pi0949), .ZN(new_n8428_));
  NAND2_X1   g05992(.A1(new_n2875_), .A2(new_n2786_), .ZN(new_n8429_));
  NOR2_X1    g05993(.A1(new_n8429_), .A2(new_n2749_), .ZN(new_n8430_));
  AOI22_X1   g05994(.A1(new_n8426_), .A2(new_n8422_), .B1(new_n8430_), .B2(new_n8428_), .ZN(new_n8431_));
  NAND2_X1   g05995(.A1(new_n8431_), .A2(new_n8417_), .ZN(new_n8432_));
  NAND2_X1   g05996(.A1(new_n8432_), .A2(new_n8421_), .ZN(new_n8433_));
  NOR2_X1    g05997(.A1(new_n8414_), .A2(new_n8254_), .ZN(new_n8434_));
  NAND4_X1   g05998(.A1(new_n8434_), .A2(new_n8427_), .A3(pi0949), .A4(new_n8420_), .ZN(new_n8435_));
  OAI21_X1   g05999(.A1(new_n8433_), .A2(pi0072), .B(new_n8435_), .ZN(new_n8436_));
  INV_X1     g06000(.I(new_n8436_), .ZN(new_n8437_));
  NOR3_X1    g06001(.A1(new_n8437_), .A2(pi0044), .A3(pi0101), .ZN(new_n8438_));
  INV_X1     g06002(.I(new_n8438_), .ZN(new_n8439_));
  NOR2_X1    g06003(.A1(new_n8377_), .A2(pi0072), .ZN(new_n8440_));
  INV_X1     g06004(.I(new_n8440_), .ZN(new_n8441_));
  NAND3_X1   g06005(.A1(new_n8415_), .A2(new_n2535_), .A3(new_n8420_), .ZN(new_n8442_));
  NAND3_X1   g06006(.A1(new_n8433_), .A2(new_n2821_), .A3(new_n8442_), .ZN(new_n8443_));
  OAI21_X1   g06007(.A1(new_n8443_), .A2(pi0044), .B(new_n8441_), .ZN(new_n8444_));
  AOI21_X1   g06008(.A1(new_n8444_), .A2(new_n8373_), .B(new_n8376_), .ZN(new_n8445_));
  AOI21_X1   g06009(.A1(new_n8439_), .A2(pi0041), .B(new_n8445_), .ZN(new_n8446_));
  NOR2_X1    g06010(.A1(new_n8446_), .A2(pi0228), .ZN(new_n8447_));
  NAND2_X1   g06011(.A1(new_n6686_), .A2(new_n6656_), .ZN(new_n8448_));
  NOR2_X1    g06012(.A1(new_n6683_), .A2(pi1093), .ZN(new_n8449_));
  AOI21_X1   g06013(.A1(new_n8449_), .A2(new_n8448_), .B(pi0044), .ZN(new_n8450_));
  INV_X1     g06014(.I(new_n8450_), .ZN(new_n8451_));
  NOR2_X1    g06015(.A1(new_n6674_), .A2(pi0097), .ZN(new_n8452_));
  OR3_X2     g06016(.A1(new_n3032_), .A2(new_n3030_), .A3(new_n8452_), .Z(new_n8453_));
  AOI21_X1   g06017(.A1(new_n8453_), .A2(new_n6720_), .B(new_n2762_), .ZN(new_n8454_));
  OAI21_X1   g06018(.A1(new_n8454_), .A2(new_n6664_), .B(new_n6665_), .ZN(new_n8455_));
  AOI21_X1   g06019(.A1(new_n8455_), .A2(new_n2744_), .B(new_n2832_), .ZN(new_n8456_));
  NOR2_X1    g06020(.A1(new_n8456_), .A2(pi0096), .ZN(new_n8457_));
  NOR2_X1    g06021(.A1(new_n6659_), .A2(new_n2536_), .ZN(new_n8458_));
  NOR2_X1    g06022(.A1(new_n6656_), .A2(pi0072), .ZN(new_n8459_));
  NAND2_X1   g06023(.A1(new_n8458_), .A2(new_n8459_), .ZN(new_n8460_));
  OAI21_X1   g06024(.A1(new_n8457_), .A2(new_n8460_), .B(new_n8448_), .ZN(new_n8461_));
  NOR2_X1    g06025(.A1(new_n8461_), .A2(new_n3041_), .ZN(new_n8462_));
  NOR2_X1    g06026(.A1(new_n8451_), .A2(new_n8462_), .ZN(new_n8463_));
  NAND2_X1   g06027(.A1(new_n8463_), .A2(new_n8373_), .ZN(new_n8464_));
  NAND2_X1   g06028(.A1(new_n8464_), .A2(pi0041), .ZN(new_n8465_));
  NAND2_X1   g06029(.A1(new_n8465_), .A2(new_n3025_), .ZN(new_n8466_));
  INV_X1     g06030(.I(new_n8458_), .ZN(new_n8467_));
  OAI21_X1   g06031(.A1(new_n6682_), .A2(new_n8467_), .B(new_n8459_), .ZN(new_n8468_));
  INV_X1     g06032(.I(new_n8468_), .ZN(new_n8469_));
  NOR3_X1    g06033(.A1(new_n6686_), .A2(pi0072), .A3(new_n6655_), .ZN(new_n8470_));
  NOR3_X1    g06034(.A1(new_n8469_), .A2(pi1093), .A3(new_n8470_), .ZN(new_n8471_));
  INV_X1     g06035(.I(new_n8471_), .ZN(new_n8472_));
  OAI21_X1   g06036(.A1(new_n8461_), .A2(pi0072), .B(pi1093), .ZN(new_n8473_));
  NAND2_X1   g06037(.A1(new_n8472_), .A2(new_n8473_), .ZN(new_n8474_));
  OAI21_X1   g06038(.A1(new_n8474_), .A2(pi0044), .B(new_n8441_), .ZN(new_n8475_));
  AOI21_X1   g06039(.A1(new_n8475_), .A2(new_n8373_), .B(new_n8376_), .ZN(new_n8476_));
  AOI21_X1   g06040(.A1(pi1093), .A2(new_n6687_), .B(new_n8451_), .ZN(new_n8477_));
  INV_X1     g06041(.I(new_n8477_), .ZN(new_n8478_));
  NOR2_X1    g06042(.A1(new_n8478_), .A2(pi0101), .ZN(new_n8479_));
  NOR3_X1    g06043(.A1(new_n8471_), .A2(pi0072), .A3(new_n6686_), .ZN(new_n8480_));
  AOI21_X1   g06044(.A1(new_n8480_), .A2(new_n8377_), .B(new_n8440_), .ZN(new_n8481_));
  INV_X1     g06045(.I(new_n8481_), .ZN(new_n8482_));
  AOI21_X1   g06046(.A1(new_n8482_), .A2(new_n8373_), .B(new_n8376_), .ZN(new_n8483_));
  INV_X1     g06047(.I(new_n8483_), .ZN(new_n8484_));
  OAI21_X1   g06048(.A1(new_n8346_), .A2(new_n8479_), .B(new_n8484_), .ZN(new_n8485_));
  OAI22_X1   g06049(.A1(new_n8485_), .A2(new_n3025_), .B1(new_n8466_), .B2(new_n8476_), .ZN(new_n8486_));
  OAI21_X1   g06050(.A1(new_n8486_), .A2(new_n2458_), .B(new_n2627_), .ZN(new_n8487_));
  OAI21_X1   g06051(.A1(new_n8487_), .A2(new_n8447_), .B(new_n8410_), .ZN(new_n8488_));
  NOR2_X1    g06052(.A1(new_n2702_), .A2(pi0038), .ZN(new_n8489_));
  NAND2_X1   g06053(.A1(new_n8370_), .A2(new_n8363_), .ZN(new_n8490_));
  INV_X1     g06054(.I(new_n8372_), .ZN(new_n8491_));
  AOI21_X1   g06055(.A1(new_n2821_), .A2(new_n8200_), .B(new_n8401_), .ZN(new_n8492_));
  INV_X1     g06056(.I(new_n8492_), .ZN(new_n8493_));
  NAND2_X1   g06057(.A1(new_n8493_), .A2(new_n8491_), .ZN(new_n8494_));
  OAI21_X1   g06058(.A1(new_n8371_), .A2(new_n8491_), .B(new_n8494_), .ZN(new_n8495_));
  NAND2_X1   g06059(.A1(new_n8390_), .A2(pi0041), .ZN(new_n8496_));
  NAND3_X1   g06060(.A1(new_n8495_), .A2(new_n8369_), .A3(new_n8496_), .ZN(new_n8497_));
  NAND3_X1   g06061(.A1(new_n8497_), .A2(new_n2627_), .A3(new_n8490_), .ZN(new_n8498_));
  NAND2_X1   g06062(.A1(new_n8498_), .A2(new_n8368_), .ZN(new_n8499_));
  OAI21_X1   g06063(.A1(new_n8365_), .A2(new_n3265_), .B(new_n3458_), .ZN(new_n8500_));
  AOI21_X1   g06064(.A1(new_n8499_), .A2(new_n8489_), .B(new_n8500_), .ZN(new_n8501_));
  AOI21_X1   g06065(.A1(new_n8488_), .A2(new_n8501_), .B(new_n8406_), .ZN(new_n8502_));
  OAI21_X1   g06066(.A1(new_n8502_), .A2(new_n8397_), .B(new_n6645_), .ZN(new_n8503_));
  AOI21_X1   g06067(.A1(new_n8503_), .A2(new_n8367_), .B(new_n8353_), .ZN(po0199));
  INV_X1     g06068(.I(pi0042), .ZN(new_n8505_));
  NOR2_X1    g06069(.A1(new_n8505_), .A2(pi0072), .ZN(new_n8506_));
  NOR2_X1    g06070(.A1(new_n8506_), .A2(pi0039), .ZN(new_n8507_));
  INV_X1     g06071(.I(new_n8507_), .ZN(new_n8508_));
  INV_X1     g06072(.I(pi0212), .ZN(new_n8509_));
  INV_X1     g06073(.I(pi0211), .ZN(new_n8510_));
  INV_X1     g06074(.I(pi0214), .ZN(new_n8511_));
  NOR2_X1    g06075(.A1(new_n8510_), .A2(new_n8511_), .ZN(new_n8512_));
  INV_X1     g06076(.I(new_n8512_), .ZN(new_n8513_));
  NOR2_X1    g06077(.A1(new_n8513_), .A2(new_n8509_), .ZN(new_n8514_));
  NOR2_X1    g06078(.A1(new_n8514_), .A2(pi0219), .ZN(new_n8515_));
  AOI21_X1   g06079(.A1(new_n6697_), .A2(new_n3361_), .B(pi0072), .ZN(new_n8516_));
  INV_X1     g06080(.I(new_n8516_), .ZN(new_n8517_));
  OAI21_X1   g06081(.A1(new_n8517_), .A2(new_n8515_), .B(pi0039), .ZN(new_n8518_));
  NAND2_X1   g06082(.A1(new_n8518_), .A2(new_n8508_), .ZN(new_n8519_));
  INV_X1     g06083(.I(new_n8515_), .ZN(new_n8520_));
  INV_X1     g06084(.I(pi0207), .ZN(new_n8521_));
  INV_X1     g06085(.I(pi0208), .ZN(new_n8522_));
  NOR2_X1    g06086(.A1(new_n8521_), .A2(new_n8522_), .ZN(new_n8523_));
  INV_X1     g06087(.I(new_n8523_), .ZN(new_n8524_));
  INV_X1     g06088(.I(pi0199), .ZN(new_n8525_));
  NOR2_X1    g06089(.A1(new_n8525_), .A2(pi0072), .ZN(new_n8526_));
  OAI21_X1   g06090(.A1(new_n8526_), .A2(pi0232), .B(new_n2628_), .ZN(new_n8527_));
  NOR2_X1    g06091(.A1(new_n8354_), .A2(pi0072), .ZN(new_n8528_));
  NAND2_X1   g06092(.A1(new_n8528_), .A2(pi0199), .ZN(new_n8529_));
  AOI21_X1   g06093(.A1(new_n8529_), .A2(pi0232), .B(new_n8527_), .ZN(new_n8530_));
  INV_X1     g06094(.I(pi0200), .ZN(new_n8531_));
  NOR2_X1    g06095(.A1(new_n8531_), .A2(pi0072), .ZN(new_n8532_));
  OAI21_X1   g06096(.A1(new_n8532_), .A2(pi0232), .B(new_n2628_), .ZN(new_n8533_));
  NAND2_X1   g06097(.A1(new_n8528_), .A2(pi0200), .ZN(new_n8534_));
  AOI21_X1   g06098(.A1(new_n8534_), .A2(pi0232), .B(new_n8533_), .ZN(new_n8535_));
  NOR2_X1    g06099(.A1(new_n8535_), .A2(new_n2627_), .ZN(new_n8536_));
  INV_X1     g06100(.I(new_n8536_), .ZN(new_n8537_));
  NOR2_X1    g06101(.A1(new_n8537_), .A2(new_n8530_), .ZN(new_n8538_));
  NOR2_X1    g06102(.A1(new_n8538_), .A2(new_n8507_), .ZN(new_n8539_));
  AOI21_X1   g06103(.A1(new_n8539_), .A2(new_n6648_), .B(new_n8524_), .ZN(new_n8540_));
  NOR2_X1    g06104(.A1(new_n3026_), .A2(pi0115), .ZN(new_n8541_));
  INV_X1     g06105(.I(new_n8541_), .ZN(new_n8542_));
  AOI21_X1   g06106(.A1(new_n8506_), .A2(new_n8542_), .B(new_n6819_), .ZN(new_n8543_));
  INV_X1     g06107(.I(new_n8543_), .ZN(new_n8544_));
  INV_X1     g06108(.I(pi0114), .ZN(new_n8545_));
  NOR2_X1    g06109(.A1(new_n8506_), .A2(new_n8545_), .ZN(new_n8546_));
  NOR2_X1    g06110(.A1(new_n8542_), .A2(new_n8546_), .ZN(new_n8547_));
  NOR2_X1    g06111(.A1(new_n8383_), .A2(new_n5313_), .ZN(new_n8548_));
  INV_X1     g06112(.I(new_n8548_), .ZN(new_n8549_));
  NOR2_X1    g06113(.A1(new_n8549_), .A2(new_n5316_), .ZN(new_n8550_));
  INV_X1     g06114(.I(new_n8550_), .ZN(new_n8551_));
  AOI21_X1   g06115(.A1(new_n8551_), .A2(new_n8506_), .B(pi0114), .ZN(new_n8552_));
  NOR2_X1    g06116(.A1(new_n8388_), .A2(new_n5311_), .ZN(new_n8553_));
  NAND2_X1   g06117(.A1(new_n8553_), .A2(new_n5315_), .ZN(new_n8554_));
  NOR2_X1    g06118(.A1(new_n8554_), .A2(new_n8200_), .ZN(new_n8555_));
  INV_X1     g06119(.I(new_n8555_), .ZN(new_n8556_));
  NOR3_X1    g06120(.A1(new_n8556_), .A2(pi0114), .A3(new_n5314_), .ZN(new_n8557_));
  INV_X1     g06121(.I(new_n8557_), .ZN(new_n8558_));
  NOR2_X1    g06122(.A1(new_n8558_), .A2(new_n6707_), .ZN(new_n8559_));
  INV_X1     g06123(.I(new_n8559_), .ZN(new_n8560_));
  OAI21_X1   g06124(.A1(pi0042), .A2(new_n8560_), .B(new_n8552_), .ZN(new_n8561_));
  AOI21_X1   g06125(.A1(new_n8561_), .A2(new_n8547_), .B(new_n8544_), .ZN(new_n8562_));
  INV_X1     g06126(.I(new_n8506_), .ZN(new_n8563_));
  NAND2_X1   g06127(.A1(new_n6819_), .A2(new_n8563_), .ZN(new_n8564_));
  NAND2_X1   g06128(.A1(new_n8564_), .A2(new_n2626_), .ZN(new_n8565_));
  AOI21_X1   g06129(.A1(new_n5792_), .A2(new_n8506_), .B(pi0039), .ZN(new_n8566_));
  OAI21_X1   g06130(.A1(new_n8562_), .A2(new_n8565_), .B(new_n8566_), .ZN(new_n8567_));
  OAI21_X1   g06131(.A1(new_n8530_), .A2(new_n8537_), .B(new_n8567_), .ZN(new_n8568_));
  AOI21_X1   g06132(.A1(new_n8568_), .A2(pi0075), .B(new_n6648_), .ZN(new_n8569_));
  NOR2_X1    g06133(.A1(new_n8539_), .A2(new_n3265_), .ZN(new_n8570_));
  NOR2_X1    g06134(.A1(new_n8570_), .A2(pi0087), .ZN(new_n8571_));
  INV_X1     g06135(.I(new_n8547_), .ZN(new_n8572_));
  NAND2_X1   g06136(.A1(new_n8558_), .A2(new_n8505_), .ZN(new_n8573_));
  NOR3_X1    g06137(.A1(new_n8379_), .A2(pi0044), .A3(new_n5313_), .ZN(new_n8574_));
  INV_X1     g06138(.I(new_n8574_), .ZN(new_n8575_));
  NOR2_X1    g06139(.A1(new_n8575_), .A2(new_n5316_), .ZN(new_n8576_));
  INV_X1     g06140(.I(new_n8576_), .ZN(new_n8577_));
  NOR2_X1    g06141(.A1(new_n8577_), .A2(new_n8200_), .ZN(new_n8578_));
  NOR2_X1    g06142(.A1(new_n8578_), .A2(pi0072), .ZN(new_n8579_));
  INV_X1     g06143(.I(new_n8579_), .ZN(new_n8580_));
  NAND2_X1   g06144(.A1(new_n8580_), .A2(pi0042), .ZN(new_n8581_));
  AOI21_X1   g06145(.A1(new_n8581_), .A2(new_n8573_), .B(pi0114), .ZN(new_n8582_));
  OAI21_X1   g06146(.A1(new_n8582_), .A2(new_n8572_), .B(new_n8543_), .ZN(new_n8583_));
  AOI21_X1   g06147(.A1(new_n8583_), .A2(new_n8564_), .B(pi0039), .ZN(new_n8584_));
  OAI21_X1   g06148(.A1(new_n8584_), .A2(new_n8538_), .B(new_n8489_), .ZN(new_n8585_));
  NAND2_X1   g06149(.A1(new_n8585_), .A2(new_n8571_), .ZN(new_n8586_));
  INV_X1     g06150(.I(pi0115), .ZN(new_n8587_));
  NOR2_X1    g06151(.A1(new_n8506_), .A2(new_n8587_), .ZN(new_n8588_));
  NOR2_X1    g06152(.A1(new_n8439_), .A2(new_n5311_), .ZN(new_n8589_));
  INV_X1     g06153(.I(new_n8589_), .ZN(new_n8590_));
  NOR2_X1    g06154(.A1(new_n8590_), .A2(new_n5316_), .ZN(new_n8591_));
  NOR2_X1    g06155(.A1(new_n8591_), .A2(pi0042), .ZN(new_n8592_));
  NOR2_X1    g06156(.A1(new_n8592_), .A2(new_n8546_), .ZN(new_n8593_));
  INV_X1     g06157(.I(pi0116), .ZN(new_n8594_));
  NOR2_X1    g06158(.A1(new_n8594_), .A2(pi0072), .ZN(new_n8595_));
  INV_X1     g06159(.I(new_n8595_), .ZN(new_n8596_));
  INV_X1     g06160(.I(pi0113), .ZN(new_n8597_));
  NOR2_X1    g06161(.A1(new_n8597_), .A2(pi0072), .ZN(new_n8598_));
  INV_X1     g06162(.I(pi0099), .ZN(new_n8599_));
  NOR2_X1    g06163(.A1(new_n8599_), .A2(pi0072), .ZN(new_n8600_));
  INV_X1     g06164(.I(new_n8600_), .ZN(new_n8601_));
  AOI22_X1   g06165(.A1(new_n8445_), .A2(new_n8601_), .B1(pi0072), .B2(new_n5311_), .ZN(new_n8602_));
  AOI21_X1   g06166(.A1(new_n8602_), .A2(new_n8597_), .B(new_n8598_), .ZN(new_n8603_));
  OAI21_X1   g06167(.A1(new_n8603_), .A2(pi0116), .B(new_n8596_), .ZN(new_n8604_));
  INV_X1     g06168(.I(new_n8604_), .ZN(new_n8605_));
  NAND3_X1   g06169(.A1(new_n8605_), .A2(pi0042), .A3(new_n8545_), .ZN(new_n8606_));
  AOI21_X1   g06170(.A1(new_n8606_), .A2(new_n8593_), .B(pi0115), .ZN(new_n8607_));
  NOR3_X1    g06171(.A1(new_n8607_), .A2(pi0228), .A3(new_n8588_), .ZN(new_n8608_));
  NOR2_X1    g06172(.A1(new_n8464_), .A2(new_n5311_), .ZN(new_n8609_));
  INV_X1     g06173(.I(new_n8609_), .ZN(new_n8610_));
  NOR2_X1    g06174(.A1(new_n8610_), .A2(new_n5316_), .ZN(new_n8611_));
  INV_X1     g06175(.I(new_n8611_), .ZN(new_n8612_));
  AOI21_X1   g06176(.A1(new_n8612_), .A2(new_n8505_), .B(new_n8546_), .ZN(new_n8613_));
  NAND3_X1   g06177(.A1(new_n8476_), .A2(new_n8599_), .A3(new_n8597_), .ZN(new_n8614_));
  OAI21_X1   g06178(.A1(new_n5311_), .A2(pi0113), .B(pi0072), .ZN(new_n8615_));
  NAND2_X1   g06179(.A1(new_n8614_), .A2(new_n8615_), .ZN(new_n8616_));
  INV_X1     g06180(.I(new_n8616_), .ZN(new_n8617_));
  AOI21_X1   g06181(.A1(new_n8617_), .A2(new_n8594_), .B(new_n8595_), .ZN(new_n8618_));
  NAND3_X1   g06182(.A1(new_n8618_), .A2(pi0042), .A3(new_n8545_), .ZN(new_n8619_));
  AOI21_X1   g06183(.A1(new_n8619_), .A2(new_n8613_), .B(new_n8542_), .ZN(new_n8620_));
  INV_X1     g06184(.I(new_n8598_), .ZN(new_n8621_));
  NAND3_X1   g06185(.A1(new_n8483_), .A2(new_n8599_), .A3(new_n8621_), .ZN(new_n8622_));
  NAND2_X1   g06186(.A1(new_n8622_), .A2(new_n8615_), .ZN(new_n8623_));
  OAI21_X1   g06187(.A1(new_n8623_), .A2(pi0116), .B(new_n8596_), .ZN(new_n8624_));
  OR2_X2     g06188(.A1(new_n8624_), .A2(new_n8505_), .Z(new_n8625_));
  INV_X1     g06189(.I(new_n8479_), .ZN(new_n8626_));
  NOR2_X1    g06190(.A1(new_n8626_), .A2(new_n5311_), .ZN(new_n8627_));
  INV_X1     g06191(.I(new_n8627_), .ZN(new_n8628_));
  NOR2_X1    g06192(.A1(new_n8628_), .A2(new_n5316_), .ZN(new_n8629_));
  INV_X1     g06193(.I(new_n8629_), .ZN(new_n8630_));
  NAND2_X1   g06194(.A1(new_n8630_), .A2(new_n8505_), .ZN(new_n8631_));
  AOI21_X1   g06195(.A1(new_n8631_), .A2(new_n8625_), .B(pi0114), .ZN(new_n8632_));
  OAI21_X1   g06196(.A1(new_n8632_), .A2(new_n8546_), .B(new_n8587_), .ZN(new_n8633_));
  NOR2_X1    g06197(.A1(new_n8633_), .A2(new_n3025_), .ZN(new_n8634_));
  NOR4_X1    g06198(.A1(new_n8634_), .A2(new_n2458_), .A3(new_n8588_), .A4(new_n8620_), .ZN(new_n8635_));
  OR3_X2     g06199(.A1(new_n8635_), .A2(pi0039), .A3(new_n8608_), .Z(new_n8636_));
  INV_X1     g06200(.I(new_n8407_), .ZN(new_n8637_));
  NOR2_X1    g06201(.A1(new_n8354_), .A2(new_n2821_), .ZN(new_n8638_));
  AOI21_X1   g06202(.A1(new_n8637_), .A2(new_n8354_), .B(new_n8638_), .ZN(new_n8639_));
  NOR2_X1    g06203(.A1(pi0199), .A2(pi0200), .ZN(new_n8640_));
  INV_X1     g06204(.I(new_n8640_), .ZN(new_n8641_));
  AOI21_X1   g06205(.A1(new_n8639_), .A2(new_n8641_), .B(new_n5666_), .ZN(new_n8642_));
  AND2_X2    g06206(.A1(new_n8527_), .A2(new_n8533_), .Z(new_n8643_));
  OAI21_X1   g06207(.A1(new_n8642_), .A2(new_n8643_), .B(pi0039), .ZN(new_n8644_));
  NAND2_X1   g06208(.A1(new_n8636_), .A2(new_n8644_), .ZN(new_n8645_));
  AOI21_X1   g06209(.A1(new_n8645_), .A2(new_n3270_), .B(new_n8586_), .ZN(new_n8646_));
  NOR2_X1    g06210(.A1(new_n8575_), .A2(new_n2458_), .ZN(new_n8647_));
  AOI21_X1   g06211(.A1(new_n8647_), .A2(new_n5319_), .B(new_n8563_), .ZN(new_n8648_));
  NOR2_X1    g06212(.A1(new_n8554_), .A2(new_n2458_), .ZN(new_n8649_));
  INV_X1     g06213(.I(new_n8649_), .ZN(new_n8650_));
  NOR2_X1    g06214(.A1(new_n8650_), .A2(new_n5318_), .ZN(new_n8651_));
  NAND2_X1   g06215(.A1(new_n8651_), .A2(new_n8505_), .ZN(new_n8652_));
  NAND2_X1   g06216(.A1(new_n8652_), .A2(new_n3272_), .ZN(new_n8653_));
  AOI21_X1   g06217(.A1(new_n8507_), .A2(new_n3271_), .B(new_n3458_), .ZN(new_n8654_));
  OAI21_X1   g06218(.A1(new_n8648_), .A2(new_n8653_), .B(new_n8654_), .ZN(new_n8655_));
  OAI21_X1   g06219(.A1(new_n8655_), .A2(new_n8538_), .B(new_n3465_), .ZN(new_n8656_));
  OAI21_X1   g06220(.A1(new_n8646_), .A2(new_n8656_), .B(new_n8569_), .ZN(new_n8657_));
  OAI21_X1   g06221(.A1(new_n2627_), .A2(new_n8530_), .B(new_n8567_), .ZN(new_n8658_));
  AOI21_X1   g06222(.A1(new_n8658_), .A2(pi0075), .B(new_n6648_), .ZN(new_n8659_));
  NOR2_X1    g06223(.A1(new_n8530_), .A2(new_n2627_), .ZN(new_n8660_));
  OAI21_X1   g06224(.A1(new_n8655_), .A2(new_n8660_), .B(new_n3465_), .ZN(new_n8661_));
  AOI21_X1   g06225(.A1(new_n8639_), .A2(pi0199), .B(new_n5666_), .ZN(new_n8662_));
  OAI21_X1   g06226(.A1(new_n8662_), .A2(new_n8527_), .B(pi0039), .ZN(new_n8663_));
  AOI21_X1   g06227(.A1(new_n8636_), .A2(new_n8663_), .B(new_n3271_), .ZN(new_n8664_));
  NOR2_X1    g06228(.A1(new_n8660_), .A2(new_n8507_), .ZN(new_n8665_));
  NOR2_X1    g06229(.A1(new_n8665_), .A2(new_n3265_), .ZN(new_n8666_));
  INV_X1     g06230(.I(new_n8489_), .ZN(new_n8667_));
  NOR2_X1    g06231(.A1(new_n8584_), .A2(new_n8660_), .ZN(new_n8668_));
  NOR2_X1    g06232(.A1(new_n8668_), .A2(new_n8667_), .ZN(new_n8669_));
  NOR4_X1    g06233(.A1(new_n8664_), .A2(pi0087), .A3(new_n8666_), .A4(new_n8669_), .ZN(new_n8670_));
  OAI21_X1   g06234(.A1(new_n8670_), .A2(new_n8661_), .B(new_n8659_), .ZN(new_n8671_));
  AOI21_X1   g06235(.A1(new_n8665_), .A2(new_n6648_), .B(new_n8523_), .ZN(new_n8672_));
  AOI22_X1   g06236(.A1(new_n8671_), .A2(new_n8672_), .B1(new_n8540_), .B2(new_n8657_), .ZN(new_n8673_));
  NOR2_X1    g06237(.A1(new_n8673_), .A2(new_n8520_), .ZN(new_n8674_));
  NOR2_X1    g06238(.A1(new_n8517_), .A2(new_n2628_), .ZN(new_n8675_));
  NOR2_X1    g06239(.A1(new_n8675_), .A2(new_n2627_), .ZN(new_n8676_));
  INV_X1     g06240(.I(new_n8676_), .ZN(new_n8677_));
  NOR2_X1    g06241(.A1(new_n8677_), .A2(new_n8530_), .ZN(new_n8678_));
  INV_X1     g06242(.I(new_n8678_), .ZN(new_n8679_));
  NAND2_X1   g06243(.A1(new_n8679_), .A2(new_n8508_), .ZN(new_n8680_));
  OAI21_X1   g06244(.A1(new_n8680_), .A2(new_n6645_), .B(new_n8520_), .ZN(new_n8681_));
  NAND2_X1   g06245(.A1(new_n8567_), .A2(new_n8679_), .ZN(new_n8682_));
  AOI21_X1   g06246(.A1(new_n8682_), .A2(pi0075), .B(new_n6648_), .ZN(new_n8683_));
  AOI21_X1   g06247(.A1(new_n8680_), .A2(pi0038), .B(pi0087), .ZN(new_n8684_));
  OAI21_X1   g06248(.A1(new_n8584_), .A2(new_n8678_), .B(new_n8489_), .ZN(new_n8685_));
  NAND2_X1   g06249(.A1(new_n8685_), .A2(new_n8684_), .ZN(new_n8686_));
  NOR2_X1    g06250(.A1(new_n5666_), .A2(new_n2628_), .ZN(new_n8687_));
  INV_X1     g06251(.I(new_n8687_), .ZN(new_n8688_));
  NOR2_X1    g06252(.A1(new_n8516_), .A2(new_n8688_), .ZN(new_n8689_));
  OAI21_X1   g06253(.A1(new_n8637_), .A2(new_n8349_), .B(new_n8689_), .ZN(new_n8690_));
  NOR2_X1    g06254(.A1(pi0199), .A2(pi0299), .ZN(new_n8691_));
  OAI21_X1   g06255(.A1(new_n8691_), .A2(pi0072), .B(new_n5666_), .ZN(new_n8692_));
  NAND2_X1   g06256(.A1(new_n8662_), .A2(new_n2628_), .ZN(new_n8693_));
  AND3_X2    g06257(.A1(new_n8693_), .A2(new_n8690_), .A3(new_n8692_), .Z(new_n8694_));
  OAI21_X1   g06258(.A1(new_n2627_), .A2(new_n8694_), .B(new_n8636_), .ZN(new_n8695_));
  AOI21_X1   g06259(.A1(new_n8695_), .A2(new_n3270_), .B(new_n8686_), .ZN(new_n8696_));
  OAI21_X1   g06260(.A1(new_n8655_), .A2(new_n8678_), .B(new_n3465_), .ZN(new_n8697_));
  OAI21_X1   g06261(.A1(new_n8696_), .A2(new_n8697_), .B(new_n8683_), .ZN(new_n8698_));
  OAI21_X1   g06262(.A1(new_n8537_), .A2(new_n8679_), .B(new_n8567_), .ZN(new_n8699_));
  AOI21_X1   g06263(.A1(new_n8699_), .A2(pi0075), .B(new_n6648_), .ZN(new_n8700_));
  NOR2_X1    g06264(.A1(new_n8679_), .A2(new_n8537_), .ZN(new_n8701_));
  NOR2_X1    g06265(.A1(new_n8584_), .A2(new_n8701_), .ZN(new_n8702_));
  OAI22_X1   g06266(.A1(new_n8702_), .A2(new_n8667_), .B1(new_n8571_), .B2(new_n8684_), .ZN(new_n8703_));
  OAI21_X1   g06267(.A1(new_n8532_), .A2(new_n8692_), .B(new_n8690_), .ZN(new_n8704_));
  AND2_X2    g06268(.A1(new_n8642_), .A2(new_n2628_), .Z(new_n8705_));
  OAI21_X1   g06269(.A1(new_n8705_), .A2(new_n8704_), .B(pi0039), .ZN(new_n8706_));
  NAND2_X1   g06270(.A1(new_n8636_), .A2(new_n8706_), .ZN(new_n8707_));
  AOI21_X1   g06271(.A1(new_n8707_), .A2(new_n3270_), .B(new_n8703_), .ZN(new_n8708_));
  OAI21_X1   g06272(.A1(new_n8655_), .A2(new_n8701_), .B(new_n3465_), .ZN(new_n8709_));
  OAI21_X1   g06273(.A1(new_n8708_), .A2(new_n8709_), .B(new_n8700_), .ZN(new_n8710_));
  AOI22_X1   g06274(.A1(new_n8698_), .A2(new_n8524_), .B1(new_n8540_), .B2(new_n8710_), .ZN(new_n8711_));
  OAI21_X1   g06275(.A1(new_n8711_), .A2(new_n8681_), .B(new_n6643_), .ZN(new_n8712_));
  OAI22_X1   g06276(.A1(new_n8712_), .A2(new_n8674_), .B1(new_n6643_), .B2(new_n8519_), .ZN(po0200));
  INV_X1     g06277(.I(pi0043), .ZN(new_n8714_));
  NOR2_X1    g06278(.A1(new_n8714_), .A2(pi0072), .ZN(new_n8715_));
  INV_X1     g06279(.I(new_n8715_), .ZN(new_n8716_));
  NAND2_X1   g06280(.A1(new_n8716_), .A2(new_n2627_), .ZN(new_n8717_));
  NOR2_X1    g06281(.A1(new_n8677_), .A2(new_n8535_), .ZN(new_n8718_));
  INV_X1     g06282(.I(new_n8718_), .ZN(new_n8719_));
  NAND2_X1   g06283(.A1(new_n8719_), .A2(new_n8717_), .ZN(new_n8720_));
  OAI21_X1   g06284(.A1(new_n8720_), .A2(new_n6645_), .B(new_n8524_), .ZN(new_n8721_));
  NOR3_X1    g06285(.A1(pi0042), .A2(pi0114), .A3(pi0115), .ZN(new_n8722_));
  INV_X1     g06286(.I(new_n8722_), .ZN(new_n8723_));
  NOR2_X1    g06287(.A1(new_n8370_), .A2(new_n8723_), .ZN(new_n8724_));
  NAND2_X1   g06288(.A1(new_n8724_), .A2(new_n2626_), .ZN(new_n8725_));
  NOR2_X1    g06289(.A1(new_n8550_), .A2(pi0072), .ZN(new_n8726_));
  INV_X1     g06290(.I(pi0052), .ZN(new_n8727_));
  NOR2_X1    g06291(.A1(new_n8727_), .A2(pi0043), .ZN(new_n8728_));
  NOR2_X1    g06292(.A1(new_n8556_), .A2(new_n6707_), .ZN(new_n8729_));
  AOI22_X1   g06293(.A1(new_n8726_), .A2(pi0043), .B1(new_n8728_), .B2(new_n8729_), .ZN(new_n8730_));
  NOR2_X1    g06294(.A1(new_n8730_), .A2(new_n8725_), .ZN(new_n8731_));
  AOI21_X1   g06295(.A1(new_n8715_), .A2(new_n8725_), .B(new_n8731_), .ZN(new_n8732_));
  NAND2_X1   g06296(.A1(new_n8732_), .A2(new_n2627_), .ZN(new_n8733_));
  NAND2_X1   g06297(.A1(new_n8733_), .A2(new_n8719_), .ZN(new_n8734_));
  AOI21_X1   g06298(.A1(new_n8734_), .A2(pi0075), .B(new_n6648_), .ZN(new_n8735_));
  AOI21_X1   g06299(.A1(new_n8720_), .A2(pi0038), .B(pi0087), .ZN(new_n8736_));
  INV_X1     g06300(.I(new_n8728_), .ZN(new_n8737_));
  OAI22_X1   g06301(.A1(new_n8580_), .A2(new_n8714_), .B1(new_n8556_), .B2(new_n8737_), .ZN(new_n8738_));
  NAND2_X1   g06302(.A1(new_n8738_), .A2(new_n8724_), .ZN(new_n8739_));
  OAI21_X1   g06303(.A1(new_n8716_), .A2(new_n8724_), .B(new_n8739_), .ZN(new_n8740_));
  NOR2_X1    g06304(.A1(new_n8740_), .A2(pi0039), .ZN(new_n8741_));
  OAI21_X1   g06305(.A1(new_n8741_), .A2(new_n8718_), .B(new_n8489_), .ZN(new_n8742_));
  NAND2_X1   g06306(.A1(new_n8742_), .A2(new_n8736_), .ZN(new_n8743_));
  NOR2_X1    g06307(.A1(new_n8609_), .A2(new_n3026_), .ZN(new_n8744_));
  NOR2_X1    g06308(.A1(new_n8627_), .A2(new_n3025_), .ZN(new_n8745_));
  NOR2_X1    g06309(.A1(new_n8745_), .A2(new_n8744_), .ZN(new_n8746_));
  INV_X1     g06310(.I(new_n8746_), .ZN(new_n8747_));
  NOR3_X1    g06311(.A1(new_n8747_), .A2(new_n2458_), .A3(new_n5316_), .ZN(new_n8748_));
  AOI21_X1   g06312(.A1(new_n2458_), .A2(new_n8591_), .B(new_n8748_), .ZN(new_n8749_));
  NAND2_X1   g06313(.A1(new_n8749_), .A2(new_n8714_), .ZN(new_n8750_));
  AOI21_X1   g06314(.A1(new_n8750_), .A2(new_n8722_), .B(new_n8715_), .ZN(new_n8751_));
  INV_X1     g06315(.I(new_n8618_), .ZN(new_n8752_));
  NAND2_X1   g06316(.A1(new_n8752_), .A2(new_n3025_), .ZN(new_n8753_));
  NAND2_X1   g06317(.A1(new_n8624_), .A2(new_n3026_), .ZN(new_n8754_));
  AOI21_X1   g06318(.A1(new_n8753_), .A2(new_n8754_), .B(new_n2458_), .ZN(new_n8755_));
  NOR2_X1    g06319(.A1(new_n8605_), .A2(pi0228), .ZN(new_n8756_));
  NOR2_X1    g06320(.A1(new_n8755_), .A2(new_n8756_), .ZN(new_n8757_));
  INV_X1     g06321(.I(new_n8757_), .ZN(new_n8758_));
  NOR3_X1    g06322(.A1(new_n8758_), .A2(new_n8714_), .A3(new_n8723_), .ZN(new_n8759_));
  OAI21_X1   g06323(.A1(new_n8759_), .A2(new_n8751_), .B(new_n2627_), .ZN(new_n8760_));
  NOR2_X1    g06324(.A1(pi0200), .A2(pi0299), .ZN(new_n8761_));
  OAI21_X1   g06325(.A1(new_n8761_), .A2(pi0072), .B(new_n5666_), .ZN(new_n8762_));
  AOI21_X1   g06326(.A1(new_n8639_), .A2(pi0200), .B(new_n5666_), .ZN(new_n8763_));
  NAND2_X1   g06327(.A1(new_n8763_), .A2(new_n2628_), .ZN(new_n8764_));
  NAND3_X1   g06328(.A1(new_n8764_), .A2(new_n8690_), .A3(new_n8762_), .ZN(new_n8765_));
  NAND2_X1   g06329(.A1(new_n8765_), .A2(pi0039), .ZN(new_n8766_));
  AOI21_X1   g06330(.A1(new_n8760_), .A2(new_n8766_), .B(new_n3271_), .ZN(new_n8767_));
  NOR2_X1    g06331(.A1(new_n8723_), .A2(new_n2458_), .ZN(new_n8768_));
  NAND2_X1   g06332(.A1(new_n8577_), .A2(new_n2821_), .ZN(new_n8769_));
  NOR2_X1    g06333(.A1(new_n8769_), .A2(new_n8714_), .ZN(new_n8770_));
  NOR2_X1    g06334(.A1(new_n8554_), .A2(pi0043), .ZN(new_n8771_));
  OAI21_X1   g06335(.A1(new_n8770_), .A2(new_n8771_), .B(new_n8768_), .ZN(new_n8772_));
  NOR2_X1    g06336(.A1(new_n8768_), .A2(new_n8716_), .ZN(new_n8773_));
  NOR2_X1    g06337(.A1(new_n8773_), .A2(new_n3273_), .ZN(new_n8774_));
  OAI21_X1   g06338(.A1(new_n8717_), .A2(new_n3270_), .B(pi0087), .ZN(new_n8775_));
  AOI21_X1   g06339(.A1(new_n8772_), .A2(new_n8774_), .B(new_n8775_), .ZN(new_n8776_));
  AOI21_X1   g06340(.A1(new_n8776_), .A2(new_n8719_), .B(pi0075), .ZN(new_n8777_));
  OAI21_X1   g06341(.A1(new_n8767_), .A2(new_n8743_), .B(new_n8777_), .ZN(new_n8778_));
  AOI21_X1   g06342(.A1(new_n8778_), .A2(new_n8735_), .B(new_n8721_), .ZN(new_n8779_));
  NOR2_X1    g06343(.A1(new_n8640_), .A2(pi0299), .ZN(new_n8780_));
  INV_X1     g06344(.I(new_n8780_), .ZN(new_n8781_));
  AOI21_X1   g06345(.A1(new_n8781_), .A2(new_n2821_), .B(pi0232), .ZN(new_n8782_));
  NOR2_X1    g06346(.A1(new_n8782_), .A2(pi0299), .ZN(new_n8783_));
  INV_X1     g06347(.I(new_n8783_), .ZN(new_n8784_));
  AOI21_X1   g06348(.A1(new_n8528_), .A2(new_n8640_), .B(new_n5666_), .ZN(new_n8785_));
  NOR2_X1    g06349(.A1(new_n8784_), .A2(new_n8785_), .ZN(new_n8786_));
  NOR2_X1    g06350(.A1(new_n8786_), .A2(new_n2627_), .ZN(new_n8787_));
  INV_X1     g06351(.I(new_n8787_), .ZN(new_n8788_));
  NOR2_X1    g06352(.A1(new_n8788_), .A2(new_n8675_), .ZN(new_n8789_));
  INV_X1     g06353(.I(new_n8789_), .ZN(new_n8790_));
  NAND2_X1   g06354(.A1(new_n8790_), .A2(new_n8717_), .ZN(new_n8791_));
  OAI21_X1   g06355(.A1(new_n8791_), .A2(new_n6645_), .B(new_n8523_), .ZN(new_n8792_));
  AOI21_X1   g06356(.A1(new_n8791_), .A2(pi0038), .B(pi0087), .ZN(new_n8793_));
  OAI21_X1   g06357(.A1(new_n8741_), .A2(new_n8789_), .B(new_n8489_), .ZN(new_n8794_));
  NAND2_X1   g06358(.A1(new_n8794_), .A2(new_n8793_), .ZN(new_n8795_));
  AOI21_X1   g06359(.A1(new_n8639_), .A2(new_n8640_), .B(new_n5666_), .ZN(new_n8796_));
  AOI21_X1   g06360(.A1(new_n8796_), .A2(new_n2628_), .B(new_n8782_), .ZN(new_n8797_));
  NAND2_X1   g06361(.A1(new_n8797_), .A2(new_n8690_), .ZN(new_n8798_));
  NAND2_X1   g06362(.A1(new_n8798_), .A2(pi0039), .ZN(new_n8799_));
  AOI21_X1   g06363(.A1(new_n8760_), .A2(new_n8799_), .B(new_n3271_), .ZN(new_n8800_));
  AOI21_X1   g06364(.A1(new_n8776_), .A2(new_n8790_), .B(pi0075), .ZN(new_n8801_));
  OAI21_X1   g06365(.A1(new_n8800_), .A2(new_n8795_), .B(new_n8801_), .ZN(new_n8802_));
  NAND2_X1   g06366(.A1(new_n8733_), .A2(new_n8790_), .ZN(new_n8803_));
  AOI21_X1   g06367(.A1(new_n8803_), .A2(pi0075), .B(new_n6648_), .ZN(new_n8804_));
  AOI21_X1   g06368(.A1(new_n8802_), .A2(new_n8804_), .B(new_n8792_), .ZN(new_n8805_));
  NOR2_X1    g06369(.A1(new_n8779_), .A2(new_n8805_), .ZN(new_n8806_));
  INV_X1     g06370(.I(pi0219), .ZN(new_n8807_));
  NOR2_X1    g06371(.A1(new_n8807_), .A2(pi0211), .ZN(new_n8808_));
  NOR2_X1    g06372(.A1(new_n8509_), .A2(new_n8511_), .ZN(new_n8809_));
  NOR2_X1    g06373(.A1(new_n8809_), .A2(pi0211), .ZN(new_n8810_));
  INV_X1     g06374(.I(new_n8809_), .ZN(new_n8811_));
  NOR2_X1    g06375(.A1(new_n8811_), .A2(new_n8510_), .ZN(new_n8812_));
  NOR2_X1    g06376(.A1(new_n8812_), .A2(new_n8810_), .ZN(new_n8813_));
  INV_X1     g06377(.I(new_n8813_), .ZN(new_n8814_));
  NOR2_X1    g06378(.A1(new_n8814_), .A2(new_n8808_), .ZN(new_n8815_));
  NAND2_X1   g06379(.A1(new_n8788_), .A2(new_n8717_), .ZN(new_n8816_));
  OAI21_X1   g06380(.A1(new_n8816_), .A2(new_n6645_), .B(new_n8523_), .ZN(new_n8817_));
  NAND2_X1   g06381(.A1(new_n8733_), .A2(new_n8788_), .ZN(new_n8818_));
  AOI21_X1   g06382(.A1(new_n8818_), .A2(pi0075), .B(new_n6648_), .ZN(new_n8819_));
  AOI21_X1   g06383(.A1(new_n8816_), .A2(pi0038), .B(pi0087), .ZN(new_n8820_));
  OAI21_X1   g06384(.A1(new_n8741_), .A2(new_n8787_), .B(new_n8489_), .ZN(new_n8821_));
  NAND2_X1   g06385(.A1(new_n8821_), .A2(new_n8820_), .ZN(new_n8822_));
  OAI21_X1   g06386(.A1(new_n8796_), .A2(new_n8784_), .B(pi0039), .ZN(new_n8823_));
  AOI21_X1   g06387(.A1(new_n8760_), .A2(new_n8823_), .B(new_n3271_), .ZN(new_n8824_));
  NAND2_X1   g06388(.A1(new_n8816_), .A2(new_n2575_), .ZN(new_n8825_));
  AOI21_X1   g06389(.A1(new_n8776_), .A2(new_n8825_), .B(pi0075), .ZN(new_n8826_));
  OAI21_X1   g06390(.A1(new_n8824_), .A2(new_n8822_), .B(new_n8826_), .ZN(new_n8827_));
  AOI21_X1   g06391(.A1(new_n8827_), .A2(new_n8819_), .B(new_n8817_), .ZN(new_n8828_));
  NAND2_X1   g06392(.A1(new_n8537_), .A2(new_n8717_), .ZN(new_n8829_));
  OAI21_X1   g06393(.A1(new_n8829_), .A2(new_n6645_), .B(new_n8524_), .ZN(new_n8830_));
  AOI21_X1   g06394(.A1(new_n8829_), .A2(pi0038), .B(pi0087), .ZN(new_n8831_));
  OAI21_X1   g06395(.A1(new_n8741_), .A2(new_n8536_), .B(new_n8489_), .ZN(new_n8832_));
  NAND2_X1   g06396(.A1(new_n8832_), .A2(new_n8831_), .ZN(new_n8833_));
  OAI21_X1   g06397(.A1(new_n8763_), .A2(new_n8533_), .B(pi0039), .ZN(new_n8834_));
  AOI21_X1   g06398(.A1(new_n8760_), .A2(new_n8834_), .B(new_n3271_), .ZN(new_n8835_));
  AOI21_X1   g06399(.A1(new_n8776_), .A2(new_n8537_), .B(pi0075), .ZN(new_n8836_));
  OAI21_X1   g06400(.A1(new_n8835_), .A2(new_n8833_), .B(new_n8836_), .ZN(new_n8837_));
  NAND2_X1   g06401(.A1(new_n8733_), .A2(new_n8537_), .ZN(new_n8838_));
  AOI21_X1   g06402(.A1(new_n8838_), .A2(pi0075), .B(new_n6648_), .ZN(new_n8839_));
  AOI21_X1   g06403(.A1(new_n8837_), .A2(new_n8839_), .B(new_n8830_), .ZN(new_n8840_));
  NOR3_X1    g06404(.A1(new_n8828_), .A2(new_n8840_), .A3(new_n8815_), .ZN(new_n8841_));
  AOI21_X1   g06405(.A1(new_n8806_), .A2(new_n8815_), .B(new_n8841_), .ZN(new_n8842_));
  NAND2_X1   g06406(.A1(po1038), .A2(new_n8717_), .ZN(new_n8843_));
  AOI21_X1   g06407(.A1(new_n8815_), .A2(new_n8516_), .B(new_n2627_), .ZN(new_n8844_));
  OAI22_X1   g06408(.A1(new_n8842_), .A2(po1038), .B1(new_n8843_), .B2(new_n8844_), .ZN(po0201));
  NOR2_X1    g06409(.A1(new_n8377_), .A2(pi0039), .ZN(new_n8846_));
  NOR2_X1    g06410(.A1(new_n3169_), .A2(new_n6698_), .ZN(new_n8847_));
  AOI21_X1   g06411(.A1(new_n8847_), .A2(pi0039), .B(new_n8846_), .ZN(new_n8848_));
  OR3_X2     g06412(.A1(new_n8848_), .A2(pi0072), .A3(new_n6643_), .Z(new_n8849_));
  NOR2_X1    g06413(.A1(new_n8224_), .A2(new_n2627_), .ZN(new_n8850_));
  OAI21_X1   g06414(.A1(new_n8850_), .A2(new_n8846_), .B(new_n2821_), .ZN(new_n8851_));
  INV_X1     g06415(.I(new_n8851_), .ZN(new_n8852_));
  OAI21_X1   g06416(.A1(new_n8852_), .A2(new_n6645_), .B(new_n6643_), .ZN(new_n8853_));
  NOR2_X1    g06417(.A1(new_n8852_), .A2(new_n2626_), .ZN(new_n8854_));
  OAI21_X1   g06418(.A1(new_n6774_), .A2(new_n8440_), .B(new_n2627_), .ZN(new_n8855_));
  AOI21_X1   g06419(.A1(new_n3026_), .A2(new_n8440_), .B(new_n6819_), .ZN(new_n8856_));
  OAI21_X1   g06420(.A1(new_n8377_), .A2(new_n2821_), .B(pi1091), .ZN(new_n8857_));
  NOR2_X1    g06421(.A1(new_n6705_), .A2(new_n8857_), .ZN(new_n8858_));
  NOR2_X1    g06422(.A1(new_n8386_), .A2(new_n8200_), .ZN(new_n8859_));
  NAND2_X1   g06423(.A1(new_n8859_), .A2(new_n6706_), .ZN(new_n8860_));
  OAI21_X1   g06424(.A1(new_n8382_), .A2(new_n8377_), .B(new_n8860_), .ZN(new_n8861_));
  NAND2_X1   g06425(.A1(new_n8861_), .A2(new_n8858_), .ZN(new_n8862_));
  AOI21_X1   g06426(.A1(new_n8862_), .A2(new_n8856_), .B(new_n8855_), .ZN(new_n8863_));
  INV_X1     g06427(.I(new_n8850_), .ZN(new_n8864_));
  NOR2_X1    g06428(.A1(new_n8864_), .A2(pi0072), .ZN(new_n8865_));
  NOR3_X1    g06429(.A1(new_n8863_), .A2(new_n5792_), .A3(new_n8865_), .ZN(new_n8866_));
  OAI21_X1   g06430(.A1(new_n8866_), .A2(new_n8854_), .B(pi0075), .ZN(new_n8867_));
  AOI21_X1   g06431(.A1(new_n8378_), .A2(pi0287), .B(pi0072), .ZN(new_n8868_));
  INV_X1     g06432(.I(new_n8868_), .ZN(new_n8869_));
  OAI21_X1   g06433(.A1(new_n8869_), .A2(new_n8864_), .B(new_n3270_), .ZN(new_n8870_));
  NAND2_X1   g06434(.A1(new_n8480_), .A2(pi0044), .ZN(new_n8871_));
  NAND2_X1   g06435(.A1(new_n8478_), .A2(new_n8871_), .ZN(new_n8872_));
  OAI21_X1   g06436(.A1(new_n8474_), .A2(new_n8377_), .B(new_n3025_), .ZN(new_n8873_));
  OAI22_X1   g06437(.A1(new_n8872_), .A2(new_n3025_), .B1(new_n8463_), .B2(new_n8873_), .ZN(new_n8874_));
  AOI21_X1   g06438(.A1(new_n8874_), .A2(pi0228), .B(pi0039), .ZN(new_n8875_));
  AOI21_X1   g06439(.A1(new_n8436_), .A2(new_n8377_), .B(pi0228), .ZN(new_n8876_));
  OAI21_X1   g06440(.A1(new_n8377_), .A2(new_n8443_), .B(new_n8876_), .ZN(new_n8877_));
  AOI21_X1   g06441(.A1(new_n8875_), .A2(new_n8877_), .B(new_n8870_), .ZN(new_n8878_));
  AOI21_X1   g06442(.A1(new_n8851_), .A2(pi0038), .B(pi0087), .ZN(new_n8879_));
  OAI21_X1   g06443(.A1(new_n8864_), .A2(pi0072), .B(new_n8489_), .ZN(new_n8880_));
  NOR2_X1    g06444(.A1(new_n8380_), .A2(new_n8377_), .ZN(new_n8881_));
  OAI21_X1   g06445(.A1(new_n8881_), .A2(new_n8859_), .B(new_n8858_), .ZN(new_n8882_));
  AOI21_X1   g06446(.A1(new_n8882_), .A2(new_n8856_), .B(new_n8855_), .ZN(new_n8883_));
  OAI21_X1   g06447(.A1(new_n8883_), .A2(new_n8880_), .B(new_n8879_), .ZN(new_n8884_));
  NAND2_X1   g06448(.A1(new_n6699_), .A2(new_n2821_), .ZN(new_n8885_));
  AOI21_X1   g06449(.A1(new_n8885_), .A2(pi0039), .B(new_n3458_), .ZN(new_n8886_));
  NOR3_X1    g06450(.A1(new_n8386_), .A2(new_n2458_), .A3(new_n3271_), .ZN(new_n8887_));
  INV_X1     g06451(.I(new_n8887_), .ZN(new_n8888_));
  NAND3_X1   g06452(.A1(new_n8378_), .A2(pi0228), .A3(new_n3270_), .ZN(new_n8889_));
  NAND2_X1   g06453(.A1(new_n8889_), .A2(new_n8440_), .ZN(new_n8890_));
  NAND3_X1   g06454(.A1(new_n8890_), .A2(new_n2627_), .A3(new_n8888_), .ZN(new_n8891_));
  AOI21_X1   g06455(.A1(new_n8891_), .A2(new_n8886_), .B(pi0075), .ZN(new_n8892_));
  OAI21_X1   g06456(.A1(new_n8878_), .A2(new_n8884_), .B(new_n8892_), .ZN(new_n8893_));
  AOI21_X1   g06457(.A1(new_n8893_), .A2(new_n8867_), .B(new_n6648_), .ZN(new_n8894_));
  OAI21_X1   g06458(.A1(new_n8894_), .A2(new_n8853_), .B(new_n8849_), .ZN(po0202));
  INV_X1     g06459(.I(new_n8150_), .ZN(new_n8896_));
  NOR2_X1    g06460(.A1(new_n8265_), .A2(new_n8896_), .ZN(new_n8897_));
  INV_X1     g06461(.I(new_n8897_), .ZN(new_n8898_));
  NOR3_X1    g06462(.A1(new_n8898_), .A2(new_n5389_), .A3(new_n8283_), .ZN(po0203));
  NAND4_X1   g06463(.A1(new_n2478_), .A2(new_n2922_), .A3(new_n2927_), .A4(new_n2482_), .ZN(new_n8900_));
  INV_X1     g06464(.I(pi0104), .ZN(new_n8901_));
  NAND3_X1   g06465(.A1(new_n2501_), .A2(new_n8901_), .A3(new_n2912_), .ZN(new_n8902_));
  NOR4_X1    g06466(.A1(new_n8900_), .A2(pi0071), .A3(new_n8902_), .A4(new_n7409_), .ZN(new_n8903_));
  INV_X1     g06467(.I(pi0083), .ZN(new_n8904_));
  NAND4_X1   g06468(.A1(new_n2911_), .A2(new_n8904_), .A3(new_n2479_), .A4(pi0061), .ZN(new_n8905_));
  NAND2_X1   g06469(.A1(new_n7305_), .A2(new_n6667_), .ZN(new_n8906_));
  NOR4_X1    g06470(.A1(new_n8906_), .A2(new_n7312_), .A3(new_n7300_), .A4(new_n8905_), .ZN(new_n8907_));
  AND3_X2    g06471(.A1(new_n8907_), .A2(new_n8317_), .A3(new_n8903_), .Z(new_n8908_));
  NAND2_X1   g06472(.A1(new_n2979_), .A2(new_n2736_), .ZN(new_n8909_));
  INV_X1     g06473(.I(new_n8909_), .ZN(new_n8910_));
  AOI22_X1   g06474(.A1(new_n8910_), .A2(pi0024), .B1(new_n3179_), .B2(new_n8908_), .ZN(new_n8911_));
  NOR2_X1    g06475(.A1(new_n8911_), .A2(new_n8262_), .ZN(po0204));
  INV_X1     g06476(.I(new_n3082_), .ZN(new_n8913_));
  OAI21_X1   g06477(.A1(new_n2885_), .A2(new_n2884_), .B(new_n6667_), .ZN(new_n8914_));
  NOR2_X1    g06478(.A1(new_n8244_), .A2(new_n7301_), .ZN(new_n8915_));
  NAND2_X1   g06479(.A1(new_n2496_), .A2(new_n8248_), .ZN(new_n8916_));
  INV_X1     g06480(.I(new_n8916_), .ZN(new_n8917_));
  INV_X1     g06481(.I(new_n2940_), .ZN(new_n8918_));
  NOR4_X1    g06482(.A1(new_n8272_), .A2(pi0084), .A3(new_n8901_), .A4(new_n2926_), .ZN(new_n8919_));
  NAND3_X1   g06483(.A1(new_n8919_), .A2(new_n8918_), .A3(new_n2911_), .ZN(new_n8920_));
  NAND2_X1   g06484(.A1(new_n8920_), .A2(new_n7416_), .ZN(new_n8921_));
  NAND4_X1   g06485(.A1(new_n8921_), .A2(new_n2887_), .A3(new_n8915_), .A4(new_n8917_), .ZN(new_n8922_));
  NOR2_X1    g06486(.A1(new_n8922_), .A2(pi0036), .ZN(new_n8923_));
  NOR2_X1    g06487(.A1(new_n8923_), .A2(pi0088), .ZN(new_n8924_));
  NOR2_X1    g06488(.A1(new_n8924_), .A2(new_n8914_), .ZN(new_n8925_));
  NAND2_X1   g06489(.A1(new_n8925_), .A2(new_n8268_), .ZN(new_n8926_));
  NOR2_X1    g06490(.A1(new_n8926_), .A2(new_n3082_), .ZN(new_n8927_));
  AOI21_X1   g06491(.A1(new_n8927_), .A2(new_n5428_), .B(new_n3044_), .ZN(new_n8928_));
  INV_X1     g06492(.I(new_n8922_), .ZN(new_n8929_));
  AOI21_X1   g06493(.A1(new_n8929_), .A2(new_n2920_), .B(pi0088), .ZN(new_n8930_));
  OR3_X2     g06494(.A1(new_n8930_), .A2(new_n2758_), .A3(new_n8914_), .Z(new_n8931_));
  OAI21_X1   g06495(.A1(new_n8931_), .A2(pi0091), .B(new_n6720_), .ZN(new_n8932_));
  NAND3_X1   g06496(.A1(new_n8932_), .A2(new_n5359_), .A3(new_n8253_), .ZN(new_n8933_));
  OAI21_X1   g06497(.A1(new_n8933_), .A2(new_n8913_), .B(new_n8928_), .ZN(new_n8934_));
  OAI21_X1   g06498(.A1(new_n8933_), .A2(new_n6258_), .B(new_n3044_), .ZN(new_n8935_));
  AOI21_X1   g06499(.A1(new_n8934_), .A2(new_n8935_), .B(pi1093), .ZN(new_n8936_));
  NOR2_X1    g06500(.A1(new_n8933_), .A2(new_n6258_), .ZN(new_n8937_));
  NOR2_X1    g06501(.A1(new_n8254_), .A2(new_n6259_), .ZN(new_n8938_));
  INV_X1     g06502(.I(new_n8938_), .ZN(new_n8939_));
  OAI22_X1   g06503(.A1(new_n8252_), .A2(new_n8939_), .B1(new_n5538_), .B2(new_n6870_), .ZN(new_n8940_));
  NOR2_X1    g06504(.A1(new_n8937_), .A2(new_n8940_), .ZN(new_n8941_));
  OR2_X2     g06505(.A1(new_n8934_), .A2(new_n3024_), .Z(new_n8942_));
  NAND2_X1   g06506(.A1(new_n8933_), .A2(new_n6781_), .ZN(new_n8943_));
  AOI21_X1   g06507(.A1(new_n8942_), .A2(new_n8943_), .B(new_n3022_), .ZN(new_n8944_));
  NOR4_X1    g06508(.A1(new_n8944_), .A2(new_n8260_), .A3(new_n8936_), .A4(new_n8941_), .ZN(po0205));
  NOR3_X1    g06509(.A1(new_n3007_), .A2(pi0072), .A3(new_n3179_), .ZN(new_n8946_));
  INV_X1     g06510(.I(new_n8946_), .ZN(new_n8947_));
  NAND4_X1   g06511(.A1(new_n8259_), .A2(new_n2519_), .A3(new_n7750_), .A4(new_n2535_), .ZN(new_n8948_));
  NOR4_X1    g06512(.A1(new_n8948_), .A2(pi0051), .A3(new_n8322_), .A4(new_n8947_), .ZN(po0206));
  NAND2_X1   g06513(.A1(new_n6227_), .A2(new_n6643_), .ZN(new_n8950_));
  NAND2_X1   g06514(.A1(new_n7334_), .A2(pi0074), .ZN(new_n8951_));
  INV_X1     g06515(.I(new_n2505_), .ZN(new_n8952_));
  NOR2_X1    g06516(.A1(new_n8952_), .A2(new_n7409_), .ZN(new_n8953_));
  NAND4_X1   g06517(.A1(new_n2925_), .A2(new_n7297_), .A3(new_n8315_), .A4(new_n2901_), .ZN(new_n8954_));
  NOR4_X1    g06518(.A1(new_n8954_), .A2(pi0068), .A3(pi0073), .A4(new_n7301_), .ZN(new_n8955_));
  INV_X1     g06519(.I(new_n8955_), .ZN(new_n8956_));
  NOR4_X1    g06520(.A1(new_n8956_), .A2(pi0045), .A3(new_n2478_), .A4(new_n8902_), .ZN(new_n8957_));
  NAND4_X1   g06521(.A1(new_n8957_), .A2(new_n2911_), .A3(new_n8918_), .A4(new_n8953_), .ZN(new_n8958_));
  NOR3_X1    g06522(.A1(new_n8958_), .A2(new_n2745_), .A3(new_n7312_), .ZN(new_n8959_));
  INV_X1     g06523(.I(new_n8959_), .ZN(new_n8960_));
  NOR2_X1    g06524(.A1(new_n8960_), .A2(new_n2536_), .ZN(new_n8961_));
  NAND4_X1   g06525(.A1(new_n8961_), .A2(new_n2625_), .A3(new_n2740_), .A4(new_n8946_), .ZN(new_n8962_));
  AOI21_X1   g06526(.A1(new_n8962_), .A2(new_n8951_), .B(new_n8950_), .ZN(po0207));
  NOR2_X1    g06527(.A1(new_n7288_), .A2(new_n2704_), .ZN(new_n8964_));
  AOI21_X1   g06528(.A1(new_n7324_), .A2(new_n2704_), .B(new_n8964_), .ZN(new_n8965_));
  NOR2_X1    g06529(.A1(new_n7276_), .A2(new_n7278_), .ZN(new_n8966_));
  AOI21_X1   g06530(.A1(new_n8966_), .A2(new_n2514_), .B(new_n8965_), .ZN(new_n8967_));
  OAI21_X1   g06531(.A1(new_n7278_), .A2(new_n7293_), .B(new_n8429_), .ZN(new_n8968_));
  NAND3_X1   g06532(.A1(new_n8968_), .A2(new_n8253_), .A3(new_n8967_), .ZN(new_n8969_));
  NOR2_X1    g06533(.A1(new_n2747_), .A2(new_n2526_), .ZN(new_n8970_));
  NAND4_X1   g06534(.A1(new_n8965_), .A2(pi0024), .A3(new_n2985_), .A4(new_n8970_), .ZN(new_n8971_));
  OR2_X2     g06535(.A1(new_n7277_), .A2(new_n8971_), .Z(new_n8972_));
  AOI21_X1   g06536(.A1(new_n8969_), .A2(new_n8972_), .B(pi0100), .ZN(new_n8973_));
  NOR3_X1    g06537(.A1(new_n5501_), .A2(new_n2702_), .A3(new_n5309_), .ZN(new_n8974_));
  NOR2_X1    g06538(.A1(new_n2565_), .A2(new_n2573_), .ZN(new_n8975_));
  OAI21_X1   g06539(.A1(new_n8973_), .A2(new_n8974_), .B(new_n8975_), .ZN(new_n8976_));
  NAND3_X1   g06540(.A1(new_n7338_), .A2(new_n5324_), .A3(new_n7288_), .ZN(new_n8977_));
  AOI21_X1   g06541(.A1(new_n8976_), .A2(new_n8977_), .B(new_n7268_), .ZN(po0208));
  NAND3_X1   g06542(.A1(new_n8261_), .A2(new_n2732_), .A3(new_n2757_), .ZN(new_n8979_));
  NAND3_X1   g06543(.A1(new_n8953_), .A2(new_n2493_), .A3(new_n8243_), .ZN(new_n8980_));
  NOR2_X1    g06544(.A1(new_n8980_), .A2(pi0103), .ZN(new_n8981_));
  NAND2_X1   g06545(.A1(new_n8981_), .A2(new_n2907_), .ZN(new_n8982_));
  NOR2_X1    g06546(.A1(new_n8982_), .A2(new_n5568_), .ZN(new_n8983_));
  INV_X1     g06547(.I(new_n8983_), .ZN(new_n8984_));
  NOR3_X1    g06548(.A1(new_n8979_), .A2(new_n2924_), .A3(new_n8984_), .ZN(po0209));
  NOR2_X1    g06549(.A1(new_n8727_), .A2(pi0072), .ZN(new_n8986_));
  INV_X1     g06550(.I(new_n8986_), .ZN(new_n8987_));
  NOR2_X1    g06551(.A1(new_n8987_), .A2(pi0039), .ZN(new_n8988_));
  INV_X1     g06552(.I(new_n8988_), .ZN(new_n8989_));
  NAND2_X1   g06553(.A1(new_n8810_), .A2(new_n8807_), .ZN(new_n8990_));
  NOR2_X1    g06554(.A1(new_n8990_), .A2(new_n2627_), .ZN(new_n8991_));
  AOI21_X1   g06555(.A1(new_n8516_), .A2(new_n8991_), .B(new_n6643_), .ZN(new_n8992_));
  NOR2_X1    g06556(.A1(new_n8986_), .A2(pi0039), .ZN(new_n8993_));
  NOR2_X1    g06557(.A1(new_n8676_), .A2(new_n8993_), .ZN(new_n8994_));
  INV_X1     g06558(.I(new_n8994_), .ZN(new_n8995_));
  AOI21_X1   g06559(.A1(new_n8995_), .A2(new_n6648_), .B(new_n8990_), .ZN(new_n8996_));
  NOR3_X1    g06560(.A1(new_n8784_), .A2(new_n8523_), .A3(new_n8785_), .ZN(new_n8997_));
  OAI21_X1   g06561(.A1(new_n8677_), .A2(new_n8997_), .B(pi0075), .ZN(new_n8998_));
  NOR3_X1    g06562(.A1(pi0042), .A2(pi0043), .A3(pi0114), .ZN(new_n8999_));
  INV_X1     g06563(.I(new_n8999_), .ZN(new_n9000_));
  NOR2_X1    g06564(.A1(new_n6819_), .A2(new_n8542_), .ZN(new_n9001_));
  INV_X1     g06565(.I(new_n9001_), .ZN(new_n9002_));
  NOR3_X1    g06566(.A1(new_n8551_), .A2(new_n9000_), .A3(new_n9002_), .ZN(new_n9003_));
  AOI21_X1   g06567(.A1(new_n9003_), .A2(new_n2626_), .B(new_n8989_), .ZN(new_n9004_));
  NOR2_X1    g06568(.A1(new_n9004_), .A2(pi0039), .ZN(new_n9005_));
  OAI21_X1   g06569(.A1(new_n9005_), .A2(new_n8998_), .B(new_n6645_), .ZN(new_n9006_));
  AOI21_X1   g06570(.A1(new_n8994_), .A2(new_n3271_), .B(new_n3458_), .ZN(new_n9007_));
  NOR2_X1    g06571(.A1(new_n8787_), .A2(new_n8993_), .ZN(new_n9008_));
  NAND2_X1   g06572(.A1(new_n9008_), .A2(new_n3271_), .ZN(new_n9009_));
  NOR2_X1    g06573(.A1(new_n9000_), .A2(pi0115), .ZN(new_n9010_));
  NAND2_X1   g06574(.A1(new_n9010_), .A2(pi0228), .ZN(new_n9011_));
  NAND2_X1   g06575(.A1(new_n9011_), .A2(new_n8987_), .ZN(new_n9012_));
  AOI21_X1   g06576(.A1(new_n8553_), .A2(new_n5315_), .B(pi0052), .ZN(new_n9013_));
  AOI21_X1   g06577(.A1(new_n8769_), .A2(pi0052), .B(new_n9013_), .ZN(new_n9014_));
  OAI21_X1   g06578(.A1(new_n9014_), .A2(new_n9011_), .B(new_n9012_), .ZN(new_n9015_));
  NAND2_X1   g06579(.A1(new_n9015_), .A2(new_n2627_), .ZN(new_n9016_));
  NAND3_X1   g06580(.A1(new_n9016_), .A2(new_n3270_), .A3(new_n8790_), .ZN(new_n9017_));
  NAND3_X1   g06581(.A1(new_n9017_), .A2(new_n9007_), .A3(new_n9009_), .ZN(new_n9018_));
  NOR2_X1    g06582(.A1(new_n9002_), .A2(new_n9000_), .ZN(new_n9019_));
  AOI21_X1   g06583(.A1(new_n8578_), .A2(new_n9019_), .B(new_n8987_), .ZN(new_n9020_));
  NOR2_X1    g06584(.A1(new_n9020_), .A2(pi0039), .ZN(new_n9021_));
  NOR2_X1    g06585(.A1(new_n9021_), .A2(new_n8789_), .ZN(new_n9022_));
  NAND2_X1   g06586(.A1(new_n8995_), .A2(pi0038), .ZN(new_n9023_));
  OAI22_X1   g06587(.A1(new_n9022_), .A2(new_n8667_), .B1(new_n9008_), .B2(new_n9023_), .ZN(new_n9024_));
  NOR2_X1    g06588(.A1(new_n9010_), .A2(new_n8986_), .ZN(new_n9025_));
  INV_X1     g06589(.I(new_n9025_), .ZN(new_n9026_));
  NOR2_X1    g06590(.A1(new_n8591_), .A2(pi0052), .ZN(new_n9027_));
  AOI21_X1   g06591(.A1(new_n8605_), .A2(pi0052), .B(new_n9027_), .ZN(new_n9028_));
  INV_X1     g06592(.I(new_n9028_), .ZN(new_n9029_));
  AOI21_X1   g06593(.A1(new_n9029_), .A2(new_n9010_), .B(pi0228), .ZN(new_n9030_));
  AOI21_X1   g06594(.A1(new_n9030_), .A2(new_n9026_), .B(pi0039), .ZN(new_n9031_));
  NOR2_X1    g06595(.A1(new_n9025_), .A2(new_n2458_), .ZN(new_n9032_));
  NOR2_X1    g06596(.A1(new_n8752_), .A2(new_n8727_), .ZN(new_n9033_));
  NOR2_X1    g06597(.A1(new_n8611_), .A2(pi0052), .ZN(new_n9034_));
  OAI21_X1   g06598(.A1(new_n9033_), .A2(new_n9034_), .B(new_n8541_), .ZN(new_n9035_));
  INV_X1     g06599(.I(new_n9035_), .ZN(new_n9036_));
  NAND2_X1   g06600(.A1(new_n8629_), .A2(new_n8727_), .ZN(new_n9037_));
  NAND3_X1   g06601(.A1(new_n9037_), .A2(new_n8587_), .A3(new_n3026_), .ZN(new_n9038_));
  AOI21_X1   g06602(.A1(new_n8624_), .A2(pi0052), .B(new_n9038_), .ZN(new_n9039_));
  NOR2_X1    g06603(.A1(new_n9036_), .A2(new_n9039_), .ZN(new_n9040_));
  OAI21_X1   g06604(.A1(new_n9040_), .A2(new_n9000_), .B(new_n9032_), .ZN(new_n9041_));
  AND2_X2    g06605(.A1(new_n9041_), .A2(new_n9031_), .Z(new_n9042_));
  INV_X1     g06606(.I(new_n9042_), .ZN(new_n9043_));
  AOI21_X1   g06607(.A1(new_n9043_), .A2(new_n8799_), .B(new_n3271_), .ZN(new_n9044_));
  OAI21_X1   g06608(.A1(new_n9044_), .A2(new_n9024_), .B(new_n3458_), .ZN(new_n9045_));
  NAND3_X1   g06609(.A1(new_n9045_), .A2(new_n8524_), .A3(new_n9018_), .ZN(new_n9046_));
  NAND3_X1   g06610(.A1(new_n9016_), .A2(new_n3270_), .A3(new_n8677_), .ZN(new_n9047_));
  AOI21_X1   g06611(.A1(new_n9047_), .A2(new_n9007_), .B(new_n8524_), .ZN(new_n9048_));
  INV_X1     g06612(.I(new_n8690_), .ZN(new_n9049_));
  OAI21_X1   g06613(.A1(new_n2821_), .A2(pi0232), .B(pi0299), .ZN(new_n9050_));
  OAI21_X1   g06614(.A1(new_n9049_), .A2(new_n9050_), .B(pi0039), .ZN(new_n9051_));
  NAND2_X1   g06615(.A1(new_n9043_), .A2(new_n9051_), .ZN(new_n9052_));
  OAI21_X1   g06616(.A1(new_n9021_), .A2(new_n8676_), .B(new_n8489_), .ZN(new_n9053_));
  NAND2_X1   g06617(.A1(new_n9053_), .A2(new_n9023_), .ZN(new_n9054_));
  AOI21_X1   g06618(.A1(new_n9052_), .A2(new_n3270_), .B(new_n9054_), .ZN(new_n9055_));
  OAI21_X1   g06619(.A1(new_n9055_), .A2(pi0087), .B(new_n9048_), .ZN(new_n9056_));
  AOI21_X1   g06620(.A1(new_n9046_), .A2(new_n9056_), .B(pi0075), .ZN(new_n9057_));
  OAI21_X1   g06621(.A1(new_n9057_), .A2(new_n9006_), .B(new_n8996_), .ZN(new_n9058_));
  OAI21_X1   g06622(.A1(new_n9008_), .A2(new_n3265_), .B(new_n3458_), .ZN(new_n9059_));
  OAI21_X1   g06623(.A1(new_n9020_), .A2(pi0039), .B(new_n8788_), .ZN(new_n9060_));
  AOI21_X1   g06624(.A1(new_n9060_), .A2(new_n8489_), .B(new_n9059_), .ZN(new_n9061_));
  NAND2_X1   g06625(.A1(new_n9043_), .A2(new_n8823_), .ZN(new_n9062_));
  NAND2_X1   g06626(.A1(new_n9062_), .A2(new_n3270_), .ZN(new_n9063_));
  NAND2_X1   g06627(.A1(new_n9063_), .A2(new_n9061_), .ZN(new_n9064_));
  INV_X1     g06628(.I(new_n9009_), .ZN(new_n9065_));
  AND3_X2    g06629(.A1(new_n9016_), .A2(new_n3270_), .A3(new_n8788_), .Z(new_n9066_));
  OAI21_X1   g06630(.A1(new_n9066_), .A2(new_n9065_), .B(pi0087), .ZN(new_n9067_));
  NAND3_X1   g06631(.A1(new_n9064_), .A2(new_n3465_), .A3(new_n9067_), .ZN(new_n9068_));
  AOI21_X1   g06632(.A1(new_n9008_), .A2(new_n5792_), .B(new_n3465_), .ZN(new_n9069_));
  NOR2_X1    g06633(.A1(new_n9003_), .A2(new_n8987_), .ZN(new_n9070_));
  NOR2_X1    g06634(.A1(new_n9070_), .A2(pi0039), .ZN(new_n9071_));
  NAND2_X1   g06635(.A1(new_n8788_), .A2(new_n2626_), .ZN(new_n9072_));
  OAI21_X1   g06636(.A1(new_n9071_), .A2(new_n9072_), .B(new_n9069_), .ZN(new_n9073_));
  NAND4_X1   g06637(.A1(new_n9068_), .A2(new_n6645_), .A3(new_n8524_), .A4(new_n9073_), .ZN(new_n9074_));
  OR2_X2     g06638(.A1(new_n9004_), .A2(new_n3465_), .Z(new_n9075_));
  NOR2_X1    g06639(.A1(new_n8989_), .A2(new_n3265_), .ZN(new_n9076_));
  NAND2_X1   g06640(.A1(new_n9043_), .A2(new_n2702_), .ZN(new_n9077_));
  NAND2_X1   g06641(.A1(new_n9020_), .A2(pi0100), .ZN(new_n9078_));
  AOI21_X1   g06642(.A1(new_n9077_), .A2(new_n9078_), .B(new_n2573_), .ZN(new_n9079_));
  OAI21_X1   g06643(.A1(new_n9079_), .A2(new_n9076_), .B(new_n3458_), .ZN(new_n9080_));
  NOR2_X1    g06644(.A1(new_n8896_), .A2(pi0100), .ZN(new_n9081_));
  NOR2_X1    g06645(.A1(new_n9081_), .A2(new_n3458_), .ZN(new_n9082_));
  INV_X1     g06646(.I(new_n9082_), .ZN(new_n9083_));
  AOI21_X1   g06647(.A1(pi0100), .A2(new_n8989_), .B(new_n9083_), .ZN(new_n9084_));
  OAI21_X1   g06648(.A1(new_n9015_), .A2(pi0038), .B(new_n2702_), .ZN(new_n9085_));
  OAI21_X1   g06649(.A1(new_n9085_), .A2(new_n9076_), .B(new_n9084_), .ZN(new_n9086_));
  NAND3_X1   g06650(.A1(new_n9080_), .A2(new_n3465_), .A3(new_n9086_), .ZN(new_n9087_));
  AOI21_X1   g06651(.A1(new_n9087_), .A2(new_n9075_), .B(new_n6648_), .ZN(new_n9088_));
  OAI21_X1   g06652(.A1(new_n8988_), .A2(new_n6645_), .B(new_n8523_), .ZN(new_n9089_));
  OAI21_X1   g06653(.A1(new_n9088_), .A2(new_n9089_), .B(new_n9074_), .ZN(new_n9090_));
  NAND3_X1   g06654(.A1(new_n9008_), .A2(new_n6648_), .A3(new_n8524_), .ZN(new_n9091_));
  NAND2_X1   g06655(.A1(new_n9091_), .A2(new_n6643_), .ZN(new_n9092_));
  AOI21_X1   g06656(.A1(new_n9090_), .A2(new_n8990_), .B(new_n9092_), .ZN(new_n9093_));
  AOI22_X1   g06657(.A1(new_n9093_), .A2(new_n9058_), .B1(new_n8989_), .B2(new_n8992_), .ZN(po0210));
  INV_X1     g06658(.I(new_n3447_), .ZN(new_n9095_));
  NOR3_X1    g06659(.A1(new_n5386_), .A2(new_n5387_), .A3(pi0979), .ZN(new_n9096_));
  AOI21_X1   g06660(.A1(new_n9096_), .A2(new_n8282_), .B(new_n2627_), .ZN(new_n9097_));
  INV_X1     g06661(.I(new_n9097_), .ZN(new_n9098_));
  NAND2_X1   g06662(.A1(new_n8280_), .A2(new_n9098_), .ZN(new_n9099_));
  NOR2_X1    g06663(.A1(new_n7571_), .A2(pi0058), .ZN(new_n9100_));
  INV_X1     g06664(.I(new_n9100_), .ZN(new_n9101_));
  NOR4_X1    g06665(.A1(new_n9101_), .A2(new_n2793_), .A3(pi0060), .A4(new_n2727_), .ZN(new_n9102_));
  NAND4_X1   g06666(.A1(new_n9102_), .A2(pi0024), .A3(new_n2627_), .A4(new_n8253_), .ZN(new_n9103_));
  AOI21_X1   g06667(.A1(new_n9103_), .A2(new_n9095_), .B(new_n9099_), .ZN(po0211));
  NAND2_X1   g06668(.A1(new_n8266_), .A2(new_n2626_), .ZN(new_n9105_));
  NOR2_X1    g06669(.A1(new_n9105_), .A2(new_n2606_), .ZN(new_n9106_));
  NAND2_X1   g06670(.A1(new_n9106_), .A2(pi0054), .ZN(new_n9107_));
  NOR2_X1    g06671(.A1(pi0060), .A2(pi0085), .ZN(new_n9108_));
  NAND4_X1   g06672(.A1(new_n2914_), .A2(pi0106), .A3(new_n7296_), .A4(new_n9108_), .ZN(new_n9109_));
  NAND2_X1   g06673(.A1(new_n8953_), .A2(new_n7302_), .ZN(new_n9110_));
  NOR4_X1    g06674(.A1(new_n9110_), .A2(new_n8900_), .A3(new_n8954_), .A4(new_n9109_), .ZN(new_n9111_));
  NOR2_X1    g06675(.A1(new_n7573_), .A2(new_n7293_), .ZN(new_n9112_));
  NAND2_X1   g06676(.A1(new_n9112_), .A2(new_n9111_), .ZN(new_n9113_));
  NAND2_X1   g06677(.A1(new_n2740_), .A2(new_n3179_), .ZN(new_n9114_));
  NOR2_X1    g06678(.A1(new_n7332_), .A2(new_n9114_), .ZN(new_n9115_));
  INV_X1     g06679(.I(new_n9115_), .ZN(new_n9116_));
  NOR3_X1    g06680(.A1(new_n9113_), .A2(new_n2745_), .A3(new_n9116_), .ZN(new_n9117_));
  NAND3_X1   g06681(.A1(new_n9117_), .A2(new_n5499_), .A3(new_n2660_), .ZN(new_n9118_));
  AOI21_X1   g06682(.A1(new_n9107_), .A2(new_n9118_), .B(new_n7266_), .ZN(po0212));
  NOR3_X1    g06683(.A1(new_n7409_), .A2(new_n2913_), .A3(new_n2933_), .ZN(new_n9120_));
  NAND3_X1   g06684(.A1(new_n8955_), .A2(new_n2934_), .A3(new_n9120_), .ZN(new_n9121_));
  INV_X1     g06685(.I(new_n9121_), .ZN(new_n9122_));
  NOR4_X1    g06686(.A1(new_n2612_), .A2(new_n7413_), .A3(new_n2536_), .A4(new_n7717_), .ZN(new_n9123_));
  AOI21_X1   g06687(.A1(new_n9123_), .A2(new_n9122_), .B(pi0055), .ZN(new_n9124_));
  NAND2_X1   g06688(.A1(new_n9106_), .A2(new_n5499_), .ZN(new_n9125_));
  INV_X1     g06689(.I(new_n9125_), .ZN(new_n9126_));
  AOI21_X1   g06690(.A1(new_n9126_), .A2(new_n2625_), .B(new_n2602_), .ZN(new_n9127_));
  NOR4_X1    g06691(.A1(new_n9127_), .A2(new_n2471_), .A3(new_n3425_), .A4(new_n9124_), .ZN(po0213));
  NAND2_X1   g06692(.A1(new_n3471_), .A2(pi0056), .ZN(new_n9129_));
  NAND2_X1   g06693(.A1(new_n8188_), .A2(pi0055), .ZN(new_n9130_));
  NOR3_X1    g06694(.A1(new_n5356_), .A2(new_n7456_), .A3(new_n2577_), .ZN(new_n9131_));
  OAI21_X1   g06695(.A1(new_n9131_), .A2(new_n3284_), .B(new_n3291_), .ZN(new_n9132_));
  AOI21_X1   g06696(.A1(new_n9129_), .A2(new_n9130_), .B(new_n9132_), .ZN(po0214));
  NOR3_X1    g06697(.A1(new_n9125_), .A2(pi0074), .A3(new_n5476_), .ZN(new_n9134_));
  NAND2_X1   g06698(.A1(new_n9134_), .A2(pi0057), .ZN(new_n9135_));
  NOR3_X1    g06699(.A1(new_n5612_), .A2(new_n7456_), .A3(new_n2577_), .ZN(new_n9136_));
  NOR2_X1    g06700(.A1(new_n3471_), .A2(pi0056), .ZN(new_n9137_));
  INV_X1     g06701(.I(new_n9137_), .ZN(new_n9138_));
  OAI21_X1   g06702(.A1(new_n9138_), .A2(pi0924), .B(new_n9129_), .ZN(new_n9139_));
  NAND3_X1   g06703(.A1(new_n9136_), .A2(new_n2582_), .A3(new_n9139_), .ZN(new_n9140_));
  AOI21_X1   g06704(.A1(new_n9135_), .A2(new_n9140_), .B(pi0059), .ZN(po0215));
  INV_X1     g06705(.I(new_n8970_), .ZN(new_n9142_));
  NOR3_X1    g06706(.A1(new_n8260_), .A2(pi0093), .A3(new_n9142_), .ZN(new_n9143_));
  AND3_X2    g06707(.A1(new_n6662_), .A2(pi0090), .A3(new_n9143_), .Z(po0216));
  NAND2_X1   g06708(.A1(new_n9134_), .A2(pi0059), .ZN(new_n9145_));
  NAND4_X1   g06709(.A1(new_n9136_), .A2(new_n2469_), .A3(pi0924), .A4(new_n9137_), .ZN(new_n9146_));
  AOI21_X1   g06710(.A1(new_n9145_), .A2(new_n9146_), .B(pi0057), .ZN(po0217));
  INV_X1     g06711(.I(pi1001), .ZN(new_n9148_));
  NOR2_X1    g06712(.A1(new_n2530_), .A2(pi0287), .ZN(new_n9149_));
  NOR3_X1    g06713(.A1(new_n5388_), .A2(new_n2627_), .A3(pi0979), .ZN(new_n9150_));
  NAND4_X1   g06714(.A1(new_n9149_), .A2(new_n2704_), .A3(new_n9148_), .A4(new_n9150_), .ZN(new_n9151_));
  NOR3_X1    g06715(.A1(new_n7573_), .A2(pi0039), .A3(new_n7293_), .ZN(new_n9152_));
  NAND4_X1   g06716(.A1(new_n9152_), .A2(pi0024), .A3(new_n2789_), .A4(new_n8253_), .ZN(new_n9153_));
  AOI21_X1   g06717(.A1(new_n9153_), .A2(new_n9151_), .B(new_n8281_), .ZN(po0218));
  NAND2_X1   g06718(.A1(new_n8908_), .A2(pi0841), .ZN(new_n9155_));
  NAND3_X1   g06719(.A1(new_n9112_), .A2(new_n7278_), .A3(new_n2789_), .ZN(new_n9156_));
  AOI21_X1   g06720(.A1(new_n9156_), .A2(new_n9155_), .B(new_n8262_), .ZN(po0219));
  NAND2_X1   g06721(.A1(new_n8190_), .A2(pi0057), .ZN(new_n9158_));
  NAND3_X1   g06722(.A1(new_n9131_), .A2(new_n2582_), .A3(new_n9137_), .ZN(new_n9159_));
  AOI21_X1   g06723(.A1(new_n9158_), .A2(new_n9159_), .B(pi0059), .ZN(po0220));
  NOR4_X1    g06724(.A1(new_n7425_), .A2(new_n2895_), .A3(pi0107), .A4(new_n7312_), .ZN(new_n9161_));
  AOI22_X1   g06725(.A1(new_n8910_), .A2(new_n7278_), .B1(pi0999), .B2(new_n9161_), .ZN(new_n9162_));
  NOR2_X1    g06726(.A1(new_n9162_), .A2(new_n8262_), .ZN(po0221));
  NAND3_X1   g06727(.A1(new_n2891_), .A2(new_n2895_), .A3(pi0107), .ZN(new_n9164_));
  NAND2_X1   g06728(.A1(new_n9164_), .A2(new_n2495_), .ZN(new_n9165_));
  NAND4_X1   g06729(.A1(new_n8277_), .A2(new_n9165_), .A3(pi0841), .A4(new_n7414_), .ZN(new_n9166_));
  NAND4_X1   g06730(.A1(new_n7424_), .A2(new_n2895_), .A3(pi0107), .A4(new_n3179_), .ZN(new_n9167_));
  AOI21_X1   g06731(.A1(new_n9166_), .A2(new_n9167_), .B(new_n8979_), .ZN(po0222));
  NAND3_X1   g06732(.A1(new_n8293_), .A2(new_n8300_), .A3(new_n8280_), .ZN(new_n9169_));
  NOR4_X1    g06733(.A1(new_n9169_), .A2(new_n2627_), .A3(new_n8297_), .A4(pi1082), .ZN(po0223));
  NOR2_X1    g06734(.A1(new_n8525_), .A2(pi0299), .ZN(new_n9171_));
  INV_X1     g06735(.I(new_n9171_), .ZN(new_n9172_));
  NOR2_X1    g06736(.A1(new_n2608_), .A2(new_n3271_), .ZN(new_n9173_));
  INV_X1     g06737(.I(new_n9173_), .ZN(new_n9174_));
  NOR4_X1    g06738(.A1(new_n7717_), .A2(new_n5590_), .A3(new_n8952_), .A4(new_n2536_), .ZN(new_n9175_));
  INV_X1     g06739(.I(new_n9175_), .ZN(new_n9176_));
  NOR2_X1    g06740(.A1(new_n2868_), .A2(new_n2500_), .ZN(new_n9177_));
  INV_X1     g06741(.I(new_n9177_), .ZN(new_n9178_));
  NOR3_X1    g06742(.A1(new_n9178_), .A2(new_n9176_), .A3(pi0102), .ZN(new_n9179_));
  INV_X1     g06743(.I(new_n9179_), .ZN(new_n9180_));
  NOR4_X1    g06744(.A1(new_n9180_), .A2(new_n7599_), .A3(new_n9172_), .A4(new_n9174_), .ZN(new_n9181_));
  OAI21_X1   g06745(.A1(new_n9181_), .A2(pi0219), .B(new_n6643_), .ZN(new_n9182_));
  INV_X1     g06746(.I(new_n8691_), .ZN(new_n9183_));
  NOR2_X1    g06747(.A1(new_n9180_), .A2(new_n2612_), .ZN(new_n9184_));
  AOI21_X1   g06748(.A1(new_n9184_), .A2(new_n9183_), .B(new_n8807_), .ZN(new_n9185_));
  NOR2_X1    g06749(.A1(new_n9182_), .A2(new_n9185_), .ZN(po0224));
  NAND2_X1   g06750(.A1(new_n8981_), .A2(pi0083), .ZN(new_n9187_));
  NOR4_X1    g06751(.A1(new_n8260_), .A2(new_n2492_), .A3(new_n9176_), .A4(new_n9187_), .ZN(po0225));
  NOR2_X1    g06752(.A1(new_n6809_), .A2(new_n5541_), .ZN(new_n9189_));
  NOR3_X1    g06753(.A1(new_n8304_), .A2(new_n2614_), .A3(pi0221), .ZN(new_n9190_));
  NOR2_X1    g06754(.A1(new_n5541_), .A2(new_n5451_), .ZN(new_n9191_));
  NOR2_X1    g06755(.A1(new_n3347_), .A2(new_n3336_), .ZN(new_n9192_));
  AOI22_X1   g06756(.A1(new_n9189_), .A2(new_n9190_), .B1(new_n9191_), .B2(new_n9192_), .ZN(new_n9193_));
  NOR2_X1    g06757(.A1(new_n9193_), .A2(new_n8898_), .ZN(po0226));
  NOR2_X1    g06758(.A1(new_n2919_), .A2(pi0083), .ZN(new_n9195_));
  NAND4_X1   g06759(.A1(new_n9195_), .A2(pi0069), .A3(new_n2901_), .A4(new_n2925_), .ZN(new_n9196_));
  NAND2_X1   g06760(.A1(new_n9196_), .A2(new_n2962_), .ZN(new_n9197_));
  NAND4_X1   g06761(.A1(new_n9197_), .A2(new_n5590_), .A3(new_n2828_), .A4(new_n5567_), .ZN(new_n9198_));
  NOR2_X1    g06762(.A1(new_n8246_), .A2(new_n6668_), .ZN(new_n9199_));
  NAND4_X1   g06763(.A1(new_n9199_), .A2(pi0071), .A3(pi0314), .A4(new_n2827_), .ZN(new_n9200_));
  AOI21_X1   g06764(.A1(new_n9198_), .A2(new_n9200_), .B(new_n8979_), .ZN(po0227));
  NOR2_X1    g06765(.A1(new_n2526_), .A2(pi0039), .ZN(new_n9202_));
  NOR3_X1    g06766(.A1(new_n2813_), .A2(new_n2835_), .A3(new_n2528_), .ZN(new_n9203_));
  NAND3_X1   g06767(.A1(new_n9203_), .A2(pi0024), .A3(new_n9202_), .ZN(new_n9204_));
  INV_X1     g06768(.I(pi0589), .ZN(new_n9205_));
  NOR2_X1    g06769(.A1(new_n2709_), .A2(new_n9205_), .ZN(new_n9206_));
  NOR3_X1    g06770(.A1(new_n6809_), .A2(new_n3304_), .A3(new_n8304_), .ZN(new_n9207_));
  NOR2_X1    g06771(.A1(new_n5451_), .A2(new_n3338_), .ZN(new_n9208_));
  NOR2_X1    g06772(.A1(new_n2672_), .A2(new_n9205_), .ZN(new_n9209_));
  AOI22_X1   g06773(.A1(new_n9207_), .A2(new_n9206_), .B1(new_n9208_), .B2(new_n9209_), .ZN(new_n9210_));
  NOR2_X1    g06774(.A1(new_n3086_), .A2(new_n5534_), .ZN(new_n9211_));
  NOR2_X1    g06775(.A1(new_n9211_), .A2(pi0593), .ZN(new_n9212_));
  NAND3_X1   g06776(.A1(new_n9212_), .A2(pi0835), .A3(new_n5391_), .ZN(new_n9213_));
  OAI21_X1   g06777(.A1(new_n9210_), .A2(new_n9213_), .B(new_n8282_), .ZN(new_n9214_));
  NAND2_X1   g06778(.A1(new_n9214_), .A2(new_n3447_), .ZN(new_n9215_));
  AOI21_X1   g06779(.A1(new_n9215_), .A2(new_n9204_), .B(new_n8281_), .ZN(po0228));
  NOR2_X1    g06780(.A1(new_n9183_), .A2(new_n8531_), .ZN(new_n9217_));
  NOR2_X1    g06781(.A1(new_n8510_), .A2(pi0219), .ZN(new_n9218_));
  INV_X1     g06782(.I(new_n9218_), .ZN(new_n9219_));
  NOR2_X1    g06783(.A1(new_n9219_), .A2(new_n2628_), .ZN(new_n9220_));
  NOR2_X1    g06784(.A1(new_n9220_), .A2(new_n9217_), .ZN(new_n9221_));
  NOR3_X1    g06785(.A1(new_n5569_), .A2(new_n2543_), .A3(new_n8916_), .ZN(new_n9222_));
  NAND4_X1   g06786(.A1(new_n9222_), .A2(new_n8915_), .A3(new_n9175_), .A4(new_n9221_), .ZN(new_n9223_));
  NAND4_X1   g06787(.A1(new_n9222_), .A2(new_n2495_), .A3(new_n2493_), .A4(new_n2907_), .ZN(new_n9224_));
  AOI21_X1   g06788(.A1(new_n9224_), .A2(new_n2500_), .B(new_n9221_), .ZN(new_n9225_));
  NOR2_X1    g06789(.A1(new_n7312_), .A2(pi0050), .ZN(new_n9226_));
  INV_X1     g06790(.I(new_n9226_), .ZN(new_n9227_));
  NOR2_X1    g06791(.A1(new_n5583_), .A2(new_n9227_), .ZN(new_n9228_));
  NAND4_X1   g06792(.A1(new_n9225_), .A2(pi0314), .A3(new_n8253_), .A4(new_n9228_), .ZN(new_n9229_));
  AOI21_X1   g06793(.A1(new_n9229_), .A2(new_n9223_), .B(new_n8260_), .ZN(po0229));
  NAND3_X1   g06794(.A1(new_n9191_), .A2(new_n2631_), .A3(new_n6806_), .ZN(new_n9231_));
  NAND2_X1   g06795(.A1(new_n9189_), .A2(new_n6810_), .ZN(new_n9232_));
  AND3_X2    g06796(.A1(new_n9232_), .A2(new_n9231_), .A3(pi0039), .Z(new_n9233_));
  INV_X1     g06797(.I(new_n2885_), .ZN(new_n9234_));
  NAND2_X1   g06798(.A1(new_n2750_), .A2(pi0024), .ZN(new_n9235_));
  NAND4_X1   g06799(.A1(new_n8251_), .A2(new_n7682_), .A3(pi0088), .A4(new_n5534_), .ZN(new_n9236_));
  OAI22_X1   g06800(.A1(new_n9235_), .A2(new_n2821_), .B1(new_n9234_), .B2(new_n9236_), .ZN(new_n9237_));
  AOI21_X1   g06801(.A1(new_n9237_), .A2(new_n2535_), .B(pi0039), .ZN(new_n9238_));
  NOR3_X1    g06802(.A1(new_n9238_), .A2(new_n8281_), .A3(new_n9233_), .ZN(po0230));
  AOI21_X1   g06803(.A1(new_n9189_), .A2(new_n7508_), .B(new_n2628_), .ZN(new_n9240_));
  NOR3_X1    g06804(.A1(new_n5541_), .A2(new_n5451_), .A3(new_n7525_), .ZN(new_n9241_));
  NOR2_X1    g06805(.A1(new_n9241_), .A2(pi0299), .ZN(new_n9242_));
  NOR2_X1    g06806(.A1(new_n9240_), .A2(new_n9242_), .ZN(new_n9243_));
  NAND2_X1   g06807(.A1(new_n9243_), .A2(pi0039), .ZN(new_n9244_));
  NOR2_X1    g06808(.A1(new_n7464_), .A2(new_n8254_), .ZN(new_n9245_));
  NAND4_X1   g06809(.A1(new_n9245_), .A2(new_n2627_), .A3(new_n5590_), .A4(pi1050), .ZN(new_n9246_));
  AOI21_X1   g06810(.A1(new_n9244_), .A2(new_n9246_), .B(new_n8281_), .ZN(po0231));
  NOR3_X1    g06811(.A1(new_n6259_), .A2(pi0096), .A3(pi1093), .ZN(new_n9248_));
  NOR3_X1    g06812(.A1(new_n3436_), .A2(new_n6648_), .A3(new_n9248_), .ZN(new_n9249_));
  AOI21_X1   g06813(.A1(new_n5350_), .A2(new_n2742_), .B(new_n2998_), .ZN(new_n9250_));
  NOR2_X1    g06814(.A1(po0840), .A2(new_n9250_), .ZN(new_n9251_));
  OAI21_X1   g06815(.A1(new_n6723_), .A2(new_n2766_), .B(new_n2742_), .ZN(new_n9252_));
  NAND4_X1   g06816(.A1(new_n6660_), .A2(new_n9249_), .A3(new_n9252_), .A4(new_n9251_), .ZN(new_n9253_));
  NAND2_X1   g06817(.A1(new_n9126_), .A2(pi0074), .ZN(new_n9254_));
  AOI21_X1   g06818(.A1(new_n9254_), .A2(new_n9253_), .B(po1038), .ZN(po0232));
  AOI21_X1   g06819(.A1(new_n8266_), .A2(new_n2626_), .B(new_n3465_), .ZN(new_n9256_));
  NAND3_X1   g06820(.A1(new_n9252_), .A2(new_n5532_), .A3(new_n3080_), .ZN(new_n9257_));
  NAND2_X1   g06821(.A1(new_n3041_), .A2(pi0096), .ZN(new_n9258_));
  AOI21_X1   g06822(.A1(new_n9257_), .A2(new_n9258_), .B(new_n2659_), .ZN(new_n9259_));
  AOI21_X1   g06823(.A1(new_n9259_), .A2(new_n6728_), .B(pi0075), .ZN(new_n9260_));
  NOR3_X1    g06824(.A1(new_n9260_), .A2(new_n7268_), .A3(new_n9256_), .ZN(po0233));
  AOI21_X1   g06825(.A1(new_n7308_), .A2(new_n2514_), .B(new_n8254_), .ZN(new_n9262_));
  NAND2_X1   g06826(.A1(new_n8429_), .A2(new_n7293_), .ZN(new_n9263_));
  NAND2_X1   g06827(.A1(new_n9263_), .A2(new_n9262_), .ZN(new_n9264_));
  NAND2_X1   g06828(.A1(new_n9264_), .A2(new_n2704_), .ZN(new_n9265_));
  NAND2_X1   g06829(.A1(new_n7307_), .A2(new_n8268_), .ZN(new_n9266_));
  NAND2_X1   g06830(.A1(new_n9266_), .A2(pi0252), .ZN(new_n9267_));
  AOI21_X1   g06831(.A1(new_n9265_), .A2(new_n9267_), .B(new_n3084_), .ZN(new_n9268_));
  INV_X1     g06832(.I(new_n9264_), .ZN(new_n9269_));
  NOR2_X1    g06833(.A1(new_n9269_), .A2(new_n3083_), .ZN(new_n9270_));
  OAI21_X1   g06834(.A1(new_n9268_), .A2(new_n9270_), .B(new_n3041_), .ZN(new_n9271_));
  NAND2_X1   g06835(.A1(new_n9264_), .A2(pi1093), .ZN(new_n9272_));
  NAND2_X1   g06836(.A1(new_n9272_), .A2(new_n3026_), .ZN(new_n9273_));
  NOR2_X1    g06837(.A1(new_n9268_), .A2(new_n9270_), .ZN(new_n9274_));
  INV_X1     g06838(.I(new_n2526_), .ZN(new_n9275_));
  NAND2_X1   g06839(.A1(new_n8430_), .A2(new_n9275_), .ZN(new_n9276_));
  OAI21_X1   g06840(.A1(new_n9276_), .A2(pi0252), .B(new_n3083_), .ZN(new_n9277_));
  OAI21_X1   g06841(.A1(new_n3083_), .A2(new_n9269_), .B(new_n9277_), .ZN(new_n9278_));
  INV_X1     g06842(.I(new_n9278_), .ZN(new_n9279_));
  OAI22_X1   g06843(.A1(new_n9279_), .A2(new_n6257_), .B1(new_n9274_), .B2(new_n6714_), .ZN(new_n9280_));
  OAI21_X1   g06844(.A1(new_n9280_), .A2(new_n3026_), .B(new_n9273_), .ZN(new_n9281_));
  NAND2_X1   g06845(.A1(new_n9281_), .A2(new_n9271_), .ZN(new_n9282_));
  NOR2_X1    g06846(.A1(new_n9266_), .A2(new_n5323_), .ZN(new_n9283_));
  OAI21_X1   g06847(.A1(new_n3026_), .A2(new_n8200_), .B(new_n9283_), .ZN(new_n9284_));
  OAI21_X1   g06848(.A1(new_n9282_), .A2(po1057), .B(new_n9284_), .ZN(new_n9285_));
  NOR2_X1    g06849(.A1(new_n9285_), .A2(new_n2709_), .ZN(new_n9286_));
  AND3_X2    g06850(.A1(po1057), .A2(new_n3016_), .A3(new_n7287_), .Z(new_n9287_));
  NAND2_X1   g06851(.A1(new_n3016_), .A2(new_n3041_), .ZN(new_n9288_));
  OAI21_X1   g06852(.A1(new_n9279_), .A2(new_n9288_), .B(new_n9272_), .ZN(new_n9289_));
  NOR2_X1    g06853(.A1(new_n9271_), .A2(new_n3016_), .ZN(new_n9290_));
  NOR2_X1    g06854(.A1(new_n9289_), .A2(new_n9290_), .ZN(new_n9291_));
  AOI21_X1   g06855(.A1(new_n9291_), .A2(new_n5323_), .B(new_n9283_), .ZN(new_n9292_));
  NOR3_X1    g06856(.A1(new_n9292_), .A2(new_n3025_), .A3(new_n9287_), .ZN(new_n9293_));
  AOI21_X1   g06857(.A1(pi0137), .A2(new_n6257_), .B(new_n3084_), .ZN(new_n9294_));
  NOR2_X1    g06858(.A1(new_n9266_), .A2(new_n9294_), .ZN(new_n9295_));
  OAI21_X1   g06859(.A1(new_n9295_), .A2(new_n5323_), .B(new_n3025_), .ZN(new_n9296_));
  NOR2_X1    g06860(.A1(new_n9280_), .A2(new_n3016_), .ZN(new_n9297_));
  AOI22_X1   g06861(.A1(new_n9297_), .A2(new_n9271_), .B1(new_n3016_), .B2(new_n9279_), .ZN(new_n9298_));
  AOI21_X1   g06862(.A1(new_n9298_), .A2(new_n5323_), .B(new_n9296_), .ZN(new_n9299_));
  NOR2_X1    g06863(.A1(new_n9299_), .A2(new_n9293_), .ZN(new_n9300_));
  AOI21_X1   g06864(.A1(new_n9300_), .A2(new_n2709_), .B(new_n9286_), .ZN(new_n9301_));
  NOR2_X1    g06865(.A1(new_n9301_), .A2(new_n2628_), .ZN(new_n9302_));
  NOR2_X1    g06866(.A1(new_n9285_), .A2(new_n2672_), .ZN(new_n9303_));
  AOI21_X1   g06867(.A1(new_n9300_), .A2(new_n2672_), .B(new_n9303_), .ZN(new_n9304_));
  NOR2_X1    g06868(.A1(new_n9304_), .A2(pi0299), .ZN(new_n9305_));
  OAI21_X1   g06869(.A1(new_n9302_), .A2(new_n9305_), .B(new_n5666_), .ZN(new_n9306_));
  NOR2_X1    g06870(.A1(new_n2670_), .A2(new_n5437_), .ZN(new_n9307_));
  AOI21_X1   g06871(.A1(new_n9281_), .A2(new_n9271_), .B(new_n2672_), .ZN(new_n9308_));
  NOR2_X1    g06872(.A1(new_n9291_), .A2(new_n3025_), .ZN(new_n9309_));
  AOI21_X1   g06873(.A1(new_n9298_), .A2(new_n3025_), .B(new_n9309_), .ZN(new_n9310_));
  NOR2_X1    g06874(.A1(new_n9310_), .A2(pi0198), .ZN(new_n9311_));
  OAI21_X1   g06875(.A1(new_n9311_), .A2(new_n9308_), .B(new_n9307_), .ZN(new_n9312_));
  OR2_X2     g06876(.A1(new_n9304_), .A2(new_n9307_), .Z(new_n9313_));
  AOI21_X1   g06877(.A1(new_n9313_), .A2(new_n9312_), .B(pi0299), .ZN(new_n9314_));
  NOR2_X1    g06878(.A1(new_n8349_), .A2(new_n2689_), .ZN(new_n9315_));
  INV_X1     g06879(.I(new_n9315_), .ZN(new_n9316_));
  NOR2_X1    g06880(.A1(new_n9282_), .A2(new_n2709_), .ZN(new_n9317_));
  AOI21_X1   g06881(.A1(new_n9310_), .A2(new_n2709_), .B(new_n9317_), .ZN(new_n9318_));
  OAI21_X1   g06882(.A1(new_n9318_), .A2(new_n9316_), .B(pi0299), .ZN(new_n9319_));
  AOI21_X1   g06883(.A1(new_n9301_), .A2(new_n9316_), .B(new_n9319_), .ZN(new_n9320_));
  OAI21_X1   g06884(.A1(new_n9314_), .A2(new_n9320_), .B(pi0232), .ZN(new_n9321_));
  NAND3_X1   g06885(.A1(new_n9321_), .A2(new_n6350_), .A3(new_n9306_), .ZN(new_n9322_));
  NOR2_X1    g06886(.A1(po0740), .A2(pi0122), .ZN(new_n9323_));
  OAI21_X1   g06887(.A1(new_n9266_), .A2(new_n9323_), .B(po1057), .ZN(new_n9324_));
  NOR2_X1    g06888(.A1(new_n9274_), .A2(new_n6714_), .ZN(new_n9325_));
  AOI21_X1   g06889(.A1(pi0252), .A2(new_n3083_), .B(new_n9276_), .ZN(new_n9326_));
  NOR2_X1    g06890(.A1(new_n9326_), .A2(pi0122), .ZN(new_n9327_));
  OAI21_X1   g06891(.A1(new_n9325_), .A2(new_n9327_), .B(pi1093), .ZN(new_n9328_));
  INV_X1     g06892(.I(new_n9268_), .ZN(new_n9329_));
  AOI22_X1   g06893(.A1(new_n9270_), .A2(new_n6258_), .B1(new_n5331_), .B2(new_n9276_), .ZN(new_n9330_));
  AOI21_X1   g06894(.A1(new_n9330_), .A2(new_n9329_), .B(pi0122), .ZN(new_n9331_));
  OAI21_X1   g06895(.A1(new_n9331_), .A2(new_n9325_), .B(new_n3041_), .ZN(new_n9332_));
  AOI21_X1   g06896(.A1(new_n9332_), .A2(new_n9328_), .B(new_n3026_), .ZN(new_n9333_));
  NAND2_X1   g06897(.A1(new_n9276_), .A2(new_n6714_), .ZN(new_n9334_));
  NOR2_X1    g06898(.A1(new_n9269_), .A2(new_n6714_), .ZN(new_n9335_));
  INV_X1     g06899(.I(new_n9335_), .ZN(new_n9336_));
  AOI21_X1   g06900(.A1(new_n9336_), .A2(new_n9334_), .B(new_n3041_), .ZN(new_n9337_));
  INV_X1     g06901(.I(new_n9337_), .ZN(new_n9338_));
  AOI21_X1   g06902(.A1(new_n9332_), .A2(new_n9338_), .B(new_n3025_), .ZN(new_n9339_));
  OAI21_X1   g06903(.A1(new_n9333_), .A2(new_n9339_), .B(new_n5323_), .ZN(new_n9340_));
  AND2_X2    g06904(.A1(new_n9340_), .A2(new_n9324_), .Z(new_n9341_));
  NAND2_X1   g06905(.A1(new_n9341_), .A2(pi0210), .ZN(new_n9342_));
  NAND2_X1   g06906(.A1(po1057), .A2(pi0137), .ZN(new_n9343_));
  NOR2_X1    g06907(.A1(new_n3025_), .A2(pi0137), .ZN(new_n9344_));
  NOR3_X1    g06908(.A1(new_n2704_), .A2(new_n3040_), .A3(pi1093), .ZN(new_n9345_));
  NAND2_X1   g06909(.A1(new_n9345_), .A2(new_n3046_), .ZN(new_n9346_));
  NAND2_X1   g06910(.A1(new_n9346_), .A2(new_n3016_), .ZN(new_n9347_));
  OAI22_X1   g06911(.A1(new_n9339_), .A2(new_n9344_), .B1(new_n9276_), .B2(new_n9347_), .ZN(new_n9348_));
  INV_X1     g06912(.I(new_n9326_), .ZN(new_n9349_));
  NOR2_X1    g06913(.A1(new_n3026_), .A2(pi0137), .ZN(new_n9350_));
  OAI22_X1   g06914(.A1(new_n9333_), .A2(new_n9350_), .B1(pi0137), .B2(new_n9349_), .ZN(new_n9351_));
  NAND2_X1   g06915(.A1(new_n9351_), .A2(new_n9348_), .ZN(new_n9352_));
  OAI21_X1   g06916(.A1(new_n9352_), .A2(po1057), .B(new_n9343_), .ZN(new_n9353_));
  NAND2_X1   g06917(.A1(new_n9353_), .A2(new_n9324_), .ZN(new_n9354_));
  OAI21_X1   g06918(.A1(new_n9354_), .A2(pi0210), .B(new_n9342_), .ZN(new_n9355_));
  NAND2_X1   g06919(.A1(new_n9355_), .A2(pi0299), .ZN(new_n9356_));
  NAND2_X1   g06920(.A1(new_n9341_), .A2(pi0198), .ZN(new_n9357_));
  OAI21_X1   g06921(.A1(new_n9354_), .A2(pi0198), .B(new_n9357_), .ZN(new_n9358_));
  NAND2_X1   g06922(.A1(new_n9358_), .A2(new_n2628_), .ZN(new_n9359_));
  AOI21_X1   g06923(.A1(new_n9356_), .A2(new_n9359_), .B(pi0232), .ZN(new_n9360_));
  INV_X1     g06924(.I(new_n9307_), .ZN(new_n9361_));
  NOR2_X1    g06925(.A1(new_n9333_), .A2(new_n9339_), .ZN(new_n9362_));
  NAND2_X1   g06926(.A1(new_n9362_), .A2(pi0198), .ZN(new_n9363_));
  INV_X1     g06927(.I(new_n9352_), .ZN(new_n9364_));
  NAND2_X1   g06928(.A1(new_n9364_), .A2(new_n2672_), .ZN(new_n9365_));
  AOI21_X1   g06929(.A1(new_n9365_), .A2(new_n9363_), .B(new_n9361_), .ZN(new_n9366_));
  AND2_X2    g06930(.A1(new_n9358_), .A2(new_n9361_), .Z(new_n9367_));
  OAI21_X1   g06931(.A1(new_n9367_), .A2(new_n9366_), .B(new_n2628_), .ZN(new_n9368_));
  NAND2_X1   g06932(.A1(new_n9362_), .A2(pi0210), .ZN(new_n9369_));
  NAND2_X1   g06933(.A1(new_n9364_), .A2(new_n2709_), .ZN(new_n9370_));
  AOI21_X1   g06934(.A1(new_n9370_), .A2(new_n9369_), .B(new_n9316_), .ZN(new_n9371_));
  AND2_X2    g06935(.A1(new_n9355_), .A2(new_n9316_), .Z(new_n9372_));
  OAI21_X1   g06936(.A1(new_n9372_), .A2(new_n9371_), .B(pi0299), .ZN(new_n9373_));
  AOI21_X1   g06937(.A1(new_n9368_), .A2(new_n9373_), .B(new_n5666_), .ZN(new_n9374_));
  OAI21_X1   g06938(.A1(new_n9374_), .A2(new_n9360_), .B(new_n6349_), .ZN(new_n9375_));
  AOI21_X1   g06939(.A1(new_n9375_), .A2(new_n9322_), .B(new_n8260_), .ZN(po0234));
  NOR3_X1    g06940(.A1(new_n2874_), .A2(new_n2879_), .A3(new_n7293_), .ZN(new_n9377_));
  NAND2_X1   g06941(.A1(new_n9377_), .A2(pi0314), .ZN(new_n9378_));
  INV_X1     g06942(.I(new_n2882_), .ZN(new_n9379_));
  OAI21_X1   g06943(.A1(new_n9379_), .A2(new_n2866_), .B(new_n2879_), .ZN(new_n9380_));
  NAND2_X1   g06944(.A1(new_n5564_), .A2(new_n9380_), .ZN(new_n9381_));
  NOR2_X1    g06945(.A1(new_n9381_), .A2(new_n2737_), .ZN(new_n9382_));
  NAND2_X1   g06946(.A1(new_n9382_), .A2(new_n5590_), .ZN(new_n9383_));
  AOI21_X1   g06947(.A1(new_n9383_), .A2(new_n9378_), .B(new_n8262_), .ZN(po0235));
  NOR3_X1    g06948(.A1(new_n6240_), .A2(new_n5666_), .A3(pi0468), .ZN(po0236));
  NAND2_X1   g06949(.A1(new_n7915_), .A2(new_n7559_), .ZN(new_n9386_));
  INV_X1     g06950(.I(new_n7916_), .ZN(new_n9387_));
  NOR3_X1    g06951(.A1(new_n8086_), .A2(new_n9387_), .A3(new_n5636_), .ZN(new_n9388_));
  NOR2_X1    g06952(.A1(pi0162), .A2(pi0197), .ZN(new_n9389_));
  NOR3_X1    g06953(.A1(new_n5437_), .A2(new_n7916_), .A3(new_n9389_), .ZN(new_n9390_));
  NOR2_X1    g06954(.A1(new_n9388_), .A2(new_n9390_), .ZN(new_n9391_));
  INV_X1     g06955(.I(pi0163), .ZN(new_n9392_));
  NOR2_X1    g06956(.A1(new_n5437_), .A2(new_n9392_), .ZN(new_n9393_));
  NAND2_X1   g06957(.A1(new_n9391_), .A2(new_n9393_), .ZN(new_n9394_));
  OAI21_X1   g06958(.A1(pi0163), .A2(new_n9391_), .B(new_n9394_), .ZN(new_n9395_));
  INV_X1     g06959(.I(new_n9395_), .ZN(new_n9396_));
  NOR2_X1    g06960(.A1(new_n9396_), .A2(new_n5666_), .ZN(new_n9397_));
  NOR2_X1    g06961(.A1(new_n9397_), .A2(new_n7342_), .ZN(new_n9398_));
  INV_X1     g06962(.I(pi0147), .ZN(new_n9399_));
  NOR2_X1    g06963(.A1(new_n6698_), .A2(new_n9399_), .ZN(new_n9400_));
  AOI21_X1   g06964(.A1(new_n7342_), .A2(new_n9400_), .B(new_n9398_), .ZN(new_n9401_));
  INV_X1     g06965(.I(new_n9401_), .ZN(new_n9402_));
  AOI21_X1   g06966(.A1(new_n9397_), .A2(new_n7348_), .B(new_n2625_), .ZN(new_n9403_));
  NOR3_X1    g06967(.A1(new_n9402_), .A2(new_n3291_), .A3(new_n9403_), .ZN(new_n9404_));
  INV_X1     g06968(.I(new_n9403_), .ZN(new_n9405_));
  NOR2_X1    g06969(.A1(new_n9401_), .A2(new_n5499_), .ZN(new_n9406_));
  INV_X1     g06970(.I(new_n9406_), .ZN(new_n9407_));
  OAI21_X1   g06971(.A1(new_n9396_), .A2(new_n5666_), .B(pi0100), .ZN(new_n9408_));
  NOR2_X1    g06972(.A1(pi0038), .A2(pi0040), .ZN(new_n9409_));
  OAI21_X1   g06973(.A1(new_n9400_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n9410_));
  OAI21_X1   g06974(.A1(new_n9409_), .A2(new_n9410_), .B(new_n9408_), .ZN(new_n9411_));
  NOR2_X1    g06975(.A1(new_n9411_), .A2(new_n7596_), .ZN(new_n9412_));
  OAI22_X1   g06976(.A1(new_n9412_), .A2(new_n8108_), .B1(new_n3465_), .B2(new_n9397_), .ZN(new_n9413_));
  INV_X1     g06977(.I(new_n9409_), .ZN(new_n9414_));
  NOR3_X1    g06978(.A1(new_n9414_), .A2(new_n3458_), .A3(new_n2496_), .ZN(new_n9415_));
  INV_X1     g06979(.I(new_n9415_), .ZN(new_n9416_));
  OAI21_X1   g06980(.A1(new_n7756_), .A2(new_n2627_), .B(new_n8170_), .ZN(new_n9417_));
  AOI21_X1   g06981(.A1(new_n7597_), .A2(new_n2496_), .B(pi0040), .ZN(new_n9418_));
  AOI21_X1   g06982(.A1(new_n7580_), .A2(new_n5437_), .B(new_n7583_), .ZN(new_n9419_));
  NAND3_X1   g06983(.A1(new_n9419_), .A2(pi0163), .A3(pi0232), .ZN(new_n9420_));
  AOI21_X1   g06984(.A1(new_n9420_), .A2(new_n9418_), .B(pi0039), .ZN(new_n9421_));
  OAI21_X1   g06985(.A1(new_n9421_), .A2(new_n9417_), .B(new_n9416_), .ZN(new_n9422_));
  OAI21_X1   g06986(.A1(new_n9422_), .A2(new_n9410_), .B(new_n9408_), .ZN(new_n9423_));
  AOI21_X1   g06987(.A1(new_n9423_), .A2(new_n2605_), .B(new_n9413_), .ZN(new_n9424_));
  OAI21_X1   g06988(.A1(new_n9424_), .A2(pi0054), .B(new_n9407_), .ZN(new_n9425_));
  AOI21_X1   g06989(.A1(new_n9425_), .A2(new_n2625_), .B(new_n2602_), .ZN(new_n9426_));
  AOI21_X1   g06990(.A1(new_n9426_), .A2(new_n9405_), .B(new_n2471_), .ZN(new_n9427_));
  AND3_X2    g06991(.A1(new_n7940_), .A2(new_n5398_), .A3(new_n7937_), .Z(new_n9428_));
  NOR2_X1    g06992(.A1(new_n9428_), .A2(pi0184), .ZN(new_n9429_));
  INV_X1     g06993(.I(new_n9429_), .ZN(new_n9430_));
  OAI21_X1   g06994(.A1(new_n9428_), .A2(new_n5437_), .B(pi0184), .ZN(new_n9431_));
  AOI21_X1   g06995(.A1(new_n9430_), .A2(new_n9431_), .B(pi0299), .ZN(new_n9432_));
  OAI21_X1   g06996(.A1(new_n9395_), .A2(new_n2628_), .B(pi0232), .ZN(new_n9433_));
  NOR2_X1    g06997(.A1(new_n9432_), .A2(new_n9433_), .ZN(new_n9434_));
  INV_X1     g06998(.I(new_n9434_), .ZN(new_n9435_));
  NOR2_X1    g06999(.A1(new_n9435_), .A2(new_n7342_), .ZN(new_n9436_));
  INV_X1     g07000(.I(new_n9436_), .ZN(new_n9437_));
  AOI21_X1   g07001(.A1(new_n9437_), .A2(pi0074), .B(pi0055), .ZN(new_n9438_));
  INV_X1     g07002(.I(new_n9438_), .ZN(new_n9439_));
  INV_X1     g07003(.I(pi0187), .ZN(new_n9440_));
  NOR2_X1    g07004(.A1(new_n9440_), .A2(pi0299), .ZN(new_n9441_));
  AOI21_X1   g07005(.A1(pi0147), .A2(pi0299), .B(new_n9441_), .ZN(new_n9442_));
  NOR2_X1    g07006(.A1(new_n6698_), .A2(new_n9442_), .ZN(new_n9443_));
  NOR2_X1    g07007(.A1(new_n9443_), .A2(new_n7348_), .ZN(new_n9444_));
  NOR3_X1    g07008(.A1(new_n9436_), .A2(new_n5499_), .A3(new_n9444_), .ZN(new_n9445_));
  INV_X1     g07009(.I(new_n9445_), .ZN(new_n9446_));
  NOR2_X1    g07010(.A1(new_n9434_), .A2(new_n2702_), .ZN(new_n9447_));
  OAI21_X1   g07011(.A1(new_n9443_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n9448_));
  NOR2_X1    g07012(.A1(new_n9448_), .A2(new_n9415_), .ZN(new_n9449_));
  AOI21_X1   g07013(.A1(pi0087), .A2(new_n9449_), .B(new_n9447_), .ZN(new_n9450_));
  NOR2_X1    g07014(.A1(new_n7398_), .A2(new_n9440_), .ZN(new_n9451_));
  NOR2_X1    g07015(.A1(new_n7401_), .A2(pi0187), .ZN(new_n9452_));
  OAI21_X1   g07016(.A1(new_n9452_), .A2(new_n9451_), .B(pi0147), .ZN(new_n9453_));
  NOR3_X1    g07017(.A1(new_n7405_), .A2(pi0147), .A3(new_n9440_), .ZN(new_n9454_));
  INV_X1     g07018(.I(new_n9454_), .ZN(new_n9455_));
  AOI21_X1   g07019(.A1(new_n9453_), .A2(new_n9455_), .B(new_n3265_), .ZN(new_n9456_));
  AOI21_X1   g07020(.A1(new_n7608_), .A2(new_n5427_), .B(new_n7409_), .ZN(new_n9457_));
  NOR2_X1    g07021(.A1(new_n9457_), .A2(pi0040), .ZN(new_n9458_));
  INV_X1     g07022(.I(new_n9458_), .ZN(new_n9459_));
  NOR2_X1    g07023(.A1(new_n9459_), .A2(new_n5446_), .ZN(new_n9460_));
  NOR2_X1    g07024(.A1(new_n7609_), .A2(pi0040), .ZN(new_n9461_));
  INV_X1     g07025(.I(new_n9461_), .ZN(new_n9462_));
  NOR2_X1    g07026(.A1(new_n9462_), .A2(new_n5445_), .ZN(new_n9463_));
  OAI21_X1   g07027(.A1(new_n9460_), .A2(new_n9463_), .B(new_n7519_), .ZN(new_n9464_));
  NAND2_X1   g07028(.A1(new_n7525_), .A2(new_n7756_), .ZN(new_n9465_));
  AOI21_X1   g07029(.A1(new_n9464_), .A2(new_n9465_), .B(pi0299), .ZN(new_n9466_));
  NOR2_X1    g07030(.A1(new_n9462_), .A2(new_n6764_), .ZN(new_n9467_));
  AOI21_X1   g07031(.A1(new_n6764_), .A2(new_n9458_), .B(new_n9467_), .ZN(new_n9468_));
  OAI21_X1   g07032(.A1(new_n9468_), .A2(new_n7637_), .B(new_n5666_), .ZN(new_n9469_));
  NOR2_X1    g07033(.A1(new_n9469_), .A2(new_n9466_), .ZN(new_n9470_));
  INV_X1     g07034(.I(pi0156), .ZN(new_n9471_));
  NOR2_X1    g07035(.A1(new_n7608_), .A2(new_n7409_), .ZN(new_n9472_));
  NOR2_X1    g07036(.A1(new_n9472_), .A2(new_n6745_), .ZN(new_n9473_));
  AOI22_X1   g07037(.A1(new_n9473_), .A2(new_n2818_), .B1(new_n5413_), .B2(new_n7756_), .ZN(new_n9474_));
  OAI21_X1   g07038(.A1(new_n7626_), .A2(new_n7409_), .B(new_n7839_), .ZN(new_n9475_));
  NAND2_X1   g07039(.A1(new_n9474_), .A2(new_n9475_), .ZN(new_n9476_));
  INV_X1     g07040(.I(new_n9476_), .ZN(new_n9477_));
  NOR3_X1    g07041(.A1(new_n9477_), .A2(pi0166), .A3(new_n5422_), .ZN(new_n9478_));
  AOI21_X1   g07042(.A1(new_n3361_), .A2(new_n6764_), .B(new_n9468_), .ZN(new_n9479_));
  OAI21_X1   g07043(.A1(new_n9479_), .A2(new_n9478_), .B(new_n7508_), .ZN(new_n9480_));
  AOI21_X1   g07044(.A1(new_n8070_), .A2(new_n7756_), .B(new_n2628_), .ZN(new_n9481_));
  NAND2_X1   g07045(.A1(new_n9480_), .A2(new_n9481_), .ZN(new_n9482_));
  NOR2_X1    g07046(.A1(new_n9461_), .A2(pi0189), .ZN(new_n9483_));
  INV_X1     g07047(.I(pi0189), .ZN(new_n9484_));
  OAI21_X1   g07048(.A1(new_n7614_), .A2(new_n7409_), .B(new_n7839_), .ZN(new_n9485_));
  NAND2_X1   g07049(.A1(new_n9474_), .A2(new_n9485_), .ZN(new_n9486_));
  NOR3_X1    g07050(.A1(new_n9486_), .A2(new_n9484_), .A3(new_n5446_), .ZN(new_n9487_));
  OAI21_X1   g07051(.A1(new_n9487_), .A2(new_n9483_), .B(pi0179), .ZN(new_n9488_));
  INV_X1     g07052(.I(new_n9463_), .ZN(new_n9489_));
  NAND2_X1   g07053(.A1(new_n9459_), .A2(pi0189), .ZN(new_n9490_));
  NAND2_X1   g07054(.A1(new_n9477_), .A2(new_n9484_), .ZN(new_n9491_));
  AOI21_X1   g07055(.A1(new_n9491_), .A2(new_n9490_), .B(pi0179), .ZN(new_n9492_));
  OAI21_X1   g07056(.A1(new_n9492_), .A2(new_n5446_), .B(new_n9489_), .ZN(new_n9493_));
  NAND3_X1   g07057(.A1(new_n9493_), .A2(new_n7519_), .A3(new_n9488_), .ZN(new_n9494_));
  NAND3_X1   g07058(.A1(new_n9494_), .A2(new_n2628_), .A3(new_n9465_), .ZN(new_n9495_));
  NAND3_X1   g07059(.A1(new_n9495_), .A2(new_n9471_), .A3(new_n9482_), .ZN(new_n9496_));
  NOR2_X1    g07060(.A1(new_n5422_), .A2(new_n3361_), .ZN(new_n9497_));
  NOR2_X1    g07061(.A1(new_n9462_), .A2(new_n9497_), .ZN(new_n9498_));
  AOI21_X1   g07062(.A1(new_n9486_), .A2(new_n9497_), .B(new_n9498_), .ZN(new_n9499_));
  OAI21_X1   g07063(.A1(new_n9499_), .A2(new_n8070_), .B(new_n9481_), .ZN(new_n9500_));
  NAND3_X1   g07064(.A1(new_n9495_), .A2(pi0156), .A3(new_n9500_), .ZN(new_n9501_));
  AND3_X2    g07065(.A1(new_n9496_), .A2(new_n9501_), .A3(pi0232), .Z(new_n9502_));
  NOR3_X1    g07066(.A1(new_n9502_), .A2(new_n2627_), .A3(new_n9470_), .ZN(new_n9503_));
  INV_X1     g07067(.I(new_n7765_), .ZN(new_n9504_));
  AOI22_X1   g07068(.A1(new_n7676_), .A2(new_n7678_), .B1(new_n3028_), .B2(new_n9504_), .ZN(new_n9505_));
  NOR2_X1    g07069(.A1(new_n7806_), .A2(pi0040), .ZN(new_n9506_));
  INV_X1     g07070(.I(new_n9506_), .ZN(new_n9507_));
  AOI21_X1   g07071(.A1(new_n9507_), .A2(new_n2462_), .B(new_n9505_), .ZN(new_n9508_));
  INV_X1     g07072(.I(new_n9508_), .ZN(new_n9509_));
  NAND2_X1   g07073(.A1(new_n9509_), .A2(pi0299), .ZN(new_n9510_));
  OAI21_X1   g07074(.A1(new_n7833_), .A2(new_n7805_), .B(new_n2818_), .ZN(new_n9511_));
  AOI21_X1   g07075(.A1(new_n9511_), .A2(new_n2462_), .B(new_n9505_), .ZN(new_n9512_));
  OR2_X2     g07076(.A1(new_n9512_), .A2(pi0299), .Z(new_n9513_));
  AOI21_X1   g07077(.A1(new_n9510_), .A2(new_n9513_), .B(pi0232), .ZN(new_n9514_));
  NAND2_X1   g07078(.A1(new_n9512_), .A2(new_n5437_), .ZN(new_n9515_));
  NOR2_X1    g07079(.A1(pi0175), .A2(pi0299), .ZN(new_n9516_));
  INV_X1     g07080(.I(pi0184), .ZN(new_n9517_));
  AOI21_X1   g07081(.A1(new_n7795_), .A2(new_n2818_), .B(pi0032), .ZN(new_n9518_));
  INV_X1     g07082(.I(new_n9518_), .ZN(new_n9519_));
  AOI21_X1   g07083(.A1(new_n9519_), .A2(new_n7758_), .B(pi0095), .ZN(new_n9520_));
  INV_X1     g07084(.I(new_n9520_), .ZN(new_n9521_));
  NAND2_X1   g07085(.A1(new_n9521_), .A2(new_n9504_), .ZN(new_n9522_));
  NOR2_X1    g07086(.A1(new_n9522_), .A2(new_n2672_), .ZN(new_n9523_));
  AOI21_X1   g07087(.A1(new_n9519_), .A2(new_n7763_), .B(pi0095), .ZN(new_n9524_));
  INV_X1     g07088(.I(new_n9524_), .ZN(new_n9525_));
  NAND2_X1   g07089(.A1(new_n9525_), .A2(new_n9504_), .ZN(new_n9526_));
  NOR2_X1    g07090(.A1(new_n9526_), .A2(pi0198), .ZN(new_n9527_));
  OAI21_X1   g07091(.A1(new_n9523_), .A2(new_n9527_), .B(new_n8354_), .ZN(new_n9528_));
  NAND3_X1   g07092(.A1(new_n9528_), .A2(pi0182), .A3(new_n9517_), .ZN(new_n9529_));
  NOR2_X1    g07093(.A1(new_n5437_), .A2(new_n9484_), .ZN(new_n9530_));
  INV_X1     g07094(.I(new_n9530_), .ZN(new_n9531_));
  NOR2_X1    g07095(.A1(new_n9511_), .A2(new_n9531_), .ZN(new_n9532_));
  OAI21_X1   g07096(.A1(new_n7701_), .A2(pi0040), .B(new_n2462_), .ZN(new_n9533_));
  NOR2_X1    g07097(.A1(new_n7710_), .A2(pi0040), .ZN(new_n9534_));
  AOI21_X1   g07098(.A1(new_n9534_), .A2(pi0189), .B(new_n9533_), .ZN(new_n9535_));
  AOI21_X1   g07099(.A1(new_n9505_), .A2(new_n5659_), .B(new_n5437_), .ZN(new_n9536_));
  OAI21_X1   g07100(.A1(new_n5659_), .A2(new_n9504_), .B(new_n9536_), .ZN(new_n9537_));
  NOR2_X1    g07101(.A1(new_n9535_), .A2(new_n9537_), .ZN(new_n9538_));
  OAI22_X1   g07102(.A1(new_n9529_), .A2(new_n9532_), .B1(new_n9517_), .B2(new_n9538_), .ZN(new_n9539_));
  NAND2_X1   g07103(.A1(new_n9539_), .A2(new_n9516_), .ZN(new_n9540_));
  INV_X1     g07104(.I(pi0175), .ZN(new_n9541_));
  NOR2_X1    g07105(.A1(new_n9541_), .A2(pi0299), .ZN(new_n9542_));
  OAI21_X1   g07106(.A1(new_n7760_), .A2(pi0095), .B(new_n9504_), .ZN(new_n9543_));
  NOR2_X1    g07107(.A1(new_n9543_), .A2(new_n2672_), .ZN(new_n9544_));
  NOR2_X1    g07108(.A1(new_n7766_), .A2(pi0198), .ZN(new_n9545_));
  OAI21_X1   g07109(.A1(new_n9544_), .A2(new_n9545_), .B(new_n9530_), .ZN(new_n9546_));
  NOR2_X1    g07110(.A1(new_n7865_), .A2(new_n8355_), .ZN(new_n9547_));
  NOR2_X1    g07111(.A1(new_n9547_), .A2(new_n5659_), .ZN(new_n9548_));
  INV_X1     g07112(.I(new_n9505_), .ZN(new_n9549_));
  OAI21_X1   g07113(.A1(new_n7760_), .A2(pi0095), .B(new_n9549_), .ZN(new_n9550_));
  NOR2_X1    g07114(.A1(new_n9550_), .A2(new_n2672_), .ZN(new_n9551_));
  OR2_X2     g07115(.A1(new_n7764_), .A2(new_n9505_), .Z(new_n9552_));
  NOR2_X1    g07116(.A1(new_n9552_), .A2(pi0198), .ZN(new_n9553_));
  OAI21_X1   g07117(.A1(new_n9551_), .A2(new_n9553_), .B(new_n9530_), .ZN(new_n9554_));
  AOI22_X1   g07118(.A1(new_n9548_), .A2(new_n9546_), .B1(new_n9554_), .B2(new_n5659_), .ZN(new_n9555_));
  NAND2_X1   g07119(.A1(new_n5659_), .A2(pi0095), .ZN(new_n9556_));
  NAND2_X1   g07120(.A1(new_n9549_), .A2(new_n8354_), .ZN(new_n9557_));
  AOI21_X1   g07121(.A1(new_n7865_), .A2(new_n9556_), .B(new_n9557_), .ZN(new_n9558_));
  OAI21_X1   g07122(.A1(new_n9555_), .A2(new_n9558_), .B(new_n9517_), .ZN(new_n9559_));
  NAND2_X1   g07123(.A1(new_n9559_), .A2(new_n9542_), .ZN(new_n9560_));
  NAND2_X1   g07124(.A1(new_n7719_), .A2(new_n2818_), .ZN(new_n9561_));
  AOI21_X1   g07125(.A1(new_n2462_), .A2(pi0189), .B(new_n7409_), .ZN(new_n9562_));
  OAI21_X1   g07126(.A1(new_n9561_), .A2(new_n9562_), .B(new_n9556_), .ZN(new_n9563_));
  AND3_X2    g07127(.A1(new_n9536_), .A2(pi0184), .A3(new_n9563_), .Z(new_n9564_));
  OAI21_X1   g07128(.A1(new_n9560_), .A2(new_n9564_), .B(new_n9540_), .ZN(new_n9565_));
  NOR3_X1    g07129(.A1(new_n9520_), .A2(new_n2672_), .A3(new_n9505_), .ZN(new_n9566_));
  NOR3_X1    g07130(.A1(new_n9524_), .A2(pi0198), .A3(new_n9505_), .ZN(new_n9567_));
  OAI21_X1   g07131(.A1(new_n9566_), .A2(new_n9567_), .B(new_n8354_), .ZN(new_n9568_));
  NAND4_X1   g07132(.A1(new_n9568_), .A2(new_n5659_), .A3(new_n9517_), .A4(new_n9516_), .ZN(new_n9569_));
  AOI21_X1   g07133(.A1(new_n9512_), .A2(new_n8355_), .B(new_n9569_), .ZN(new_n9570_));
  AOI21_X1   g07134(.A1(new_n9565_), .A2(new_n9515_), .B(new_n9570_), .ZN(new_n9571_));
  AOI21_X1   g07135(.A1(new_n9508_), .A2(new_n5437_), .B(new_n2628_), .ZN(new_n9572_));
  NAND2_X1   g07136(.A1(new_n7862_), .A2(pi0210), .ZN(new_n9573_));
  NOR2_X1    g07137(.A1(new_n7863_), .A2(new_n7765_), .ZN(new_n9574_));
  NAND2_X1   g07138(.A1(new_n9574_), .A2(new_n2709_), .ZN(new_n9575_));
  AOI21_X1   g07139(.A1(new_n9573_), .A2(new_n9575_), .B(new_n8349_), .ZN(new_n9576_));
  NOR2_X1    g07140(.A1(new_n5437_), .A2(new_n3361_), .ZN(new_n9577_));
  NOR2_X1    g07141(.A1(new_n9543_), .A2(new_n2709_), .ZN(new_n9578_));
  NOR2_X1    g07142(.A1(new_n7766_), .A2(pi0210), .ZN(new_n9579_));
  OAI21_X1   g07143(.A1(new_n9578_), .A2(new_n9579_), .B(new_n9577_), .ZN(new_n9580_));
  NAND2_X1   g07144(.A1(new_n9580_), .A2(pi0153), .ZN(new_n9581_));
  OAI21_X1   g07145(.A1(new_n9581_), .A2(new_n9576_), .B(pi0160), .ZN(new_n9582_));
  NOR2_X1    g07146(.A1(new_n9522_), .A2(new_n2709_), .ZN(new_n9583_));
  NOR2_X1    g07147(.A1(new_n9526_), .A2(pi0210), .ZN(new_n9584_));
  OAI21_X1   g07148(.A1(new_n9583_), .A2(new_n9584_), .B(new_n8348_), .ZN(new_n9585_));
  NAND2_X1   g07149(.A1(new_n9585_), .A2(new_n2455_), .ZN(new_n9586_));
  AOI21_X1   g07150(.A1(new_n9506_), .A2(new_n9577_), .B(new_n9586_), .ZN(new_n9587_));
  NOR2_X1    g07151(.A1(new_n9587_), .A2(new_n9582_), .ZN(new_n9588_));
  OAI21_X1   g07152(.A1(new_n7861_), .A2(new_n9505_), .B(pi0210), .ZN(new_n9589_));
  OAI21_X1   g07153(.A1(new_n7863_), .A2(new_n9505_), .B(new_n2709_), .ZN(new_n9590_));
  AND3_X2    g07154(.A1(new_n9589_), .A2(new_n9590_), .A3(new_n8348_), .Z(new_n9591_));
  NOR2_X1    g07155(.A1(new_n9550_), .A2(new_n2709_), .ZN(new_n9592_));
  NOR2_X1    g07156(.A1(new_n9552_), .A2(pi0210), .ZN(new_n9593_));
  OAI21_X1   g07157(.A1(new_n9592_), .A2(new_n9593_), .B(new_n9577_), .ZN(new_n9594_));
  NAND2_X1   g07158(.A1(new_n9594_), .A2(pi0153), .ZN(new_n9595_));
  OAI21_X1   g07159(.A1(new_n9595_), .A2(new_n9591_), .B(new_n5635_), .ZN(new_n9596_));
  NAND3_X1   g07160(.A1(new_n9521_), .A2(pi0210), .A3(new_n9549_), .ZN(new_n9597_));
  NAND3_X1   g07161(.A1(new_n9525_), .A2(new_n2709_), .A3(new_n9549_), .ZN(new_n9598_));
  AOI21_X1   g07162(.A1(new_n9597_), .A2(new_n9598_), .B(new_n8349_), .ZN(new_n9599_));
  NOR2_X1    g07163(.A1(new_n9509_), .A2(new_n3361_), .ZN(new_n9600_));
  NOR3_X1    g07164(.A1(new_n9600_), .A2(pi0153), .A3(new_n9599_), .ZN(new_n9601_));
  OAI21_X1   g07165(.A1(new_n9601_), .A2(new_n9596_), .B(new_n9392_), .ZN(new_n9602_));
  NAND2_X1   g07166(.A1(new_n9561_), .A2(new_n2462_), .ZN(new_n9603_));
  NAND2_X1   g07167(.A1(new_n9245_), .A2(new_n3361_), .ZN(new_n9604_));
  AOI21_X1   g07168(.A1(new_n9603_), .A2(new_n9604_), .B(new_n2455_), .ZN(new_n9605_));
  NOR4_X1    g07169(.A1(new_n9505_), .A2(new_n9605_), .A3(pi0160), .A4(new_n5437_), .ZN(new_n9606_));
  AOI21_X1   g07170(.A1(new_n9534_), .A2(pi0166), .B(new_n9533_), .ZN(new_n9607_));
  NAND2_X1   g07171(.A1(new_n9607_), .A2(new_n2455_), .ZN(new_n9608_));
  AOI21_X1   g07172(.A1(new_n9608_), .A2(new_n9606_), .B(new_n9392_), .ZN(new_n9609_));
  NOR2_X1    g07173(.A1(new_n9607_), .A2(new_n5437_), .ZN(new_n9610_));
  AOI21_X1   g07174(.A1(new_n9610_), .A2(new_n9504_), .B(pi0153), .ZN(new_n9611_));
  AOI21_X1   g07175(.A1(new_n8348_), .A2(new_n7756_), .B(new_n2455_), .ZN(new_n9612_));
  NAND3_X1   g07176(.A1(new_n9603_), .A2(new_n9504_), .A3(new_n9577_), .ZN(new_n9613_));
  NAND2_X1   g07177(.A1(new_n9613_), .A2(new_n9612_), .ZN(new_n9614_));
  NAND2_X1   g07178(.A1(new_n9614_), .A2(pi0160), .ZN(new_n9615_));
  OAI21_X1   g07179(.A1(new_n9611_), .A2(new_n9615_), .B(new_n9609_), .ZN(new_n9616_));
  OAI21_X1   g07180(.A1(new_n9602_), .A2(new_n9588_), .B(new_n9616_), .ZN(new_n9617_));
  NAND2_X1   g07181(.A1(new_n9617_), .A2(new_n9572_), .ZN(new_n9618_));
  AOI21_X1   g07182(.A1(new_n9571_), .A2(new_n9618_), .B(new_n5666_), .ZN(new_n9619_));
  NOR3_X1    g07183(.A1(new_n9619_), .A2(pi0039), .A3(new_n9514_), .ZN(new_n9620_));
  NOR3_X1    g07184(.A1(new_n9620_), .A2(pi0038), .A3(new_n9503_), .ZN(new_n9621_));
  OAI21_X1   g07185(.A1(new_n9621_), .A2(new_n9456_), .B(new_n2603_), .ZN(new_n9622_));
  AOI21_X1   g07186(.A1(new_n9622_), .A2(new_n9450_), .B(new_n2606_), .ZN(new_n9623_));
  INV_X1     g07187(.I(new_n9417_), .ZN(new_n9624_));
  INV_X1     g07188(.I(new_n9418_), .ZN(new_n9625_));
  NOR2_X1    g07189(.A1(new_n9471_), .A2(new_n2628_), .ZN(new_n9626_));
  INV_X1     g07190(.I(pi0179), .ZN(new_n9627_));
  NOR2_X1    g07191(.A1(new_n9627_), .A2(pi0299), .ZN(new_n9628_));
  OAI21_X1   g07192(.A1(new_n9626_), .A2(new_n9628_), .B(new_n6697_), .ZN(new_n9629_));
  NOR2_X1    g07193(.A1(new_n9629_), .A2(new_n7409_), .ZN(new_n9630_));
  OAI21_X1   g07194(.A1(new_n9625_), .A2(new_n9630_), .B(new_n2627_), .ZN(new_n9631_));
  NAND2_X1   g07195(.A1(new_n9631_), .A2(new_n9624_), .ZN(new_n9632_));
  AOI21_X1   g07196(.A1(new_n9632_), .A2(new_n9449_), .B(new_n9447_), .ZN(new_n9633_));
  OAI22_X1   g07197(.A1(new_n9633_), .A2(new_n8108_), .B1(new_n3465_), .B2(new_n9434_), .ZN(new_n9634_));
  OAI21_X1   g07198(.A1(new_n9623_), .A2(new_n9634_), .B(new_n5499_), .ZN(new_n9635_));
  AOI21_X1   g07199(.A1(new_n9635_), .A2(new_n9446_), .B(pi0074), .ZN(new_n9636_));
  OAI21_X1   g07200(.A1(new_n9636_), .A2(new_n9439_), .B(new_n9427_), .ZN(new_n9637_));
  NOR2_X1    g07201(.A1(new_n9397_), .A2(new_n3465_), .ZN(new_n9638_));
  AOI21_X1   g07202(.A1(new_n9411_), .A2(new_n3465_), .B(new_n9638_), .ZN(new_n9639_));
  OAI21_X1   g07203(.A1(new_n9639_), .A2(pi0054), .B(new_n9407_), .ZN(new_n9640_));
  AOI21_X1   g07204(.A1(new_n9640_), .A2(new_n2625_), .B(new_n9403_), .ZN(new_n9641_));
  OAI21_X1   g07205(.A1(new_n9641_), .A2(new_n2470_), .B(new_n3291_), .ZN(new_n9642_));
  NOR2_X1    g07206(.A1(new_n9642_), .A2(new_n7906_), .ZN(new_n9643_));
  AOI21_X1   g07207(.A1(new_n9637_), .A2(new_n9643_), .B(new_n9404_), .ZN(new_n9644_));
  INV_X1     g07208(.I(new_n9404_), .ZN(new_n9645_));
  INV_X1     g07209(.I(new_n9447_), .ZN(new_n9646_));
  INV_X1     g07210(.I(new_n9448_), .ZN(new_n9647_));
  NOR4_X1    g07211(.A1(new_n2553_), .A2(new_n7456_), .A3(new_n7599_), .A4(new_n9629_), .ZN(new_n9648_));
  OAI21_X1   g07212(.A1(new_n9648_), .A2(new_n9414_), .B(new_n9647_), .ZN(new_n9649_));
  NAND2_X1   g07213(.A1(new_n9649_), .A2(new_n9646_), .ZN(new_n9650_));
  AOI22_X1   g07214(.A1(new_n9650_), .A2(new_n7387_), .B1(pi0075), .B2(new_n9435_), .ZN(new_n9651_));
  NAND3_X1   g07215(.A1(new_n9647_), .A2(pi0087), .A3(new_n9414_), .ZN(new_n9652_));
  NAND2_X1   g07216(.A1(new_n9646_), .A2(new_n9652_), .ZN(new_n9653_));
  INV_X1     g07217(.I(new_n9456_), .ZN(new_n9654_));
  NOR2_X1    g07218(.A1(new_n7456_), .A2(new_n5437_), .ZN(new_n9655_));
  NAND2_X1   g07219(.A1(new_n2552_), .A2(new_n9655_), .ZN(new_n9656_));
  AOI22_X1   g07220(.A1(new_n7606_), .A2(new_n9484_), .B1(pi0179), .B2(new_n5397_), .ZN(new_n9657_));
  NOR4_X1    g07221(.A1(new_n9657_), .A2(new_n5446_), .A3(new_n7525_), .A4(new_n9656_), .ZN(new_n9658_));
  NOR3_X1    g07222(.A1(new_n9658_), .A2(pi0040), .A3(pi0299), .ZN(new_n9659_));
  AOI22_X1   g07223(.A1(new_n7606_), .A2(new_n3361_), .B1(pi0156), .B2(new_n5397_), .ZN(new_n9660_));
  NOR4_X1    g07224(.A1(new_n9660_), .A2(new_n5422_), .A3(new_n8070_), .A4(new_n9656_), .ZN(new_n9661_));
  NOR3_X1    g07225(.A1(new_n9661_), .A2(pi0040), .A3(new_n2628_), .ZN(new_n9662_));
  NOR3_X1    g07226(.A1(new_n9659_), .A2(new_n9662_), .A3(new_n2627_), .ZN(new_n9663_));
  INV_X1     g07227(.I(new_n9516_), .ZN(new_n9664_));
  OAI21_X1   g07228(.A1(new_n7435_), .A2(new_n5647_), .B(pi0184), .ZN(new_n9665_));
  NAND2_X1   g07229(.A1(new_n7472_), .A2(new_n9517_), .ZN(new_n9666_));
  AOI21_X1   g07230(.A1(new_n9665_), .A2(new_n9666_), .B(pi0189), .ZN(new_n9667_));
  NAND2_X1   g07231(.A1(new_n7482_), .A2(pi0184), .ZN(new_n9668_));
  NOR3_X1    g07232(.A1(new_n2553_), .A2(pi0032), .A3(new_n3028_), .ZN(new_n9669_));
  INV_X1     g07233(.I(new_n9669_), .ZN(new_n9670_));
  OAI22_X1   g07234(.A1(new_n9668_), .A2(new_n9484_), .B1(new_n5659_), .B2(new_n9670_), .ZN(new_n9671_));
  OAI21_X1   g07235(.A1(new_n9667_), .A2(new_n9671_), .B(new_n5398_), .ZN(new_n9672_));
  AOI21_X1   g07236(.A1(new_n9672_), .A2(new_n2818_), .B(new_n9664_), .ZN(new_n9673_));
  INV_X1     g07237(.I(new_n9542_), .ZN(new_n9674_));
  NOR2_X1    g07238(.A1(new_n9669_), .A2(pi0040), .ZN(new_n9675_));
  AOI21_X1   g07239(.A1(new_n7489_), .A2(new_n9675_), .B(new_n9531_), .ZN(new_n9676_));
  NAND2_X1   g07240(.A1(new_n5437_), .A2(pi0040), .ZN(new_n9677_));
  NAND2_X1   g07241(.A1(new_n9677_), .A2(pi0184), .ZN(new_n9678_));
  INV_X1     g07242(.I(new_n7497_), .ZN(new_n9679_));
  INV_X1     g07243(.I(new_n9675_), .ZN(new_n9680_));
  NOR2_X1    g07244(.A1(new_n7442_), .A2(new_n9680_), .ZN(new_n9681_));
  AOI21_X1   g07245(.A1(new_n9679_), .A2(new_n9681_), .B(new_n8355_), .ZN(new_n9682_));
  NOR4_X1    g07246(.A1(new_n9682_), .A2(new_n5659_), .A3(new_n9676_), .A4(new_n9678_), .ZN(new_n9683_));
  NAND2_X1   g07247(.A1(new_n7490_), .A2(pi0189), .ZN(new_n9684_));
  INV_X1     g07248(.I(new_n7498_), .ZN(new_n9685_));
  NAND2_X1   g07249(.A1(new_n9685_), .A2(new_n8354_), .ZN(new_n9686_));
  NAND4_X1   g07250(.A1(new_n9686_), .A2(new_n5659_), .A3(pi0184), .A4(new_n9684_), .ZN(new_n9687_));
  NOR2_X1    g07251(.A1(new_n9670_), .A2(new_n5659_), .ZN(new_n9688_));
  NAND2_X1   g07252(.A1(new_n7460_), .A2(pi0189), .ZN(new_n9689_));
  NAND2_X1   g07253(.A1(new_n7465_), .A2(new_n9484_), .ZN(new_n9690_));
  AOI21_X1   g07254(.A1(new_n9690_), .A2(new_n9689_), .B(new_n7456_), .ZN(new_n9691_));
  OAI21_X1   g07255(.A1(new_n9691_), .A2(new_n9688_), .B(new_n5398_), .ZN(new_n9692_));
  NAND2_X1   g07256(.A1(new_n9692_), .A2(new_n9517_), .ZN(new_n9693_));
  AOI21_X1   g07257(.A1(new_n9687_), .A2(new_n9693_), .B(pi0040), .ZN(new_n9694_));
  NOR3_X1    g07258(.A1(new_n9694_), .A2(new_n9674_), .A3(new_n9683_), .ZN(new_n9695_));
  NAND2_X1   g07259(.A1(new_n7472_), .A2(new_n8348_), .ZN(new_n9696_));
  NAND3_X1   g07260(.A1(new_n7460_), .A2(pi0153), .A3(new_n9655_), .ZN(new_n9697_));
  NAND4_X1   g07261(.A1(new_n9697_), .A2(new_n2818_), .A3(new_n9392_), .A4(new_n9696_), .ZN(new_n9698_));
  NOR2_X1    g07262(.A1(new_n9670_), .A2(new_n5437_), .ZN(new_n9699_));
  OAI21_X1   g07263(.A1(new_n9698_), .A2(new_n9699_), .B(pi0299), .ZN(new_n9700_));
  OAI21_X1   g07264(.A1(new_n2455_), .A2(new_n7441_), .B(new_n7436_), .ZN(new_n9701_));
  NAND2_X1   g07265(.A1(new_n9701_), .A2(new_n8348_), .ZN(new_n9702_));
  NOR2_X1    g07266(.A1(new_n8123_), .A2(new_n2455_), .ZN(new_n9703_));
  OAI21_X1   g07267(.A1(new_n9703_), .A2(new_n8122_), .B(new_n9577_), .ZN(new_n9704_));
  NAND4_X1   g07268(.A1(new_n9702_), .A2(new_n2818_), .A3(pi0163), .A4(new_n9704_), .ZN(new_n9705_));
  NAND3_X1   g07269(.A1(new_n9705_), .A2(new_n5635_), .A3(new_n9698_), .ZN(new_n9706_));
  OAI21_X1   g07270(.A1(new_n7435_), .A2(new_n5615_), .B(new_n2709_), .ZN(new_n9707_));
  AOI21_X1   g07271(.A1(new_n9681_), .A2(new_n9707_), .B(new_n8349_), .ZN(new_n9708_));
  INV_X1     g07272(.I(new_n9577_), .ZN(new_n9709_));
  NOR2_X1    g07273(.A1(new_n8122_), .A2(new_n9680_), .ZN(new_n9710_));
  AOI21_X1   g07274(.A1(new_n9710_), .A2(new_n8123_), .B(new_n9709_), .ZN(new_n9711_));
  NOR3_X1    g07275(.A1(new_n9708_), .A2(new_n2455_), .A3(new_n9711_), .ZN(new_n9712_));
  NAND2_X1   g07276(.A1(new_n7436_), .A2(new_n9675_), .ZN(new_n9713_));
  OAI21_X1   g07277(.A1(new_n9710_), .A2(new_n9709_), .B(new_n2455_), .ZN(new_n9714_));
  AOI21_X1   g07278(.A1(new_n9713_), .A2(new_n8348_), .B(new_n9714_), .ZN(new_n9715_));
  NOR2_X1    g07279(.A1(new_n9712_), .A2(new_n9715_), .ZN(new_n9716_));
  NAND2_X1   g07280(.A1(new_n9677_), .A2(pi0163), .ZN(new_n9717_));
  OAI21_X1   g07281(.A1(new_n9716_), .A2(new_n9717_), .B(pi0160), .ZN(new_n9718_));
  AOI21_X1   g07282(.A1(new_n9718_), .A2(new_n9706_), .B(new_n9700_), .ZN(new_n9719_));
  NOR3_X1    g07283(.A1(new_n9719_), .A2(new_n9695_), .A3(new_n9673_), .ZN(new_n9720_));
  OAI21_X1   g07284(.A1(new_n9720_), .A2(pi0039), .B(pi0232), .ZN(new_n9721_));
  AOI21_X1   g07285(.A1(new_n2818_), .A2(new_n5666_), .B(pi0038), .ZN(new_n9722_));
  OAI21_X1   g07286(.A1(new_n9721_), .A2(new_n9663_), .B(new_n9722_), .ZN(new_n9723_));
  AOI21_X1   g07287(.A1(new_n9723_), .A2(new_n9654_), .B(new_n2604_), .ZN(new_n9724_));
  OAI21_X1   g07288(.A1(new_n9724_), .A2(new_n9653_), .B(new_n2605_), .ZN(new_n9725_));
  AOI21_X1   g07289(.A1(new_n9725_), .A2(new_n9651_), .B(pi0054), .ZN(new_n9726_));
  OAI21_X1   g07290(.A1(new_n9726_), .A2(new_n9445_), .B(new_n2625_), .ZN(new_n9727_));
  NAND4_X1   g07291(.A1(new_n7598_), .A2(new_n3444_), .A3(pi0163), .A4(pi0232), .ZN(new_n9728_));
  OAI21_X1   g07292(.A1(new_n9656_), .A2(new_n9728_), .B(new_n9409_), .ZN(new_n9729_));
  NOR2_X1    g07293(.A1(new_n9410_), .A2(pi0075), .ZN(new_n9730_));
  AOI21_X1   g07294(.A1(new_n9729_), .A2(new_n9730_), .B(new_n9398_), .ZN(new_n9731_));
  NOR2_X1    g07295(.A1(new_n9731_), .A2(pi0054), .ZN(new_n9732_));
  OAI21_X1   g07296(.A1(new_n9732_), .A2(new_n9406_), .B(new_n2625_), .ZN(new_n9733_));
  NAND3_X1   g07297(.A1(new_n9733_), .A2(pi0055), .A3(new_n9405_), .ZN(new_n9734_));
  NAND2_X1   g07298(.A1(new_n9734_), .A2(new_n2470_), .ZN(new_n9735_));
  AOI21_X1   g07299(.A1(new_n9727_), .A2(new_n9438_), .B(new_n9735_), .ZN(new_n9736_));
  OAI21_X1   g07300(.A1(new_n9736_), .A2(new_n9642_), .B(new_n9645_), .ZN(new_n9737_));
  NAND2_X1   g07301(.A1(new_n9737_), .A2(pi0079), .ZN(new_n9738_));
  OAI21_X1   g07302(.A1(new_n9644_), .A2(pi0079), .B(new_n9738_), .ZN(new_n9739_));
  NAND2_X1   g07303(.A1(new_n9739_), .A2(new_n9386_), .ZN(new_n9740_));
  NOR2_X1    g07304(.A1(new_n7563_), .A2(pi0079), .ZN(new_n9741_));
  NOR2_X1    g07305(.A1(new_n9644_), .A2(new_n9741_), .ZN(new_n9742_));
  AOI21_X1   g07306(.A1(new_n9737_), .A2(new_n9741_), .B(new_n9742_), .ZN(new_n9743_));
  OAI21_X1   g07307(.A1(new_n9743_), .A2(new_n9386_), .B(new_n9740_), .ZN(po0237));
  NOR2_X1    g07308(.A1(new_n2887_), .A2(new_n3040_), .ZN(new_n9745_));
  INV_X1     g07309(.I(new_n9745_), .ZN(new_n9746_));
  NOR2_X1    g07310(.A1(new_n9746_), .A2(new_n3041_), .ZN(new_n9747_));
  NOR2_X1    g07311(.A1(new_n3043_), .A2(pi0567), .ZN(new_n9748_));
  NOR2_X1    g07312(.A1(new_n9747_), .A2(new_n9748_), .ZN(new_n9749_));
  OAI21_X1   g07313(.A1(new_n9749_), .A2(pi0080), .B(pi0217), .ZN(new_n9750_));
  INV_X1     g07314(.I(pi0217), .ZN(new_n9751_));
  INV_X1     g07315(.I(new_n9749_), .ZN(new_n9752_));
  OAI21_X1   g07316(.A1(new_n9752_), .A2(new_n6350_), .B(po1038), .ZN(new_n9753_));
  NOR2_X1    g07317(.A1(new_n9753_), .A2(pi0080), .ZN(new_n9754_));
  AOI21_X1   g07318(.A1(new_n6301_), .A2(pi0592), .B(new_n6269_), .ZN(new_n9755_));
  NAND2_X1   g07319(.A1(new_n6320_), .A2(new_n9755_), .ZN(new_n9756_));
  NAND2_X1   g07320(.A1(new_n9756_), .A2(new_n9749_), .ZN(new_n9757_));
  AOI21_X1   g07321(.A1(new_n9757_), .A2(new_n6380_), .B(new_n6254_), .ZN(new_n9758_));
  INV_X1     g07322(.I(new_n6331_), .ZN(new_n9759_));
  INV_X1     g07323(.I(pi0448), .ZN(new_n9760_));
  INV_X1     g07324(.I(new_n9757_), .ZN(new_n9761_));
  NOR2_X1    g07325(.A1(new_n6271_), .A2(new_n9752_), .ZN(new_n9762_));
  AOI22_X1   g07326(.A1(new_n9761_), .A2(new_n6849_), .B1(new_n6851_), .B2(new_n9762_), .ZN(new_n9763_));
  AOI22_X1   g07327(.A1(new_n9761_), .A2(new_n6851_), .B1(new_n6849_), .B2(new_n9762_), .ZN(new_n9764_));
  OAI22_X1   g07328(.A1(new_n6853_), .A2(new_n9764_), .B1(new_n9763_), .B2(new_n6856_), .ZN(new_n9765_));
  AND2_X2    g07329(.A1(new_n9765_), .A2(pi0445), .Z(new_n9766_));
  OAI22_X1   g07330(.A1(new_n6853_), .A2(new_n9763_), .B1(new_n9764_), .B2(new_n6856_), .ZN(new_n9767_));
  AOI21_X1   g07331(.A1(new_n6859_), .A2(new_n9767_), .B(new_n9766_), .ZN(new_n9768_));
  NOR2_X1    g07332(.A1(new_n9768_), .A2(new_n9760_), .ZN(new_n9769_));
  AND2_X2    g07333(.A1(new_n9767_), .A2(pi0445), .Z(new_n9770_));
  AOI21_X1   g07334(.A1(new_n6859_), .A2(new_n9765_), .B(new_n9770_), .ZN(new_n9771_));
  NOR2_X1    g07335(.A1(new_n9771_), .A2(pi0448), .ZN(new_n9772_));
  OAI21_X1   g07336(.A1(new_n9769_), .A2(new_n9772_), .B(new_n9759_), .ZN(new_n9773_));
  NOR2_X1    g07337(.A1(new_n9771_), .A2(new_n9760_), .ZN(new_n9774_));
  NOR2_X1    g07338(.A1(new_n9768_), .A2(pi0448), .ZN(new_n9775_));
  OAI21_X1   g07339(.A1(new_n9774_), .A2(new_n9775_), .B(new_n6331_), .ZN(new_n9776_));
  NAND3_X1   g07340(.A1(new_n9773_), .A2(new_n9776_), .A3(pi1199), .ZN(new_n9777_));
  AOI21_X1   g07341(.A1(new_n9749_), .A2(new_n6254_), .B(new_n6251_), .ZN(new_n9778_));
  INV_X1     g07342(.I(new_n9778_), .ZN(new_n9779_));
  AOI21_X1   g07343(.A1(new_n9777_), .A2(new_n9758_), .B(new_n9779_), .ZN(new_n9780_));
  AOI21_X1   g07344(.A1(new_n9752_), .A2(pi0591), .B(new_n6352_), .ZN(new_n9781_));
  INV_X1     g07345(.I(new_n9781_), .ZN(new_n9782_));
  INV_X1     g07346(.I(new_n6546_), .ZN(new_n9783_));
  INV_X1     g07347(.I(pi0354), .ZN(new_n9784_));
  INV_X1     g07348(.I(pi0356), .ZN(new_n9785_));
  NAND3_X1   g07349(.A1(new_n6529_), .A2(new_n6381_), .A3(new_n9749_), .ZN(new_n9786_));
  NOR2_X1    g07350(.A1(new_n9786_), .A2(new_n6534_), .ZN(new_n9787_));
  NOR2_X1    g07351(.A1(new_n9787_), .A2(new_n9762_), .ZN(new_n9788_));
  NOR2_X1    g07352(.A1(new_n9786_), .A2(new_n6444_), .ZN(new_n9789_));
  NOR2_X1    g07353(.A1(new_n9789_), .A2(new_n9762_), .ZN(new_n9790_));
  AOI22_X1   g07354(.A1(new_n6442_), .A2(new_n9788_), .B1(new_n9790_), .B2(new_n6533_), .ZN(new_n9791_));
  NOR2_X1    g07355(.A1(new_n9791_), .A2(new_n9785_), .ZN(new_n9792_));
  NAND2_X1   g07356(.A1(new_n9790_), .A2(new_n6442_), .ZN(new_n9793_));
  NAND2_X1   g07357(.A1(new_n9788_), .A2(new_n6533_), .ZN(new_n9794_));
  NAND2_X1   g07358(.A1(new_n9793_), .A2(new_n9794_), .ZN(new_n9795_));
  AOI21_X1   g07359(.A1(new_n9785_), .A2(new_n9795_), .B(new_n9792_), .ZN(new_n9796_));
  NAND2_X1   g07360(.A1(new_n9796_), .A2(new_n9784_), .ZN(new_n9797_));
  NAND2_X1   g07361(.A1(new_n9795_), .A2(pi0356), .ZN(new_n9798_));
  OAI21_X1   g07362(.A1(pi0356), .A2(new_n9791_), .B(new_n9798_), .ZN(new_n9799_));
  OR2_X2     g07363(.A1(new_n9799_), .A2(new_n9784_), .Z(new_n9800_));
  AOI21_X1   g07364(.A1(new_n9800_), .A2(new_n9797_), .B(new_n9783_), .ZN(new_n9801_));
  AND2_X2    g07365(.A1(new_n9796_), .A2(pi0354), .Z(new_n9802_));
  NOR2_X1    g07366(.A1(new_n9799_), .A2(pi0354), .ZN(new_n9803_));
  OAI21_X1   g07367(.A1(new_n9802_), .A2(new_n9803_), .B(new_n9783_), .ZN(new_n9804_));
  NAND2_X1   g07368(.A1(new_n9804_), .A2(new_n6440_), .ZN(new_n9805_));
  NOR2_X1    g07369(.A1(new_n9805_), .A2(new_n9801_), .ZN(new_n9806_));
  NAND2_X1   g07370(.A1(new_n6614_), .A2(new_n6274_), .ZN(new_n9807_));
  NAND2_X1   g07371(.A1(pi0592), .A2(pi1198), .ZN(new_n9808_));
  AOI21_X1   g07372(.A1(new_n9807_), .A2(new_n9808_), .B(new_n6269_), .ZN(new_n9809_));
  AOI21_X1   g07373(.A1(new_n6638_), .A2(new_n9809_), .B(new_n9752_), .ZN(new_n9810_));
  OAI21_X1   g07374(.A1(new_n9810_), .A2(pi0591), .B(new_n6352_), .ZN(new_n9811_));
  XOR2_X1    g07375(.A1(new_n6364_), .A2(pi0392), .Z(new_n9812_));
  NOR3_X1    g07376(.A1(new_n6924_), .A2(new_n6271_), .A3(new_n9752_), .ZN(new_n9813_));
  NOR2_X1    g07377(.A1(new_n6960_), .A2(new_n6259_), .ZN(new_n9814_));
  NOR2_X1    g07378(.A1(new_n9814_), .A2(pi0122), .ZN(new_n9815_));
  INV_X1     g07379(.I(new_n9747_), .ZN(new_n9816_));
  NOR2_X1    g07380(.A1(new_n9816_), .A2(new_n3022_), .ZN(new_n9817_));
  INV_X1     g07381(.I(new_n9817_), .ZN(new_n9818_));
  AOI22_X1   g07382(.A1(new_n9815_), .A2(new_n9746_), .B1(new_n6871_), .B2(new_n9818_), .ZN(new_n9819_));
  INV_X1     g07383(.I(new_n9819_), .ZN(new_n9820_));
  NOR2_X1    g07384(.A1(new_n6259_), .A2(pi0122), .ZN(new_n9821_));
  INV_X1     g07385(.I(new_n9821_), .ZN(new_n9822_));
  AOI21_X1   g07386(.A1(new_n9746_), .A2(new_n9822_), .B(new_n9820_), .ZN(new_n9823_));
  NAND2_X1   g07387(.A1(new_n3043_), .A2(new_n6255_), .ZN(new_n9824_));
  OAI21_X1   g07388(.A1(new_n9823_), .A2(new_n6255_), .B(new_n9824_), .ZN(new_n9825_));
  NAND2_X1   g07389(.A1(new_n9752_), .A2(pi0592), .ZN(new_n9826_));
  OAI21_X1   g07390(.A1(new_n9825_), .A2(new_n6961_), .B(new_n9826_), .ZN(new_n9827_));
  NOR2_X1    g07391(.A1(pi0404), .A2(pi0411), .ZN(new_n9828_));
  INV_X1     g07392(.I(pi0404), .ZN(new_n9829_));
  NOR2_X1    g07393(.A1(new_n9829_), .A2(new_n6382_), .ZN(new_n9830_));
  OAI21_X1   g07394(.A1(new_n9830_), .A2(new_n9828_), .B(pi0397), .ZN(new_n9831_));
  INV_X1     g07395(.I(pi0397), .ZN(new_n9832_));
  NOR2_X1    g07396(.A1(new_n6382_), .A2(pi0404), .ZN(new_n9833_));
  NOR2_X1    g07397(.A1(new_n9829_), .A2(pi0411), .ZN(new_n9834_));
  OAI21_X1   g07398(.A1(new_n9833_), .A2(new_n9834_), .B(new_n9832_), .ZN(new_n9835_));
  NAND2_X1   g07399(.A1(new_n9831_), .A2(new_n9835_), .ZN(new_n9836_));
  NOR2_X1    g07400(.A1(new_n9836_), .A2(new_n6396_), .ZN(new_n9837_));
  AOI21_X1   g07401(.A1(new_n6399_), .A2(new_n9836_), .B(new_n9837_), .ZN(new_n9838_));
  NAND2_X1   g07402(.A1(new_n9838_), .A2(new_n6258_), .ZN(new_n9839_));
  XOR2_X1    g07403(.A1(new_n6393_), .A2(pi0412), .Z(new_n9840_));
  AND3_X2    g07404(.A1(new_n9839_), .A2(new_n9746_), .A3(new_n9840_), .Z(new_n9841_));
  OAI21_X1   g07405(.A1(new_n9838_), .A2(new_n6259_), .B(new_n9746_), .ZN(new_n9842_));
  NOR2_X1    g07406(.A1(new_n9842_), .A2(new_n9840_), .ZN(new_n9843_));
  NOR3_X1    g07407(.A1(new_n9841_), .A2(new_n9843_), .A3(pi0122), .ZN(new_n9844_));
  INV_X1     g07408(.I(new_n9844_), .ZN(new_n9845_));
  AOI21_X1   g07409(.A1(new_n9845_), .A2(new_n9746_), .B(new_n6871_), .ZN(new_n9846_));
  NOR2_X1    g07410(.A1(new_n9846_), .A2(new_n9817_), .ZN(new_n9847_));
  INV_X1     g07411(.I(new_n9847_), .ZN(new_n9848_));
  NAND2_X1   g07412(.A1(new_n9848_), .A2(pi0567), .ZN(new_n9849_));
  AND2_X2    g07413(.A1(new_n9825_), .A2(new_n9849_), .Z(new_n9850_));
  NOR2_X1    g07414(.A1(new_n9850_), .A2(new_n6304_), .ZN(new_n9851_));
  NOR3_X1    g07415(.A1(new_n9851_), .A2(new_n6380_), .A3(new_n9827_), .ZN(new_n9852_));
  OAI21_X1   g07416(.A1(new_n9749_), .A2(new_n6303_), .B(new_n6380_), .ZN(new_n9853_));
  INV_X1     g07417(.I(new_n9748_), .ZN(new_n9854_));
  NAND2_X1   g07418(.A1(new_n9849_), .A2(new_n9854_), .ZN(new_n9855_));
  AOI21_X1   g07419(.A1(new_n9855_), .A2(new_n6303_), .B(new_n9853_), .ZN(new_n9856_));
  OR2_X2     g07420(.A1(new_n9852_), .A2(new_n9856_), .Z(new_n9857_));
  AOI21_X1   g07421(.A1(new_n9857_), .A2(new_n6924_), .B(new_n9813_), .ZN(new_n9858_));
  OR2_X2     g07422(.A1(new_n9858_), .A2(new_n6422_), .Z(new_n9859_));
  NOR2_X1    g07423(.A1(new_n7035_), .A2(pi1197), .ZN(new_n9860_));
  NOR3_X1    g07424(.A1(new_n9860_), .A2(new_n6271_), .A3(new_n9752_), .ZN(new_n9861_));
  AOI21_X1   g07425(.A1(new_n9857_), .A2(new_n9860_), .B(new_n9861_), .ZN(new_n9862_));
  OAI21_X1   g07426(.A1(pi0333), .A2(new_n9862_), .B(new_n9859_), .ZN(new_n9863_));
  NAND2_X1   g07427(.A1(new_n9863_), .A2(pi0391), .ZN(new_n9864_));
  INV_X1     g07428(.I(pi0391), .ZN(new_n9865_));
  OR2_X2     g07429(.A1(new_n9862_), .A2(new_n6422_), .Z(new_n9866_));
  OAI21_X1   g07430(.A1(pi0333), .A2(new_n9858_), .B(new_n9866_), .ZN(new_n9867_));
  NAND2_X1   g07431(.A1(new_n9867_), .A2(new_n9865_), .ZN(new_n9868_));
  AOI21_X1   g07432(.A1(new_n9864_), .A2(new_n9868_), .B(new_n9812_), .ZN(new_n9869_));
  INV_X1     g07433(.I(new_n9812_), .ZN(new_n9870_));
  NAND2_X1   g07434(.A1(new_n9867_), .A2(pi0391), .ZN(new_n9871_));
  NAND2_X1   g07435(.A1(new_n9863_), .A2(new_n9865_), .ZN(new_n9872_));
  AOI21_X1   g07436(.A1(new_n9871_), .A2(new_n9872_), .B(new_n9870_), .ZN(new_n9873_));
  NOR3_X1    g07437(.A1(new_n9869_), .A2(new_n9873_), .A3(new_n6440_), .ZN(new_n9874_));
  OAI22_X1   g07438(.A1(new_n9874_), .A2(new_n9811_), .B1(new_n9782_), .B2(new_n9806_), .ZN(new_n9875_));
  OAI21_X1   g07439(.A1(new_n9875_), .A2(pi0588), .B(new_n6350_), .ZN(new_n9876_));
  OAI21_X1   g07440(.A1(new_n9876_), .A2(new_n9780_), .B(new_n9754_), .ZN(new_n9877_));
  INV_X1     g07441(.I(pi0080), .ZN(new_n9878_));
  INV_X1     g07442(.I(new_n7048_), .ZN(new_n9879_));
  NOR2_X1    g07443(.A1(new_n9879_), .A2(new_n7227_), .ZN(new_n9880_));
  NOR2_X1    g07444(.A1(new_n7048_), .A2(new_n7231_), .ZN(new_n9881_));
  INV_X1     g07445(.I(pi0369), .ZN(new_n9882_));
  INV_X1     g07446(.I(new_n7052_), .ZN(new_n9883_));
  NOR2_X1    g07447(.A1(new_n9752_), .A2(new_n6645_), .ZN(new_n9884_));
  NAND2_X1   g07448(.A1(new_n9816_), .A2(pi0075), .ZN(new_n9885_));
  NOR2_X1    g07449(.A1(new_n2733_), .A2(new_n3130_), .ZN(new_n9886_));
  NOR2_X1    g07450(.A1(new_n6673_), .A2(new_n8423_), .ZN(new_n9887_));
  NAND4_X1   g07451(.A1(new_n2869_), .A2(new_n6669_), .A3(new_n9886_), .A4(new_n9887_), .ZN(new_n9888_));
  NAND2_X1   g07452(.A1(new_n2985_), .A2(pi0093), .ZN(new_n9889_));
  NAND2_X1   g07453(.A1(new_n2771_), .A2(pi0090), .ZN(new_n9890_));
  AOI21_X1   g07454(.A1(new_n9889_), .A2(new_n9890_), .B(new_n2761_), .ZN(new_n9891_));
  AOI22_X1   g07455(.A1(new_n9891_), .A2(new_n3179_), .B1(pi0051), .B2(new_n6678_), .ZN(new_n9892_));
  NOR2_X1    g07456(.A1(new_n5428_), .A2(new_n3045_), .ZN(new_n9893_));
  INV_X1     g07457(.I(new_n9893_), .ZN(new_n9894_));
  NOR4_X1    g07458(.A1(new_n9888_), .A2(new_n6685_), .A3(new_n9892_), .A4(new_n9894_), .ZN(new_n9895_));
  OAI21_X1   g07459(.A1(new_n9895_), .A2(pi0098), .B(pi1092), .ZN(new_n9896_));
  OAI21_X1   g07460(.A1(new_n9896_), .A2(new_n6871_), .B(new_n9818_), .ZN(new_n9897_));
  NAND2_X1   g07461(.A1(new_n9897_), .A2(new_n2658_), .ZN(new_n9898_));
  INV_X1     g07462(.I(new_n2529_), .ZN(new_n9899_));
  NOR4_X1    g07463(.A1(new_n9888_), .A2(new_n9899_), .A3(new_n6679_), .A4(new_n9894_), .ZN(new_n9900_));
  OAI21_X1   g07464(.A1(new_n9900_), .A2(pi0098), .B(pi1092), .ZN(new_n9901_));
  OAI21_X1   g07465(.A1(new_n9901_), .A2(new_n6871_), .B(new_n9818_), .ZN(new_n9902_));
  NAND2_X1   g07466(.A1(new_n9902_), .A2(new_n6802_), .ZN(new_n9903_));
  NAND2_X1   g07467(.A1(new_n9747_), .A2(new_n3273_), .ZN(new_n9904_));
  NAND4_X1   g07468(.A1(new_n9903_), .A2(new_n9898_), .A3(new_n3465_), .A4(new_n9904_), .ZN(new_n9905_));
  NAND3_X1   g07469(.A1(new_n9905_), .A2(pi0567), .A3(new_n9885_), .ZN(new_n9906_));
  NOR2_X1    g07470(.A1(new_n9748_), .A2(new_n6648_), .ZN(new_n9907_));
  AOI21_X1   g07471(.A1(new_n9906_), .A2(new_n9907_), .B(new_n9884_), .ZN(new_n9908_));
  NAND2_X1   g07472(.A1(new_n9749_), .A2(new_n6268_), .ZN(new_n9909_));
  OAI21_X1   g07473(.A1(new_n9908_), .A2(new_n6268_), .B(new_n9909_), .ZN(new_n9910_));
  AND2_X2    g07474(.A1(new_n9910_), .A2(new_n7052_), .Z(new_n9911_));
  INV_X1     g07475(.I(new_n6611_), .ZN(new_n9912_));
  NOR2_X1    g07476(.A1(new_n9912_), .A2(new_n9749_), .ZN(new_n9913_));
  INV_X1     g07477(.I(new_n9913_), .ZN(new_n9914_));
  OAI21_X1   g07478(.A1(new_n9910_), .A2(new_n6611_), .B(new_n9914_), .ZN(new_n9915_));
  AOI21_X1   g07479(.A1(new_n9910_), .A2(new_n6571_), .B(pi1199), .ZN(new_n9916_));
  MUX2_X1    g07480(.I0(new_n9749_), .I1(new_n9910_), .S(new_n6589_), .Z(new_n9917_));
  NOR2_X1    g07481(.A1(new_n9917_), .A2(new_n6273_), .ZN(new_n9918_));
  INV_X1     g07482(.I(new_n6571_), .ZN(new_n9919_));
  OAI21_X1   g07483(.A1(pi1197), .A2(new_n9749_), .B(new_n9919_), .ZN(new_n9920_));
  OR2_X2     g07484(.A1(new_n9918_), .A2(new_n9920_), .Z(new_n9921_));
  AOI22_X1   g07485(.A1(new_n9921_), .A2(new_n9916_), .B1(pi1199), .B2(new_n9915_), .ZN(new_n9922_));
  AOI21_X1   g07486(.A1(new_n9922_), .A2(new_n9883_), .B(new_n9911_), .ZN(new_n9923_));
  NOR2_X1    g07487(.A1(new_n9923_), .A2(new_n9882_), .ZN(new_n9924_));
  INV_X1     g07488(.I(new_n7071_), .ZN(new_n9925_));
  AND2_X2    g07489(.A1(new_n9910_), .A2(new_n7071_), .Z(new_n9926_));
  AOI21_X1   g07490(.A1(new_n9922_), .A2(new_n9925_), .B(new_n9926_), .ZN(new_n9927_));
  NOR2_X1    g07491(.A1(new_n9927_), .A2(pi0369), .ZN(new_n9928_));
  OAI22_X1   g07492(.A1(new_n9924_), .A2(new_n9928_), .B1(new_n9880_), .B2(new_n9881_), .ZN(new_n9929_));
  NOR2_X1    g07493(.A1(new_n9880_), .A2(new_n9881_), .ZN(new_n9930_));
  NOR2_X1    g07494(.A1(new_n9927_), .A2(new_n9882_), .ZN(new_n9931_));
  NOR2_X1    g07495(.A1(new_n9923_), .A2(pi0369), .ZN(new_n9932_));
  OAI21_X1   g07496(.A1(new_n9931_), .A2(new_n9932_), .B(new_n9930_), .ZN(new_n9933_));
  NAND3_X1   g07497(.A1(new_n9929_), .A2(new_n9933_), .A3(new_n6440_), .ZN(new_n9934_));
  INV_X1     g07498(.I(new_n6363_), .ZN(new_n9935_));
  INV_X1     g07499(.I(pi0392), .ZN(new_n9936_));
  XNOR2_X1   g07500(.A1(pi0333), .A2(pi0391), .ZN(new_n9937_));
  INV_X1     g07501(.I(new_n9907_), .ZN(new_n9938_));
  NOR2_X1    g07502(.A1(new_n9938_), .A2(new_n7170_), .ZN(new_n9939_));
  OAI21_X1   g07503(.A1(new_n9939_), .A2(new_n9749_), .B(pi1199), .ZN(new_n9940_));
  NOR2_X1    g07504(.A1(new_n6416_), .A2(new_n9745_), .ZN(new_n9941_));
  AOI21_X1   g07505(.A1(new_n9896_), .A2(new_n6416_), .B(new_n9941_), .ZN(new_n9942_));
  INV_X1     g07506(.I(new_n9942_), .ZN(new_n9943_));
  NOR2_X1    g07507(.A1(new_n9943_), .A2(new_n9898_), .ZN(new_n9944_));
  AOI21_X1   g07508(.A1(new_n9901_), .A2(new_n6416_), .B(new_n9941_), .ZN(new_n9945_));
  INV_X1     g07509(.I(new_n9945_), .ZN(new_n9946_));
  OAI21_X1   g07510(.A1(new_n9946_), .A2(new_n9903_), .B(new_n9904_), .ZN(new_n9947_));
  NOR2_X1    g07511(.A1(new_n9884_), .A2(new_n6961_), .ZN(new_n9948_));
  OAI21_X1   g07512(.A1(new_n9947_), .A2(new_n9944_), .B(new_n9948_), .ZN(new_n9949_));
  NOR2_X1    g07513(.A1(new_n9884_), .A2(new_n6304_), .ZN(new_n9950_));
  INV_X1     g07514(.I(new_n9950_), .ZN(new_n9951_));
  NOR2_X1    g07515(.A1(new_n6403_), .A2(new_n9746_), .ZN(new_n9952_));
  NOR2_X1    g07516(.A1(new_n6404_), .A2(new_n9896_), .ZN(new_n9953_));
  NOR2_X1    g07517(.A1(new_n9953_), .A2(new_n9952_), .ZN(new_n9954_));
  OAI21_X1   g07518(.A1(new_n9954_), .A2(new_n6871_), .B(new_n9818_), .ZN(new_n9955_));
  NAND2_X1   g07519(.A1(new_n9955_), .A2(new_n2658_), .ZN(new_n9956_));
  INV_X1     g07520(.I(new_n9901_), .ZN(new_n9957_));
  AOI21_X1   g07521(.A1(new_n6403_), .A2(new_n9957_), .B(new_n9952_), .ZN(new_n9958_));
  NOR2_X1    g07522(.A1(new_n9958_), .A2(new_n6871_), .ZN(new_n9959_));
  OAI21_X1   g07523(.A1(new_n9959_), .A2(new_n9817_), .B(new_n6802_), .ZN(new_n9960_));
  NAND3_X1   g07524(.A1(new_n9956_), .A2(new_n9960_), .A3(new_n9904_), .ZN(new_n9961_));
  NOR2_X1    g07525(.A1(new_n9903_), .A2(new_n6960_), .ZN(new_n9962_));
  NOR3_X1    g07526(.A1(new_n9961_), .A2(new_n9944_), .A3(new_n9962_), .ZN(new_n9963_));
  OAI21_X1   g07527(.A1(new_n9963_), .A2(new_n9951_), .B(new_n9949_), .ZN(new_n9964_));
  NOR2_X1    g07528(.A1(new_n6255_), .A2(pi0075), .ZN(new_n9965_));
  AOI21_X1   g07529(.A1(new_n9964_), .A2(new_n9965_), .B(new_n9940_), .ZN(new_n9966_));
  NAND4_X1   g07530(.A1(new_n9956_), .A2(new_n3465_), .A3(new_n9960_), .A4(new_n9904_), .ZN(new_n9967_));
  NAND3_X1   g07531(.A1(new_n9967_), .A2(pi0567), .A3(new_n9885_), .ZN(new_n9968_));
  NAND2_X1   g07532(.A1(new_n9968_), .A2(new_n9907_), .ZN(new_n9969_));
  AOI21_X1   g07533(.A1(new_n9969_), .A2(new_n9950_), .B(new_n9853_), .ZN(new_n9970_));
  NOR3_X1    g07534(.A1(new_n9966_), .A2(new_n9970_), .A3(new_n7035_), .ZN(new_n9971_));
  NAND2_X1   g07535(.A1(new_n9971_), .A2(new_n6273_), .ZN(new_n9972_));
  OR2_X2     g07536(.A1(new_n9908_), .A2(pi0592), .Z(new_n9973_));
  NOR2_X1    g07537(.A1(new_n9752_), .A2(new_n6268_), .ZN(new_n9974_));
  INV_X1     g07538(.I(new_n9974_), .ZN(new_n9975_));
  NAND2_X1   g07539(.A1(new_n9973_), .A2(new_n9975_), .ZN(new_n9976_));
  OAI21_X1   g07540(.A1(new_n9860_), .A2(new_n9976_), .B(new_n9972_), .ZN(new_n9977_));
  NOR2_X1    g07541(.A1(new_n9976_), .A2(new_n6924_), .ZN(new_n9978_));
  OR2_X2     g07542(.A1(new_n9971_), .A2(new_n9978_), .Z(new_n9979_));
  XOR2_X1    g07543(.A1(pi0333), .A2(pi0391), .Z(new_n9980_));
  OAI22_X1   g07544(.A1(new_n9977_), .A2(new_n9937_), .B1(new_n9979_), .B2(new_n9980_), .ZN(new_n9981_));
  AND2_X2    g07545(.A1(new_n9981_), .A2(pi0392), .Z(new_n9982_));
  OAI22_X1   g07546(.A1(new_n9977_), .A2(new_n9980_), .B1(new_n9937_), .B2(new_n9979_), .ZN(new_n9983_));
  AOI21_X1   g07547(.A1(new_n9936_), .A2(new_n9983_), .B(new_n9982_), .ZN(new_n9984_));
  NOR2_X1    g07548(.A1(new_n9984_), .A2(new_n7158_), .ZN(new_n9985_));
  AND2_X2    g07549(.A1(new_n9983_), .A2(pi0392), .Z(new_n9986_));
  AOI21_X1   g07550(.A1(new_n9936_), .A2(new_n9981_), .B(new_n9986_), .ZN(new_n9987_));
  NOR2_X1    g07551(.A1(new_n9987_), .A2(pi0393), .ZN(new_n9988_));
  OAI21_X1   g07552(.A1(new_n9985_), .A2(new_n9988_), .B(new_n9935_), .ZN(new_n9989_));
  NOR2_X1    g07553(.A1(new_n9987_), .A2(new_n7158_), .ZN(new_n9990_));
  NOR2_X1    g07554(.A1(new_n9984_), .A2(pi0393), .ZN(new_n9991_));
  OAI21_X1   g07555(.A1(new_n9990_), .A2(new_n9991_), .B(new_n6363_), .ZN(new_n9992_));
  NAND3_X1   g07556(.A1(new_n9989_), .A2(new_n9992_), .A3(pi0591), .ZN(new_n9993_));
  NAND3_X1   g07557(.A1(new_n9993_), .A2(new_n6352_), .A3(new_n9934_), .ZN(new_n9994_));
  INV_X1     g07558(.I(new_n9976_), .ZN(new_n9995_));
  NAND2_X1   g07559(.A1(new_n6516_), .A2(new_n9749_), .ZN(new_n9996_));
  NAND2_X1   g07560(.A1(new_n9976_), .A2(new_n6515_), .ZN(new_n9997_));
  AOI21_X1   g07561(.A1(new_n9997_), .A2(new_n9996_), .B(new_n6274_), .ZN(new_n9998_));
  OAI21_X1   g07562(.A1(new_n9749_), .A2(pi1196), .B(new_n6274_), .ZN(new_n9999_));
  INV_X1     g07563(.I(new_n6483_), .ZN(new_n10000_));
  INV_X1     g07564(.I(new_n6490_), .ZN(new_n10001_));
  INV_X1     g07565(.I(new_n7131_), .ZN(new_n10002_));
  AOI22_X1   g07566(.A1(new_n9976_), .A2(new_n10001_), .B1(new_n10002_), .B2(new_n9749_), .ZN(new_n10003_));
  NAND2_X1   g07567(.A1(new_n9752_), .A2(new_n10001_), .ZN(new_n10004_));
  OAI21_X1   g07568(.A1(new_n9976_), .A2(new_n10001_), .B(new_n10004_), .ZN(new_n10005_));
  AND2_X2    g07569(.A1(new_n10005_), .A2(pi0355), .Z(new_n10006_));
  AOI21_X1   g07570(.A1(new_n6485_), .A2(new_n10003_), .B(new_n10006_), .ZN(new_n10007_));
  AND2_X2    g07571(.A1(new_n10007_), .A2(pi0458), .Z(new_n10008_));
  NAND2_X1   g07572(.A1(new_n10003_), .A2(pi0355), .ZN(new_n10009_));
  NAND2_X1   g07573(.A1(new_n10005_), .A2(new_n6485_), .ZN(new_n10010_));
  NAND2_X1   g07574(.A1(new_n10009_), .A2(new_n10010_), .ZN(new_n10011_));
  NOR2_X1    g07575(.A1(new_n10011_), .A2(pi0458), .ZN(new_n10012_));
  OAI21_X1   g07576(.A1(new_n10008_), .A2(new_n10012_), .B(new_n10000_), .ZN(new_n10013_));
  NAND2_X1   g07577(.A1(new_n10007_), .A2(new_n7136_), .ZN(new_n10014_));
  OAI21_X1   g07578(.A1(new_n7136_), .A2(new_n10011_), .B(new_n10014_), .ZN(new_n10015_));
  AOI21_X1   g07579(.A1(new_n10015_), .A2(new_n6483_), .B(new_n6302_), .ZN(new_n10016_));
  AOI21_X1   g07580(.A1(new_n10016_), .A2(new_n10013_), .B(new_n9999_), .ZN(new_n10017_));
  NOR3_X1    g07581(.A1(new_n10017_), .A2(new_n6467_), .A3(new_n9998_), .ZN(new_n10018_));
  AOI21_X1   g07582(.A1(new_n6467_), .A2(new_n9995_), .B(new_n10018_), .ZN(new_n10019_));
  INV_X1     g07583(.I(new_n10019_), .ZN(new_n10020_));
  NOR2_X1    g07584(.A1(new_n10020_), .A2(new_n6444_), .ZN(new_n10021_));
  AOI21_X1   g07585(.A1(new_n6444_), .A2(new_n9976_), .B(new_n10021_), .ZN(new_n10022_));
  INV_X1     g07586(.I(new_n10022_), .ZN(new_n10023_));
  NOR2_X1    g07587(.A1(new_n10020_), .A2(new_n6534_), .ZN(new_n10024_));
  AOI21_X1   g07588(.A1(new_n6534_), .A2(new_n9976_), .B(new_n10024_), .ZN(new_n10025_));
  INV_X1     g07589(.I(new_n10025_), .ZN(new_n10026_));
  AOI22_X1   g07590(.A1(new_n6442_), .A2(new_n10023_), .B1(new_n10026_), .B2(new_n6533_), .ZN(new_n10027_));
  NOR2_X1    g07591(.A1(new_n10027_), .A2(new_n9785_), .ZN(new_n10028_));
  AOI22_X1   g07592(.A1(new_n6442_), .A2(new_n10026_), .B1(new_n10023_), .B2(new_n6533_), .ZN(new_n10029_));
  NOR2_X1    g07593(.A1(new_n10029_), .A2(pi0356), .ZN(new_n10030_));
  OAI21_X1   g07594(.A1(new_n10028_), .A2(new_n10030_), .B(pi0354), .ZN(new_n10031_));
  NOR2_X1    g07595(.A1(new_n10029_), .A2(new_n9785_), .ZN(new_n10032_));
  NOR2_X1    g07596(.A1(new_n10027_), .A2(pi0356), .ZN(new_n10033_));
  OAI21_X1   g07597(.A1(new_n10032_), .A2(new_n10033_), .B(new_n9784_), .ZN(new_n10034_));
  AOI21_X1   g07598(.A1(new_n10031_), .A2(new_n10034_), .B(new_n9783_), .ZN(new_n10035_));
  NOR2_X1    g07599(.A1(new_n10032_), .A2(new_n10033_), .ZN(new_n10036_));
  NOR2_X1    g07600(.A1(new_n10036_), .A2(new_n9784_), .ZN(new_n10037_));
  NOR2_X1    g07601(.A1(new_n10028_), .A2(new_n10030_), .ZN(new_n10038_));
  NOR2_X1    g07602(.A1(new_n10038_), .A2(pi0354), .ZN(new_n10039_));
  OAI21_X1   g07603(.A1(new_n10039_), .A2(new_n10037_), .B(new_n9783_), .ZN(new_n10040_));
  NAND2_X1   g07604(.A1(new_n10040_), .A2(new_n6440_), .ZN(new_n10041_));
  OAI21_X1   g07605(.A1(new_n10041_), .A2(new_n10035_), .B(new_n9781_), .ZN(new_n10042_));
  NAND3_X1   g07606(.A1(new_n10042_), .A2(new_n6251_), .A3(new_n9994_), .ZN(new_n10043_));
  NAND2_X1   g07607(.A1(new_n9976_), .A2(new_n6301_), .ZN(new_n10044_));
  INV_X1     g07608(.I(pi0435), .ZN(new_n10045_));
  NOR2_X1    g07609(.A1(new_n9752_), .A2(pi0443), .ZN(new_n10046_));
  AOI21_X1   g07610(.A1(new_n9976_), .A2(pi0443), .B(new_n10046_), .ZN(new_n10047_));
  INV_X1     g07611(.I(new_n10047_), .ZN(new_n10048_));
  XOR2_X1    g07612(.A1(pi0436), .A2(pi0444), .Z(new_n10049_));
  INV_X1     g07613(.I(pi0443), .ZN(new_n10050_));
  NOR2_X1    g07614(.A1(new_n9752_), .A2(new_n10050_), .ZN(new_n10051_));
  INV_X1     g07615(.I(new_n10051_), .ZN(new_n10052_));
  OAI21_X1   g07616(.A1(new_n9995_), .A2(pi0443), .B(new_n10052_), .ZN(new_n10053_));
  AOI22_X1   g07617(.A1(new_n10048_), .A2(new_n10049_), .B1(new_n10053_), .B2(new_n6830_), .ZN(new_n10054_));
  NAND2_X1   g07618(.A1(new_n10054_), .A2(new_n10045_), .ZN(new_n10055_));
  NAND2_X1   g07619(.A1(new_n10047_), .A2(new_n6830_), .ZN(new_n10056_));
  OAI21_X1   g07620(.A1(new_n6830_), .A2(new_n10053_), .B(new_n10056_), .ZN(new_n10057_));
  NAND2_X1   g07621(.A1(new_n10057_), .A2(pi0435), .ZN(new_n10058_));
  INV_X1     g07622(.I(pi0429), .ZN(new_n10059_));
  XOR2_X1    g07623(.A1(new_n6315_), .A2(new_n10059_), .Z(new_n10060_));
  NAND3_X1   g07624(.A1(new_n10055_), .A2(new_n10058_), .A3(new_n10060_), .ZN(new_n10061_));
  INV_X1     g07625(.I(new_n10060_), .ZN(new_n10062_));
  NAND2_X1   g07626(.A1(new_n10054_), .A2(pi0435), .ZN(new_n10063_));
  NAND2_X1   g07627(.A1(new_n10057_), .A2(new_n10045_), .ZN(new_n10064_));
  NAND3_X1   g07628(.A1(new_n10063_), .A2(new_n10064_), .A3(new_n10062_), .ZN(new_n10065_));
  NAND3_X1   g07629(.A1(new_n10061_), .A2(new_n10065_), .A3(pi1196), .ZN(new_n10066_));
  NOR2_X1    g07630(.A1(new_n9749_), .A2(pi1196), .ZN(new_n10067_));
  NOR2_X1    g07631(.A1(new_n6301_), .A2(new_n10067_), .ZN(new_n10068_));
  NAND2_X1   g07632(.A1(new_n10066_), .A2(new_n10068_), .ZN(new_n10069_));
  NAND2_X1   g07633(.A1(new_n10069_), .A2(new_n10044_), .ZN(new_n10070_));
  OAI21_X1   g07634(.A1(new_n10070_), .A2(pi1199), .B(new_n6253_), .ZN(new_n10071_));
  NOR2_X1    g07635(.A1(new_n10070_), .A2(new_n6850_), .ZN(new_n10072_));
  AOI21_X1   g07636(.A1(new_n6849_), .A2(new_n9995_), .B(new_n10072_), .ZN(new_n10073_));
  NOR2_X1    g07637(.A1(new_n10070_), .A2(new_n6848_), .ZN(new_n10074_));
  AOI21_X1   g07638(.A1(new_n6851_), .A2(new_n9995_), .B(new_n10074_), .ZN(new_n10075_));
  OAI22_X1   g07639(.A1(new_n6853_), .A2(new_n10075_), .B1(new_n10073_), .B2(new_n6856_), .ZN(new_n10076_));
  AND2_X2    g07640(.A1(new_n10076_), .A2(pi0445), .Z(new_n10077_));
  OAI22_X1   g07641(.A1(new_n6853_), .A2(new_n10073_), .B1(new_n10075_), .B2(new_n6856_), .ZN(new_n10078_));
  AOI21_X1   g07642(.A1(new_n6859_), .A2(new_n10078_), .B(new_n10077_), .ZN(new_n10079_));
  NAND2_X1   g07643(.A1(new_n10079_), .A2(new_n9760_), .ZN(new_n10080_));
  AND2_X2    g07644(.A1(new_n10078_), .A2(pi0445), .Z(new_n10081_));
  AOI21_X1   g07645(.A1(new_n6859_), .A2(new_n10076_), .B(new_n10081_), .ZN(new_n10082_));
  NAND2_X1   g07646(.A1(new_n10082_), .A2(pi0448), .ZN(new_n10083_));
  AOI21_X1   g07647(.A1(new_n10080_), .A2(new_n10083_), .B(new_n6331_), .ZN(new_n10084_));
  NAND2_X1   g07648(.A1(new_n10079_), .A2(pi0448), .ZN(new_n10085_));
  NAND2_X1   g07649(.A1(new_n10082_), .A2(new_n9760_), .ZN(new_n10086_));
  AOI21_X1   g07650(.A1(new_n10085_), .A2(new_n10086_), .B(new_n9759_), .ZN(new_n10087_));
  NOR3_X1    g07651(.A1(new_n10084_), .A2(new_n10087_), .A3(new_n6380_), .ZN(new_n10088_));
  OAI21_X1   g07652(.A1(new_n10088_), .A2(new_n10071_), .B(new_n9778_), .ZN(new_n10089_));
  NAND3_X1   g07653(.A1(new_n10043_), .A2(new_n6349_), .A3(new_n10089_), .ZN(new_n10090_));
  NOR2_X1    g07654(.A1(new_n6259_), .A2(new_n6257_), .ZN(new_n10091_));
  INV_X1     g07655(.I(new_n10091_), .ZN(new_n10092_));
  NOR2_X1    g07656(.A1(new_n10092_), .A2(pi1091), .ZN(new_n10093_));
  NOR2_X1    g07657(.A1(new_n10093_), .A2(new_n9747_), .ZN(new_n10094_));
  OAI21_X1   g07658(.A1(new_n10094_), .A2(new_n6645_), .B(new_n9854_), .ZN(new_n10095_));
  NOR2_X1    g07659(.A1(new_n6648_), .A2(new_n6255_), .ZN(new_n10096_));
  NAND2_X1   g07660(.A1(new_n10094_), .A2(new_n6650_), .ZN(new_n10097_));
  NAND2_X1   g07661(.A1(new_n10097_), .A2(new_n10096_), .ZN(new_n10098_));
  NOR2_X1    g07662(.A1(new_n9817_), .A2(new_n3273_), .ZN(new_n10099_));
  INV_X1     g07663(.I(new_n10099_), .ZN(new_n10100_));
  AOI21_X1   g07664(.A1(new_n10094_), .A2(new_n6714_), .B(new_n6871_), .ZN(new_n10101_));
  AND2_X2    g07665(.A1(new_n9896_), .A2(new_n3458_), .Z(new_n10102_));
  NOR2_X1    g07666(.A1(new_n9957_), .A2(new_n3458_), .ZN(new_n10103_));
  OAI21_X1   g07667(.A1(new_n10103_), .A2(new_n10102_), .B(pi0122), .ZN(new_n10104_));
  AOI21_X1   g07668(.A1(new_n10104_), .A2(new_n10101_), .B(new_n10100_), .ZN(new_n10105_));
  AOI21_X1   g07669(.A1(new_n10105_), .A2(new_n3465_), .B(new_n10098_), .ZN(new_n10106_));
  NOR2_X1    g07670(.A1(new_n10106_), .A2(new_n10095_), .ZN(new_n10107_));
  NAND2_X1   g07671(.A1(new_n10107_), .A2(pi0592), .ZN(new_n10108_));
  NAND2_X1   g07672(.A1(new_n10108_), .A2(new_n9909_), .ZN(new_n10109_));
  OAI22_X1   g07673(.A1(new_n10109_), .A2(new_n6586_), .B1(new_n6585_), .B2(new_n9749_), .ZN(new_n10110_));
  NOR2_X1    g07674(.A1(new_n10110_), .A2(new_n6572_), .ZN(new_n10111_));
  INV_X1     g07675(.I(new_n10109_), .ZN(new_n10112_));
  OAI22_X1   g07676(.A1(new_n10112_), .A2(new_n6585_), .B1(new_n6586_), .B2(new_n9752_), .ZN(new_n10113_));
  AND2_X2    g07677(.A1(new_n10113_), .A2(new_n6572_), .Z(new_n10114_));
  OAI21_X1   g07678(.A1(new_n10114_), .A2(new_n10111_), .B(new_n6581_), .ZN(new_n10115_));
  INV_X1     g07679(.I(new_n6581_), .ZN(new_n10116_));
  INV_X1     g07680(.I(new_n6572_), .ZN(new_n10117_));
  NAND2_X1   g07681(.A1(new_n10113_), .A2(new_n10117_), .ZN(new_n10118_));
  OAI21_X1   g07682(.A1(new_n10117_), .A2(new_n10110_), .B(new_n10118_), .ZN(new_n10119_));
  AOI21_X1   g07683(.A1(new_n10119_), .A2(new_n10116_), .B(new_n6273_), .ZN(new_n10120_));
  AOI21_X1   g07684(.A1(new_n10120_), .A2(new_n10115_), .B(new_n9920_), .ZN(new_n10121_));
  OAI21_X1   g07685(.A1(new_n10112_), .A2(new_n9919_), .B(new_n6380_), .ZN(new_n10122_));
  AOI21_X1   g07686(.A1(new_n10112_), .A2(new_n9912_), .B(new_n9913_), .ZN(new_n10123_));
  OAI22_X1   g07687(.A1(new_n10121_), .A2(new_n10122_), .B1(new_n6380_), .B2(new_n10123_), .ZN(new_n10124_));
  NOR2_X1    g07688(.A1(new_n10124_), .A2(new_n7051_), .ZN(new_n10125_));
  OAI22_X1   g07689(.A1(new_n10123_), .A2(new_n7219_), .B1(new_n6274_), .B2(new_n10109_), .ZN(new_n10126_));
  NOR3_X1    g07690(.A1(new_n10121_), .A2(pi1198), .A3(new_n10122_), .ZN(new_n10127_));
  OR2_X2     g07691(.A1(new_n10127_), .A2(new_n10126_), .Z(new_n10128_));
  NOR2_X1    g07692(.A1(new_n10128_), .A2(pi0374), .ZN(new_n10129_));
  XOR2_X1    g07693(.A1(new_n9930_), .A2(new_n9882_), .Z(new_n10130_));
  INV_X1     g07694(.I(new_n10130_), .ZN(new_n10131_));
  NOR3_X1    g07695(.A1(new_n10129_), .A2(new_n10125_), .A3(new_n10131_), .ZN(new_n10132_));
  NOR2_X1    g07696(.A1(new_n10128_), .A2(new_n7051_), .ZN(new_n10133_));
  NOR2_X1    g07697(.A1(new_n10124_), .A2(pi0374), .ZN(new_n10134_));
  NOR3_X1    g07698(.A1(new_n10133_), .A2(new_n10130_), .A3(new_n10134_), .ZN(new_n10135_));
  OAI21_X1   g07699(.A1(new_n10132_), .A2(new_n10135_), .B(new_n6440_), .ZN(new_n10136_));
  NAND2_X1   g07700(.A1(new_n10107_), .A2(new_n6268_), .ZN(new_n10137_));
  NAND2_X1   g07701(.A1(new_n10137_), .A2(new_n9975_), .ZN(new_n10138_));
  INV_X1     g07702(.I(new_n10138_), .ZN(new_n10139_));
  NOR2_X1    g07703(.A1(new_n10139_), .A2(new_n6924_), .ZN(new_n10140_));
  NOR2_X1    g07704(.A1(new_n9823_), .A2(new_n6649_), .ZN(new_n10141_));
  NAND2_X1   g07705(.A1(new_n9820_), .A2(new_n3272_), .ZN(new_n10142_));
  NAND2_X1   g07706(.A1(new_n10099_), .A2(new_n3458_), .ZN(new_n10143_));
  NOR2_X1    g07707(.A1(new_n10100_), .A2(new_n3458_), .ZN(new_n10144_));
  INV_X1     g07708(.I(new_n10144_), .ZN(new_n10145_));
  OAI22_X1   g07709(.A1(new_n9942_), .A2(new_n10143_), .B1(new_n9945_), .B2(new_n10145_), .ZN(new_n10146_));
  NAND2_X1   g07710(.A1(new_n10146_), .A2(pi0122), .ZN(new_n10147_));
  AOI21_X1   g07711(.A1(new_n10142_), .A2(new_n10147_), .B(pi0075), .ZN(new_n10148_));
  NOR4_X1    g07712(.A1(new_n10141_), .A2(new_n6255_), .A3(new_n10148_), .A4(new_n6648_), .ZN(new_n10149_));
  NOR2_X1    g07713(.A1(new_n9825_), .A2(new_n9907_), .ZN(new_n10150_));
  OAI21_X1   g07714(.A1(new_n10149_), .A2(new_n10150_), .B(new_n6302_), .ZN(new_n10151_));
  NOR2_X1    g07715(.A1(new_n9850_), .A2(new_n9907_), .ZN(new_n10152_));
  AOI21_X1   g07716(.A1(new_n9814_), .A2(new_n6714_), .B(new_n9844_), .ZN(new_n10153_));
  NAND2_X1   g07717(.A1(new_n6416_), .A2(new_n9957_), .ZN(new_n10154_));
  AND3_X2    g07718(.A1(new_n9958_), .A2(new_n10144_), .A3(new_n10154_), .Z(new_n10155_));
  NOR3_X1    g07719(.A1(new_n6400_), .A2(pi0411), .A3(new_n9746_), .ZN(new_n10156_));
  NOR4_X1    g07720(.A1(new_n9953_), .A2(new_n9942_), .A3(new_n10143_), .A4(new_n10156_), .ZN(new_n10157_));
  OAI21_X1   g07721(.A1(new_n10155_), .A2(new_n10157_), .B(new_n10153_), .ZN(new_n10158_));
  OAI21_X1   g07722(.A1(new_n9846_), .A2(new_n10142_), .B(new_n10158_), .ZN(new_n10159_));
  INV_X1     g07723(.I(new_n10141_), .ZN(new_n10160_));
  OAI21_X1   g07724(.A1(new_n10160_), .A2(new_n9846_), .B(new_n10096_), .ZN(new_n10161_));
  AOI21_X1   g07725(.A1(new_n10159_), .A2(new_n3465_), .B(new_n10161_), .ZN(new_n10162_));
  OAI21_X1   g07726(.A1(new_n10162_), .A2(new_n10152_), .B(pi1196), .ZN(new_n10163_));
  NAND2_X1   g07727(.A1(new_n10163_), .A2(new_n10151_), .ZN(new_n10164_));
  NAND3_X1   g07728(.A1(new_n10164_), .A2(new_n6268_), .A3(pi1199), .ZN(new_n10165_));
  NOR2_X1    g07729(.A1(new_n9847_), .A2(new_n3465_), .ZN(new_n10166_));
  NOR2_X1    g07730(.A1(new_n9848_), .A2(new_n3272_), .ZN(new_n10167_));
  OAI21_X1   g07731(.A1(new_n9958_), .A2(new_n6714_), .B(new_n9845_), .ZN(new_n10168_));
  AOI21_X1   g07732(.A1(new_n10168_), .A2(new_n6870_), .B(new_n10145_), .ZN(new_n10169_));
  OAI21_X1   g07733(.A1(new_n9954_), .A2(new_n6714_), .B(new_n9845_), .ZN(new_n10170_));
  AOI21_X1   g07734(.A1(new_n10170_), .A2(new_n6870_), .B(new_n10143_), .ZN(new_n10171_));
  NOR4_X1    g07735(.A1(new_n10171_), .A2(pi0075), .A3(new_n10169_), .A4(new_n10167_), .ZN(new_n10172_));
  OAI21_X1   g07736(.A1(new_n10172_), .A2(new_n10166_), .B(new_n10096_), .ZN(new_n10173_));
  NAND2_X1   g07737(.A1(new_n9855_), .A2(new_n9938_), .ZN(new_n10174_));
  AOI21_X1   g07738(.A1(new_n10173_), .A2(new_n10174_), .B(new_n6304_), .ZN(new_n10175_));
  OAI21_X1   g07739(.A1(new_n10175_), .A2(new_n10067_), .B(new_n6380_), .ZN(new_n10176_));
  AND3_X2    g07740(.A1(new_n10165_), .A2(new_n9826_), .A3(new_n10176_), .Z(new_n10177_));
  AOI21_X1   g07741(.A1(new_n10177_), .A2(new_n6924_), .B(new_n10140_), .ZN(new_n10178_));
  INV_X1     g07742(.I(new_n9860_), .ZN(new_n10179_));
  NAND2_X1   g07743(.A1(new_n10139_), .A2(new_n10179_), .ZN(new_n10180_));
  OAI21_X1   g07744(.A1(new_n10177_), .A2(new_n10179_), .B(new_n10180_), .ZN(new_n10181_));
  OAI22_X1   g07745(.A1(new_n9980_), .A2(new_n10178_), .B1(new_n10181_), .B2(new_n9937_), .ZN(new_n10182_));
  XOR2_X1    g07746(.A1(pi0392), .A2(pi0393), .Z(new_n10183_));
  INV_X1     g07747(.I(new_n9937_), .ZN(new_n10184_));
  INV_X1     g07748(.I(new_n9980_), .ZN(new_n10185_));
  AOI22_X1   g07749(.A1(new_n10184_), .A2(new_n10178_), .B1(new_n10181_), .B2(new_n10185_), .ZN(new_n10186_));
  XNOR2_X1   g07750(.A1(pi0392), .A2(pi0393), .ZN(new_n10187_));
  OAI22_X1   g07751(.A1(new_n10182_), .A2(new_n10183_), .B1(new_n10186_), .B2(new_n10187_), .ZN(new_n10188_));
  NAND2_X1   g07752(.A1(new_n10188_), .A2(new_n9935_), .ZN(new_n10189_));
  OAI22_X1   g07753(.A1(new_n10182_), .A2(new_n10187_), .B1(new_n10186_), .B2(new_n10183_), .ZN(new_n10190_));
  NAND2_X1   g07754(.A1(new_n10190_), .A2(new_n6363_), .ZN(new_n10191_));
  NAND2_X1   g07755(.A1(new_n10189_), .A2(new_n10191_), .ZN(new_n10192_));
  AOI21_X1   g07756(.A1(new_n10192_), .A2(pi0591), .B(pi0590), .ZN(new_n10193_));
  AOI21_X1   g07757(.A1(new_n10193_), .A2(new_n10136_), .B(pi0588), .ZN(new_n10194_));
  NAND2_X1   g07758(.A1(new_n10138_), .A2(new_n6515_), .ZN(new_n10195_));
  AOI21_X1   g07759(.A1(new_n10195_), .A2(new_n9996_), .B(new_n6274_), .ZN(new_n10196_));
  OAI22_X1   g07760(.A1(new_n10139_), .A2(new_n6490_), .B1(new_n7131_), .B2(new_n9752_), .ZN(new_n10197_));
  NOR2_X1    g07761(.A1(new_n10197_), .A2(new_n6485_), .ZN(new_n10198_));
  OAI21_X1   g07762(.A1(new_n10138_), .A2(new_n10001_), .B(new_n10004_), .ZN(new_n10199_));
  AOI21_X1   g07763(.A1(new_n6485_), .A2(new_n10199_), .B(new_n10198_), .ZN(new_n10200_));
  AND2_X2    g07764(.A1(new_n10200_), .A2(pi0458), .Z(new_n10201_));
  NAND2_X1   g07765(.A1(new_n10199_), .A2(pi0355), .ZN(new_n10202_));
  OAI21_X1   g07766(.A1(pi0355), .A2(new_n10197_), .B(new_n10202_), .ZN(new_n10203_));
  NOR2_X1    g07767(.A1(new_n10203_), .A2(pi0458), .ZN(new_n10204_));
  OAI21_X1   g07768(.A1(new_n10201_), .A2(new_n10204_), .B(new_n6483_), .ZN(new_n10205_));
  NAND2_X1   g07769(.A1(new_n10200_), .A2(new_n7136_), .ZN(new_n10206_));
  OAI21_X1   g07770(.A1(new_n7136_), .A2(new_n10203_), .B(new_n10206_), .ZN(new_n10207_));
  AOI21_X1   g07771(.A1(new_n10207_), .A2(new_n10000_), .B(new_n6302_), .ZN(new_n10208_));
  AND2_X2    g07772(.A1(new_n10208_), .A2(new_n10205_), .Z(new_n10209_));
  OAI21_X1   g07773(.A1(new_n10209_), .A2(new_n9999_), .B(new_n7085_), .ZN(new_n10210_));
  OAI22_X1   g07774(.A1(new_n10210_), .A2(new_n10196_), .B1(new_n7085_), .B2(new_n10138_), .ZN(new_n10211_));
  NAND2_X1   g07775(.A1(new_n10138_), .A2(new_n6444_), .ZN(new_n10212_));
  OAI21_X1   g07776(.A1(new_n10211_), .A2(new_n6444_), .B(new_n10212_), .ZN(new_n10213_));
  NAND2_X1   g07777(.A1(new_n10138_), .A2(new_n6534_), .ZN(new_n10214_));
  OAI21_X1   g07778(.A1(new_n10211_), .A2(new_n6534_), .B(new_n10214_), .ZN(new_n10215_));
  AOI22_X1   g07779(.A1(new_n6442_), .A2(new_n10213_), .B1(new_n10215_), .B2(new_n6533_), .ZN(new_n10216_));
  OR2_X2     g07780(.A1(new_n10216_), .A2(new_n9785_), .Z(new_n10217_));
  AOI22_X1   g07781(.A1(new_n6442_), .A2(new_n10215_), .B1(new_n10213_), .B2(new_n6533_), .ZN(new_n10218_));
  OAI21_X1   g07782(.A1(pi0356), .A2(new_n10218_), .B(new_n10217_), .ZN(new_n10219_));
  NAND2_X1   g07783(.A1(new_n10219_), .A2(pi0354), .ZN(new_n10220_));
  OR2_X2     g07784(.A1(new_n10218_), .A2(new_n9785_), .Z(new_n10221_));
  OAI21_X1   g07785(.A1(pi0356), .A2(new_n10216_), .B(new_n10221_), .ZN(new_n10222_));
  NAND2_X1   g07786(.A1(new_n10222_), .A2(new_n9784_), .ZN(new_n10223_));
  AOI21_X1   g07787(.A1(new_n10220_), .A2(new_n10223_), .B(new_n9783_), .ZN(new_n10224_));
  NAND2_X1   g07788(.A1(new_n10222_), .A2(pi0354), .ZN(new_n10225_));
  NAND2_X1   g07789(.A1(new_n10219_), .A2(new_n9784_), .ZN(new_n10226_));
  AOI21_X1   g07790(.A1(new_n10225_), .A2(new_n10226_), .B(new_n6546_), .ZN(new_n10227_));
  NOR3_X1    g07791(.A1(new_n10224_), .A2(new_n10227_), .A3(pi0591), .ZN(new_n10228_));
  OAI21_X1   g07792(.A1(new_n10228_), .A2(new_n9782_), .B(new_n10194_), .ZN(new_n10229_));
  NAND2_X1   g07793(.A1(new_n10138_), .A2(new_n6301_), .ZN(new_n10230_));
  AOI21_X1   g07794(.A1(new_n10138_), .A2(pi0443), .B(new_n10046_), .ZN(new_n10231_));
  INV_X1     g07795(.I(new_n10231_), .ZN(new_n10232_));
  AOI21_X1   g07796(.A1(new_n10138_), .A2(new_n10050_), .B(new_n10051_), .ZN(new_n10233_));
  INV_X1     g07797(.I(new_n10233_), .ZN(new_n10234_));
  AOI22_X1   g07798(.A1(new_n6830_), .A2(new_n10234_), .B1(new_n10232_), .B2(new_n10049_), .ZN(new_n10235_));
  NAND2_X1   g07799(.A1(new_n10235_), .A2(new_n10045_), .ZN(new_n10236_));
  NAND2_X1   g07800(.A1(new_n10231_), .A2(new_n6830_), .ZN(new_n10237_));
  OAI21_X1   g07801(.A1(new_n6830_), .A2(new_n10234_), .B(new_n10237_), .ZN(new_n10238_));
  NAND2_X1   g07802(.A1(new_n10238_), .A2(pi0435), .ZN(new_n10239_));
  NAND3_X1   g07803(.A1(new_n10236_), .A2(new_n10239_), .A3(new_n10060_), .ZN(new_n10240_));
  NAND2_X1   g07804(.A1(new_n10235_), .A2(pi0435), .ZN(new_n10241_));
  NAND2_X1   g07805(.A1(new_n10238_), .A2(new_n10045_), .ZN(new_n10242_));
  NAND3_X1   g07806(.A1(new_n10241_), .A2(new_n10242_), .A3(new_n10062_), .ZN(new_n10243_));
  NAND3_X1   g07807(.A1(new_n10240_), .A2(new_n10243_), .A3(pi1196), .ZN(new_n10244_));
  NAND2_X1   g07808(.A1(new_n10244_), .A2(new_n10068_), .ZN(new_n10245_));
  NAND2_X1   g07809(.A1(new_n10245_), .A2(new_n10230_), .ZN(new_n10246_));
  OAI21_X1   g07810(.A1(new_n10246_), .A2(pi1199), .B(new_n6253_), .ZN(new_n10247_));
  NOR2_X1    g07811(.A1(new_n10246_), .A2(new_n6848_), .ZN(new_n10248_));
  AOI21_X1   g07812(.A1(new_n6851_), .A2(new_n10139_), .B(new_n10248_), .ZN(new_n10249_));
  NOR2_X1    g07813(.A1(new_n10246_), .A2(new_n6850_), .ZN(new_n10250_));
  AOI21_X1   g07814(.A1(new_n6849_), .A2(new_n10139_), .B(new_n10250_), .ZN(new_n10251_));
  OAI22_X1   g07815(.A1(new_n6853_), .A2(new_n10251_), .B1(new_n10249_), .B2(new_n6856_), .ZN(new_n10252_));
  AND2_X2    g07816(.A1(new_n10252_), .A2(pi0445), .Z(new_n10253_));
  OAI22_X1   g07817(.A1(new_n6853_), .A2(new_n10249_), .B1(new_n10251_), .B2(new_n6856_), .ZN(new_n10254_));
  AOI21_X1   g07818(.A1(new_n6859_), .A2(new_n10254_), .B(new_n10253_), .ZN(new_n10255_));
  NAND2_X1   g07819(.A1(new_n10255_), .A2(new_n9760_), .ZN(new_n10256_));
  AND2_X2    g07820(.A1(new_n10254_), .A2(pi0445), .Z(new_n10257_));
  AOI21_X1   g07821(.A1(new_n6859_), .A2(new_n10252_), .B(new_n10257_), .ZN(new_n10258_));
  NAND2_X1   g07822(.A1(new_n10258_), .A2(pi0448), .ZN(new_n10259_));
  AOI21_X1   g07823(.A1(new_n10256_), .A2(new_n10259_), .B(new_n9759_), .ZN(new_n10260_));
  NAND2_X1   g07824(.A1(new_n10255_), .A2(pi0448), .ZN(new_n10261_));
  NAND2_X1   g07825(.A1(new_n10258_), .A2(new_n9760_), .ZN(new_n10262_));
  AOI21_X1   g07826(.A1(new_n10261_), .A2(new_n10262_), .B(new_n6331_), .ZN(new_n10263_));
  NOR3_X1    g07827(.A1(new_n10260_), .A2(new_n10263_), .A3(new_n6380_), .ZN(new_n10264_));
  OAI21_X1   g07828(.A1(new_n10264_), .A2(new_n10247_), .B(new_n9778_), .ZN(new_n10265_));
  NAND3_X1   g07829(.A1(new_n10229_), .A2(new_n6350_), .A3(new_n10265_), .ZN(new_n10266_));
  NAND4_X1   g07830(.A1(new_n10090_), .A2(new_n9878_), .A3(new_n6643_), .A4(new_n10266_), .ZN(new_n10267_));
  NAND3_X1   g07831(.A1(new_n10267_), .A2(new_n9751_), .A3(new_n9877_), .ZN(new_n10268_));
  AND3_X2    g07832(.A1(new_n10268_), .A2(new_n7253_), .A3(new_n9750_), .Z(po0238));
  NAND3_X1   g07833(.A1(new_n2542_), .A2(pi0068), .A3(new_n2500_), .ZN(new_n10270_));
  NOR4_X1    g07834(.A1(new_n10270_), .A2(new_n7301_), .A3(new_n8916_), .A4(pi0064), .ZN(new_n10271_));
  AOI22_X1   g07835(.A1(new_n9177_), .A2(new_n5590_), .B1(new_n2923_), .B2(new_n10271_), .ZN(new_n10272_));
  NAND2_X1   g07836(.A1(new_n9123_), .A2(new_n6643_), .ZN(new_n10273_));
  NOR2_X1    g07837(.A1(new_n10273_), .A2(new_n10272_), .ZN(po0239));
  NOR2_X1    g07838(.A1(new_n2905_), .A2(new_n2908_), .ZN(new_n10275_));
  NOR4_X1    g07839(.A1(new_n2825_), .A2(new_n2929_), .A3(pi0073), .A4(new_n2824_), .ZN(new_n10276_));
  AOI21_X1   g07840(.A1(new_n10275_), .A2(pi0314), .B(new_n10276_), .ZN(new_n10277_));
  NOR4_X1    g07841(.A1(new_n8979_), .A2(new_n2475_), .A3(new_n8980_), .A4(new_n10277_), .ZN(po0240));
  NAND2_X1   g07842(.A1(new_n2916_), .A2(new_n2542_), .ZN(new_n10279_));
  INV_X1     g07843(.I(new_n10279_), .ZN(new_n10280_));
  NAND3_X1   g07844(.A1(new_n10280_), .A2(pi0084), .A3(new_n7417_), .ZN(new_n10281_));
  INV_X1     g07845(.I(new_n10281_), .ZN(new_n10282_));
  NOR2_X1    g07846(.A1(new_n8980_), .A2(new_n7312_), .ZN(new_n10283_));
  NAND4_X1   g07847(.A1(new_n10282_), .A2(pi0314), .A3(new_n2474_), .A4(new_n10283_), .ZN(new_n10284_));
  NAND2_X1   g07848(.A1(new_n10281_), .A2(new_n8904_), .ZN(new_n10285_));
  NAND4_X1   g07849(.A1(new_n10285_), .A2(new_n5590_), .A3(new_n2909_), .A4(new_n10283_), .ZN(new_n10286_));
  AOI21_X1   g07850(.A1(new_n10286_), .A2(new_n10284_), .B(new_n8262_), .ZN(po0241));
  NOR2_X1    g07851(.A1(new_n8641_), .A2(pi0299), .ZN(new_n10288_));
  NOR2_X1    g07852(.A1(new_n2628_), .A2(pi0219), .ZN(new_n10289_));
  AOI21_X1   g07853(.A1(new_n8510_), .A2(new_n10289_), .B(new_n10288_), .ZN(new_n10290_));
  NOR4_X1    g07854(.A1(new_n9180_), .A2(new_n2612_), .A3(po1038), .A4(new_n10290_), .ZN(po0242));
  NOR2_X1    g07855(.A1(new_n5569_), .A2(new_n2543_), .ZN(new_n10292_));
  NAND3_X1   g07856(.A1(new_n10292_), .A2(new_n5590_), .A3(new_n8983_), .ZN(new_n10293_));
  NAND4_X1   g07857(.A1(new_n8981_), .A2(pi0067), .A3(new_n2902_), .A4(new_n2907_), .ZN(new_n10294_));
  AOI21_X1   g07858(.A1(new_n10293_), .A2(new_n10294_), .B(new_n8979_), .ZN(po0243));
  NOR2_X1    g07859(.A1(new_n6751_), .A2(new_n6809_), .ZN(new_n10296_));
  AOI22_X1   g07860(.A1(new_n6805_), .A2(new_n9192_), .B1(new_n10296_), .B2(new_n9190_), .ZN(new_n10297_));
  NOR2_X1    g07861(.A1(new_n10297_), .A2(new_n8898_), .ZN(po0244));
  INV_X1     g07862(.I(new_n8980_), .ZN(new_n10299_));
  NAND3_X1   g07863(.A1(new_n2906_), .A2(new_n2728_), .A3(new_n10299_), .ZN(new_n10300_));
  NOR4_X1    g07864(.A1(new_n8262_), .A2(new_n5590_), .A3(new_n2737_), .A4(new_n10300_), .ZN(po0245));
  INV_X1     g07865(.I(new_n8218_), .ZN(new_n10302_));
  INV_X1     g07866(.I(new_n9886_), .ZN(new_n10303_));
  NAND3_X1   g07867(.A1(new_n8923_), .A2(new_n6669_), .A3(new_n9887_), .ZN(new_n10304_));
  NOR3_X1    g07868(.A1(new_n10304_), .A2(new_n8939_), .A3(new_n10303_), .ZN(new_n10305_));
  NOR2_X1    g07869(.A1(new_n10305_), .A2(new_n3041_), .ZN(new_n10306_));
  NOR2_X1    g07870(.A1(new_n10306_), .A2(new_n2612_), .ZN(new_n10307_));
  OAI21_X1   g07871(.A1(new_n8926_), .A2(new_n6259_), .B(new_n3041_), .ZN(new_n10308_));
  NAND4_X1   g07872(.A1(new_n10307_), .A2(new_n10308_), .A3(new_n6349_), .A4(new_n10302_), .ZN(new_n10309_));
  NAND4_X1   g07873(.A1(new_n2748_), .A2(new_n3041_), .A3(new_n9275_), .A4(new_n6258_), .ZN(new_n10310_));
  NOR3_X1    g07874(.A1(new_n2612_), .A2(new_n9234_), .A3(new_n10310_), .ZN(new_n10311_));
  NAND4_X1   g07875(.A1(new_n10311_), .A2(pi0088), .A3(new_n6350_), .A4(new_n8251_), .ZN(new_n10312_));
  AOI21_X1   g07876(.A1(new_n10309_), .A2(new_n10312_), .B(po1038), .ZN(po0246));
  NOR4_X1    g07877(.A1(new_n8275_), .A2(new_n7413_), .A3(new_n8242_), .A4(new_n7312_), .ZN(new_n10314_));
  NAND3_X1   g07878(.A1(new_n10314_), .A2(pi0841), .A3(new_n6676_), .ZN(new_n10315_));
  NAND2_X1   g07879(.A1(new_n10315_), .A2(new_n2835_), .ZN(new_n10316_));
  NAND3_X1   g07880(.A1(new_n10316_), .A2(new_n2529_), .A3(new_n8259_), .ZN(new_n10317_));
  AOI21_X1   g07881(.A1(pi0070), .A2(new_n7333_), .B(new_n10317_), .ZN(po0247));
  OAI21_X1   g07882(.A1(new_n7464_), .A2(pi1050), .B(new_n2985_), .ZN(new_n10319_));
  OAI21_X1   g07883(.A1(new_n2739_), .A2(new_n3179_), .B(pi0090), .ZN(new_n10320_));
  AND3_X2    g07884(.A1(new_n10320_), .A2(new_n10319_), .A3(new_n9143_), .Z(po0248));
  NAND3_X1   g07885(.A1(new_n3188_), .A2(pi0024), .A3(new_n2763_), .ZN(new_n10322_));
  NAND2_X1   g07886(.A1(new_n2839_), .A2(new_n8970_), .ZN(new_n10323_));
  OAI21_X1   g07887(.A1(new_n10323_), .A2(new_n10322_), .B(new_n2627_), .ZN(new_n10324_));
  INV_X1     g07888(.I(new_n8250_), .ZN(new_n10325_));
  INV_X1     g07889(.I(new_n8251_), .ZN(new_n10326_));
  OAI22_X1   g07890(.A1(new_n6718_), .A2(pi0058), .B1(new_n10325_), .B2(new_n10326_), .ZN(new_n10327_));
  NOR2_X1    g07891(.A1(new_n3188_), .A2(new_n8254_), .ZN(new_n10328_));
  AOI21_X1   g07892(.A1(new_n10327_), .A2(new_n10328_), .B(new_n10324_), .ZN(new_n10329_));
  NOR3_X1    g07893(.A1(new_n6813_), .A2(new_n8265_), .A3(new_n10329_), .ZN(po0249));
  INV_X1     g07894(.I(new_n9081_), .ZN(new_n10331_));
  NOR2_X1    g07895(.A1(new_n5756_), .A2(new_n2614_), .ZN(new_n10332_));
  NOR2_X1    g07896(.A1(new_n7525_), .A2(pi0299), .ZN(new_n10333_));
  AOI22_X1   g07897(.A1(new_n6805_), .A2(new_n10333_), .B1(new_n10296_), .B2(new_n10332_), .ZN(new_n10334_));
  OR3_X2     g07898(.A1(new_n10334_), .A2(new_n2567_), .A3(new_n10331_), .Z(new_n10335_));
  NOR2_X1    g07899(.A1(new_n2530_), .A2(new_n3444_), .ZN(new_n10336_));
  NAND4_X1   g07900(.A1(new_n10336_), .A2(new_n5590_), .A3(pi1050), .A4(new_n3415_), .ZN(new_n10337_));
  AOI21_X1   g07901(.A1(new_n10335_), .A2(new_n10337_), .B(new_n8256_), .ZN(po0250));
  INV_X1     g07902(.I(pi1050), .ZN(new_n10339_));
  AOI21_X1   g07903(.A1(new_n2531_), .A2(new_n10339_), .B(new_n3444_), .ZN(new_n10340_));
  NOR4_X1    g07904(.A1(new_n2548_), .A2(new_n2771_), .A3(new_n3179_), .A4(new_n9142_), .ZN(new_n10341_));
  OAI21_X1   g07905(.A1(new_n10341_), .A2(pi0092), .B(new_n8257_), .ZN(new_n10342_));
  NOR2_X1    g07906(.A1(new_n10342_), .A2(new_n10340_), .ZN(po0251));
  NOR2_X1    g07907(.A1(new_n8960_), .A2(new_n9116_), .ZN(new_n10344_));
  NAND2_X1   g07908(.A1(new_n7324_), .A2(pi0252), .ZN(new_n10345_));
  NAND2_X1   g07909(.A1(new_n10344_), .A2(new_n10345_), .ZN(new_n10346_));
  AOI21_X1   g07910(.A1(new_n10344_), .A2(new_n3025_), .B(new_n3041_), .ZN(new_n10347_));
  NOR2_X1    g07911(.A1(new_n8958_), .A2(new_n8328_), .ZN(new_n10348_));
  NOR2_X1    g07912(.A1(new_n2875_), .A2(new_n10348_), .ZN(new_n10349_));
  NAND3_X1   g07913(.A1(new_n8253_), .A2(new_n2786_), .A3(pi0252), .ZN(new_n10350_));
  OAI22_X1   g07914(.A1(new_n10349_), .A2(new_n10350_), .B1(new_n3084_), .B2(new_n10347_), .ZN(new_n10351_));
  OAI21_X1   g07915(.A1(new_n8960_), .A2(new_n9116_), .B(po0840), .ZN(new_n10352_));
  NAND3_X1   g07916(.A1(new_n10351_), .A2(new_n7324_), .A3(new_n10352_), .ZN(new_n10353_));
  AOI21_X1   g07917(.A1(new_n10353_), .A2(new_n10346_), .B(new_n8260_), .ZN(po0252));
  INV_X1     g07918(.I(new_n10314_), .ZN(new_n10355_));
  NAND2_X1   g07919(.A1(new_n8253_), .A2(new_n2630_), .ZN(new_n10356_));
  NOR3_X1    g07920(.A1(new_n10355_), .A2(new_n9114_), .A3(new_n10356_), .ZN(new_n10357_));
  NAND3_X1   g07921(.A1(new_n2524_), .A2(new_n2725_), .A3(pi0095), .ZN(new_n10358_));
  OAI21_X1   g07922(.A1(new_n9235_), .A2(new_n10358_), .B(new_n2627_), .ZN(new_n10359_));
  OAI21_X1   g07923(.A1(new_n10359_), .A2(new_n10357_), .B(new_n8280_), .ZN(new_n10360_));
  INV_X1     g07924(.I(new_n9207_), .ZN(new_n10361_));
  NOR3_X1    g07925(.A1(new_n10361_), .A2(new_n5551_), .A3(new_n9206_), .ZN(new_n10362_));
  NAND2_X1   g07926(.A1(new_n5536_), .A2(new_n5452_), .ZN(new_n10363_));
  NOR3_X1    g07927(.A1(new_n10363_), .A2(new_n3338_), .A3(new_n9209_), .ZN(new_n10364_));
  NOR3_X1    g07928(.A1(new_n10362_), .A2(new_n2627_), .A3(new_n10364_), .ZN(new_n10365_));
  NOR2_X1    g07929(.A1(new_n10360_), .A2(new_n10365_), .ZN(po0253));
  NAND4_X1   g07930(.A1(new_n2533_), .A2(new_n2743_), .A3(new_n2835_), .A4(pi0096), .ZN(new_n10367_));
  NOR2_X1    g07931(.A1(po0840), .A2(new_n2998_), .ZN(new_n10368_));
  NOR4_X1    g07932(.A1(new_n3009_), .A2(new_n3010_), .A3(new_n10367_), .A4(new_n10368_), .ZN(new_n10369_));
  INV_X1     g07933(.I(new_n10368_), .ZN(new_n10370_));
  NOR4_X1    g07934(.A1(new_n2811_), .A2(pi0032), .A3(new_n2726_), .A4(new_n10370_), .ZN(new_n10371_));
  OAI21_X1   g07935(.A1(new_n10371_), .A2(new_n10369_), .B(new_n2462_), .ZN(new_n10372_));
  NOR2_X1    g07936(.A1(new_n2751_), .A2(pi0024), .ZN(new_n10373_));
  NAND4_X1   g07937(.A1(new_n10373_), .A2(new_n2725_), .A3(pi0095), .A4(new_n2524_), .ZN(new_n10374_));
  AOI21_X1   g07938(.A1(new_n10372_), .A2(new_n10374_), .B(new_n8260_), .ZN(po0254));
  INV_X1     g07939(.I(new_n9210_), .ZN(new_n10376_));
  NAND4_X1   g07940(.A1(new_n10376_), .A2(pi0039), .A3(new_n5536_), .A4(pi0593), .ZN(new_n10377_));
  NOR2_X1    g07941(.A1(new_n6723_), .A2(new_n2766_), .ZN(new_n10378_));
  OAI21_X1   g07942(.A1(new_n10370_), .A2(new_n5350_), .B(new_n8241_), .ZN(new_n10379_));
  NAND4_X1   g07943(.A1(new_n10378_), .A2(new_n2742_), .A3(new_n9202_), .A4(new_n10379_), .ZN(new_n10380_));
  AOI21_X1   g07944(.A1(new_n10377_), .A2(new_n10380_), .B(new_n8281_), .ZN(po0255));
  AOI21_X1   g07945(.A1(new_n9245_), .A2(new_n3444_), .B(new_n10336_), .ZN(new_n10382_));
  NOR4_X1    g07946(.A1(new_n10382_), .A2(new_n5590_), .A3(new_n10339_), .A4(new_n8258_), .ZN(po0256));
  NOR4_X1    g07947(.A1(new_n8349_), .A2(pi0072), .A3(new_n3369_), .A4(new_n3360_), .ZN(new_n10384_));
  AOI22_X1   g07948(.A1(new_n10384_), .A2(new_n7506_), .B1(new_n2627_), .B2(new_n8600_), .ZN(new_n10385_));
  INV_X1     g07949(.I(new_n8356_), .ZN(new_n10386_));
  INV_X1     g07950(.I(new_n10384_), .ZN(new_n10387_));
  NAND3_X1   g07951(.A1(new_n2821_), .A2(new_n2628_), .A3(pi0174), .ZN(new_n10388_));
  OAI22_X1   g07952(.A1(new_n10387_), .A2(new_n2628_), .B1(new_n10386_), .B2(new_n10388_), .ZN(new_n10389_));
  AOI21_X1   g07953(.A1(new_n10389_), .A2(pi0232), .B(new_n2627_), .ZN(new_n10390_));
  AOI21_X1   g07954(.A1(new_n2627_), .A2(new_n8601_), .B(new_n10390_), .ZN(new_n10391_));
  OAI21_X1   g07955(.A1(new_n10391_), .A2(new_n6645_), .B(new_n6643_), .ZN(new_n10392_));
  NOR2_X1    g07956(.A1(new_n8369_), .A2(new_n8601_), .ZN(new_n10393_));
  INV_X1     g07957(.I(new_n10393_), .ZN(new_n10394_));
  NOR2_X1    g07958(.A1(new_n8860_), .A2(new_n5313_), .ZN(new_n10395_));
  INV_X1     g07959(.I(new_n8383_), .ZN(new_n10396_));
  AOI21_X1   g07960(.A1(new_n10396_), .A2(new_n8375_), .B(new_n8601_), .ZN(new_n10397_));
  OAI21_X1   g07961(.A1(new_n10397_), .A2(new_n10395_), .B(new_n8491_), .ZN(new_n10398_));
  OAI21_X1   g07962(.A1(new_n10398_), .A2(new_n8370_), .B(new_n10394_), .ZN(new_n10399_));
  OAI21_X1   g07963(.A1(new_n10399_), .A2(pi0039), .B(new_n2626_), .ZN(new_n10400_));
  AOI21_X1   g07964(.A1(new_n10391_), .A2(new_n5792_), .B(new_n3465_), .ZN(new_n10401_));
  OAI21_X1   g07965(.A1(new_n10400_), .A2(new_n10390_), .B(new_n10401_), .ZN(new_n10402_));
  AOI22_X1   g07966(.A1(new_n8493_), .A2(new_n8600_), .B1(new_n5310_), .B2(new_n8389_), .ZN(new_n10403_));
  NOR2_X1    g07967(.A1(new_n10403_), .A2(new_n8372_), .ZN(new_n10404_));
  AOI21_X1   g07968(.A1(new_n10404_), .A2(new_n8369_), .B(new_n10393_), .ZN(new_n10405_));
  AOI21_X1   g07969(.A1(new_n10405_), .A2(new_n2627_), .B(new_n10390_), .ZN(new_n10406_));
  INV_X1     g07970(.I(new_n10391_), .ZN(new_n10407_));
  AOI21_X1   g07971(.A1(new_n10407_), .A2(pi0038), .B(pi0087), .ZN(new_n10408_));
  OAI21_X1   g07972(.A1(new_n10406_), .A2(new_n8667_), .B(new_n10408_), .ZN(new_n10409_));
  OAI21_X1   g07973(.A1(new_n8346_), .A2(new_n2821_), .B(pi0099), .ZN(new_n10410_));
  NOR2_X1    g07974(.A1(new_n8445_), .A2(new_n10410_), .ZN(new_n10411_));
  NOR2_X1    g07975(.A1(new_n10411_), .A2(pi0228), .ZN(new_n10412_));
  OAI21_X1   g07976(.A1(new_n8483_), .A2(new_n10410_), .B(new_n8745_), .ZN(new_n10413_));
  OAI21_X1   g07977(.A1(new_n8476_), .A2(new_n10410_), .B(new_n8744_), .ZN(new_n10414_));
  NAND2_X1   g07978(.A1(new_n10413_), .A2(new_n10414_), .ZN(new_n10415_));
  AOI22_X1   g07979(.A1(new_n10415_), .A2(pi0228), .B1(new_n8590_), .B2(new_n10412_), .ZN(new_n10416_));
  INV_X1     g07980(.I(new_n10389_), .ZN(new_n10417_));
  OAI21_X1   g07981(.A1(new_n8379_), .A2(new_n8282_), .B(new_n7506_), .ZN(new_n10418_));
  OAI21_X1   g07982(.A1(new_n10418_), .A2(new_n10417_), .B(new_n3270_), .ZN(new_n10419_));
  AOI21_X1   g07983(.A1(new_n10416_), .A2(new_n2627_), .B(new_n10419_), .ZN(new_n10420_));
  AOI21_X1   g07984(.A1(new_n10407_), .A2(new_n2575_), .B(new_n3458_), .ZN(new_n10421_));
  NAND2_X1   g07985(.A1(new_n8553_), .A2(pi0228), .ZN(new_n10422_));
  NAND2_X1   g07986(.A1(new_n8400_), .A2(pi0228), .ZN(new_n10423_));
  NAND2_X1   g07987(.A1(new_n10423_), .A2(new_n8600_), .ZN(new_n10424_));
  NAND3_X1   g07988(.A1(new_n10424_), .A2(new_n2574_), .A3(new_n10422_), .ZN(new_n10425_));
  AOI21_X1   g07989(.A1(new_n10425_), .A2(new_n10421_), .B(pi0075), .ZN(new_n10426_));
  OAI21_X1   g07990(.A1(new_n10420_), .A2(new_n10409_), .B(new_n10426_), .ZN(new_n10427_));
  AOI21_X1   g07991(.A1(new_n10427_), .A2(new_n10402_), .B(new_n6648_), .ZN(new_n10428_));
  OAI22_X1   g07992(.A1(new_n10428_), .A2(new_n10392_), .B1(new_n6643_), .B2(new_n10385_), .ZN(po0257));
  NOR4_X1    g07993(.A1(new_n7325_), .A2(pi0024), .A3(new_n7288_), .A4(new_n7337_), .ZN(new_n10430_));
  NAND2_X1   g07994(.A1(new_n8222_), .A2(new_n6698_), .ZN(new_n10431_));
  AOI21_X1   g07995(.A1(new_n10431_), .A2(pi0129), .B(new_n6696_), .ZN(new_n10432_));
  NOR2_X1    g07996(.A1(new_n8222_), .A2(new_n7322_), .ZN(new_n10433_));
  OAI22_X1   g07997(.A1(new_n10433_), .A2(new_n8225_), .B1(new_n5335_), .B2(new_n5309_), .ZN(new_n10434_));
  NOR2_X1    g07998(.A1(new_n10434_), .A2(new_n10432_), .ZN(new_n10435_));
  NOR4_X1    g07999(.A1(new_n10435_), .A2(pi0075), .A3(new_n7599_), .A4(new_n8667_), .ZN(new_n10436_));
  OAI21_X1   g08000(.A1(new_n10436_), .A2(new_n10430_), .B(new_n7267_), .ZN(new_n10437_));
  NOR2_X1    g08001(.A1(new_n10437_), .A2(new_n2530_), .ZN(po0258));
  INV_X1     g08002(.I(new_n8374_), .ZN(new_n10439_));
  NOR4_X1    g08003(.A1(new_n5437_), .A2(new_n3369_), .A3(pi0161), .A4(pi0166), .ZN(new_n10440_));
  NAND2_X1   g08004(.A1(new_n10440_), .A2(new_n2821_), .ZN(new_n10441_));
  OAI22_X1   g08005(.A1(new_n10441_), .A2(new_n7507_), .B1(pi0039), .B2(new_n10439_), .ZN(new_n10442_));
  NAND2_X1   g08006(.A1(new_n10442_), .A2(po1038), .ZN(new_n10443_));
  NAND4_X1   g08007(.A1(new_n8354_), .A2(new_n2821_), .A3(new_n8058_), .A4(pi0174), .ZN(new_n10444_));
  AOI21_X1   g08008(.A1(new_n10444_), .A2(new_n2628_), .B(new_n5666_), .ZN(new_n10445_));
  NAND2_X1   g08009(.A1(new_n10441_), .A2(pi0299), .ZN(new_n10446_));
  AOI21_X1   g08010(.A1(new_n10445_), .A2(new_n10446_), .B(new_n2627_), .ZN(new_n10447_));
  AOI21_X1   g08011(.A1(new_n2627_), .A2(new_n10439_), .B(new_n10447_), .ZN(new_n10448_));
  OAI21_X1   g08012(.A1(new_n10448_), .A2(new_n6645_), .B(new_n6643_), .ZN(new_n10449_));
  NOR2_X1    g08013(.A1(new_n8369_), .A2(new_n10439_), .ZN(new_n10450_));
  INV_X1     g08014(.I(new_n10450_), .ZN(new_n10451_));
  NOR2_X1    g08015(.A1(new_n10396_), .A2(new_n10439_), .ZN(new_n10452_));
  OAI21_X1   g08016(.A1(new_n10452_), .A2(new_n8391_), .B(new_n5322_), .ZN(new_n10453_));
  OAI21_X1   g08017(.A1(new_n10453_), .A2(new_n8370_), .B(new_n10451_), .ZN(new_n10454_));
  OAI21_X1   g08018(.A1(new_n10454_), .A2(pi0039), .B(new_n2626_), .ZN(new_n10455_));
  AOI21_X1   g08019(.A1(new_n10448_), .A2(new_n5792_), .B(new_n3465_), .ZN(new_n10456_));
  OAI21_X1   g08020(.A1(new_n10455_), .A2(new_n10447_), .B(new_n10456_), .ZN(new_n10457_));
  INV_X1     g08021(.I(new_n10447_), .ZN(new_n10458_));
  NAND4_X1   g08022(.A1(new_n8378_), .A2(new_n8377_), .A3(pi0228), .A4(new_n3270_), .ZN(new_n10459_));
  AOI22_X1   g08023(.A1(new_n10459_), .A2(new_n8374_), .B1(new_n8373_), .B2(new_n8887_), .ZN(new_n10460_));
  AOI21_X1   g08024(.A1(new_n10460_), .A2(new_n2627_), .B(new_n3458_), .ZN(new_n10461_));
  AOI21_X1   g08025(.A1(new_n10461_), .A2(new_n10458_), .B(pi0075), .ZN(new_n10462_));
  NOR4_X1    g08026(.A1(new_n8869_), .A2(pi0144), .A3(new_n7488_), .A4(new_n8355_), .ZN(new_n10463_));
  OAI21_X1   g08027(.A1(new_n10463_), .A2(pi0299), .B(new_n7506_), .ZN(new_n10464_));
  AOI21_X1   g08028(.A1(new_n8868_), .A2(new_n10440_), .B(new_n2628_), .ZN(new_n10465_));
  OAI21_X1   g08029(.A1(new_n10464_), .A2(new_n10465_), .B(new_n3270_), .ZN(new_n10466_));
  NAND2_X1   g08030(.A1(new_n8444_), .A2(pi0101), .ZN(new_n10467_));
  NAND3_X1   g08031(.A1(new_n8439_), .A2(new_n2458_), .A3(new_n10467_), .ZN(new_n10468_));
  NAND2_X1   g08032(.A1(new_n8482_), .A2(pi0101), .ZN(new_n10469_));
  NAND3_X1   g08033(.A1(new_n8626_), .A2(new_n3026_), .A3(new_n10469_), .ZN(new_n10470_));
  NAND2_X1   g08034(.A1(new_n8475_), .A2(pi0101), .ZN(new_n10471_));
  NAND3_X1   g08035(.A1(new_n10471_), .A2(new_n3025_), .A3(new_n8464_), .ZN(new_n10472_));
  NAND2_X1   g08036(.A1(new_n10470_), .A2(new_n10472_), .ZN(new_n10473_));
  AOI21_X1   g08037(.A1(new_n10473_), .A2(pi0228), .B(pi0039), .ZN(new_n10474_));
  AOI21_X1   g08038(.A1(new_n10474_), .A2(new_n10468_), .B(new_n10466_), .ZN(new_n10475_));
  OAI21_X1   g08039(.A1(new_n8381_), .A2(pi0044), .B(new_n8374_), .ZN(new_n10476_));
  AOI21_X1   g08040(.A1(new_n10476_), .A2(new_n8390_), .B(new_n5321_), .ZN(new_n10477_));
  AOI21_X1   g08041(.A1(new_n10477_), .A2(new_n8369_), .B(new_n10450_), .ZN(new_n10478_));
  AOI21_X1   g08042(.A1(new_n10478_), .A2(new_n2627_), .B(new_n10447_), .ZN(new_n10479_));
  NOR2_X1    g08043(.A1(new_n10448_), .A2(new_n3265_), .ZN(new_n10480_));
  NOR2_X1    g08044(.A1(new_n10480_), .A2(pi0087), .ZN(new_n10481_));
  OAI21_X1   g08045(.A1(new_n10479_), .A2(new_n8667_), .B(new_n10481_), .ZN(new_n10482_));
  OAI21_X1   g08046(.A1(new_n10475_), .A2(new_n10482_), .B(new_n10462_), .ZN(new_n10483_));
  AOI21_X1   g08047(.A1(new_n10483_), .A2(new_n10457_), .B(new_n6648_), .ZN(new_n10484_));
  OAI21_X1   g08048(.A1(new_n10484_), .A2(new_n10449_), .B(new_n10443_), .ZN(po0259));
  NAND3_X1   g08049(.A1(new_n2963_), .A2(new_n2496_), .A3(new_n7297_), .ZN(new_n10486_));
  NOR2_X1    g08050(.A1(new_n10273_), .A2(new_n10486_), .ZN(po0260));
  NAND2_X1   g08051(.A1(new_n10300_), .A2(new_n2508_), .ZN(new_n10488_));
  AOI21_X1   g08052(.A1(new_n10488_), .A2(new_n5562_), .B(pi0314), .ZN(new_n10489_));
  NOR2_X1    g08053(.A1(new_n2731_), .A2(new_n2508_), .ZN(new_n10490_));
  AOI21_X1   g08054(.A1(new_n10490_), .A2(new_n2847_), .B(new_n5590_), .ZN(new_n10491_));
  NOR4_X1    g08055(.A1(new_n10489_), .A2(new_n2733_), .A3(new_n8262_), .A4(new_n10491_), .ZN(po0261));
  OAI21_X1   g08056(.A1(new_n7324_), .A2(new_n6350_), .B(new_n8219_), .ZN(new_n10493_));
  NAND2_X1   g08057(.A1(new_n8434_), .A2(new_n10493_), .ZN(new_n10494_));
  NOR2_X1    g08058(.A1(new_n10305_), .A2(new_n5323_), .ZN(new_n10495_));
  AOI21_X1   g08059(.A1(new_n10495_), .A2(new_n8224_), .B(new_n8218_), .ZN(new_n10496_));
  NAND2_X1   g08060(.A1(new_n10304_), .A2(new_n2509_), .ZN(new_n10497_));
  NOR2_X1    g08061(.A1(new_n8939_), .A2(pi0047), .ZN(new_n10498_));
  NAND4_X1   g08062(.A1(new_n5365_), .A2(new_n2732_), .A3(new_n10497_), .A4(new_n10498_), .ZN(new_n10499_));
  NAND4_X1   g08063(.A1(new_n10305_), .A2(po1057), .A3(new_n8224_), .A4(new_n10302_), .ZN(new_n10500_));
  NAND2_X1   g08064(.A1(new_n10499_), .A2(new_n10500_), .ZN(new_n10501_));
  NAND3_X1   g08065(.A1(new_n10501_), .A2(new_n6350_), .A3(new_n10496_), .ZN(new_n10502_));
  AOI21_X1   g08066(.A1(new_n10502_), .A2(new_n10494_), .B(new_n8260_), .ZN(po0262));
  NOR2_X1    g08067(.A1(new_n9113_), .A2(new_n7278_), .ZN(new_n10504_));
  OAI21_X1   g08068(.A1(pi0053), .A2(new_n9111_), .B(new_n2795_), .ZN(new_n10505_));
  NOR3_X1    g08069(.A1(new_n10505_), .A2(pi0024), .A3(new_n2787_), .ZN(new_n10506_));
  OAI21_X1   g08070(.A1(new_n10506_), .A2(new_n10504_), .B(pi0841), .ZN(new_n10507_));
  NAND3_X1   g08071(.A1(new_n9102_), .A2(new_n7278_), .A3(new_n3179_), .ZN(new_n10508_));
  AOI21_X1   g08072(.A1(new_n10507_), .A2(new_n10508_), .B(new_n8262_), .ZN(po0264));
  INV_X1     g08073(.I(new_n9161_), .ZN(new_n10510_));
  NOR3_X1    g08074(.A1(new_n8262_), .A2(pi0999), .A3(new_n10510_), .ZN(po0265));
  AOI21_X1   g08075(.A1(new_n6674_), .A2(new_n2864_), .B(pi0108), .ZN(new_n10512_));
  OR3_X2     g08076(.A1(new_n10512_), .A2(new_n8327_), .A3(new_n7273_), .Z(new_n10513_));
  NOR2_X1    g08077(.A1(new_n10513_), .A2(new_n6679_), .ZN(new_n10514_));
  AOI21_X1   g08078(.A1(new_n10514_), .A2(new_n8312_), .B(pi0051), .ZN(new_n10515_));
  NOR2_X1    g08079(.A1(new_n8312_), .A2(new_n6679_), .ZN(new_n10516_));
  NOR2_X1    g08080(.A1(new_n6675_), .A2(new_n5590_), .ZN(new_n10517_));
  NOR2_X1    g08081(.A1(new_n10513_), .A2(pi0314), .ZN(new_n10518_));
  OAI21_X1   g08082(.A1(new_n10518_), .A2(new_n10517_), .B(new_n10516_), .ZN(new_n10519_));
  AOI21_X1   g08083(.A1(new_n10515_), .A2(new_n10519_), .B(new_n3273_), .ZN(new_n10520_));
  AOI21_X1   g08084(.A1(new_n10520_), .A2(new_n6715_), .B(pi0087), .ZN(new_n10521_));
  NOR3_X1    g08085(.A1(new_n10521_), .A2(new_n5304_), .A3(new_n7268_), .ZN(po0266));
  NOR4_X1    g08086(.A1(new_n8262_), .A2(new_n5590_), .A3(new_n9379_), .A4(new_n9227_), .ZN(po0267));
  NOR2_X1    g08087(.A1(new_n8217_), .A2(new_n8220_), .ZN(new_n10524_));
  NOR4_X1    g08088(.A1(new_n10303_), .A2(pi0082), .A3(pi0109), .A4(new_n2912_), .ZN(new_n10525_));
  NOR3_X1    g08089(.A1(new_n8984_), .A2(pi0068), .A3(new_n2917_), .ZN(new_n10526_));
  NAND3_X1   g08090(.A1(new_n10526_), .A2(new_n2728_), .A3(new_n10525_), .ZN(new_n10527_));
  INV_X1     g08091(.I(new_n10527_), .ZN(new_n10528_));
  AOI22_X1   g08092(.A1(new_n10528_), .A2(pi0314), .B1(new_n8413_), .B2(new_n10524_), .ZN(new_n10529_));
  NOR2_X1    g08093(.A1(new_n10529_), .A2(new_n8262_), .ZN(po0268));
  NOR2_X1    g08094(.A1(new_n10527_), .A2(pi0314), .ZN(new_n10531_));
  AOI22_X1   g08095(.A1(new_n10373_), .A2(pi0072), .B1(new_n10531_), .B2(new_n7682_), .ZN(new_n10532_));
  NOR3_X1    g08096(.A1(new_n10532_), .A2(new_n2536_), .A3(new_n8260_), .ZN(po0269));
  INV_X1     g08097(.I(pi0468), .ZN(new_n10534_));
  NAND2_X1   g08098(.A1(new_n10534_), .A2(pi0124), .ZN(po0270));
  NAND2_X1   g08099(.A1(new_n8598_), .A2(new_n2627_), .ZN(new_n10536_));
  AOI21_X1   g08100(.A1(new_n8549_), .A2(new_n5320_), .B(new_n8370_), .ZN(new_n10537_));
  NAND2_X1   g08101(.A1(new_n8369_), .A2(new_n5320_), .ZN(new_n10538_));
  NOR4_X1    g08102(.A1(new_n8390_), .A2(pi0113), .A3(new_n5311_), .A4(new_n10538_), .ZN(new_n10539_));
  INV_X1     g08103(.I(new_n10539_), .ZN(new_n10540_));
  OAI22_X1   g08104(.A1(new_n10537_), .A2(new_n8621_), .B1(new_n6707_), .B2(new_n10540_), .ZN(new_n10541_));
  OAI21_X1   g08105(.A1(new_n2626_), .A2(new_n10536_), .B(pi0075), .ZN(new_n10542_));
  AOI21_X1   g08106(.A1(new_n10541_), .A2(new_n2658_), .B(new_n10542_), .ZN(new_n10543_));
  OAI22_X1   g08107(.A1(new_n8647_), .A2(new_n8621_), .B1(pi0113), .B2(new_n10422_), .ZN(new_n10544_));
  OAI21_X1   g08108(.A1(new_n10536_), .A2(new_n3270_), .B(pi0087), .ZN(new_n10545_));
  AOI21_X1   g08109(.A1(new_n10544_), .A2(new_n2574_), .B(new_n10545_), .ZN(new_n10546_));
  OR2_X2     g08110(.A1(new_n8602_), .A2(new_n8597_), .Z(new_n10547_));
  NAND2_X1   g08111(.A1(new_n8590_), .A2(new_n8597_), .ZN(new_n10548_));
  AOI21_X1   g08112(.A1(new_n10548_), .A2(new_n10547_), .B(pi0228), .ZN(new_n10549_));
  AND2_X2    g08113(.A1(new_n8476_), .A2(new_n3025_), .Z(new_n10550_));
  NOR2_X1    g08114(.A1(new_n8484_), .A2(new_n3025_), .ZN(new_n10551_));
  OAI21_X1   g08115(.A1(new_n10551_), .A2(new_n10550_), .B(new_n8599_), .ZN(new_n10552_));
  AOI21_X1   g08116(.A1(new_n5311_), .A2(pi0072), .B(new_n8597_), .ZN(new_n10553_));
  OAI21_X1   g08117(.A1(new_n8747_), .A2(pi0113), .B(pi0228), .ZN(new_n10554_));
  AOI21_X1   g08118(.A1(new_n10552_), .A2(new_n10553_), .B(new_n10554_), .ZN(new_n10555_));
  NOR3_X1    g08119(.A1(new_n10555_), .A2(pi0039), .A3(new_n10549_), .ZN(new_n10556_));
  NAND2_X1   g08120(.A1(new_n8574_), .A2(new_n6703_), .ZN(new_n10557_));
  NAND2_X1   g08121(.A1(new_n10557_), .A2(new_n5320_), .ZN(new_n10558_));
  AOI21_X1   g08122(.A1(new_n10558_), .A2(new_n8369_), .B(new_n8621_), .ZN(new_n10559_));
  OAI21_X1   g08123(.A1(new_n10559_), .A2(new_n10539_), .B(new_n2627_), .ZN(new_n10560_));
  AOI22_X1   g08124(.A1(new_n10560_), .A2(new_n8489_), .B1(pi0038), .B2(new_n10536_), .ZN(new_n10561_));
  OAI21_X1   g08125(.A1(new_n10556_), .A2(new_n3271_), .B(new_n10561_), .ZN(new_n10562_));
  AOI21_X1   g08126(.A1(new_n10562_), .A2(new_n3458_), .B(new_n10546_), .ZN(new_n10563_));
  OAI21_X1   g08127(.A1(new_n10563_), .A2(pi0075), .B(new_n7267_), .ZN(new_n10564_));
  OAI22_X1   g08128(.A1(new_n10564_), .A2(new_n10543_), .B1(new_n7267_), .B2(new_n10536_), .ZN(po0271));
  NOR2_X1    g08129(.A1(new_n8545_), .A2(pi0072), .ZN(new_n10566_));
  NAND2_X1   g08130(.A1(new_n10566_), .A2(new_n2627_), .ZN(new_n10567_));
  NAND2_X1   g08131(.A1(new_n8726_), .A2(pi0114), .ZN(new_n10568_));
  NAND3_X1   g08132(.A1(new_n10568_), .A2(new_n8560_), .A3(new_n9001_), .ZN(new_n10569_));
  INV_X1     g08133(.I(new_n10566_), .ZN(new_n10570_));
  AOI21_X1   g08134(.A1(new_n9002_), .A2(new_n10570_), .B(new_n2659_), .ZN(new_n10571_));
  OAI21_X1   g08135(.A1(new_n2626_), .A2(new_n10567_), .B(pi0075), .ZN(new_n10572_));
  AOI21_X1   g08136(.A1(new_n10569_), .A2(new_n10571_), .B(new_n10572_), .ZN(new_n10573_));
  AOI21_X1   g08137(.A1(new_n3271_), .A2(new_n10567_), .B(new_n9083_), .ZN(new_n10574_));
  NOR3_X1    g08138(.A1(new_n8577_), .A2(pi0115), .A3(new_n2458_), .ZN(new_n10575_));
  OAI21_X1   g08139(.A1(new_n10575_), .A2(new_n10570_), .B(new_n3270_), .ZN(new_n10576_));
  OAI21_X1   g08140(.A1(new_n10576_), .A2(new_n8651_), .B(new_n10574_), .ZN(new_n10577_));
  NAND2_X1   g08141(.A1(new_n10577_), .A2(new_n3465_), .ZN(new_n10578_));
  AOI21_X1   g08142(.A1(new_n10567_), .A2(pi0038), .B(pi0087), .ZN(new_n10579_));
  AOI21_X1   g08143(.A1(new_n8579_), .A2(pi0114), .B(new_n9002_), .ZN(new_n10580_));
  OAI21_X1   g08144(.A1(new_n9001_), .A2(new_n10566_), .B(new_n2627_), .ZN(new_n10581_));
  AOI21_X1   g08145(.A1(new_n10580_), .A2(new_n8558_), .B(new_n10581_), .ZN(new_n10582_));
  OAI21_X1   g08146(.A1(new_n10582_), .A2(new_n8667_), .B(new_n10579_), .ZN(new_n10583_));
  NOR2_X1    g08147(.A1(new_n10570_), .A2(new_n8587_), .ZN(new_n10584_));
  NAND2_X1   g08148(.A1(new_n8758_), .A2(pi0114), .ZN(new_n10585_));
  OR2_X2     g08149(.A1(new_n8749_), .A2(pi0114), .Z(new_n10586_));
  AOI21_X1   g08150(.A1(new_n10585_), .A2(new_n10586_), .B(pi0115), .ZN(new_n10587_));
  OAI21_X1   g08151(.A1(new_n10587_), .A2(new_n10584_), .B(new_n2627_), .ZN(new_n10588_));
  AOI21_X1   g08152(.A1(new_n10588_), .A2(new_n3270_), .B(new_n10583_), .ZN(new_n10589_));
  OAI21_X1   g08153(.A1(new_n10589_), .A2(new_n10578_), .B(new_n7267_), .ZN(new_n10590_));
  OAI22_X1   g08154(.A1(new_n10590_), .A2(new_n10573_), .B1(new_n7267_), .B2(new_n10567_), .ZN(po0272));
  NOR3_X1    g08155(.A1(new_n8587_), .A2(pi0039), .A3(pi0072), .ZN(new_n10592_));
  INV_X1     g08156(.I(new_n10592_), .ZN(new_n10593_));
  OAI21_X1   g08157(.A1(new_n2626_), .A2(new_n10593_), .B(pi0075), .ZN(new_n10594_));
  NAND2_X1   g08158(.A1(new_n2821_), .A2(pi0115), .ZN(new_n10595_));
  NAND2_X1   g08159(.A1(new_n8370_), .A2(new_n10595_), .ZN(new_n10596_));
  AOI21_X1   g08160(.A1(new_n8726_), .A2(pi0115), .B(new_n8370_), .ZN(new_n10597_));
  NOR2_X1    g08161(.A1(new_n9000_), .A2(pi0052), .ZN(new_n10598_));
  NOR3_X1    g08162(.A1(new_n8556_), .A2(pi0115), .A3(new_n10598_), .ZN(new_n10599_));
  NAND2_X1   g08163(.A1(new_n10599_), .A2(new_n6706_), .ZN(new_n10600_));
  AOI21_X1   g08164(.A1(new_n10597_), .A2(new_n10600_), .B(new_n2659_), .ZN(new_n10601_));
  AOI21_X1   g08165(.A1(new_n10601_), .A2(new_n10596_), .B(new_n10594_), .ZN(new_n10602_));
  NOR2_X1    g08166(.A1(new_n10592_), .A2(new_n3270_), .ZN(new_n10603_));
  NOR2_X1    g08167(.A1(new_n8577_), .A2(new_n2458_), .ZN(new_n10604_));
  OAI21_X1   g08168(.A1(new_n10604_), .A2(new_n10595_), .B(new_n3270_), .ZN(new_n10605_));
  NOR2_X1    g08169(.A1(new_n8650_), .A2(pi0115), .ZN(new_n10606_));
  OAI21_X1   g08170(.A1(new_n10605_), .A2(new_n10606_), .B(new_n9082_), .ZN(new_n10607_));
  OAI21_X1   g08171(.A1(new_n10607_), .A2(new_n10603_), .B(new_n3465_), .ZN(new_n10608_));
  OAI21_X1   g08172(.A1(new_n8580_), .A2(new_n8587_), .B(new_n8369_), .ZN(new_n10609_));
  OAI21_X1   g08173(.A1(new_n10609_), .A2(new_n10599_), .B(new_n2627_), .ZN(new_n10610_));
  AOI21_X1   g08174(.A1(new_n8370_), .A2(new_n10595_), .B(new_n10610_), .ZN(new_n10611_));
  AOI21_X1   g08175(.A1(new_n10593_), .A2(pi0038), .B(pi0087), .ZN(new_n10612_));
  OAI21_X1   g08176(.A1(new_n10611_), .A2(new_n8667_), .B(new_n10612_), .ZN(new_n10613_));
  NOR2_X1    g08177(.A1(new_n8757_), .A2(new_n8587_), .ZN(new_n10614_));
  NOR2_X1    g08178(.A1(new_n8749_), .A2(pi0115), .ZN(new_n10615_));
  OAI21_X1   g08179(.A1(new_n10614_), .A2(new_n10615_), .B(new_n2627_), .ZN(new_n10616_));
  AOI21_X1   g08180(.A1(new_n10616_), .A2(new_n3270_), .B(new_n10613_), .ZN(new_n10617_));
  OAI21_X1   g08181(.A1(new_n10617_), .A2(new_n10608_), .B(new_n7267_), .ZN(new_n10618_));
  OAI22_X1   g08182(.A1(new_n10618_), .A2(new_n10602_), .B1(new_n7267_), .B2(new_n10593_), .ZN(po0273));
  NOR2_X1    g08183(.A1(new_n8596_), .A2(pi0039), .ZN(new_n10620_));
  INV_X1     g08184(.I(new_n10620_), .ZN(new_n10621_));
  INV_X1     g08185(.I(new_n10538_), .ZN(new_n10622_));
  NOR2_X1    g08186(.A1(new_n8549_), .A2(pi0113), .ZN(new_n10623_));
  OAI22_X1   g08187(.A1(new_n10623_), .A2(new_n8596_), .B1(new_n6707_), .B2(new_n8556_), .ZN(new_n10624_));
  NOR2_X1    g08188(.A1(new_n8369_), .A2(new_n8596_), .ZN(new_n10625_));
  AOI21_X1   g08189(.A1(new_n10624_), .A2(new_n10622_), .B(new_n10625_), .ZN(new_n10626_));
  AOI21_X1   g08190(.A1(new_n5792_), .A2(new_n10620_), .B(new_n3465_), .ZN(new_n10627_));
  OAI21_X1   g08191(.A1(new_n10626_), .A2(new_n2659_), .B(new_n10627_), .ZN(new_n10628_));
  NAND2_X1   g08192(.A1(new_n10621_), .A2(new_n3271_), .ZN(new_n10629_));
  NAND2_X1   g08193(.A1(new_n8647_), .A2(new_n8597_), .ZN(new_n10630_));
  NAND2_X1   g08194(.A1(new_n10630_), .A2(new_n8595_), .ZN(new_n10631_));
  NAND4_X1   g08195(.A1(new_n10631_), .A2(new_n3265_), .A3(new_n2702_), .A4(new_n8650_), .ZN(new_n10632_));
  NAND3_X1   g08196(.A1(new_n10632_), .A2(new_n9082_), .A3(new_n10629_), .ZN(new_n10633_));
  OAI21_X1   g08197(.A1(new_n10620_), .A2(new_n3265_), .B(new_n3458_), .ZN(new_n10634_));
  OAI21_X1   g08198(.A1(new_n10557_), .A2(pi0113), .B(new_n8595_), .ZN(new_n10635_));
  AOI21_X1   g08199(.A1(new_n10635_), .A2(new_n8556_), .B(new_n10538_), .ZN(new_n10636_));
  OAI21_X1   g08200(.A1(new_n10636_), .A2(new_n10625_), .B(new_n2627_), .ZN(new_n10637_));
  AOI21_X1   g08201(.A1(new_n10637_), .A2(new_n8489_), .B(new_n10634_), .ZN(new_n10638_));
  OAI21_X1   g08202(.A1(new_n8603_), .A2(new_n8594_), .B(new_n2458_), .ZN(new_n10639_));
  NOR2_X1    g08203(.A1(new_n10639_), .A2(new_n8591_), .ZN(new_n10640_));
  OAI21_X1   g08204(.A1(new_n8617_), .A2(new_n3026_), .B(pi0116), .ZN(new_n10641_));
  NAND2_X1   g08205(.A1(new_n10641_), .A2(new_n8612_), .ZN(new_n10642_));
  OAI21_X1   g08206(.A1(new_n8623_), .A2(new_n8594_), .B(new_n3026_), .ZN(new_n10643_));
  OAI21_X1   g08207(.A1(new_n8630_), .A2(new_n3025_), .B(pi0228), .ZN(new_n10644_));
  AOI21_X1   g08208(.A1(new_n10642_), .A2(new_n10643_), .B(new_n10644_), .ZN(new_n10645_));
  NOR3_X1    g08209(.A1(new_n10645_), .A2(pi0039), .A3(new_n10640_), .ZN(new_n10646_));
  OAI21_X1   g08210(.A1(new_n10646_), .A2(new_n3271_), .B(new_n10638_), .ZN(new_n10647_));
  NAND3_X1   g08211(.A1(new_n10647_), .A2(new_n3465_), .A3(new_n10633_), .ZN(new_n10648_));
  NAND3_X1   g08212(.A1(new_n10648_), .A2(new_n7267_), .A3(new_n10628_), .ZN(new_n10649_));
  OAI21_X1   g08213(.A1(new_n7267_), .A2(new_n10621_), .B(new_n10649_), .ZN(po0274));
  INV_X1     g08214(.I(new_n5298_), .ZN(new_n10651_));
  NOR2_X1    g08215(.A1(new_n6179_), .A2(pi0054), .ZN(new_n10652_));
  INV_X1     g08216(.I(new_n6214_), .ZN(new_n10653_));
  OAI22_X1   g08217(.A1(new_n3452_), .A2(pi0100), .B1(pi0039), .B2(new_n10653_), .ZN(new_n10654_));
  AOI21_X1   g08218(.A1(new_n10654_), .A2(new_n3265_), .B(pi0087), .ZN(new_n10655_));
  OAI21_X1   g08219(.A1(new_n10655_), .A2(new_n5304_), .B(new_n3444_), .ZN(new_n10656_));
  NAND3_X1   g08220(.A1(new_n10656_), .A2(new_n7263_), .A3(new_n10652_), .ZN(new_n10657_));
  NAND2_X1   g08221(.A1(new_n6169_), .A2(pi0055), .ZN(new_n10658_));
  NAND3_X1   g08222(.A1(new_n10657_), .A2(new_n3284_), .A3(new_n10658_), .ZN(new_n10659_));
  AOI21_X1   g08223(.A1(new_n10659_), .A2(new_n10651_), .B(pi0062), .ZN(new_n10660_));
  NOR3_X1    g08224(.A1(new_n10660_), .A2(new_n3425_), .A3(new_n5464_), .ZN(po0275));
  NOR2_X1    g08225(.A1(new_n9386_), .A2(pi0079), .ZN(new_n10662_));
  INV_X1     g08226(.I(new_n10662_), .ZN(new_n10663_));
  INV_X1     g08227(.I(pi0118), .ZN(new_n10664_));
  INV_X1     g08228(.I(pi0165), .ZN(new_n10665_));
  NOR2_X1    g08229(.A1(new_n6698_), .A2(new_n10665_), .ZN(new_n10666_));
  NAND2_X1   g08230(.A1(new_n10666_), .A2(new_n7342_), .ZN(new_n10667_));
  NAND2_X1   g08231(.A1(new_n10667_), .A2(new_n3425_), .ZN(new_n10668_));
  INV_X1     g08232(.I(new_n9388_), .ZN(new_n10669_));
  NOR2_X1    g08233(.A1(new_n9390_), .A2(new_n5437_), .ZN(new_n10670_));
  NAND4_X1   g08234(.A1(new_n10670_), .A2(new_n10669_), .A3(pi0150), .A4(new_n9392_), .ZN(new_n10671_));
  INV_X1     g08235(.I(pi0150), .ZN(new_n10672_));
  OAI21_X1   g08236(.A1(new_n9395_), .A2(new_n9393_), .B(new_n10672_), .ZN(new_n10673_));
  NAND2_X1   g08237(.A1(new_n10673_), .A2(new_n10671_), .ZN(new_n10674_));
  NAND3_X1   g08238(.A1(new_n10674_), .A2(pi0232), .A3(new_n7348_), .ZN(new_n10675_));
  NAND2_X1   g08239(.A1(new_n7342_), .A2(new_n2625_), .ZN(new_n10676_));
  AOI21_X1   g08240(.A1(new_n10675_), .A2(new_n10676_), .B(new_n10668_), .ZN(new_n10677_));
  INV_X1     g08241(.I(new_n10675_), .ZN(new_n10678_));
  AOI21_X1   g08242(.A1(new_n3265_), .A2(new_n5499_), .B(new_n10666_), .ZN(new_n10679_));
  INV_X1     g08243(.I(new_n10679_), .ZN(new_n10680_));
  NOR2_X1    g08244(.A1(new_n6698_), .A2(new_n10672_), .ZN(new_n10681_));
  NOR2_X1    g08245(.A1(new_n7601_), .A2(pi0092), .ZN(new_n10682_));
  NAND2_X1   g08246(.A1(new_n10682_), .A2(new_n10681_), .ZN(new_n10683_));
  NAND4_X1   g08247(.A1(new_n10683_), .A2(new_n3265_), .A3(new_n5499_), .A4(new_n7568_), .ZN(new_n10684_));
  AOI21_X1   g08248(.A1(new_n10684_), .A2(new_n10680_), .B(new_n10676_), .ZN(new_n10685_));
  OAI21_X1   g08249(.A1(new_n10685_), .A2(new_n10678_), .B(pi0055), .ZN(new_n10686_));
  NAND2_X1   g08250(.A1(new_n10674_), .A2(pi0299), .ZN(new_n10687_));
  INV_X1     g08251(.I(pi0185), .ZN(new_n10688_));
  XOR2_X1    g08252(.A1(new_n9429_), .A2(new_n10688_), .Z(new_n10689_));
  NAND3_X1   g08253(.A1(new_n10689_), .A2(new_n2628_), .A3(new_n5398_), .ZN(new_n10690_));
  NAND2_X1   g08254(.A1(new_n10690_), .A2(new_n10687_), .ZN(new_n10691_));
  NAND3_X1   g08255(.A1(new_n10691_), .A2(pi0232), .A3(new_n7348_), .ZN(new_n10692_));
  AOI21_X1   g08256(.A1(new_n10692_), .A2(pi0074), .B(pi0055), .ZN(new_n10693_));
  NOR2_X1    g08257(.A1(new_n10665_), .A2(new_n2628_), .ZN(new_n10694_));
  INV_X1     g08258(.I(pi0143), .ZN(new_n10695_));
  NOR2_X1    g08259(.A1(new_n10695_), .A2(pi0299), .ZN(new_n10696_));
  OAI21_X1   g08260(.A1(new_n10694_), .A2(new_n10696_), .B(new_n6697_), .ZN(new_n10697_));
  INV_X1     g08261(.I(new_n10697_), .ZN(new_n10698_));
  OAI21_X1   g08262(.A1(new_n7348_), .A2(new_n10698_), .B(new_n10692_), .ZN(new_n10699_));
  NOR2_X1    g08263(.A1(new_n10699_), .A2(new_n5499_), .ZN(new_n10700_));
  NAND2_X1   g08264(.A1(new_n10691_), .A2(pi0232), .ZN(new_n10701_));
  NAND2_X1   g08265(.A1(new_n10701_), .A2(pi0100), .ZN(new_n10702_));
  NOR2_X1    g08266(.A1(new_n10698_), .A2(new_n3265_), .ZN(new_n10703_));
  NOR2_X1    g08267(.A1(new_n10703_), .A2(pi0100), .ZN(new_n10704_));
  INV_X1     g08268(.I(new_n10704_), .ZN(new_n10705_));
  NOR2_X1    g08269(.A1(pi0178), .A2(pi0299), .ZN(new_n10706_));
  NOR2_X1    g08270(.A1(new_n2628_), .A2(pi0157), .ZN(new_n10707_));
  NOR3_X1    g08271(.A1(new_n6698_), .A2(new_n10706_), .A3(new_n10707_), .ZN(new_n10708_));
  AOI21_X1   g08272(.A1(new_n7600_), .A2(new_n10708_), .B(new_n7585_), .ZN(new_n10709_));
  OAI21_X1   g08273(.A1(new_n10709_), .A2(new_n10705_), .B(new_n10702_), .ZN(new_n10710_));
  AOI22_X1   g08274(.A1(new_n10710_), .A2(new_n7387_), .B1(pi0075), .B2(new_n10701_), .ZN(new_n10711_));
  NOR2_X1    g08275(.A1(new_n7405_), .A2(new_n10695_), .ZN(new_n10712_));
  AOI21_X1   g08276(.A1(new_n10712_), .A2(new_n10665_), .B(new_n3265_), .ZN(new_n10713_));
  NOR2_X1    g08277(.A1(new_n7398_), .A2(new_n10695_), .ZN(new_n10714_));
  NOR2_X1    g08278(.A1(new_n7401_), .A2(pi0143), .ZN(new_n10715_));
  OAI21_X1   g08279(.A1(new_n10715_), .A2(new_n10714_), .B(pi0165), .ZN(new_n10716_));
  AOI21_X1   g08280(.A1(new_n10713_), .A2(new_n10716_), .B(new_n2604_), .ZN(new_n10717_));
  AOI21_X1   g08281(.A1(new_n7568_), .A2(new_n5666_), .B(new_n2627_), .ZN(new_n10718_));
  AOI21_X1   g08282(.A1(new_n5446_), .A2(new_n7583_), .B(new_n7525_), .ZN(new_n10719_));
  NAND3_X1   g08283(.A1(new_n7639_), .A2(pi0178), .A3(new_n10719_), .ZN(new_n10720_));
  INV_X1     g08284(.I(pi0190), .ZN(new_n10721_));
  NOR2_X1    g08285(.A1(new_n10721_), .A2(pi0299), .ZN(new_n10722_));
  NAND3_X1   g08286(.A1(new_n10720_), .A2(new_n7613_), .A3(new_n10722_), .ZN(new_n10723_));
  INV_X1     g08287(.I(pi0178), .ZN(new_n10724_));
  NAND2_X1   g08288(.A1(new_n10719_), .A2(new_n10724_), .ZN(new_n10725_));
  NOR2_X1    g08289(.A1(new_n7616_), .A2(new_n10725_), .ZN(new_n10726_));
  OAI21_X1   g08290(.A1(new_n10723_), .A2(new_n10726_), .B(pi0232), .ZN(new_n10727_));
  NAND2_X1   g08291(.A1(new_n7647_), .A2(pi0178), .ZN(new_n10728_));
  NAND2_X1   g08292(.A1(new_n10728_), .A2(new_n10721_), .ZN(new_n10729_));
  INV_X1     g08293(.I(new_n10706_), .ZN(new_n10730_));
  AOI22_X1   g08294(.A1(pi0157), .A2(new_n7626_), .B1(new_n7614_), .B2(pi0168), .ZN(new_n10731_));
  NOR4_X1    g08295(.A1(new_n10731_), .A2(new_n5437_), .A3(new_n5422_), .A4(new_n8070_), .ZN(new_n10732_));
  OAI21_X1   g08296(.A1(new_n10732_), .A2(new_n2628_), .B(new_n10730_), .ZN(new_n10733_));
  AOI22_X1   g08297(.A1(new_n10729_), .A2(new_n2628_), .B1(new_n7568_), .B2(new_n10733_), .ZN(new_n10734_));
  OAI21_X1   g08298(.A1(new_n10727_), .A2(new_n10734_), .B(new_n10718_), .ZN(new_n10735_));
  INV_X1     g08299(.I(pi0173), .ZN(new_n10736_));
  NOR2_X1    g08300(.A1(new_n7726_), .A2(new_n5398_), .ZN(new_n10737_));
  NOR2_X1    g08301(.A1(new_n7704_), .A2(new_n10737_), .ZN(new_n10738_));
  NOR2_X1    g08302(.A1(new_n10738_), .A2(new_n10736_), .ZN(new_n10739_));
  NOR2_X1    g08303(.A1(new_n7726_), .A2(pi0173), .ZN(new_n10740_));
  OAI21_X1   g08304(.A1(new_n10739_), .A2(new_n10740_), .B(new_n10688_), .ZN(new_n10741_));
  NAND2_X1   g08305(.A1(new_n7726_), .A2(new_n5437_), .ZN(new_n10742_));
  INV_X1     g08306(.I(new_n10742_), .ZN(new_n10743_));
  NAND2_X1   g08307(.A1(new_n7883_), .A2(new_n10736_), .ZN(new_n10744_));
  OAI21_X1   g08308(.A1(new_n10736_), .A2(new_n8002_), .B(new_n10744_), .ZN(new_n10745_));
  AOI21_X1   g08309(.A1(new_n10745_), .A2(new_n5398_), .B(new_n10743_), .ZN(new_n10746_));
  AOI21_X1   g08310(.A1(new_n10746_), .A2(pi0185), .B(pi0190), .ZN(new_n10747_));
  AOI21_X1   g08311(.A1(new_n10747_), .A2(new_n10741_), .B(pi0299), .ZN(new_n10748_));
  AOI21_X1   g08312(.A1(new_n7880_), .A2(new_n10742_), .B(pi0173), .ZN(new_n10749_));
  NOR2_X1    g08313(.A1(new_n7834_), .A2(new_n5437_), .ZN(new_n10750_));
  NOR3_X1    g08314(.A1(new_n10750_), .A2(new_n10736_), .A3(new_n10737_), .ZN(new_n10751_));
  NOR3_X1    g08315(.A1(new_n10749_), .A2(new_n10688_), .A3(new_n10751_), .ZN(new_n10752_));
  NOR3_X1    g08316(.A1(new_n10743_), .A2(new_n7877_), .A3(pi0173), .ZN(new_n10753_));
  OR2_X2     g08317(.A1(new_n7713_), .A2(new_n10737_), .Z(new_n10754_));
  AOI21_X1   g08318(.A1(new_n10754_), .A2(pi0173), .B(new_n10753_), .ZN(new_n10755_));
  OAI21_X1   g08319(.A1(new_n10755_), .A2(pi0185), .B(pi0190), .ZN(new_n10756_));
  OAI21_X1   g08320(.A1(new_n10752_), .A2(new_n10756_), .B(new_n10748_), .ZN(new_n10757_));
  NAND2_X1   g08321(.A1(new_n7877_), .A2(pi0168), .ZN(new_n10758_));
  NOR2_X1    g08322(.A1(new_n5437_), .A2(new_n4571_), .ZN(new_n10759_));
  INV_X1     g08323(.I(new_n10759_), .ZN(new_n10760_));
  NAND2_X1   g08324(.A1(new_n7726_), .A2(new_n10760_), .ZN(new_n10761_));
  NAND3_X1   g08325(.A1(new_n10758_), .A2(new_n3533_), .A3(new_n10761_), .ZN(new_n10762_));
  NAND2_X1   g08326(.A1(new_n10754_), .A2(pi0168), .ZN(new_n10763_));
  OAI21_X1   g08327(.A1(pi0168), .A2(new_n10738_), .B(new_n10763_), .ZN(new_n10764_));
  AOI21_X1   g08328(.A1(new_n10764_), .A2(pi0151), .B(pi0150), .ZN(new_n10765_));
  AOI21_X1   g08329(.A1(new_n10765_), .A2(new_n10762_), .B(new_n2628_), .ZN(new_n10766_));
  NOR2_X1    g08330(.A1(new_n7691_), .A2(new_n5437_), .ZN(new_n10767_));
  OAI21_X1   g08331(.A1(new_n10767_), .A2(new_n10737_), .B(pi0151), .ZN(new_n10768_));
  NOR2_X1    g08332(.A1(new_n10768_), .A2(new_n4571_), .ZN(new_n10769_));
  NAND2_X1   g08333(.A1(new_n7821_), .A2(pi0168), .ZN(new_n10770_));
  NAND2_X1   g08334(.A1(new_n7827_), .A2(new_n4571_), .ZN(new_n10771_));
  AOI21_X1   g08335(.A1(new_n10770_), .A2(new_n10771_), .B(pi0151), .ZN(new_n10772_));
  NOR3_X1    g08336(.A1(new_n8035_), .A2(new_n3533_), .A3(pi0168), .ZN(new_n10773_));
  OAI21_X1   g08337(.A1(new_n10772_), .A2(new_n10773_), .B(new_n10742_), .ZN(new_n10774_));
  NAND2_X1   g08338(.A1(new_n10774_), .A2(pi0150), .ZN(new_n10775_));
  OAI21_X1   g08339(.A1(new_n10775_), .A2(new_n10769_), .B(new_n10766_), .ZN(new_n10776_));
  NAND3_X1   g08340(.A1(new_n10776_), .A2(pi0232), .A3(new_n10757_), .ZN(new_n10777_));
  NAND2_X1   g08341(.A1(new_n7726_), .A2(new_n5666_), .ZN(new_n10778_));
  NAND3_X1   g08342(.A1(new_n10777_), .A2(new_n2627_), .A3(new_n10778_), .ZN(new_n10779_));
  NAND3_X1   g08343(.A1(new_n10779_), .A2(new_n3265_), .A3(new_n10735_), .ZN(new_n10780_));
  OAI21_X1   g08344(.A1(new_n10698_), .A2(new_n3265_), .B(new_n6800_), .ZN(new_n10781_));
  OAI21_X1   g08345(.A1(new_n7584_), .A2(new_n10781_), .B(new_n10702_), .ZN(new_n10782_));
  AOI21_X1   g08346(.A1(new_n10780_), .A2(new_n10717_), .B(new_n10782_), .ZN(new_n10783_));
  OAI21_X1   g08347(.A1(new_n10783_), .A2(new_n2606_), .B(new_n10711_), .ZN(new_n10784_));
  AOI21_X1   g08348(.A1(new_n10784_), .A2(new_n5499_), .B(new_n10700_), .ZN(new_n10785_));
  OAI21_X1   g08349(.A1(new_n10785_), .A2(pi0074), .B(new_n10693_), .ZN(new_n10786_));
  NAND3_X1   g08350(.A1(new_n10786_), .A2(new_n2470_), .A3(new_n10686_), .ZN(new_n10787_));
  INV_X1     g08351(.I(new_n8103_), .ZN(new_n10788_));
  NAND2_X1   g08352(.A1(new_n10679_), .A2(new_n7342_), .ZN(new_n10789_));
  OAI21_X1   g08353(.A1(pi0074), .A2(new_n10789_), .B(new_n10675_), .ZN(new_n10790_));
  OAI21_X1   g08354(.A1(new_n10790_), .A2(new_n2470_), .B(new_n3291_), .ZN(new_n10791_));
  NAND2_X1   g08355(.A1(new_n10791_), .A2(new_n10788_), .ZN(new_n10792_));
  AOI21_X1   g08356(.A1(new_n10787_), .A2(new_n10792_), .B(new_n10677_), .ZN(new_n10793_));
  NAND2_X1   g08357(.A1(new_n10675_), .A2(pi0074), .ZN(new_n10794_));
  NOR4_X1    g08358(.A1(new_n10681_), .A2(pi0092), .A3(new_n2657_), .A4(new_n7348_), .ZN(new_n10795_));
  NAND2_X1   g08359(.A1(new_n10666_), .A2(pi0054), .ZN(new_n10796_));
  NAND3_X1   g08360(.A1(new_n2531_), .A2(new_n10795_), .A3(new_n10796_), .ZN(new_n10797_));
  NAND4_X1   g08361(.A1(new_n10675_), .A2(new_n2625_), .A3(new_n10789_), .A4(new_n10797_), .ZN(new_n10798_));
  NAND3_X1   g08362(.A1(new_n10798_), .A2(pi0055), .A3(new_n10794_), .ZN(new_n10799_));
  NAND2_X1   g08363(.A1(new_n10701_), .A2(pi0075), .ZN(new_n10800_));
  NOR3_X1    g08364(.A1(new_n2530_), .A2(new_n2657_), .A3(new_n10708_), .ZN(new_n10801_));
  OAI21_X1   g08365(.A1(new_n10705_), .A2(new_n10801_), .B(new_n10702_), .ZN(new_n10802_));
  NOR2_X1    g08366(.A1(new_n7496_), .A2(new_n5351_), .ZN(new_n10803_));
  NOR2_X1    g08367(.A1(new_n10803_), .A2(pi0232), .ZN(new_n10804_));
  NAND3_X1   g08368(.A1(new_n7462_), .A2(new_n10736_), .A3(pi0190), .ZN(new_n10805_));
  NAND2_X1   g08369(.A1(new_n7465_), .A2(new_n10736_), .ZN(new_n10806_));
  OAI21_X1   g08370(.A1(new_n10736_), .A2(new_n7471_), .B(new_n10806_), .ZN(new_n10807_));
  NAND4_X1   g08371(.A1(new_n10807_), .A2(new_n10721_), .A3(new_n2535_), .A4(new_n5398_), .ZN(new_n10808_));
  NAND3_X1   g08372(.A1(new_n10808_), .A2(pi0185), .A3(new_n10805_), .ZN(new_n10809_));
  NAND2_X1   g08373(.A1(new_n7442_), .A2(new_n10736_), .ZN(new_n10810_));
  AOI21_X1   g08374(.A1(new_n10810_), .A2(new_n7481_), .B(pi0190), .ZN(new_n10811_));
  OAI21_X1   g08375(.A1(new_n7482_), .A2(new_n10736_), .B(pi0190), .ZN(new_n10812_));
  OAI21_X1   g08376(.A1(new_n7491_), .A2(new_n10812_), .B(new_n10688_), .ZN(new_n10813_));
  OAI21_X1   g08377(.A1(new_n10811_), .A2(new_n10813_), .B(new_n10809_), .ZN(new_n10814_));
  AOI21_X1   g08378(.A1(new_n9685_), .A2(new_n5437_), .B(pi0299), .ZN(new_n10815_));
  NAND2_X1   g08379(.A1(new_n10814_), .A2(new_n10815_), .ZN(new_n10816_));
  NAND2_X1   g08380(.A1(new_n7442_), .A2(new_n3533_), .ZN(new_n10817_));
  NAND2_X1   g08381(.A1(new_n10817_), .A2(new_n7436_), .ZN(new_n10818_));
  NOR2_X1    g08382(.A1(new_n8123_), .A2(pi0151), .ZN(new_n10819_));
  OAI21_X1   g08383(.A1(new_n10819_), .A2(new_n8122_), .B(new_n10759_), .ZN(new_n10820_));
  NAND2_X1   g08384(.A1(new_n10820_), .A2(new_n10672_), .ZN(new_n10821_));
  AOI21_X1   g08385(.A1(new_n10818_), .A2(new_n4571_), .B(new_n10821_), .ZN(new_n10822_));
  NAND2_X1   g08386(.A1(new_n7460_), .A2(pi0168), .ZN(new_n10823_));
  NAND2_X1   g08387(.A1(new_n7465_), .A2(new_n4571_), .ZN(new_n10824_));
  AOI21_X1   g08388(.A1(new_n10824_), .A2(new_n10823_), .B(pi0151), .ZN(new_n10825_));
  NOR3_X1    g08389(.A1(new_n7471_), .A2(new_n3533_), .A3(pi0168), .ZN(new_n10826_));
  OAI21_X1   g08390(.A1(new_n10825_), .A2(new_n10826_), .B(new_n7457_), .ZN(new_n10827_));
  AOI21_X1   g08391(.A1(pi0150), .A2(new_n10827_), .B(new_n10822_), .ZN(new_n10828_));
  AOI21_X1   g08392(.A1(new_n9707_), .A2(new_n7441_), .B(new_n5398_), .ZN(new_n10829_));
  OR3_X2     g08393(.A1(new_n10828_), .A2(new_n2628_), .A3(new_n10829_), .Z(new_n10830_));
  NAND2_X1   g08394(.A1(new_n10830_), .A2(new_n10816_), .ZN(new_n10831_));
  AOI22_X1   g08395(.A1(new_n10831_), .A2(pi0232), .B1(new_n7441_), .B2(new_n10804_), .ZN(new_n10832_));
  NOR2_X1    g08396(.A1(new_n5551_), .A2(new_n6745_), .ZN(new_n10833_));
  INV_X1     g08397(.I(pi0157), .ZN(new_n10834_));
  NAND2_X1   g08398(.A1(new_n10834_), .A2(new_n4571_), .ZN(new_n10835_));
  OAI22_X1   g08399(.A1(new_n7509_), .A2(new_n10835_), .B1(new_n10834_), .B2(new_n7511_), .ZN(new_n10836_));
  AOI21_X1   g08400(.A1(new_n7514_), .A2(new_n10834_), .B(new_n4571_), .ZN(new_n10837_));
  NOR2_X1    g08401(.A1(new_n10837_), .A2(new_n10836_), .ZN(new_n10838_));
  OAI21_X1   g08402(.A1(new_n10838_), .A2(new_n10833_), .B(new_n10332_), .ZN(new_n10839_));
  NAND2_X1   g08403(.A1(new_n10363_), .A2(new_n10724_), .ZN(new_n10840_));
  NAND2_X1   g08404(.A1(new_n10840_), .A2(new_n10721_), .ZN(new_n10841_));
  NOR3_X1    g08405(.A1(new_n10833_), .A2(new_n10724_), .A3(new_n7521_), .ZN(new_n10842_));
  NOR2_X1    g08406(.A1(new_n6751_), .A2(new_n7520_), .ZN(new_n10843_));
  AOI21_X1   g08407(.A1(new_n10843_), .A2(new_n10724_), .B(new_n10833_), .ZN(new_n10844_));
  OAI22_X1   g08408(.A1(new_n10844_), .A2(new_n10721_), .B1(new_n10841_), .B2(new_n10842_), .ZN(new_n10845_));
  AOI21_X1   g08409(.A1(new_n10845_), .A2(new_n10333_), .B(new_n5666_), .ZN(new_n10846_));
  NAND3_X1   g08410(.A1(new_n5536_), .A2(new_n5423_), .A3(new_n10332_), .ZN(new_n10847_));
  NAND2_X1   g08411(.A1(new_n10847_), .A2(new_n5666_), .ZN(new_n10848_));
  INV_X1     g08412(.I(new_n10333_), .ZN(new_n10849_));
  NOR2_X1    g08413(.A1(new_n10363_), .A2(new_n10849_), .ZN(new_n10850_));
  OAI21_X1   g08414(.A1(new_n10848_), .A2(new_n10850_), .B(pi0039), .ZN(new_n10851_));
  AOI21_X1   g08415(.A1(new_n10846_), .A2(new_n10839_), .B(new_n10851_), .ZN(new_n10852_));
  AOI21_X1   g08416(.A1(new_n10832_), .A2(new_n2627_), .B(new_n10852_), .ZN(new_n10853_));
  OAI21_X1   g08417(.A1(new_n10853_), .A2(pi0038), .B(new_n10717_), .ZN(new_n10854_));
  NAND3_X1   g08418(.A1(new_n10854_), .A2(new_n10702_), .A3(new_n10781_), .ZN(new_n10855_));
  AOI22_X1   g08419(.A1(new_n10855_), .A2(new_n2605_), .B1(new_n7387_), .B2(new_n10802_), .ZN(new_n10856_));
  AOI21_X1   g08420(.A1(new_n10856_), .A2(new_n10800_), .B(pi0054), .ZN(new_n10857_));
  OAI21_X1   g08421(.A1(new_n10857_), .A2(new_n10700_), .B(new_n2625_), .ZN(new_n10858_));
  AOI21_X1   g08422(.A1(new_n10858_), .A2(new_n10693_), .B(new_n2471_), .ZN(new_n10859_));
  AOI21_X1   g08423(.A1(new_n10859_), .A2(new_n10799_), .B(new_n10791_), .ZN(new_n10860_));
  OR2_X2     g08424(.A1(new_n10860_), .A2(new_n10677_), .Z(new_n10861_));
  NAND2_X1   g08425(.A1(new_n10861_), .A2(new_n10664_), .ZN(new_n10862_));
  OAI21_X1   g08426(.A1(new_n10793_), .A2(new_n10664_), .B(new_n10862_), .ZN(new_n10863_));
  NAND2_X1   g08427(.A1(new_n10863_), .A2(new_n10663_), .ZN(new_n10864_));
  NAND2_X1   g08428(.A1(new_n7562_), .A2(new_n10664_), .ZN(new_n10865_));
  NOR2_X1    g08429(.A1(new_n10793_), .A2(new_n10865_), .ZN(new_n10866_));
  AOI21_X1   g08430(.A1(new_n10861_), .A2(new_n10865_), .B(new_n10866_), .ZN(new_n10867_));
  OAI21_X1   g08431(.A1(new_n10867_), .A2(new_n10663_), .B(new_n10864_), .ZN(po0276));
  NAND2_X1   g08432(.A1(pi0128), .A2(pi0228), .ZN(new_n10869_));
  INV_X1     g08433(.I(new_n6207_), .ZN(new_n10870_));
  AND3_X2    g08434(.A1(new_n10870_), .A2(pi0092), .A3(new_n10869_), .Z(new_n10871_));
  NOR2_X1    g08435(.A1(new_n3487_), .A2(new_n2659_), .ZN(new_n10872_));
  AOI21_X1   g08436(.A1(pi0128), .A2(pi0228), .B(new_n10872_), .ZN(new_n10873_));
  OAI21_X1   g08437(.A1(new_n10873_), .A2(new_n3465_), .B(new_n3444_), .ZN(new_n10874_));
  INV_X1     g08438(.I(new_n5562_), .ZN(new_n10875_));
  NAND2_X1   g08439(.A1(new_n5639_), .A2(pi0299), .ZN(new_n10876_));
  AOI21_X1   g08440(.A1(new_n10876_), .A2(new_n5664_), .B(new_n6698_), .ZN(new_n10877_));
  NAND2_X1   g08441(.A1(new_n10877_), .A2(new_n2734_), .ZN(new_n10878_));
  OAI21_X1   g08442(.A1(new_n10875_), .A2(new_n10877_), .B(new_n10878_), .ZN(new_n10879_));
  OAI22_X1   g08443(.A1(new_n9381_), .A2(new_n3086_), .B1(new_n2508_), .B2(new_n10877_), .ZN(new_n10880_));
  NOR2_X1    g08444(.A1(new_n10325_), .A2(new_n2856_), .ZN(new_n10881_));
  OAI21_X1   g08445(.A1(new_n9380_), .A2(new_n10881_), .B(new_n2878_), .ZN(new_n10882_));
  INV_X1     g08446(.I(new_n2865_), .ZN(new_n10883_));
  NAND4_X1   g08447(.A1(new_n10883_), .A2(new_n2511_), .A3(new_n2849_), .A4(new_n3086_), .ZN(new_n10884_));
  AOI21_X1   g08448(.A1(new_n10882_), .A2(new_n2864_), .B(new_n10884_), .ZN(new_n10885_));
  OAI21_X1   g08449(.A1(new_n10880_), .A2(new_n10885_), .B(new_n10879_), .ZN(new_n10886_));
  OAI21_X1   g08450(.A1(new_n10886_), .A2(pi0091), .B(new_n6718_), .ZN(new_n10887_));
  AOI21_X1   g08451(.A1(new_n10887_), .A2(new_n2763_), .B(new_n2989_), .ZN(new_n10888_));
  NOR3_X1    g08452(.A1(new_n10888_), .A2(pi0039), .A3(new_n9142_), .ZN(new_n10889_));
  NAND3_X1   g08453(.A1(new_n6805_), .A2(new_n2642_), .A3(new_n3335_), .ZN(new_n10890_));
  NAND3_X1   g08454(.A1(new_n10296_), .A2(new_n3304_), .A3(new_n5113_), .ZN(new_n10891_));
  AOI21_X1   g08455(.A1(new_n10890_), .A2(new_n10891_), .B(new_n2627_), .ZN(new_n10892_));
  OAI21_X1   g08456(.A1(new_n10889_), .A2(new_n10892_), .B(new_n3265_), .ZN(new_n10893_));
  OAI21_X1   g08457(.A1(new_n10893_), .A2(pi0228), .B(new_n2702_), .ZN(new_n10894_));
  OAI21_X1   g08458(.A1(new_n3487_), .A2(new_n2573_), .B(pi0100), .ZN(new_n10895_));
  NAND3_X1   g08459(.A1(new_n10894_), .A2(new_n3458_), .A3(new_n10895_), .ZN(new_n10896_));
  AOI21_X1   g08460(.A1(new_n10896_), .A2(new_n10869_), .B(pi0075), .ZN(new_n10897_));
  OAI21_X1   g08461(.A1(new_n10897_), .A2(new_n10874_), .B(new_n8255_), .ZN(new_n10898_));
  OAI22_X1   g08462(.A1(new_n10898_), .A2(new_n10871_), .B1(new_n8255_), .B2(new_n10869_), .ZN(po0277));
  INV_X1     g08463(.I(pi0031), .ZN(new_n10900_));
  NAND3_X1   g08464(.A1(new_n10900_), .A2(new_n9878_), .A3(pi0818), .ZN(new_n10901_));
  INV_X1     g08465(.I(new_n10901_), .ZN(new_n10902_));
  INV_X1     g08466(.I(pi0120), .ZN(new_n10903_));
  NOR2_X1    g08467(.A1(new_n10093_), .A2(new_n10903_), .ZN(new_n10904_));
  NOR2_X1    g08468(.A1(new_n3041_), .A2(pi0120), .ZN(new_n10905_));
  OAI21_X1   g08469(.A1(new_n9822_), .A2(pi1091), .B(new_n10905_), .ZN(new_n10906_));
  INV_X1     g08470(.I(new_n10906_), .ZN(new_n10907_));
  NOR2_X1    g08471(.A1(new_n10904_), .A2(new_n10907_), .ZN(new_n10908_));
  INV_X1     g08472(.I(new_n10908_), .ZN(new_n10909_));
  NOR2_X1    g08473(.A1(new_n10909_), .A2(new_n6349_), .ZN(new_n10910_));
  NOR2_X1    g08474(.A1(pi0120), .A2(pi1093), .ZN(new_n10911_));
  INV_X1     g08475(.I(new_n10911_), .ZN(new_n10912_));
  NAND2_X1   g08476(.A1(new_n10902_), .A2(new_n10912_), .ZN(new_n10913_));
  OAI21_X1   g08477(.A1(new_n10910_), .A2(new_n10913_), .B(po1038), .ZN(new_n10914_));
  NAND3_X1   g08478(.A1(pi0951), .A2(pi0982), .A3(pi1092), .ZN(new_n10915_));
  NOR2_X1    g08479(.A1(new_n10915_), .A2(new_n3041_), .ZN(new_n10916_));
  NOR2_X1    g08480(.A1(new_n10916_), .A2(pi0120), .ZN(new_n10917_));
  NOR2_X1    g08481(.A1(new_n10910_), .A2(new_n10917_), .ZN(new_n10918_));
  OAI21_X1   g08482(.A1(new_n10914_), .A2(new_n10918_), .B(new_n7253_), .ZN(new_n10919_));
  INV_X1     g08483(.I(new_n7253_), .ZN(new_n10920_));
  NOR2_X1    g08484(.A1(new_n10910_), .A2(new_n10903_), .ZN(new_n10921_));
  OAI21_X1   g08485(.A1(new_n10914_), .A2(new_n10921_), .B(new_n10920_), .ZN(new_n10922_));
  NAND2_X1   g08486(.A1(new_n10919_), .A2(new_n10922_), .ZN(new_n10923_));
  AOI21_X1   g08487(.A1(new_n10093_), .A2(new_n6648_), .B(new_n6349_), .ZN(new_n10924_));
  INV_X1     g08488(.I(new_n10924_), .ZN(new_n10925_));
  NOR2_X1    g08489(.A1(new_n6645_), .A2(new_n10912_), .ZN(new_n10926_));
  NOR2_X1    g08490(.A1(new_n10925_), .A2(new_n10926_), .ZN(new_n10927_));
  NOR2_X1    g08491(.A1(new_n10909_), .A2(new_n6700_), .ZN(new_n10928_));
  AOI21_X1   g08492(.A1(new_n3022_), .A2(new_n10092_), .B(new_n6709_), .ZN(new_n10929_));
  OAI21_X1   g08493(.A1(new_n10929_), .A2(new_n10903_), .B(new_n8224_), .ZN(new_n10930_));
  AND2_X2    g08494(.A1(new_n6797_), .A2(new_n10907_), .Z(new_n10931_));
  NOR3_X1    g08495(.A1(new_n10930_), .A2(new_n2659_), .A3(new_n10931_), .ZN(new_n10932_));
  NOR3_X1    g08496(.A1(new_n10932_), .A2(new_n3465_), .A3(new_n10928_), .ZN(new_n10933_));
  NOR2_X1    g08497(.A1(new_n6776_), .A2(new_n10903_), .ZN(new_n10934_));
  NAND2_X1   g08498(.A1(new_n6775_), .A2(pi1091), .ZN(new_n10935_));
  AOI21_X1   g08499(.A1(new_n6776_), .A2(new_n10904_), .B(new_n10935_), .ZN(new_n10936_));
  OAI21_X1   g08500(.A1(new_n10936_), .A2(new_n10934_), .B(new_n6820_), .ZN(new_n10937_));
  NAND2_X1   g08501(.A1(new_n10937_), .A2(pi0100), .ZN(new_n10938_));
  NAND3_X1   g08502(.A1(new_n6748_), .A2(pi1091), .A3(pi1092), .ZN(new_n10939_));
  AOI22_X1   g08503(.A1(new_n6751_), .A2(new_n10904_), .B1(new_n10907_), .B2(new_n10939_), .ZN(new_n10940_));
  NAND2_X1   g08504(.A1(new_n10909_), .A2(new_n6745_), .ZN(new_n10941_));
  OAI21_X1   g08505(.A1(new_n10940_), .A2(new_n6745_), .B(new_n10941_), .ZN(new_n10942_));
  NOR2_X1    g08506(.A1(new_n10942_), .A2(new_n6764_), .ZN(new_n10943_));
  NOR2_X1    g08507(.A1(new_n10909_), .A2(new_n5427_), .ZN(new_n10944_));
  AOI21_X1   g08508(.A1(new_n10940_), .A2(new_n5427_), .B(new_n10944_), .ZN(new_n10945_));
  NOR2_X1    g08509(.A1(new_n10945_), .A2(new_n5422_), .ZN(new_n10946_));
  OAI21_X1   g08510(.A1(new_n10946_), .A2(new_n10943_), .B(new_n6761_), .ZN(new_n10947_));
  AOI21_X1   g08511(.A1(new_n10908_), .A2(new_n6762_), .B(new_n2628_), .ZN(new_n10948_));
  NOR2_X1    g08512(.A1(new_n10942_), .A2(new_n5445_), .ZN(new_n10949_));
  NOR2_X1    g08513(.A1(new_n10945_), .A2(new_n5446_), .ZN(new_n10950_));
  OAI21_X1   g08514(.A1(new_n10950_), .A2(new_n10949_), .B(new_n6744_), .ZN(new_n10951_));
  AOI21_X1   g08515(.A1(new_n10908_), .A2(new_n6759_), .B(pi0299), .ZN(new_n10952_));
  AOI22_X1   g08516(.A1(new_n10947_), .A2(new_n10948_), .B1(new_n10951_), .B2(new_n10952_), .ZN(new_n10953_));
  NOR2_X1    g08517(.A1(new_n6688_), .A2(new_n6714_), .ZN(new_n10954_));
  NOR2_X1    g08518(.A1(new_n10954_), .A2(new_n3024_), .ZN(new_n10955_));
  NOR2_X1    g08519(.A1(new_n6687_), .A2(new_n6259_), .ZN(new_n10956_));
  AOI21_X1   g08520(.A1(new_n10956_), .A2(new_n3044_), .B(pi0122), .ZN(new_n10957_));
  OAI21_X1   g08521(.A1(new_n6729_), .A2(new_n8457_), .B(new_n10957_), .ZN(new_n10958_));
  AOI21_X1   g08522(.A1(new_n10958_), .A2(new_n10955_), .B(new_n3081_), .ZN(new_n10959_));
  NOR2_X1    g08523(.A1(new_n10956_), .A2(new_n6871_), .ZN(new_n10960_));
  AOI21_X1   g08524(.A1(new_n9822_), .A2(new_n10960_), .B(new_n10959_), .ZN(new_n10961_));
  NAND2_X1   g08525(.A1(new_n6689_), .A2(new_n3041_), .ZN(new_n10962_));
  INV_X1     g08526(.I(new_n10962_), .ZN(new_n10963_));
  AOI21_X1   g08527(.A1(new_n10963_), .A2(pi0120), .B(pi0039), .ZN(new_n10964_));
  AOI22_X1   g08528(.A1(new_n10961_), .A2(new_n10964_), .B1(pi0039), .B2(new_n10953_), .ZN(new_n10965_));
  NOR2_X1    g08529(.A1(new_n10965_), .A2(pi0038), .ZN(new_n10966_));
  OAI21_X1   g08530(.A1(new_n10093_), .A2(new_n10911_), .B(pi0038), .ZN(new_n10967_));
  NAND2_X1   g08531(.A1(new_n10967_), .A2(new_n2702_), .ZN(new_n10968_));
  OAI22_X1   g08532(.A1(new_n10966_), .A2(new_n10968_), .B1(new_n10908_), .B2(new_n10938_), .ZN(new_n10969_));
  OAI21_X1   g08533(.A1(new_n2531_), .A2(new_n6714_), .B(new_n6258_), .ZN(new_n10970_));
  NAND2_X1   g08534(.A1(new_n10970_), .A2(new_n6870_), .ZN(new_n10971_));
  NAND3_X1   g08535(.A1(new_n6873_), .A2(new_n10971_), .A3(new_n3272_), .ZN(new_n10972_));
  AOI21_X1   g08536(.A1(new_n10093_), .A2(new_n3273_), .B(new_n3458_), .ZN(new_n10973_));
  NAND2_X1   g08537(.A1(new_n10972_), .A2(new_n10973_), .ZN(new_n10974_));
  OR2_X2     g08538(.A1(new_n6875_), .A2(new_n10911_), .Z(new_n10975_));
  NOR2_X1    g08539(.A1(new_n10975_), .A2(new_n10974_), .ZN(new_n10976_));
  AOI21_X1   g08540(.A1(new_n10969_), .A2(new_n3458_), .B(new_n10976_), .ZN(new_n10977_));
  OAI21_X1   g08541(.A1(new_n10977_), .A2(pi0075), .B(new_n6645_), .ZN(new_n10978_));
  OAI21_X1   g08542(.A1(new_n10978_), .A2(new_n10933_), .B(new_n10927_), .ZN(new_n10979_));
  AOI21_X1   g08543(.A1(new_n3041_), .A2(new_n5422_), .B(new_n5423_), .ZN(new_n10980_));
  NOR2_X1    g08544(.A1(new_n10980_), .A2(new_n6762_), .ZN(new_n10981_));
  AOI21_X1   g08545(.A1(new_n6750_), .A2(new_n10981_), .B(new_n2628_), .ZN(new_n10982_));
  OAI21_X1   g08546(.A1(pi1093), .A2(new_n5445_), .B(new_n5451_), .ZN(new_n10983_));
  NAND3_X1   g08547(.A1(new_n6750_), .A2(new_n6744_), .A3(new_n10983_), .ZN(new_n10984_));
  AOI21_X1   g08548(.A1(new_n2628_), .A2(new_n10984_), .B(new_n10982_), .ZN(new_n10985_));
  OAI21_X1   g08549(.A1(new_n10985_), .A2(new_n10911_), .B(pi0039), .ZN(new_n10986_));
  NOR2_X1    g08550(.A1(new_n10959_), .A2(new_n10960_), .ZN(new_n10987_));
  NAND2_X1   g08551(.A1(new_n10987_), .A2(new_n10964_), .ZN(new_n10988_));
  NAND3_X1   g08552(.A1(new_n10988_), .A2(new_n3265_), .A3(new_n10986_), .ZN(new_n10989_));
  NAND2_X1   g08553(.A1(new_n10912_), .A2(pi0038), .ZN(new_n10990_));
  AOI21_X1   g08554(.A1(new_n10989_), .A2(new_n10990_), .B(pi0100), .ZN(new_n10991_));
  INV_X1     g08555(.I(new_n10934_), .ZN(new_n10992_));
  OAI21_X1   g08556(.A1(new_n10935_), .A2(pi0120), .B(new_n10992_), .ZN(new_n10993_));
  NAND2_X1   g08557(.A1(new_n10912_), .A2(pi0100), .ZN(new_n10994_));
  AOI21_X1   g08558(.A1(new_n10993_), .A2(new_n6820_), .B(new_n10994_), .ZN(new_n10995_));
  OAI21_X1   g08559(.A1(new_n10991_), .A2(new_n10995_), .B(new_n3458_), .ZN(new_n10996_));
  AOI21_X1   g08560(.A1(new_n10996_), .A2(new_n10975_), .B(pi0075), .ZN(new_n10997_));
  OAI21_X1   g08561(.A1(new_n6869_), .A2(new_n10911_), .B(new_n6645_), .ZN(new_n10998_));
  NOR2_X1    g08562(.A1(new_n10926_), .A2(new_n6350_), .ZN(new_n10999_));
  OAI21_X1   g08563(.A1(new_n10997_), .A2(new_n10998_), .B(new_n10999_), .ZN(new_n11000_));
  AOI21_X1   g08564(.A1(new_n10979_), .A2(new_n11000_), .B(new_n10901_), .ZN(new_n11001_));
  OAI21_X1   g08565(.A1(new_n11001_), .A2(po1038), .B(new_n10923_), .ZN(new_n11002_));
  AOI21_X1   g08566(.A1(new_n6648_), .A2(new_n10917_), .B(new_n10919_), .ZN(new_n11003_));
  INV_X1     g08567(.I(new_n10927_), .ZN(new_n11004_));
  NOR2_X1    g08568(.A1(new_n3081_), .A2(new_n10915_), .ZN(new_n11005_));
  NAND3_X1   g08569(.A1(new_n2549_), .A2(new_n2771_), .A3(new_n6714_), .ZN(new_n11006_));
  NOR4_X1    g08570(.A1(new_n2536_), .A2(new_n3047_), .A3(new_n7279_), .A4(new_n11006_), .ZN(new_n11007_));
  NAND4_X1   g08571(.A1(new_n2738_), .A2(pi0252), .A3(new_n2746_), .A4(new_n11007_), .ZN(new_n11008_));
  OAI21_X1   g08572(.A1(new_n11008_), .A2(new_n6705_), .B(new_n11005_), .ZN(new_n11009_));
  INV_X1     g08573(.I(new_n10916_), .ZN(new_n11010_));
  NOR2_X1    g08574(.A1(new_n11010_), .A2(pi1091), .ZN(new_n11011_));
  NOR2_X1    g08575(.A1(new_n11011_), .A2(pi0120), .ZN(new_n11012_));
  AOI22_X1   g08576(.A1(new_n6798_), .A2(pi0120), .B1(new_n11009_), .B2(new_n11012_), .ZN(new_n11013_));
  NAND2_X1   g08577(.A1(new_n11013_), .A2(new_n8224_), .ZN(new_n11014_));
  OAI21_X1   g08578(.A1(new_n8224_), .A2(new_n10917_), .B(new_n11014_), .ZN(new_n11015_));
  NAND2_X1   g08579(.A1(new_n11015_), .A2(new_n2658_), .ZN(new_n11016_));
  INV_X1     g08580(.I(new_n10917_), .ZN(new_n11017_));
  AOI21_X1   g08581(.A1(new_n2659_), .A2(new_n11017_), .B(new_n3465_), .ZN(new_n11018_));
  OAI21_X1   g08582(.A1(new_n11017_), .A2(new_n3272_), .B(pi0087), .ZN(new_n11019_));
  AOI21_X1   g08583(.A1(new_n6874_), .A2(pi0120), .B(new_n3273_), .ZN(new_n11020_));
  INV_X1     g08584(.I(new_n11005_), .ZN(new_n11021_));
  NOR3_X1    g08585(.A1(new_n3024_), .A2(new_n3045_), .A3(new_n5329_), .ZN(new_n11022_));
  AOI21_X1   g08586(.A1(new_n2531_), .A2(new_n11022_), .B(new_n11021_), .ZN(new_n11023_));
  INV_X1     g08587(.I(new_n11011_), .ZN(new_n11024_));
  AOI21_X1   g08588(.A1(new_n2531_), .A2(new_n9893_), .B(new_n11024_), .ZN(new_n11025_));
  OAI21_X1   g08589(.A1(new_n11023_), .A2(new_n11025_), .B(new_n10903_), .ZN(new_n11026_));
  AOI21_X1   g08590(.A1(new_n11020_), .A2(new_n11026_), .B(new_n11019_), .ZN(new_n11027_));
  NOR4_X1    g08591(.A1(new_n6705_), .A2(new_n3045_), .A3(new_n2530_), .A4(new_n6654_), .ZN(new_n11028_));
  OAI21_X1   g08592(.A1(new_n11028_), .A2(new_n11021_), .B(new_n11012_), .ZN(new_n11029_));
  AOI21_X1   g08593(.A1(new_n10992_), .A2(new_n11029_), .B(new_n6819_), .ZN(new_n11030_));
  AOI21_X1   g08594(.A1(new_n11030_), .A2(new_n2627_), .B(new_n2702_), .ZN(new_n11031_));
  OAI22_X1   g08595(.A1(new_n11031_), .A2(pi0038), .B1(new_n6820_), .B2(new_n11017_), .ZN(new_n11032_));
  AOI21_X1   g08596(.A1(new_n6756_), .A2(new_n11017_), .B(new_n5446_), .ZN(new_n11033_));
  AOI21_X1   g08597(.A1(new_n6753_), .A2(new_n11017_), .B(new_n5445_), .ZN(new_n11034_));
  OAI21_X1   g08598(.A1(new_n11033_), .A2(new_n11034_), .B(new_n6744_), .ZN(new_n11035_));
  AOI21_X1   g08599(.A1(new_n6759_), .A2(new_n10917_), .B(pi0299), .ZN(new_n11036_));
  AOI21_X1   g08600(.A1(new_n6762_), .A2(new_n10917_), .B(new_n2628_), .ZN(new_n11037_));
  AOI21_X1   g08601(.A1(new_n6756_), .A2(new_n11017_), .B(new_n5422_), .ZN(new_n11038_));
  AOI21_X1   g08602(.A1(new_n6753_), .A2(new_n11017_), .B(new_n6764_), .ZN(new_n11039_));
  OAI21_X1   g08603(.A1(new_n11038_), .A2(new_n11039_), .B(new_n6761_), .ZN(new_n11040_));
  AOI22_X1   g08604(.A1(new_n11035_), .A2(new_n11036_), .B1(new_n11040_), .B2(new_n11037_), .ZN(new_n11041_));
  NOR2_X1    g08605(.A1(new_n11041_), .A2(new_n2627_), .ZN(new_n11042_));
  INV_X1     g08606(.I(new_n10915_), .ZN(new_n11043_));
  INV_X1     g08607(.I(new_n6666_), .ZN(new_n11044_));
  NOR4_X1    g08608(.A1(new_n2870_), .A2(pi0088), .A3(new_n2887_), .A4(new_n2858_), .ZN(new_n11045_));
  AND4_X2    g08609(.A1(new_n2985_), .A2(new_n6665_), .A3(new_n2786_), .A4(new_n11045_), .Z(new_n11046_));
  OAI21_X1   g08610(.A1(new_n11044_), .A2(new_n11046_), .B(pi0950), .ZN(new_n11047_));
  NOR2_X1    g08611(.A1(new_n11047_), .A2(new_n6716_), .ZN(new_n11048_));
  NAND3_X1   g08612(.A1(new_n11043_), .A2(pi0122), .A3(pi0829), .ZN(new_n11049_));
  NAND2_X1   g08613(.A1(new_n11048_), .A2(pi0824), .ZN(new_n11050_));
  NAND2_X1   g08614(.A1(new_n11050_), .A2(new_n11043_), .ZN(new_n11051_));
  OAI22_X1   g08615(.A1(new_n11051_), .A2(pi0829), .B1(new_n11048_), .B2(new_n11049_), .ZN(new_n11052_));
  NOR3_X1    g08616(.A1(new_n8467_), .A2(pi0072), .A3(new_n3045_), .ZN(new_n11053_));
  NOR2_X1    g08617(.A1(new_n11045_), .A2(pi0097), .ZN(new_n11054_));
  NOR3_X1    g08618(.A1(new_n3032_), .A2(new_n11054_), .A3(new_n3030_), .ZN(new_n11055_));
  OAI21_X1   g08619(.A1(new_n11055_), .A2(new_n6719_), .B(new_n2520_), .ZN(new_n11056_));
  NAND2_X1   g08620(.A1(new_n11056_), .A2(new_n6663_), .ZN(new_n11057_));
  AOI21_X1   g08621(.A1(new_n11057_), .A2(new_n6665_), .B(pi0051), .ZN(new_n11058_));
  OAI21_X1   g08622(.A1(new_n11058_), .A2(new_n2832_), .B(new_n2742_), .ZN(new_n11059_));
  AOI21_X1   g08623(.A1(new_n11059_), .A2(new_n11053_), .B(new_n6654_), .ZN(new_n11060_));
  AOI21_X1   g08624(.A1(new_n11043_), .A2(new_n11060_), .B(new_n11052_), .ZN(new_n11061_));
  OAI22_X1   g08625(.A1(new_n11061_), .A2(new_n6713_), .B1(new_n5532_), .B2(new_n11010_), .ZN(new_n11062_));
  NAND2_X1   g08626(.A1(new_n11062_), .A2(pi1091), .ZN(new_n11063_));
  AOI21_X1   g08627(.A1(new_n11050_), .A2(new_n11011_), .B(pi0120), .ZN(new_n11064_));
  NOR3_X1    g08628(.A1(new_n10959_), .A2(new_n10960_), .A3(new_n10963_), .ZN(new_n11065_));
  AOI22_X1   g08629(.A1(new_n11065_), .A2(pi0120), .B1(new_n11063_), .B2(new_n11064_), .ZN(new_n11066_));
  AOI21_X1   g08630(.A1(new_n11066_), .A2(new_n2627_), .B(new_n11042_), .ZN(new_n11067_));
  OAI21_X1   g08631(.A1(new_n11067_), .A2(new_n3271_), .B(new_n11032_), .ZN(new_n11068_));
  AOI21_X1   g08632(.A1(new_n11068_), .A2(new_n3458_), .B(new_n11027_), .ZN(new_n11069_));
  AOI22_X1   g08633(.A1(new_n11069_), .A2(new_n3465_), .B1(new_n11016_), .B2(new_n11018_), .ZN(new_n11070_));
  NOR2_X1    g08634(.A1(new_n11070_), .A2(new_n6648_), .ZN(new_n11071_));
  NOR2_X1    g08635(.A1(new_n10908_), .A2(new_n10917_), .ZN(new_n11072_));
  NOR2_X1    g08636(.A1(new_n11072_), .A2(new_n6700_), .ZN(new_n11073_));
  NOR2_X1    g08637(.A1(new_n11024_), .A2(new_n9821_), .ZN(new_n11074_));
  INV_X1     g08638(.I(new_n11074_), .ZN(new_n11075_));
  AOI21_X1   g08639(.A1(new_n11009_), .A2(new_n11075_), .B(pi0120), .ZN(new_n11076_));
  NOR3_X1    g08640(.A1(new_n10930_), .A2(new_n2659_), .A3(new_n11076_), .ZN(new_n11077_));
  NOR3_X1    g08641(.A1(new_n11077_), .A2(new_n3465_), .A3(new_n11073_), .ZN(new_n11078_));
  AOI21_X1   g08642(.A1(new_n10093_), .A2(new_n3273_), .B(new_n11019_), .ZN(new_n11079_));
  INV_X1     g08643(.I(new_n10972_), .ZN(new_n11080_));
  NOR2_X1    g08644(.A1(new_n11023_), .A2(new_n11074_), .ZN(new_n11081_));
  OAI22_X1   g08645(.A1(new_n11020_), .A2(new_n11080_), .B1(new_n11026_), .B2(new_n11081_), .ZN(new_n11082_));
  NAND2_X1   g08646(.A1(new_n11082_), .A2(new_n11079_), .ZN(new_n11083_));
  INV_X1     g08647(.I(new_n11072_), .ZN(new_n11084_));
  NAND2_X1   g08648(.A1(new_n11084_), .A2(new_n6819_), .ZN(new_n11085_));
  INV_X1     g08649(.I(new_n10904_), .ZN(new_n11086_));
  NOR2_X1    g08650(.A1(new_n11028_), .A2(new_n11021_), .ZN(new_n11087_));
  NOR2_X1    g08651(.A1(new_n11087_), .A2(new_n11074_), .ZN(new_n11088_));
  OAI22_X1   g08652(.A1(new_n11088_), .A2(pi0120), .B1(new_n6777_), .B2(new_n11086_), .ZN(new_n11089_));
  OAI21_X1   g08653(.A1(new_n11089_), .A2(new_n6819_), .B(new_n11085_), .ZN(new_n11090_));
  OAI21_X1   g08654(.A1(new_n11072_), .A2(new_n2572_), .B(pi0100), .ZN(new_n11091_));
  AOI21_X1   g08655(.A1(new_n11090_), .A2(new_n2572_), .B(new_n11091_), .ZN(new_n11092_));
  NAND2_X1   g08656(.A1(new_n11072_), .A2(pi0038), .ZN(new_n11093_));
  NOR2_X1    g08657(.A1(new_n11072_), .A2(new_n5449_), .ZN(new_n11094_));
  OAI21_X1   g08658(.A1(new_n6748_), .A2(new_n11021_), .B(new_n11075_), .ZN(new_n11095_));
  AOI22_X1   g08659(.A1(new_n6751_), .A2(new_n10904_), .B1(new_n10903_), .B2(new_n11095_), .ZN(new_n11096_));
  AOI21_X1   g08660(.A1(new_n11096_), .A2(new_n5449_), .B(new_n11094_), .ZN(new_n11097_));
  NOR2_X1    g08661(.A1(new_n11097_), .A2(new_n5445_), .ZN(new_n11098_));
  NOR2_X1    g08662(.A1(new_n11072_), .A2(new_n5427_), .ZN(new_n11099_));
  AOI21_X1   g08663(.A1(new_n11096_), .A2(new_n5427_), .B(new_n11099_), .ZN(new_n11100_));
  NOR2_X1    g08664(.A1(new_n11100_), .A2(new_n5446_), .ZN(new_n11101_));
  OAI21_X1   g08665(.A1(new_n11098_), .A2(new_n11101_), .B(new_n6744_), .ZN(new_n11102_));
  AOI21_X1   g08666(.A1(new_n11084_), .A2(new_n6759_), .B(pi0299), .ZN(new_n11103_));
  NAND2_X1   g08667(.A1(new_n11102_), .A2(new_n11103_), .ZN(new_n11104_));
  NOR2_X1    g08668(.A1(new_n11097_), .A2(new_n6764_), .ZN(new_n11105_));
  NOR2_X1    g08669(.A1(new_n11100_), .A2(new_n5422_), .ZN(new_n11106_));
  OAI21_X1   g08670(.A1(new_n11105_), .A2(new_n11106_), .B(new_n6761_), .ZN(new_n11107_));
  NAND2_X1   g08671(.A1(new_n10093_), .A2(new_n6762_), .ZN(new_n11108_));
  NAND3_X1   g08672(.A1(new_n11107_), .A2(new_n11037_), .A3(new_n11108_), .ZN(new_n11109_));
  NAND3_X1   g08673(.A1(new_n11109_), .A2(new_n11104_), .A3(pi0039), .ZN(new_n11110_));
  NAND2_X1   g08674(.A1(new_n10961_), .A2(new_n10962_), .ZN(new_n11111_));
  NOR2_X1    g08675(.A1(new_n11111_), .A2(new_n10903_), .ZN(new_n11112_));
  NAND4_X1   g08676(.A1(new_n11050_), .A2(new_n6870_), .A3(new_n9822_), .A4(new_n11043_), .ZN(new_n11113_));
  AND3_X2    g08677(.A1(new_n11063_), .A2(new_n10903_), .A3(new_n11113_), .Z(new_n11114_));
  OAI21_X1   g08678(.A1(new_n11112_), .A2(new_n11114_), .B(new_n2627_), .ZN(new_n11115_));
  NAND3_X1   g08679(.A1(new_n11115_), .A2(new_n3265_), .A3(new_n11110_), .ZN(new_n11116_));
  AOI21_X1   g08680(.A1(new_n11116_), .A2(new_n11093_), .B(pi0100), .ZN(new_n11117_));
  OAI21_X1   g08681(.A1(new_n11117_), .A2(new_n11092_), .B(new_n3458_), .ZN(new_n11118_));
  AOI21_X1   g08682(.A1(new_n11118_), .A2(new_n11083_), .B(pi0075), .ZN(new_n11119_));
  NOR3_X1    g08683(.A1(new_n11119_), .A2(new_n6648_), .A3(new_n11078_), .ZN(new_n11120_));
  OAI22_X1   g08684(.A1(new_n11120_), .A2(new_n11004_), .B1(new_n6350_), .B2(new_n11071_), .ZN(new_n11121_));
  OAI21_X1   g08685(.A1(new_n11065_), .A2(pi0039), .B(new_n6876_), .ZN(new_n11122_));
  AOI21_X1   g08686(.A1(new_n11122_), .A2(new_n2702_), .B(new_n6821_), .ZN(new_n11123_));
  OAI21_X1   g08687(.A1(new_n11123_), .A2(pi0087), .B(new_n6875_), .ZN(new_n11124_));
  AOI21_X1   g08688(.A1(new_n11124_), .A2(new_n3465_), .B(new_n6799_), .ZN(new_n11125_));
  OAI21_X1   g08689(.A1(pi0120), .A2(new_n6645_), .B(new_n6349_), .ZN(new_n11126_));
  OAI22_X1   g08690(.A1(new_n11125_), .A2(new_n11126_), .B1(new_n6645_), .B2(new_n10910_), .ZN(new_n11127_));
  OR2_X2     g08691(.A1(new_n10929_), .A2(new_n6701_), .Z(new_n11128_));
  INV_X1     g08692(.I(new_n10093_), .ZN(new_n11129_));
  NAND2_X1   g08693(.A1(new_n6701_), .A2(new_n11129_), .ZN(new_n11130_));
  AOI21_X1   g08694(.A1(new_n11128_), .A2(new_n11130_), .B(new_n3465_), .ZN(new_n11131_));
  NOR2_X1    g08695(.A1(new_n6752_), .A2(new_n10093_), .ZN(new_n11132_));
  INV_X1     g08696(.I(new_n11132_), .ZN(new_n11133_));
  NAND2_X1   g08697(.A1(new_n11133_), .A2(new_n5446_), .ZN(new_n11134_));
  NOR2_X1    g08698(.A1(new_n6755_), .A2(new_n10093_), .ZN(new_n11135_));
  OAI21_X1   g08699(.A1(new_n5446_), .A2(new_n11135_), .B(new_n11134_), .ZN(new_n11136_));
  OAI21_X1   g08700(.A1(new_n11129_), .A2(new_n6744_), .B(new_n2628_), .ZN(new_n11137_));
  AOI21_X1   g08701(.A1(new_n11136_), .A2(new_n6744_), .B(new_n11137_), .ZN(new_n11138_));
  NAND2_X1   g08702(.A1(new_n11133_), .A2(new_n5422_), .ZN(new_n11139_));
  OAI21_X1   g08703(.A1(new_n5422_), .A2(new_n11135_), .B(new_n11139_), .ZN(new_n11140_));
  NAND2_X1   g08704(.A1(new_n11108_), .A2(pi0299), .ZN(new_n11141_));
  AOI21_X1   g08705(.A1(new_n11140_), .A2(new_n6761_), .B(new_n11141_), .ZN(new_n11142_));
  NOR3_X1    g08706(.A1(new_n11138_), .A2(new_n11142_), .A3(new_n2627_), .ZN(new_n11143_));
  NOR2_X1    g08707(.A1(new_n11111_), .A2(pi0039), .ZN(new_n11144_));
  OAI21_X1   g08708(.A1(new_n11144_), .A2(new_n11143_), .B(new_n3265_), .ZN(new_n11145_));
  AOI21_X1   g08709(.A1(new_n10093_), .A2(pi0038), .B(pi0100), .ZN(new_n11146_));
  AOI22_X1   g08710(.A1(new_n11145_), .A2(new_n11146_), .B1(new_n6821_), .B2(new_n11129_), .ZN(new_n11147_));
  OAI21_X1   g08711(.A1(new_n11147_), .A2(pi0087), .B(new_n10974_), .ZN(new_n11148_));
  AOI21_X1   g08712(.A1(new_n11148_), .A2(new_n3465_), .B(new_n11131_), .ZN(new_n11149_));
  NOR2_X1    g08713(.A1(new_n11149_), .A2(new_n10925_), .ZN(new_n11150_));
  OAI21_X1   g08714(.A1(new_n11150_), .A2(new_n11127_), .B(pi0120), .ZN(new_n11151_));
  NOR2_X1    g08715(.A1(new_n11151_), .A2(new_n10922_), .ZN(new_n11152_));
  AOI21_X1   g08716(.A1(new_n11121_), .A2(new_n11003_), .B(new_n11152_), .ZN(new_n11153_));
  OAI21_X1   g08717(.A1(new_n11153_), .A2(new_n10902_), .B(new_n11002_), .ZN(po0278));
  INV_X1     g08718(.I(new_n9393_), .ZN(new_n11155_));
  NOR2_X1    g08719(.A1(new_n11155_), .A2(new_n3458_), .ZN(new_n11156_));
  NOR2_X1    g08720(.A1(new_n5437_), .A2(new_n2744_), .ZN(new_n11157_));
  INV_X1     g08721(.I(new_n11157_), .ZN(new_n11158_));
  NOR2_X1    g08722(.A1(new_n11158_), .A2(pi0146), .ZN(new_n11159_));
  NOR2_X1    g08723(.A1(new_n11159_), .A2(new_n3360_), .ZN(new_n11160_));
  NOR3_X1    g08724(.A1(new_n2488_), .A2(pi0067), .A3(pi0071), .ZN(new_n11161_));
  INV_X1     g08725(.I(new_n11161_), .ZN(new_n11162_));
  NOR2_X1    g08726(.A1(new_n11162_), .A2(pi0051), .ZN(new_n11163_));
  NOR2_X1    g08727(.A1(new_n11163_), .A2(new_n5437_), .ZN(new_n11164_));
  INV_X1     g08728(.I(new_n11164_), .ZN(new_n11165_));
  NOR2_X1    g08729(.A1(new_n2744_), .A2(new_n3107_), .ZN(new_n11166_));
  NOR3_X1    g08730(.A1(new_n11165_), .A2(new_n11160_), .A3(new_n11166_), .ZN(new_n11167_));
  INV_X1     g08731(.I(new_n11167_), .ZN(new_n11168_));
  NOR2_X1    g08732(.A1(new_n11168_), .A2(pi0087), .ZN(new_n11169_));
  OAI21_X1   g08733(.A1(new_n11169_), .A2(new_n11156_), .B(pi0232), .ZN(new_n11170_));
  INV_X1     g08734(.I(new_n11163_), .ZN(new_n11171_));
  NOR2_X1    g08735(.A1(new_n11171_), .A2(pi0087), .ZN(new_n11172_));
  INV_X1     g08736(.I(pi0130), .ZN(new_n11173_));
  INV_X1     g08737(.I(pi0132), .ZN(new_n11174_));
  INV_X1     g08738(.I(pi0136), .ZN(new_n11175_));
  NOR2_X1    g08739(.A1(pi0134), .A2(pi0135), .ZN(new_n11176_));
  NAND4_X1   g08740(.A1(new_n11176_), .A2(new_n11173_), .A3(new_n11174_), .A4(new_n11175_), .ZN(new_n11177_));
  NOR3_X1    g08741(.A1(new_n11177_), .A2(pi0121), .A3(pi0126), .ZN(new_n11178_));
  INV_X1     g08742(.I(new_n11178_), .ZN(new_n11179_));
  NOR2_X1    g08743(.A1(pi0125), .A2(pi0133), .ZN(new_n11180_));
  OR2_X2     g08744(.A1(new_n11180_), .A2(pi0121), .Z(new_n11181_));
  NAND2_X1   g08745(.A1(new_n11180_), .A2(pi0121), .ZN(new_n11182_));
  NAND3_X1   g08746(.A1(new_n11179_), .A2(new_n11181_), .A3(new_n11182_), .ZN(new_n11183_));
  AOI21_X1   g08747(.A1(new_n11172_), .A2(new_n11183_), .B(new_n6643_), .ZN(new_n11184_));
  NAND2_X1   g08748(.A1(new_n11170_), .A2(new_n11184_), .ZN(new_n11185_));
  NOR2_X1    g08749(.A1(new_n9517_), .A2(pi0299), .ZN(new_n11186_));
  AOI21_X1   g08750(.A1(pi0163), .A2(pi0299), .B(new_n11186_), .ZN(new_n11187_));
  OAI21_X1   g08751(.A1(new_n6698_), .A2(new_n11187_), .B(pi0087), .ZN(new_n11188_));
  NAND2_X1   g08752(.A1(new_n11168_), .A2(pi0299), .ZN(new_n11189_));
  NOR2_X1    g08753(.A1(new_n11158_), .A2(pi0142), .ZN(new_n11190_));
  NOR2_X1    g08754(.A1(new_n11190_), .A2(new_n8058_), .ZN(new_n11191_));
  NOR2_X1    g08755(.A1(new_n2744_), .A2(new_n2724_), .ZN(new_n11192_));
  NOR2_X1    g08756(.A1(new_n11165_), .A2(new_n11192_), .ZN(new_n11193_));
  INV_X1     g08757(.I(new_n11193_), .ZN(new_n11194_));
  NOR2_X1    g08758(.A1(new_n11194_), .A2(new_n11191_), .ZN(new_n11195_));
  INV_X1     g08759(.I(new_n11195_), .ZN(new_n11196_));
  NAND2_X1   g08760(.A1(new_n11196_), .A2(new_n2628_), .ZN(new_n11197_));
  NAND3_X1   g08761(.A1(new_n11197_), .A2(pi0232), .A3(new_n11189_), .ZN(new_n11198_));
  NOR2_X1    g08762(.A1(new_n2607_), .A2(pi0087), .ZN(new_n11199_));
  AOI21_X1   g08763(.A1(new_n11198_), .A2(new_n11199_), .B(new_n11183_), .ZN(new_n11200_));
  NAND2_X1   g08764(.A1(new_n11200_), .A2(new_n11188_), .ZN(new_n11201_));
  NOR2_X1    g08765(.A1(new_n11198_), .A2(new_n2702_), .ZN(new_n11202_));
  AND2_X2    g08766(.A1(new_n11198_), .A2(pi0038), .Z(new_n11203_));
  NOR2_X1    g08767(.A1(new_n11203_), .A2(pi0100), .ZN(new_n11204_));
  INV_X1     g08768(.I(new_n11160_), .ZN(new_n11205_));
  NOR2_X1    g08769(.A1(new_n5437_), .A2(pi0051), .ZN(new_n11206_));
  INV_X1     g08770(.I(new_n11206_), .ZN(new_n11207_));
  NAND3_X1   g08771(.A1(new_n8247_), .A2(new_n2474_), .A3(new_n10280_), .ZN(new_n11208_));
  INV_X1     g08772(.I(new_n11208_), .ZN(new_n11209_));
  NAND4_X1   g08773(.A1(new_n11209_), .A2(new_n7275_), .A3(pi0077), .A4(new_n2515_), .ZN(new_n11210_));
  NOR2_X1    g08774(.A1(new_n6677_), .A2(new_n3007_), .ZN(new_n11211_));
  INV_X1     g08775(.I(new_n11211_), .ZN(new_n11212_));
  NOR3_X1    g08776(.A1(new_n11212_), .A2(pi0024), .A3(new_n5590_), .ZN(new_n11213_));
  INV_X1     g08777(.I(new_n11213_), .ZN(new_n11214_));
  NOR3_X1    g08778(.A1(new_n11210_), .A2(new_n7293_), .A3(new_n11214_), .ZN(new_n11215_));
  INV_X1     g08779(.I(new_n11215_), .ZN(new_n11216_));
  NOR2_X1    g08780(.A1(new_n11216_), .A2(new_n2526_), .ZN(new_n11217_));
  INV_X1     g08781(.I(new_n11217_), .ZN(new_n11218_));
  AOI21_X1   g08782(.A1(new_n11218_), .A2(new_n11161_), .B(new_n11207_), .ZN(new_n11219_));
  NOR2_X1    g08783(.A1(new_n11219_), .A2(new_n3107_), .ZN(new_n11220_));
  NOR2_X1    g08784(.A1(new_n11217_), .A2(new_n11171_), .ZN(new_n11221_));
  NOR2_X1    g08785(.A1(new_n11221_), .A2(new_n5437_), .ZN(new_n11222_));
  INV_X1     g08786(.I(new_n11222_), .ZN(new_n11223_));
  AOI21_X1   g08787(.A1(new_n3107_), .A2(new_n11223_), .B(new_n11220_), .ZN(new_n11224_));
  NAND4_X1   g08788(.A1(new_n2882_), .A2(new_n2744_), .A3(new_n9226_), .A4(new_n11213_), .ZN(new_n11225_));
  NOR2_X1    g08789(.A1(new_n2526_), .A2(new_n5437_), .ZN(new_n11226_));
  INV_X1     g08790(.I(new_n11226_), .ZN(new_n11227_));
  NOR2_X1    g08791(.A1(new_n11225_), .A2(new_n11227_), .ZN(new_n11228_));
  OAI22_X1   g08792(.A1(new_n11224_), .A2(pi0161), .B1(new_n11205_), .B2(new_n11228_), .ZN(new_n11229_));
  OAI21_X1   g08793(.A1(new_n11189_), .A2(pi0158), .B(pi0232), .ZN(new_n11230_));
  AOI21_X1   g08794(.A1(new_n11229_), .A2(new_n7731_), .B(new_n11230_), .ZN(new_n11231_));
  NAND2_X1   g08795(.A1(new_n2572_), .A2(new_n9471_), .ZN(new_n11232_));
  OAI21_X1   g08796(.A1(new_n11231_), .A2(new_n11232_), .B(new_n11204_), .ZN(new_n11233_));
  NOR2_X1    g08797(.A1(new_n11161_), .A2(pi0051), .ZN(new_n11234_));
  INV_X1     g08798(.I(new_n11234_), .ZN(new_n11235_));
  NOR2_X1    g08799(.A1(new_n11235_), .A2(new_n8282_), .ZN(new_n11236_));
  NOR2_X1    g08800(.A1(new_n11208_), .A2(new_n2856_), .ZN(new_n11237_));
  NAND3_X1   g08801(.A1(new_n11237_), .A2(new_n9100_), .A3(new_n11211_), .ZN(new_n11238_));
  NOR2_X1    g08802(.A1(new_n11238_), .A2(new_n2526_), .ZN(new_n11239_));
  NOR2_X1    g08803(.A1(new_n11239_), .A2(new_n11171_), .ZN(new_n11240_));
  NOR2_X1    g08804(.A1(new_n11240_), .A2(pi0051), .ZN(new_n11241_));
  AOI21_X1   g08805(.A1(new_n11241_), .A2(new_n8282_), .B(new_n11236_), .ZN(new_n11242_));
  NOR2_X1    g08806(.A1(new_n11242_), .A2(new_n5437_), .ZN(new_n11243_));
  NOR3_X1    g08807(.A1(new_n11243_), .A2(pi0161), .A3(new_n11159_), .ZN(new_n11244_));
  NOR2_X1    g08808(.A1(new_n8283_), .A2(new_n5437_), .ZN(new_n11245_));
  OAI21_X1   g08809(.A1(new_n11245_), .A2(new_n11205_), .B(new_n7508_), .ZN(new_n11246_));
  AOI21_X1   g08810(.A1(new_n11167_), .A2(new_n8070_), .B(new_n7981_), .ZN(new_n11247_));
  OAI21_X1   g08811(.A1(new_n11244_), .A2(new_n11246_), .B(new_n11247_), .ZN(new_n11248_));
  NAND2_X1   g08812(.A1(new_n11243_), .A2(new_n7519_), .ZN(new_n11249_));
  NAND3_X1   g08813(.A1(new_n11249_), .A2(new_n8058_), .A3(new_n11194_), .ZN(new_n11250_));
  NOR2_X1    g08814(.A1(new_n5437_), .A2(pi0287), .ZN(new_n11251_));
  INV_X1     g08815(.I(new_n11251_), .ZN(new_n11252_));
  NOR2_X1    g08816(.A1(new_n7525_), .A2(new_n11252_), .ZN(new_n11253_));
  NOR2_X1    g08817(.A1(new_n2530_), .A2(new_n2724_), .ZN(new_n11254_));
  NAND2_X1   g08818(.A1(new_n2831_), .A2(new_n6684_), .ZN(new_n11255_));
  NOR2_X1    g08819(.A1(new_n11255_), .A2(pi0142), .ZN(new_n11256_));
  OAI21_X1   g08820(.A1(new_n11256_), .A2(new_n11254_), .B(new_n11253_), .ZN(new_n11257_));
  AOI21_X1   g08821(.A1(new_n11257_), .A2(new_n11191_), .B(new_n5658_), .ZN(new_n11258_));
  NAND2_X1   g08822(.A1(new_n11250_), .A2(new_n11258_), .ZN(new_n11259_));
  AOI21_X1   g08823(.A1(new_n11195_), .A2(new_n5658_), .B(pi0299), .ZN(new_n11260_));
  OAI21_X1   g08824(.A1(new_n11189_), .A2(pi0159), .B(new_n7506_), .ZN(new_n11261_));
  AOI21_X1   g08825(.A1(new_n11259_), .A2(new_n11260_), .B(new_n11261_), .ZN(new_n11262_));
  AOI21_X1   g08826(.A1(new_n11262_), .A2(new_n11248_), .B(pi0038), .ZN(new_n11263_));
  INV_X1     g08827(.I(new_n11219_), .ZN(new_n11264_));
  NAND2_X1   g08828(.A1(new_n11264_), .A2(pi0142), .ZN(new_n11265_));
  NAND2_X1   g08829(.A1(new_n11223_), .A2(new_n2724_), .ZN(new_n11266_));
  AOI21_X1   g08830(.A1(new_n11266_), .A2(new_n11265_), .B(pi0144), .ZN(new_n11267_));
  INV_X1     g08831(.I(new_n11191_), .ZN(new_n11268_));
  OAI21_X1   g08832(.A1(new_n11228_), .A2(new_n11268_), .B(pi0180), .ZN(new_n11269_));
  OAI22_X1   g08833(.A1(new_n11267_), .A2(new_n11269_), .B1(pi0180), .B2(new_n11196_), .ZN(new_n11270_));
  NOR2_X1    g08834(.A1(new_n11270_), .A2(pi0179), .ZN(new_n11271_));
  INV_X1     g08835(.I(new_n11237_), .ZN(new_n11272_));
  OAI22_X1   g08836(.A1(new_n11210_), .A2(new_n7278_), .B1(new_n11272_), .B2(new_n2879_), .ZN(new_n11273_));
  NAND2_X1   g08837(.A1(new_n11273_), .A2(new_n7274_), .ZN(new_n11274_));
  AOI21_X1   g08838(.A1(new_n11212_), .A2(new_n11161_), .B(pi0051), .ZN(new_n11275_));
  INV_X1     g08839(.I(new_n11275_), .ZN(new_n11276_));
  AOI21_X1   g08840(.A1(new_n11274_), .A2(new_n11161_), .B(new_n11276_), .ZN(new_n11277_));
  NAND2_X1   g08841(.A1(new_n11277_), .A2(new_n9275_), .ZN(new_n11278_));
  INV_X1     g08842(.I(new_n11278_), .ZN(new_n11279_));
  NOR2_X1    g08843(.A1(new_n11235_), .A2(new_n9275_), .ZN(new_n11280_));
  OAI21_X1   g08844(.A1(new_n11279_), .A2(new_n11280_), .B(new_n5398_), .ZN(new_n11281_));
  NOR2_X1    g08845(.A1(new_n11279_), .A2(new_n11171_), .ZN(new_n11282_));
  NOR2_X1    g08846(.A1(new_n11282_), .A2(new_n5437_), .ZN(new_n11283_));
  NAND2_X1   g08847(.A1(new_n11283_), .A2(new_n2724_), .ZN(new_n11284_));
  OAI21_X1   g08848(.A1(new_n2724_), .A2(new_n11281_), .B(new_n11284_), .ZN(new_n11285_));
  OAI21_X1   g08849(.A1(new_n11285_), .A2(pi0144), .B(new_n5657_), .ZN(new_n11286_));
  NAND2_X1   g08850(.A1(new_n9382_), .A2(pi0024), .ZN(new_n11287_));
  NAND2_X1   g08851(.A1(new_n9377_), .A2(new_n7278_), .ZN(new_n11288_));
  AOI21_X1   g08852(.A1(new_n11287_), .A2(new_n11288_), .B(new_n2749_), .ZN(new_n11289_));
  NAND2_X1   g08853(.A1(new_n11289_), .A2(new_n11226_), .ZN(new_n11290_));
  INV_X1     g08854(.I(new_n11290_), .ZN(new_n11291_));
  NOR2_X1    g08855(.A1(new_n11291_), .A2(new_n11268_), .ZN(new_n11292_));
  OAI21_X1   g08856(.A1(new_n11292_), .A2(new_n11286_), .B(pi0179), .ZN(new_n11293_));
  NOR2_X1    g08857(.A1(pi0024), .A2(pi0314), .ZN(new_n11294_));
  NOR3_X1    g08858(.A1(new_n9381_), .A2(new_n2737_), .A3(new_n11294_), .ZN(new_n11295_));
  AOI21_X1   g08859(.A1(new_n9377_), .A2(new_n11294_), .B(new_n11295_), .ZN(new_n11296_));
  NOR3_X1    g08860(.A1(new_n11296_), .A2(new_n6677_), .A3(new_n7332_), .ZN(new_n11297_));
  NOR2_X1    g08861(.A1(new_n11297_), .A2(pi0051), .ZN(new_n11298_));
  NOR2_X1    g08862(.A1(new_n11298_), .A2(new_n5437_), .ZN(new_n11299_));
  INV_X1     g08863(.I(new_n11299_), .ZN(new_n11300_));
  OAI21_X1   g08864(.A1(new_n11300_), .A2(new_n11192_), .B(pi0144), .ZN(new_n11301_));
  INV_X1     g08865(.I(new_n11221_), .ZN(new_n11302_));
  NOR2_X1    g08866(.A1(new_n11279_), .A2(new_n11302_), .ZN(new_n11303_));
  OAI21_X1   g08867(.A1(new_n11303_), .A2(new_n5437_), .B(new_n2724_), .ZN(new_n11304_));
  NAND4_X1   g08868(.A1(new_n11274_), .A2(new_n11161_), .A3(new_n11216_), .A4(new_n11211_), .ZN(new_n11305_));
  AND3_X2    g08869(.A1(new_n11305_), .A2(new_n9275_), .A3(new_n11275_), .Z(new_n11306_));
  OAI21_X1   g08870(.A1(new_n11306_), .A2(new_n11280_), .B(new_n5398_), .ZN(new_n11307_));
  INV_X1     g08871(.I(new_n11307_), .ZN(new_n11308_));
  OAI21_X1   g08872(.A1(new_n2724_), .A2(new_n11308_), .B(new_n11304_), .ZN(new_n11309_));
  AOI21_X1   g08873(.A1(new_n11309_), .A2(new_n8058_), .B(new_n5657_), .ZN(new_n11310_));
  AOI21_X1   g08874(.A1(new_n11301_), .A2(new_n11310_), .B(new_n11293_), .ZN(new_n11311_));
  OAI21_X1   g08875(.A1(new_n11311_), .A2(new_n11271_), .B(new_n2628_), .ZN(new_n11312_));
  INV_X1     g08876(.I(new_n7731_), .ZN(new_n11313_));
  INV_X1     g08877(.I(new_n11303_), .ZN(new_n11314_));
  AOI21_X1   g08878(.A1(new_n11314_), .A2(new_n5398_), .B(pi0146), .ZN(new_n11315_));
  NOR2_X1    g08879(.A1(new_n11308_), .A2(new_n3107_), .ZN(new_n11316_));
  OAI21_X1   g08880(.A1(new_n11316_), .A2(new_n11315_), .B(new_n3360_), .ZN(new_n11317_));
  OAI21_X1   g08881(.A1(new_n11300_), .A2(new_n11166_), .B(pi0161), .ZN(new_n11318_));
  AOI21_X1   g08882(.A1(new_n11318_), .A2(new_n11317_), .B(new_n11313_), .ZN(new_n11319_));
  NAND2_X1   g08883(.A1(new_n11283_), .A2(new_n3107_), .ZN(new_n11320_));
  OAI21_X1   g08884(.A1(new_n3107_), .A2(new_n11281_), .B(new_n11320_), .ZN(new_n11321_));
  OAI22_X1   g08885(.A1(new_n11291_), .A2(new_n11205_), .B1(pi0161), .B2(new_n11321_), .ZN(new_n11322_));
  NAND2_X1   g08886(.A1(new_n11322_), .A2(new_n7689_), .ZN(new_n11323_));
  NAND2_X1   g08887(.A1(new_n11323_), .A2(pi0232), .ZN(new_n11324_));
  OAI21_X1   g08888(.A1(new_n11319_), .A2(new_n11324_), .B(pi0156), .ZN(new_n11325_));
  NAND3_X1   g08889(.A1(new_n11312_), .A2(new_n11325_), .A3(new_n2627_), .ZN(new_n11326_));
  AOI21_X1   g08890(.A1(new_n11326_), .A2(new_n11263_), .B(new_n11233_), .ZN(new_n11327_));
  NOR3_X1    g08891(.A1(new_n11327_), .A2(new_n2569_), .A3(new_n11202_), .ZN(new_n11328_));
  OAI21_X1   g08892(.A1(new_n11328_), .A2(new_n11201_), .B(new_n6643_), .ZN(new_n11329_));
  INV_X1     g08893(.I(new_n11202_), .ZN(new_n11330_));
  NOR2_X1    g08894(.A1(new_n11171_), .A2(new_n2702_), .ZN(new_n11331_));
  NOR2_X1    g08895(.A1(new_n11331_), .A2(new_n2569_), .ZN(new_n11332_));
  INV_X1     g08896(.I(new_n11332_), .ZN(new_n11333_));
  AOI21_X1   g08897(.A1(new_n11203_), .A2(new_n11171_), .B(pi0100), .ZN(new_n11334_));
  INV_X1     g08898(.I(new_n6806_), .ZN(new_n11335_));
  INV_X1     g08899(.I(new_n11239_), .ZN(new_n11336_));
  AOI21_X1   g08900(.A1(new_n5756_), .A2(new_n11335_), .B(new_n11336_), .ZN(new_n11337_));
  NAND2_X1   g08901(.A1(new_n11163_), .A2(new_n5666_), .ZN(new_n11338_));
  OAI21_X1   g08902(.A1(new_n11337_), .A2(new_n11338_), .B(pi0039), .ZN(new_n11339_));
  OAI21_X1   g08903(.A1(new_n11167_), .A2(new_n11163_), .B(new_n5550_), .ZN(new_n11340_));
  INV_X1     g08904(.I(new_n11159_), .ZN(new_n11341_));
  INV_X1     g08905(.I(new_n11255_), .ZN(new_n11342_));
  NOR2_X1    g08906(.A1(new_n11342_), .A2(pi0051), .ZN(new_n11343_));
  INV_X1     g08907(.I(new_n11343_), .ZN(new_n11344_));
  NOR2_X1    g08908(.A1(new_n11344_), .A2(new_n5437_), .ZN(new_n11345_));
  INV_X1     g08909(.I(new_n11240_), .ZN(new_n11346_));
  NOR2_X1    g08910(.A1(new_n11346_), .A2(new_n5398_), .ZN(new_n11347_));
  NOR2_X1    g08911(.A1(new_n11347_), .A2(new_n11345_), .ZN(new_n11348_));
  INV_X1     g08912(.I(new_n11348_), .ZN(new_n11349_));
  NOR2_X1    g08913(.A1(new_n11252_), .A2(pi0051), .ZN(new_n11350_));
  NOR2_X1    g08914(.A1(new_n11349_), .A2(new_n11350_), .ZN(new_n11351_));
  INV_X1     g08915(.I(new_n11351_), .ZN(new_n11352_));
  AOI21_X1   g08916(.A1(new_n11239_), .A2(new_n11252_), .B(new_n11171_), .ZN(new_n11353_));
  INV_X1     g08917(.I(new_n11353_), .ZN(new_n11354_));
  NAND2_X1   g08918(.A1(new_n11354_), .A2(pi0161), .ZN(new_n11355_));
  OAI21_X1   g08919(.A1(new_n11352_), .A2(pi0161), .B(new_n11355_), .ZN(new_n11356_));
  NAND2_X1   g08920(.A1(new_n11356_), .A2(new_n11341_), .ZN(new_n11357_));
  OAI21_X1   g08921(.A1(new_n11240_), .A2(new_n11159_), .B(pi0161), .ZN(new_n11358_));
  NOR2_X1    g08922(.A1(new_n11348_), .A2(new_n3107_), .ZN(new_n11359_));
  AOI21_X1   g08923(.A1(new_n2587_), .A2(new_n5398_), .B(new_n11347_), .ZN(new_n11360_));
  NOR2_X1    g08924(.A1(new_n11360_), .A2(pi0146), .ZN(new_n11361_));
  OAI21_X1   g08925(.A1(new_n11361_), .A2(new_n11359_), .B(new_n3360_), .ZN(new_n11362_));
  AOI21_X1   g08926(.A1(new_n11362_), .A2(new_n11358_), .B(new_n5550_), .ZN(new_n11363_));
  OAI22_X1   g08927(.A1(new_n11357_), .A2(new_n2614_), .B1(new_n7508_), .B2(new_n11363_), .ZN(new_n11364_));
  NAND4_X1   g08928(.A1(new_n11364_), .A2(pi0159), .A3(pi0299), .A4(new_n11340_), .ZN(new_n11365_));
  OAI21_X1   g08929(.A1(new_n11163_), .A2(new_n11190_), .B(new_n5525_), .ZN(new_n11366_));
  INV_X1     g08930(.I(new_n11366_), .ZN(new_n11367_));
  NOR2_X1    g08931(.A1(new_n11240_), .A2(new_n11157_), .ZN(new_n11368_));
  NOR3_X1    g08932(.A1(new_n11368_), .A2(new_n5525_), .A3(new_n11192_), .ZN(new_n11369_));
  NOR3_X1    g08933(.A1(new_n11369_), .A2(new_n8058_), .A3(new_n11367_), .ZN(new_n11370_));
  INV_X1     g08934(.I(new_n11370_), .ZN(new_n11371_));
  NOR2_X1    g08935(.A1(new_n11348_), .A2(new_n2724_), .ZN(new_n11372_));
  NOR2_X1    g08936(.A1(new_n11360_), .A2(pi0142), .ZN(new_n11373_));
  OAI21_X1   g08937(.A1(new_n11373_), .A2(new_n11372_), .B(new_n5524_), .ZN(new_n11374_));
  NOR2_X1    g08938(.A1(new_n11235_), .A2(new_n5437_), .ZN(new_n11375_));
  INV_X1     g08939(.I(new_n11375_), .ZN(new_n11376_));
  NOR2_X1    g08940(.A1(new_n11376_), .A2(new_n5524_), .ZN(new_n11377_));
  NOR3_X1    g08941(.A1(new_n11377_), .A2(pi0144), .A3(new_n11367_), .ZN(new_n11378_));
  NAND2_X1   g08942(.A1(new_n11374_), .A2(new_n11378_), .ZN(new_n11379_));
  NAND3_X1   g08943(.A1(new_n11379_), .A2(new_n5658_), .A3(new_n11371_), .ZN(new_n11380_));
  INV_X1     g08944(.I(new_n11378_), .ZN(new_n11381_));
  INV_X1     g08945(.I(new_n11243_), .ZN(new_n11382_));
  NAND2_X1   g08946(.A1(new_n11382_), .A2(new_n11194_), .ZN(new_n11383_));
  NAND3_X1   g08947(.A1(new_n11383_), .A2(new_n7519_), .A3(new_n11161_), .ZN(new_n11384_));
  AOI21_X1   g08948(.A1(new_n11384_), .A2(new_n11370_), .B(new_n5658_), .ZN(new_n11385_));
  NOR2_X1    g08949(.A1(new_n11190_), .A2(new_n2631_), .ZN(new_n11386_));
  AOI22_X1   g08950(.A1(new_n11374_), .A2(new_n7525_), .B1(new_n11351_), .B2(new_n11386_), .ZN(new_n11387_));
  OAI21_X1   g08951(.A1(new_n11381_), .A2(new_n11387_), .B(new_n11385_), .ZN(new_n11388_));
  NAND3_X1   g08952(.A1(new_n11388_), .A2(new_n2628_), .A3(new_n11380_), .ZN(new_n11389_));
  INV_X1     g08953(.I(new_n8033_), .ZN(new_n11390_));
  NOR2_X1    g08954(.A1(new_n11363_), .A2(new_n11390_), .ZN(new_n11391_));
  AOI21_X1   g08955(.A1(new_n11391_), .A2(new_n11340_), .B(new_n5666_), .ZN(new_n11392_));
  AND3_X2    g08956(.A1(new_n11365_), .A2(new_n11389_), .A3(new_n11392_), .Z(new_n11393_));
  NOR3_X1    g08957(.A1(new_n11238_), .A2(new_n2821_), .A3(new_n2536_), .ZN(new_n11394_));
  INV_X1     g08958(.I(new_n11394_), .ZN(new_n11395_));
  NAND2_X1   g08959(.A1(new_n11282_), .A2(new_n11395_), .ZN(new_n11396_));
  NOR2_X1    g08960(.A1(new_n11396_), .A2(new_n11217_), .ZN(new_n11397_));
  NAND2_X1   g08961(.A1(new_n2627_), .A2(new_n5666_), .ZN(new_n11398_));
  OAI22_X1   g08962(.A1(new_n11393_), .A2(new_n11339_), .B1(new_n11397_), .B2(new_n11398_), .ZN(new_n11399_));
  INV_X1     g08963(.I(new_n7504_), .ZN(new_n11400_));
  INV_X1     g08964(.I(new_n11397_), .ZN(new_n11401_));
  NAND3_X1   g08965(.A1(new_n11401_), .A2(new_n7689_), .A3(new_n11341_), .ZN(new_n11402_));
  NOR2_X1    g08966(.A1(new_n11397_), .A2(new_n5398_), .ZN(new_n11403_));
  INV_X1     g08967(.I(new_n11396_), .ZN(new_n11404_));
  NOR2_X1    g08968(.A1(new_n11404_), .A2(new_n11207_), .ZN(new_n11405_));
  NOR2_X1    g08969(.A1(new_n11403_), .A2(new_n11405_), .ZN(new_n11406_));
  NOR2_X1    g08970(.A1(new_n11303_), .A2(new_n5398_), .ZN(new_n11407_));
  NOR2_X1    g08971(.A1(new_n11407_), .A2(new_n11164_), .ZN(new_n11408_));
  OAI21_X1   g08972(.A1(new_n11321_), .A2(new_n11408_), .B(new_n11406_), .ZN(new_n11409_));
  AOI21_X1   g08973(.A1(new_n11409_), .A2(new_n7731_), .B(new_n3360_), .ZN(new_n11410_));
  AOI21_X1   g08974(.A1(new_n11410_), .A2(new_n11402_), .B(pi0156), .ZN(new_n11411_));
  INV_X1     g08975(.I(new_n11403_), .ZN(new_n11412_));
  NOR2_X1    g08976(.A1(new_n8379_), .A2(new_n2821_), .ZN(new_n11413_));
  INV_X1     g08977(.I(new_n11413_), .ZN(new_n11414_));
  AOI21_X1   g08978(.A1(new_n11414_), .A2(new_n2744_), .B(new_n5437_), .ZN(new_n11415_));
  NOR2_X1    g08979(.A1(new_n11291_), .A2(new_n11415_), .ZN(new_n11416_));
  AOI21_X1   g08980(.A1(new_n11416_), .A2(new_n11412_), .B(new_n3107_), .ZN(new_n11417_));
  OAI21_X1   g08981(.A1(new_n11289_), .A2(pi0072), .B(new_n5558_), .ZN(new_n11418_));
  NOR2_X1    g08982(.A1(new_n11418_), .A2(new_n5437_), .ZN(new_n11419_));
  INV_X1     g08983(.I(new_n11419_), .ZN(new_n11420_));
  AOI21_X1   g08984(.A1(new_n11420_), .A2(new_n11412_), .B(pi0146), .ZN(new_n11421_));
  OAI21_X1   g08985(.A1(new_n11421_), .A2(new_n11417_), .B(new_n7731_), .ZN(new_n11422_));
  NOR2_X1    g08986(.A1(new_n11401_), .A2(new_n5398_), .ZN(new_n11423_));
  INV_X1     g08987(.I(new_n11298_), .ZN(new_n11424_));
  NOR2_X1    g08988(.A1(new_n11424_), .A2(new_n11413_), .ZN(new_n11425_));
  INV_X1     g08989(.I(new_n11425_), .ZN(new_n11426_));
  NOR2_X1    g08990(.A1(new_n11426_), .A2(new_n5437_), .ZN(new_n11427_));
  NOR3_X1    g08991(.A1(new_n11427_), .A2(new_n3107_), .A3(new_n11423_), .ZN(new_n11428_));
  NOR2_X1    g08992(.A1(new_n11296_), .A2(new_n2749_), .ZN(new_n11429_));
  NOR2_X1    g08993(.A1(new_n11429_), .A2(pi0072), .ZN(new_n11430_));
  NOR2_X1    g08994(.A1(new_n11430_), .A2(new_n5559_), .ZN(new_n11431_));
  NAND2_X1   g08995(.A1(new_n11431_), .A2(new_n5398_), .ZN(new_n11432_));
  INV_X1     g08996(.I(new_n11432_), .ZN(new_n11433_));
  NOR2_X1    g08997(.A1(new_n11433_), .A2(new_n11403_), .ZN(new_n11434_));
  NOR2_X1    g08998(.A1(new_n11434_), .A2(pi0146), .ZN(new_n11435_));
  OAI21_X1   g08999(.A1(new_n11428_), .A2(new_n11435_), .B(new_n7689_), .ZN(new_n11436_));
  NAND3_X1   g09000(.A1(new_n11436_), .A2(new_n3360_), .A3(new_n11422_), .ZN(new_n11437_));
  NAND2_X1   g09001(.A1(new_n11437_), .A2(new_n11411_), .ZN(new_n11438_));
  INV_X1     g09002(.I(new_n11408_), .ZN(new_n11439_));
  NOR2_X1    g09003(.A1(new_n11439_), .A2(new_n11394_), .ZN(new_n11440_));
  NAND2_X1   g09004(.A1(new_n11440_), .A2(pi0144), .ZN(new_n11441_));
  NOR2_X1    g09005(.A1(new_n11403_), .A2(new_n11415_), .ZN(new_n11442_));
  INV_X1     g09006(.I(new_n11442_), .ZN(new_n11443_));
  OAI21_X1   g09007(.A1(pi0144), .A2(new_n11443_), .B(new_n11441_), .ZN(new_n11444_));
  OAI21_X1   g09008(.A1(new_n11444_), .A2(new_n11190_), .B(pi0180), .ZN(new_n11445_));
  NAND2_X1   g09009(.A1(new_n11440_), .A2(new_n11218_), .ZN(new_n11446_));
  AOI21_X1   g09010(.A1(new_n11446_), .A2(new_n11191_), .B(pi0180), .ZN(new_n11447_));
  INV_X1     g09011(.I(new_n11228_), .ZN(new_n11448_));
  AOI21_X1   g09012(.A1(new_n11442_), .A2(new_n11448_), .B(new_n2724_), .ZN(new_n11449_));
  AOI21_X1   g09013(.A1(new_n2821_), .A2(new_n11225_), .B(new_n5559_), .ZN(new_n11450_));
  INV_X1     g09014(.I(new_n11450_), .ZN(new_n11451_));
  NOR2_X1    g09015(.A1(new_n11451_), .A2(new_n5437_), .ZN(new_n11452_));
  INV_X1     g09016(.I(new_n11452_), .ZN(new_n11453_));
  AOI21_X1   g09017(.A1(new_n11412_), .A2(new_n11453_), .B(pi0142), .ZN(new_n11454_));
  OAI21_X1   g09018(.A1(new_n11449_), .A2(new_n11454_), .B(new_n8058_), .ZN(new_n11455_));
  AOI21_X1   g09019(.A1(new_n11455_), .A2(new_n11447_), .B(new_n9627_), .ZN(new_n11456_));
  NAND2_X1   g09020(.A1(new_n11456_), .A2(new_n11445_), .ZN(new_n11457_));
  OR3_X2     g09021(.A1(new_n11427_), .A2(new_n2724_), .A3(new_n11423_), .Z(new_n11458_));
  OAI21_X1   g09022(.A1(pi0142), .A2(new_n11434_), .B(new_n11458_), .ZN(new_n11459_));
  OAI21_X1   g09023(.A1(new_n11397_), .A2(new_n11268_), .B(new_n5657_), .ZN(new_n11460_));
  AOI21_X1   g09024(.A1(new_n11459_), .A2(new_n8058_), .B(new_n11460_), .ZN(new_n11461_));
  OAI21_X1   g09025(.A1(new_n11285_), .A2(new_n11408_), .B(new_n11406_), .ZN(new_n11462_));
  NAND2_X1   g09026(.A1(new_n11462_), .A2(pi0144), .ZN(new_n11463_));
  AOI21_X1   g09027(.A1(new_n11416_), .A2(new_n11412_), .B(new_n2724_), .ZN(new_n11464_));
  AOI21_X1   g09028(.A1(new_n11420_), .A2(new_n11412_), .B(pi0142), .ZN(new_n11465_));
  OAI21_X1   g09029(.A1(new_n11465_), .A2(new_n11464_), .B(new_n8058_), .ZN(new_n11466_));
  NAND3_X1   g09030(.A1(new_n11466_), .A2(pi0180), .A3(new_n11463_), .ZN(new_n11467_));
  NAND2_X1   g09031(.A1(new_n11467_), .A2(new_n9627_), .ZN(new_n11468_));
  OAI21_X1   g09032(.A1(new_n11461_), .A2(new_n11468_), .B(new_n11457_), .ZN(new_n11469_));
  INV_X1     g09033(.I(new_n7689_), .ZN(new_n11470_));
  NAND2_X1   g09034(.A1(new_n11395_), .A2(new_n11161_), .ZN(new_n11471_));
  NOR2_X1    g09035(.A1(new_n11471_), .A2(new_n11207_), .ZN(new_n11472_));
  AOI21_X1   g09036(.A1(new_n11472_), .A2(new_n11218_), .B(new_n11157_), .ZN(new_n11473_));
  AOI21_X1   g09037(.A1(pi0146), .A2(new_n11171_), .B(new_n11473_), .ZN(new_n11474_));
  NOR3_X1    g09038(.A1(new_n11423_), .A2(new_n3360_), .A3(new_n11474_), .ZN(new_n11475_));
  OAI21_X1   g09039(.A1(new_n11443_), .A2(new_n11228_), .B(pi0146), .ZN(new_n11476_));
  OAI21_X1   g09040(.A1(new_n11403_), .A2(new_n11452_), .B(new_n3107_), .ZN(new_n11477_));
  AOI21_X1   g09041(.A1(new_n11476_), .A2(new_n11477_), .B(pi0161), .ZN(new_n11478_));
  NOR2_X1    g09042(.A1(new_n11478_), .A2(new_n11475_), .ZN(new_n11479_));
  NAND2_X1   g09043(.A1(new_n11471_), .A2(new_n11206_), .ZN(new_n11480_));
  INV_X1     g09044(.I(new_n11480_), .ZN(new_n11481_));
  NOR3_X1    g09045(.A1(new_n11403_), .A2(pi0146), .A3(new_n11481_), .ZN(new_n11482_));
  NOR3_X1    g09046(.A1(new_n11439_), .A2(new_n3107_), .A3(new_n11394_), .ZN(new_n11483_));
  NOR3_X1    g09047(.A1(new_n11482_), .A2(new_n11483_), .A3(new_n3360_), .ZN(new_n11484_));
  NOR3_X1    g09048(.A1(new_n11442_), .A2(pi0161), .A3(new_n11159_), .ZN(new_n11485_));
  NOR2_X1    g09049(.A1(new_n11484_), .A2(new_n11485_), .ZN(new_n11486_));
  OAI22_X1   g09050(.A1(new_n11479_), .A2(new_n11470_), .B1(new_n11486_), .B2(new_n11313_), .ZN(new_n11487_));
  AOI22_X1   g09051(.A1(new_n11469_), .A2(new_n2628_), .B1(pi0156), .B2(new_n11487_), .ZN(new_n11488_));
  AOI21_X1   g09052(.A1(new_n11488_), .A2(new_n11438_), .B(new_n11400_), .ZN(new_n11489_));
  OAI21_X1   g09053(.A1(new_n11489_), .A2(new_n11399_), .B(new_n3265_), .ZN(new_n11490_));
  AOI21_X1   g09054(.A1(new_n11490_), .A2(new_n11334_), .B(new_n11333_), .ZN(new_n11491_));
  INV_X1     g09055(.I(new_n11199_), .ZN(new_n11492_));
  NOR2_X1    g09056(.A1(new_n11492_), .A2(new_n11163_), .ZN(new_n11493_));
  NAND2_X1   g09057(.A1(new_n11198_), .A2(new_n11493_), .ZN(new_n11494_));
  NAND3_X1   g09058(.A1(new_n11494_), .A2(new_n11183_), .A3(new_n11188_), .ZN(new_n11495_));
  AOI21_X1   g09059(.A1(new_n11491_), .A2(new_n11330_), .B(new_n11495_), .ZN(new_n11496_));
  OAI21_X1   g09060(.A1(new_n11496_), .A2(new_n11329_), .B(new_n11185_), .ZN(po0279));
  AND2_X2    g09061(.A1(new_n11125_), .A2(new_n6645_), .Z(new_n11498_));
  OAI21_X1   g09062(.A1(new_n11498_), .A2(new_n6350_), .B(new_n6643_), .ZN(new_n11499_));
  AOI21_X1   g09063(.A1(new_n11149_), .A2(new_n6645_), .B(new_n10925_), .ZN(new_n11500_));
  NAND2_X1   g09064(.A1(new_n10093_), .A2(po1038), .ZN(new_n11501_));
  OAI22_X1   g09065(.A1(new_n11500_), .A2(new_n11499_), .B1(new_n6349_), .B2(new_n11501_), .ZN(po0280));
  NOR2_X1    g09066(.A1(new_n2610_), .A2(pi0038), .ZN(new_n11503_));
  NOR4_X1    g09067(.A1(new_n7607_), .A2(pi0110), .A3(new_n5451_), .A4(new_n11335_), .ZN(new_n11504_));
  NAND4_X1   g09068(.A1(new_n7606_), .A2(new_n5423_), .A3(new_n2509_), .A4(new_n5549_), .ZN(new_n11505_));
  OAI21_X1   g09069(.A1(new_n11505_), .A2(new_n2628_), .B(pi0039), .ZN(new_n11506_));
  INV_X1     g09070(.I(new_n10524_), .ZN(new_n11507_));
  OAI21_X1   g09071(.A1(new_n11507_), .A2(new_n2509_), .B(new_n2627_), .ZN(new_n11508_));
  OAI22_X1   g09072(.A1(new_n11508_), .A2(new_n11503_), .B1(new_n11506_), .B2(new_n11504_), .ZN(new_n11509_));
  INV_X1     g09073(.I(new_n5567_), .ZN(new_n11510_));
  NOR2_X1    g09074(.A1(new_n5574_), .A2(pi0111), .ZN(new_n11511_));
  NOR2_X1    g09075(.A1(new_n11511_), .A2(new_n2949_), .ZN(new_n11512_));
  NAND3_X1   g09076(.A1(new_n11512_), .A2(new_n7416_), .A3(new_n2476_), .ZN(new_n11513_));
  NAND2_X1   g09077(.A1(pi0067), .A2(pi0069), .ZN(new_n11514_));
  NAND3_X1   g09078(.A1(new_n2902_), .A2(new_n2824_), .A3(new_n11514_), .ZN(new_n11515_));
  NAND3_X1   g09079(.A1(new_n11513_), .A2(new_n8904_), .A3(new_n11515_), .ZN(new_n11516_));
  AOI21_X1   g09080(.A1(new_n11516_), .A2(new_n2909_), .B(pi0071), .ZN(new_n11517_));
  OAI21_X1   g09081(.A1(new_n11517_), .A2(new_n11510_), .B(new_n2500_), .ZN(new_n11518_));
  AOI21_X1   g09082(.A1(new_n11518_), .A2(new_n9228_), .B(pi0090), .ZN(new_n11519_));
  OR2_X2     g09083(.A1(new_n11519_), .A2(new_n2747_), .Z(new_n11520_));
  NOR3_X1    g09084(.A1(new_n11520_), .A2(pi0093), .A3(new_n2986_), .ZN(new_n11521_));
  OAI21_X1   g09085(.A1(new_n11521_), .A2(pi0072), .B(new_n5558_), .ZN(new_n11522_));
  OAI21_X1   g09086(.A1(new_n11522_), .A2(new_n10524_), .B(new_n2627_), .ZN(new_n11523_));
  AOI21_X1   g09087(.A1(new_n2842_), .A2(new_n7272_), .B(new_n2985_), .ZN(new_n11524_));
  NOR4_X1    g09088(.A1(new_n11520_), .A2(pi0072), .A3(pi0093), .A4(new_n11524_), .ZN(new_n11525_));
  NOR3_X1    g09089(.A1(new_n8412_), .A2(new_n2821_), .A3(new_n2749_), .ZN(new_n11526_));
  OAI21_X1   g09090(.A1(new_n11525_), .A2(new_n11526_), .B(new_n2535_), .ZN(new_n11527_));
  AOI21_X1   g09091(.A1(new_n11527_), .A2(new_n2509_), .B(new_n11507_), .ZN(new_n11528_));
  NOR2_X1    g09092(.A1(new_n11528_), .A2(new_n11523_), .ZN(new_n11529_));
  AOI21_X1   g09093(.A1(new_n11529_), .A2(new_n11503_), .B(new_n11509_), .ZN(new_n11530_));
  NOR4_X1    g09094(.A1(new_n5323_), .A2(new_n2509_), .A3(new_n8220_), .A4(new_n8847_), .ZN(new_n11531_));
  OAI21_X1   g09095(.A1(new_n11531_), .A2(pi0039), .B(po1038), .ZN(new_n11532_));
  AOI21_X1   g09096(.A1(new_n11505_), .A2(pi0039), .B(new_n11532_), .ZN(new_n11533_));
  AOI21_X1   g09097(.A1(new_n11530_), .A2(new_n6643_), .B(new_n11533_), .ZN(po0281));
  NOR2_X1    g09098(.A1(new_n7985_), .A2(new_n2628_), .ZN(new_n11535_));
  AOI21_X1   g09099(.A1(pi0140), .A2(new_n2628_), .B(new_n11535_), .ZN(new_n11536_));
  OAI21_X1   g09100(.A1(new_n6698_), .A2(new_n11536_), .B(pi0087), .ZN(new_n11537_));
  AND2_X2    g09101(.A1(pi0125), .A2(pi0133), .Z(new_n11538_));
  AOI21_X1   g09102(.A1(new_n11179_), .A2(new_n11180_), .B(new_n11538_), .ZN(new_n11539_));
  NOR2_X1    g09103(.A1(new_n11158_), .A2(new_n7858_), .ZN(new_n11540_));
  OAI21_X1   g09104(.A1(new_n11376_), .A2(pi0174), .B(new_n2628_), .ZN(new_n11541_));
  NOR2_X1    g09105(.A1(new_n11541_), .A2(new_n11540_), .ZN(new_n11542_));
  NOR2_X1    g09106(.A1(new_n11158_), .A2(new_n3778_), .ZN(new_n11543_));
  NOR2_X1    g09107(.A1(new_n11376_), .A2(pi0152), .ZN(new_n11544_));
  NOR2_X1    g09108(.A1(new_n11544_), .A2(new_n11543_), .ZN(new_n11545_));
  INV_X1     g09109(.I(new_n11545_), .ZN(new_n11546_));
  NOR2_X1    g09110(.A1(new_n11546_), .A2(new_n2628_), .ZN(new_n11547_));
  NOR3_X1    g09111(.A1(new_n11547_), .A2(new_n5666_), .A3(new_n11542_), .ZN(new_n11548_));
  INV_X1     g09112(.I(new_n11548_), .ZN(new_n11549_));
  AOI21_X1   g09113(.A1(new_n11549_), .A2(new_n11199_), .B(new_n11539_), .ZN(new_n11550_));
  NAND2_X1   g09114(.A1(new_n11550_), .A2(new_n11537_), .ZN(new_n11551_));
  NOR2_X1    g09115(.A1(new_n11549_), .A2(new_n2702_), .ZN(new_n11552_));
  INV_X1     g09116(.I(new_n11552_), .ZN(new_n11553_));
  AOI21_X1   g09117(.A1(new_n11414_), .A2(new_n5666_), .B(pi0039), .ZN(new_n11554_));
  NOR2_X1    g09118(.A1(new_n11554_), .A2(pi0038), .ZN(new_n11555_));
  AOI21_X1   g09119(.A1(new_n2628_), .A2(new_n6744_), .B(new_n6810_), .ZN(new_n11556_));
  INV_X1     g09120(.I(new_n11556_), .ZN(new_n11557_));
  NAND2_X1   g09121(.A1(new_n2531_), .A2(new_n11557_), .ZN(new_n11558_));
  AOI21_X1   g09122(.A1(new_n11558_), .A2(new_n5666_), .B(new_n2627_), .ZN(new_n11559_));
  INV_X1     g09123(.I(new_n11241_), .ZN(new_n11560_));
  NOR2_X1    g09124(.A1(new_n2531_), .A2(new_n5398_), .ZN(new_n11561_));
  AOI21_X1   g09125(.A1(new_n11560_), .A2(new_n5398_), .B(new_n11561_), .ZN(new_n11562_));
  OAI21_X1   g09126(.A1(new_n6744_), .A2(new_n11164_), .B(new_n11562_), .ZN(new_n11563_));
  NAND2_X1   g09127(.A1(new_n11563_), .A2(new_n7488_), .ZN(new_n11564_));
  NAND2_X1   g09128(.A1(new_n2531_), .A2(new_n6744_), .ZN(new_n11565_));
  NAND2_X1   g09129(.A1(new_n11565_), .A2(pi0174), .ZN(new_n11566_));
  AOI21_X1   g09130(.A1(new_n11564_), .A2(new_n11566_), .B(new_n11540_), .ZN(new_n11567_));
  OAI21_X1   g09131(.A1(new_n11567_), .A2(pi0180), .B(new_n2628_), .ZN(new_n11568_));
  INV_X1     g09132(.I(new_n11377_), .ZN(new_n11569_));
  INV_X1     g09133(.I(new_n11562_), .ZN(new_n11570_));
  NOR2_X1    g09134(.A1(new_n11570_), .A2(pi0224), .ZN(new_n11571_));
  NOR2_X1    g09135(.A1(new_n11382_), .A2(new_n2631_), .ZN(new_n11572_));
  OAI21_X1   g09136(.A1(new_n11572_), .A2(new_n11571_), .B(new_n5524_), .ZN(new_n11573_));
  NAND2_X1   g09137(.A1(new_n11573_), .A2(new_n11569_), .ZN(new_n11574_));
  NOR2_X1    g09138(.A1(new_n11574_), .A2(pi0174), .ZN(new_n11575_));
  INV_X1     g09139(.I(new_n11253_), .ZN(new_n11576_));
  AOI21_X1   g09140(.A1(new_n6759_), .A2(new_n11576_), .B(new_n2530_), .ZN(new_n11577_));
  NOR2_X1    g09141(.A1(new_n11577_), .A2(new_n7488_), .ZN(new_n11578_));
  OAI21_X1   g09142(.A1(new_n11575_), .A2(new_n11578_), .B(new_n7858_), .ZN(new_n11579_));
  NOR2_X1    g09143(.A1(new_n11346_), .A2(new_n5437_), .ZN(new_n11580_));
  NOR2_X1    g09144(.A1(new_n11580_), .A2(new_n11561_), .ZN(new_n11581_));
  NOR2_X1    g09145(.A1(new_n11581_), .A2(new_n6759_), .ZN(new_n11582_));
  OAI21_X1   g09146(.A1(new_n11336_), .A2(new_n11252_), .B(pi0224), .ZN(new_n11583_));
  AOI21_X1   g09147(.A1(new_n11583_), .A2(new_n5524_), .B(new_n11164_), .ZN(new_n11584_));
  NOR2_X1    g09148(.A1(new_n11582_), .A2(new_n11584_), .ZN(new_n11585_));
  NOR2_X1    g09149(.A1(new_n11255_), .A2(new_n11252_), .ZN(new_n11586_));
  NOR2_X1    g09150(.A1(new_n11586_), .A2(new_n11157_), .ZN(new_n11587_));
  AOI21_X1   g09151(.A1(new_n11587_), .A2(pi0224), .B(new_n5525_), .ZN(new_n11588_));
  INV_X1     g09152(.I(new_n11588_), .ZN(new_n11589_));
  NOR2_X1    g09153(.A1(new_n11345_), .A2(new_n11561_), .ZN(new_n11590_));
  NOR2_X1    g09154(.A1(new_n11590_), .A2(new_n6759_), .ZN(new_n11591_));
  OAI21_X1   g09155(.A1(new_n11591_), .A2(new_n11589_), .B(new_n11158_), .ZN(new_n11592_));
  INV_X1     g09156(.I(new_n11592_), .ZN(new_n11593_));
  NAND2_X1   g09157(.A1(new_n11593_), .A2(pi0174), .ZN(new_n11594_));
  OAI21_X1   g09158(.A1(pi0174), .A2(new_n11585_), .B(new_n11594_), .ZN(new_n11595_));
  AOI21_X1   g09159(.A1(new_n11595_), .A2(pi0193), .B(new_n5657_), .ZN(new_n11596_));
  AOI21_X1   g09160(.A1(new_n11579_), .A2(new_n11596_), .B(new_n11568_), .ZN(new_n11597_));
  OAI21_X1   g09161(.A1(new_n11545_), .A2(new_n5549_), .B(new_n7731_), .ZN(new_n11598_));
  INV_X1     g09162(.I(new_n11590_), .ZN(new_n11599_));
  NAND2_X1   g09163(.A1(new_n11599_), .A2(pi0152), .ZN(new_n11600_));
  INV_X1     g09164(.I(new_n11581_), .ZN(new_n11601_));
  NAND2_X1   g09165(.A1(new_n11601_), .A2(new_n3369_), .ZN(new_n11602_));
  NAND2_X1   g09166(.A1(new_n3778_), .A2(pi0051), .ZN(new_n11603_));
  NAND3_X1   g09167(.A1(new_n11602_), .A2(new_n11600_), .A3(new_n11603_), .ZN(new_n11604_));
  NAND2_X1   g09168(.A1(new_n11604_), .A2(new_n2614_), .ZN(new_n11605_));
  AOI21_X1   g09169(.A1(new_n11239_), .A2(new_n11251_), .B(new_n11164_), .ZN(new_n11606_));
  NOR2_X1    g09170(.A1(new_n11606_), .A2(pi0152), .ZN(new_n11607_));
  NOR2_X1    g09171(.A1(new_n11587_), .A2(new_n3369_), .ZN(new_n11608_));
  OAI21_X1   g09172(.A1(new_n11607_), .A2(new_n11608_), .B(pi0172), .ZN(new_n11609_));
  NAND2_X1   g09173(.A1(new_n11245_), .A2(pi0152), .ZN(new_n11610_));
  OAI21_X1   g09174(.A1(new_n11382_), .A2(pi0152), .B(new_n11610_), .ZN(new_n11611_));
  AOI21_X1   g09175(.A1(new_n11611_), .A2(new_n3778_), .B(new_n2614_), .ZN(new_n11612_));
  AOI21_X1   g09176(.A1(new_n11612_), .A2(new_n11609_), .B(new_n5550_), .ZN(new_n11613_));
  AOI21_X1   g09177(.A1(new_n11613_), .A2(new_n11605_), .B(new_n11598_), .ZN(new_n11614_));
  NOR2_X1    g09178(.A1(new_n11545_), .A2(new_n5549_), .ZN(new_n11615_));
  OR2_X2     g09179(.A1(new_n11605_), .A2(new_n11615_), .Z(new_n11616_));
  NAND2_X1   g09180(.A1(new_n11545_), .A2(new_n6762_), .ZN(new_n11617_));
  AOI21_X1   g09181(.A1(new_n11616_), .A2(new_n11617_), .B(new_n11470_), .ZN(new_n11618_));
  NOR3_X1    g09182(.A1(new_n11597_), .A2(new_n11614_), .A3(new_n11618_), .ZN(new_n11619_));
  OAI21_X1   g09183(.A1(new_n11619_), .A2(new_n5666_), .B(new_n11559_), .ZN(new_n11620_));
  OAI21_X1   g09184(.A1(new_n11548_), .A2(new_n3265_), .B(new_n2702_), .ZN(new_n11621_));
  AOI21_X1   g09185(.A1(new_n11620_), .A2(new_n11555_), .B(new_n11621_), .ZN(new_n11622_));
  NAND2_X1   g09186(.A1(pi0152), .A2(pi0197), .ZN(new_n11623_));
  NOR2_X1    g09187(.A1(new_n11414_), .A2(new_n5398_), .ZN(new_n11624_));
  NOR2_X1    g09188(.A1(new_n11452_), .A2(new_n11624_), .ZN(new_n11625_));
  NAND2_X1   g09189(.A1(new_n11625_), .A2(new_n3778_), .ZN(new_n11626_));
  NOR3_X1    g09190(.A1(new_n11413_), .A2(new_n11157_), .A3(new_n11228_), .ZN(new_n11627_));
  NAND2_X1   g09191(.A1(new_n11627_), .A2(pi0172), .ZN(new_n11628_));
  AOI21_X1   g09192(.A1(new_n11626_), .A2(new_n11628_), .B(new_n11623_), .ZN(new_n11629_));
  AOI21_X1   g09193(.A1(new_n11481_), .A2(new_n3369_), .B(pi0197), .ZN(new_n11630_));
  NOR2_X1    g09194(.A1(new_n5437_), .A2(pi0152), .ZN(new_n11631_));
  OAI21_X1   g09195(.A1(new_n11414_), .A2(new_n11631_), .B(new_n11630_), .ZN(new_n11632_));
  NOR2_X1    g09196(.A1(new_n11413_), .A2(new_n5398_), .ZN(new_n11633_));
  INV_X1     g09197(.I(new_n11633_), .ZN(new_n11634_));
  NAND2_X1   g09198(.A1(new_n11634_), .A2(new_n11473_), .ZN(new_n11635_));
  NAND3_X1   g09199(.A1(new_n11635_), .A2(new_n3369_), .A3(pi0197), .ZN(new_n11636_));
  AOI21_X1   g09200(.A1(new_n11636_), .A2(new_n11632_), .B(new_n11543_), .ZN(new_n11637_));
  OAI21_X1   g09201(.A1(new_n11629_), .A2(new_n11637_), .B(new_n8066_), .ZN(new_n11638_));
  INV_X1     g09202(.I(new_n11472_), .ZN(new_n11639_));
  NOR2_X1    g09203(.A1(new_n11396_), .A2(new_n11639_), .ZN(new_n11640_));
  NOR2_X1    g09204(.A1(new_n11640_), .A2(new_n11633_), .ZN(new_n11641_));
  NOR2_X1    g09205(.A1(new_n11641_), .A2(pi0152), .ZN(new_n11642_));
  NOR3_X1    g09206(.A1(new_n11291_), .A2(new_n11157_), .A3(new_n11413_), .ZN(new_n11643_));
  INV_X1     g09207(.I(new_n11643_), .ZN(new_n11644_));
  NOR2_X1    g09208(.A1(new_n11644_), .A2(new_n3369_), .ZN(new_n11645_));
  OAI21_X1   g09209(.A1(new_n11645_), .A2(new_n11642_), .B(pi0172), .ZN(new_n11646_));
  NOR2_X1    g09210(.A1(new_n11419_), .A2(new_n11624_), .ZN(new_n11647_));
  INV_X1     g09211(.I(new_n11647_), .ZN(new_n11648_));
  NOR2_X1    g09212(.A1(new_n11648_), .A2(new_n3369_), .ZN(new_n11649_));
  NOR2_X1    g09213(.A1(new_n11405_), .A2(new_n11624_), .ZN(new_n11650_));
  INV_X1     g09214(.I(new_n11650_), .ZN(new_n11651_));
  NOR2_X1    g09215(.A1(new_n11651_), .A2(pi0152), .ZN(new_n11652_));
  OAI21_X1   g09216(.A1(new_n11649_), .A2(new_n11652_), .B(new_n3778_), .ZN(new_n11653_));
  NAND3_X1   g09217(.A1(new_n11653_), .A2(new_n11646_), .A3(new_n5636_), .ZN(new_n11654_));
  NOR2_X1    g09218(.A1(new_n11433_), .A2(new_n11624_), .ZN(new_n11655_));
  INV_X1     g09219(.I(new_n11655_), .ZN(new_n11656_));
  NOR2_X1    g09220(.A1(new_n11656_), .A2(pi0172), .ZN(new_n11657_));
  NOR2_X1    g09221(.A1(new_n11299_), .A2(new_n11413_), .ZN(new_n11658_));
  INV_X1     g09222(.I(new_n11658_), .ZN(new_n11659_));
  NOR2_X1    g09223(.A1(new_n11659_), .A2(new_n3778_), .ZN(new_n11660_));
  OAI21_X1   g09224(.A1(new_n11657_), .A2(new_n11660_), .B(pi0152), .ZN(new_n11661_));
  AOI21_X1   g09225(.A1(new_n11401_), .A2(new_n11206_), .B(new_n11624_), .ZN(new_n11662_));
  INV_X1     g09226(.I(new_n11662_), .ZN(new_n11663_));
  NOR3_X1    g09227(.A1(new_n11663_), .A2(pi0152), .A3(new_n11543_), .ZN(new_n11664_));
  NOR2_X1    g09228(.A1(new_n11664_), .A2(new_n5636_), .ZN(new_n11665_));
  NAND2_X1   g09229(.A1(new_n11661_), .A2(new_n11665_), .ZN(new_n11666_));
  NAND4_X1   g09230(.A1(new_n11666_), .A2(new_n3265_), .A3(pi0155), .A4(new_n11654_), .ZN(new_n11667_));
  AOI21_X1   g09231(.A1(new_n11667_), .A2(new_n11638_), .B(new_n2628_), .ZN(new_n11668_));
  INV_X1     g09232(.I(new_n8057_), .ZN(new_n11669_));
  OR3_X2     g09233(.A1(new_n11663_), .A2(new_n5656_), .A3(new_n11540_), .Z(new_n11670_));
  NAND2_X1   g09234(.A1(new_n11650_), .A2(new_n7858_), .ZN(new_n11671_));
  OAI21_X1   g09235(.A1(new_n7858_), .A2(new_n11641_), .B(new_n11671_), .ZN(new_n11672_));
  AOI21_X1   g09236(.A1(new_n11672_), .A2(new_n5656_), .B(pi0174), .ZN(new_n11673_));
  AOI21_X1   g09237(.A1(new_n11673_), .A2(new_n11670_), .B(new_n11669_), .ZN(new_n11674_));
  NAND2_X1   g09238(.A1(new_n11655_), .A2(pi0145), .ZN(new_n11675_));
  NAND2_X1   g09239(.A1(new_n11647_), .A2(new_n5656_), .ZN(new_n11676_));
  AOI21_X1   g09240(.A1(new_n11675_), .A2(new_n11676_), .B(pi0193), .ZN(new_n11677_));
  NOR2_X1    g09241(.A1(new_n11644_), .A2(pi0145), .ZN(new_n11678_));
  AOI21_X1   g09242(.A1(pi0145), .A2(new_n11658_), .B(new_n11678_), .ZN(new_n11679_));
  OAI21_X1   g09243(.A1(new_n11679_), .A2(new_n7858_), .B(pi0174), .ZN(new_n11680_));
  OAI21_X1   g09244(.A1(new_n11677_), .A2(new_n11680_), .B(new_n11674_), .ZN(new_n11681_));
  AOI21_X1   g09245(.A1(new_n11218_), .A2(new_n11158_), .B(new_n5656_), .ZN(new_n11682_));
  NOR2_X1    g09246(.A1(new_n11682_), .A2(new_n11639_), .ZN(new_n11683_));
  NOR3_X1    g09247(.A1(new_n11633_), .A2(new_n11683_), .A3(pi0174), .ZN(new_n11684_));
  NAND2_X1   g09248(.A1(new_n11228_), .A2(new_n5656_), .ZN(new_n11685_));
  OAI21_X1   g09249(.A1(new_n11157_), .A2(new_n11228_), .B(new_n11685_), .ZN(new_n11686_));
  AOI21_X1   g09250(.A1(new_n11414_), .A2(new_n11686_), .B(new_n7488_), .ZN(new_n11687_));
  NOR3_X1    g09251(.A1(new_n11684_), .A2(new_n7858_), .A3(new_n11687_), .ZN(new_n11688_));
  INV_X1     g09252(.I(new_n11635_), .ZN(new_n11689_));
  NOR2_X1    g09253(.A1(new_n11689_), .A2(new_n5656_), .ZN(new_n11690_));
  NOR2_X1    g09254(.A1(new_n11624_), .A2(new_n11481_), .ZN(new_n11691_));
  INV_X1     g09255(.I(new_n11691_), .ZN(new_n11692_));
  NOR2_X1    g09256(.A1(new_n11692_), .A2(pi0145), .ZN(new_n11693_));
  OAI21_X1   g09257(.A1(new_n11693_), .A2(new_n11690_), .B(new_n7488_), .ZN(new_n11694_));
  INV_X1     g09258(.I(new_n11625_), .ZN(new_n11695_));
  NOR2_X1    g09259(.A1(new_n11695_), .A2(new_n5656_), .ZN(new_n11696_));
  NOR2_X1    g09260(.A1(new_n11413_), .A2(pi0145), .ZN(new_n11697_));
  OAI21_X1   g09261(.A1(new_n11696_), .A2(new_n11697_), .B(pi0174), .ZN(new_n11698_));
  AOI21_X1   g09262(.A1(new_n11698_), .A2(new_n11694_), .B(pi0193), .ZN(new_n11699_));
  OAI21_X1   g09263(.A1(new_n11699_), .A2(new_n11688_), .B(new_n7969_), .ZN(new_n11700_));
  AOI21_X1   g09264(.A1(new_n11681_), .A2(new_n11700_), .B(pi0038), .ZN(new_n11701_));
  OAI21_X1   g09265(.A1(new_n11668_), .A2(new_n11701_), .B(new_n7504_), .ZN(new_n11702_));
  AOI21_X1   g09266(.A1(new_n11702_), .A2(new_n11622_), .B(new_n2569_), .ZN(new_n11703_));
  AOI21_X1   g09267(.A1(new_n11703_), .A2(new_n11553_), .B(new_n11551_), .ZN(new_n11704_));
  NAND2_X1   g09268(.A1(new_n11549_), .A2(new_n11493_), .ZN(new_n11705_));
  NAND3_X1   g09269(.A1(new_n11705_), .A2(new_n11537_), .A3(new_n11539_), .ZN(new_n11706_));
  NAND3_X1   g09270(.A1(new_n11549_), .A2(pi0038), .A3(new_n11171_), .ZN(new_n11707_));
  AOI21_X1   g09271(.A1(new_n11314_), .A2(new_n5666_), .B(pi0039), .ZN(new_n11708_));
  AOI21_X1   g09272(.A1(new_n11239_), .A2(new_n7519_), .B(new_n11171_), .ZN(new_n11709_));
  INV_X1     g09273(.I(new_n11709_), .ZN(new_n11710_));
  NOR2_X1    g09274(.A1(new_n11336_), .A2(new_n8070_), .ZN(new_n11711_));
  NAND2_X1   g09275(.A1(new_n11163_), .A2(pi0299), .ZN(new_n11712_));
  OAI22_X1   g09276(.A1(new_n11710_), .A2(pi0299), .B1(new_n11711_), .B2(new_n11712_), .ZN(new_n11713_));
  NOR2_X1    g09277(.A1(new_n11713_), .A2(pi0232), .ZN(new_n11714_));
  NOR2_X1    g09278(.A1(new_n11714_), .A2(new_n2627_), .ZN(new_n11715_));
  INV_X1     g09279(.I(new_n11715_), .ZN(new_n11716_));
  NAND2_X1   g09280(.A1(new_n11353_), .A2(pi0180), .ZN(new_n11717_));
  NAND3_X1   g09281(.A1(new_n11717_), .A2(new_n11710_), .A3(pi0174), .ZN(new_n11718_));
  NOR2_X1    g09282(.A1(new_n11348_), .A2(new_n7525_), .ZN(new_n11719_));
  NOR2_X1    g09283(.A1(new_n11161_), .A2(new_n5398_), .ZN(new_n11720_));
  NOR3_X1    g09284(.A1(new_n11720_), .A2(new_n7519_), .A3(pi0051), .ZN(new_n11721_));
  NOR2_X1    g09285(.A1(new_n11719_), .A2(new_n11721_), .ZN(new_n11722_));
  INV_X1     g09286(.I(new_n11722_), .ZN(new_n11723_));
  AOI21_X1   g09287(.A1(pi0180), .A2(new_n11350_), .B(new_n11723_), .ZN(new_n11724_));
  NAND2_X1   g09288(.A1(new_n11724_), .A2(new_n7488_), .ZN(new_n11725_));
  NAND3_X1   g09289(.A1(new_n11725_), .A2(new_n7858_), .A3(new_n11718_), .ZN(new_n11726_));
  NOR2_X1    g09290(.A1(new_n11353_), .A2(pi0051), .ZN(new_n11727_));
  NOR2_X1    g09291(.A1(new_n11727_), .A2(new_n5437_), .ZN(new_n11728_));
  NOR3_X1    g09292(.A1(new_n11728_), .A2(new_n7488_), .A3(new_n11709_), .ZN(new_n11729_));
  AOI21_X1   g09293(.A1(new_n5398_), .A2(new_n8637_), .B(new_n11347_), .ZN(new_n11730_));
  AOI21_X1   g09294(.A1(new_n11171_), .A2(new_n5437_), .B(new_n7519_), .ZN(new_n11731_));
  INV_X1     g09295(.I(new_n11731_), .ZN(new_n11732_));
  OAI21_X1   g09296(.A1(new_n11730_), .A2(new_n7525_), .B(new_n11732_), .ZN(new_n11733_));
  NOR2_X1    g09297(.A1(new_n11733_), .A2(pi0174), .ZN(new_n11734_));
  OAI21_X1   g09298(.A1(new_n11734_), .A2(new_n11729_), .B(pi0180), .ZN(new_n11735_));
  NOR3_X1    g09299(.A1(new_n11709_), .A2(new_n7488_), .A3(new_n11157_), .ZN(new_n11736_));
  OAI21_X1   g09300(.A1(new_n11360_), .A2(new_n7525_), .B(new_n11732_), .ZN(new_n11737_));
  NOR2_X1    g09301(.A1(new_n11737_), .A2(pi0174), .ZN(new_n11738_));
  OAI21_X1   g09302(.A1(new_n11738_), .A2(new_n11736_), .B(new_n5657_), .ZN(new_n11739_));
  NAND3_X1   g09303(.A1(new_n11739_), .A2(new_n11735_), .A3(pi0193), .ZN(new_n11740_));
  NAND3_X1   g09304(.A1(new_n11726_), .A2(new_n2628_), .A3(new_n11740_), .ZN(new_n11741_));
  NAND2_X1   g09305(.A1(new_n11360_), .A2(new_n3369_), .ZN(new_n11742_));
  NAND2_X1   g09306(.A1(new_n11368_), .A2(pi0152), .ZN(new_n11743_));
  AOI21_X1   g09307(.A1(new_n11742_), .A2(new_n11743_), .B(new_n3778_), .ZN(new_n11744_));
  NAND2_X1   g09308(.A1(new_n11343_), .A2(new_n11631_), .ZN(new_n11745_));
  OAI21_X1   g09309(.A1(pi0152), .A2(new_n5437_), .B(new_n11240_), .ZN(new_n11746_));
  NAND3_X1   g09310(.A1(new_n11746_), .A2(new_n3778_), .A3(new_n11745_), .ZN(new_n11747_));
  NAND2_X1   g09311(.A1(new_n11747_), .A2(new_n7508_), .ZN(new_n11748_));
  OAI21_X1   g09312(.A1(new_n11744_), .A2(new_n11748_), .B(new_n5631_), .ZN(new_n11749_));
  NAND2_X1   g09313(.A1(new_n11354_), .A2(pi0152), .ZN(new_n11750_));
  NAND2_X1   g09314(.A1(new_n11351_), .A2(new_n3369_), .ZN(new_n11751_));
  AOI21_X1   g09315(.A1(new_n11751_), .A2(new_n11750_), .B(new_n11543_), .ZN(new_n11752_));
  OAI21_X1   g09316(.A1(new_n11752_), .A2(new_n8070_), .B(pi0158), .ZN(new_n11753_));
  NAND2_X1   g09317(.A1(new_n11753_), .A2(new_n11749_), .ZN(new_n11754_));
  OAI21_X1   g09318(.A1(new_n11546_), .A2(new_n11163_), .B(new_n8070_), .ZN(new_n11755_));
  NAND3_X1   g09319(.A1(new_n11754_), .A2(pi0299), .A3(new_n11755_), .ZN(new_n11756_));
  NAND2_X1   g09320(.A1(new_n11741_), .A2(new_n11756_), .ZN(new_n11757_));
  AOI21_X1   g09321(.A1(new_n11757_), .A2(pi0232), .B(new_n11716_), .ZN(new_n11758_));
  OR3_X2     g09322(.A1(new_n11758_), .A2(pi0038), .A3(new_n11708_), .Z(new_n11759_));
  NAND3_X1   g09323(.A1(new_n11759_), .A2(new_n2702_), .A3(new_n11707_), .ZN(new_n11760_));
  NOR3_X1    g09324(.A1(new_n11408_), .A2(pi0172), .A3(new_n11544_), .ZN(new_n11761_));
  NOR2_X1    g09325(.A1(new_n11376_), .A2(new_n3369_), .ZN(new_n11762_));
  NOR2_X1    g09326(.A1(new_n11407_), .A2(new_n11762_), .ZN(new_n11763_));
  NOR2_X1    g09327(.A1(new_n11763_), .A2(new_n3778_), .ZN(new_n11764_));
  NOR3_X1    g09328(.A1(new_n11761_), .A2(new_n11764_), .A3(new_n5636_), .ZN(new_n11765_));
  INV_X1     g09329(.I(new_n11407_), .ZN(new_n11766_));
  NAND2_X1   g09330(.A1(new_n11766_), .A2(new_n11448_), .ZN(new_n11767_));
  NOR3_X1    g09331(.A1(new_n11767_), .A2(pi0152), .A3(new_n11157_), .ZN(new_n11768_));
  NOR3_X1    g09332(.A1(new_n11407_), .A2(new_n3369_), .A3(new_n11222_), .ZN(new_n11769_));
  NOR3_X1    g09333(.A1(new_n11768_), .A2(pi0172), .A3(new_n11769_), .ZN(new_n11770_));
  NAND2_X1   g09334(.A1(new_n11767_), .A2(new_n3369_), .ZN(new_n11771_));
  NAND2_X1   g09335(.A1(new_n11766_), .A2(new_n11264_), .ZN(new_n11772_));
  NAND2_X1   g09336(.A1(new_n11772_), .A2(pi0152), .ZN(new_n11773_));
  AOI21_X1   g09337(.A1(new_n11771_), .A2(new_n11773_), .B(new_n3778_), .ZN(new_n11774_));
  NOR3_X1    g09338(.A1(new_n11770_), .A2(new_n11774_), .A3(pi0197), .ZN(new_n11775_));
  NOR4_X1    g09339(.A1(new_n11775_), .A2(new_n2628_), .A3(new_n8073_), .A4(new_n11765_), .ZN(new_n11776_));
  NAND2_X1   g09340(.A1(new_n11766_), .A2(new_n11281_), .ZN(new_n11777_));
  NOR2_X1    g09341(.A1(new_n11221_), .A2(new_n5398_), .ZN(new_n11778_));
  NOR2_X1    g09342(.A1(new_n11778_), .A2(new_n11164_), .ZN(new_n11779_));
  INV_X1     g09343(.I(new_n11779_), .ZN(new_n11780_));
  NOR2_X1    g09344(.A1(new_n11780_), .A2(new_n11279_), .ZN(new_n11781_));
  NOR2_X1    g09345(.A1(new_n11781_), .A2(pi0172), .ZN(new_n11782_));
  AOI21_X1   g09346(.A1(new_n11777_), .A2(pi0172), .B(new_n11782_), .ZN(new_n11783_));
  AOI21_X1   g09347(.A1(new_n11157_), .A2(new_n3778_), .B(new_n5636_), .ZN(new_n11784_));
  OAI21_X1   g09348(.A1(new_n11783_), .A2(new_n3369_), .B(new_n11784_), .ZN(new_n11785_));
  NOR2_X1    g09349(.A1(new_n11291_), .A2(new_n11407_), .ZN(new_n11786_));
  NOR2_X1    g09350(.A1(new_n11786_), .A2(pi0152), .ZN(new_n11787_));
  OAI21_X1   g09351(.A1(new_n11787_), .A2(new_n11785_), .B(new_n8066_), .ZN(new_n11788_));
  NOR2_X1    g09352(.A1(new_n11788_), .A2(new_n2628_), .ZN(new_n11789_));
  NOR2_X1    g09353(.A1(new_n11308_), .A2(new_n11407_), .ZN(new_n11790_));
  NAND2_X1   g09354(.A1(new_n11790_), .A2(pi0152), .ZN(new_n11791_));
  AOI21_X1   g09355(.A1(new_n11429_), .A2(new_n11226_), .B(new_n11407_), .ZN(new_n11792_));
  NAND2_X1   g09356(.A1(new_n11792_), .A2(new_n3369_), .ZN(new_n11793_));
  AOI21_X1   g09357(.A1(new_n11793_), .A2(new_n11791_), .B(new_n3778_), .ZN(new_n11794_));
  OAI21_X1   g09358(.A1(new_n11303_), .A2(new_n11631_), .B(new_n3778_), .ZN(new_n11795_));
  AOI21_X1   g09359(.A1(new_n11299_), .A2(new_n3369_), .B(new_n11795_), .ZN(new_n11796_));
  OAI21_X1   g09360(.A1(new_n11796_), .A2(new_n11794_), .B(new_n5636_), .ZN(new_n11797_));
  AOI21_X1   g09361(.A1(new_n11789_), .A2(new_n11797_), .B(new_n11776_), .ZN(new_n11798_));
  NAND2_X1   g09362(.A1(new_n11685_), .A2(new_n7488_), .ZN(new_n11799_));
  OAI21_X1   g09363(.A1(new_n5656_), .A2(new_n11162_), .B(new_n11799_), .ZN(new_n11800_));
  NAND3_X1   g09364(.A1(new_n11766_), .A2(new_n11158_), .A3(new_n11800_), .ZN(new_n11801_));
  NOR2_X1    g09365(.A1(new_n11407_), .A2(new_n11222_), .ZN(new_n11802_));
  NAND2_X1   g09366(.A1(new_n11802_), .A2(pi0174), .ZN(new_n11803_));
  AOI21_X1   g09367(.A1(new_n11803_), .A2(new_n11801_), .B(pi0193), .ZN(new_n11804_));
  NOR2_X1    g09368(.A1(new_n7488_), .A2(pi0145), .ZN(new_n11805_));
  AOI22_X1   g09369(.A1(new_n11264_), .A2(new_n11805_), .B1(pi0145), .B2(new_n11376_), .ZN(new_n11806_));
  NAND2_X1   g09370(.A1(new_n11806_), .A2(new_n11799_), .ZN(new_n11807_));
  AND3_X2    g09371(.A1(new_n11807_), .A2(new_n11766_), .A3(pi0193), .Z(new_n11808_));
  NOR3_X1    g09372(.A1(new_n11804_), .A2(new_n11669_), .A3(new_n11808_), .ZN(new_n11809_));
  NOR3_X1    g09373(.A1(new_n11291_), .A2(new_n5656_), .A3(new_n11407_), .ZN(new_n11810_));
  AOI21_X1   g09374(.A1(new_n11810_), .A2(new_n2744_), .B(pi0174), .ZN(new_n11811_));
  NAND3_X1   g09375(.A1(new_n11300_), .A2(new_n5656_), .A3(new_n11766_), .ZN(new_n11812_));
  INV_X1     g09376(.I(new_n11781_), .ZN(new_n11813_));
  AOI21_X1   g09377(.A1(new_n5656_), .A2(new_n11302_), .B(new_n11813_), .ZN(new_n11814_));
  OAI21_X1   g09378(.A1(new_n11814_), .A2(new_n7488_), .B(new_n7858_), .ZN(new_n11815_));
  AOI21_X1   g09379(.A1(new_n11812_), .A2(new_n11811_), .B(new_n11815_), .ZN(new_n11816_));
  INV_X1     g09380(.I(new_n11790_), .ZN(new_n11817_));
  NAND2_X1   g09381(.A1(new_n11814_), .A2(new_n9275_), .ZN(new_n11818_));
  AND3_X2    g09382(.A1(new_n11818_), .A2(pi0174), .A3(new_n11817_), .Z(new_n11819_));
  INV_X1     g09383(.I(new_n11792_), .ZN(new_n11820_));
  OAI21_X1   g09384(.A1(new_n11820_), .A2(pi0145), .B(new_n7488_), .ZN(new_n11821_));
  NOR2_X1    g09385(.A1(new_n11821_), .A2(new_n11810_), .ZN(new_n11822_));
  NOR3_X1    g09386(.A1(new_n11822_), .A2(new_n7858_), .A3(new_n11819_), .ZN(new_n11823_));
  NOR4_X1    g09387(.A1(new_n11823_), .A2(new_n11816_), .A3(pi0177), .A4(pi0299), .ZN(new_n11824_));
  OAI21_X1   g09388(.A1(new_n11824_), .A2(new_n11809_), .B(new_n3265_), .ZN(new_n11825_));
  AOI21_X1   g09389(.A1(new_n11825_), .A2(new_n11798_), .B(new_n11400_), .ZN(new_n11826_));
  OAI21_X1   g09390(.A1(new_n11826_), .A2(new_n11760_), .B(new_n11332_), .ZN(new_n11827_));
  NOR2_X1    g09391(.A1(new_n11827_), .A2(new_n11552_), .ZN(new_n11828_));
  OAI21_X1   g09392(.A1(new_n11828_), .A2(new_n11706_), .B(new_n6643_), .ZN(new_n11829_));
  NOR3_X1    g09393(.A1(new_n6698_), .A2(new_n3458_), .A3(new_n7985_), .ZN(new_n11830_));
  NOR2_X1    g09394(.A1(new_n11830_), .A2(new_n6643_), .ZN(new_n11831_));
  AOI22_X1   g09395(.A1(new_n11546_), .A2(pi0232), .B1(new_n11163_), .B2(new_n11539_), .ZN(new_n11832_));
  OAI21_X1   g09396(.A1(new_n11832_), .A2(pi0087), .B(new_n11831_), .ZN(new_n11833_));
  OAI21_X1   g09397(.A1(new_n11704_), .A2(new_n11829_), .B(new_n11833_), .ZN(po0282));
  NAND2_X1   g09398(.A1(new_n10681_), .A2(pi0087), .ZN(new_n11835_));
  INV_X1     g09399(.I(pi0126), .ZN(new_n11836_));
  NOR3_X1    g09400(.A1(pi0121), .A2(pi0125), .A3(pi0133), .ZN(new_n11837_));
  NOR2_X1    g09401(.A1(new_n11837_), .A2(new_n11836_), .ZN(new_n11838_));
  NAND2_X1   g09402(.A1(new_n11837_), .A2(new_n11836_), .ZN(new_n11839_));
  INV_X1     g09403(.I(new_n11839_), .ZN(new_n11840_));
  AOI21_X1   g09404(.A1(new_n11840_), .A2(new_n11177_), .B(new_n11838_), .ZN(new_n11841_));
  INV_X1     g09405(.I(new_n11841_), .ZN(new_n11842_));
  NOR2_X1    g09406(.A1(new_n11375_), .A2(pi0051), .ZN(new_n11843_));
  OAI21_X1   g09407(.A1(new_n11843_), .A2(new_n5666_), .B(new_n11842_), .ZN(new_n11844_));
  NAND2_X1   g09408(.A1(new_n11162_), .A2(new_n8349_), .ZN(new_n11845_));
  NOR2_X1    g09409(.A1(new_n11158_), .A2(new_n2455_), .ZN(new_n11846_));
  AOI21_X1   g09410(.A1(new_n11845_), .A2(new_n2744_), .B(new_n11846_), .ZN(new_n11847_));
  AOI21_X1   g09411(.A1(new_n5666_), .A2(new_n11171_), .B(new_n11847_), .ZN(new_n11848_));
  NAND3_X1   g09412(.A1(new_n11844_), .A2(new_n11848_), .A3(new_n3458_), .ZN(new_n11849_));
  NAND2_X1   g09413(.A1(new_n11849_), .A2(new_n11835_), .ZN(new_n11850_));
  INV_X1     g09414(.I(new_n11172_), .ZN(new_n11851_));
  OAI21_X1   g09415(.A1(new_n11376_), .A2(pi0189), .B(new_n2628_), .ZN(new_n11852_));
  AOI21_X1   g09416(.A1(pi0175), .A2(new_n11157_), .B(new_n11852_), .ZN(new_n11853_));
  NOR2_X1    g09417(.A1(new_n11843_), .A2(new_n11847_), .ZN(new_n11854_));
  OAI21_X1   g09418(.A1(new_n11854_), .A2(new_n2628_), .B(pi0232), .ZN(new_n11855_));
  NOR2_X1    g09419(.A1(new_n11853_), .A2(new_n11855_), .ZN(new_n11856_));
  NOR2_X1    g09420(.A1(new_n11856_), .A2(new_n11492_), .ZN(new_n11857_));
  NOR2_X1    g09421(.A1(new_n10672_), .A2(new_n2628_), .ZN(new_n11858_));
  INV_X1     g09422(.I(new_n11858_), .ZN(new_n11859_));
  OAI21_X1   g09423(.A1(new_n10688_), .A2(pi0299), .B(new_n11859_), .ZN(new_n11860_));
  AOI21_X1   g09424(.A1(new_n11860_), .A2(new_n6697_), .B(new_n3458_), .ZN(new_n11861_));
  OAI22_X1   g09425(.A1(new_n11857_), .A2(new_n11861_), .B1(new_n11851_), .B2(new_n11842_), .ZN(new_n11862_));
  OAI21_X1   g09426(.A1(new_n11847_), .A2(new_n7508_), .B(pi0299), .ZN(new_n11863_));
  NAND2_X1   g09427(.A1(new_n11360_), .A2(new_n3361_), .ZN(new_n11864_));
  NAND2_X1   g09428(.A1(new_n11368_), .A2(pi0166), .ZN(new_n11865_));
  AOI21_X1   g09429(.A1(new_n11864_), .A2(new_n11865_), .B(new_n2455_), .ZN(new_n11866_));
  NOR2_X1    g09430(.A1(new_n11344_), .A2(new_n8349_), .ZN(new_n11867_));
  NOR2_X1    g09431(.A1(new_n11346_), .A2(new_n8348_), .ZN(new_n11868_));
  NOR3_X1    g09432(.A1(new_n11868_), .A2(pi0153), .A3(new_n11867_), .ZN(new_n11869_));
  OAI21_X1   g09433(.A1(new_n11866_), .A2(new_n11869_), .B(new_n5635_), .ZN(new_n11870_));
  NOR2_X1    g09434(.A1(new_n11846_), .A2(new_n5635_), .ZN(new_n11871_));
  NAND2_X1   g09435(.A1(new_n11354_), .A2(pi0166), .ZN(new_n11872_));
  OAI21_X1   g09436(.A1(new_n11352_), .A2(pi0166), .B(new_n11872_), .ZN(new_n11873_));
  AOI21_X1   g09437(.A1(new_n11873_), .A2(new_n11871_), .B(new_n8070_), .ZN(new_n11874_));
  AOI21_X1   g09438(.A1(new_n11874_), .A2(new_n11870_), .B(new_n11863_), .ZN(new_n11875_));
  NAND2_X1   g09439(.A1(new_n11353_), .A2(pi0182), .ZN(new_n11876_));
  NAND3_X1   g09440(.A1(new_n11876_), .A2(new_n11710_), .A3(pi0189), .ZN(new_n11877_));
  AOI21_X1   g09441(.A1(new_n11350_), .A2(pi0182), .B(pi0189), .ZN(new_n11878_));
  NAND2_X1   g09442(.A1(new_n11722_), .A2(new_n11878_), .ZN(new_n11879_));
  AOI21_X1   g09443(.A1(new_n11879_), .A2(new_n11877_), .B(new_n9664_), .ZN(new_n11880_));
  NOR3_X1    g09444(.A1(new_n11709_), .A2(new_n9484_), .A3(new_n11157_), .ZN(new_n11881_));
  NOR2_X1    g09445(.A1(new_n11737_), .A2(pi0189), .ZN(new_n11882_));
  OAI21_X1   g09446(.A1(new_n11882_), .A2(new_n11881_), .B(new_n5659_), .ZN(new_n11883_));
  NOR3_X1    g09447(.A1(new_n11728_), .A2(new_n9484_), .A3(new_n11709_), .ZN(new_n11884_));
  NOR2_X1    g09448(.A1(new_n11733_), .A2(pi0189), .ZN(new_n11885_));
  OAI21_X1   g09449(.A1(new_n11885_), .A2(new_n11884_), .B(pi0182), .ZN(new_n11886_));
  AOI21_X1   g09450(.A1(new_n11883_), .A2(new_n11886_), .B(new_n9674_), .ZN(new_n11887_));
  NOR3_X1    g09451(.A1(new_n11875_), .A2(new_n11880_), .A3(new_n11887_), .ZN(new_n11888_));
  OAI21_X1   g09452(.A1(new_n11888_), .A2(new_n5666_), .B(new_n11715_), .ZN(new_n11889_));
  NOR2_X1    g09453(.A1(new_n11376_), .A2(new_n3361_), .ZN(new_n11890_));
  OAI21_X1   g09454(.A1(new_n11407_), .A2(new_n11890_), .B(pi0153), .ZN(new_n11891_));
  NOR3_X1    g09455(.A1(new_n11408_), .A2(pi0153), .A3(new_n11854_), .ZN(new_n11892_));
  NOR2_X1    g09456(.A1(new_n11892_), .A2(new_n10834_), .ZN(new_n11893_));
  AOI21_X1   g09457(.A1(new_n11893_), .A2(new_n11891_), .B(new_n7981_), .ZN(new_n11894_));
  NOR2_X1    g09458(.A1(new_n11158_), .A2(pi0166), .ZN(new_n11895_));
  AOI21_X1   g09459(.A1(new_n11813_), .A2(pi0166), .B(new_n11895_), .ZN(new_n11896_));
  OAI21_X1   g09460(.A1(new_n11896_), .A2(pi0153), .B(new_n10834_), .ZN(new_n11897_));
  NOR2_X1    g09461(.A1(new_n2455_), .A2(new_n3361_), .ZN(new_n11898_));
  AOI21_X1   g09462(.A1(new_n11777_), .A2(new_n11898_), .B(new_n11897_), .ZN(new_n11899_));
  OAI21_X1   g09463(.A1(pi0166), .A2(new_n11786_), .B(new_n11899_), .ZN(new_n11900_));
  NAND2_X1   g09464(.A1(new_n11900_), .A2(new_n11894_), .ZN(new_n11901_));
  NOR2_X1    g09465(.A1(new_n11281_), .A2(new_n9484_), .ZN(new_n11902_));
  NOR2_X1    g09466(.A1(new_n11290_), .A2(pi0189), .ZN(new_n11903_));
  OAI21_X1   g09467(.A1(new_n11903_), .A2(new_n11902_), .B(new_n10724_), .ZN(new_n11904_));
  NAND3_X1   g09468(.A1(new_n11234_), .A2(pi0178), .A3(new_n9530_), .ZN(new_n11905_));
  NAND4_X1   g09469(.A1(new_n11904_), .A2(pi0181), .A3(new_n11766_), .A4(new_n11905_), .ZN(new_n11906_));
  NAND2_X1   g09470(.A1(new_n11906_), .A2(new_n9542_), .ZN(new_n11907_));
  NAND2_X1   g09471(.A1(new_n11817_), .A2(pi0189), .ZN(new_n11908_));
  OAI21_X1   g09472(.A1(new_n11792_), .A2(pi0189), .B(new_n11908_), .ZN(new_n11909_));
  OAI21_X1   g09473(.A1(new_n11767_), .A2(pi0189), .B(pi0178), .ZN(new_n11910_));
  NOR2_X1    g09474(.A1(new_n11772_), .A2(new_n9484_), .ZN(new_n11911_));
  OAI21_X1   g09475(.A1(new_n11910_), .A2(new_n11911_), .B(new_n5658_), .ZN(new_n11912_));
  AOI21_X1   g09476(.A1(new_n11909_), .A2(new_n10724_), .B(new_n11912_), .ZN(new_n11913_));
  OAI21_X1   g09477(.A1(new_n11907_), .A2(new_n11913_), .B(new_n11901_), .ZN(new_n11914_));
  NAND2_X1   g09478(.A1(new_n11772_), .A2(new_n11898_), .ZN(new_n11915_));
  NOR2_X1    g09479(.A1(new_n11802_), .A2(new_n3361_), .ZN(new_n11916_));
  OAI21_X1   g09480(.A1(new_n11916_), .A2(new_n11895_), .B(new_n2455_), .ZN(new_n11917_));
  NAND2_X1   g09481(.A1(new_n11767_), .A2(new_n3361_), .ZN(new_n11918_));
  NAND4_X1   g09482(.A1(new_n11917_), .A2(pi0157), .A3(new_n11915_), .A4(new_n11918_), .ZN(new_n11919_));
  NAND2_X1   g09483(.A1(new_n11919_), .A2(new_n8033_), .ZN(new_n11920_));
  NOR2_X1    g09484(.A1(new_n11817_), .A2(new_n3361_), .ZN(new_n11921_));
  AOI21_X1   g09485(.A1(new_n11792_), .A2(new_n3361_), .B(new_n11921_), .ZN(new_n11922_));
  OAI21_X1   g09486(.A1(new_n11303_), .A2(new_n8348_), .B(new_n2455_), .ZN(new_n11923_));
  NOR2_X1    g09487(.A1(new_n11300_), .A2(pi0166), .ZN(new_n11924_));
  OAI22_X1   g09488(.A1(new_n11924_), .A2(new_n11923_), .B1(new_n2455_), .B2(new_n11922_), .ZN(new_n11925_));
  AOI21_X1   g09489(.A1(new_n11925_), .A2(new_n10834_), .B(new_n11920_), .ZN(new_n11926_));
  NOR3_X1    g09490(.A1(new_n11407_), .A2(pi0189), .A3(new_n11157_), .ZN(new_n11927_));
  NOR2_X1    g09491(.A1(new_n11927_), .A2(new_n10724_), .ZN(new_n11928_));
  INV_X1     g09492(.I(new_n11928_), .ZN(new_n11929_));
  AOI22_X1   g09493(.A1(new_n11929_), .A2(new_n11910_), .B1(pi0189), .B2(new_n11802_), .ZN(new_n11930_));
  NOR2_X1    g09494(.A1(new_n11424_), .A2(new_n8355_), .ZN(new_n11931_));
  NOR2_X1    g09495(.A1(new_n11314_), .A2(new_n8354_), .ZN(new_n11932_));
  NOR3_X1    g09496(.A1(new_n11931_), .A2(pi0178), .A3(new_n11932_), .ZN(new_n11933_));
  NOR3_X1    g09497(.A1(new_n11933_), .A2(pi0181), .A3(new_n11930_), .ZN(new_n11934_));
  OAI21_X1   g09498(.A1(new_n9484_), .A2(new_n11439_), .B(new_n11928_), .ZN(new_n11935_));
  INV_X1     g09499(.I(new_n11927_), .ZN(new_n11936_));
  AOI21_X1   g09500(.A1(new_n11781_), .A2(pi0189), .B(pi0178), .ZN(new_n11937_));
  OAI21_X1   g09501(.A1(new_n11291_), .A2(new_n11936_), .B(new_n11937_), .ZN(new_n11938_));
  AND3_X2    g09502(.A1(new_n11938_), .A2(pi0181), .A3(new_n11935_), .Z(new_n11939_));
  NOR3_X1    g09503(.A1(new_n11934_), .A2(new_n9664_), .A3(new_n11939_), .ZN(new_n11940_));
  NOR3_X1    g09504(.A1(new_n11926_), .A2(new_n11940_), .A3(new_n11914_), .ZN(new_n11941_));
  OAI21_X1   g09505(.A1(new_n11941_), .A2(new_n5666_), .B(new_n11708_), .ZN(new_n11942_));
  NAND3_X1   g09506(.A1(new_n11942_), .A2(new_n11841_), .A3(new_n11889_), .ZN(new_n11943_));
  INV_X1     g09507(.I(new_n11554_), .ZN(new_n11944_));
  NOR2_X1    g09508(.A1(new_n11585_), .A2(pi0189), .ZN(new_n11945_));
  NOR2_X1    g09509(.A1(new_n11592_), .A2(new_n9484_), .ZN(new_n11946_));
  OAI21_X1   g09510(.A1(new_n11945_), .A2(new_n11946_), .B(pi0182), .ZN(new_n11947_));
  NAND2_X1   g09511(.A1(new_n11563_), .A2(new_n9484_), .ZN(new_n11948_));
  NAND2_X1   g09512(.A1(new_n11565_), .A2(pi0189), .ZN(new_n11949_));
  AOI21_X1   g09513(.A1(new_n11948_), .A2(new_n11949_), .B(pi0182), .ZN(new_n11950_));
  NAND2_X1   g09514(.A1(new_n11950_), .A2(new_n11158_), .ZN(new_n11951_));
  AOI21_X1   g09515(.A1(new_n11951_), .A2(new_n11947_), .B(new_n9674_), .ZN(new_n11952_));
  OR2_X2     g09516(.A1(new_n11577_), .A2(new_n9484_), .Z(new_n11953_));
  INV_X1     g09517(.I(new_n11574_), .ZN(new_n11954_));
  NAND2_X1   g09518(.A1(new_n11954_), .A2(new_n9484_), .ZN(new_n11955_));
  AOI21_X1   g09519(.A1(new_n11955_), .A2(new_n11953_), .B(new_n5659_), .ZN(new_n11956_));
  OAI21_X1   g09520(.A1(new_n11956_), .A2(new_n11950_), .B(new_n9516_), .ZN(new_n11957_));
  NAND2_X1   g09521(.A1(new_n11382_), .A2(new_n3361_), .ZN(new_n11958_));
  INV_X1     g09522(.I(new_n11245_), .ZN(new_n11959_));
  NAND2_X1   g09523(.A1(new_n11959_), .A2(pi0166), .ZN(new_n11960_));
  AOI21_X1   g09524(.A1(new_n11958_), .A2(new_n11960_), .B(pi0153), .ZN(new_n11961_));
  NAND2_X1   g09525(.A1(new_n11587_), .A2(pi0166), .ZN(new_n11962_));
  NAND2_X1   g09526(.A1(new_n11606_), .A2(new_n3361_), .ZN(new_n11963_));
  AOI21_X1   g09527(.A1(new_n11963_), .A2(new_n11962_), .B(new_n2455_), .ZN(new_n11964_));
  NOR4_X1    g09528(.A1(new_n11961_), .A2(new_n5635_), .A3(new_n2614_), .A4(new_n11964_), .ZN(new_n11965_));
  NOR2_X1    g09529(.A1(new_n11590_), .A2(new_n3361_), .ZN(new_n11966_));
  NOR2_X1    g09530(.A1(new_n11581_), .A2(pi0166), .ZN(new_n11967_));
  NOR2_X1    g09531(.A1(new_n2744_), .A2(pi0153), .ZN(new_n11968_));
  NOR4_X1    g09532(.A1(new_n11967_), .A2(pi0216), .A3(new_n11966_), .A4(new_n11968_), .ZN(new_n11969_));
  OAI21_X1   g09533(.A1(new_n11965_), .A2(new_n11969_), .B(new_n5549_), .ZN(new_n11970_));
  OAI21_X1   g09534(.A1(pi0160), .A2(new_n2614_), .B(new_n5549_), .ZN(new_n11971_));
  AOI21_X1   g09535(.A1(new_n11854_), .A2(new_n11971_), .B(new_n2628_), .ZN(new_n11972_));
  NAND2_X1   g09536(.A1(new_n11970_), .A2(new_n11972_), .ZN(new_n11973_));
  NAND2_X1   g09537(.A1(new_n11957_), .A2(new_n11973_), .ZN(new_n11974_));
  OAI21_X1   g09538(.A1(new_n11974_), .A2(new_n11952_), .B(pi0232), .ZN(new_n11975_));
  AOI21_X1   g09539(.A1(new_n11975_), .A2(new_n11559_), .B(new_n11841_), .ZN(new_n11976_));
  NOR2_X1    g09540(.A1(new_n11414_), .A2(new_n9484_), .ZN(new_n11977_));
  OR3_X2     g09541(.A1(new_n11692_), .A2(pi0178), .A3(new_n11977_), .Z(new_n11978_));
  NOR2_X1    g09542(.A1(new_n11648_), .A2(new_n9484_), .ZN(new_n11979_));
  NOR2_X1    g09543(.A1(new_n11651_), .A2(pi0189), .ZN(new_n11980_));
  OAI21_X1   g09544(.A1(new_n11979_), .A2(new_n11980_), .B(pi0178), .ZN(new_n11981_));
  NOR3_X1    g09545(.A1(new_n11977_), .A2(pi0178), .A3(new_n11157_), .ZN(new_n11982_));
  NOR2_X1    g09546(.A1(new_n11691_), .A2(pi0189), .ZN(new_n11983_));
  INV_X1     g09547(.I(new_n11983_), .ZN(new_n11984_));
  AOI21_X1   g09548(.A1(new_n11984_), .A2(new_n11982_), .B(pi0181), .ZN(new_n11985_));
  NAND3_X1   g09549(.A1(new_n11981_), .A2(new_n11978_), .A3(new_n11985_), .ZN(new_n11986_));
  NAND2_X1   g09550(.A1(new_n11695_), .A2(pi0189), .ZN(new_n11987_));
  NAND2_X1   g09551(.A1(new_n11689_), .A2(new_n9484_), .ZN(new_n11988_));
  AOI21_X1   g09552(.A1(new_n11987_), .A2(new_n11988_), .B(pi0178), .ZN(new_n11989_));
  NAND2_X1   g09553(.A1(new_n11656_), .A2(pi0189), .ZN(new_n11990_));
  NAND2_X1   g09554(.A1(new_n11663_), .A2(new_n9484_), .ZN(new_n11991_));
  AOI21_X1   g09555(.A1(new_n11990_), .A2(new_n11991_), .B(new_n10724_), .ZN(new_n11992_));
  OAI21_X1   g09556(.A1(new_n11992_), .A2(new_n11989_), .B(pi0181), .ZN(new_n11993_));
  NAND3_X1   g09557(.A1(new_n11993_), .A2(new_n9516_), .A3(new_n11986_), .ZN(new_n11994_));
  NAND2_X1   g09558(.A1(new_n11659_), .A2(new_n11936_), .ZN(new_n11995_));
  AOI21_X1   g09559(.A1(new_n11663_), .A2(new_n9484_), .B(new_n10724_), .ZN(new_n11996_));
  NOR4_X1    g09560(.A1(new_n11413_), .A2(new_n9484_), .A3(new_n11157_), .A4(new_n11228_), .ZN(new_n11997_));
  NOR3_X1    g09561(.A1(new_n11689_), .A2(pi0189), .A3(new_n11157_), .ZN(new_n11998_));
  OAI21_X1   g09562(.A1(new_n11998_), .A2(new_n11997_), .B(new_n10724_), .ZN(new_n11999_));
  NAND2_X1   g09563(.A1(new_n11999_), .A2(pi0181), .ZN(new_n12000_));
  AOI21_X1   g09564(.A1(new_n11995_), .A2(new_n11996_), .B(new_n12000_), .ZN(new_n12001_));
  INV_X1     g09565(.I(new_n11985_), .ZN(new_n12002_));
  INV_X1     g09566(.I(new_n11641_), .ZN(new_n12003_));
  NAND2_X1   g09567(.A1(new_n12003_), .A2(new_n9484_), .ZN(new_n12004_));
  NAND2_X1   g09568(.A1(new_n11643_), .A2(pi0189), .ZN(new_n12005_));
  AOI21_X1   g09569(.A1(new_n12005_), .A2(new_n12004_), .B(new_n10724_), .ZN(new_n12006_));
  OAI21_X1   g09570(.A1(new_n12006_), .A2(new_n12002_), .B(new_n9542_), .ZN(new_n12007_));
  NOR2_X1    g09571(.A1(new_n12001_), .A2(new_n12007_), .ZN(new_n12008_));
  NOR2_X1    g09572(.A1(new_n11846_), .A2(pi0157), .ZN(new_n12009_));
  NOR2_X1    g09573(.A1(new_n11413_), .A2(new_n3361_), .ZN(new_n12010_));
  NOR2_X1    g09574(.A1(new_n11692_), .A2(pi0166), .ZN(new_n12011_));
  OAI21_X1   g09575(.A1(new_n12011_), .A2(new_n12010_), .B(new_n12009_), .ZN(new_n12012_));
  NAND2_X1   g09576(.A1(new_n11647_), .A2(pi0166), .ZN(new_n12013_));
  NAND2_X1   g09577(.A1(new_n11650_), .A2(new_n3361_), .ZN(new_n12014_));
  AOI21_X1   g09578(.A1(new_n12013_), .A2(new_n12014_), .B(pi0153), .ZN(new_n12015_));
  NAND2_X1   g09579(.A1(new_n12003_), .A2(new_n3361_), .ZN(new_n12016_));
  NAND2_X1   g09580(.A1(new_n11643_), .A2(pi0166), .ZN(new_n12017_));
  AOI21_X1   g09581(.A1(new_n12017_), .A2(new_n12016_), .B(new_n2455_), .ZN(new_n12018_));
  OAI21_X1   g09582(.A1(new_n12015_), .A2(new_n12018_), .B(pi0157), .ZN(new_n12019_));
  AOI21_X1   g09583(.A1(new_n12019_), .A2(new_n12012_), .B(new_n11390_), .ZN(new_n12020_));
  NOR2_X1    g09584(.A1(new_n11689_), .A2(pi0157), .ZN(new_n12021_));
  AOI21_X1   g09585(.A1(new_n11662_), .A2(pi0157), .B(new_n12021_), .ZN(new_n12022_));
  OR3_X2     g09586(.A1(new_n12022_), .A2(pi0166), .A3(new_n11846_), .Z(new_n12023_));
  NAND2_X1   g09587(.A1(new_n11625_), .A2(new_n2455_), .ZN(new_n12024_));
  NAND2_X1   g09588(.A1(new_n11627_), .A2(pi0153), .ZN(new_n12025_));
  AOI21_X1   g09589(.A1(new_n12024_), .A2(new_n12025_), .B(pi0157), .ZN(new_n12026_));
  NAND2_X1   g09590(.A1(new_n11655_), .A2(new_n2455_), .ZN(new_n12027_));
  NAND2_X1   g09591(.A1(new_n11658_), .A2(pi0153), .ZN(new_n12028_));
  AOI21_X1   g09592(.A1(new_n12027_), .A2(new_n12028_), .B(new_n10834_), .ZN(new_n12029_));
  OAI21_X1   g09593(.A1(new_n12029_), .A2(new_n12026_), .B(pi0166), .ZN(new_n12030_));
  AOI21_X1   g09594(.A1(new_n12030_), .A2(new_n12023_), .B(new_n7981_), .ZN(new_n12031_));
  NOR3_X1    g09595(.A1(new_n12031_), .A2(new_n12008_), .A3(new_n12020_), .ZN(new_n12032_));
  AOI21_X1   g09596(.A1(new_n12032_), .A2(new_n11994_), .B(new_n5666_), .ZN(new_n12033_));
  OAI21_X1   g09597(.A1(new_n12033_), .A2(new_n11944_), .B(new_n11976_), .ZN(new_n12034_));
  NAND3_X1   g09598(.A1(new_n12034_), .A2(new_n3270_), .A3(new_n11943_), .ZN(new_n12035_));
  NAND2_X1   g09599(.A1(new_n11163_), .A2(new_n3271_), .ZN(new_n12036_));
  OAI21_X1   g09600(.A1(new_n12036_), .A2(new_n11842_), .B(new_n2568_), .ZN(new_n12037_));
  AOI21_X1   g09601(.A1(new_n11856_), .A2(new_n3271_), .B(new_n12037_), .ZN(new_n12038_));
  AOI21_X1   g09602(.A1(new_n12035_), .A2(new_n12038_), .B(po1038), .ZN(new_n12039_));
  AOI22_X1   g09603(.A1(new_n12039_), .A2(new_n11862_), .B1(po1038), .B2(new_n11850_), .ZN(po0283));
  NOR2_X1    g09604(.A1(new_n8216_), .A2(new_n2577_), .ZN(new_n12041_));
  NAND2_X1   g09605(.A1(new_n9138_), .A2(new_n9129_), .ZN(new_n12042_));
  INV_X1     g09606(.I(new_n6177_), .ZN(new_n12043_));
  NOR2_X1    g09607(.A1(new_n12043_), .A2(new_n7322_), .ZN(new_n12044_));
  NAND2_X1   g09608(.A1(new_n12044_), .A2(new_n2607_), .ZN(new_n12045_));
  NOR4_X1    g09609(.A1(new_n12043_), .A2(pi0054), .A3(new_n7322_), .A4(new_n2606_), .ZN(new_n12046_));
  OAI21_X1   g09610(.A1(new_n12046_), .A2(new_n2625_), .B(new_n2602_), .ZN(new_n12047_));
  OAI21_X1   g09611(.A1(new_n5345_), .A2(new_n3265_), .B(pi0129), .ZN(new_n12048_));
  XNOR2_X1   g09612(.A1(pi0035), .A2(pi0093), .ZN(new_n12049_));
  INV_X1     g09613(.I(new_n12049_), .ZN(new_n12050_));
  INV_X1     g09614(.I(new_n2987_), .ZN(new_n12051_));
  INV_X1     g09615(.I(new_n2846_), .ZN(new_n12052_));
  NAND2_X1   g09616(.A1(new_n2966_), .A2(new_n2851_), .ZN(new_n12053_));
  AOI21_X1   g09617(.A1(new_n12053_), .A2(new_n2971_), .B(new_n2850_), .ZN(new_n12054_));
  OAI21_X1   g09618(.A1(new_n12054_), .A2(new_n2890_), .B(new_n2883_), .ZN(new_n12055_));
  NAND2_X1   g09619(.A1(new_n12055_), .A2(new_n2881_), .ZN(new_n12056_));
  NAND2_X1   g09620(.A1(new_n12056_), .A2(new_n2790_), .ZN(new_n12057_));
  AOI21_X1   g09621(.A1(new_n12057_), .A2(new_n5566_), .B(pi0086), .ZN(new_n12058_));
  NOR2_X1    g09622(.A1(new_n12058_), .A2(new_n5563_), .ZN(new_n12059_));
  OAI21_X1   g09623(.A1(new_n12059_), .A2(pi0097), .B(new_n10883_), .ZN(new_n12060_));
  NAND2_X1   g09624(.A1(new_n12060_), .A2(new_n2849_), .ZN(new_n12061_));
  NAND2_X1   g09625(.A1(new_n12061_), .A2(new_n2863_), .ZN(new_n12062_));
  NAND2_X1   g09626(.A1(new_n12062_), .A2(new_n2980_), .ZN(new_n12063_));
  AOI21_X1   g09627(.A1(new_n12063_), .A2(new_n5366_), .B(new_n3130_), .ZN(new_n12064_));
  NOR2_X1    g09628(.A1(new_n12064_), .A2(new_n12052_), .ZN(new_n12065_));
  OAI21_X1   g09629(.A1(new_n12059_), .A2(new_n2877_), .B(new_n10883_), .ZN(new_n12066_));
  NAND2_X1   g09630(.A1(new_n12066_), .A2(new_n2849_), .ZN(new_n12067_));
  NAND2_X1   g09631(.A1(new_n12067_), .A2(new_n2863_), .ZN(new_n12068_));
  NAND2_X1   g09632(.A1(new_n12068_), .A2(new_n2980_), .ZN(new_n12069_));
  AOI21_X1   g09633(.A1(new_n12069_), .A2(new_n5366_), .B(new_n3130_), .ZN(new_n12070_));
  NOR2_X1    g09634(.A1(new_n12070_), .A2(new_n12052_), .ZN(new_n12071_));
  MUX2_X1    g09635(.I0(new_n12065_), .I1(new_n12071_), .S(pi0127), .Z(new_n12072_));
  NOR2_X1    g09636(.A1(new_n10345_), .A2(new_n5327_), .ZN(new_n12073_));
  NOR2_X1    g09637(.A1(new_n12065_), .A2(new_n8241_), .ZN(new_n12074_));
  NOR2_X1    g09638(.A1(new_n12071_), .A2(po0740), .ZN(new_n12075_));
  OAI21_X1   g09639(.A1(new_n12074_), .A2(new_n12075_), .B(new_n12073_), .ZN(new_n12076_));
  OAI21_X1   g09640(.A1(new_n12072_), .A2(new_n12073_), .B(new_n12076_), .ZN(new_n12077_));
  AOI21_X1   g09641(.A1(new_n12077_), .A2(new_n2840_), .B(new_n12051_), .ZN(new_n12078_));
  AOI22_X1   g09642(.A1(new_n12078_), .A2(new_n2521_), .B1(new_n5375_), .B2(new_n12050_), .ZN(new_n12079_));
  AOI21_X1   g09643(.A1(new_n12079_), .A2(new_n2835_), .B(new_n3170_), .ZN(new_n12080_));
  OAI21_X1   g09644(.A1(new_n12080_), .A2(pi0051), .B(new_n2833_), .ZN(new_n12081_));
  AOI21_X1   g09645(.A1(new_n12081_), .A2(new_n3190_), .B(new_n2822_), .ZN(new_n12082_));
  OAI21_X1   g09646(.A1(new_n12082_), .A2(new_n2534_), .B(new_n3401_), .ZN(new_n12083_));
  AOI21_X1   g09647(.A1(new_n12083_), .A2(new_n2462_), .B(new_n3000_), .ZN(new_n12084_));
  AOI21_X1   g09648(.A1(new_n12084_), .A2(new_n2627_), .B(new_n3447_), .ZN(new_n12085_));
  AOI21_X1   g09649(.A1(new_n12085_), .A2(new_n3265_), .B(new_n12048_), .ZN(new_n12086_));
  NOR2_X1    g09650(.A1(new_n2656_), .A2(new_n3272_), .ZN(new_n12087_));
  NOR3_X1    g09651(.A1(new_n8216_), .A2(new_n2603_), .A3(new_n12087_), .ZN(new_n12088_));
  AOI21_X1   g09652(.A1(new_n12086_), .A2(new_n2603_), .B(new_n12088_), .ZN(new_n12089_));
  AOI21_X1   g09653(.A1(new_n12044_), .A2(pi0075), .B(pi0092), .ZN(new_n12090_));
  OAI21_X1   g09654(.A1(new_n12089_), .A2(pi0075), .B(new_n12090_), .ZN(new_n12091_));
  INV_X1     g09655(.I(new_n10652_), .ZN(new_n12092_));
  AOI21_X1   g09656(.A1(pi0092), .A2(new_n7322_), .B(new_n12092_), .ZN(new_n12093_));
  NOR2_X1    g09657(.A1(new_n2661_), .A2(new_n5499_), .ZN(new_n12094_));
  INV_X1     g09658(.I(new_n12094_), .ZN(new_n12095_));
  OAI21_X1   g09659(.A1(new_n8216_), .A2(new_n12095_), .B(new_n2625_), .ZN(new_n12096_));
  AOI21_X1   g09660(.A1(new_n12091_), .A2(new_n12093_), .B(new_n12096_), .ZN(new_n12097_));
  OAI22_X1   g09661(.A1(new_n12097_), .A2(new_n12047_), .B1(new_n2602_), .B2(new_n12045_), .ZN(new_n12098_));
  AOI22_X1   g09662(.A1(new_n12098_), .A2(new_n2470_), .B1(new_n12041_), .B2(new_n12042_), .ZN(new_n12099_));
  NAND4_X1   g09663(.A1(new_n12041_), .A2(new_n2470_), .A3(new_n3425_), .A4(new_n5295_), .ZN(new_n12100_));
  OAI21_X1   g09664(.A1(new_n12099_), .A2(new_n3425_), .B(new_n12100_), .ZN(po0284));
  NOR2_X1    g09665(.A1(new_n6170_), .A2(new_n5300_), .ZN(new_n12102_));
  NOR3_X1    g09666(.A1(new_n8217_), .A2(po0740), .A3(new_n8420_), .ZN(new_n12103_));
  AOI21_X1   g09667(.A1(new_n7324_), .A2(new_n8419_), .B(new_n7322_), .ZN(new_n12104_));
  OAI21_X1   g09668(.A1(new_n12103_), .A2(new_n12104_), .B(new_n7336_), .ZN(new_n12105_));
  OAI21_X1   g09669(.A1(new_n12105_), .A2(new_n2530_), .B(new_n5305_), .ZN(new_n12106_));
  AOI21_X1   g09670(.A1(new_n3453_), .A2(new_n3265_), .B(new_n5347_), .ZN(new_n12107_));
  AOI21_X1   g09671(.A1(new_n5338_), .A2(new_n5333_), .B(pi0087), .ZN(new_n12108_));
  OAI21_X1   g09672(.A1(new_n12107_), .A2(pi0100), .B(new_n12108_), .ZN(new_n12109_));
  AOI21_X1   g09673(.A1(new_n12109_), .A2(new_n5303_), .B(new_n12106_), .ZN(new_n12110_));
  NOR3_X1    g09674(.A1(new_n12110_), .A2(new_n6175_), .A3(new_n6179_), .ZN(new_n12111_));
  OAI21_X1   g09675(.A1(new_n12111_), .A2(new_n7264_), .B(new_n12102_), .ZN(new_n12112_));
  AOI21_X1   g09676(.A1(new_n12112_), .A2(new_n3284_), .B(new_n5298_), .ZN(new_n12113_));
  OAI21_X1   g09677(.A1(new_n12113_), .A2(pi0062), .B(new_n5465_), .ZN(new_n12114_));
  AOI21_X1   g09678(.A1(new_n12114_), .A2(new_n3291_), .B(new_n5296_), .ZN(po0286));
  NOR2_X1    g09679(.A1(new_n6698_), .A2(new_n4414_), .ZN(new_n12116_));
  NOR3_X1    g09680(.A1(new_n11235_), .A2(new_n12116_), .A3(pi0087), .ZN(new_n12117_));
  AOI21_X1   g09681(.A1(pi0087), .A2(new_n8089_), .B(new_n6643_), .ZN(new_n12118_));
  NAND3_X1   g09682(.A1(new_n11176_), .A2(new_n11173_), .A3(new_n11175_), .ZN(new_n12119_));
  NOR2_X1    g09683(.A1(new_n11839_), .A2(pi0132), .ZN(new_n12120_));
  NOR2_X1    g09684(.A1(new_n12120_), .A2(new_n11173_), .ZN(new_n12121_));
  NAND2_X1   g09685(.A1(new_n12120_), .A2(new_n11173_), .ZN(new_n12122_));
  INV_X1     g09686(.I(new_n12122_), .ZN(new_n12123_));
  OAI21_X1   g09687(.A1(new_n12123_), .A2(new_n12121_), .B(new_n12119_), .ZN(new_n12124_));
  AOI21_X1   g09688(.A1(new_n11375_), .A2(pi0169), .B(pi0051), .ZN(new_n12125_));
  NAND2_X1   g09689(.A1(new_n12125_), .A2(new_n3458_), .ZN(new_n12126_));
  OAI21_X1   g09690(.A1(new_n12126_), .A2(new_n12124_), .B(new_n12118_), .ZN(new_n12127_));
  NOR2_X1    g09691(.A1(new_n12127_), .A2(new_n12117_), .ZN(new_n12128_));
  NOR2_X1    g09692(.A1(new_n6698_), .A2(new_n7378_), .ZN(new_n12129_));
  NOR2_X1    g09693(.A1(new_n11235_), .A2(new_n12129_), .ZN(new_n12130_));
  NOR2_X1    g09694(.A1(new_n11843_), .A2(new_n12130_), .ZN(new_n12131_));
  OAI22_X1   g09695(.A1(new_n12131_), .A2(new_n11492_), .B1(new_n3458_), .B2(new_n7961_), .ZN(new_n12132_));
  NAND2_X1   g09696(.A1(new_n12130_), .A2(new_n8896_), .ZN(new_n12133_));
  NAND2_X1   g09697(.A1(new_n12133_), .A2(new_n2702_), .ZN(new_n12134_));
  INV_X1     g09698(.I(new_n11713_), .ZN(new_n12135_));
  AOI21_X1   g09699(.A1(new_n12135_), .A2(new_n2744_), .B(pi0232), .ZN(new_n12136_));
  NOR2_X1    g09700(.A1(new_n12136_), .A2(new_n8896_), .ZN(new_n12137_));
  NAND2_X1   g09701(.A1(new_n2628_), .A2(pi0191), .ZN(new_n12138_));
  NOR2_X1    g09702(.A1(new_n11723_), .A2(pi0051), .ZN(new_n12139_));
  NAND2_X1   g09703(.A1(new_n11251_), .A2(pi0140), .ZN(new_n12140_));
  AOI21_X1   g09704(.A1(new_n12139_), .A2(new_n12140_), .B(new_n12138_), .ZN(new_n12141_));
  INV_X1     g09705(.I(new_n7376_), .ZN(new_n12142_));
  NOR2_X1    g09706(.A1(new_n11709_), .A2(pi0051), .ZN(new_n12143_));
  INV_X1     g09707(.I(new_n12143_), .ZN(new_n12144_));
  AOI21_X1   g09708(.A1(new_n11728_), .A2(pi0140), .B(new_n12144_), .ZN(new_n12145_));
  NAND2_X1   g09709(.A1(new_n7508_), .A2(new_n7985_), .ZN(new_n12146_));
  NOR2_X1    g09710(.A1(new_n5437_), .A2(new_n4414_), .ZN(new_n12147_));
  INV_X1     g09711(.I(new_n12147_), .ZN(new_n12148_));
  NOR2_X1    g09712(.A1(new_n2530_), .A2(new_n12148_), .ZN(new_n12149_));
  AOI21_X1   g09713(.A1(new_n11241_), .A2(new_n12148_), .B(new_n12149_), .ZN(new_n12150_));
  NOR2_X1    g09714(.A1(new_n11235_), .A2(new_n7508_), .ZN(new_n12151_));
  AOI21_X1   g09715(.A1(new_n12151_), .A2(new_n12148_), .B(new_n2628_), .ZN(new_n12152_));
  OAI21_X1   g09716(.A1(new_n12150_), .A2(new_n12146_), .B(new_n12152_), .ZN(new_n12153_));
  NAND2_X1   g09717(.A1(new_n7508_), .A2(pi0162), .ZN(new_n12154_));
  NOR3_X1    g09718(.A1(new_n11349_), .A2(pi0051), .A3(new_n11251_), .ZN(new_n12155_));
  NAND2_X1   g09719(.A1(new_n12155_), .A2(pi0169), .ZN(new_n12156_));
  NAND2_X1   g09720(.A1(new_n11727_), .A2(new_n4414_), .ZN(new_n12157_));
  AOI21_X1   g09721(.A1(new_n12156_), .A2(new_n12157_), .B(new_n12154_), .ZN(new_n12158_));
  OAI22_X1   g09722(.A1(new_n12158_), .A2(new_n12153_), .B1(new_n12142_), .B2(new_n12145_), .ZN(new_n12159_));
  OAI21_X1   g09723(.A1(new_n12159_), .A2(new_n12141_), .B(pi0232), .ZN(new_n12160_));
  AOI21_X1   g09724(.A1(new_n12160_), .A2(new_n12137_), .B(new_n12134_), .ZN(new_n12161_));
  AOI21_X1   g09725(.A1(new_n12131_), .A2(pi0100), .B(new_n2569_), .ZN(new_n12162_));
  OAI21_X1   g09726(.A1(new_n2702_), .A2(new_n11171_), .B(new_n12162_), .ZN(new_n12163_));
  INV_X1     g09727(.I(new_n12124_), .ZN(new_n12164_));
  AOI21_X1   g09728(.A1(new_n12132_), .A2(new_n11851_), .B(new_n12164_), .ZN(new_n12165_));
  OAI21_X1   g09729(.A1(new_n12161_), .A2(new_n12163_), .B(new_n12165_), .ZN(new_n12166_));
  INV_X1     g09730(.I(new_n12162_), .ZN(new_n12167_));
  NAND2_X1   g09731(.A1(new_n12131_), .A2(pi0038), .ZN(new_n12168_));
  INV_X1     g09732(.I(new_n12125_), .ZN(new_n12169_));
  NAND3_X1   g09733(.A1(new_n12169_), .A2(new_n6762_), .A3(new_n12154_), .ZN(new_n12170_));
  NOR2_X1    g09734(.A1(new_n11346_), .A2(new_n12148_), .ZN(new_n12171_));
  NOR2_X1    g09735(.A1(new_n11344_), .A2(new_n12147_), .ZN(new_n12172_));
  NOR3_X1    g09736(.A1(new_n12171_), .A2(pi0216), .A3(new_n12172_), .ZN(new_n12173_));
  NOR2_X1    g09737(.A1(new_n11586_), .A2(pi0051), .ZN(new_n12174_));
  OAI21_X1   g09738(.A1(new_n2744_), .A2(new_n5398_), .B(new_n11606_), .ZN(new_n12175_));
  INV_X1     g09739(.I(new_n12175_), .ZN(new_n12176_));
  NAND2_X1   g09740(.A1(new_n12176_), .A2(pi0169), .ZN(new_n12177_));
  NAND3_X1   g09741(.A1(new_n12177_), .A2(pi0162), .A3(pi0216), .ZN(new_n12178_));
  AOI21_X1   g09742(.A1(new_n4414_), .A2(new_n12174_), .B(new_n12178_), .ZN(new_n12179_));
  OAI21_X1   g09743(.A1(new_n12179_), .A2(new_n12173_), .B(new_n5549_), .ZN(new_n12180_));
  AOI21_X1   g09744(.A1(new_n12180_), .A2(new_n12170_), .B(new_n2628_), .ZN(new_n12181_));
  AOI21_X1   g09745(.A1(new_n11588_), .A2(new_n11342_), .B(pi0051), .ZN(new_n12182_));
  INV_X1     g09746(.I(new_n12182_), .ZN(new_n12183_));
  NAND2_X1   g09747(.A1(new_n12183_), .A2(pi0140), .ZN(new_n12184_));
  AOI21_X1   g09748(.A1(new_n11342_), .A2(new_n6744_), .B(pi0051), .ZN(new_n12185_));
  INV_X1     g09749(.I(new_n12185_), .ZN(new_n12186_));
  NAND2_X1   g09750(.A1(new_n12186_), .A2(new_n7934_), .ZN(new_n12187_));
  AOI21_X1   g09751(.A1(new_n12184_), .A2(new_n12187_), .B(new_n12142_), .ZN(new_n12188_));
  AOI21_X1   g09752(.A1(new_n5437_), .A2(new_n11343_), .B(new_n11580_), .ZN(new_n12189_));
  NOR2_X1    g09753(.A1(new_n12189_), .A2(pi0224), .ZN(new_n12190_));
  AOI21_X1   g09754(.A1(pi0224), .A2(new_n12176_), .B(new_n12190_), .ZN(new_n12191_));
  NOR2_X1    g09755(.A1(new_n12191_), .A2(new_n5525_), .ZN(new_n12192_));
  AOI21_X1   g09756(.A1(new_n5525_), .A2(new_n11843_), .B(new_n12192_), .ZN(new_n12193_));
  NAND2_X1   g09757(.A1(new_n12193_), .A2(pi0140), .ZN(new_n12194_));
  NOR2_X1    g09758(.A1(new_n12189_), .A2(new_n6759_), .ZN(new_n12195_));
  AOI21_X1   g09759(.A1(new_n6759_), .A2(new_n11843_), .B(new_n12195_), .ZN(new_n12196_));
  NAND2_X1   g09760(.A1(new_n12196_), .A2(new_n7934_), .ZN(new_n12197_));
  AOI21_X1   g09761(.A1(new_n12194_), .A2(new_n12197_), .B(new_n12138_), .ZN(new_n12198_));
  NOR3_X1    g09762(.A1(new_n12198_), .A2(new_n12181_), .A3(new_n12188_), .ZN(new_n12199_));
  OAI21_X1   g09763(.A1(new_n11255_), .A2(new_n11556_), .B(new_n2744_), .ZN(new_n12200_));
  AOI21_X1   g09764(.A1(new_n12200_), .A2(new_n5666_), .B(new_n2627_), .ZN(new_n12201_));
  OAI21_X1   g09765(.A1(new_n12199_), .A2(new_n5666_), .B(new_n12201_), .ZN(new_n12202_));
  NOR2_X1    g09766(.A1(new_n11425_), .A2(new_n7377_), .ZN(new_n12203_));
  NOR2_X1    g09767(.A1(new_n11397_), .A2(new_n5437_), .ZN(new_n12204_));
  AOI21_X1   g09768(.A1(new_n11426_), .A2(new_n5437_), .B(new_n12204_), .ZN(new_n12205_));
  INV_X1     g09769(.I(new_n12205_), .ZN(new_n12206_));
  AOI21_X1   g09770(.A1(new_n12206_), .A2(new_n7377_), .B(new_n12203_), .ZN(new_n12207_));
  AOI21_X1   g09771(.A1(new_n11426_), .A2(new_n5666_), .B(pi0039), .ZN(new_n12208_));
  OAI21_X1   g09772(.A1(new_n12207_), .A2(new_n5666_), .B(new_n12208_), .ZN(new_n12209_));
  NAND3_X1   g09773(.A1(new_n12209_), .A2(new_n12202_), .A3(new_n3265_), .ZN(new_n12210_));
  AOI21_X1   g09774(.A1(new_n12210_), .A2(new_n12168_), .B(pi0100), .ZN(new_n12211_));
  OAI21_X1   g09775(.A1(new_n12211_), .A2(new_n12167_), .B(new_n12164_), .ZN(new_n12212_));
  OAI21_X1   g09776(.A1(new_n12212_), .A2(new_n12132_), .B(new_n12166_), .ZN(new_n12213_));
  AOI21_X1   g09777(.A1(new_n12213_), .A2(new_n6643_), .B(new_n12128_), .ZN(po0287));
  NOR2_X1    g09778(.A1(new_n12043_), .A2(new_n3465_), .ZN(new_n12215_));
  OR2_X2     g09779(.A1(new_n10893_), .A2(pi0100), .Z(new_n12216_));
  AOI21_X1   g09780(.A1(new_n12216_), .A2(new_n5339_), .B(new_n2565_), .ZN(new_n12217_));
  NOR3_X1    g09781(.A1(new_n12217_), .A2(pi0092), .A3(new_n12215_), .ZN(new_n12218_));
  NOR3_X1    g09782(.A1(new_n12218_), .A2(new_n7266_), .A3(new_n12092_), .ZN(po0288));
  NOR2_X1    g09783(.A1(new_n11158_), .A2(new_n10736_), .ZN(new_n12220_));
  OAI21_X1   g09784(.A1(new_n11376_), .A2(new_n10721_), .B(new_n2628_), .ZN(new_n12221_));
  NOR2_X1    g09785(.A1(new_n12221_), .A2(new_n12220_), .ZN(new_n12222_));
  NAND2_X1   g09786(.A1(new_n3533_), .A2(pi0051), .ZN(new_n12223_));
  OAI21_X1   g09787(.A1(new_n10759_), .A2(new_n11157_), .B(new_n12223_), .ZN(new_n12224_));
  NOR2_X1    g09788(.A1(new_n11165_), .A2(new_n12224_), .ZN(new_n12225_));
  NOR2_X1    g09789(.A1(new_n12225_), .A2(new_n2628_), .ZN(new_n12226_));
  INV_X1     g09790(.I(new_n12226_), .ZN(new_n12227_));
  NAND2_X1   g09791(.A1(new_n12227_), .A2(pi0232), .ZN(new_n12228_));
  NOR2_X1    g09792(.A1(new_n12228_), .A2(new_n12222_), .ZN(new_n12229_));
  INV_X1     g09793(.I(new_n12229_), .ZN(new_n12230_));
  NAND2_X1   g09794(.A1(new_n12230_), .A2(new_n3271_), .ZN(new_n12231_));
  NOR2_X1    g09795(.A1(new_n11418_), .A2(new_n5398_), .ZN(new_n12232_));
  OAI21_X1   g09796(.A1(new_n2744_), .A2(pi0173), .B(new_n5398_), .ZN(new_n12233_));
  NAND2_X1   g09797(.A1(new_n11217_), .A2(pi0182), .ZN(new_n12234_));
  AOI21_X1   g09798(.A1(new_n11404_), .A2(new_n12234_), .B(new_n12233_), .ZN(new_n12235_));
  NOR4_X1    g09799(.A1(new_n12232_), .A2(new_n10721_), .A3(pi0299), .A4(new_n12235_), .ZN(new_n12236_));
  AND2_X2    g09800(.A1(new_n11418_), .A2(new_n5437_), .Z(new_n12237_));
  NAND2_X1   g09801(.A1(new_n12223_), .A2(pi0168), .ZN(new_n12238_));
  OAI21_X1   g09802(.A1(new_n11397_), .A2(new_n12238_), .B(new_n5398_), .ZN(new_n12239_));
  NAND2_X1   g09803(.A1(new_n11431_), .A2(new_n3533_), .ZN(new_n12240_));
  OAI21_X1   g09804(.A1(new_n3533_), .A2(new_n11425_), .B(new_n12240_), .ZN(new_n12241_));
  AOI21_X1   g09805(.A1(new_n12241_), .A2(new_n4571_), .B(new_n12239_), .ZN(new_n12242_));
  NOR3_X1    g09806(.A1(new_n12242_), .A2(new_n5635_), .A3(new_n12237_), .ZN(new_n12243_));
  NAND2_X1   g09807(.A1(new_n11405_), .A2(pi0168), .ZN(new_n12244_));
  NAND2_X1   g09808(.A1(new_n12244_), .A2(new_n3533_), .ZN(new_n12245_));
  NOR2_X1    g09809(.A1(new_n11418_), .A2(new_n10759_), .ZN(new_n12246_));
  OAI21_X1   g09810(.A1(new_n12246_), .A2(new_n12245_), .B(new_n5635_), .ZN(new_n12247_));
  NOR3_X1    g09811(.A1(new_n12237_), .A2(new_n4571_), .A3(new_n11640_), .ZN(new_n12248_));
  INV_X1     g09812(.I(new_n12232_), .ZN(new_n12249_));
  AOI21_X1   g09813(.A1(new_n12249_), .A2(new_n11416_), .B(pi0168), .ZN(new_n12250_));
  NOR3_X1    g09814(.A1(new_n12250_), .A2(new_n12248_), .A3(new_n3533_), .ZN(new_n12251_));
  OAI21_X1   g09815(.A1(new_n12251_), .A2(new_n12247_), .B(pi0299), .ZN(new_n12252_));
  OAI21_X1   g09816(.A1(new_n11427_), .A2(new_n12237_), .B(pi0182), .ZN(new_n12253_));
  NAND3_X1   g09817(.A1(new_n12249_), .A2(new_n11416_), .A3(new_n5659_), .ZN(new_n12254_));
  AOI21_X1   g09818(.A1(new_n12253_), .A2(new_n12254_), .B(new_n10736_), .ZN(new_n12255_));
  AOI21_X1   g09819(.A1(new_n11432_), .A2(new_n12249_), .B(new_n5659_), .ZN(new_n12256_));
  NOR2_X1    g09820(.A1(new_n11418_), .A2(pi0182), .ZN(new_n12257_));
  NOR3_X1    g09821(.A1(new_n12256_), .A2(pi0173), .A3(new_n12257_), .ZN(new_n12258_));
  OAI21_X1   g09822(.A1(new_n12255_), .A2(new_n12258_), .B(new_n2628_), .ZN(new_n12259_));
  OAI22_X1   g09823(.A1(new_n12259_), .A2(pi0190), .B1(new_n12243_), .B2(new_n12252_), .ZN(new_n12260_));
  NOR3_X1    g09824(.A1(new_n12260_), .A2(new_n5666_), .A3(new_n12236_), .ZN(new_n12261_));
  NOR2_X1    g09825(.A1(new_n11418_), .A2(pi0232), .ZN(new_n12262_));
  OAI21_X1   g09826(.A1(new_n12261_), .A2(new_n12262_), .B(new_n2627_), .ZN(new_n12263_));
  NAND3_X1   g09827(.A1(new_n11565_), .A2(new_n7479_), .A3(new_n11158_), .ZN(new_n12264_));
  NAND2_X1   g09828(.A1(new_n11593_), .A2(pi0183), .ZN(new_n12265_));
  NAND3_X1   g09829(.A1(new_n12265_), .A2(pi0173), .A3(new_n12264_), .ZN(new_n12266_));
  NAND2_X1   g09830(.A1(new_n6759_), .A2(new_n7479_), .ZN(new_n12267_));
  NAND3_X1   g09831(.A1(new_n11577_), .A2(new_n10736_), .A3(new_n12267_), .ZN(new_n12268_));
  NAND4_X1   g09832(.A1(new_n12266_), .A2(new_n10721_), .A3(new_n2628_), .A4(new_n12268_), .ZN(new_n12269_));
  NAND2_X1   g09833(.A1(new_n11954_), .A2(pi0183), .ZN(new_n12270_));
  NAND2_X1   g09834(.A1(new_n11570_), .A2(new_n7479_), .ZN(new_n12271_));
  AOI21_X1   g09835(.A1(new_n12270_), .A2(new_n12271_), .B(pi0173), .ZN(new_n12272_));
  OAI21_X1   g09836(.A1(new_n11582_), .A2(pi0183), .B(pi0173), .ZN(new_n12273_));
  OAI22_X1   g09837(.A1(new_n12273_), .A2(new_n11585_), .B1(new_n11164_), .B2(new_n12267_), .ZN(new_n12274_));
  OAI21_X1   g09838(.A1(new_n12272_), .A2(new_n12274_), .B(new_n10722_), .ZN(new_n12275_));
  NAND2_X1   g09839(.A1(new_n12275_), .A2(new_n12269_), .ZN(new_n12276_));
  NAND2_X1   g09840(.A1(new_n11382_), .A2(pi0168), .ZN(new_n12277_));
  NAND2_X1   g09841(.A1(new_n11959_), .A2(new_n4571_), .ZN(new_n12278_));
  AOI21_X1   g09842(.A1(new_n12277_), .A2(new_n12278_), .B(pi0151), .ZN(new_n12279_));
  NAND2_X1   g09843(.A1(new_n11606_), .A2(pi0168), .ZN(new_n12280_));
  NAND2_X1   g09844(.A1(new_n11587_), .A2(new_n4571_), .ZN(new_n12281_));
  AOI21_X1   g09845(.A1(new_n12280_), .A2(new_n12281_), .B(new_n3533_), .ZN(new_n12282_));
  NOR4_X1    g09846(.A1(new_n12279_), .A2(new_n7455_), .A3(new_n2614_), .A4(new_n12282_), .ZN(new_n12283_));
  NOR2_X1    g09847(.A1(new_n11601_), .A2(new_n4571_), .ZN(new_n12284_));
  NOR2_X1    g09848(.A1(new_n11599_), .A2(pi0168), .ZN(new_n12285_));
  OAI21_X1   g09849(.A1(new_n12284_), .A2(new_n12285_), .B(new_n12223_), .ZN(new_n12286_));
  NOR2_X1    g09850(.A1(new_n12286_), .A2(pi0216), .ZN(new_n12287_));
  OAI21_X1   g09851(.A1(new_n12283_), .A2(new_n12287_), .B(new_n5549_), .ZN(new_n12288_));
  OAI21_X1   g09852(.A1(pi0149), .A2(new_n2614_), .B(new_n5549_), .ZN(new_n12289_));
  AOI21_X1   g09853(.A1(new_n12225_), .A2(new_n12289_), .B(new_n2628_), .ZN(new_n12290_));
  AOI21_X1   g09854(.A1(new_n12288_), .A2(new_n12290_), .B(new_n12276_), .ZN(new_n12291_));
  OAI21_X1   g09855(.A1(new_n12291_), .A2(new_n5666_), .B(new_n11559_), .ZN(new_n12292_));
  NAND3_X1   g09856(.A1(new_n12263_), .A2(new_n3270_), .A3(new_n12292_), .ZN(new_n12293_));
  AOI21_X1   g09857(.A1(new_n12293_), .A2(new_n12231_), .B(new_n2569_), .ZN(new_n12294_));
  NOR2_X1    g09858(.A1(new_n11840_), .A2(new_n11174_), .ZN(new_n12295_));
  AOI21_X1   g09859(.A1(new_n12119_), .A2(new_n12120_), .B(new_n12295_), .ZN(new_n12296_));
  NOR2_X1    g09860(.A1(new_n7384_), .A2(new_n3458_), .ZN(new_n12297_));
  NOR2_X1    g09861(.A1(new_n12297_), .A2(new_n12296_), .ZN(new_n12298_));
  OAI21_X1   g09862(.A1(new_n12229_), .A2(new_n11492_), .B(new_n12298_), .ZN(new_n12299_));
  OAI21_X1   g09863(.A1(new_n3458_), .A2(new_n7384_), .B(new_n12296_), .ZN(new_n12300_));
  AOI21_X1   g09864(.A1(new_n12230_), .A2(new_n11493_), .B(new_n12300_), .ZN(new_n12301_));
  NAND2_X1   g09865(.A1(new_n12230_), .A2(new_n11171_), .ZN(new_n12302_));
  AOI21_X1   g09866(.A1(new_n12302_), .A2(new_n3271_), .B(new_n2569_), .ZN(new_n12303_));
  NOR3_X1    g09867(.A1(new_n12220_), .A2(pi0190), .A3(pi0299), .ZN(new_n12304_));
  INV_X1     g09868(.I(new_n12304_), .ZN(new_n12305_));
  AOI21_X1   g09869(.A1(new_n11779_), .A2(pi0182), .B(new_n12305_), .ZN(new_n12306_));
  OAI21_X1   g09870(.A1(new_n12306_), .A2(new_n5666_), .B(new_n11302_), .ZN(new_n12307_));
  AOI21_X1   g09871(.A1(new_n11157_), .A2(new_n3533_), .B(new_n4571_), .ZN(new_n12308_));
  NAND2_X1   g09872(.A1(new_n11221_), .A2(new_n3533_), .ZN(new_n12309_));
  OAI21_X1   g09873(.A1(new_n3533_), .A2(new_n11219_), .B(new_n12309_), .ZN(new_n12310_));
  AOI22_X1   g09874(.A1(new_n12310_), .A2(new_n4571_), .B1(new_n11448_), .B2(new_n12308_), .ZN(new_n12311_));
  NOR3_X1    g09875(.A1(new_n12311_), .A2(pi0160), .A3(new_n11778_), .ZN(new_n12312_));
  INV_X1     g09876(.I(new_n11778_), .ZN(new_n12313_));
  NAND2_X1   g09877(.A1(new_n11375_), .A2(new_n4571_), .ZN(new_n12314_));
  AOI21_X1   g09878(.A1(new_n12313_), .A2(new_n12314_), .B(new_n3533_), .ZN(new_n12315_));
  INV_X1     g09879(.I(new_n12225_), .ZN(new_n12316_));
  NAND3_X1   g09880(.A1(new_n11780_), .A2(new_n3533_), .A3(new_n12316_), .ZN(new_n12317_));
  NAND2_X1   g09881(.A1(new_n12317_), .A2(pi0160), .ZN(new_n12318_));
  OAI21_X1   g09882(.A1(new_n12318_), .A2(new_n12315_), .B(pi0299), .ZN(new_n12319_));
  OAI21_X1   g09883(.A1(new_n2744_), .A2(pi0173), .B(new_n12313_), .ZN(new_n12320_));
  NOR2_X1    g09884(.A1(new_n11448_), .A2(pi0182), .ZN(new_n12321_));
  OAI21_X1   g09885(.A1(new_n12320_), .A2(new_n12321_), .B(new_n10722_), .ZN(new_n12322_));
  OAI21_X1   g09886(.A1(new_n12319_), .A2(new_n12312_), .B(new_n12322_), .ZN(new_n12323_));
  NAND2_X1   g09887(.A1(new_n12323_), .A2(pi0232), .ZN(new_n12324_));
  AOI21_X1   g09888(.A1(new_n12324_), .A2(new_n12307_), .B(pi0039), .ZN(new_n12325_));
  NAND2_X1   g09889(.A1(new_n11353_), .A2(pi0183), .ZN(new_n12326_));
  NAND3_X1   g09890(.A1(new_n12326_), .A2(new_n11710_), .A3(new_n12304_), .ZN(new_n12327_));
  NAND2_X1   g09891(.A1(new_n11350_), .A2(pi0183), .ZN(new_n12328_));
  AND3_X2    g09892(.A1(new_n11722_), .A2(new_n10736_), .A3(new_n12328_), .Z(new_n12329_));
  OR2_X2     g09893(.A1(new_n11733_), .A2(new_n7479_), .Z(new_n12330_));
  OR2_X2     g09894(.A1(new_n11737_), .A2(pi0183), .Z(new_n12331_));
  AOI21_X1   g09895(.A1(new_n12330_), .A2(new_n12331_), .B(new_n10736_), .ZN(new_n12332_));
  OAI21_X1   g09896(.A1(new_n12332_), .A2(new_n12329_), .B(new_n10722_), .ZN(new_n12333_));
  NOR2_X1    g09897(.A1(new_n12227_), .A2(new_n11163_), .ZN(new_n12334_));
  INV_X1     g09898(.I(new_n12224_), .ZN(new_n12335_));
  OAI21_X1   g09899(.A1(new_n11353_), .A2(new_n12335_), .B(new_n4571_), .ZN(new_n12336_));
  NAND2_X1   g09900(.A1(new_n12336_), .A2(pi0149), .ZN(new_n12337_));
  OAI21_X1   g09901(.A1(new_n11586_), .A2(new_n11157_), .B(new_n12223_), .ZN(new_n12338_));
  AOI21_X1   g09902(.A1(new_n11348_), .A2(new_n12338_), .B(new_n4571_), .ZN(new_n12339_));
  OAI21_X1   g09903(.A1(new_n12339_), .A2(new_n12337_), .B(new_n7508_), .ZN(new_n12340_));
  OAI21_X1   g09904(.A1(new_n11240_), .A2(new_n11157_), .B(new_n4571_), .ZN(new_n12341_));
  OAI21_X1   g09905(.A1(new_n11360_), .A2(new_n4571_), .B(new_n12341_), .ZN(new_n12342_));
  OAI21_X1   g09906(.A1(new_n11240_), .A2(new_n10759_), .B(new_n3533_), .ZN(new_n12343_));
  NOR2_X1    g09907(.A1(new_n11343_), .A2(new_n10760_), .ZN(new_n12344_));
  OAI21_X1   g09908(.A1(new_n12343_), .A2(new_n12344_), .B(new_n7455_), .ZN(new_n12345_));
  AOI21_X1   g09909(.A1(new_n12342_), .A2(pi0151), .B(new_n12345_), .ZN(new_n12346_));
  OAI22_X1   g09910(.A1(new_n12346_), .A2(new_n12340_), .B1(new_n10332_), .B2(new_n12334_), .ZN(new_n12347_));
  NAND3_X1   g09911(.A1(new_n12333_), .A2(new_n12347_), .A3(new_n12327_), .ZN(new_n12348_));
  AOI21_X1   g09912(.A1(new_n12348_), .A2(pi0232), .B(new_n11714_), .ZN(new_n12349_));
  OAI21_X1   g09913(.A1(new_n12349_), .A2(new_n2627_), .B(new_n3270_), .ZN(new_n12350_));
  OAI21_X1   g09914(.A1(new_n12350_), .A2(new_n12325_), .B(new_n12303_), .ZN(new_n12351_));
  AOI21_X1   g09915(.A1(new_n12351_), .A2(new_n12301_), .B(po1038), .ZN(new_n12352_));
  OAI21_X1   g09916(.A1(new_n12294_), .A2(new_n12299_), .B(new_n12352_), .ZN(new_n12353_));
  AOI21_X1   g09917(.A1(pi0087), .A2(new_n7360_), .B(new_n6643_), .ZN(new_n12354_));
  AND2_X2    g09918(.A1(new_n12296_), .A2(new_n11163_), .Z(new_n12355_));
  NOR2_X1    g09919(.A1(new_n12316_), .A2(new_n5666_), .ZN(new_n12356_));
  OAI21_X1   g09920(.A1(new_n12356_), .A2(new_n12355_), .B(new_n3458_), .ZN(new_n12357_));
  NAND2_X1   g09921(.A1(new_n12357_), .A2(new_n12354_), .ZN(new_n12358_));
  NAND2_X1   g09922(.A1(new_n12353_), .A2(new_n12358_), .ZN(po0289));
  OAI21_X1   g09923(.A1(new_n7547_), .A2(new_n3458_), .B(po1038), .ZN(new_n12360_));
  INV_X1     g09924(.I(pi0125), .ZN(new_n12361_));
  AOI21_X1   g09925(.A1(new_n11178_), .A2(new_n12361_), .B(pi0133), .ZN(new_n12362_));
  NOR2_X1    g09926(.A1(new_n11851_), .A2(new_n12362_), .ZN(new_n12363_));
  INV_X1     g09927(.I(new_n12362_), .ZN(new_n12364_));
  NOR3_X1    g09928(.A1(new_n3321_), .A2(new_n5666_), .A3(new_n2628_), .ZN(new_n12365_));
  OAI21_X1   g09929(.A1(new_n11451_), .A2(new_n12365_), .B(new_n7518_), .ZN(new_n12366_));
  NOR2_X1    g09930(.A1(new_n12366_), .A2(pi0039), .ZN(new_n12367_));
  OAI21_X1   g09931(.A1(new_n5398_), .A2(new_n11451_), .B(new_n11432_), .ZN(new_n12368_));
  NAND2_X1   g09932(.A1(new_n12368_), .A2(new_n12365_), .ZN(new_n12369_));
  AOI21_X1   g09933(.A1(new_n11253_), .A2(pi0145), .B(new_n6744_), .ZN(new_n12370_));
  NOR2_X1    g09934(.A1(new_n11252_), .A2(new_n5636_), .ZN(new_n12371_));
  NOR2_X1    g09935(.A1(new_n12371_), .A2(new_n5056_), .ZN(new_n12372_));
  OAI22_X1   g09936(.A1(new_n12370_), .A2(pi0299), .B1(new_n5756_), .B2(new_n12372_), .ZN(new_n12373_));
  NAND2_X1   g09937(.A1(new_n12373_), .A2(pi0232), .ZN(new_n12374_));
  NAND2_X1   g09938(.A1(new_n11557_), .A2(new_n5666_), .ZN(new_n12375_));
  AOI21_X1   g09939(.A1(new_n12374_), .A2(new_n12375_), .B(new_n2530_), .ZN(new_n12376_));
  OAI21_X1   g09940(.A1(new_n12376_), .A2(new_n2627_), .B(new_n9173_), .ZN(new_n12377_));
  AOI21_X1   g09941(.A1(new_n12369_), .A2(new_n12367_), .B(new_n12377_), .ZN(new_n12378_));
  NOR2_X1    g09942(.A1(new_n7518_), .A2(pi0039), .ZN(new_n12379_));
  NOR2_X1    g09943(.A1(new_n12368_), .A2(new_n7392_), .ZN(new_n12380_));
  NOR2_X1    g09944(.A1(new_n11450_), .A2(new_n7391_), .ZN(new_n12381_));
  OAI21_X1   g09945(.A1(new_n12380_), .A2(new_n12381_), .B(new_n12379_), .ZN(new_n12382_));
  AOI21_X1   g09946(.A1(new_n12382_), .A2(new_n12378_), .B(new_n12364_), .ZN(new_n12383_));
  NOR2_X1    g09947(.A1(new_n7479_), .A2(pi0299), .ZN(new_n12384_));
  AOI21_X1   g09948(.A1(pi0149), .A2(pi0299), .B(new_n12384_), .ZN(new_n12385_));
  NOR2_X1    g09949(.A1(new_n6698_), .A2(new_n12385_), .ZN(new_n12386_));
  OAI21_X1   g09950(.A1(new_n11278_), .A2(new_n7394_), .B(new_n11163_), .ZN(new_n12387_));
  NOR2_X1    g09951(.A1(new_n12387_), .A2(pi0039), .ZN(new_n12388_));
  NAND2_X1   g09952(.A1(new_n11353_), .A2(pi0145), .ZN(new_n12389_));
  NAND3_X1   g09953(.A1(new_n12389_), .A2(new_n11710_), .A3(new_n2628_), .ZN(new_n12390_));
  NOR3_X1    g09954(.A1(new_n11336_), .A2(new_n8070_), .A3(new_n12371_), .ZN(new_n12391_));
  OAI21_X1   g09955(.A1(new_n12391_), .A2(new_n11171_), .B(pi0299), .ZN(new_n12392_));
  AOI21_X1   g09956(.A1(new_n12390_), .A2(new_n12392_), .B(new_n5666_), .ZN(new_n12393_));
  OAI21_X1   g09957(.A1(new_n11716_), .A2(new_n12393_), .B(new_n3265_), .ZN(new_n12394_));
  AOI21_X1   g09958(.A1(new_n11171_), .A2(pi0038), .B(pi0100), .ZN(new_n12395_));
  OAI21_X1   g09959(.A1(new_n12394_), .A2(new_n12388_), .B(new_n12395_), .ZN(new_n12396_));
  AOI21_X1   g09960(.A1(new_n12396_), .A2(new_n11332_), .B(new_n11493_), .ZN(new_n12397_));
  OAI22_X1   g09961(.A1(new_n12397_), .A2(new_n12362_), .B1(new_n3458_), .B2(new_n12386_), .ZN(new_n12398_));
  AOI21_X1   g09962(.A1(new_n12383_), .A2(new_n3458_), .B(new_n12398_), .ZN(new_n12399_));
  OAI22_X1   g09963(.A1(new_n12399_), .A2(po1038), .B1(new_n12360_), .B2(new_n12363_), .ZN(po0290));
  NOR2_X1    g09964(.A1(new_n5437_), .A2(new_n3932_), .ZN(new_n12401_));
  INV_X1     g09965(.I(new_n12401_), .ZN(new_n12402_));
  NOR2_X1    g09966(.A1(new_n12402_), .A2(new_n11161_), .ZN(new_n12403_));
  NAND2_X1   g09967(.A1(new_n12403_), .A2(pi0232), .ZN(new_n12404_));
  NOR3_X1    g09968(.A1(new_n6643_), .A2(pi0051), .A3(pi0087), .ZN(new_n12405_));
  NOR2_X1    g09969(.A1(new_n12122_), .A2(pi0136), .ZN(new_n12406_));
  INV_X1     g09970(.I(new_n12406_), .ZN(new_n12407_));
  OAI21_X1   g09971(.A1(new_n12407_), .A2(pi0135), .B(pi0134), .ZN(new_n12408_));
  NAND2_X1   g09972(.A1(new_n12408_), .A2(new_n11161_), .ZN(new_n12409_));
  NAND3_X1   g09973(.A1(new_n12409_), .A2(new_n12404_), .A3(new_n12405_), .ZN(new_n12410_));
  NOR2_X1    g09974(.A1(new_n3932_), .A2(new_n2628_), .ZN(new_n12411_));
  INV_X1     g09975(.I(pi0192), .ZN(new_n12412_));
  NOR2_X1    g09976(.A1(new_n12412_), .A2(pi0299), .ZN(new_n12413_));
  NOR2_X1    g09977(.A1(new_n12411_), .A2(new_n12413_), .ZN(new_n12414_));
  NOR2_X1    g09978(.A1(new_n6698_), .A2(new_n12414_), .ZN(new_n12415_));
  NOR2_X1    g09979(.A1(new_n11235_), .A2(new_n12415_), .ZN(new_n12416_));
  NOR2_X1    g09980(.A1(new_n11843_), .A2(new_n12416_), .ZN(new_n12417_));
  NOR2_X1    g09981(.A1(new_n12417_), .A2(new_n11492_), .ZN(new_n12418_));
  AOI21_X1   g09982(.A1(new_n12417_), .A2(new_n3271_), .B(new_n2569_), .ZN(new_n12419_));
  INV_X1     g09983(.I(new_n12419_), .ZN(new_n12420_));
  NOR3_X1    g09984(.A1(new_n12206_), .A2(new_n5666_), .A3(new_n12414_), .ZN(new_n12421_));
  NOR2_X1    g09985(.A1(new_n12414_), .A2(new_n5666_), .ZN(new_n12422_));
  NOR2_X1    g09986(.A1(new_n11426_), .A2(new_n12422_), .ZN(new_n12423_));
  OAI21_X1   g09987(.A1(new_n12421_), .A2(new_n12423_), .B(new_n2627_), .ZN(new_n12424_));
  NOR2_X1    g09988(.A1(new_n2614_), .A2(pi0164), .ZN(new_n12425_));
  OAI22_X1   g09989(.A1(new_n12403_), .A2(pi0051), .B1(new_n5550_), .B2(new_n12425_), .ZN(new_n12426_));
  NOR2_X1    g09990(.A1(new_n11346_), .A2(new_n12402_), .ZN(new_n12427_));
  NOR2_X1    g09991(.A1(new_n11344_), .A2(new_n12401_), .ZN(new_n12428_));
  NOR3_X1    g09992(.A1(new_n12427_), .A2(pi0216), .A3(new_n12428_), .ZN(new_n12429_));
  NAND2_X1   g09993(.A1(new_n12176_), .A2(pi0171), .ZN(new_n12430_));
  NAND3_X1   g09994(.A1(new_n12430_), .A2(pi0164), .A3(pi0216), .ZN(new_n12431_));
  AOI21_X1   g09995(.A1(new_n3932_), .A2(new_n12174_), .B(new_n12431_), .ZN(new_n12432_));
  OAI21_X1   g09996(.A1(new_n12432_), .A2(new_n12429_), .B(new_n5549_), .ZN(new_n12433_));
  AOI21_X1   g09997(.A1(new_n12433_), .A2(new_n12426_), .B(new_n2628_), .ZN(new_n12434_));
  NOR2_X1    g09998(.A1(pi0192), .A2(pi0299), .ZN(new_n12435_));
  AOI21_X1   g09999(.A1(new_n12183_), .A2(new_n12435_), .B(new_n7381_), .ZN(new_n12436_));
  NAND2_X1   g10000(.A1(new_n12193_), .A2(new_n12413_), .ZN(new_n12437_));
  NOR2_X1    g10001(.A1(new_n2627_), .A2(new_n7381_), .ZN(new_n12438_));
  AOI21_X1   g10002(.A1(new_n12186_), .A2(new_n12435_), .B(new_n12438_), .ZN(new_n12439_));
  NAND2_X1   g10003(.A1(new_n12196_), .A2(new_n12413_), .ZN(new_n12440_));
  AOI22_X1   g10004(.A1(new_n12437_), .A2(new_n12436_), .B1(new_n12439_), .B2(new_n12440_), .ZN(new_n12441_));
  OAI21_X1   g10005(.A1(new_n12441_), .A2(new_n12434_), .B(pi0232), .ZN(new_n12442_));
  AOI21_X1   g10006(.A1(new_n12442_), .A2(new_n12201_), .B(new_n3271_), .ZN(new_n12443_));
  AOI21_X1   g10007(.A1(new_n12424_), .A2(new_n12443_), .B(new_n12420_), .ZN(new_n12444_));
  NOR3_X1    g10008(.A1(new_n12444_), .A2(new_n12408_), .A3(new_n12418_), .ZN(new_n12445_));
  NAND2_X1   g10009(.A1(new_n12419_), .A2(new_n12036_), .ZN(new_n12446_));
  NOR2_X1    g10010(.A1(new_n12416_), .A2(pi0039), .ZN(new_n12447_));
  INV_X1     g10011(.I(new_n12447_), .ZN(new_n12448_));
  NOR2_X1    g10012(.A1(new_n2627_), .A2(pi0186), .ZN(new_n12449_));
  INV_X1     g10013(.I(new_n11727_), .ZN(new_n12450_));
  NOR2_X1    g10014(.A1(new_n12450_), .A2(pi0171), .ZN(new_n12451_));
  AOI21_X1   g10015(.A1(new_n12155_), .A2(pi0171), .B(new_n12451_), .ZN(new_n12452_));
  AOI21_X1   g10016(.A1(new_n12151_), .A2(new_n12402_), .B(new_n2628_), .ZN(new_n12453_));
  OAI21_X1   g10017(.A1(new_n12452_), .A2(new_n8070_), .B(new_n12453_), .ZN(new_n12454_));
  NOR2_X1    g10018(.A1(new_n12139_), .A2(new_n12412_), .ZN(new_n12455_));
  NOR2_X1    g10019(.A1(new_n12143_), .A2(pi0192), .ZN(new_n12456_));
  OAI21_X1   g10020(.A1(new_n12455_), .A2(new_n12456_), .B(new_n2628_), .ZN(new_n12457_));
  AOI21_X1   g10021(.A1(new_n12457_), .A2(new_n12454_), .B(new_n5666_), .ZN(new_n12458_));
  OAI21_X1   g10022(.A1(new_n12458_), .A2(new_n12136_), .B(new_n12449_), .ZN(new_n12459_));
  NOR3_X1    g10023(.A1(new_n11723_), .A2(pi0051), .A3(new_n11251_), .ZN(new_n12460_));
  OAI21_X1   g10024(.A1(new_n11728_), .A2(new_n12144_), .B(new_n12412_), .ZN(new_n12461_));
  OAI21_X1   g10025(.A1(new_n12460_), .A2(new_n12412_), .B(new_n12461_), .ZN(new_n12462_));
  NAND2_X1   g10026(.A1(new_n12462_), .A2(new_n2628_), .ZN(new_n12463_));
  AOI21_X1   g10027(.A1(new_n12463_), .A2(new_n12454_), .B(new_n5666_), .ZN(new_n12464_));
  OAI21_X1   g10028(.A1(new_n12464_), .A2(new_n12136_), .B(new_n12438_), .ZN(new_n12465_));
  NAND4_X1   g10029(.A1(new_n12465_), .A2(new_n12459_), .A3(pi0164), .A4(new_n12448_), .ZN(new_n12466_));
  NAND2_X1   g10030(.A1(new_n2530_), .A2(new_n5398_), .ZN(new_n12467_));
  AOI21_X1   g10031(.A1(new_n11560_), .A2(new_n12402_), .B(new_n8070_), .ZN(new_n12468_));
  OAI21_X1   g10032(.A1(new_n3932_), .A2(new_n12467_), .B(new_n12468_), .ZN(new_n12469_));
  AND2_X2    g10033(.A1(new_n12469_), .A2(new_n12453_), .Z(new_n12470_));
  INV_X1     g10034(.I(new_n12470_), .ZN(new_n12471_));
  NAND2_X1   g10035(.A1(new_n12457_), .A2(new_n12471_), .ZN(new_n12472_));
  AOI21_X1   g10036(.A1(new_n12472_), .A2(pi0232), .B(new_n12136_), .ZN(new_n12473_));
  NOR3_X1    g10037(.A1(new_n12473_), .A2(new_n2627_), .A3(pi0186), .ZN(new_n12474_));
  NOR3_X1    g10038(.A1(new_n12474_), .A2(pi0164), .A3(new_n12447_), .ZN(new_n12475_));
  AOI21_X1   g10039(.A1(new_n12463_), .A2(new_n12471_), .B(new_n5666_), .ZN(new_n12476_));
  OAI21_X1   g10040(.A1(new_n12476_), .A2(new_n12136_), .B(new_n12438_), .ZN(new_n12477_));
  AOI21_X1   g10041(.A1(new_n12475_), .A2(new_n12477_), .B(new_n3271_), .ZN(new_n12478_));
  AOI21_X1   g10042(.A1(new_n12478_), .A2(new_n12466_), .B(new_n12446_), .ZN(new_n12479_));
  NAND2_X1   g10043(.A1(new_n12416_), .A2(new_n11199_), .ZN(new_n12480_));
  NAND2_X1   g10044(.A1(new_n12408_), .A2(new_n12480_), .ZN(new_n12481_));
  OAI21_X1   g10045(.A1(new_n12479_), .A2(new_n12481_), .B(new_n6643_), .ZN(new_n12482_));
  OAI21_X1   g10046(.A1(new_n12445_), .A2(new_n12482_), .B(new_n12410_), .ZN(po0291));
  NOR2_X1    g10047(.A1(new_n12407_), .A2(pi0135), .ZN(new_n12484_));
  INV_X1     g10048(.I(pi0135), .ZN(new_n12485_));
  NOR2_X1    g10049(.A1(new_n12406_), .A2(new_n12485_), .ZN(new_n12486_));
  AOI21_X1   g10050(.A1(new_n12484_), .A2(pi0134), .B(new_n12486_), .ZN(new_n12487_));
  NOR2_X1    g10051(.A1(new_n12487_), .A2(new_n11162_), .ZN(new_n12488_));
  AOI21_X1   g10052(.A1(new_n6697_), .A2(pi0170), .B(new_n11161_), .ZN(new_n12489_));
  OAI21_X1   g10053(.A1(new_n12488_), .A2(new_n12489_), .B(new_n12405_), .ZN(new_n12490_));
  NOR2_X1    g10054(.A1(new_n5437_), .A2(new_n4089_), .ZN(new_n12491_));
  INV_X1     g10055(.I(new_n12491_), .ZN(new_n12492_));
  NOR2_X1    g10056(.A1(new_n12492_), .A2(new_n8688_), .ZN(new_n12493_));
  INV_X1     g10057(.I(pi0194), .ZN(new_n12494_));
  NOR3_X1    g10058(.A1(new_n6698_), .A2(new_n12494_), .A3(pi0299), .ZN(new_n12495_));
  NOR3_X1    g10059(.A1(new_n12495_), .A2(new_n11235_), .A3(new_n12493_), .ZN(new_n12496_));
  NOR2_X1    g10060(.A1(new_n11843_), .A2(new_n12496_), .ZN(new_n12497_));
  AOI21_X1   g10061(.A1(new_n12497_), .A2(pi0100), .B(new_n2569_), .ZN(new_n12498_));
  NOR2_X1    g10062(.A1(new_n11235_), .A2(new_n12493_), .ZN(new_n12499_));
  AOI21_X1   g10063(.A1(new_n12499_), .A2(new_n8896_), .B(pi0194), .ZN(new_n12500_));
  AOI21_X1   g10064(.A1(new_n4089_), .A2(pi0299), .B(new_n6698_), .ZN(new_n12501_));
  NOR2_X1    g10065(.A1(new_n12501_), .A2(new_n11235_), .ZN(new_n12502_));
  AOI21_X1   g10066(.A1(new_n12502_), .A2(new_n8896_), .B(new_n12494_), .ZN(new_n12503_));
  NOR2_X1    g10067(.A1(new_n12503_), .A2(new_n12500_), .ZN(new_n12504_));
  NOR2_X1    g10068(.A1(new_n12450_), .A2(pi0170), .ZN(new_n12505_));
  AOI21_X1   g10069(.A1(new_n12155_), .A2(pi0170), .B(new_n12505_), .ZN(new_n12506_));
  OAI21_X1   g10070(.A1(new_n12506_), .A2(new_n8070_), .B(pi0150), .ZN(new_n12507_));
  NOR2_X1    g10071(.A1(new_n12467_), .A2(new_n4089_), .ZN(new_n12508_));
  OAI21_X1   g10072(.A1(new_n11241_), .A2(new_n12491_), .B(new_n7508_), .ZN(new_n12509_));
  OAI21_X1   g10073(.A1(new_n12509_), .A2(new_n12508_), .B(new_n10672_), .ZN(new_n12510_));
  AOI21_X1   g10074(.A1(new_n12507_), .A2(new_n12510_), .B(new_n2628_), .ZN(new_n12511_));
  AOI21_X1   g10075(.A1(new_n12151_), .A2(new_n12492_), .B(new_n12504_), .ZN(new_n12512_));
  OAI21_X1   g10076(.A1(new_n10688_), .A2(new_n11252_), .B(new_n12139_), .ZN(new_n12513_));
  NAND2_X1   g10077(.A1(new_n12513_), .A2(new_n12503_), .ZN(new_n12514_));
  NOR3_X1    g10078(.A1(new_n11727_), .A2(new_n10688_), .A3(new_n5437_), .ZN(new_n12515_));
  OAI21_X1   g10079(.A1(new_n12515_), .A2(new_n12144_), .B(new_n12500_), .ZN(new_n12516_));
  NAND2_X1   g10080(.A1(new_n12514_), .A2(new_n12516_), .ZN(new_n12517_));
  AOI22_X1   g10081(.A1(new_n12517_), .A2(new_n2628_), .B1(new_n12511_), .B2(new_n12512_), .ZN(new_n12518_));
  OAI22_X1   g10082(.A1(new_n12518_), .A2(new_n5666_), .B1(new_n12137_), .B2(new_n12504_), .ZN(new_n12519_));
  AOI21_X1   g10083(.A1(new_n12519_), .A2(new_n2702_), .B(new_n11331_), .ZN(new_n12520_));
  NAND2_X1   g10084(.A1(new_n12496_), .A2(new_n11199_), .ZN(new_n12521_));
  NAND2_X1   g10085(.A1(new_n12487_), .A2(new_n12521_), .ZN(new_n12522_));
  AOI21_X1   g10086(.A1(new_n12520_), .A2(new_n12498_), .B(new_n12522_), .ZN(new_n12523_));
  INV_X1     g10087(.I(new_n12487_), .ZN(new_n12524_));
  OAI21_X1   g10088(.A1(new_n11492_), .A2(new_n12497_), .B(new_n12524_), .ZN(new_n12525_));
  INV_X1     g10089(.I(new_n12498_), .ZN(new_n12526_));
  OAI21_X1   g10090(.A1(new_n11843_), .A2(new_n12502_), .B(pi0038), .ZN(new_n12527_));
  NAND2_X1   g10091(.A1(new_n12527_), .A2(pi0194), .ZN(new_n12528_));
  AOI21_X1   g10092(.A1(new_n11346_), .A2(new_n12491_), .B(new_n6762_), .ZN(new_n12529_));
  OAI21_X1   g10093(.A1(new_n11343_), .A2(new_n12491_), .B(new_n12529_), .ZN(new_n12530_));
  AOI21_X1   g10094(.A1(new_n11162_), .A2(new_n12491_), .B(pi0051), .ZN(new_n12531_));
  NAND2_X1   g10095(.A1(new_n12531_), .A2(new_n6762_), .ZN(new_n12532_));
  NAND4_X1   g10096(.A1(new_n12530_), .A2(new_n10672_), .A3(pi0299), .A4(new_n12532_), .ZN(new_n12533_));
  NAND2_X1   g10097(.A1(new_n12175_), .A2(pi0170), .ZN(new_n12534_));
  OAI21_X1   g10098(.A1(pi0170), .A2(new_n12174_), .B(new_n12534_), .ZN(new_n12535_));
  AOI22_X1   g10099(.A1(new_n12535_), .A2(pi0216), .B1(new_n8070_), .B2(new_n12530_), .ZN(new_n12536_));
  NAND2_X1   g10100(.A1(new_n12531_), .A2(new_n5550_), .ZN(new_n12537_));
  NAND2_X1   g10101(.A1(new_n12537_), .A2(new_n11858_), .ZN(new_n12538_));
  OAI21_X1   g10102(.A1(new_n12536_), .A2(new_n12538_), .B(new_n12533_), .ZN(new_n12539_));
  NAND2_X1   g10103(.A1(new_n12193_), .A2(pi0185), .ZN(new_n12540_));
  NAND2_X1   g10104(.A1(new_n12196_), .A2(new_n10688_), .ZN(new_n12541_));
  AOI21_X1   g10105(.A1(new_n12540_), .A2(new_n12541_), .B(pi0299), .ZN(new_n12542_));
  OAI21_X1   g10106(.A1(new_n12542_), .A2(new_n12539_), .B(pi0232), .ZN(new_n12543_));
  AOI21_X1   g10107(.A1(new_n11425_), .A2(new_n4089_), .B(new_n8688_), .ZN(new_n12544_));
  OAI21_X1   g10108(.A1(new_n12206_), .A2(new_n4089_), .B(new_n12544_), .ZN(new_n12545_));
  AND2_X2    g10109(.A1(new_n12545_), .A2(new_n12208_), .Z(new_n12546_));
  NAND3_X1   g10110(.A1(new_n12206_), .A2(pi0232), .A3(new_n2628_), .ZN(new_n12547_));
  AOI22_X1   g10111(.A1(new_n12546_), .A2(new_n12547_), .B1(new_n12201_), .B2(new_n12543_), .ZN(new_n12548_));
  NOR2_X1    g10112(.A1(new_n12548_), .A2(pi0038), .ZN(new_n12549_));
  OAI21_X1   g10113(.A1(new_n11843_), .A2(new_n12499_), .B(pi0038), .ZN(new_n12550_));
  NAND2_X1   g10114(.A1(new_n12550_), .A2(new_n12494_), .ZN(new_n12551_));
  NAND2_X1   g10115(.A1(new_n12186_), .A2(new_n10688_), .ZN(new_n12552_));
  OAI21_X1   g10116(.A1(new_n12182_), .A2(new_n10688_), .B(new_n12552_), .ZN(new_n12553_));
  AOI21_X1   g10117(.A1(new_n2628_), .A2(new_n12553_), .B(new_n12539_), .ZN(new_n12554_));
  OAI21_X1   g10118(.A1(new_n12554_), .A2(new_n5666_), .B(new_n12201_), .ZN(new_n12555_));
  OAI21_X1   g10119(.A1(pi0299), .A2(new_n11425_), .B(new_n12546_), .ZN(new_n12556_));
  AOI21_X1   g10120(.A1(new_n12556_), .A2(new_n12555_), .B(pi0038), .ZN(new_n12557_));
  OAI22_X1   g10121(.A1(new_n12557_), .A2(new_n12551_), .B1(new_n12549_), .B2(new_n12528_), .ZN(new_n12558_));
  AOI21_X1   g10122(.A1(new_n12558_), .A2(new_n2702_), .B(new_n12526_), .ZN(new_n12559_));
  OAI21_X1   g10123(.A1(new_n12559_), .A2(new_n12525_), .B(new_n6643_), .ZN(new_n12560_));
  OAI21_X1   g10124(.A1(new_n12560_), .A2(new_n12523_), .B(new_n12490_), .ZN(po0292));
  AOI21_X1   g10125(.A1(new_n6697_), .A2(pi0148), .B(new_n11161_), .ZN(new_n12562_));
  NOR2_X1    g10126(.A1(new_n12407_), .A2(new_n11176_), .ZN(new_n12563_));
  AOI21_X1   g10127(.A1(pi0136), .A2(new_n12122_), .B(new_n12563_), .ZN(new_n12564_));
  NOR2_X1    g10128(.A1(new_n12564_), .A2(new_n11234_), .ZN(new_n12565_));
  OAI21_X1   g10129(.A1(new_n12565_), .A2(new_n12562_), .B(new_n12405_), .ZN(new_n12566_));
  AOI21_X1   g10130(.A1(new_n7955_), .A2(new_n11162_), .B(pi0051), .ZN(new_n12567_));
  NAND2_X1   g10131(.A1(new_n12567_), .A2(new_n11199_), .ZN(new_n12568_));
  OAI21_X1   g10132(.A1(new_n11161_), .A2(new_n12568_), .B(new_n12564_), .ZN(new_n12569_));
  NAND2_X1   g10133(.A1(new_n12567_), .A2(new_n10331_), .ZN(new_n12570_));
  INV_X1     g10134(.I(new_n7952_), .ZN(new_n12571_));
  NAND2_X1   g10135(.A1(new_n11728_), .A2(pi0184), .ZN(new_n12572_));
  AOI21_X1   g10136(.A1(new_n12572_), .A2(new_n12143_), .B(new_n12571_), .ZN(new_n12573_));
  NAND2_X1   g10137(.A1(new_n2628_), .A2(pi0141), .ZN(new_n12574_));
  NAND2_X1   g10138(.A1(new_n11251_), .A2(pi0184), .ZN(new_n12575_));
  AOI21_X1   g10139(.A1(new_n12139_), .A2(new_n12575_), .B(new_n12574_), .ZN(new_n12576_));
  AOI21_X1   g10140(.A1(new_n12151_), .A2(new_n5437_), .B(new_n4257_), .ZN(new_n12577_));
  NAND2_X1   g10141(.A1(new_n7508_), .A2(new_n2744_), .ZN(new_n12578_));
  OAI21_X1   g10142(.A1(new_n11349_), .A2(new_n12578_), .B(new_n12577_), .ZN(new_n12579_));
  AOI21_X1   g10143(.A1(new_n11711_), .A2(new_n2744_), .B(pi0148), .ZN(new_n12580_));
  NOR2_X1    g10144(.A1(new_n11155_), .A2(pi0287), .ZN(new_n12581_));
  OAI22_X1   g10145(.A1(new_n12580_), .A2(new_n12581_), .B1(pi0148), .B2(new_n11235_), .ZN(new_n12582_));
  AOI21_X1   g10146(.A1(new_n12579_), .A2(new_n12582_), .B(new_n2628_), .ZN(new_n12583_));
  NOR3_X1    g10147(.A1(new_n12576_), .A2(new_n12583_), .A3(new_n12573_), .ZN(new_n12584_));
  OAI21_X1   g10148(.A1(new_n12584_), .A2(new_n5666_), .B(new_n12137_), .ZN(new_n12585_));
  OAI22_X1   g10149(.A1(new_n12585_), .A2(pi0100), .B1(new_n11161_), .B2(new_n12570_), .ZN(new_n12586_));
  AOI21_X1   g10150(.A1(new_n12586_), .A2(new_n2568_), .B(new_n12569_), .ZN(new_n12587_));
  NAND2_X1   g10151(.A1(new_n12193_), .A2(pi0184), .ZN(new_n12588_));
  NAND2_X1   g10152(.A1(new_n12196_), .A2(new_n9517_), .ZN(new_n12589_));
  AOI21_X1   g10153(.A1(new_n12588_), .A2(new_n12589_), .B(new_n12574_), .ZN(new_n12590_));
  NOR2_X1    g10154(.A1(new_n12185_), .A2(pi0184), .ZN(new_n12591_));
  AOI21_X1   g10155(.A1(new_n12183_), .A2(pi0184), .B(new_n12591_), .ZN(new_n12592_));
  NAND2_X1   g10156(.A1(new_n5549_), .A2(pi0163), .ZN(new_n12593_));
  OAI21_X1   g10157(.A1(new_n11843_), .A2(new_n6761_), .B(new_n12593_), .ZN(new_n12594_));
  OAI21_X1   g10158(.A1(new_n12175_), .A2(new_n12593_), .B(new_n12594_), .ZN(new_n12595_));
  NAND2_X1   g10159(.A1(new_n12189_), .A2(new_n6761_), .ZN(new_n12596_));
  NAND3_X1   g10160(.A1(new_n12596_), .A2(pi0148), .A3(new_n12595_), .ZN(new_n12597_));
  NOR2_X1    g10161(.A1(new_n12581_), .A2(new_n2614_), .ZN(new_n12598_));
  NOR2_X1    g10162(.A1(new_n12598_), .A2(new_n5550_), .ZN(new_n12599_));
  AOI21_X1   g10163(.A1(new_n11342_), .A2(new_n12599_), .B(pi0148), .ZN(new_n12600_));
  AOI21_X1   g10164(.A1(new_n12600_), .A2(new_n2744_), .B(new_n2628_), .ZN(new_n12601_));
  NAND2_X1   g10165(.A1(new_n12597_), .A2(new_n12601_), .ZN(new_n12602_));
  OAI21_X1   g10166(.A1(new_n12571_), .A2(new_n12592_), .B(new_n12602_), .ZN(new_n12603_));
  OAI21_X1   g10167(.A1(new_n12590_), .A2(new_n12603_), .B(pi0232), .ZN(new_n12604_));
  NAND2_X1   g10168(.A1(new_n12604_), .A2(new_n12201_), .ZN(new_n12605_));
  NOR2_X1    g10169(.A1(new_n11425_), .A2(new_n7953_), .ZN(new_n12606_));
  NOR2_X1    g10170(.A1(new_n12205_), .A2(new_n7954_), .ZN(new_n12607_));
  OAI21_X1   g10171(.A1(new_n12607_), .A2(new_n12606_), .B(pi0232), .ZN(new_n12608_));
  AOI21_X1   g10172(.A1(new_n12608_), .A2(new_n12208_), .B(new_n3271_), .ZN(new_n12609_));
  OAI21_X1   g10173(.A1(new_n12567_), .A2(new_n3270_), .B(new_n2568_), .ZN(new_n12610_));
  AOI21_X1   g10174(.A1(new_n12609_), .A2(new_n12605_), .B(new_n12610_), .ZN(new_n12611_));
  INV_X1     g10175(.I(new_n12564_), .ZN(new_n12612_));
  NAND2_X1   g10176(.A1(new_n12612_), .A2(new_n12568_), .ZN(new_n12613_));
  OAI21_X1   g10177(.A1(new_n12611_), .A2(new_n12613_), .B(new_n6643_), .ZN(new_n12614_));
  OAI21_X1   g10178(.A1(new_n12614_), .A2(new_n12587_), .B(new_n12566_), .ZN(po0293));
  NOR2_X1    g10179(.A1(new_n9316_), .A2(pi0210), .ZN(new_n12616_));
  INV_X1     g10180(.I(new_n12616_), .ZN(new_n12617_));
  NOR2_X1    g10181(.A1(po1038), .A2(pi0299), .ZN(new_n12618_));
  NAND2_X1   g10182(.A1(new_n12618_), .A2(new_n9307_), .ZN(new_n12619_));
  OAI22_X1   g10183(.A1(new_n12617_), .A2(new_n2628_), .B1(pi0198), .B2(new_n12619_), .ZN(new_n12620_));
  NAND2_X1   g10184(.A1(new_n8407_), .A2(new_n11503_), .ZN(new_n12621_));
  AOI22_X1   g10185(.A1(new_n12621_), .A2(new_n12620_), .B1(po1038), .B2(new_n12616_), .ZN(new_n12622_));
  OAI22_X1   g10186(.A1(new_n12622_), .A2(new_n7507_), .B1(pi0039), .B2(new_n3016_), .ZN(po0294));
  NOR2_X1    g10187(.A1(new_n10663_), .A2(pi0118), .ZN(new_n12624_));
  INV_X1     g10188(.I(new_n12624_), .ZN(new_n12625_));
  NOR2_X1    g10189(.A1(new_n12625_), .A2(pi0139), .ZN(new_n12626_));
  OAI21_X1   g10190(.A1(new_n10682_), .A2(new_n7905_), .B(pi0055), .ZN(new_n12627_));
  INV_X1     g10191(.I(new_n12627_), .ZN(new_n12628_));
  NAND2_X1   g10192(.A1(new_n7898_), .A2(new_n3465_), .ZN(new_n12629_));
  NOR2_X1    g10193(.A1(new_n8001_), .A2(pi0299), .ZN(new_n12630_));
  INV_X1     g10194(.I(new_n12630_), .ZN(new_n12631_));
  NAND2_X1   g10195(.A1(new_n7815_), .A2(pi0299), .ZN(new_n12632_));
  NAND3_X1   g10196(.A1(new_n12631_), .A2(new_n12632_), .A3(new_n5666_), .ZN(new_n12633_));
  NAND2_X1   g10197(.A1(new_n12633_), .A2(new_n2627_), .ZN(new_n12634_));
  INV_X1     g10198(.I(new_n12634_), .ZN(new_n12635_));
  NAND2_X1   g10199(.A1(new_n5398_), .A2(pi0148), .ZN(new_n12636_));
  AOI22_X1   g10200(.A1(new_n7815_), .A2(new_n12636_), .B1(pi0148), .B2(new_n10767_), .ZN(new_n12637_));
  INV_X1     g10201(.I(pi0141), .ZN(new_n12638_));
  AOI21_X1   g10202(.A1(new_n12630_), .A2(new_n12638_), .B(new_n5666_), .ZN(new_n12639_));
  OAI21_X1   g10203(.A1(new_n12637_), .A2(new_n2628_), .B(new_n12639_), .ZN(new_n12640_));
  INV_X1     g10204(.I(new_n10750_), .ZN(new_n12641_));
  NAND2_X1   g10205(.A1(new_n8002_), .A2(new_n5437_), .ZN(new_n12642_));
  AOI21_X1   g10206(.A1(new_n12642_), .A2(new_n12641_), .B(pi0299), .ZN(new_n12643_));
  AND2_X2    g10207(.A1(new_n12643_), .A2(pi0141), .Z(new_n12644_));
  OAI21_X1   g10208(.A1(new_n12644_), .A2(new_n12640_), .B(new_n12635_), .ZN(new_n12645_));
  NOR2_X1    g10209(.A1(new_n7627_), .A2(new_n9419_), .ZN(new_n12646_));
  NOR4_X1    g10210(.A1(new_n12646_), .A2(new_n7525_), .A3(new_n7583_), .A4(new_n7646_), .ZN(new_n12647_));
  NOR3_X1    g10211(.A1(new_n12647_), .A2(pi0299), .A3(new_n7610_), .ZN(new_n12648_));
  INV_X1     g10212(.I(new_n9419_), .ZN(new_n12649_));
  OAI21_X1   g10213(.A1(new_n6764_), .A2(new_n12649_), .B(new_n7628_), .ZN(new_n12650_));
  AOI21_X1   g10214(.A1(new_n12650_), .A2(new_n7508_), .B(new_n7637_), .ZN(new_n12651_));
  OAI21_X1   g10215(.A1(new_n12648_), .A2(new_n12651_), .B(new_n5666_), .ZN(new_n12652_));
  INV_X1     g10216(.I(new_n12652_), .ZN(new_n12653_));
  INV_X1     g10217(.I(new_n12648_), .ZN(new_n12654_));
  NAND2_X1   g10218(.A1(new_n12654_), .A2(new_n12638_), .ZN(new_n12655_));
  NAND2_X1   g10219(.A1(new_n12647_), .A2(new_n7639_), .ZN(new_n12656_));
  NAND3_X1   g10220(.A1(new_n12656_), .A2(new_n2628_), .A3(new_n7613_), .ZN(new_n12657_));
  INV_X1     g10221(.I(new_n12657_), .ZN(new_n12658_));
  OAI21_X1   g10222(.A1(new_n12638_), .A2(new_n12658_), .B(new_n12655_), .ZN(new_n12659_));
  NOR2_X1    g10223(.A1(new_n7631_), .A2(new_n12646_), .ZN(new_n12660_));
  NOR2_X1    g10224(.A1(new_n12660_), .A2(new_n7619_), .ZN(new_n12661_));
  NOR2_X1    g10225(.A1(new_n4257_), .A2(new_n2628_), .ZN(new_n12662_));
  OAI22_X1   g10226(.A1(new_n4257_), .A2(new_n12661_), .B1(new_n12651_), .B2(new_n12662_), .ZN(new_n12663_));
  AOI21_X1   g10227(.A1(new_n12659_), .A2(new_n12663_), .B(new_n5666_), .ZN(new_n12664_));
  OAI21_X1   g10228(.A1(new_n12664_), .A2(new_n12653_), .B(pi0039), .ZN(new_n12665_));
  NAND3_X1   g10229(.A1(new_n12645_), .A2(new_n3270_), .A3(new_n12665_), .ZN(new_n12666_));
  AOI21_X1   g10230(.A1(new_n12666_), .A2(new_n3458_), .B(new_n12629_), .ZN(new_n12667_));
  NAND2_X1   g10231(.A1(new_n7601_), .A2(new_n8092_), .ZN(new_n12668_));
  AOI21_X1   g10232(.A1(new_n12668_), .A2(pi0092), .B(new_n2563_), .ZN(new_n12669_));
  OAI21_X1   g10233(.A1(new_n12667_), .A2(pi0092), .B(new_n12669_), .ZN(new_n12670_));
  AOI21_X1   g10234(.A1(new_n12670_), .A2(new_n2602_), .B(new_n12628_), .ZN(new_n12671_));
  OAI21_X1   g10235(.A1(new_n12671_), .A2(new_n2471_), .B(new_n8103_), .ZN(new_n12672_));
  NOR2_X1    g10236(.A1(new_n5541_), .A2(new_n6745_), .ZN(new_n12673_));
  INV_X1     g10237(.I(new_n12673_), .ZN(new_n12674_));
  NOR2_X1    g10238(.A1(new_n12674_), .A2(new_n7525_), .ZN(new_n12675_));
  NOR2_X1    g10239(.A1(new_n12675_), .A2(new_n12574_), .ZN(new_n12676_));
  NOR3_X1    g10240(.A1(new_n5449_), .A2(new_n4257_), .A3(new_n2628_), .ZN(new_n12677_));
  OAI21_X1   g10241(.A1(new_n12676_), .A2(new_n12677_), .B(pi0232), .ZN(new_n12678_));
  INV_X1     g10242(.I(new_n9243_), .ZN(new_n12679_));
  OAI21_X1   g10243(.A1(new_n5666_), .A2(new_n12574_), .B(new_n12679_), .ZN(new_n12680_));
  NAND3_X1   g10244(.A1(new_n12680_), .A2(pi0039), .A3(new_n12678_), .ZN(new_n12681_));
  NOR2_X1    g10245(.A1(new_n7471_), .A2(new_n2536_), .ZN(new_n12682_));
  INV_X1     g10246(.I(new_n12682_), .ZN(new_n12683_));
  OR3_X2     g10247(.A1(new_n12683_), .A2(pi0039), .A3(new_n7955_), .Z(new_n12684_));
  AOI21_X1   g10248(.A1(new_n12681_), .A2(new_n12684_), .B(new_n8281_), .ZN(new_n12685_));
  NOR2_X1    g10249(.A1(new_n12685_), .A2(pi0138), .ZN(new_n12686_));
  AOI21_X1   g10250(.A1(new_n12672_), .A2(pi0138), .B(new_n12686_), .ZN(new_n12687_));
  NOR2_X1    g10251(.A1(new_n12687_), .A2(new_n12626_), .ZN(new_n12688_));
  INV_X1     g10252(.I(pi0195), .ZN(new_n12689_));
  INV_X1     g10253(.I(pi0196), .ZN(new_n12690_));
  AOI21_X1   g10254(.A1(new_n12689_), .A2(new_n12690_), .B(pi0138), .ZN(new_n12691_));
  NAND2_X1   g10255(.A1(new_n12672_), .A2(new_n12691_), .ZN(new_n12692_));
  OAI21_X1   g10256(.A1(new_n12685_), .A2(new_n12691_), .B(new_n12692_), .ZN(new_n12693_));
  AOI21_X1   g10257(.A1(new_n12693_), .A2(new_n12626_), .B(new_n12688_), .ZN(po0295));
  INV_X1     g10258(.I(new_n12669_), .ZN(new_n12695_));
  INV_X1     g10259(.I(new_n12629_), .ZN(new_n12696_));
  INV_X1     g10260(.I(new_n10767_), .ZN(new_n12697_));
  OAI22_X1   g10261(.A1(new_n12697_), .A2(new_n4414_), .B1(new_n7814_), .B2(new_n12147_), .ZN(new_n12698_));
  OAI21_X1   g10262(.A1(new_n12631_), .A2(pi0191), .B(pi0232), .ZN(new_n12699_));
  AOI21_X1   g10263(.A1(new_n12698_), .A2(pi0299), .B(new_n12699_), .ZN(new_n12700_));
  NAND2_X1   g10264(.A1(new_n12643_), .A2(pi0191), .ZN(new_n12701_));
  AOI21_X1   g10265(.A1(new_n12700_), .A2(new_n12701_), .B(new_n12634_), .ZN(new_n12702_));
  NOR2_X1    g10266(.A1(new_n12648_), .A2(pi0191), .ZN(new_n12703_));
  INV_X1     g10267(.I(pi0191), .ZN(new_n12704_));
  NOR2_X1    g10268(.A1(new_n12658_), .A2(new_n12704_), .ZN(new_n12705_));
  AOI21_X1   g10269(.A1(new_n4414_), .A2(new_n7627_), .B(new_n12660_), .ZN(new_n12706_));
  NOR2_X1    g10270(.A1(new_n12706_), .A2(new_n8070_), .ZN(new_n12707_));
  OAI22_X1   g10271(.A1(new_n12705_), .A2(new_n12703_), .B1(new_n7637_), .B2(new_n12707_), .ZN(new_n12708_));
  AOI21_X1   g10272(.A1(new_n12708_), .A2(pi0232), .B(new_n12653_), .ZN(new_n12709_));
  OAI21_X1   g10273(.A1(new_n12709_), .A2(new_n2627_), .B(new_n3270_), .ZN(new_n12710_));
  OAI21_X1   g10274(.A1(new_n12702_), .A2(new_n12710_), .B(new_n3458_), .ZN(new_n12711_));
  AOI21_X1   g10275(.A1(new_n12711_), .A2(new_n12696_), .B(pi0092), .ZN(new_n12712_));
  OAI21_X1   g10276(.A1(new_n12712_), .A2(new_n12695_), .B(new_n2602_), .ZN(new_n12713_));
  NAND2_X1   g10277(.A1(new_n12713_), .A2(new_n12627_), .ZN(new_n12714_));
  NAND2_X1   g10278(.A1(new_n12714_), .A2(new_n2470_), .ZN(new_n12715_));
  NAND2_X1   g10279(.A1(new_n12715_), .A2(new_n8103_), .ZN(new_n12716_));
  NAND2_X1   g10280(.A1(new_n12716_), .A2(pi0139), .ZN(new_n12717_));
  INV_X1     g10281(.I(pi0139), .ZN(new_n12718_));
  NOR2_X1    g10282(.A1(new_n12679_), .A2(pi0232), .ZN(new_n12719_));
  INV_X1     g10283(.I(new_n12719_), .ZN(new_n12720_));
  INV_X1     g10284(.I(new_n9240_), .ZN(new_n12721_));
  NAND3_X1   g10285(.A1(new_n6745_), .A2(pi0169), .A3(pi0299), .ZN(new_n12722_));
  NOR2_X1    g10286(.A1(new_n9241_), .A2(pi0191), .ZN(new_n12723_));
  NOR2_X1    g10287(.A1(new_n12675_), .A2(new_n12704_), .ZN(new_n12724_));
  OAI21_X1   g10288(.A1(new_n12724_), .A2(new_n12723_), .B(new_n2628_), .ZN(new_n12725_));
  NAND4_X1   g10289(.A1(new_n12725_), .A2(pi0232), .A3(new_n12721_), .A4(new_n12722_), .ZN(new_n12726_));
  AOI21_X1   g10290(.A1(new_n12726_), .A2(new_n12720_), .B(new_n2627_), .ZN(new_n12727_));
  NOR3_X1    g10291(.A1(new_n12683_), .A2(pi0039), .A3(new_n12129_), .ZN(new_n12728_));
  OAI21_X1   g10292(.A1(new_n12727_), .A2(new_n12728_), .B(new_n8280_), .ZN(new_n12729_));
  NAND2_X1   g10293(.A1(new_n12729_), .A2(new_n12718_), .ZN(new_n12730_));
  AOI21_X1   g10294(.A1(new_n12717_), .A2(new_n12730_), .B(new_n12624_), .ZN(new_n12731_));
  NOR3_X1    g10295(.A1(pi0138), .A2(pi0195), .A3(pi0196), .ZN(new_n12732_));
  NOR2_X1    g10296(.A1(new_n12732_), .A2(pi0139), .ZN(new_n12733_));
  NAND2_X1   g10297(.A1(new_n12716_), .A2(new_n12733_), .ZN(new_n12734_));
  OAI21_X1   g10298(.A1(pi0139), .A2(new_n12732_), .B(new_n12729_), .ZN(new_n12735_));
  AOI21_X1   g10299(.A1(new_n12734_), .A2(new_n12735_), .B(new_n12625_), .ZN(new_n12736_));
  NOR2_X1    g10300(.A1(new_n12731_), .A2(new_n12736_), .ZN(po0296));
  INV_X1     g10301(.I(pi0832), .ZN(new_n12738_));
  INV_X1     g10302(.I(pi1160), .ZN(new_n12739_));
  INV_X1     g10303(.I(pi0715), .ZN(new_n12740_));
  INV_X1     g10304(.I(pi0647), .ZN(new_n12741_));
  INV_X1     g10305(.I(pi1156), .ZN(new_n12742_));
  NOR2_X1    g10306(.A1(new_n3042_), .A2(pi0140), .ZN(new_n12743_));
  INV_X1     g10307(.I(new_n12743_), .ZN(new_n12744_));
  INV_X1     g10308(.I(pi1158), .ZN(new_n12745_));
  NOR2_X1    g10309(.A1(new_n12745_), .A2(pi0626), .ZN(new_n12746_));
  INV_X1     g10310(.I(pi0626), .ZN(new_n12747_));
  NOR2_X1    g10311(.A1(new_n12747_), .A2(pi1158), .ZN(new_n12748_));
  NOR2_X1    g10312(.A1(new_n12746_), .A2(new_n12748_), .ZN(new_n12749_));
  INV_X1     g10313(.I(pi0761), .ZN(new_n12750_));
  INV_X1     g10314(.I(pi0603), .ZN(new_n12751_));
  INV_X1     g10315(.I(pi0621), .ZN(new_n12752_));
  NOR2_X1    g10316(.A1(new_n12752_), .A2(new_n3022_), .ZN(new_n12753_));
  NOR2_X1    g10317(.A1(new_n12753_), .A2(new_n12751_), .ZN(new_n12754_));
  INV_X1     g10318(.I(new_n12754_), .ZN(new_n12755_));
  NOR2_X1    g10319(.A1(new_n12755_), .A2(new_n3043_), .ZN(new_n12756_));
  AOI21_X1   g10320(.A1(new_n12756_), .A2(new_n12750_), .B(new_n12743_), .ZN(new_n12757_));
  INV_X1     g10321(.I(pi0778), .ZN(new_n12758_));
  XNOR2_X1   g10322(.A1(pi0608), .A2(pi1153), .ZN(new_n12759_));
  NOR2_X1    g10323(.A1(new_n12759_), .A2(new_n12758_), .ZN(new_n12760_));
  INV_X1     g10324(.I(new_n12760_), .ZN(new_n12761_));
  NOR2_X1    g10325(.A1(new_n12761_), .A2(new_n3043_), .ZN(new_n12762_));
  NOR3_X1    g10326(.A1(new_n12757_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n12763_));
  INV_X1     g10327(.I(pi0785), .ZN(new_n12764_));
  NOR2_X1    g10328(.A1(new_n12757_), .A2(new_n12762_), .ZN(new_n12765_));
  INV_X1     g10329(.I(pi0609), .ZN(new_n12766_));
  NOR2_X1    g10330(.A1(new_n3043_), .A2(new_n12766_), .ZN(new_n12767_));
  INV_X1     g10331(.I(new_n12767_), .ZN(new_n12768_));
  AOI21_X1   g10332(.A1(new_n12765_), .A2(new_n12768_), .B(pi1155), .ZN(new_n12769_));
  INV_X1     g10333(.I(pi1155), .ZN(new_n12770_));
  INV_X1     g10334(.I(new_n12757_), .ZN(new_n12771_));
  NOR2_X1    g10335(.A1(new_n12760_), .A2(new_n12766_), .ZN(new_n12772_));
  NOR2_X1    g10336(.A1(new_n12772_), .A2(new_n3043_), .ZN(new_n12773_));
  INV_X1     g10337(.I(new_n12773_), .ZN(new_n12774_));
  AOI21_X1   g10338(.A1(new_n12771_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n12775_));
  NOR3_X1    g10339(.A1(new_n12769_), .A2(new_n12775_), .A3(new_n12764_), .ZN(new_n12776_));
  NOR2_X1    g10340(.A1(new_n12776_), .A2(new_n12763_), .ZN(new_n12777_));
  NOR2_X1    g10341(.A1(new_n12777_), .A2(pi0781), .ZN(new_n12778_));
  INV_X1     g10342(.I(pi0781), .ZN(new_n12779_));
  INV_X1     g10343(.I(new_n12777_), .ZN(new_n12780_));
  INV_X1     g10344(.I(pi0618), .ZN(new_n12781_));
  NOR2_X1    g10345(.A1(new_n3043_), .A2(new_n12781_), .ZN(new_n12782_));
  INV_X1     g10346(.I(new_n12782_), .ZN(new_n12783_));
  AOI21_X1   g10347(.A1(new_n12780_), .A2(new_n12783_), .B(pi1154), .ZN(new_n12784_));
  INV_X1     g10348(.I(pi1154), .ZN(new_n12785_));
  NOR2_X1    g10349(.A1(new_n3043_), .A2(pi0618), .ZN(new_n12786_));
  INV_X1     g10350(.I(new_n12786_), .ZN(new_n12787_));
  AOI21_X1   g10351(.A1(new_n12780_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n12788_));
  NOR3_X1    g10352(.A1(new_n12784_), .A2(new_n12788_), .A3(new_n12779_), .ZN(new_n12789_));
  NOR2_X1    g10353(.A1(new_n12789_), .A2(new_n12778_), .ZN(new_n12790_));
  INV_X1     g10354(.I(pi1159), .ZN(new_n12791_));
  NOR3_X1    g10355(.A1(new_n12789_), .A2(pi0619), .A3(new_n12778_), .ZN(new_n12792_));
  INV_X1     g10356(.I(pi0619), .ZN(new_n12793_));
  NOR2_X1    g10357(.A1(new_n12743_), .A2(new_n12793_), .ZN(new_n12794_));
  OAI21_X1   g10358(.A1(new_n12792_), .A2(new_n12794_), .B(new_n12791_), .ZN(new_n12795_));
  INV_X1     g10359(.I(pi0789), .ZN(new_n12796_));
  NAND2_X1   g10360(.A1(new_n12790_), .A2(pi0619), .ZN(new_n12797_));
  NAND2_X1   g10361(.A1(new_n12744_), .A2(new_n12793_), .ZN(new_n12798_));
  AOI21_X1   g10362(.A1(new_n12797_), .A2(new_n12798_), .B(new_n12791_), .ZN(new_n12799_));
  NOR2_X1    g10363(.A1(new_n12799_), .A2(new_n12796_), .ZN(new_n12800_));
  NAND2_X1   g10364(.A1(new_n12800_), .A2(new_n12795_), .ZN(new_n12801_));
  OAI21_X1   g10365(.A1(pi0789), .A2(new_n12790_), .B(new_n12801_), .ZN(new_n12802_));
  XOR2_X1    g10366(.A1(pi0626), .A2(pi1158), .Z(new_n12803_));
  INV_X1     g10367(.I(new_n12803_), .ZN(new_n12804_));
  NAND2_X1   g10368(.A1(new_n12802_), .A2(new_n12804_), .ZN(new_n12805_));
  OAI21_X1   g10369(.A1(new_n12744_), .A2(new_n12749_), .B(new_n12805_), .ZN(new_n12806_));
  NAND2_X1   g10370(.A1(new_n12806_), .A2(pi0788), .ZN(new_n12807_));
  INV_X1     g10371(.I(pi0788), .ZN(new_n12808_));
  NAND2_X1   g10372(.A1(new_n12802_), .A2(new_n12808_), .ZN(new_n12809_));
  NAND2_X1   g10373(.A1(new_n12807_), .A2(new_n12809_), .ZN(new_n12810_));
  NOR2_X1    g10374(.A1(new_n12810_), .A2(pi0628), .ZN(new_n12811_));
  NOR2_X1    g10375(.A1(new_n12745_), .A2(pi0641), .ZN(new_n12812_));
  INV_X1     g10376(.I(new_n12812_), .ZN(new_n12813_));
  INV_X1     g10377(.I(pi0641), .ZN(new_n12814_));
  NOR2_X1    g10378(.A1(new_n12814_), .A2(pi1158), .ZN(new_n12815_));
  INV_X1     g10379(.I(new_n12815_), .ZN(new_n12816_));
  AOI21_X1   g10380(.A1(new_n12813_), .A2(new_n12816_), .B(new_n12808_), .ZN(new_n12817_));
  NOR2_X1    g10381(.A1(new_n12749_), .A2(new_n12808_), .ZN(new_n12818_));
  NOR2_X1    g10382(.A1(new_n12818_), .A2(new_n12817_), .ZN(new_n12819_));
  INV_X1     g10383(.I(pi0738), .ZN(new_n12820_));
  INV_X1     g10384(.I(pi0680), .ZN(new_n12821_));
  INV_X1     g10385(.I(pi0665), .ZN(new_n12822_));
  NOR2_X1    g10386(.A1(new_n12822_), .A2(new_n3022_), .ZN(new_n12823_));
  NOR2_X1    g10387(.A1(new_n12823_), .A2(new_n12821_), .ZN(new_n12824_));
  INV_X1     g10388(.I(new_n12824_), .ZN(new_n12825_));
  NOR2_X1    g10389(.A1(new_n12825_), .A2(new_n3043_), .ZN(new_n12826_));
  AOI21_X1   g10390(.A1(new_n12826_), .A2(new_n12820_), .B(new_n12743_), .ZN(new_n12827_));
  NOR2_X1    g10391(.A1(new_n12827_), .A2(new_n12754_), .ZN(new_n12828_));
  NOR2_X1    g10392(.A1(new_n12828_), .A2(new_n12771_), .ZN(new_n12829_));
  NAND2_X1   g10393(.A1(new_n12829_), .A2(new_n12758_), .ZN(new_n12830_));
  NOR2_X1    g10394(.A1(new_n12743_), .A2(pi1153), .ZN(new_n12831_));
  INV_X1     g10395(.I(new_n12826_), .ZN(new_n12832_));
  NOR2_X1    g10396(.A1(new_n12832_), .A2(pi0625), .ZN(new_n12833_));
  INV_X1     g10397(.I(new_n12833_), .ZN(new_n12834_));
  NOR2_X1    g10398(.A1(new_n12834_), .A2(pi0738), .ZN(new_n12835_));
  INV_X1     g10399(.I(new_n12835_), .ZN(new_n12836_));
  NAND2_X1   g10400(.A1(new_n12836_), .A2(new_n12831_), .ZN(new_n12837_));
  NAND2_X1   g10401(.A1(new_n12828_), .A2(pi0625), .ZN(new_n12838_));
  NAND3_X1   g10402(.A1(new_n12838_), .A2(pi1153), .A3(new_n12757_), .ZN(new_n12839_));
  AND3_X2    g10403(.A1(new_n12837_), .A2(pi0608), .A3(new_n12839_), .Z(new_n12840_));
  INV_X1     g10404(.I(pi1153), .ZN(new_n12841_));
  NOR2_X1    g10405(.A1(new_n12835_), .A2(new_n12827_), .ZN(new_n12842_));
  NOR2_X1    g10406(.A1(new_n12842_), .A2(new_n12841_), .ZN(new_n12843_));
  NOR2_X1    g10407(.A1(new_n12843_), .A2(pi0608), .ZN(new_n12844_));
  INV_X1     g10408(.I(new_n12838_), .ZN(new_n12845_));
  OAI21_X1   g10409(.A1(new_n12845_), .A2(new_n12829_), .B(new_n12831_), .ZN(new_n12846_));
  NAND2_X1   g10410(.A1(new_n12844_), .A2(new_n12846_), .ZN(new_n12847_));
  NAND2_X1   g10411(.A1(new_n12847_), .A2(pi0778), .ZN(new_n12848_));
  OAI21_X1   g10412(.A1(new_n12848_), .A2(new_n12840_), .B(new_n12830_), .ZN(new_n12849_));
  INV_X1     g10413(.I(new_n12849_), .ZN(new_n12850_));
  NOR2_X1    g10414(.A1(new_n12827_), .A2(pi0778), .ZN(new_n12851_));
  INV_X1     g10415(.I(new_n12837_), .ZN(new_n12852_));
  NOR3_X1    g10416(.A1(new_n12852_), .A2(new_n12758_), .A3(new_n12843_), .ZN(new_n12853_));
  NOR2_X1    g10417(.A1(new_n12853_), .A2(new_n12851_), .ZN(new_n12854_));
  INV_X1     g10418(.I(new_n12854_), .ZN(new_n12855_));
  NOR2_X1    g10419(.A1(new_n12855_), .A2(pi0609), .ZN(new_n12856_));
  AOI21_X1   g10420(.A1(new_n12849_), .A2(pi0609), .B(new_n12856_), .ZN(new_n12857_));
  NOR2_X1    g10421(.A1(new_n12857_), .A2(new_n12770_), .ZN(new_n12858_));
  NOR2_X1    g10422(.A1(new_n12858_), .A2(new_n12769_), .ZN(new_n12859_));
  NOR2_X1    g10423(.A1(new_n12850_), .A2(pi0609), .ZN(new_n12860_));
  NOR2_X1    g10424(.A1(new_n12855_), .A2(new_n12766_), .ZN(new_n12861_));
  OAI21_X1   g10425(.A1(new_n12860_), .A2(new_n12861_), .B(new_n12770_), .ZN(new_n12862_));
  NOR2_X1    g10426(.A1(new_n12775_), .A2(pi0660), .ZN(new_n12863_));
  AOI22_X1   g10427(.A1(new_n12859_), .A2(pi0660), .B1(new_n12862_), .B2(new_n12863_), .ZN(new_n12864_));
  NAND2_X1   g10428(.A1(new_n12864_), .A2(pi0785), .ZN(new_n12865_));
  OAI21_X1   g10429(.A1(pi0785), .A2(new_n12850_), .B(new_n12865_), .ZN(new_n12866_));
  INV_X1     g10430(.I(new_n12788_), .ZN(new_n12867_));
  XNOR2_X1   g10431(.A1(pi0660), .A2(pi1155), .ZN(new_n12868_));
  NOR2_X1    g10432(.A1(new_n12868_), .A2(new_n12764_), .ZN(new_n12869_));
  INV_X1     g10433(.I(new_n12869_), .ZN(new_n12870_));
  NOR2_X1    g10434(.A1(new_n12870_), .A2(new_n3043_), .ZN(new_n12871_));
  NOR2_X1    g10435(.A1(new_n12854_), .A2(new_n12871_), .ZN(new_n12872_));
  NOR2_X1    g10436(.A1(new_n12872_), .A2(new_n12781_), .ZN(new_n12873_));
  AOI21_X1   g10437(.A1(new_n12866_), .A2(new_n12781_), .B(new_n12873_), .ZN(new_n12874_));
  OAI21_X1   g10438(.A1(new_n12874_), .A2(pi1154), .B(new_n12867_), .ZN(new_n12875_));
  INV_X1     g10439(.I(new_n12872_), .ZN(new_n12876_));
  NAND2_X1   g10440(.A1(new_n12876_), .A2(new_n12781_), .ZN(new_n12877_));
  NAND2_X1   g10441(.A1(new_n12866_), .A2(pi0618), .ZN(new_n12878_));
  AOI21_X1   g10442(.A1(new_n12878_), .A2(new_n12877_), .B(new_n12785_), .ZN(new_n12879_));
  INV_X1     g10443(.I(pi0627), .ZN(new_n12880_));
  OR2_X2     g10444(.A1(new_n12784_), .A2(new_n12880_), .Z(new_n12881_));
  OAI22_X1   g10445(.A1(new_n12875_), .A2(pi0627), .B1(new_n12879_), .B2(new_n12881_), .ZN(new_n12882_));
  NOR2_X1    g10446(.A1(new_n12882_), .A2(new_n12779_), .ZN(new_n12883_));
  AOI21_X1   g10447(.A1(new_n12779_), .A2(new_n12866_), .B(new_n12883_), .ZN(new_n12884_));
  OAI21_X1   g10448(.A1(new_n12884_), .A2(pi0789), .B(new_n12819_), .ZN(new_n12885_));
  XNOR2_X1   g10449(.A1(pi0627), .A2(pi1154), .ZN(new_n12886_));
  NOR2_X1    g10450(.A1(new_n12886_), .A2(new_n12779_), .ZN(new_n12887_));
  INV_X1     g10451(.I(new_n12887_), .ZN(new_n12888_));
  NOR2_X1    g10452(.A1(new_n12888_), .A2(new_n3043_), .ZN(new_n12889_));
  NOR2_X1    g10453(.A1(new_n12876_), .A2(new_n12889_), .ZN(new_n12890_));
  NOR2_X1    g10454(.A1(new_n12890_), .A2(pi0619), .ZN(new_n12891_));
  NOR2_X1    g10455(.A1(new_n12884_), .A2(new_n12793_), .ZN(new_n12892_));
  OAI21_X1   g10456(.A1(new_n12892_), .A2(new_n12891_), .B(pi1159), .ZN(new_n12893_));
  NAND3_X1   g10457(.A1(new_n12893_), .A2(pi0648), .A3(new_n12795_), .ZN(new_n12894_));
  INV_X1     g10458(.I(pi0648), .ZN(new_n12895_));
  INV_X1     g10459(.I(new_n12890_), .ZN(new_n12896_));
  NAND2_X1   g10460(.A1(new_n12896_), .A2(pi0619), .ZN(new_n12897_));
  OAI21_X1   g10461(.A1(new_n12884_), .A2(pi0619), .B(new_n12897_), .ZN(new_n12898_));
  AOI21_X1   g10462(.A1(new_n12898_), .A2(new_n12791_), .B(new_n12799_), .ZN(new_n12899_));
  AOI21_X1   g10463(.A1(new_n12899_), .A2(new_n12895_), .B(new_n12796_), .ZN(new_n12900_));
  AOI21_X1   g10464(.A1(new_n12900_), .A2(new_n12894_), .B(new_n12885_), .ZN(new_n12901_));
  NOR2_X1    g10465(.A1(new_n12814_), .A2(new_n12745_), .ZN(new_n12902_));
  NOR2_X1    g10466(.A1(pi0641), .A2(pi1158), .ZN(new_n12903_));
  INV_X1     g10467(.I(new_n12903_), .ZN(new_n12904_));
  NOR2_X1    g10468(.A1(new_n12904_), .A2(new_n12747_), .ZN(new_n12905_));
  AOI21_X1   g10469(.A1(new_n12747_), .A2(new_n12902_), .B(new_n12905_), .ZN(new_n12906_));
  NOR2_X1    g10470(.A1(new_n12791_), .A2(pi0648), .ZN(new_n12907_));
  NOR2_X1    g10471(.A1(new_n12895_), .A2(pi1159), .ZN(new_n12908_));
  NOR2_X1    g10472(.A1(new_n12907_), .A2(new_n12908_), .ZN(new_n12909_));
  NOR2_X1    g10473(.A1(new_n12909_), .A2(new_n12796_), .ZN(new_n12910_));
  INV_X1     g10474(.I(new_n12910_), .ZN(new_n12911_));
  NOR2_X1    g10475(.A1(new_n12911_), .A2(new_n3043_), .ZN(new_n12912_));
  NOR2_X1    g10476(.A1(new_n12912_), .A2(new_n12906_), .ZN(new_n12913_));
  NOR2_X1    g10477(.A1(new_n12902_), .A2(new_n12903_), .ZN(new_n12914_));
  AOI22_X1   g10478(.A1(new_n12806_), .A2(new_n12914_), .B1(new_n12890_), .B2(new_n12913_), .ZN(new_n12915_));
  NOR2_X1    g10479(.A1(new_n12915_), .A2(new_n12808_), .ZN(new_n12916_));
  NOR2_X1    g10480(.A1(new_n12901_), .A2(new_n12916_), .ZN(new_n12917_));
  AOI21_X1   g10481(.A1(new_n12917_), .A2(pi0628), .B(new_n12811_), .ZN(new_n12918_));
  INV_X1     g10482(.I(pi0629), .ZN(new_n12919_));
  INV_X1     g10483(.I(pi0628), .ZN(new_n12920_));
  NOR2_X1    g10484(.A1(new_n3043_), .A2(new_n12920_), .ZN(new_n12921_));
  INV_X1     g10485(.I(new_n12921_), .ZN(new_n12922_));
  NOR2_X1    g10486(.A1(new_n12910_), .A2(new_n12817_), .ZN(new_n12923_));
  NOR2_X1    g10487(.A1(new_n12923_), .A2(new_n3043_), .ZN(new_n12924_));
  NOR2_X1    g10488(.A1(new_n12896_), .A2(new_n12924_), .ZN(new_n12925_));
  NAND2_X1   g10489(.A1(new_n12925_), .A2(new_n12922_), .ZN(new_n12926_));
  AOI21_X1   g10490(.A1(new_n12926_), .A2(new_n12742_), .B(new_n12919_), .ZN(new_n12927_));
  OAI21_X1   g10491(.A1(new_n12918_), .A2(new_n12742_), .B(new_n12927_), .ZN(new_n12928_));
  NOR2_X1    g10492(.A1(new_n12810_), .A2(new_n12920_), .ZN(new_n12929_));
  AOI21_X1   g10493(.A1(new_n12917_), .A2(new_n12920_), .B(new_n12929_), .ZN(new_n12930_));
  NOR2_X1    g10494(.A1(new_n3043_), .A2(pi0628), .ZN(new_n12931_));
  INV_X1     g10495(.I(new_n12931_), .ZN(new_n12932_));
  NAND2_X1   g10496(.A1(new_n12925_), .A2(new_n12932_), .ZN(new_n12933_));
  AOI21_X1   g10497(.A1(new_n12933_), .A2(pi1156), .B(pi0629), .ZN(new_n12934_));
  OAI21_X1   g10498(.A1(new_n12930_), .A2(pi1156), .B(new_n12934_), .ZN(new_n12935_));
  NAND3_X1   g10499(.A1(new_n12928_), .A2(new_n12935_), .A3(pi0792), .ZN(new_n12936_));
  INV_X1     g10500(.I(pi0792), .ZN(new_n12937_));
  NAND2_X1   g10501(.A1(new_n12917_), .A2(new_n12937_), .ZN(new_n12938_));
  AOI21_X1   g10502(.A1(new_n12936_), .A2(new_n12938_), .B(new_n12741_), .ZN(new_n12939_));
  NOR2_X1    g10503(.A1(new_n12742_), .A2(pi0629), .ZN(new_n12940_));
  NOR2_X1    g10504(.A1(new_n12919_), .A2(pi1156), .ZN(new_n12941_));
  NOR2_X1    g10505(.A1(new_n12940_), .A2(new_n12941_), .ZN(new_n12942_));
  NOR2_X1    g10506(.A1(new_n12942_), .A2(new_n12937_), .ZN(new_n12943_));
  NOR2_X1    g10507(.A1(new_n12810_), .A2(new_n12943_), .ZN(new_n12944_));
  AOI21_X1   g10508(.A1(new_n12744_), .A2(new_n12943_), .B(new_n12944_), .ZN(new_n12945_));
  NOR2_X1    g10509(.A1(new_n12945_), .A2(pi0647), .ZN(new_n12946_));
  OAI21_X1   g10510(.A1(new_n12939_), .A2(new_n12946_), .B(pi1157), .ZN(new_n12947_));
  NOR2_X1    g10511(.A1(new_n12742_), .A2(pi0628), .ZN(new_n12948_));
  NOR2_X1    g10512(.A1(new_n12920_), .A2(pi1156), .ZN(new_n12949_));
  NOR2_X1    g10513(.A1(new_n12948_), .A2(new_n12949_), .ZN(new_n12950_));
  NOR2_X1    g10514(.A1(new_n12950_), .A2(new_n12937_), .ZN(new_n12951_));
  INV_X1     g10515(.I(new_n12951_), .ZN(new_n12952_));
  NOR2_X1    g10516(.A1(new_n12952_), .A2(new_n3043_), .ZN(new_n12953_));
  INV_X1     g10517(.I(new_n12953_), .ZN(new_n12954_));
  NAND2_X1   g10518(.A1(new_n12925_), .A2(new_n12954_), .ZN(new_n12955_));
  NAND2_X1   g10519(.A1(new_n12955_), .A2(new_n12741_), .ZN(new_n12956_));
  NOR2_X1    g10520(.A1(new_n12743_), .A2(new_n12741_), .ZN(new_n12957_));
  INV_X1     g10521(.I(new_n12957_), .ZN(new_n12958_));
  AOI21_X1   g10522(.A1(new_n12956_), .A2(new_n12958_), .B(pi1157), .ZN(new_n12959_));
  INV_X1     g10523(.I(new_n12959_), .ZN(new_n12960_));
  NAND3_X1   g10524(.A1(new_n12947_), .A2(pi0630), .A3(new_n12960_), .ZN(new_n12961_));
  NAND2_X1   g10525(.A1(new_n12936_), .A2(new_n12938_), .ZN(new_n12962_));
  NOR2_X1    g10526(.A1(new_n12945_), .A2(new_n12741_), .ZN(new_n12963_));
  AOI21_X1   g10527(.A1(new_n12962_), .A2(new_n12741_), .B(new_n12963_), .ZN(new_n12964_));
  INV_X1     g10528(.I(pi1157), .ZN(new_n12965_));
  NAND2_X1   g10529(.A1(new_n12955_), .A2(pi0647), .ZN(new_n12966_));
  NAND2_X1   g10530(.A1(new_n12744_), .A2(new_n12741_), .ZN(new_n12967_));
  AOI21_X1   g10531(.A1(new_n12966_), .A2(new_n12967_), .B(new_n12965_), .ZN(new_n12968_));
  NOR2_X1    g10532(.A1(new_n12968_), .A2(pi0630), .ZN(new_n12969_));
  OAI21_X1   g10533(.A1(new_n12964_), .A2(pi1157), .B(new_n12969_), .ZN(new_n12970_));
  NAND3_X1   g10534(.A1(new_n12961_), .A2(new_n12970_), .A3(pi0787), .ZN(new_n12971_));
  INV_X1     g10535(.I(pi0787), .ZN(new_n12972_));
  NAND2_X1   g10536(.A1(new_n12962_), .A2(new_n12972_), .ZN(new_n12973_));
  AOI21_X1   g10537(.A1(new_n12971_), .A2(new_n12973_), .B(pi0644), .ZN(new_n12974_));
  INV_X1     g10538(.I(pi0644), .ZN(new_n12975_));
  OR2_X2     g10539(.A1(new_n12968_), .A2(new_n12972_), .Z(new_n12976_));
  OAI22_X1   g10540(.A1(new_n12976_), .A2(new_n12959_), .B1(pi0787), .B2(new_n12955_), .ZN(new_n12977_));
  NOR2_X1    g10541(.A1(new_n12977_), .A2(new_n12975_), .ZN(new_n12978_));
  OAI21_X1   g10542(.A1(new_n12974_), .A2(new_n12978_), .B(new_n12740_), .ZN(new_n12979_));
  NOR2_X1    g10543(.A1(new_n12965_), .A2(pi0630), .ZN(new_n12980_));
  INV_X1     g10544(.I(pi0630), .ZN(new_n12981_));
  NOR2_X1    g10545(.A1(new_n12981_), .A2(pi1157), .ZN(new_n12982_));
  NOR2_X1    g10546(.A1(new_n12980_), .A2(new_n12982_), .ZN(new_n12983_));
  NOR2_X1    g10547(.A1(new_n12983_), .A2(new_n12972_), .ZN(new_n12984_));
  INV_X1     g10548(.I(new_n12984_), .ZN(new_n12985_));
  NAND2_X1   g10549(.A1(new_n12945_), .A2(new_n12985_), .ZN(new_n12986_));
  OAI21_X1   g10550(.A1(new_n12744_), .A2(new_n12985_), .B(new_n12986_), .ZN(new_n12987_));
  NOR2_X1    g10551(.A1(new_n12987_), .A2(pi0644), .ZN(new_n12988_));
  NOR2_X1    g10552(.A1(new_n12743_), .A2(new_n12975_), .ZN(new_n12989_));
  OAI21_X1   g10553(.A1(new_n12988_), .A2(new_n12989_), .B(pi0715), .ZN(new_n12990_));
  NAND3_X1   g10554(.A1(new_n12979_), .A2(new_n12739_), .A3(new_n12990_), .ZN(new_n12991_));
  NAND2_X1   g10555(.A1(new_n12971_), .A2(new_n12973_), .ZN(new_n12992_));
  NOR2_X1    g10556(.A1(new_n12977_), .A2(pi0644), .ZN(new_n12993_));
  AOI21_X1   g10557(.A1(new_n12992_), .A2(pi0644), .B(new_n12993_), .ZN(new_n12994_));
  NAND2_X1   g10558(.A1(new_n12744_), .A2(new_n12975_), .ZN(new_n12995_));
  OAI21_X1   g10559(.A1(new_n12987_), .A2(new_n12975_), .B(new_n12995_), .ZN(new_n12996_));
  AOI21_X1   g10560(.A1(new_n12996_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n12997_));
  OAI21_X1   g10561(.A1(new_n12994_), .A2(new_n12740_), .B(new_n12997_), .ZN(new_n12998_));
  NAND3_X1   g10562(.A1(new_n12991_), .A2(new_n12998_), .A3(pi0790), .ZN(new_n12999_));
  INV_X1     g10563(.I(pi0790), .ZN(new_n13000_));
  NAND2_X1   g10564(.A1(new_n12992_), .A2(new_n13000_), .ZN(new_n13001_));
  AOI21_X1   g10565(.A1(new_n12999_), .A2(new_n13001_), .B(new_n12738_), .ZN(new_n13002_));
  AOI21_X1   g10566(.A1(po1038), .A2(new_n7934_), .B(pi0832), .ZN(new_n13003_));
  NOR2_X1    g10567(.A1(new_n5346_), .A2(new_n3043_), .ZN(new_n13004_));
  NOR2_X1    g10568(.A1(new_n13004_), .A2(new_n3265_), .ZN(new_n13005_));
  NOR2_X1    g10569(.A1(new_n10302_), .A2(new_n3040_), .ZN(po1106));
  NAND2_X1   g10570(.A1(new_n9121_), .A2(new_n2501_), .ZN(new_n13007_));
  AOI21_X1   g10571(.A1(new_n2970_), .A2(pi0102), .B(pi0098), .ZN(new_n13008_));
  NAND2_X1   g10572(.A1(new_n13008_), .A2(new_n13007_), .ZN(new_n13009_));
  NAND2_X1   g10573(.A1(new_n6672_), .A2(new_n6667_), .ZN(new_n13010_));
  NOR4_X1    g10574(.A1(new_n13009_), .A2(new_n7293_), .A3(new_n7469_), .A4(new_n13010_), .ZN(new_n13011_));
  NOR2_X1    g10575(.A1(new_n13011_), .A2(pi0040), .ZN(new_n13012_));
  OAI21_X1   g10576(.A1(new_n13012_), .A2(new_n8342_), .B(new_n2704_), .ZN(new_n13013_));
  OAI21_X1   g10577(.A1(new_n2553_), .A2(new_n2818_), .B(pi0252), .ZN(new_n13014_));
  NAND3_X1   g10578(.A1(new_n8309_), .A2(new_n2818_), .A3(new_n7569_), .ZN(new_n13015_));
  NOR3_X1    g10579(.A1(new_n2845_), .A2(pi0091), .A3(new_n2764_), .ZN(new_n13016_));
  NAND4_X1   g10580(.A1(new_n2853_), .A2(new_n2864_), .A3(new_n2857_), .A4(new_n8330_), .ZN(new_n13017_));
  OAI21_X1   g10581(.A1(new_n13017_), .A2(new_n5590_), .B(new_n2844_), .ZN(new_n13018_));
  NOR3_X1    g10582(.A1(new_n13009_), .A2(new_n7271_), .A3(new_n13010_), .ZN(new_n13019_));
  OAI21_X1   g10583(.A1(new_n13018_), .A2(new_n13019_), .B(new_n13016_), .ZN(new_n13020_));
  AOI21_X1   g10584(.A1(new_n13020_), .A2(new_n2743_), .B(new_n13015_), .ZN(new_n13021_));
  OAI21_X1   g10585(.A1(new_n13021_), .A2(new_n13014_), .B(new_n13013_), .ZN(new_n13022_));
  NOR2_X1    g10586(.A1(new_n13022_), .A2(new_n7456_), .ZN(new_n13023_));
  AOI21_X1   g10587(.A1(new_n13023_), .A2(po1106), .B(new_n3025_), .ZN(new_n13024_));
  INV_X1     g10588(.I(new_n13024_), .ZN(new_n13025_));
  NOR4_X1    g10589(.A1(new_n13022_), .A2(new_n3040_), .A3(new_n7456_), .A4(new_n9893_), .ZN(new_n13026_));
  AOI21_X1   g10590(.A1(new_n13008_), .A2(new_n13007_), .B(pi0088), .ZN(new_n13027_));
  OR3_X2     g10591(.A1(new_n13027_), .A2(new_n7717_), .A3(new_n8914_), .Z(new_n13028_));
  OAI21_X1   g10592(.A1(new_n13028_), .A2(pi0252), .B(new_n2818_), .ZN(new_n13029_));
  NOR3_X1    g10593(.A1(new_n13027_), .A2(new_n8914_), .A3(new_n2756_), .ZN(new_n13030_));
  OAI21_X1   g10594(.A1(new_n13030_), .A2(new_n13018_), .B(new_n13016_), .ZN(new_n13031_));
  NAND3_X1   g10595(.A1(new_n8309_), .A2(pi0252), .A3(new_n7569_), .ZN(new_n13032_));
  AOI21_X1   g10596(.A1(new_n13031_), .A2(new_n2743_), .B(new_n13032_), .ZN(new_n13033_));
  NOR2_X1    g10597(.A1(new_n13033_), .A2(new_n13029_), .ZN(new_n13034_));
  NOR3_X1    g10598(.A1(new_n13034_), .A2(new_n6259_), .A3(new_n8342_), .ZN(new_n13035_));
  OAI21_X1   g10599(.A1(new_n13026_), .A2(new_n13035_), .B(pi1093), .ZN(new_n13036_));
  NAND2_X1   g10600(.A1(new_n13036_), .A2(new_n5532_), .ZN(new_n13037_));
  NAND2_X1   g10601(.A1(new_n13037_), .A2(new_n13025_), .ZN(new_n13038_));
  OR2_X2     g10602(.A1(new_n13036_), .A2(pi1091), .Z(new_n13039_));
  AOI21_X1   g10603(.A1(new_n13038_), .A2(new_n13039_), .B(pi0210), .ZN(new_n13040_));
  NOR2_X1    g10604(.A1(new_n9893_), .A2(new_n3040_), .ZN(new_n13041_));
  NAND2_X1   g10605(.A1(new_n5612_), .A2(pi0032), .ZN(new_n13042_));
  NAND3_X1   g10606(.A1(new_n13042_), .A2(new_n2462_), .A3(new_n8913_), .ZN(new_n13043_));
  INV_X1     g10607(.I(new_n3400_), .ZN(new_n13044_));
  OAI21_X1   g10608(.A1(new_n13033_), .A2(new_n13029_), .B(new_n13044_), .ZN(new_n13045_));
  AOI21_X1   g10609(.A1(new_n13045_), .A2(new_n2725_), .B(new_n13043_), .ZN(new_n13046_));
  AOI22_X1   g10610(.A1(new_n13046_), .A2(pi0824), .B1(new_n13023_), .B2(new_n13041_), .ZN(new_n13047_));
  NOR2_X1    g10611(.A1(new_n13047_), .A2(new_n6871_), .ZN(new_n13048_));
  INV_X1     g10612(.I(new_n13048_), .ZN(new_n13049_));
  AOI21_X1   g10613(.A1(new_n13022_), .A2(new_n2725_), .B(new_n13043_), .ZN(new_n13050_));
  NAND3_X1   g10614(.A1(new_n13050_), .A2(new_n5428_), .A3(pi0829), .ZN(new_n13051_));
  AOI21_X1   g10615(.A1(new_n13047_), .A2(new_n13051_), .B(new_n3041_), .ZN(new_n13052_));
  OAI21_X1   g10616(.A1(new_n13052_), .A2(new_n3024_), .B(new_n13025_), .ZN(new_n13053_));
  NAND2_X1   g10617(.A1(new_n13053_), .A2(new_n13049_), .ZN(new_n13054_));
  AOI21_X1   g10618(.A1(new_n13054_), .A2(pi0210), .B(new_n13040_), .ZN(new_n13055_));
  NOR2_X1    g10619(.A1(new_n13055_), .A2(new_n2628_), .ZN(new_n13056_));
  AOI21_X1   g10620(.A1(new_n13038_), .A2(new_n13039_), .B(pi0198), .ZN(new_n13057_));
  AOI21_X1   g10621(.A1(new_n13054_), .A2(pi0198), .B(new_n13057_), .ZN(new_n13058_));
  NOR2_X1    g10622(.A1(new_n13058_), .A2(pi0299), .ZN(new_n13059_));
  NOR2_X1    g10623(.A1(new_n13056_), .A2(new_n13059_), .ZN(new_n13060_));
  NOR2_X1    g10624(.A1(new_n13060_), .A2(pi0039), .ZN(new_n13061_));
  OAI21_X1   g10625(.A1(new_n2530_), .A2(new_n3043_), .B(pi0120), .ZN(new_n13062_));
  INV_X1     g10626(.I(new_n13062_), .ZN(new_n13063_));
  NAND2_X1   g10627(.A1(new_n13062_), .A2(new_n3022_), .ZN(new_n13064_));
  NOR2_X1    g10628(.A1(new_n3045_), .A2(pi0824), .ZN(new_n13065_));
  INV_X1     g10629(.I(new_n13065_), .ZN(new_n13066_));
  NAND2_X1   g10630(.A1(new_n8285_), .A2(new_n8282_), .ZN(new_n13067_));
  INV_X1     g10631(.I(new_n13067_), .ZN(new_n13068_));
  NAND4_X1   g10632(.A1(new_n2547_), .A2(new_n2523_), .A3(new_n2529_), .A4(new_n13068_), .ZN(new_n13069_));
  AOI21_X1   g10633(.A1(new_n13069_), .A2(new_n13066_), .B(new_n3040_), .ZN(new_n13070_));
  OAI21_X1   g10634(.A1(new_n8283_), .A2(new_n5391_), .B(new_n5428_), .ZN(new_n13071_));
  NAND3_X1   g10635(.A1(new_n13070_), .A2(new_n13071_), .A3(pi1093), .ZN(new_n13072_));
  AOI21_X1   g10636(.A1(new_n13072_), .A2(new_n10903_), .B(new_n13064_), .ZN(new_n13073_));
  INV_X1     g10637(.I(new_n13073_), .ZN(new_n13074_));
  OAI21_X1   g10638(.A1(new_n13069_), .A2(new_n3040_), .B(pi0829), .ZN(new_n13075_));
  NAND2_X1   g10639(.A1(new_n13075_), .A2(new_n6712_), .ZN(new_n13076_));
  AOI21_X1   g10640(.A1(new_n13070_), .A2(new_n13071_), .B(pi0829), .ZN(new_n13077_));
  NOR4_X1    g10641(.A1(new_n8283_), .A2(new_n5532_), .A3(new_n3043_), .A4(new_n5391_), .ZN(new_n13078_));
  INV_X1     g10642(.I(new_n13078_), .ZN(new_n13079_));
  OAI21_X1   g10643(.A1(new_n13077_), .A2(new_n13076_), .B(new_n13079_), .ZN(new_n13080_));
  AOI21_X1   g10644(.A1(new_n13080_), .A2(pi1091), .B(pi0120), .ZN(new_n13081_));
  OAI21_X1   g10645(.A1(new_n13081_), .A2(new_n13063_), .B(new_n13074_), .ZN(new_n13082_));
  NAND2_X1   g10646(.A1(new_n13082_), .A2(new_n5402_), .ZN(new_n13083_));
  NAND2_X1   g10647(.A1(new_n2531_), .A2(pi0120), .ZN(new_n13084_));
  NOR2_X1    g10648(.A1(new_n8283_), .A2(new_n5391_), .ZN(new_n13085_));
  NAND2_X1   g10649(.A1(new_n13085_), .A2(new_n10903_), .ZN(new_n13086_));
  NAND2_X1   g10650(.A1(new_n13086_), .A2(new_n13084_), .ZN(new_n13087_));
  NAND2_X1   g10651(.A1(new_n13087_), .A2(new_n3042_), .ZN(new_n13088_));
  NOR2_X1    g10652(.A1(new_n13088_), .A2(new_n5691_), .ZN(new_n13089_));
  AOI21_X1   g10653(.A1(new_n13082_), .A2(new_n5691_), .B(new_n13089_), .ZN(new_n13090_));
  OAI21_X1   g10654(.A1(new_n13090_), .A2(new_n5402_), .B(new_n13083_), .ZN(new_n13091_));
  NAND2_X1   g10655(.A1(new_n13090_), .A2(pi0681), .ZN(new_n13092_));
  OAI21_X1   g10656(.A1(new_n13091_), .A2(pi0681), .B(new_n13092_), .ZN(new_n13093_));
  AOI21_X1   g10657(.A1(new_n13093_), .A2(new_n5419_), .B(new_n5421_), .ZN(new_n13094_));
  NOR2_X1    g10658(.A1(pi0614), .A2(pi0616), .ZN(new_n13095_));
  INV_X1     g10659(.I(new_n13095_), .ZN(new_n13096_));
  NOR3_X1    g10660(.A1(new_n5398_), .A2(new_n12751_), .A3(pi0642), .ZN(new_n13097_));
  AOI21_X1   g10661(.A1(new_n13086_), .A2(new_n13084_), .B(new_n3043_), .ZN(new_n13098_));
  INV_X1     g10662(.I(new_n13097_), .ZN(new_n13099_));
  NAND2_X1   g10663(.A1(new_n13098_), .A2(new_n13099_), .ZN(new_n13100_));
  INV_X1     g10664(.I(new_n13100_), .ZN(new_n13101_));
  AOI21_X1   g10665(.A1(new_n13082_), .A2(new_n13097_), .B(new_n13101_), .ZN(new_n13102_));
  NOR2_X1    g10666(.A1(new_n13102_), .A2(new_n13096_), .ZN(new_n13103_));
  NAND2_X1   g10667(.A1(new_n13098_), .A2(new_n13096_), .ZN(new_n13104_));
  INV_X1     g10668(.I(new_n13104_), .ZN(new_n13105_));
  NOR3_X1    g10669(.A1(new_n13103_), .A2(new_n5399_), .A3(new_n13105_), .ZN(new_n13106_));
  NOR2_X1    g10670(.A1(new_n13098_), .A2(new_n5437_), .ZN(new_n13107_));
  INV_X1     g10671(.I(new_n13107_), .ZN(new_n13108_));
  OAI21_X1   g10672(.A1(new_n13082_), .A2(new_n5398_), .B(new_n13108_), .ZN(new_n13109_));
  NOR3_X1    g10673(.A1(new_n13109_), .A2(pi0614), .A3(new_n5403_), .ZN(new_n13110_));
  INV_X1     g10674(.I(pi0616), .ZN(new_n13111_));
  NAND2_X1   g10675(.A1(new_n13088_), .A2(pi0616), .ZN(new_n13112_));
  NAND3_X1   g10676(.A1(new_n13112_), .A2(new_n5405_), .A3(new_n5403_), .ZN(new_n13113_));
  AOI21_X1   g10677(.A1(new_n13102_), .A2(new_n13111_), .B(new_n13113_), .ZN(new_n13114_));
  NOR2_X1    g10678(.A1(new_n13110_), .A2(new_n13114_), .ZN(new_n13115_));
  NOR2_X1    g10679(.A1(pi0661), .A2(pi0681), .ZN(new_n13116_));
  INV_X1     g10680(.I(new_n13116_), .ZN(new_n13117_));
  NOR2_X1    g10681(.A1(new_n13117_), .A2(pi0662), .ZN(new_n13118_));
  INV_X1     g10682(.I(new_n13118_), .ZN(new_n13119_));
  NAND2_X1   g10683(.A1(new_n13098_), .A2(new_n13119_), .ZN(new_n13120_));
  NOR2_X1    g10684(.A1(new_n13120_), .A2(new_n5405_), .ZN(new_n13121_));
  AOI21_X1   g10685(.A1(new_n13088_), .A2(new_n12821_), .B(new_n13119_), .ZN(new_n13122_));
  NAND2_X1   g10686(.A1(new_n13122_), .A2(pi0614), .ZN(new_n13123_));
  AOI21_X1   g10687(.A1(new_n13109_), .A2(pi0680), .B(new_n13123_), .ZN(new_n13124_));
  NOR3_X1    g10688(.A1(new_n13124_), .A2(pi0681), .A3(new_n13121_), .ZN(new_n13125_));
  AOI21_X1   g10689(.A1(new_n13125_), .A2(new_n13115_), .B(new_n13106_), .ZN(new_n13126_));
  OAI21_X1   g10690(.A1(new_n13126_), .A2(new_n5419_), .B(new_n13094_), .ZN(new_n13127_));
  OAI21_X1   g10691(.A1(new_n13093_), .A2(new_n5420_), .B(new_n3304_), .ZN(new_n13128_));
  NOR2_X1    g10692(.A1(new_n13098_), .A2(new_n3304_), .ZN(new_n13129_));
  INV_X1     g10693(.I(new_n13129_), .ZN(new_n13130_));
  AOI21_X1   g10694(.A1(new_n13128_), .A2(new_n13130_), .B(pi0215), .ZN(new_n13131_));
  OAI21_X1   g10695(.A1(new_n13127_), .A2(new_n3303_), .B(new_n13131_), .ZN(new_n13132_));
  NAND2_X1   g10696(.A1(new_n9149_), .A2(new_n5392_), .ZN(new_n13133_));
  OAI21_X1   g10697(.A1(new_n13133_), .A2(new_n3043_), .B(new_n10903_), .ZN(new_n13134_));
  NOR3_X1    g10698(.A1(new_n5396_), .A2(new_n10903_), .A3(new_n5428_), .ZN(new_n13135_));
  NOR2_X1    g10699(.A1(new_n2530_), .A2(new_n3043_), .ZN(new_n13136_));
  INV_X1     g10700(.I(new_n5329_), .ZN(new_n13137_));
  NAND4_X1   g10701(.A1(new_n5395_), .A2(pi0950), .A3(new_n5532_), .A4(new_n13137_), .ZN(new_n13138_));
  AOI21_X1   g10702(.A1(new_n13136_), .A2(new_n13138_), .B(new_n10903_), .ZN(new_n13139_));
  OAI22_X1   g10703(.A1(new_n3022_), .A2(new_n13139_), .B1(new_n13064_), .B2(new_n13135_), .ZN(new_n13140_));
  NAND3_X1   g10704(.A1(new_n13140_), .A2(new_n13097_), .A3(new_n13134_), .ZN(new_n13141_));
  NAND2_X1   g10705(.A1(new_n13141_), .A2(new_n13100_), .ZN(new_n13142_));
  AOI21_X1   g10706(.A1(new_n13142_), .A2(new_n13095_), .B(new_n13105_), .ZN(new_n13143_));
  INV_X1     g10707(.I(new_n13143_), .ZN(new_n13144_));
  NOR2_X1    g10708(.A1(new_n13144_), .A2(new_n5399_), .ZN(new_n13145_));
  NAND2_X1   g10709(.A1(new_n13122_), .A2(pi0616), .ZN(new_n13146_));
  NOR2_X1    g10710(.A1(new_n13064_), .A2(new_n13135_), .ZN(new_n13147_));
  NOR2_X1    g10711(.A1(new_n13139_), .A2(new_n3022_), .ZN(new_n13148_));
  OAI21_X1   g10712(.A1(new_n13147_), .A2(new_n13148_), .B(new_n13134_), .ZN(new_n13149_));
  AOI21_X1   g10713(.A1(new_n13149_), .A2(new_n5437_), .B(new_n13107_), .ZN(new_n13150_));
  NOR2_X1    g10714(.A1(new_n13150_), .A2(new_n12821_), .ZN(new_n13151_));
  OAI22_X1   g10715(.A1(new_n13151_), .A2(new_n13146_), .B1(new_n13111_), .B2(new_n13120_), .ZN(new_n13152_));
  NOR2_X1    g10716(.A1(new_n13088_), .A2(new_n5405_), .ZN(new_n13153_));
  AOI21_X1   g10717(.A1(new_n13141_), .A2(new_n13100_), .B(pi0614), .ZN(new_n13154_));
  NOR2_X1    g10718(.A1(new_n13154_), .A2(new_n13153_), .ZN(new_n13155_));
  NOR3_X1    g10719(.A1(new_n13155_), .A2(pi0616), .A3(new_n13118_), .ZN(new_n13156_));
  NOR2_X1    g10720(.A1(new_n13119_), .A2(pi0616), .ZN(new_n13157_));
  OAI21_X1   g10721(.A1(new_n13150_), .A2(new_n12821_), .B(new_n13157_), .ZN(new_n13158_));
  NOR3_X1    g10722(.A1(new_n13154_), .A2(pi0616), .A3(new_n13153_), .ZN(new_n13159_));
  AOI21_X1   g10723(.A1(new_n13159_), .A2(new_n12821_), .B(new_n13158_), .ZN(new_n13160_));
  NOR4_X1    g10724(.A1(new_n13160_), .A2(new_n13152_), .A3(new_n13156_), .A4(pi0681), .ZN(new_n13161_));
  NOR3_X1    g10725(.A1(new_n13161_), .A2(new_n5419_), .A3(new_n13145_), .ZN(new_n13162_));
  INV_X1     g10726(.I(new_n5401_), .ZN(new_n13163_));
  OAI21_X1   g10727(.A1(new_n5398_), .A2(new_n13163_), .B(new_n13149_), .ZN(new_n13164_));
  NAND3_X1   g10728(.A1(new_n13143_), .A2(new_n5437_), .A3(new_n5401_), .ZN(new_n13165_));
  AOI21_X1   g10729(.A1(new_n13165_), .A2(new_n13164_), .B(new_n13117_), .ZN(new_n13166_));
  NOR2_X1    g10730(.A1(new_n13142_), .A2(pi0614), .ZN(new_n13167_));
  NAND2_X1   g10731(.A1(new_n13098_), .A2(new_n5437_), .ZN(new_n13168_));
  OAI21_X1   g10732(.A1(new_n13149_), .A2(new_n5437_), .B(new_n13168_), .ZN(new_n13169_));
  INV_X1     g10733(.I(new_n13169_), .ZN(new_n13170_));
  AOI21_X1   g10734(.A1(new_n13167_), .A2(new_n13111_), .B(new_n13170_), .ZN(new_n13171_));
  NOR2_X1    g10735(.A1(new_n13171_), .A2(new_n13116_), .ZN(new_n13172_));
  NOR3_X1    g10736(.A1(new_n13166_), .A2(new_n13172_), .A3(new_n5418_), .ZN(new_n13173_));
  OAI21_X1   g10737(.A1(new_n13162_), .A2(new_n13173_), .B(new_n5420_), .ZN(new_n13174_));
  NOR2_X1    g10738(.A1(new_n13166_), .A2(new_n13172_), .ZN(new_n13175_));
  AOI21_X1   g10739(.A1(new_n13175_), .A2(new_n5421_), .B(new_n2436_), .ZN(new_n13176_));
  NAND2_X1   g10740(.A1(new_n13174_), .A2(new_n13176_), .ZN(new_n13177_));
  AOI21_X1   g10741(.A1(new_n13132_), .A2(new_n13177_), .B(new_n2628_), .ZN(new_n13178_));
  NOR2_X1    g10742(.A1(new_n13161_), .A2(new_n13145_), .ZN(new_n13179_));
  NAND2_X1   g10743(.A1(new_n13179_), .A2(new_n5446_), .ZN(new_n13180_));
  NAND2_X1   g10744(.A1(new_n13175_), .A2(new_n5445_), .ZN(new_n13181_));
  NAND3_X1   g10745(.A1(new_n13180_), .A2(pi0223), .A3(new_n13181_), .ZN(new_n13182_));
  NOR2_X1    g10746(.A1(new_n13093_), .A2(new_n5446_), .ZN(new_n13183_));
  AOI21_X1   g10747(.A1(new_n13126_), .A2(new_n5446_), .B(new_n13183_), .ZN(new_n13184_));
  NOR2_X1    g10748(.A1(new_n13088_), .A2(new_n2642_), .ZN(new_n13185_));
  NOR2_X1    g10749(.A1(new_n13185_), .A2(pi0223), .ZN(new_n13186_));
  OAI21_X1   g10750(.A1(new_n13184_), .A2(new_n2641_), .B(new_n13186_), .ZN(new_n13187_));
  AOI21_X1   g10751(.A1(new_n13187_), .A2(new_n13182_), .B(pi0299), .ZN(new_n13188_));
  NOR3_X1    g10752(.A1(new_n13178_), .A2(new_n13188_), .A3(new_n2627_), .ZN(new_n13189_));
  NOR3_X1    g10753(.A1(new_n13189_), .A2(pi0038), .A3(new_n13061_), .ZN(new_n13190_));
  NOR2_X1    g10754(.A1(new_n13190_), .A2(new_n13005_), .ZN(new_n13191_));
  NAND2_X1   g10755(.A1(new_n13191_), .A2(new_n2609_), .ZN(new_n13192_));
  INV_X1     g10756(.I(new_n13192_), .ZN(new_n13193_));
  NOR2_X1    g10757(.A1(new_n13193_), .A2(pi0140), .ZN(new_n13194_));
  AOI21_X1   g10758(.A1(new_n13194_), .A2(pi0644), .B(new_n12740_), .ZN(new_n13195_));
  INV_X1     g10759(.I(new_n13194_), .ZN(new_n13196_));
  NOR2_X1    g10760(.A1(new_n2609_), .A2(new_n7934_), .ZN(new_n13197_));
  OAI21_X1   g10761(.A1(new_n13053_), .A2(pi0621), .B(new_n13049_), .ZN(new_n13198_));
  NAND3_X1   g10762(.A1(new_n13037_), .A2(new_n13025_), .A3(new_n12752_), .ZN(new_n13199_));
  AOI21_X1   g10763(.A1(new_n13199_), .A2(new_n13039_), .B(pi0210), .ZN(new_n13200_));
  AOI21_X1   g10764(.A1(new_n13198_), .A2(pi0210), .B(new_n13200_), .ZN(new_n13201_));
  NOR3_X1    g10765(.A1(new_n13201_), .A2(new_n2628_), .A3(new_n12751_), .ZN(new_n13202_));
  AOI21_X1   g10766(.A1(new_n13199_), .A2(new_n13039_), .B(pi0198), .ZN(new_n13203_));
  OAI21_X1   g10767(.A1(new_n13048_), .A2(new_n12752_), .B(pi0198), .ZN(new_n13204_));
  AOI21_X1   g10768(.A1(new_n13053_), .A2(new_n13049_), .B(new_n13204_), .ZN(new_n13205_));
  NOR2_X1    g10769(.A1(new_n13205_), .A2(new_n13203_), .ZN(new_n13206_));
  NOR3_X1    g10770(.A1(new_n13206_), .A2(pi0299), .A3(new_n12751_), .ZN(new_n13207_));
  NOR3_X1    g10771(.A1(new_n13202_), .A2(new_n13207_), .A3(pi0039), .ZN(new_n13208_));
  NAND2_X1   g10772(.A1(new_n13149_), .A2(new_n5437_), .ZN(new_n13209_));
  NOR2_X1    g10773(.A1(new_n13088_), .A2(new_n12755_), .ZN(new_n13210_));
  NAND2_X1   g10774(.A1(new_n13209_), .A2(new_n13210_), .ZN(new_n13211_));
  INV_X1     g10775(.I(new_n13209_), .ZN(new_n13212_));
  NAND2_X1   g10776(.A1(new_n13212_), .A2(new_n5408_), .ZN(new_n13213_));
  NAND2_X1   g10777(.A1(new_n13098_), .A2(new_n12754_), .ZN(new_n13214_));
  NOR2_X1    g10778(.A1(new_n13170_), .A2(new_n13214_), .ZN(new_n13215_));
  NAND3_X1   g10779(.A1(new_n13215_), .A2(new_n13213_), .A3(new_n5403_), .ZN(new_n13216_));
  NAND2_X1   g10780(.A1(new_n13216_), .A2(new_n13211_), .ZN(new_n13217_));
  NOR2_X1    g10781(.A1(new_n13169_), .A2(new_n5422_), .ZN(new_n13218_));
  INV_X1     g10782(.I(new_n13218_), .ZN(new_n13219_));
  AOI21_X1   g10783(.A1(new_n13217_), .A2(new_n13219_), .B(new_n2436_), .ZN(new_n13220_));
  INV_X1     g10784(.I(new_n13087_), .ZN(new_n13221_));
  NOR2_X1    g10785(.A1(new_n13221_), .A2(new_n3304_), .ZN(new_n13222_));
  AOI21_X1   g10786(.A1(new_n13222_), .A2(new_n12756_), .B(pi0215), .ZN(new_n13223_));
  INV_X1     g10787(.I(new_n13223_), .ZN(new_n13224_));
  NAND2_X1   g10788(.A1(new_n13082_), .A2(new_n5404_), .ZN(new_n13225_));
  OAI21_X1   g10789(.A1(new_n13090_), .A2(new_n5404_), .B(new_n13225_), .ZN(new_n13226_));
  NAND3_X1   g10790(.A1(new_n13226_), .A2(new_n6764_), .A3(new_n12754_), .ZN(new_n13227_));
  NOR2_X1    g10791(.A1(new_n13109_), .A2(new_n12755_), .ZN(new_n13228_));
  NOR2_X1    g10792(.A1(new_n5404_), .A2(new_n5408_), .ZN(new_n13229_));
  NAND2_X1   g10793(.A1(new_n13214_), .A2(new_n13229_), .ZN(new_n13230_));
  OAI21_X1   g10794(.A1(new_n13228_), .A2(new_n13229_), .B(new_n13230_), .ZN(new_n13231_));
  OAI21_X1   g10795(.A1(new_n6764_), .A2(new_n13231_), .B(new_n13227_), .ZN(new_n13232_));
  AOI21_X1   g10796(.A1(new_n13232_), .A2(new_n3304_), .B(new_n13224_), .ZN(new_n13233_));
  NOR3_X1    g10797(.A1(new_n13233_), .A2(new_n2628_), .A3(new_n13220_), .ZN(new_n13234_));
  NOR2_X1    g10798(.A1(new_n13169_), .A2(new_n5446_), .ZN(new_n13235_));
  AOI21_X1   g10799(.A1(new_n13216_), .A2(new_n13211_), .B(new_n13235_), .ZN(new_n13236_));
  OAI21_X1   g10800(.A1(new_n13236_), .A2(new_n2668_), .B(new_n2628_), .ZN(new_n13237_));
  AOI21_X1   g10801(.A1(new_n13185_), .A2(new_n12754_), .B(pi0223), .ZN(new_n13238_));
  NAND2_X1   g10802(.A1(new_n13226_), .A2(new_n12754_), .ZN(new_n13239_));
  NOR2_X1    g10803(.A1(new_n13239_), .A2(new_n5446_), .ZN(new_n13240_));
  NOR2_X1    g10804(.A1(new_n13231_), .A2(new_n5445_), .ZN(new_n13241_));
  OAI21_X1   g10805(.A1(new_n13240_), .A2(new_n13241_), .B(new_n2642_), .ZN(new_n13242_));
  AOI21_X1   g10806(.A1(new_n13242_), .A2(new_n13238_), .B(new_n13237_), .ZN(new_n13243_));
  NOR3_X1    g10807(.A1(new_n13234_), .A2(new_n2627_), .A3(new_n13243_), .ZN(new_n13244_));
  NOR2_X1    g10808(.A1(new_n13208_), .A2(new_n13244_), .ZN(new_n13245_));
  NAND3_X1   g10809(.A1(new_n13245_), .A2(pi0140), .A3(new_n12750_), .ZN(new_n13246_));
  NAND3_X1   g10810(.A1(new_n13037_), .A2(new_n13025_), .A3(new_n2709_), .ZN(new_n13247_));
  OAI21_X1   g10811(.A1(new_n13053_), .A2(new_n2709_), .B(new_n13247_), .ZN(new_n13248_));
  AOI21_X1   g10812(.A1(new_n13248_), .A2(pi0621), .B(new_n12751_), .ZN(new_n13249_));
  OAI21_X1   g10813(.A1(new_n13249_), .A2(new_n13055_), .B(pi0299), .ZN(new_n13250_));
  OAI21_X1   g10814(.A1(new_n13205_), .A2(new_n13203_), .B(new_n12751_), .ZN(new_n13251_));
  NAND3_X1   g10815(.A1(new_n13037_), .A2(new_n13025_), .A3(new_n2672_), .ZN(new_n13252_));
  OAI21_X1   g10816(.A1(new_n13053_), .A2(new_n2672_), .B(new_n13252_), .ZN(new_n13253_));
  NAND2_X1   g10817(.A1(new_n13253_), .A2(pi0621), .ZN(new_n13254_));
  NAND3_X1   g10818(.A1(new_n13251_), .A2(new_n2628_), .A3(new_n13254_), .ZN(new_n13255_));
  NAND2_X1   g10819(.A1(new_n13255_), .A2(new_n13250_), .ZN(new_n13256_));
  NAND2_X1   g10820(.A1(new_n13256_), .A2(new_n2627_), .ZN(new_n13257_));
  AOI21_X1   g10821(.A1(new_n13098_), .A2(new_n12753_), .B(new_n5437_), .ZN(new_n13258_));
  AOI21_X1   g10822(.A1(new_n13085_), .A2(new_n3042_), .B(pi0120), .ZN(new_n13259_));
  NOR2_X1    g10823(.A1(new_n13259_), .A2(new_n13139_), .ZN(new_n13260_));
  NAND2_X1   g10824(.A1(new_n13260_), .A2(new_n12753_), .ZN(new_n13261_));
  AOI21_X1   g10825(.A1(new_n5437_), .A2(new_n13261_), .B(new_n13258_), .ZN(new_n13262_));
  NOR2_X1    g10826(.A1(new_n13262_), .A2(new_n12751_), .ZN(new_n13263_));
  INV_X1     g10827(.I(new_n5408_), .ZN(new_n13264_));
  NOR2_X1    g10828(.A1(new_n13088_), .A2(new_n12754_), .ZN(new_n13265_));
  NAND2_X1   g10829(.A1(new_n13265_), .A2(new_n13264_), .ZN(new_n13266_));
  AOI21_X1   g10830(.A1(new_n13088_), .A2(new_n12751_), .B(new_n13264_), .ZN(new_n13267_));
  OAI21_X1   g10831(.A1(new_n13262_), .A2(new_n12751_), .B(new_n13267_), .ZN(new_n13268_));
  NAND2_X1   g10832(.A1(new_n13268_), .A2(new_n13266_), .ZN(new_n13269_));
  NAND2_X1   g10833(.A1(new_n13269_), .A2(new_n5403_), .ZN(new_n13270_));
  NAND2_X1   g10834(.A1(new_n13150_), .A2(new_n5404_), .ZN(new_n13271_));
  OAI21_X1   g10835(.A1(new_n13263_), .A2(new_n13271_), .B(new_n13270_), .ZN(new_n13272_));
  NAND2_X1   g10836(.A1(new_n13272_), .A2(new_n5446_), .ZN(new_n13273_));
  INV_X1     g10837(.I(new_n13149_), .ZN(new_n13274_));
  NOR2_X1    g10838(.A1(new_n12754_), .A2(new_n3043_), .ZN(new_n13275_));
  AOI21_X1   g10839(.A1(new_n13274_), .A2(new_n13275_), .B(new_n5403_), .ZN(new_n13276_));
  NAND2_X1   g10840(.A1(new_n13169_), .A2(new_n13275_), .ZN(new_n13277_));
  AOI21_X1   g10841(.A1(new_n13260_), .A2(pi1091), .B(new_n5409_), .ZN(new_n13278_));
  NOR2_X1    g10842(.A1(new_n13277_), .A2(new_n13278_), .ZN(new_n13279_));
  NOR2_X1    g10843(.A1(new_n13279_), .A2(new_n5404_), .ZN(new_n13280_));
  NOR2_X1    g10844(.A1(new_n13280_), .A2(new_n13276_), .ZN(new_n13281_));
  NAND2_X1   g10845(.A1(new_n13281_), .A2(new_n5445_), .ZN(new_n13282_));
  AOI21_X1   g10846(.A1(new_n13273_), .A2(new_n13282_), .B(new_n2668_), .ZN(new_n13283_));
  INV_X1     g10847(.I(new_n13265_), .ZN(new_n13284_));
  NOR2_X1    g10848(.A1(new_n13284_), .A2(new_n2642_), .ZN(new_n13285_));
  INV_X1     g10849(.I(new_n13285_), .ZN(new_n13286_));
  INV_X1     g10850(.I(new_n13266_), .ZN(new_n13287_));
  INV_X1     g10851(.I(new_n13267_), .ZN(new_n13288_));
  INV_X1     g10852(.I(new_n13258_), .ZN(new_n13289_));
  INV_X1     g10853(.I(new_n12753_), .ZN(new_n13290_));
  NOR3_X1    g10854(.A1(new_n13081_), .A2(new_n13290_), .A3(new_n13063_), .ZN(new_n13291_));
  OAI21_X1   g10855(.A1(new_n13291_), .A2(new_n5398_), .B(new_n13289_), .ZN(new_n13292_));
  AOI21_X1   g10856(.A1(new_n13292_), .A2(pi0603), .B(new_n13288_), .ZN(new_n13293_));
  NOR3_X1    g10857(.A1(new_n13293_), .A2(new_n5404_), .A3(new_n13287_), .ZN(new_n13294_));
  NOR4_X1    g10858(.A1(new_n2829_), .A2(new_n2830_), .A3(new_n9899_), .A4(new_n13067_), .ZN(new_n13295_));
  NAND2_X1   g10859(.A1(new_n13295_), .A2(pi1092), .ZN(new_n13296_));
  AOI21_X1   g10860(.A1(new_n13296_), .A2(pi0829), .B(new_n6713_), .ZN(new_n13297_));
  OAI21_X1   g10861(.A1(new_n13295_), .A2(new_n13065_), .B(pi1092), .ZN(new_n13298_));
  AOI21_X1   g10862(.A1(new_n9149_), .A2(new_n5392_), .B(pi0824), .ZN(new_n13299_));
  OAI21_X1   g10863(.A1(new_n13299_), .A2(new_n13298_), .B(new_n3044_), .ZN(new_n13300_));
  AOI21_X1   g10864(.A1(new_n13300_), .A2(new_n13297_), .B(new_n13078_), .ZN(new_n13301_));
  OAI21_X1   g10865(.A1(new_n13301_), .A2(new_n3022_), .B(new_n10903_), .ZN(new_n13302_));
  AOI21_X1   g10866(.A1(new_n13302_), .A2(new_n13062_), .B(new_n13073_), .ZN(new_n13303_));
  AOI21_X1   g10867(.A1(new_n13303_), .A2(new_n5437_), .B(new_n13107_), .ZN(new_n13304_));
  NAND2_X1   g10868(.A1(new_n13292_), .A2(pi0603), .ZN(new_n13305_));
  AOI21_X1   g10869(.A1(new_n13305_), .A2(new_n13304_), .B(new_n5403_), .ZN(new_n13306_));
  OAI21_X1   g10870(.A1(new_n13294_), .A2(new_n13306_), .B(new_n5446_), .ZN(new_n13307_));
  INV_X1     g10871(.I(new_n13226_), .ZN(new_n13308_));
  NAND3_X1   g10872(.A1(new_n13302_), .A2(new_n12753_), .A3(new_n13062_), .ZN(new_n13309_));
  NOR2_X1    g10873(.A1(new_n13081_), .A2(new_n13063_), .ZN(new_n13310_));
  AOI21_X1   g10874(.A1(new_n13310_), .A2(new_n12752_), .B(new_n13073_), .ZN(new_n13311_));
  OAI21_X1   g10875(.A1(new_n13311_), .A2(pi0603), .B(new_n13309_), .ZN(new_n13312_));
  INV_X1     g10876(.I(new_n13168_), .ZN(new_n13313_));
  NAND2_X1   g10877(.A1(new_n13313_), .A2(new_n12753_), .ZN(new_n13314_));
  AOI21_X1   g10878(.A1(new_n13291_), .A2(new_n5398_), .B(new_n12751_), .ZN(new_n13315_));
  AOI21_X1   g10879(.A1(new_n13082_), .A2(new_n5398_), .B(new_n13313_), .ZN(new_n13316_));
  AOI22_X1   g10880(.A1(new_n13314_), .A2(new_n13315_), .B1(new_n13316_), .B2(new_n12751_), .ZN(new_n13317_));
  NOR2_X1    g10881(.A1(new_n13317_), .A2(new_n13312_), .ZN(new_n13318_));
  OAI21_X1   g10882(.A1(new_n13318_), .A2(new_n13308_), .B(new_n5445_), .ZN(new_n13319_));
  NAND3_X1   g10883(.A1(new_n13319_), .A2(new_n13307_), .A3(new_n2642_), .ZN(new_n13320_));
  AOI21_X1   g10884(.A1(new_n13320_), .A2(new_n13286_), .B(pi0223), .ZN(new_n13321_));
  OAI21_X1   g10885(.A1(new_n13321_), .A2(new_n13283_), .B(new_n2628_), .ZN(new_n13322_));
  NAND2_X1   g10886(.A1(new_n13272_), .A2(new_n5422_), .ZN(new_n13323_));
  NAND2_X1   g10887(.A1(new_n13281_), .A2(new_n6764_), .ZN(new_n13324_));
  AOI21_X1   g10888(.A1(new_n13323_), .A2(new_n13324_), .B(new_n2436_), .ZN(new_n13325_));
  NOR2_X1    g10889(.A1(new_n13284_), .A2(new_n3304_), .ZN(new_n13326_));
  INV_X1     g10890(.I(new_n13326_), .ZN(new_n13327_));
  OAI21_X1   g10891(.A1(new_n13294_), .A2(new_n13306_), .B(new_n5422_), .ZN(new_n13328_));
  OAI21_X1   g10892(.A1(new_n13318_), .A2(new_n13308_), .B(new_n6764_), .ZN(new_n13329_));
  NAND3_X1   g10893(.A1(new_n13329_), .A2(new_n13328_), .A3(new_n3304_), .ZN(new_n13330_));
  AOI21_X1   g10894(.A1(new_n13330_), .A2(new_n13327_), .B(pi0215), .ZN(new_n13331_));
  OAI21_X1   g10895(.A1(new_n13331_), .A2(new_n13325_), .B(pi0299), .ZN(new_n13332_));
  NAND3_X1   g10896(.A1(new_n13322_), .A2(new_n13332_), .A3(pi0039), .ZN(new_n13333_));
  NAND2_X1   g10897(.A1(new_n13333_), .A2(new_n13257_), .ZN(new_n13334_));
  OAI21_X1   g10898(.A1(new_n13334_), .A2(pi0761), .B(new_n7934_), .ZN(new_n13335_));
  INV_X1     g10899(.I(new_n13061_), .ZN(new_n13336_));
  INV_X1     g10900(.I(new_n13189_), .ZN(new_n13337_));
  AOI21_X1   g10901(.A1(new_n13337_), .A2(new_n13336_), .B(new_n12750_), .ZN(new_n13338_));
  OAI21_X1   g10902(.A1(new_n13335_), .A2(new_n13338_), .B(new_n13246_), .ZN(new_n13339_));
  INV_X1     g10903(.I(new_n12756_), .ZN(new_n13340_));
  NOR2_X1    g10904(.A1(new_n5337_), .A2(new_n13340_), .ZN(new_n13341_));
  INV_X1     g10905(.I(new_n13341_), .ZN(new_n13342_));
  NOR2_X1    g10906(.A1(new_n13342_), .A2(pi0761), .ZN(new_n13343_));
  NOR2_X1    g10907(.A1(new_n5337_), .A2(new_n3043_), .ZN(new_n13344_));
  NOR2_X1    g10908(.A1(new_n13344_), .A2(pi0140), .ZN(new_n13345_));
  OAI21_X1   g10909(.A1(new_n13343_), .A2(new_n13345_), .B(pi0038), .ZN(new_n13346_));
  INV_X1     g10910(.I(new_n13346_), .ZN(new_n13347_));
  AOI21_X1   g10911(.A1(new_n13339_), .A2(new_n3265_), .B(new_n13347_), .ZN(new_n13348_));
  AOI21_X1   g10912(.A1(new_n13348_), .A2(new_n2609_), .B(new_n13197_), .ZN(new_n13349_));
  NOR2_X1    g10913(.A1(new_n13349_), .A2(new_n12760_), .ZN(new_n13350_));
  AOI21_X1   g10914(.A1(new_n12760_), .A2(new_n13196_), .B(new_n13350_), .ZN(new_n13351_));
  NAND2_X1   g10915(.A1(new_n13351_), .A2(new_n12764_), .ZN(new_n13352_));
  NOR2_X1    g10916(.A1(new_n12760_), .A2(pi0609), .ZN(new_n13353_));
  INV_X1     g10917(.I(new_n13353_), .ZN(new_n13354_));
  AOI22_X1   g10918(.A1(new_n13350_), .A2(new_n12766_), .B1(new_n13196_), .B2(new_n13354_), .ZN(new_n13355_));
  NOR2_X1    g10919(.A1(new_n13355_), .A2(pi1155), .ZN(new_n13356_));
  INV_X1     g10920(.I(new_n12772_), .ZN(new_n13357_));
  AOI22_X1   g10921(.A1(new_n13350_), .A2(pi0609), .B1(new_n13357_), .B2(new_n13196_), .ZN(new_n13358_));
  OAI21_X1   g10922(.A1(new_n13358_), .A2(new_n12770_), .B(pi0785), .ZN(new_n13359_));
  OAI21_X1   g10923(.A1(new_n13359_), .A2(new_n13356_), .B(new_n13352_), .ZN(new_n13360_));
  NAND2_X1   g10924(.A1(new_n13360_), .A2(new_n12779_), .ZN(new_n13361_));
  NAND2_X1   g10925(.A1(new_n13196_), .A2(pi0618), .ZN(new_n13362_));
  OAI21_X1   g10926(.A1(new_n13360_), .A2(pi0618), .B(new_n13362_), .ZN(new_n13363_));
  NAND2_X1   g10927(.A1(new_n13363_), .A2(new_n12785_), .ZN(new_n13364_));
  NOR2_X1    g10928(.A1(new_n13360_), .A2(new_n12781_), .ZN(new_n13365_));
  NOR2_X1    g10929(.A1(new_n13194_), .A2(pi0618), .ZN(new_n13366_));
  OAI21_X1   g10930(.A1(new_n13365_), .A2(new_n13366_), .B(pi1154), .ZN(new_n13367_));
  NAND3_X1   g10931(.A1(new_n13367_), .A2(new_n13364_), .A3(pi0781), .ZN(new_n13368_));
  NAND2_X1   g10932(.A1(new_n13368_), .A2(new_n13361_), .ZN(new_n13369_));
  NAND2_X1   g10933(.A1(new_n13196_), .A2(pi0619), .ZN(new_n13370_));
  OAI21_X1   g10934(.A1(new_n13369_), .A2(pi0619), .B(new_n13370_), .ZN(new_n13371_));
  NAND2_X1   g10935(.A1(new_n13371_), .A2(new_n12791_), .ZN(new_n13372_));
  NAND2_X1   g10936(.A1(new_n13196_), .A2(new_n12793_), .ZN(new_n13373_));
  OAI21_X1   g10937(.A1(new_n13369_), .A2(new_n12793_), .B(new_n13373_), .ZN(new_n13374_));
  AOI21_X1   g10938(.A1(new_n13374_), .A2(pi1159), .B(new_n12796_), .ZN(new_n13375_));
  AOI22_X1   g10939(.A1(new_n13375_), .A2(new_n13372_), .B1(new_n12796_), .B2(new_n13369_), .ZN(new_n13376_));
  NOR2_X1    g10940(.A1(new_n13194_), .A2(pi0626), .ZN(new_n13377_));
  AOI21_X1   g10941(.A1(new_n13376_), .A2(pi0626), .B(new_n13377_), .ZN(new_n13378_));
  NOR2_X1    g10942(.A1(new_n13378_), .A2(new_n12745_), .ZN(new_n13379_));
  NOR2_X1    g10943(.A1(new_n13194_), .A2(new_n12747_), .ZN(new_n13380_));
  AOI21_X1   g10944(.A1(new_n13376_), .A2(new_n12747_), .B(new_n13380_), .ZN(new_n13381_));
  OAI21_X1   g10945(.A1(new_n13381_), .A2(pi1158), .B(pi0788), .ZN(new_n13382_));
  OAI22_X1   g10946(.A1(new_n13382_), .A2(new_n13379_), .B1(pi0788), .B2(new_n13376_), .ZN(new_n13383_));
  INV_X1     g10947(.I(new_n12943_), .ZN(new_n13384_));
  NOR2_X1    g10948(.A1(new_n13194_), .A2(new_n13384_), .ZN(new_n13385_));
  INV_X1     g10949(.I(new_n13385_), .ZN(new_n13386_));
  OAI21_X1   g10950(.A1(new_n13383_), .A2(new_n12943_), .B(new_n13386_), .ZN(new_n13387_));
  NAND2_X1   g10951(.A1(new_n13194_), .A2(new_n12984_), .ZN(new_n13388_));
  OAI21_X1   g10952(.A1(new_n13387_), .A2(new_n12984_), .B(new_n13388_), .ZN(new_n13389_));
  NAND2_X1   g10953(.A1(new_n13389_), .A2(new_n12975_), .ZN(new_n13390_));
  AOI21_X1   g10954(.A1(new_n13390_), .A2(new_n13195_), .B(pi1160), .ZN(new_n13391_));
  INV_X1     g10955(.I(new_n12817_), .ZN(new_n13392_));
  NOR2_X1    g10956(.A1(new_n13196_), .A2(new_n12870_), .ZN(new_n13393_));
  INV_X1     g10957(.I(new_n13197_), .ZN(new_n13394_));
  INV_X1     g10958(.I(new_n13191_), .ZN(new_n13395_));
  NAND3_X1   g10959(.A1(new_n13395_), .A2(new_n7934_), .A3(pi0738), .ZN(new_n13396_));
  INV_X1     g10960(.I(new_n13344_), .ZN(new_n13397_));
  NOR2_X1    g10961(.A1(new_n13397_), .A2(new_n12825_), .ZN(new_n13398_));
  NOR2_X1    g10962(.A1(new_n13398_), .A2(new_n3265_), .ZN(new_n13399_));
  OAI21_X1   g10963(.A1(pi0140), .A2(new_n13344_), .B(new_n13399_), .ZN(new_n13400_));
  AOI21_X1   g10964(.A1(new_n13253_), .A2(pi0665), .B(new_n12821_), .ZN(new_n13401_));
  OAI21_X1   g10965(.A1(new_n13401_), .A2(new_n13058_), .B(new_n2628_), .ZN(new_n13402_));
  AOI21_X1   g10966(.A1(new_n13248_), .A2(pi0665), .B(new_n12821_), .ZN(new_n13403_));
  OAI21_X1   g10967(.A1(new_n13403_), .A2(new_n13055_), .B(pi0299), .ZN(new_n13404_));
  NAND2_X1   g10968(.A1(new_n13402_), .A2(new_n13404_), .ZN(new_n13405_));
  INV_X1     g10969(.I(new_n13405_), .ZN(new_n13406_));
  NAND2_X1   g10970(.A1(new_n13406_), .A2(new_n7934_), .ZN(new_n13407_));
  OAI21_X1   g10971(.A1(new_n13053_), .A2(pi0665), .B(new_n13049_), .ZN(new_n13408_));
  NAND3_X1   g10972(.A1(new_n13037_), .A2(new_n13025_), .A3(new_n12822_), .ZN(new_n13409_));
  AOI21_X1   g10973(.A1(new_n13409_), .A2(new_n13039_), .B(pi0210), .ZN(new_n13410_));
  AOI21_X1   g10974(.A1(new_n13408_), .A2(pi0210), .B(new_n13410_), .ZN(new_n13411_));
  NOR2_X1    g10975(.A1(new_n13411_), .A2(new_n2628_), .ZN(new_n13412_));
  AOI21_X1   g10976(.A1(new_n13409_), .A2(new_n13039_), .B(pi0198), .ZN(new_n13413_));
  AOI21_X1   g10977(.A1(new_n13408_), .A2(pi0198), .B(new_n13413_), .ZN(new_n13414_));
  NOR2_X1    g10978(.A1(new_n13414_), .A2(pi0299), .ZN(new_n13415_));
  OAI21_X1   g10979(.A1(new_n13412_), .A2(new_n13415_), .B(pi0680), .ZN(new_n13416_));
  NAND2_X1   g10980(.A1(new_n13416_), .A2(pi0140), .ZN(new_n13417_));
  AOI21_X1   g10981(.A1(new_n13407_), .A2(new_n13417_), .B(pi0039), .ZN(new_n13418_));
  INV_X1     g10982(.I(new_n12823_), .ZN(new_n13419_));
  NAND2_X1   g10983(.A1(new_n13098_), .A2(new_n13419_), .ZN(new_n13420_));
  INV_X1     g10984(.I(new_n13420_), .ZN(new_n13421_));
  AOI21_X1   g10985(.A1(new_n13209_), .A2(new_n13421_), .B(new_n13119_), .ZN(new_n13422_));
  OAI21_X1   g10986(.A1(new_n13209_), .A2(new_n5409_), .B(new_n13421_), .ZN(new_n13423_));
  NOR3_X1    g10987(.A1(new_n13235_), .A2(new_n13423_), .A3(new_n12821_), .ZN(new_n13424_));
  INV_X1     g10988(.I(new_n13424_), .ZN(new_n13425_));
  OR3_X2     g10989(.A1(new_n13425_), .A2(new_n2668_), .A3(new_n13422_), .Z(new_n13426_));
  NOR3_X1    g10990(.A1(new_n13081_), .A2(pi0665), .A3(new_n13063_), .ZN(new_n13427_));
  NOR2_X1    g10991(.A1(new_n13427_), .A2(new_n13073_), .ZN(new_n13428_));
  NOR2_X1    g10992(.A1(new_n13428_), .A2(new_n5403_), .ZN(new_n13429_));
  NOR2_X1    g10993(.A1(new_n13090_), .A2(new_n12825_), .ZN(new_n13430_));
  AOI21_X1   g10994(.A1(new_n13430_), .A2(new_n13119_), .B(new_n13429_), .ZN(new_n13431_));
  AOI21_X1   g10995(.A1(new_n13431_), .A2(new_n5445_), .B(new_n2641_), .ZN(new_n13432_));
  NOR3_X1    g10996(.A1(new_n13427_), .A2(new_n13073_), .A3(new_n13421_), .ZN(new_n13433_));
  OAI21_X1   g10997(.A1(new_n13433_), .A2(new_n13109_), .B(new_n13118_), .ZN(new_n13434_));
  NAND2_X1   g10998(.A1(new_n13434_), .A2(pi0680), .ZN(new_n13435_));
  OAI21_X1   g10999(.A1(new_n13433_), .A2(new_n13109_), .B(new_n5410_), .ZN(new_n13436_));
  NAND2_X1   g11000(.A1(new_n13420_), .A2(new_n5409_), .ZN(new_n13437_));
  AOI21_X1   g11001(.A1(new_n13436_), .A2(new_n13437_), .B(new_n13118_), .ZN(new_n13438_));
  OAI21_X1   g11002(.A1(new_n13438_), .A2(new_n13435_), .B(new_n5446_), .ZN(new_n13439_));
  AOI22_X1   g11003(.A1(new_n13439_), .A2(new_n13432_), .B1(new_n12824_), .B2(new_n13185_), .ZN(new_n13440_));
  OAI21_X1   g11004(.A1(new_n13440_), .A2(pi0223), .B(new_n13426_), .ZN(new_n13441_));
  NAND2_X1   g11005(.A1(new_n13441_), .A2(new_n2628_), .ZN(new_n13442_));
  NOR3_X1    g11006(.A1(new_n13218_), .A2(new_n13423_), .A3(new_n12821_), .ZN(new_n13443_));
  INV_X1     g11007(.I(new_n13443_), .ZN(new_n13444_));
  NOR3_X1    g11008(.A1(new_n13444_), .A2(new_n2436_), .A3(new_n13422_), .ZN(new_n13445_));
  NOR2_X1    g11009(.A1(new_n13088_), .A2(new_n12825_), .ZN(new_n13446_));
  NAND2_X1   g11010(.A1(new_n13446_), .A2(new_n3303_), .ZN(new_n13447_));
  NAND2_X1   g11011(.A1(new_n13431_), .A2(new_n6764_), .ZN(new_n13448_));
  OAI21_X1   g11012(.A1(new_n13438_), .A2(new_n13435_), .B(new_n5422_), .ZN(new_n13449_));
  NAND3_X1   g11013(.A1(new_n13449_), .A2(new_n3304_), .A3(new_n13448_), .ZN(new_n13450_));
  AOI21_X1   g11014(.A1(new_n13450_), .A2(new_n13447_), .B(pi0215), .ZN(new_n13451_));
  OAI21_X1   g11015(.A1(new_n13451_), .A2(new_n13445_), .B(pi0299), .ZN(new_n13452_));
  NAND3_X1   g11016(.A1(new_n13442_), .A2(new_n13452_), .A3(pi0140), .ZN(new_n13453_));
  NAND2_X1   g11017(.A1(new_n13098_), .A2(new_n12823_), .ZN(new_n13454_));
  OAI21_X1   g11018(.A1(new_n13454_), .A2(new_n5410_), .B(pi0680), .ZN(new_n13455_));
  NAND2_X1   g11019(.A1(new_n13454_), .A2(new_n5398_), .ZN(new_n13456_));
  NAND3_X1   g11020(.A1(new_n13260_), .A2(pi0665), .A3(pi1091), .ZN(new_n13457_));
  INV_X1     g11021(.I(new_n13457_), .ZN(new_n13458_));
  OAI21_X1   g11022(.A1(new_n5398_), .A2(new_n13458_), .B(new_n13456_), .ZN(new_n13459_));
  INV_X1     g11023(.I(new_n13459_), .ZN(new_n13460_));
  AOI21_X1   g11024(.A1(new_n5403_), .A2(new_n13455_), .B(new_n13460_), .ZN(new_n13461_));
  NOR2_X1    g11025(.A1(new_n13168_), .A2(new_n13419_), .ZN(new_n13462_));
  NAND2_X1   g11026(.A1(new_n13462_), .A2(new_n5409_), .ZN(new_n13463_));
  NAND3_X1   g11027(.A1(new_n13463_), .A2(pi0680), .A3(new_n13457_), .ZN(new_n13464_));
  NAND2_X1   g11028(.A1(new_n13167_), .A2(new_n13111_), .ZN(new_n13465_));
  NAND2_X1   g11029(.A1(new_n13465_), .A2(new_n13169_), .ZN(new_n13466_));
  NAND2_X1   g11030(.A1(new_n13466_), .A2(new_n12821_), .ZN(new_n13467_));
  NAND2_X1   g11031(.A1(new_n13467_), .A2(new_n13464_), .ZN(new_n13468_));
  NOR2_X1    g11032(.A1(new_n13468_), .A2(new_n13461_), .ZN(new_n13469_));
  NOR2_X1    g11033(.A1(new_n13469_), .A2(new_n5446_), .ZN(new_n13470_));
  INV_X1     g11034(.I(new_n13461_), .ZN(new_n13471_));
  NAND2_X1   g11035(.A1(new_n13143_), .A2(new_n12821_), .ZN(new_n13472_));
  NAND2_X1   g11036(.A1(new_n13471_), .A2(new_n13472_), .ZN(new_n13473_));
  NAND2_X1   g11037(.A1(new_n13473_), .A2(new_n5446_), .ZN(new_n13474_));
  INV_X1     g11038(.I(new_n13474_), .ZN(new_n13475_));
  OAI21_X1   g11039(.A1(new_n13470_), .A2(new_n13475_), .B(pi0223), .ZN(new_n13476_));
  INV_X1     g11040(.I(new_n13476_), .ZN(new_n13477_));
  NOR3_X1    g11041(.A1(new_n13081_), .A2(new_n13419_), .A3(new_n13063_), .ZN(new_n13478_));
  INV_X1     g11042(.I(new_n13478_), .ZN(new_n13479_));
  NAND2_X1   g11043(.A1(new_n13479_), .A2(new_n13118_), .ZN(new_n13480_));
  AOI22_X1   g11044(.A1(new_n13478_), .A2(new_n5691_), .B1(new_n5409_), .B2(new_n13462_), .ZN(new_n13481_));
  NAND2_X1   g11045(.A1(new_n13481_), .A2(new_n13119_), .ZN(new_n13482_));
  AOI21_X1   g11046(.A1(new_n13482_), .A2(new_n13480_), .B(new_n12821_), .ZN(new_n13483_));
  INV_X1     g11047(.I(new_n13089_), .ZN(new_n13484_));
  OAI21_X1   g11048(.A1(new_n13303_), .A2(new_n5724_), .B(new_n13484_), .ZN(new_n13485_));
  NOR2_X1    g11049(.A1(new_n13485_), .A2(pi0680), .ZN(new_n13486_));
  OR2_X2     g11050(.A1(new_n13483_), .A2(new_n13486_), .Z(new_n13487_));
  AOI21_X1   g11051(.A1(new_n13487_), .A2(new_n5445_), .B(new_n2641_), .ZN(new_n13488_));
  NOR3_X1    g11052(.A1(new_n13103_), .A2(pi0680), .A3(new_n13105_), .ZN(new_n13489_));
  INV_X1     g11053(.I(new_n13456_), .ZN(new_n13490_));
  NOR2_X1    g11054(.A1(new_n13478_), .A2(new_n5398_), .ZN(new_n13491_));
  NOR2_X1    g11055(.A1(new_n13491_), .A2(new_n13490_), .ZN(new_n13492_));
  NOR2_X1    g11056(.A1(new_n13492_), .A2(new_n12821_), .ZN(new_n13493_));
  OR3_X2     g11057(.A1(new_n13489_), .A2(new_n13119_), .A3(new_n13493_), .Z(new_n13494_));
  AOI21_X1   g11058(.A1(new_n13492_), .A2(new_n5410_), .B(new_n13455_), .ZN(new_n13495_));
  NOR2_X1    g11059(.A1(new_n13489_), .A2(new_n13495_), .ZN(new_n13496_));
  NAND2_X1   g11060(.A1(new_n13496_), .A2(new_n13119_), .ZN(new_n13497_));
  NAND3_X1   g11061(.A1(new_n13497_), .A2(new_n13494_), .A3(new_n5446_), .ZN(new_n13498_));
  AOI21_X1   g11062(.A1(new_n13185_), .A2(new_n12825_), .B(pi0223), .ZN(new_n13499_));
  INV_X1     g11063(.I(new_n13499_), .ZN(new_n13500_));
  AOI21_X1   g11064(.A1(new_n13498_), .A2(new_n13488_), .B(new_n13500_), .ZN(new_n13501_));
  OAI21_X1   g11065(.A1(new_n13477_), .A2(new_n13501_), .B(new_n2628_), .ZN(new_n13502_));
  NOR2_X1    g11066(.A1(new_n13469_), .A2(new_n5422_), .ZN(new_n13503_));
  NAND2_X1   g11067(.A1(new_n13473_), .A2(new_n5422_), .ZN(new_n13504_));
  INV_X1     g11068(.I(new_n13504_), .ZN(new_n13505_));
  OAI21_X1   g11069(.A1(new_n13503_), .A2(new_n13505_), .B(pi0215), .ZN(new_n13506_));
  INV_X1     g11070(.I(new_n13506_), .ZN(new_n13507_));
  AOI21_X1   g11071(.A1(new_n13487_), .A2(new_n6764_), .B(new_n3303_), .ZN(new_n13508_));
  NAND3_X1   g11072(.A1(new_n13497_), .A2(new_n13494_), .A3(new_n5422_), .ZN(new_n13509_));
  NOR2_X1    g11073(.A1(new_n12824_), .A2(new_n3043_), .ZN(new_n13510_));
  AOI21_X1   g11074(.A1(new_n13222_), .A2(new_n13510_), .B(pi0215), .ZN(new_n13511_));
  INV_X1     g11075(.I(new_n13511_), .ZN(new_n13512_));
  AOI21_X1   g11076(.A1(new_n13509_), .A2(new_n13508_), .B(new_n13512_), .ZN(new_n13513_));
  OAI21_X1   g11077(.A1(new_n13507_), .A2(new_n13513_), .B(pi0299), .ZN(new_n13514_));
  NAND3_X1   g11078(.A1(new_n13502_), .A2(new_n13514_), .A3(new_n7934_), .ZN(new_n13515_));
  AOI21_X1   g11079(.A1(new_n13515_), .A2(new_n13453_), .B(new_n2627_), .ZN(new_n13516_));
  OAI21_X1   g11080(.A1(new_n13516_), .A2(new_n13418_), .B(new_n3265_), .ZN(new_n13517_));
  NAND3_X1   g11081(.A1(new_n13517_), .A2(new_n12820_), .A3(new_n13400_), .ZN(new_n13518_));
  NAND3_X1   g11082(.A1(new_n13518_), .A2(new_n13396_), .A3(new_n2609_), .ZN(new_n13519_));
  NAND2_X1   g11083(.A1(new_n13519_), .A2(new_n13394_), .ZN(new_n13520_));
  INV_X1     g11084(.I(pi0625), .ZN(new_n13521_));
  NAND2_X1   g11085(.A1(new_n13520_), .A2(new_n13521_), .ZN(new_n13522_));
  NAND2_X1   g11086(.A1(new_n13196_), .A2(pi0625), .ZN(new_n13523_));
  AOI21_X1   g11087(.A1(new_n13522_), .A2(new_n13523_), .B(pi1153), .ZN(new_n13524_));
  AOI21_X1   g11088(.A1(new_n13519_), .A2(new_n13394_), .B(new_n13521_), .ZN(new_n13525_));
  NOR2_X1    g11089(.A1(new_n13194_), .A2(pi0625), .ZN(new_n13526_));
  OAI21_X1   g11090(.A1(new_n13525_), .A2(new_n13526_), .B(pi1153), .ZN(new_n13527_));
  NAND2_X1   g11091(.A1(new_n13527_), .A2(pi0778), .ZN(new_n13528_));
  OAI22_X1   g11092(.A1(new_n13528_), .A2(new_n13524_), .B1(pi0778), .B2(new_n13520_), .ZN(new_n13529_));
  AOI21_X1   g11093(.A1(new_n13529_), .A2(new_n12870_), .B(new_n13393_), .ZN(new_n13530_));
  NOR2_X1    g11094(.A1(new_n13194_), .A2(new_n12888_), .ZN(new_n13531_));
  AOI21_X1   g11095(.A1(new_n13530_), .A2(new_n12888_), .B(new_n13531_), .ZN(new_n13532_));
  NOR2_X1    g11096(.A1(new_n13196_), .A2(new_n12911_), .ZN(new_n13533_));
  AOI21_X1   g11097(.A1(new_n13532_), .A2(new_n12911_), .B(new_n13533_), .ZN(new_n13534_));
  NAND2_X1   g11098(.A1(new_n13534_), .A2(new_n13392_), .ZN(new_n13535_));
  OAI21_X1   g11099(.A1(new_n13392_), .A2(new_n13194_), .B(new_n13535_), .ZN(new_n13536_));
  NAND2_X1   g11100(.A1(new_n13536_), .A2(new_n12920_), .ZN(new_n13537_));
  NAND2_X1   g11101(.A1(new_n13196_), .A2(pi0628), .ZN(new_n13538_));
  AOI21_X1   g11102(.A1(new_n13537_), .A2(new_n13538_), .B(pi1156), .ZN(new_n13539_));
  NAND2_X1   g11103(.A1(new_n13196_), .A2(new_n12920_), .ZN(new_n13540_));
  NAND2_X1   g11104(.A1(new_n13536_), .A2(pi0628), .ZN(new_n13541_));
  AOI21_X1   g11105(.A1(new_n13541_), .A2(new_n13540_), .B(new_n12742_), .ZN(new_n13542_));
  NOR3_X1    g11106(.A1(new_n13539_), .A2(new_n13542_), .A3(new_n12937_), .ZN(new_n13543_));
  NOR2_X1    g11107(.A1(new_n13536_), .A2(pi0792), .ZN(new_n13544_));
  NOR2_X1    g11108(.A1(new_n13543_), .A2(new_n13544_), .ZN(new_n13545_));
  NAND2_X1   g11109(.A1(new_n13545_), .A2(new_n12741_), .ZN(new_n13546_));
  NAND2_X1   g11110(.A1(new_n13196_), .A2(pi0647), .ZN(new_n13547_));
  AOI21_X1   g11111(.A1(new_n13546_), .A2(new_n13547_), .B(pi1157), .ZN(new_n13548_));
  NAND2_X1   g11112(.A1(new_n13545_), .A2(pi0647), .ZN(new_n13549_));
  OAI21_X1   g11113(.A1(pi0647), .A2(new_n13194_), .B(new_n13549_), .ZN(new_n13550_));
  NAND2_X1   g11114(.A1(new_n13550_), .A2(pi1157), .ZN(new_n13551_));
  NAND2_X1   g11115(.A1(new_n13551_), .A2(pi0787), .ZN(new_n13552_));
  OAI22_X1   g11116(.A1(new_n13552_), .A2(new_n13548_), .B1(pi0787), .B2(new_n13545_), .ZN(new_n13553_));
  AOI21_X1   g11117(.A1(new_n13553_), .A2(pi0644), .B(pi0715), .ZN(new_n13554_));
  NOR2_X1    g11118(.A1(new_n13539_), .A2(new_n12919_), .ZN(new_n13555_));
  AOI21_X1   g11119(.A1(new_n13383_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n13556_));
  INV_X1     g11120(.I(new_n12902_), .ZN(new_n13557_));
  OAI21_X1   g11121(.A1(new_n13378_), .A2(new_n12745_), .B(new_n13557_), .ZN(new_n13558_));
  AOI21_X1   g11122(.A1(new_n13534_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n13559_));
  INV_X1     g11123(.I(pi0608), .ZN(new_n13560_));
  NOR2_X1    g11124(.A1(new_n2627_), .A2(pi0140), .ZN(new_n13561_));
  NOR2_X1    g11125(.A1(new_n12832_), .A2(new_n12754_), .ZN(new_n13562_));
  NOR2_X1    g11126(.A1(new_n13562_), .A2(new_n12756_), .ZN(new_n13563_));
  NAND2_X1   g11127(.A1(new_n2531_), .A2(pi0140), .ZN(new_n13564_));
  OAI21_X1   g11128(.A1(new_n13564_), .A2(new_n13563_), .B(new_n12750_), .ZN(new_n13565_));
  NAND3_X1   g11129(.A1(new_n13136_), .A2(new_n12755_), .A3(new_n12825_), .ZN(new_n13566_));
  AOI21_X1   g11130(.A1(new_n7934_), .A2(new_n13566_), .B(new_n13565_), .ZN(new_n13567_));
  INV_X1     g11131(.I(new_n13136_), .ZN(new_n13568_));
  NOR2_X1    g11132(.A1(new_n12754_), .A2(new_n12823_), .ZN(new_n13569_));
  INV_X1     g11133(.I(new_n13569_), .ZN(new_n13570_));
  NOR2_X1    g11134(.A1(new_n13570_), .A2(new_n12821_), .ZN(new_n13571_));
  INV_X1     g11135(.I(new_n13571_), .ZN(new_n13572_));
  NOR2_X1    g11136(.A1(new_n13568_), .A2(new_n13572_), .ZN(new_n13573_));
  OAI21_X1   g11137(.A1(new_n13136_), .A2(pi0140), .B(pi0761), .ZN(new_n13574_));
  NOR2_X1    g11138(.A1(new_n13573_), .A2(new_n13574_), .ZN(new_n13575_));
  NOR3_X1    g11139(.A1(new_n13567_), .A2(pi0039), .A3(new_n13575_), .ZN(new_n13576_));
  OAI21_X1   g11140(.A1(new_n13576_), .A2(new_n13561_), .B(pi0038), .ZN(new_n13577_));
  NOR2_X1    g11141(.A1(new_n13170_), .A2(new_n13420_), .ZN(new_n13578_));
  INV_X1     g11142(.I(new_n13578_), .ZN(new_n13579_));
  NOR4_X1    g11143(.A1(new_n13579_), .A2(new_n13422_), .A3(new_n13423_), .A4(new_n12821_), .ZN(new_n13580_));
  OAI21_X1   g11144(.A1(new_n13149_), .A2(new_n13214_), .B(new_n13216_), .ZN(new_n13581_));
  NOR2_X1    g11145(.A1(new_n13581_), .A2(new_n13580_), .ZN(new_n13582_));
  AOI21_X1   g11146(.A1(new_n13582_), .A2(new_n5445_), .B(new_n2668_), .ZN(new_n13583_));
  NOR2_X1    g11147(.A1(new_n13118_), .A2(new_n12821_), .ZN(new_n13584_));
  INV_X1     g11148(.I(new_n13584_), .ZN(new_n13585_));
  NOR2_X1    g11149(.A1(new_n12751_), .A2(pi0621), .ZN(new_n13586_));
  NOR2_X1    g11150(.A1(new_n13419_), .A2(new_n13586_), .ZN(new_n13587_));
  NOR2_X1    g11151(.A1(new_n13088_), .A2(new_n13587_), .ZN(new_n13588_));
  AOI21_X1   g11152(.A1(new_n13588_), .A2(new_n13264_), .B(new_n13585_), .ZN(new_n13589_));
  INV_X1     g11153(.I(new_n13589_), .ZN(new_n13590_));
  AOI21_X1   g11154(.A1(new_n13423_), .A2(new_n13211_), .B(new_n13264_), .ZN(new_n13591_));
  NOR2_X1    g11155(.A1(new_n13422_), .A2(new_n12821_), .ZN(new_n13592_));
  OAI22_X1   g11156(.A1(new_n13217_), .A2(new_n13592_), .B1(new_n13590_), .B2(new_n13591_), .ZN(new_n13593_));
  NAND2_X1   g11157(.A1(new_n13593_), .A2(new_n5446_), .ZN(new_n13594_));
  AOI21_X1   g11158(.A1(new_n13583_), .A2(new_n13594_), .B(pi0299), .ZN(new_n13595_));
  INV_X1     g11159(.I(new_n13595_), .ZN(new_n13596_));
  INV_X1     g11160(.I(new_n13563_), .ZN(new_n13597_));
  AOI21_X1   g11161(.A1(new_n13098_), .A2(new_n13597_), .B(new_n2642_), .ZN(new_n13598_));
  NOR2_X1    g11162(.A1(new_n13598_), .A2(pi0223), .ZN(new_n13599_));
  NAND2_X1   g11163(.A1(new_n13485_), .A2(new_n5403_), .ZN(new_n13600_));
  AOI21_X1   g11164(.A1(new_n13600_), .A2(new_n13225_), .B(new_n12755_), .ZN(new_n13601_));
  NOR3_X1    g11165(.A1(new_n13601_), .A2(new_n13429_), .A3(new_n13584_), .ZN(new_n13602_));
  OAI21_X1   g11166(.A1(new_n13303_), .A2(new_n5437_), .B(new_n13168_), .ZN(new_n13603_));
  NAND3_X1   g11167(.A1(new_n13302_), .A2(new_n12822_), .A3(new_n13062_), .ZN(new_n13604_));
  NAND3_X1   g11168(.A1(new_n13604_), .A2(new_n13074_), .A3(new_n13420_), .ZN(new_n13605_));
  AOI21_X1   g11169(.A1(new_n13603_), .A2(new_n13605_), .B(pi0603), .ZN(new_n13606_));
  NOR2_X1    g11170(.A1(new_n13073_), .A2(new_n12752_), .ZN(new_n13607_));
  NOR2_X1    g11171(.A1(new_n13303_), .A2(new_n13607_), .ZN(new_n13608_));
  OAI21_X1   g11172(.A1(new_n13309_), .A2(pi0665), .B(pi0603), .ZN(new_n13609_));
  NOR2_X1    g11173(.A1(new_n13609_), .A2(new_n13608_), .ZN(new_n13610_));
  OAI21_X1   g11174(.A1(new_n13606_), .A2(new_n13610_), .B(new_n5408_), .ZN(new_n13611_));
  NOR2_X1    g11175(.A1(new_n13605_), .A2(new_n12754_), .ZN(new_n13612_));
  OAI21_X1   g11176(.A1(new_n13612_), .A2(new_n13316_), .B(new_n13264_), .ZN(new_n13613_));
  AOI21_X1   g11177(.A1(new_n13611_), .A2(new_n13613_), .B(new_n13585_), .ZN(new_n13614_));
  NOR2_X1    g11178(.A1(new_n13614_), .A2(new_n13602_), .ZN(new_n13615_));
  NAND2_X1   g11179(.A1(new_n13615_), .A2(new_n5445_), .ZN(new_n13616_));
  NAND2_X1   g11180(.A1(new_n13433_), .A2(new_n12755_), .ZN(new_n13617_));
  AOI21_X1   g11181(.A1(new_n13617_), .A2(new_n13304_), .B(new_n5403_), .ZN(new_n13618_));
  INV_X1     g11182(.I(new_n13618_), .ZN(new_n13619_));
  OAI21_X1   g11183(.A1(new_n13109_), .A2(new_n12755_), .B(new_n5408_), .ZN(new_n13620_));
  NOR2_X1    g11184(.A1(new_n13210_), .A2(new_n5408_), .ZN(new_n13621_));
  INV_X1     g11185(.I(new_n13621_), .ZN(new_n13622_));
  AOI21_X1   g11186(.A1(new_n13620_), .A2(new_n13622_), .B(pi0680), .ZN(new_n13623_));
  INV_X1     g11187(.I(new_n13623_), .ZN(new_n13624_));
  NOR2_X1    g11188(.A1(new_n12751_), .A2(pi0665), .ZN(new_n13625_));
  INV_X1     g11189(.I(new_n13625_), .ZN(new_n13626_));
  OAI21_X1   g11190(.A1(new_n13420_), .A2(pi0603), .B(new_n13626_), .ZN(new_n13627_));
  INV_X1     g11191(.I(new_n13627_), .ZN(new_n13628_));
  AOI21_X1   g11192(.A1(new_n13292_), .A2(pi0603), .B(new_n13628_), .ZN(new_n13629_));
  OAI21_X1   g11193(.A1(new_n13629_), .A2(new_n13228_), .B(new_n5408_), .ZN(new_n13630_));
  NAND2_X1   g11194(.A1(new_n13630_), .A2(new_n13589_), .ZN(new_n13631_));
  NAND4_X1   g11195(.A1(new_n13631_), .A2(new_n13624_), .A3(new_n13619_), .A4(new_n5446_), .ZN(new_n13632_));
  NAND3_X1   g11196(.A1(new_n13616_), .A2(new_n2642_), .A3(new_n13632_), .ZN(new_n13633_));
  AOI21_X1   g11197(.A1(new_n13633_), .A2(new_n13599_), .B(new_n13596_), .ZN(new_n13634_));
  NAND2_X1   g11198(.A1(new_n13593_), .A2(new_n5422_), .ZN(new_n13635_));
  NAND2_X1   g11199(.A1(new_n13582_), .A2(new_n6764_), .ZN(new_n13636_));
  AOI21_X1   g11200(.A1(new_n13636_), .A2(new_n13635_), .B(new_n2436_), .ZN(new_n13637_));
  INV_X1     g11201(.I(new_n13637_), .ZN(new_n13638_));
  NOR2_X1    g11202(.A1(new_n13088_), .A2(new_n3304_), .ZN(new_n13639_));
  AOI21_X1   g11203(.A1(new_n13639_), .A2(new_n13597_), .B(pi0215), .ZN(new_n13640_));
  NAND2_X1   g11204(.A1(new_n13303_), .A2(new_n5437_), .ZN(new_n13641_));
  NAND3_X1   g11205(.A1(new_n13641_), .A2(new_n12754_), .A3(new_n13108_), .ZN(new_n13642_));
  AOI21_X1   g11206(.A1(new_n13309_), .A2(new_n5437_), .B(new_n13258_), .ZN(new_n13643_));
  OAI21_X1   g11207(.A1(new_n13643_), .A2(new_n12751_), .B(new_n13627_), .ZN(new_n13644_));
  NAND2_X1   g11208(.A1(new_n13644_), .A2(new_n13642_), .ZN(new_n13645_));
  AOI21_X1   g11209(.A1(new_n13645_), .A2(new_n5408_), .B(new_n13590_), .ZN(new_n13646_));
  NOR4_X1    g11210(.A1(new_n13646_), .A2(new_n6764_), .A3(new_n13618_), .A4(new_n13623_), .ZN(new_n13647_));
  NOR3_X1    g11211(.A1(new_n13614_), .A2(new_n5422_), .A3(new_n13602_), .ZN(new_n13648_));
  OAI21_X1   g11212(.A1(new_n13648_), .A2(new_n13647_), .B(new_n3304_), .ZN(new_n13649_));
  NAND2_X1   g11213(.A1(new_n13649_), .A2(new_n13640_), .ZN(new_n13650_));
  AOI21_X1   g11214(.A1(new_n13650_), .A2(new_n13638_), .B(new_n2628_), .ZN(new_n13651_));
  OAI21_X1   g11215(.A1(new_n13651_), .A2(new_n13634_), .B(pi0140), .ZN(new_n13652_));
  INV_X1     g11216(.I(new_n13462_), .ZN(new_n13653_));
  NAND2_X1   g11217(.A1(new_n13653_), .A2(new_n13457_), .ZN(new_n13654_));
  AOI21_X1   g11218(.A1(new_n13269_), .A2(new_n13654_), .B(new_n13585_), .ZN(new_n13655_));
  AOI21_X1   g11219(.A1(new_n13457_), .A2(pi0680), .B(new_n13586_), .ZN(new_n13656_));
  OAI22_X1   g11220(.A1(new_n13279_), .A2(pi0680), .B1(new_n5403_), .B2(new_n13656_), .ZN(new_n13657_));
  OAI21_X1   g11221(.A1(new_n13655_), .A2(new_n13657_), .B(new_n5445_), .ZN(new_n13658_));
  INV_X1     g11222(.I(new_n13586_), .ZN(new_n13659_));
  NAND3_X1   g11223(.A1(new_n13460_), .A2(new_n5404_), .A3(new_n13659_), .ZN(new_n13660_));
  NAND3_X1   g11224(.A1(new_n13269_), .A2(new_n5403_), .A3(new_n12825_), .ZN(new_n13661_));
  NAND3_X1   g11225(.A1(new_n13661_), .A2(new_n5446_), .A3(new_n13660_), .ZN(new_n13662_));
  AOI21_X1   g11226(.A1(new_n13658_), .A2(new_n13662_), .B(new_n2668_), .ZN(new_n13663_));
  NOR3_X1    g11227(.A1(new_n13293_), .A2(pi0680), .A3(new_n13287_), .ZN(new_n13664_));
  NOR2_X1    g11228(.A1(new_n13454_), .A2(new_n13586_), .ZN(new_n13665_));
  AOI21_X1   g11229(.A1(new_n13665_), .A2(new_n13264_), .B(new_n13585_), .ZN(new_n13666_));
  INV_X1     g11230(.I(new_n13666_), .ZN(new_n13667_));
  AOI21_X1   g11231(.A1(new_n13293_), .A2(new_n12823_), .B(new_n13667_), .ZN(new_n13668_));
  AOI21_X1   g11232(.A1(new_n13492_), .A2(new_n13587_), .B(new_n5403_), .ZN(new_n13669_));
  NOR4_X1    g11233(.A1(new_n13664_), .A2(new_n13668_), .A3(new_n5445_), .A4(new_n13669_), .ZN(new_n13670_));
  OAI21_X1   g11234(.A1(new_n13479_), .A2(new_n13586_), .B(new_n5404_), .ZN(new_n13671_));
  INV_X1     g11235(.I(new_n13587_), .ZN(new_n13672_));
  OAI21_X1   g11236(.A1(new_n13481_), .A2(new_n13672_), .B(new_n13584_), .ZN(new_n13673_));
  NAND2_X1   g11237(.A1(new_n13673_), .A2(new_n13671_), .ZN(new_n13674_));
  AOI21_X1   g11238(.A1(new_n13485_), .A2(new_n12755_), .B(pi0680), .ZN(new_n13675_));
  NOR3_X1    g11239(.A1(new_n13674_), .A2(new_n5446_), .A3(new_n13675_), .ZN(new_n13676_));
  OAI21_X1   g11240(.A1(new_n13670_), .A2(new_n13676_), .B(new_n2642_), .ZN(new_n13677_));
  NOR2_X1    g11241(.A1(new_n13085_), .A2(pi0120), .ZN(new_n13678_));
  INV_X1     g11242(.I(new_n13678_), .ZN(new_n13679_));
  NOR2_X1    g11243(.A1(new_n13566_), .A2(new_n2642_), .ZN(new_n13680_));
  AOI21_X1   g11244(.A1(new_n13680_), .A2(new_n13679_), .B(pi0223), .ZN(new_n13681_));
  AOI21_X1   g11245(.A1(new_n13677_), .A2(new_n13681_), .B(new_n13663_), .ZN(new_n13682_));
  OAI21_X1   g11246(.A1(new_n13655_), .A2(new_n13657_), .B(new_n6764_), .ZN(new_n13683_));
  NAND3_X1   g11247(.A1(new_n13661_), .A2(new_n5422_), .A3(new_n13660_), .ZN(new_n13684_));
  AOI21_X1   g11248(.A1(new_n13683_), .A2(new_n13684_), .B(new_n2436_), .ZN(new_n13685_));
  NOR4_X1    g11249(.A1(new_n13664_), .A2(new_n13668_), .A3(new_n6764_), .A4(new_n13669_), .ZN(new_n13686_));
  NOR3_X1    g11250(.A1(new_n13674_), .A2(new_n5422_), .A3(new_n13675_), .ZN(new_n13687_));
  OAI21_X1   g11251(.A1(new_n13686_), .A2(new_n13687_), .B(new_n3304_), .ZN(new_n13688_));
  NOR2_X1    g11252(.A1(new_n13566_), .A2(new_n3304_), .ZN(new_n13689_));
  AOI21_X1   g11253(.A1(new_n13689_), .A2(new_n13679_), .B(pi0215), .ZN(new_n13690_));
  AOI21_X1   g11254(.A1(new_n13688_), .A2(new_n13690_), .B(new_n13685_), .ZN(new_n13691_));
  MUX2_X1    g11255(.I0(new_n13691_), .I1(new_n13682_), .S(new_n2628_), .Z(new_n13692_));
  NAND2_X1   g11256(.A1(new_n13692_), .A2(new_n7934_), .ZN(new_n13693_));
  AOI21_X1   g11257(.A1(new_n13652_), .A2(new_n13693_), .B(pi0761), .ZN(new_n13694_));
  NAND3_X1   g11258(.A1(new_n13459_), .A2(new_n5404_), .A3(new_n13211_), .ZN(new_n13695_));
  NAND2_X1   g11259(.A1(new_n13695_), .A2(new_n13472_), .ZN(new_n13696_));
  NAND2_X1   g11260(.A1(new_n13098_), .A2(new_n13570_), .ZN(new_n13697_));
  INV_X1     g11261(.I(new_n13697_), .ZN(new_n13698_));
  NOR2_X1    g11262(.A1(new_n13698_), .A2(new_n13111_), .ZN(new_n13699_));
  INV_X1     g11263(.I(new_n13699_), .ZN(new_n13700_));
  NOR2_X1    g11264(.A1(new_n13698_), .A2(new_n5405_), .ZN(new_n13701_));
  NAND2_X1   g11265(.A1(new_n13697_), .A2(pi0642), .ZN(new_n13702_));
  NOR2_X1    g11266(.A1(new_n13149_), .A2(new_n13214_), .ZN(new_n13703_));
  NOR3_X1    g11267(.A1(new_n13168_), .A2(pi0603), .A3(new_n13419_), .ZN(new_n13704_));
  NOR3_X1    g11268(.A1(new_n13704_), .A2(new_n13703_), .A3(new_n13458_), .ZN(new_n13705_));
  NAND4_X1   g11269(.A1(new_n13705_), .A2(new_n13459_), .A3(new_n5406_), .A4(new_n13211_), .ZN(new_n13706_));
  AOI21_X1   g11270(.A1(new_n13706_), .A2(new_n13702_), .B(pi0614), .ZN(new_n13707_));
  OAI21_X1   g11271(.A1(new_n13707_), .A2(new_n13701_), .B(new_n13111_), .ZN(new_n13708_));
  AOI21_X1   g11272(.A1(new_n13708_), .A2(new_n13700_), .B(new_n13585_), .ZN(new_n13709_));
  NOR3_X1    g11273(.A1(new_n13709_), .A2(new_n5445_), .A3(new_n13696_), .ZN(new_n13710_));
  INV_X1     g11274(.I(new_n13467_), .ZN(new_n13711_));
  NOR2_X1    g11275(.A1(new_n13703_), .A2(new_n13458_), .ZN(new_n13712_));
  INV_X1     g11276(.I(new_n13712_), .ZN(new_n13713_));
  NOR3_X1    g11277(.A1(new_n13713_), .A2(new_n13264_), .A3(new_n13704_), .ZN(new_n13714_));
  NOR3_X1    g11278(.A1(new_n13215_), .A2(new_n5408_), .A3(new_n13654_), .ZN(new_n13715_));
  NOR2_X1    g11279(.A1(new_n13715_), .A2(new_n13714_), .ZN(new_n13716_));
  NOR2_X1    g11280(.A1(new_n13716_), .A2(new_n13585_), .ZN(new_n13717_));
  NOR2_X1    g11281(.A1(new_n13713_), .A2(new_n5403_), .ZN(new_n13718_));
  NOR4_X1    g11282(.A1(new_n13717_), .A2(new_n13711_), .A3(new_n5446_), .A4(new_n13718_), .ZN(new_n13719_));
  OAI21_X1   g11283(.A1(new_n13710_), .A2(new_n13719_), .B(pi0223), .ZN(new_n13720_));
  NOR3_X1    g11284(.A1(new_n13303_), .A2(new_n12751_), .A3(new_n13607_), .ZN(new_n13721_));
  NOR2_X1    g11285(.A1(new_n13671_), .A2(new_n13721_), .ZN(new_n13722_));
  AOI21_X1   g11286(.A1(new_n13485_), .A2(new_n13570_), .B(new_n13585_), .ZN(new_n13723_));
  NOR3_X1    g11287(.A1(new_n13722_), .A2(new_n13723_), .A3(new_n13486_), .ZN(new_n13724_));
  INV_X1     g11288(.I(new_n13724_), .ZN(new_n13725_));
  OAI21_X1   g11289(.A1(new_n13725_), .A2(new_n5446_), .B(new_n2642_), .ZN(new_n13726_));
  NAND2_X1   g11290(.A1(new_n13098_), .A2(pi0642), .ZN(new_n13727_));
  NOR2_X1    g11291(.A1(new_n5398_), .A2(new_n12751_), .ZN(new_n13728_));
  NOR2_X1    g11292(.A1(new_n13088_), .A2(new_n13728_), .ZN(new_n13729_));
  AOI21_X1   g11293(.A1(new_n13082_), .A2(new_n13728_), .B(new_n13729_), .ZN(new_n13730_));
  OAI21_X1   g11294(.A1(new_n13730_), .A2(pi0642), .B(new_n13727_), .ZN(new_n13731_));
  AOI21_X1   g11295(.A1(new_n13731_), .A2(new_n13570_), .B(pi0614), .ZN(new_n13732_));
  OAI21_X1   g11296(.A1(new_n13732_), .A2(new_n13701_), .B(new_n13111_), .ZN(new_n13733_));
  AOI21_X1   g11297(.A1(new_n13733_), .A2(new_n13700_), .B(new_n13585_), .ZN(new_n13734_));
  INV_X1     g11298(.I(new_n13489_), .ZN(new_n13735_));
  NOR2_X1    g11299(.A1(new_n13492_), .A2(pi0603), .ZN(new_n13736_));
  OAI22_X1   g11300(.A1(new_n13304_), .A2(new_n12751_), .B1(new_n13290_), .B2(new_n13626_), .ZN(new_n13737_));
  OAI21_X1   g11301(.A1(new_n13737_), .A2(new_n13736_), .B(new_n5404_), .ZN(new_n13738_));
  NAND2_X1   g11302(.A1(new_n13738_), .A2(new_n13735_), .ZN(new_n13739_));
  NOR3_X1    g11303(.A1(new_n13734_), .A2(new_n5445_), .A3(new_n13739_), .ZN(new_n13740_));
  NOR2_X1    g11304(.A1(new_n13088_), .A2(new_n13571_), .ZN(new_n13741_));
  INV_X1     g11305(.I(new_n13741_), .ZN(new_n13742_));
  AOI21_X1   g11306(.A1(new_n13742_), .A2(new_n2641_), .B(pi0223), .ZN(new_n13743_));
  OAI21_X1   g11307(.A1(new_n13740_), .A2(new_n13726_), .B(new_n13743_), .ZN(new_n13744_));
  AOI21_X1   g11308(.A1(new_n13744_), .A2(new_n13720_), .B(pi0299), .ZN(new_n13745_));
  NOR3_X1    g11309(.A1(new_n13709_), .A2(new_n6764_), .A3(new_n13696_), .ZN(new_n13746_));
  NOR4_X1    g11310(.A1(new_n13717_), .A2(new_n13711_), .A3(new_n5422_), .A4(new_n13718_), .ZN(new_n13747_));
  OAI21_X1   g11311(.A1(new_n13746_), .A2(new_n13747_), .B(pi0215), .ZN(new_n13748_));
  AOI21_X1   g11312(.A1(new_n13742_), .A2(new_n3303_), .B(pi0215), .ZN(new_n13749_));
  NAND2_X1   g11313(.A1(new_n13724_), .A2(new_n6764_), .ZN(new_n13750_));
  NAND3_X1   g11314(.A1(new_n13738_), .A2(new_n13735_), .A3(new_n5422_), .ZN(new_n13751_));
  OAI21_X1   g11315(.A1(new_n13734_), .A2(new_n13751_), .B(new_n13750_), .ZN(new_n13752_));
  OAI21_X1   g11316(.A1(new_n13752_), .A2(new_n3303_), .B(new_n13749_), .ZN(new_n13753_));
  AOI21_X1   g11317(.A1(new_n13753_), .A2(new_n13748_), .B(new_n2628_), .ZN(new_n13754_));
  NOR3_X1    g11318(.A1(new_n13745_), .A2(new_n13754_), .A3(pi0140), .ZN(new_n13755_));
  INV_X1     g11319(.I(new_n13238_), .ZN(new_n13756_));
  NOR2_X1    g11320(.A1(new_n13756_), .A2(new_n13598_), .ZN(new_n13757_));
  INV_X1     g11321(.I(new_n5407_), .ZN(new_n13758_));
  NAND2_X1   g11322(.A1(new_n13265_), .A2(new_n13419_), .ZN(new_n13759_));
  OAI21_X1   g11323(.A1(new_n13759_), .A2(new_n13758_), .B(new_n13111_), .ZN(new_n13760_));
  AOI21_X1   g11324(.A1(new_n13629_), .A2(new_n13758_), .B(new_n13760_), .ZN(new_n13761_));
  AOI21_X1   g11325(.A1(new_n13759_), .A2(pi0616), .B(new_n13585_), .ZN(new_n13762_));
  INV_X1     g11326(.I(new_n13762_), .ZN(new_n13763_));
  OAI22_X1   g11327(.A1(new_n13738_), .A2(new_n13109_), .B1(new_n13761_), .B2(new_n13763_), .ZN(new_n13764_));
  NAND2_X1   g11328(.A1(new_n13764_), .A2(new_n5446_), .ZN(new_n13765_));
  NAND2_X1   g11329(.A1(new_n13429_), .A2(new_n13609_), .ZN(new_n13766_));
  NAND2_X1   g11330(.A1(new_n13766_), .A2(new_n13585_), .ZN(new_n13767_));
  OAI21_X1   g11331(.A1(new_n13433_), .A2(new_n13316_), .B(new_n12751_), .ZN(new_n13768_));
  AOI21_X1   g11332(.A1(new_n13768_), .A2(new_n13609_), .B(new_n13264_), .ZN(new_n13769_));
  AOI21_X1   g11333(.A1(new_n13317_), .A2(new_n13605_), .B(new_n5408_), .ZN(new_n13770_));
  OAI21_X1   g11334(.A1(new_n13770_), .A2(new_n13769_), .B(new_n13119_), .ZN(new_n13771_));
  NAND3_X1   g11335(.A1(new_n13771_), .A2(new_n5445_), .A3(new_n13767_), .ZN(new_n13772_));
  NAND3_X1   g11336(.A1(new_n13765_), .A2(new_n13772_), .A3(new_n2642_), .ZN(new_n13773_));
  AOI21_X1   g11337(.A1(new_n13268_), .A2(new_n13266_), .B(new_n12823_), .ZN(new_n13774_));
  OAI21_X1   g11338(.A1(new_n13774_), .A2(pi0616), .B(new_n13762_), .ZN(new_n13775_));
  OR3_X2     g11339(.A1(new_n13263_), .A2(new_n13271_), .A3(new_n13628_), .Z(new_n13776_));
  AOI21_X1   g11340(.A1(new_n13775_), .A2(new_n13776_), .B(new_n5445_), .ZN(new_n13777_));
  NAND2_X1   g11341(.A1(new_n13274_), .A2(new_n13571_), .ZN(new_n13778_));
  NOR2_X1    g11342(.A1(new_n13277_), .A2(new_n13628_), .ZN(new_n13779_));
  OAI21_X1   g11343(.A1(new_n13262_), .A2(new_n12751_), .B(new_n13627_), .ZN(new_n13780_));
  NAND3_X1   g11344(.A1(new_n13780_), .A2(new_n5405_), .A3(new_n5406_), .ZN(new_n13781_));
  OAI21_X1   g11345(.A1(new_n13781_), .A2(pi0616), .B(new_n13779_), .ZN(new_n13782_));
  AOI22_X1   g11346(.A1(new_n13782_), .A2(new_n13119_), .B1(new_n13585_), .B2(new_n13778_), .ZN(new_n13783_));
  AOI21_X1   g11347(.A1(new_n13783_), .A2(new_n5445_), .B(new_n13777_), .ZN(new_n13784_));
  OAI21_X1   g11348(.A1(new_n13784_), .A2(new_n2668_), .B(new_n2628_), .ZN(new_n13785_));
  AOI21_X1   g11349(.A1(new_n13773_), .A2(new_n13757_), .B(new_n13785_), .ZN(new_n13786_));
  NOR2_X1    g11350(.A1(new_n13783_), .A2(new_n5422_), .ZN(new_n13787_));
  AND3_X2    g11351(.A1(new_n13775_), .A2(new_n5422_), .A3(new_n13776_), .Z(new_n13788_));
  OAI21_X1   g11352(.A1(new_n13787_), .A2(new_n13788_), .B(pi0215), .ZN(new_n13789_));
  AOI21_X1   g11353(.A1(new_n13639_), .A2(new_n13571_), .B(pi0215), .ZN(new_n13790_));
  AOI21_X1   g11354(.A1(new_n13771_), .A2(new_n13767_), .B(new_n5422_), .ZN(new_n13791_));
  OAI21_X1   g11355(.A1(new_n13764_), .A2(new_n6764_), .B(new_n3304_), .ZN(new_n13792_));
  OAI21_X1   g11356(.A1(new_n13792_), .A2(new_n13791_), .B(new_n13790_), .ZN(new_n13793_));
  AOI21_X1   g11357(.A1(new_n13793_), .A2(new_n13789_), .B(new_n2628_), .ZN(new_n13794_));
  NOR3_X1    g11358(.A1(new_n13794_), .A2(new_n13786_), .A3(new_n7934_), .ZN(new_n13795_));
  NOR3_X1    g11359(.A1(new_n13755_), .A2(new_n12750_), .A3(new_n13795_), .ZN(new_n13796_));
  OAI21_X1   g11360(.A1(new_n13694_), .A2(new_n13796_), .B(pi0039), .ZN(new_n13797_));
  NOR2_X1    g11361(.A1(new_n13202_), .A2(new_n13207_), .ZN(new_n13798_));
  AOI21_X1   g11362(.A1(new_n13416_), .A2(new_n13798_), .B(new_n7934_), .ZN(new_n13799_));
  NOR2_X1    g11363(.A1(new_n13256_), .A2(new_n13405_), .ZN(new_n13800_));
  NOR2_X1    g11364(.A1(new_n13800_), .A2(pi0140), .ZN(new_n13801_));
  OAI21_X1   g11365(.A1(new_n13801_), .A2(new_n13799_), .B(new_n12750_), .ZN(new_n13802_));
  NAND2_X1   g11366(.A1(new_n13248_), .A2(pi0621), .ZN(new_n13803_));
  OAI22_X1   g11367(.A1(new_n13411_), .A2(pi0603), .B1(new_n13803_), .B2(new_n13626_), .ZN(new_n13804_));
  NAND3_X1   g11368(.A1(new_n13804_), .A2(pi0299), .A3(pi0680), .ZN(new_n13805_));
  OAI22_X1   g11369(.A1(new_n13414_), .A2(pi0603), .B1(new_n13254_), .B2(new_n13626_), .ZN(new_n13806_));
  NAND3_X1   g11370(.A1(new_n13806_), .A2(new_n2628_), .A3(pi0680), .ZN(new_n13807_));
  AOI21_X1   g11371(.A1(new_n13805_), .A2(new_n13807_), .B(new_n7934_), .ZN(new_n13808_));
  NOR2_X1    g11372(.A1(new_n13798_), .A2(new_n12821_), .ZN(new_n13809_));
  NOR3_X1    g11373(.A1(new_n13809_), .A2(new_n13406_), .A3(pi0140), .ZN(new_n13810_));
  OAI21_X1   g11374(.A1(new_n13810_), .A2(new_n13808_), .B(pi0761), .ZN(new_n13811_));
  NAND3_X1   g11375(.A1(new_n13802_), .A2(new_n13811_), .A3(new_n2627_), .ZN(new_n13812_));
  NAND3_X1   g11376(.A1(new_n13797_), .A2(new_n3265_), .A3(new_n13812_), .ZN(new_n13813_));
  AOI21_X1   g11377(.A1(new_n13813_), .A2(new_n13577_), .B(pi0738), .ZN(new_n13814_));
  OAI21_X1   g11378(.A1(new_n13348_), .A2(new_n12820_), .B(new_n2609_), .ZN(new_n13815_));
  OAI21_X1   g11379(.A1(new_n13814_), .A2(new_n13815_), .B(new_n13394_), .ZN(new_n13816_));
  NAND2_X1   g11380(.A1(new_n13816_), .A2(pi0625), .ZN(new_n13817_));
  OR2_X2     g11381(.A1(new_n13349_), .A2(pi0625), .Z(new_n13818_));
  AOI21_X1   g11382(.A1(new_n13817_), .A2(new_n13818_), .B(new_n12841_), .ZN(new_n13819_));
  NOR3_X1    g11383(.A1(new_n13819_), .A2(new_n13560_), .A3(new_n13524_), .ZN(new_n13820_));
  NOR2_X1    g11384(.A1(new_n13349_), .A2(new_n13521_), .ZN(new_n13821_));
  AOI21_X1   g11385(.A1(new_n13816_), .A2(new_n13521_), .B(new_n13821_), .ZN(new_n13822_));
  OAI21_X1   g11386(.A1(new_n13822_), .A2(pi1153), .B(new_n13527_), .ZN(new_n13823_));
  OAI21_X1   g11387(.A1(new_n13823_), .A2(pi0608), .B(pi0778), .ZN(new_n13824_));
  NAND2_X1   g11388(.A1(new_n13816_), .A2(new_n12758_), .ZN(new_n13825_));
  OAI21_X1   g11389(.A1(new_n13824_), .A2(new_n13820_), .B(new_n13825_), .ZN(new_n13826_));
  NAND2_X1   g11390(.A1(new_n13826_), .A2(new_n12764_), .ZN(new_n13827_));
  INV_X1     g11391(.I(new_n13827_), .ZN(new_n13828_));
  INV_X1     g11392(.I(pi0660), .ZN(new_n13829_));
  NOR2_X1    g11393(.A1(new_n13356_), .A2(new_n13829_), .ZN(new_n13830_));
  AOI21_X1   g11394(.A1(new_n13529_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n13831_));
  OAI21_X1   g11395(.A1(new_n13826_), .A2(new_n12766_), .B(new_n13831_), .ZN(new_n13832_));
  NAND2_X1   g11396(.A1(new_n13832_), .A2(new_n13830_), .ZN(new_n13833_));
  NOR2_X1    g11397(.A1(new_n13358_), .A2(new_n12770_), .ZN(new_n13834_));
  NOR2_X1    g11398(.A1(new_n13834_), .A2(pi0660), .ZN(new_n13835_));
  AOI21_X1   g11399(.A1(new_n13529_), .A2(pi0609), .B(pi1155), .ZN(new_n13836_));
  OAI21_X1   g11400(.A1(new_n13826_), .A2(pi0609), .B(new_n13836_), .ZN(new_n13837_));
  AOI21_X1   g11401(.A1(new_n13837_), .A2(new_n13835_), .B(new_n12764_), .ZN(new_n13838_));
  AOI21_X1   g11402(.A1(new_n13838_), .A2(new_n13833_), .B(new_n13828_), .ZN(new_n13839_));
  OR2_X2     g11403(.A1(new_n13839_), .A2(pi0781), .Z(new_n13840_));
  NAND2_X1   g11404(.A1(new_n13364_), .A2(pi0627), .ZN(new_n13841_));
  NOR2_X1    g11405(.A1(new_n13530_), .A2(pi0618), .ZN(new_n13842_));
  NOR2_X1    g11406(.A1(new_n13842_), .A2(new_n12785_), .ZN(new_n13843_));
  NAND2_X1   g11407(.A1(new_n13839_), .A2(pi0618), .ZN(new_n13844_));
  AOI21_X1   g11408(.A1(new_n13844_), .A2(new_n13843_), .B(new_n13841_), .ZN(new_n13845_));
  NAND2_X1   g11409(.A1(new_n13367_), .A2(new_n12880_), .ZN(new_n13846_));
  OAI21_X1   g11410(.A1(new_n13530_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n13847_));
  AOI21_X1   g11411(.A1(new_n13839_), .A2(new_n12781_), .B(new_n13847_), .ZN(new_n13848_));
  OAI21_X1   g11412(.A1(new_n13848_), .A2(new_n13846_), .B(pi0781), .ZN(new_n13849_));
  OAI21_X1   g11413(.A1(new_n13849_), .A2(new_n13845_), .B(new_n13840_), .ZN(new_n13850_));
  AND2_X2    g11414(.A1(new_n13850_), .A2(new_n12796_), .Z(new_n13851_));
  AOI21_X1   g11415(.A1(new_n13371_), .A2(new_n12791_), .B(new_n12895_), .ZN(new_n13852_));
  AOI21_X1   g11416(.A1(new_n13532_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n13853_));
  OAI21_X1   g11417(.A1(new_n13850_), .A2(new_n12793_), .B(new_n13853_), .ZN(new_n13854_));
  NAND2_X1   g11418(.A1(new_n13854_), .A2(new_n13852_), .ZN(new_n13855_));
  AOI21_X1   g11419(.A1(new_n13374_), .A2(pi1159), .B(pi0648), .ZN(new_n13856_));
  AOI21_X1   g11420(.A1(new_n13532_), .A2(pi0619), .B(pi1159), .ZN(new_n13857_));
  OAI21_X1   g11421(.A1(new_n13850_), .A2(pi0619), .B(new_n13857_), .ZN(new_n13858_));
  AOI21_X1   g11422(.A1(new_n13858_), .A2(new_n13856_), .B(new_n12796_), .ZN(new_n13859_));
  AOI21_X1   g11423(.A1(new_n13859_), .A2(new_n13855_), .B(new_n13851_), .ZN(new_n13860_));
  OAI21_X1   g11424(.A1(new_n13860_), .A2(new_n12747_), .B(new_n13559_), .ZN(new_n13861_));
  NAND2_X1   g11425(.A1(new_n13861_), .A2(new_n13558_), .ZN(new_n13862_));
  OAI21_X1   g11426(.A1(new_n13381_), .A2(pi1158), .B(new_n12904_), .ZN(new_n13863_));
  AOI21_X1   g11427(.A1(new_n13534_), .A2(pi0626), .B(pi0641), .ZN(new_n13864_));
  OAI21_X1   g11428(.A1(new_n13860_), .A2(pi0626), .B(new_n13864_), .ZN(new_n13865_));
  AOI21_X1   g11429(.A1(new_n13865_), .A2(new_n13863_), .B(new_n12808_), .ZN(new_n13866_));
  AND2_X2    g11430(.A1(new_n13860_), .A2(new_n12808_), .Z(new_n13867_));
  AOI21_X1   g11431(.A1(new_n13866_), .A2(new_n13862_), .B(new_n13867_), .ZN(new_n13868_));
  OAI21_X1   g11432(.A1(new_n13868_), .A2(new_n12920_), .B(new_n13556_), .ZN(new_n13869_));
  NAND2_X1   g11433(.A1(new_n13869_), .A2(new_n13555_), .ZN(new_n13870_));
  NOR2_X1    g11434(.A1(new_n13542_), .A2(pi0629), .ZN(new_n13871_));
  AOI21_X1   g11435(.A1(new_n13383_), .A2(pi0628), .B(pi1156), .ZN(new_n13872_));
  OAI21_X1   g11436(.A1(new_n13868_), .A2(pi0628), .B(new_n13872_), .ZN(new_n13873_));
  AOI21_X1   g11437(.A1(new_n13873_), .A2(new_n13871_), .B(new_n12937_), .ZN(new_n13874_));
  AND2_X2    g11438(.A1(new_n13868_), .A2(new_n12937_), .Z(new_n13875_));
  AOI21_X1   g11439(.A1(new_n13874_), .A2(new_n13870_), .B(new_n13875_), .ZN(new_n13876_));
  OR2_X2     g11440(.A1(new_n13876_), .A2(pi0787), .Z(new_n13877_));
  OR2_X2     g11441(.A1(new_n13548_), .A2(new_n12981_), .Z(new_n13878_));
  NOR2_X1    g11442(.A1(new_n13387_), .A2(pi0647), .ZN(new_n13879_));
  NOR2_X1    g11443(.A1(new_n13879_), .A2(new_n12965_), .ZN(new_n13880_));
  NAND2_X1   g11444(.A1(new_n13876_), .A2(pi0647), .ZN(new_n13881_));
  AOI21_X1   g11445(.A1(new_n13881_), .A2(new_n13880_), .B(new_n13878_), .ZN(new_n13882_));
  NAND2_X1   g11446(.A1(new_n13551_), .A2(new_n12981_), .ZN(new_n13883_));
  OAI21_X1   g11447(.A1(new_n13387_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n13884_));
  AOI21_X1   g11448(.A1(new_n13876_), .A2(new_n12741_), .B(new_n13884_), .ZN(new_n13885_));
  OAI21_X1   g11449(.A1(new_n13885_), .A2(new_n13883_), .B(pi0787), .ZN(new_n13886_));
  OAI21_X1   g11450(.A1(new_n13886_), .A2(new_n13882_), .B(new_n13877_), .ZN(new_n13887_));
  OAI21_X1   g11451(.A1(new_n13887_), .A2(pi0644), .B(new_n13554_), .ZN(new_n13888_));
  NAND2_X1   g11452(.A1(new_n13888_), .A2(new_n13391_), .ZN(new_n13889_));
  AOI21_X1   g11453(.A1(new_n13194_), .A2(new_n12975_), .B(pi0715), .ZN(new_n13890_));
  NAND2_X1   g11454(.A1(new_n13389_), .A2(pi0644), .ZN(new_n13891_));
  AOI21_X1   g11455(.A1(new_n13891_), .A2(new_n13890_), .B(new_n12739_), .ZN(new_n13892_));
  NOR2_X1    g11456(.A1(new_n13553_), .A2(pi0644), .ZN(new_n13893_));
  AOI21_X1   g11457(.A1(new_n13887_), .A2(pi0644), .B(new_n13893_), .ZN(new_n13894_));
  OAI21_X1   g11458(.A1(new_n13894_), .A2(new_n12740_), .B(new_n13892_), .ZN(new_n13895_));
  NAND3_X1   g11459(.A1(new_n13895_), .A2(new_n13889_), .A3(pi0790), .ZN(new_n13896_));
  AOI21_X1   g11460(.A1(new_n13887_), .A2(new_n13000_), .B(po1038), .ZN(new_n13897_));
  NAND2_X1   g11461(.A1(new_n13896_), .A2(new_n13897_), .ZN(new_n13898_));
  AOI21_X1   g11462(.A1(new_n13898_), .A2(new_n13003_), .B(new_n13002_), .ZN(po0297));
  NOR2_X1    g11463(.A1(new_n3042_), .A2(pi0141), .ZN(new_n13900_));
  INV_X1     g11464(.I(new_n13900_), .ZN(new_n13901_));
  AOI21_X1   g11465(.A1(new_n12756_), .A2(pi0749), .B(new_n13900_), .ZN(new_n13902_));
  NOR3_X1    g11466(.A1(new_n13902_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n13903_));
  NOR2_X1    g11467(.A1(new_n13902_), .A2(new_n12762_), .ZN(new_n13904_));
  AOI21_X1   g11468(.A1(new_n13904_), .A2(new_n12768_), .B(pi1155), .ZN(new_n13905_));
  INV_X1     g11469(.I(new_n13902_), .ZN(new_n13906_));
  AOI21_X1   g11470(.A1(new_n13906_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n13907_));
  NOR3_X1    g11471(.A1(new_n13905_), .A2(new_n13907_), .A3(new_n12764_), .ZN(new_n13908_));
  NOR2_X1    g11472(.A1(new_n13908_), .A2(new_n13903_), .ZN(new_n13909_));
  NOR2_X1    g11473(.A1(new_n13909_), .A2(pi0781), .ZN(new_n13910_));
  INV_X1     g11474(.I(new_n13909_), .ZN(new_n13911_));
  AOI21_X1   g11475(.A1(new_n13911_), .A2(new_n12783_), .B(pi1154), .ZN(new_n13912_));
  AOI21_X1   g11476(.A1(new_n13911_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n13913_));
  NOR3_X1    g11477(.A1(new_n13912_), .A2(new_n13913_), .A3(new_n12779_), .ZN(new_n13914_));
  NOR2_X1    g11478(.A1(new_n13914_), .A2(new_n13910_), .ZN(new_n13915_));
  NOR3_X1    g11479(.A1(new_n13914_), .A2(pi0619), .A3(new_n13910_), .ZN(new_n13916_));
  NOR2_X1    g11480(.A1(new_n13900_), .A2(new_n12793_), .ZN(new_n13917_));
  OAI21_X1   g11481(.A1(new_n13916_), .A2(new_n13917_), .B(new_n12791_), .ZN(new_n13918_));
  NAND2_X1   g11482(.A1(new_n13915_), .A2(pi0619), .ZN(new_n13919_));
  NAND2_X1   g11483(.A1(new_n13901_), .A2(new_n12793_), .ZN(new_n13920_));
  AOI21_X1   g11484(.A1(new_n13919_), .A2(new_n13920_), .B(new_n12791_), .ZN(new_n13921_));
  NOR2_X1    g11485(.A1(new_n13921_), .A2(new_n12796_), .ZN(new_n13922_));
  NAND2_X1   g11486(.A1(new_n13922_), .A2(new_n13918_), .ZN(new_n13923_));
  OAI21_X1   g11487(.A1(pi0789), .A2(new_n13915_), .B(new_n13923_), .ZN(new_n13924_));
  NAND2_X1   g11488(.A1(new_n13924_), .A2(new_n12804_), .ZN(new_n13925_));
  OAI21_X1   g11489(.A1(new_n12749_), .A2(new_n13901_), .B(new_n13925_), .ZN(new_n13926_));
  NAND2_X1   g11490(.A1(new_n13926_), .A2(pi0788), .ZN(new_n13927_));
  NAND2_X1   g11491(.A1(new_n13924_), .A2(new_n12808_), .ZN(new_n13928_));
  NAND2_X1   g11492(.A1(new_n13927_), .A2(new_n13928_), .ZN(new_n13929_));
  NOR2_X1    g11493(.A1(new_n13929_), .A2(pi0628), .ZN(new_n13930_));
  AOI21_X1   g11494(.A1(new_n12826_), .A2(pi0706), .B(new_n13900_), .ZN(new_n13931_));
  NOR2_X1    g11495(.A1(new_n13931_), .A2(new_n12754_), .ZN(new_n13932_));
  NOR2_X1    g11496(.A1(new_n13932_), .A2(new_n13906_), .ZN(new_n13933_));
  NAND2_X1   g11497(.A1(new_n13933_), .A2(new_n12758_), .ZN(new_n13934_));
  INV_X1     g11498(.I(pi0706), .ZN(new_n13935_));
  NOR2_X1    g11499(.A1(new_n12834_), .A2(new_n13935_), .ZN(new_n13936_));
  INV_X1     g11500(.I(new_n13936_), .ZN(new_n13937_));
  NOR2_X1    g11501(.A1(new_n13900_), .A2(pi1153), .ZN(new_n13938_));
  NAND2_X1   g11502(.A1(new_n13937_), .A2(new_n13938_), .ZN(new_n13939_));
  NAND2_X1   g11503(.A1(new_n13932_), .A2(pi0625), .ZN(new_n13940_));
  NAND3_X1   g11504(.A1(new_n13940_), .A2(pi1153), .A3(new_n13902_), .ZN(new_n13941_));
  AND3_X2    g11505(.A1(new_n13939_), .A2(pi0608), .A3(new_n13941_), .Z(new_n13942_));
  NOR2_X1    g11506(.A1(new_n13936_), .A2(new_n13931_), .ZN(new_n13943_));
  NOR2_X1    g11507(.A1(new_n13943_), .A2(new_n12841_), .ZN(new_n13944_));
  NOR2_X1    g11508(.A1(new_n13944_), .A2(pi0608), .ZN(new_n13945_));
  INV_X1     g11509(.I(new_n13940_), .ZN(new_n13946_));
  OAI21_X1   g11510(.A1(new_n13946_), .A2(new_n13933_), .B(new_n13938_), .ZN(new_n13947_));
  NAND2_X1   g11511(.A1(new_n13945_), .A2(new_n13947_), .ZN(new_n13948_));
  NAND2_X1   g11512(.A1(new_n13948_), .A2(pi0778), .ZN(new_n13949_));
  OAI21_X1   g11513(.A1(new_n13949_), .A2(new_n13942_), .B(new_n13934_), .ZN(new_n13950_));
  INV_X1     g11514(.I(new_n13950_), .ZN(new_n13951_));
  NOR2_X1    g11515(.A1(new_n13931_), .A2(pi0778), .ZN(new_n13952_));
  INV_X1     g11516(.I(new_n13939_), .ZN(new_n13953_));
  NOR3_X1    g11517(.A1(new_n13953_), .A2(new_n12758_), .A3(new_n13944_), .ZN(new_n13954_));
  NOR2_X1    g11518(.A1(new_n13954_), .A2(new_n13952_), .ZN(new_n13955_));
  INV_X1     g11519(.I(new_n13955_), .ZN(new_n13956_));
  NOR2_X1    g11520(.A1(new_n13956_), .A2(pi0609), .ZN(new_n13957_));
  AOI21_X1   g11521(.A1(new_n13950_), .A2(pi0609), .B(new_n13957_), .ZN(new_n13958_));
  NOR2_X1    g11522(.A1(new_n13958_), .A2(new_n12770_), .ZN(new_n13959_));
  NOR2_X1    g11523(.A1(new_n13959_), .A2(new_n13905_), .ZN(new_n13960_));
  NOR2_X1    g11524(.A1(new_n13951_), .A2(pi0609), .ZN(new_n13961_));
  NOR2_X1    g11525(.A1(new_n13956_), .A2(new_n12766_), .ZN(new_n13962_));
  OAI21_X1   g11526(.A1(new_n13961_), .A2(new_n13962_), .B(new_n12770_), .ZN(new_n13963_));
  NOR2_X1    g11527(.A1(new_n13907_), .A2(pi0660), .ZN(new_n13964_));
  AOI22_X1   g11528(.A1(new_n13960_), .A2(pi0660), .B1(new_n13963_), .B2(new_n13964_), .ZN(new_n13965_));
  NAND2_X1   g11529(.A1(new_n13965_), .A2(pi0785), .ZN(new_n13966_));
  OAI21_X1   g11530(.A1(pi0785), .A2(new_n13951_), .B(new_n13966_), .ZN(new_n13967_));
  INV_X1     g11531(.I(new_n13913_), .ZN(new_n13968_));
  NOR2_X1    g11532(.A1(new_n13955_), .A2(new_n12871_), .ZN(new_n13969_));
  NOR2_X1    g11533(.A1(new_n13969_), .A2(new_n12781_), .ZN(new_n13970_));
  AOI21_X1   g11534(.A1(new_n13967_), .A2(new_n12781_), .B(new_n13970_), .ZN(new_n13971_));
  OAI21_X1   g11535(.A1(new_n13971_), .A2(pi1154), .B(new_n13968_), .ZN(new_n13972_));
  INV_X1     g11536(.I(new_n13969_), .ZN(new_n13973_));
  NAND2_X1   g11537(.A1(new_n13973_), .A2(new_n12781_), .ZN(new_n13974_));
  NAND2_X1   g11538(.A1(new_n13967_), .A2(pi0618), .ZN(new_n13975_));
  AOI21_X1   g11539(.A1(new_n13975_), .A2(new_n13974_), .B(new_n12785_), .ZN(new_n13976_));
  OR2_X2     g11540(.A1(new_n13912_), .A2(new_n12880_), .Z(new_n13977_));
  OAI22_X1   g11541(.A1(new_n13972_), .A2(pi0627), .B1(new_n13976_), .B2(new_n13977_), .ZN(new_n13978_));
  NOR2_X1    g11542(.A1(new_n13978_), .A2(new_n12779_), .ZN(new_n13979_));
  AOI21_X1   g11543(.A1(new_n12779_), .A2(new_n13967_), .B(new_n13979_), .ZN(new_n13980_));
  OAI21_X1   g11544(.A1(new_n13980_), .A2(pi0789), .B(new_n12819_), .ZN(new_n13981_));
  NOR2_X1    g11545(.A1(new_n13973_), .A2(new_n12889_), .ZN(new_n13982_));
  NOR2_X1    g11546(.A1(new_n13982_), .A2(pi0619), .ZN(new_n13983_));
  NOR2_X1    g11547(.A1(new_n13980_), .A2(new_n12793_), .ZN(new_n13984_));
  OAI21_X1   g11548(.A1(new_n13984_), .A2(new_n13983_), .B(pi1159), .ZN(new_n13985_));
  NAND3_X1   g11549(.A1(new_n13985_), .A2(pi0648), .A3(new_n13918_), .ZN(new_n13986_));
  INV_X1     g11550(.I(new_n13982_), .ZN(new_n13987_));
  NAND2_X1   g11551(.A1(new_n13987_), .A2(pi0619), .ZN(new_n13988_));
  OAI21_X1   g11552(.A1(new_n13980_), .A2(pi0619), .B(new_n13988_), .ZN(new_n13989_));
  AOI21_X1   g11553(.A1(new_n13989_), .A2(new_n12791_), .B(new_n13921_), .ZN(new_n13990_));
  AOI21_X1   g11554(.A1(new_n13990_), .A2(new_n12895_), .B(new_n12796_), .ZN(new_n13991_));
  AOI21_X1   g11555(.A1(new_n13991_), .A2(new_n13986_), .B(new_n13981_), .ZN(new_n13992_));
  AOI22_X1   g11556(.A1(new_n13926_), .A2(new_n12914_), .B1(new_n12913_), .B2(new_n13982_), .ZN(new_n13993_));
  NOR2_X1    g11557(.A1(new_n13993_), .A2(new_n12808_), .ZN(new_n13994_));
  NOR2_X1    g11558(.A1(new_n13992_), .A2(new_n13994_), .ZN(new_n13995_));
  AOI21_X1   g11559(.A1(new_n13995_), .A2(pi0628), .B(new_n13930_), .ZN(new_n13996_));
  NOR2_X1    g11560(.A1(new_n13987_), .A2(new_n12924_), .ZN(new_n13997_));
  NAND2_X1   g11561(.A1(new_n13997_), .A2(new_n12922_), .ZN(new_n13998_));
  AOI21_X1   g11562(.A1(new_n13998_), .A2(new_n12742_), .B(new_n12919_), .ZN(new_n13999_));
  OAI21_X1   g11563(.A1(new_n13996_), .A2(new_n12742_), .B(new_n13999_), .ZN(new_n14000_));
  NOR2_X1    g11564(.A1(new_n13929_), .A2(new_n12920_), .ZN(new_n14001_));
  AOI21_X1   g11565(.A1(new_n13995_), .A2(new_n12920_), .B(new_n14001_), .ZN(new_n14002_));
  NAND2_X1   g11566(.A1(new_n13997_), .A2(new_n12932_), .ZN(new_n14003_));
  AOI21_X1   g11567(.A1(new_n14003_), .A2(pi1156), .B(pi0629), .ZN(new_n14004_));
  OAI21_X1   g11568(.A1(new_n14002_), .A2(pi1156), .B(new_n14004_), .ZN(new_n14005_));
  NAND3_X1   g11569(.A1(new_n14000_), .A2(new_n14005_), .A3(pi0792), .ZN(new_n14006_));
  NAND2_X1   g11570(.A1(new_n13995_), .A2(new_n12937_), .ZN(new_n14007_));
  AOI21_X1   g11571(.A1(new_n14006_), .A2(new_n14007_), .B(new_n12741_), .ZN(new_n14008_));
  NOR2_X1    g11572(.A1(new_n13929_), .A2(new_n12943_), .ZN(new_n14009_));
  AOI21_X1   g11573(.A1(new_n12943_), .A2(new_n13901_), .B(new_n14009_), .ZN(new_n14010_));
  NOR2_X1    g11574(.A1(new_n14010_), .A2(pi0647), .ZN(new_n14011_));
  OAI21_X1   g11575(.A1(new_n14008_), .A2(new_n14011_), .B(pi1157), .ZN(new_n14012_));
  NAND2_X1   g11576(.A1(new_n13997_), .A2(new_n12954_), .ZN(new_n14013_));
  NAND2_X1   g11577(.A1(new_n14013_), .A2(new_n12741_), .ZN(new_n14014_));
  NOR2_X1    g11578(.A1(new_n13900_), .A2(new_n12741_), .ZN(new_n14015_));
  INV_X1     g11579(.I(new_n14015_), .ZN(new_n14016_));
  AOI21_X1   g11580(.A1(new_n14014_), .A2(new_n14016_), .B(pi1157), .ZN(new_n14017_));
  INV_X1     g11581(.I(new_n14017_), .ZN(new_n14018_));
  NAND3_X1   g11582(.A1(new_n14012_), .A2(pi0630), .A3(new_n14018_), .ZN(new_n14019_));
  NAND2_X1   g11583(.A1(new_n14006_), .A2(new_n14007_), .ZN(new_n14020_));
  NOR2_X1    g11584(.A1(new_n14010_), .A2(new_n12741_), .ZN(new_n14021_));
  AOI21_X1   g11585(.A1(new_n14020_), .A2(new_n12741_), .B(new_n14021_), .ZN(new_n14022_));
  NAND2_X1   g11586(.A1(new_n14013_), .A2(pi0647), .ZN(new_n14023_));
  NAND2_X1   g11587(.A1(new_n13901_), .A2(new_n12741_), .ZN(new_n14024_));
  AOI21_X1   g11588(.A1(new_n14023_), .A2(new_n14024_), .B(new_n12965_), .ZN(new_n14025_));
  NOR2_X1    g11589(.A1(new_n14025_), .A2(pi0630), .ZN(new_n14026_));
  OAI21_X1   g11590(.A1(new_n14022_), .A2(pi1157), .B(new_n14026_), .ZN(new_n14027_));
  NAND3_X1   g11591(.A1(new_n14019_), .A2(new_n14027_), .A3(pi0787), .ZN(new_n14028_));
  NAND2_X1   g11592(.A1(new_n14020_), .A2(new_n12972_), .ZN(new_n14029_));
  AOI21_X1   g11593(.A1(new_n14028_), .A2(new_n14029_), .B(pi0644), .ZN(new_n14030_));
  OR2_X2     g11594(.A1(new_n14025_), .A2(new_n12972_), .Z(new_n14031_));
  OAI22_X1   g11595(.A1(new_n14031_), .A2(new_n14017_), .B1(pi0787), .B2(new_n14013_), .ZN(new_n14032_));
  NOR2_X1    g11596(.A1(new_n14032_), .A2(new_n12975_), .ZN(new_n14033_));
  OAI21_X1   g11597(.A1(new_n14030_), .A2(new_n14033_), .B(new_n12740_), .ZN(new_n14034_));
  NAND2_X1   g11598(.A1(new_n14010_), .A2(new_n12985_), .ZN(new_n14035_));
  OAI21_X1   g11599(.A1(new_n12985_), .A2(new_n13901_), .B(new_n14035_), .ZN(new_n14036_));
  NOR2_X1    g11600(.A1(new_n14036_), .A2(pi0644), .ZN(new_n14037_));
  NOR2_X1    g11601(.A1(new_n13900_), .A2(new_n12975_), .ZN(new_n14038_));
  OAI21_X1   g11602(.A1(new_n14037_), .A2(new_n14038_), .B(pi0715), .ZN(new_n14039_));
  NAND3_X1   g11603(.A1(new_n14034_), .A2(new_n12739_), .A3(new_n14039_), .ZN(new_n14040_));
  NAND2_X1   g11604(.A1(new_n14028_), .A2(new_n14029_), .ZN(new_n14041_));
  NOR2_X1    g11605(.A1(new_n14032_), .A2(pi0644), .ZN(new_n14042_));
  AOI21_X1   g11606(.A1(new_n14041_), .A2(pi0644), .B(new_n14042_), .ZN(new_n14043_));
  NAND2_X1   g11607(.A1(new_n13901_), .A2(new_n12975_), .ZN(new_n14044_));
  OAI21_X1   g11608(.A1(new_n14036_), .A2(new_n12975_), .B(new_n14044_), .ZN(new_n14045_));
  AOI21_X1   g11609(.A1(new_n14045_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n14046_));
  OAI21_X1   g11610(.A1(new_n14043_), .A2(new_n12740_), .B(new_n14046_), .ZN(new_n14047_));
  NAND3_X1   g11611(.A1(new_n14040_), .A2(new_n14047_), .A3(pi0790), .ZN(new_n14048_));
  NAND2_X1   g11612(.A1(new_n14041_), .A2(new_n13000_), .ZN(new_n14049_));
  AOI21_X1   g11613(.A1(new_n14048_), .A2(new_n14049_), .B(new_n12738_), .ZN(new_n14050_));
  AOI21_X1   g11614(.A1(po1038), .A2(new_n12638_), .B(pi0832), .ZN(new_n14051_));
  NOR2_X1    g11615(.A1(new_n13193_), .A2(pi0141), .ZN(new_n14052_));
  AOI21_X1   g11616(.A1(new_n14052_), .A2(pi0644), .B(new_n12740_), .ZN(new_n14053_));
  NOR2_X1    g11617(.A1(new_n2609_), .A2(new_n12638_), .ZN(new_n14054_));
  INV_X1     g11618(.I(new_n14054_), .ZN(new_n14055_));
  NOR2_X1    g11619(.A1(new_n13344_), .A2(pi0141), .ZN(new_n14056_));
  AOI21_X1   g11620(.A1(pi0749), .A2(new_n13341_), .B(new_n14056_), .ZN(new_n14057_));
  OR2_X2     g11621(.A1(new_n14057_), .A2(new_n3265_), .Z(new_n14058_));
  INV_X1     g11622(.I(pi0749), .ZN(new_n14059_));
  NOR2_X1    g11623(.A1(new_n13208_), .A2(new_n12638_), .ZN(new_n14060_));
  AOI21_X1   g11624(.A1(new_n13334_), .A2(new_n12638_), .B(new_n14060_), .ZN(new_n14061_));
  NAND3_X1   g11625(.A1(new_n13336_), .A2(new_n12638_), .A3(new_n14059_), .ZN(new_n14062_));
  OAI21_X1   g11626(.A1(new_n14061_), .A2(new_n14059_), .B(new_n14062_), .ZN(new_n14063_));
  NOR2_X1    g11627(.A1(new_n13178_), .A2(new_n13188_), .ZN(new_n14064_));
  INV_X1     g11628(.I(new_n14064_), .ZN(new_n14065_));
  NOR2_X1    g11629(.A1(new_n13234_), .A2(new_n13243_), .ZN(new_n14066_));
  INV_X1     g11630(.I(new_n14066_), .ZN(new_n14067_));
  OAI22_X1   g11631(.A1(new_n14065_), .A2(pi0749), .B1(new_n12638_), .B2(new_n14067_), .ZN(new_n14068_));
  NAND2_X1   g11632(.A1(new_n14068_), .A2(pi0039), .ZN(new_n14069_));
  NAND3_X1   g11633(.A1(new_n14063_), .A2(new_n3265_), .A3(new_n14069_), .ZN(new_n14070_));
  NAND3_X1   g11634(.A1(new_n14070_), .A2(new_n2609_), .A3(new_n14058_), .ZN(new_n14071_));
  NAND2_X1   g11635(.A1(new_n14071_), .A2(new_n14055_), .ZN(new_n14072_));
  NAND2_X1   g11636(.A1(new_n14072_), .A2(new_n12761_), .ZN(new_n14073_));
  INV_X1     g11637(.I(new_n14052_), .ZN(new_n14074_));
  NAND2_X1   g11638(.A1(new_n14074_), .A2(new_n12760_), .ZN(new_n14075_));
  NAND3_X1   g11639(.A1(new_n14073_), .A2(new_n12764_), .A3(new_n14075_), .ZN(new_n14076_));
  OAI22_X1   g11640(.A1(new_n14073_), .A2(pi0609), .B1(new_n13353_), .B2(new_n14052_), .ZN(new_n14077_));
  NAND2_X1   g11641(.A1(new_n14077_), .A2(new_n12770_), .ZN(new_n14078_));
  OAI22_X1   g11642(.A1(new_n14073_), .A2(new_n12766_), .B1(new_n12772_), .B2(new_n14052_), .ZN(new_n14079_));
  NAND2_X1   g11643(.A1(new_n14079_), .A2(pi1155), .ZN(new_n14080_));
  NAND3_X1   g11644(.A1(new_n14078_), .A2(new_n14080_), .A3(pi0785), .ZN(new_n14081_));
  NAND2_X1   g11645(.A1(new_n14081_), .A2(new_n14076_), .ZN(new_n14082_));
  NAND2_X1   g11646(.A1(new_n14082_), .A2(new_n12779_), .ZN(new_n14083_));
  NAND2_X1   g11647(.A1(new_n14074_), .A2(pi0618), .ZN(new_n14084_));
  OAI21_X1   g11648(.A1(new_n14082_), .A2(pi0618), .B(new_n14084_), .ZN(new_n14085_));
  NAND2_X1   g11649(.A1(new_n14085_), .A2(new_n12785_), .ZN(new_n14086_));
  NOR2_X1    g11650(.A1(new_n14082_), .A2(new_n12781_), .ZN(new_n14087_));
  NOR2_X1    g11651(.A1(new_n14052_), .A2(pi0618), .ZN(new_n14088_));
  OAI21_X1   g11652(.A1(new_n14087_), .A2(new_n14088_), .B(pi1154), .ZN(new_n14089_));
  NAND3_X1   g11653(.A1(new_n14089_), .A2(new_n14086_), .A3(pi0781), .ZN(new_n14090_));
  NAND2_X1   g11654(.A1(new_n14090_), .A2(new_n14083_), .ZN(new_n14091_));
  NOR2_X1    g11655(.A1(new_n14091_), .A2(pi0619), .ZN(new_n14092_));
  NOR2_X1    g11656(.A1(new_n14052_), .A2(new_n12793_), .ZN(new_n14093_));
  OAI21_X1   g11657(.A1(new_n14092_), .A2(new_n14093_), .B(new_n12791_), .ZN(new_n14094_));
  NAND2_X1   g11658(.A1(new_n14074_), .A2(new_n12793_), .ZN(new_n14095_));
  OAI21_X1   g11659(.A1(new_n14091_), .A2(new_n12793_), .B(new_n14095_), .ZN(new_n14096_));
  AOI21_X1   g11660(.A1(new_n14096_), .A2(pi1159), .B(new_n12796_), .ZN(new_n14097_));
  AOI22_X1   g11661(.A1(new_n14097_), .A2(new_n14094_), .B1(new_n12796_), .B2(new_n14091_), .ZN(new_n14098_));
  NOR2_X1    g11662(.A1(new_n14052_), .A2(pi0626), .ZN(new_n14099_));
  AOI21_X1   g11663(.A1(new_n14098_), .A2(pi0626), .B(new_n14099_), .ZN(new_n14100_));
  NOR2_X1    g11664(.A1(new_n14100_), .A2(new_n12745_), .ZN(new_n14101_));
  NOR2_X1    g11665(.A1(new_n14052_), .A2(new_n12747_), .ZN(new_n14102_));
  AOI21_X1   g11666(.A1(new_n14098_), .A2(new_n12747_), .B(new_n14102_), .ZN(new_n14103_));
  OAI21_X1   g11667(.A1(new_n14103_), .A2(pi1158), .B(pi0788), .ZN(new_n14104_));
  OAI22_X1   g11668(.A1(new_n14104_), .A2(new_n14101_), .B1(pi0788), .B2(new_n14098_), .ZN(new_n14105_));
  NAND2_X1   g11669(.A1(new_n14074_), .A2(new_n12943_), .ZN(new_n14106_));
  OAI21_X1   g11670(.A1(new_n14105_), .A2(new_n12943_), .B(new_n14106_), .ZN(new_n14107_));
  NAND2_X1   g11671(.A1(new_n14052_), .A2(new_n12984_), .ZN(new_n14108_));
  OAI21_X1   g11672(.A1(new_n14107_), .A2(new_n12984_), .B(new_n14108_), .ZN(new_n14109_));
  NAND2_X1   g11673(.A1(new_n14109_), .A2(new_n12975_), .ZN(new_n14110_));
  AOI21_X1   g11674(.A1(new_n14110_), .A2(new_n14053_), .B(pi1160), .ZN(new_n14111_));
  NOR2_X1    g11675(.A1(new_n14074_), .A2(new_n12870_), .ZN(new_n14112_));
  NOR2_X1    g11676(.A1(pi0141), .A2(pi0706), .ZN(new_n14113_));
  AOI21_X1   g11677(.A1(new_n13395_), .A2(new_n14113_), .B(new_n2610_), .ZN(new_n14114_));
  NOR2_X1    g11678(.A1(new_n13405_), .A2(pi0039), .ZN(new_n14115_));
  INV_X1     g11679(.I(new_n14115_), .ZN(new_n14116_));
  NAND3_X1   g11680(.A1(new_n13502_), .A2(new_n13514_), .A3(pi0039), .ZN(new_n14117_));
  NAND2_X1   g11681(.A1(new_n14117_), .A2(new_n14116_), .ZN(new_n14118_));
  NAND2_X1   g11682(.A1(new_n14118_), .A2(new_n12638_), .ZN(new_n14119_));
  NAND2_X1   g11683(.A1(new_n13416_), .A2(new_n2627_), .ZN(new_n14120_));
  NAND3_X1   g11684(.A1(new_n13442_), .A2(new_n13452_), .A3(pi0039), .ZN(new_n14121_));
  NAND2_X1   g11685(.A1(new_n14121_), .A2(new_n14120_), .ZN(new_n14122_));
  NAND2_X1   g11686(.A1(new_n14122_), .A2(pi0141), .ZN(new_n14123_));
  AOI21_X1   g11687(.A1(new_n14119_), .A2(new_n14123_), .B(pi0038), .ZN(new_n14124_));
  INV_X1     g11688(.I(new_n13399_), .ZN(new_n14125_));
  OAI21_X1   g11689(.A1(new_n14125_), .A2(new_n14056_), .B(pi0706), .ZN(new_n14126_));
  OAI21_X1   g11690(.A1(new_n14124_), .A2(new_n14126_), .B(new_n14114_), .ZN(new_n14127_));
  NAND2_X1   g11691(.A1(new_n14127_), .A2(new_n14055_), .ZN(new_n14128_));
  NOR2_X1    g11692(.A1(new_n13521_), .A2(new_n12841_), .ZN(new_n14129_));
  NOR2_X1    g11693(.A1(pi0625), .A2(pi1153), .ZN(new_n14130_));
  NOR3_X1    g11694(.A1(new_n14129_), .A2(new_n12758_), .A3(new_n14130_), .ZN(new_n14131_));
  XNOR2_X1   g11695(.A1(pi0625), .A2(pi1153), .ZN(new_n14132_));
  INV_X1     g11696(.I(new_n14132_), .ZN(new_n14133_));
  NAND2_X1   g11697(.A1(new_n14052_), .A2(new_n14133_), .ZN(new_n14134_));
  OAI22_X1   g11698(.A1(new_n14128_), .A2(new_n14131_), .B1(new_n12758_), .B2(new_n14134_), .ZN(new_n14135_));
  AOI21_X1   g11699(.A1(new_n14135_), .A2(new_n12870_), .B(new_n14112_), .ZN(new_n14136_));
  NOR2_X1    g11700(.A1(new_n14052_), .A2(new_n12888_), .ZN(new_n14137_));
  AOI21_X1   g11701(.A1(new_n14136_), .A2(new_n12888_), .B(new_n14137_), .ZN(new_n14138_));
  NOR2_X1    g11702(.A1(new_n14074_), .A2(new_n12911_), .ZN(new_n14139_));
  AOI21_X1   g11703(.A1(new_n14138_), .A2(new_n12911_), .B(new_n14139_), .ZN(new_n14140_));
  NOR2_X1    g11704(.A1(new_n14052_), .A2(new_n13392_), .ZN(new_n14141_));
  AOI21_X1   g11705(.A1(new_n14140_), .A2(new_n13392_), .B(new_n14141_), .ZN(new_n14142_));
  NOR2_X1    g11706(.A1(new_n14142_), .A2(pi0628), .ZN(new_n14143_));
  NOR2_X1    g11707(.A1(new_n14052_), .A2(new_n12920_), .ZN(new_n14144_));
  OAI21_X1   g11708(.A1(new_n14143_), .A2(new_n14144_), .B(new_n12742_), .ZN(new_n14145_));
  NOR2_X1    g11709(.A1(new_n14142_), .A2(new_n12920_), .ZN(new_n14146_));
  AOI21_X1   g11710(.A1(new_n12920_), .A2(new_n14074_), .B(new_n14146_), .ZN(new_n14147_));
  NOR2_X1    g11711(.A1(new_n14147_), .A2(new_n12742_), .ZN(new_n14148_));
  NOR2_X1    g11712(.A1(new_n14148_), .A2(new_n12937_), .ZN(new_n14149_));
  AOI22_X1   g11713(.A1(new_n14149_), .A2(new_n14145_), .B1(new_n12937_), .B2(new_n14142_), .ZN(new_n14150_));
  NAND2_X1   g11714(.A1(new_n14150_), .A2(new_n12741_), .ZN(new_n14151_));
  NAND2_X1   g11715(.A1(new_n14074_), .A2(pi0647), .ZN(new_n14152_));
  AOI21_X1   g11716(.A1(new_n14151_), .A2(new_n14152_), .B(pi1157), .ZN(new_n14153_));
  NAND2_X1   g11717(.A1(new_n14150_), .A2(pi0647), .ZN(new_n14154_));
  OAI21_X1   g11718(.A1(pi0647), .A2(new_n14052_), .B(new_n14154_), .ZN(new_n14155_));
  NAND2_X1   g11719(.A1(new_n14155_), .A2(pi1157), .ZN(new_n14156_));
  NAND2_X1   g11720(.A1(new_n14156_), .A2(pi0787), .ZN(new_n14157_));
  OAI22_X1   g11721(.A1(new_n14157_), .A2(new_n14153_), .B1(pi0787), .B2(new_n14150_), .ZN(new_n14158_));
  AOI21_X1   g11722(.A1(new_n14158_), .A2(pi0644), .B(pi0715), .ZN(new_n14159_));
  AOI21_X1   g11723(.A1(new_n14105_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n14160_));
  OAI21_X1   g11724(.A1(new_n14100_), .A2(new_n12745_), .B(new_n13557_), .ZN(new_n14161_));
  AOI21_X1   g11725(.A1(new_n14140_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n14162_));
  AOI21_X1   g11726(.A1(new_n13191_), .A2(new_n2609_), .B(new_n13521_), .ZN(new_n14163_));
  AOI21_X1   g11727(.A1(new_n14163_), .A2(new_n12638_), .B(pi1153), .ZN(new_n14164_));
  OAI21_X1   g11728(.A1(new_n14128_), .A2(pi0625), .B(new_n14164_), .ZN(new_n14165_));
  NAND2_X1   g11729(.A1(new_n14165_), .A2(pi0608), .ZN(new_n14166_));
  NOR2_X1    g11730(.A1(new_n14072_), .A2(pi0625), .ZN(new_n14167_));
  NOR2_X1    g11731(.A1(new_n14167_), .A2(new_n12841_), .ZN(new_n14168_));
  AOI21_X1   g11732(.A1(new_n13573_), .A2(new_n2627_), .B(new_n3265_), .ZN(new_n14169_));
  AOI21_X1   g11733(.A1(new_n14057_), .A2(new_n14169_), .B(new_n13935_), .ZN(new_n14170_));
  INV_X1     g11734(.I(new_n14170_), .ZN(new_n14171_));
  NAND2_X1   g11735(.A1(new_n13416_), .A2(new_n13798_), .ZN(new_n14172_));
  NOR2_X1    g11736(.A1(new_n14172_), .A2(new_n12638_), .ZN(new_n14173_));
  NAND4_X1   g11737(.A1(new_n13250_), .A2(new_n13255_), .A3(new_n13402_), .A4(new_n13404_), .ZN(new_n14174_));
  NOR2_X1    g11738(.A1(new_n14174_), .A2(pi0141), .ZN(new_n14175_));
  OAI21_X1   g11739(.A1(new_n14173_), .A2(new_n14175_), .B(pi0749), .ZN(new_n14176_));
  NOR2_X1    g11740(.A1(new_n13809_), .A2(new_n13406_), .ZN(new_n14177_));
  NAND3_X1   g11741(.A1(new_n13805_), .A2(new_n13807_), .A3(pi0141), .ZN(new_n14178_));
  OAI21_X1   g11742(.A1(new_n14177_), .A2(pi0141), .B(new_n14178_), .ZN(new_n14179_));
  AOI21_X1   g11743(.A1(new_n14179_), .A2(new_n14059_), .B(pi0039), .ZN(new_n14180_));
  AOI21_X1   g11744(.A1(new_n14180_), .A2(new_n14176_), .B(pi0038), .ZN(new_n14181_));
  NOR2_X1    g11745(.A1(new_n13745_), .A2(new_n13754_), .ZN(new_n14182_));
  NOR2_X1    g11746(.A1(new_n14182_), .A2(pi0141), .ZN(new_n14183_));
  NOR2_X1    g11747(.A1(new_n13794_), .A2(new_n13786_), .ZN(new_n14184_));
  NOR2_X1    g11748(.A1(new_n14184_), .A2(new_n12638_), .ZN(new_n14185_));
  OAI21_X1   g11749(.A1(new_n14183_), .A2(new_n14185_), .B(new_n14059_), .ZN(new_n14186_));
  NOR2_X1    g11750(.A1(new_n13651_), .A2(new_n13634_), .ZN(new_n14187_));
  NOR2_X1    g11751(.A1(new_n14187_), .A2(new_n12638_), .ZN(new_n14188_));
  INV_X1     g11752(.I(new_n13692_), .ZN(new_n14189_));
  NOR2_X1    g11753(.A1(new_n14189_), .A2(pi0141), .ZN(new_n14190_));
  OAI21_X1   g11754(.A1(new_n14188_), .A2(new_n14190_), .B(pi0749), .ZN(new_n14191_));
  NAND3_X1   g11755(.A1(new_n14191_), .A2(new_n14186_), .A3(pi0039), .ZN(new_n14192_));
  AOI21_X1   g11756(.A1(new_n14192_), .A2(new_n14181_), .B(new_n14171_), .ZN(new_n14193_));
  AOI21_X1   g11757(.A1(new_n14070_), .A2(new_n14058_), .B(pi0706), .ZN(new_n14194_));
  NOR3_X1    g11758(.A1(new_n14194_), .A2(new_n14193_), .A3(new_n2610_), .ZN(new_n14195_));
  INV_X1     g11759(.I(new_n14195_), .ZN(new_n14196_));
  NAND3_X1   g11760(.A1(new_n14196_), .A2(pi0625), .A3(new_n14055_), .ZN(new_n14197_));
  AOI21_X1   g11761(.A1(new_n14197_), .A2(new_n14168_), .B(new_n14166_), .ZN(new_n14198_));
  AOI21_X1   g11762(.A1(new_n13191_), .A2(new_n2609_), .B(pi0625), .ZN(new_n14199_));
  AOI21_X1   g11763(.A1(new_n14199_), .A2(new_n12638_), .B(new_n12841_), .ZN(new_n14200_));
  NAND3_X1   g11764(.A1(new_n14127_), .A2(pi0625), .A3(new_n14055_), .ZN(new_n14201_));
  AOI21_X1   g11765(.A1(new_n14201_), .A2(new_n14200_), .B(pi0608), .ZN(new_n14202_));
  OAI21_X1   g11766(.A1(new_n14072_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n14203_));
  NOR3_X1    g11767(.A1(new_n14195_), .A2(pi0625), .A3(new_n14054_), .ZN(new_n14204_));
  OAI21_X1   g11768(.A1(new_n14204_), .A2(new_n14203_), .B(new_n14202_), .ZN(new_n14205_));
  NAND2_X1   g11769(.A1(new_n14205_), .A2(pi0778), .ZN(new_n14206_));
  AOI21_X1   g11770(.A1(new_n14196_), .A2(new_n14055_), .B(pi0778), .ZN(new_n14207_));
  INV_X1     g11771(.I(new_n14207_), .ZN(new_n14208_));
  OAI21_X1   g11772(.A1(new_n14206_), .A2(new_n14198_), .B(new_n14208_), .ZN(new_n14209_));
  NAND2_X1   g11773(.A1(new_n14209_), .A2(new_n12764_), .ZN(new_n14210_));
  INV_X1     g11774(.I(new_n14210_), .ZN(new_n14211_));
  AOI21_X1   g11775(.A1(new_n14077_), .A2(new_n12770_), .B(new_n13829_), .ZN(new_n14212_));
  AOI21_X1   g11776(.A1(new_n14135_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n14213_));
  OAI21_X1   g11777(.A1(new_n14209_), .A2(new_n12766_), .B(new_n14213_), .ZN(new_n14214_));
  NAND2_X1   g11778(.A1(new_n14214_), .A2(new_n14212_), .ZN(new_n14215_));
  AOI21_X1   g11779(.A1(new_n14079_), .A2(pi1155), .B(pi0660), .ZN(new_n14216_));
  AOI21_X1   g11780(.A1(new_n14135_), .A2(pi0609), .B(pi1155), .ZN(new_n14217_));
  OAI21_X1   g11781(.A1(new_n14209_), .A2(pi0609), .B(new_n14217_), .ZN(new_n14218_));
  AOI21_X1   g11782(.A1(new_n14218_), .A2(new_n14216_), .B(new_n12764_), .ZN(new_n14219_));
  AOI21_X1   g11783(.A1(new_n14219_), .A2(new_n14215_), .B(new_n14211_), .ZN(new_n14220_));
  OR2_X2     g11784(.A1(new_n14220_), .A2(pi0781), .Z(new_n14221_));
  NAND2_X1   g11785(.A1(new_n14086_), .A2(pi0627), .ZN(new_n14222_));
  INV_X1     g11786(.I(new_n14136_), .ZN(new_n14223_));
  AOI21_X1   g11787(.A1(new_n14223_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n14224_));
  NAND2_X1   g11788(.A1(new_n14220_), .A2(pi0618), .ZN(new_n14225_));
  AOI21_X1   g11789(.A1(new_n14225_), .A2(new_n14224_), .B(new_n14222_), .ZN(new_n14226_));
  NAND2_X1   g11790(.A1(new_n14089_), .A2(new_n12880_), .ZN(new_n14227_));
  AOI21_X1   g11791(.A1(new_n14223_), .A2(pi0618), .B(pi1154), .ZN(new_n14228_));
  INV_X1     g11792(.I(new_n14228_), .ZN(new_n14229_));
  AOI21_X1   g11793(.A1(new_n14220_), .A2(new_n12781_), .B(new_n14229_), .ZN(new_n14230_));
  OAI21_X1   g11794(.A1(new_n14230_), .A2(new_n14227_), .B(pi0781), .ZN(new_n14231_));
  OAI21_X1   g11795(.A1(new_n14231_), .A2(new_n14226_), .B(new_n14221_), .ZN(new_n14232_));
  AND2_X2    g11796(.A1(new_n14232_), .A2(new_n12796_), .Z(new_n14233_));
  AOI21_X1   g11797(.A1(new_n14138_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n14234_));
  OAI21_X1   g11798(.A1(new_n14232_), .A2(new_n12793_), .B(new_n14234_), .ZN(new_n14235_));
  NAND3_X1   g11799(.A1(new_n14235_), .A2(pi0648), .A3(new_n14094_), .ZN(new_n14236_));
  AOI21_X1   g11800(.A1(new_n14096_), .A2(pi1159), .B(pi0648), .ZN(new_n14237_));
  AOI21_X1   g11801(.A1(new_n14138_), .A2(pi0619), .B(pi1159), .ZN(new_n14238_));
  OAI21_X1   g11802(.A1(new_n14232_), .A2(pi0619), .B(new_n14238_), .ZN(new_n14239_));
  AOI21_X1   g11803(.A1(new_n14239_), .A2(new_n14237_), .B(new_n12796_), .ZN(new_n14240_));
  AOI21_X1   g11804(.A1(new_n14240_), .A2(new_n14236_), .B(new_n14233_), .ZN(new_n14241_));
  OAI21_X1   g11805(.A1(new_n14241_), .A2(new_n12747_), .B(new_n14162_), .ZN(new_n14242_));
  NAND2_X1   g11806(.A1(new_n14242_), .A2(new_n14161_), .ZN(new_n14243_));
  OAI21_X1   g11807(.A1(new_n14103_), .A2(pi1158), .B(new_n12904_), .ZN(new_n14244_));
  AOI21_X1   g11808(.A1(new_n14140_), .A2(pi0626), .B(pi0641), .ZN(new_n14245_));
  OAI21_X1   g11809(.A1(new_n14241_), .A2(pi0626), .B(new_n14245_), .ZN(new_n14246_));
  AOI21_X1   g11810(.A1(new_n14246_), .A2(new_n14244_), .B(new_n12808_), .ZN(new_n14247_));
  AND2_X2    g11811(.A1(new_n14241_), .A2(new_n12808_), .Z(new_n14248_));
  AOI21_X1   g11812(.A1(new_n14247_), .A2(new_n14243_), .B(new_n14248_), .ZN(new_n14249_));
  OAI21_X1   g11813(.A1(new_n14249_), .A2(new_n12920_), .B(new_n14160_), .ZN(new_n14250_));
  NAND3_X1   g11814(.A1(new_n14250_), .A2(pi0629), .A3(new_n14145_), .ZN(new_n14251_));
  NOR2_X1    g11815(.A1(new_n14148_), .A2(pi0629), .ZN(new_n14252_));
  AOI21_X1   g11816(.A1(new_n14105_), .A2(pi0628), .B(pi1156), .ZN(new_n14253_));
  OAI21_X1   g11817(.A1(new_n14249_), .A2(pi0628), .B(new_n14253_), .ZN(new_n14254_));
  AOI21_X1   g11818(.A1(new_n14254_), .A2(new_n14252_), .B(new_n12937_), .ZN(new_n14255_));
  AND2_X2    g11819(.A1(new_n14249_), .A2(new_n12937_), .Z(new_n14256_));
  AOI21_X1   g11820(.A1(new_n14255_), .A2(new_n14251_), .B(new_n14256_), .ZN(new_n14257_));
  OR2_X2     g11821(.A1(new_n14257_), .A2(pi0787), .Z(new_n14258_));
  OR2_X2     g11822(.A1(new_n14153_), .A2(new_n12981_), .Z(new_n14259_));
  NOR2_X1    g11823(.A1(new_n14107_), .A2(pi0647), .ZN(new_n14260_));
  NOR2_X1    g11824(.A1(new_n14260_), .A2(new_n12965_), .ZN(new_n14261_));
  NAND2_X1   g11825(.A1(new_n14257_), .A2(pi0647), .ZN(new_n14262_));
  AOI21_X1   g11826(.A1(new_n14262_), .A2(new_n14261_), .B(new_n14259_), .ZN(new_n14263_));
  NAND2_X1   g11827(.A1(new_n14156_), .A2(new_n12981_), .ZN(new_n14264_));
  OAI21_X1   g11828(.A1(new_n14107_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n14265_));
  AOI21_X1   g11829(.A1(new_n14257_), .A2(new_n12741_), .B(new_n14265_), .ZN(new_n14266_));
  OAI21_X1   g11830(.A1(new_n14266_), .A2(new_n14264_), .B(pi0787), .ZN(new_n14267_));
  OAI21_X1   g11831(.A1(new_n14267_), .A2(new_n14263_), .B(new_n14258_), .ZN(new_n14268_));
  OAI21_X1   g11832(.A1(new_n14268_), .A2(pi0644), .B(new_n14159_), .ZN(new_n14269_));
  NAND2_X1   g11833(.A1(new_n14269_), .A2(new_n14111_), .ZN(new_n14270_));
  AOI21_X1   g11834(.A1(new_n14052_), .A2(new_n12975_), .B(pi0715), .ZN(new_n14271_));
  NAND2_X1   g11835(.A1(new_n14109_), .A2(pi0644), .ZN(new_n14272_));
  AOI21_X1   g11836(.A1(new_n14272_), .A2(new_n14271_), .B(new_n12739_), .ZN(new_n14273_));
  NOR2_X1    g11837(.A1(new_n14158_), .A2(pi0644), .ZN(new_n14274_));
  AOI21_X1   g11838(.A1(new_n14268_), .A2(pi0644), .B(new_n14274_), .ZN(new_n14275_));
  OAI21_X1   g11839(.A1(new_n14275_), .A2(new_n12740_), .B(new_n14273_), .ZN(new_n14276_));
  NAND3_X1   g11840(.A1(new_n14276_), .A2(new_n14270_), .A3(pi0790), .ZN(new_n14277_));
  AOI21_X1   g11841(.A1(new_n14268_), .A2(new_n13000_), .B(po1038), .ZN(new_n14278_));
  NAND2_X1   g11842(.A1(new_n14277_), .A2(new_n14278_), .ZN(new_n14279_));
  AOI21_X1   g11843(.A1(new_n14279_), .A2(new_n14051_), .B(new_n14050_), .ZN(po0298));
  NOR2_X1    g11844(.A1(new_n3042_), .A2(new_n2724_), .ZN(new_n14281_));
  INV_X1     g11845(.I(new_n14281_), .ZN(new_n14282_));
  INV_X1     g11846(.I(pi0735), .ZN(new_n14283_));
  NOR2_X1    g11847(.A1(new_n12832_), .A2(new_n14283_), .ZN(new_n14284_));
  NOR2_X1    g11848(.A1(new_n14132_), .A2(new_n12758_), .ZN(new_n14285_));
  INV_X1     g11849(.I(new_n14285_), .ZN(new_n14286_));
  AOI21_X1   g11850(.A1(new_n14284_), .A2(new_n14286_), .B(new_n14281_), .ZN(new_n14287_));
  INV_X1     g11851(.I(new_n12923_), .ZN(new_n14288_));
  NOR2_X1    g11852(.A1(new_n12869_), .A2(new_n12887_), .ZN(new_n14289_));
  INV_X1     g11853(.I(new_n14289_), .ZN(new_n14290_));
  NOR2_X1    g11854(.A1(new_n14288_), .A2(new_n14290_), .ZN(new_n14291_));
  INV_X1     g11855(.I(new_n14291_), .ZN(new_n14292_));
  NOR2_X1    g11856(.A1(new_n14287_), .A2(new_n14292_), .ZN(new_n14293_));
  INV_X1     g11857(.I(new_n14293_), .ZN(new_n14294_));
  NOR2_X1    g11858(.A1(new_n14294_), .A2(new_n12951_), .ZN(new_n14295_));
  INV_X1     g11859(.I(new_n14295_), .ZN(new_n14296_));
  NOR2_X1    g11860(.A1(new_n12965_), .A2(pi0647), .ZN(new_n14297_));
  NOR2_X1    g11861(.A1(new_n12741_), .A2(pi1157), .ZN(new_n14298_));
  NOR2_X1    g11862(.A1(new_n14297_), .A2(new_n14298_), .ZN(new_n14299_));
  NOR2_X1    g11863(.A1(new_n14299_), .A2(new_n12972_), .ZN(new_n14300_));
  OAI21_X1   g11864(.A1(new_n14296_), .A2(new_n14300_), .B(new_n14282_), .ZN(new_n14301_));
  NOR2_X1    g11865(.A1(new_n14301_), .A2(new_n12975_), .ZN(new_n14302_));
  INV_X1     g11866(.I(new_n12819_), .ZN(new_n14303_));
  INV_X1     g11867(.I(pi0743), .ZN(new_n14304_));
  NOR2_X1    g11868(.A1(new_n13340_), .A2(new_n14304_), .ZN(new_n14305_));
  INV_X1     g11869(.I(new_n14305_), .ZN(new_n14306_));
  NOR2_X1    g11870(.A1(new_n14306_), .A2(new_n12760_), .ZN(new_n14307_));
  INV_X1     g11871(.I(new_n14307_), .ZN(new_n14308_));
  NOR2_X1    g11872(.A1(new_n14281_), .A2(pi0785), .ZN(new_n14309_));
  OAI21_X1   g11873(.A1(new_n14308_), .A2(new_n12766_), .B(pi1155), .ZN(new_n14310_));
  NOR2_X1    g11874(.A1(new_n14310_), .A2(new_n14281_), .ZN(new_n14311_));
  INV_X1     g11875(.I(new_n14311_), .ZN(new_n14312_));
  OAI21_X1   g11876(.A1(new_n14308_), .A2(pi0609), .B(new_n12770_), .ZN(new_n14313_));
  NOR2_X1    g11877(.A1(new_n14313_), .A2(new_n14281_), .ZN(new_n14314_));
  INV_X1     g11878(.I(new_n14314_), .ZN(new_n14315_));
  NAND2_X1   g11879(.A1(new_n14312_), .A2(new_n14315_), .ZN(new_n14316_));
  AOI22_X1   g11880(.A1(new_n14316_), .A2(pi0785), .B1(new_n14308_), .B2(new_n14309_), .ZN(new_n14317_));
  INV_X1     g11881(.I(new_n14317_), .ZN(new_n14318_));
  NAND2_X1   g11882(.A1(new_n14318_), .A2(pi0618), .ZN(new_n14319_));
  NAND2_X1   g11883(.A1(new_n14282_), .A2(new_n12781_), .ZN(new_n14320_));
  AOI21_X1   g11884(.A1(new_n14319_), .A2(new_n14320_), .B(new_n12785_), .ZN(new_n14321_));
  INV_X1     g11885(.I(new_n14287_), .ZN(new_n14322_));
  AOI21_X1   g11886(.A1(new_n14322_), .A2(new_n12870_), .B(new_n14281_), .ZN(new_n14323_));
  NAND2_X1   g11887(.A1(new_n14323_), .A2(pi0618), .ZN(new_n14324_));
  NOR2_X1    g11888(.A1(new_n14322_), .A2(new_n12766_), .ZN(new_n14325_));
  NAND2_X1   g11889(.A1(new_n13562_), .A2(pi0735), .ZN(new_n14326_));
  NAND3_X1   g11890(.A1(new_n14326_), .A2(new_n14306_), .A3(new_n14282_), .ZN(new_n14327_));
  INV_X1     g11891(.I(new_n13562_), .ZN(new_n14328_));
  NOR2_X1    g11892(.A1(new_n14328_), .A2(new_n13521_), .ZN(new_n14329_));
  INV_X1     g11893(.I(new_n14329_), .ZN(new_n14330_));
  OAI21_X1   g11894(.A1(new_n14330_), .A2(new_n14283_), .B(new_n14327_), .ZN(new_n14331_));
  INV_X1     g11895(.I(new_n14284_), .ZN(new_n14332_));
  OAI21_X1   g11896(.A1(new_n14332_), .A2(new_n13521_), .B(pi1153), .ZN(new_n14333_));
  OAI21_X1   g11897(.A1(new_n14333_), .A2(new_n14281_), .B(new_n13560_), .ZN(new_n14334_));
  AOI21_X1   g11898(.A1(new_n14331_), .A2(new_n12841_), .B(new_n14334_), .ZN(new_n14335_));
  AOI21_X1   g11899(.A1(new_n14284_), .A2(new_n14130_), .B(new_n14281_), .ZN(new_n14336_));
  OAI21_X1   g11900(.A1(new_n14330_), .A2(new_n14283_), .B(new_n14306_), .ZN(new_n14337_));
  NAND2_X1   g11901(.A1(new_n14337_), .A2(pi1153), .ZN(new_n14338_));
  AOI21_X1   g11902(.A1(new_n14338_), .A2(new_n14336_), .B(new_n13560_), .ZN(new_n14339_));
  NOR2_X1    g11903(.A1(new_n14339_), .A2(new_n14335_), .ZN(new_n14340_));
  NOR2_X1    g11904(.A1(new_n14327_), .A2(pi0778), .ZN(new_n14341_));
  AOI21_X1   g11905(.A1(new_n14340_), .A2(pi0778), .B(new_n14341_), .ZN(new_n14342_));
  INV_X1     g11906(.I(new_n14342_), .ZN(new_n14343_));
  AOI21_X1   g11907(.A1(new_n14343_), .A2(new_n12766_), .B(new_n14325_), .ZN(new_n14344_));
  OAI21_X1   g11908(.A1(new_n14344_), .A2(pi1155), .B(new_n14312_), .ZN(new_n14345_));
  NAND2_X1   g11909(.A1(new_n14343_), .A2(pi0609), .ZN(new_n14346_));
  NAND2_X1   g11910(.A1(new_n14287_), .A2(new_n12766_), .ZN(new_n14347_));
  AOI21_X1   g11911(.A1(new_n14346_), .A2(new_n14347_), .B(new_n12770_), .ZN(new_n14348_));
  NAND2_X1   g11912(.A1(new_n14315_), .A2(pi0660), .ZN(new_n14349_));
  OAI22_X1   g11913(.A1(new_n14345_), .A2(pi0660), .B1(new_n14348_), .B2(new_n14349_), .ZN(new_n14350_));
  NAND2_X1   g11914(.A1(new_n14343_), .A2(new_n12764_), .ZN(new_n14351_));
  OAI21_X1   g11915(.A1(new_n14350_), .A2(new_n12764_), .B(new_n14351_), .ZN(new_n14352_));
  NAND2_X1   g11916(.A1(new_n14352_), .A2(new_n12781_), .ZN(new_n14353_));
  AOI21_X1   g11917(.A1(new_n14353_), .A2(new_n14324_), .B(pi1154), .ZN(new_n14354_));
  NOR3_X1    g11918(.A1(new_n14354_), .A2(pi0627), .A3(new_n14321_), .ZN(new_n14355_));
  NAND2_X1   g11919(.A1(new_n14352_), .A2(pi0618), .ZN(new_n14356_));
  NAND2_X1   g11920(.A1(new_n14323_), .A2(new_n12781_), .ZN(new_n14357_));
  AOI21_X1   g11921(.A1(new_n14356_), .A2(new_n14357_), .B(new_n12785_), .ZN(new_n14358_));
  NAND2_X1   g11922(.A1(new_n14318_), .A2(new_n12781_), .ZN(new_n14359_));
  NAND2_X1   g11923(.A1(new_n14282_), .A2(pi0618), .ZN(new_n14360_));
  AOI21_X1   g11924(.A1(new_n14359_), .A2(new_n14360_), .B(pi1154), .ZN(new_n14361_));
  NOR3_X1    g11925(.A1(new_n14358_), .A2(new_n12880_), .A3(new_n14361_), .ZN(new_n14362_));
  OR3_X2     g11926(.A1(new_n14355_), .A2(new_n14362_), .A3(new_n12779_), .Z(new_n14363_));
  NAND2_X1   g11927(.A1(new_n14352_), .A2(new_n12779_), .ZN(new_n14364_));
  NAND2_X1   g11928(.A1(new_n14363_), .A2(new_n14364_), .ZN(new_n14365_));
  AOI21_X1   g11929(.A1(new_n14365_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n14366_));
  NOR3_X1    g11930(.A1(new_n14321_), .A2(new_n14361_), .A3(new_n12779_), .ZN(new_n14367_));
  AOI21_X1   g11931(.A1(new_n12779_), .A2(new_n14317_), .B(new_n14367_), .ZN(new_n14368_));
  NAND2_X1   g11932(.A1(new_n14368_), .A2(new_n12793_), .ZN(new_n14369_));
  NAND2_X1   g11933(.A1(new_n14282_), .A2(pi0619), .ZN(new_n14370_));
  AOI21_X1   g11934(.A1(new_n14369_), .A2(new_n14370_), .B(pi1159), .ZN(new_n14371_));
  NAND2_X1   g11935(.A1(new_n14365_), .A2(pi0619), .ZN(new_n14372_));
  AOI21_X1   g11936(.A1(new_n14322_), .A2(new_n14289_), .B(new_n14281_), .ZN(new_n14373_));
  NAND2_X1   g11937(.A1(new_n14373_), .A2(new_n12793_), .ZN(new_n14374_));
  AOI21_X1   g11938(.A1(new_n14372_), .A2(new_n14374_), .B(new_n12791_), .ZN(new_n14375_));
  NOR3_X1    g11939(.A1(new_n14375_), .A2(new_n12895_), .A3(new_n14371_), .ZN(new_n14376_));
  NAND2_X1   g11940(.A1(new_n14368_), .A2(pi0619), .ZN(new_n14377_));
  NAND2_X1   g11941(.A1(new_n14282_), .A2(new_n12793_), .ZN(new_n14378_));
  AOI21_X1   g11942(.A1(new_n14377_), .A2(new_n14378_), .B(new_n12791_), .ZN(new_n14379_));
  NAND2_X1   g11943(.A1(new_n14373_), .A2(pi0619), .ZN(new_n14380_));
  NAND2_X1   g11944(.A1(new_n14365_), .A2(new_n12793_), .ZN(new_n14381_));
  AOI21_X1   g11945(.A1(new_n14381_), .A2(new_n14380_), .B(pi1159), .ZN(new_n14382_));
  OR3_X2     g11946(.A1(new_n14382_), .A2(pi0648), .A3(new_n14379_), .Z(new_n14383_));
  NAND2_X1   g11947(.A1(new_n14383_), .A2(pi0789), .ZN(new_n14384_));
  OAI21_X1   g11948(.A1(new_n14384_), .A2(new_n14376_), .B(new_n14366_), .ZN(new_n14385_));
  INV_X1     g11949(.I(new_n12906_), .ZN(new_n14386_));
  OAI21_X1   g11950(.A1(new_n12911_), .A2(new_n14281_), .B(new_n14386_), .ZN(new_n14387_));
  NOR2_X1    g11951(.A1(new_n14373_), .A2(new_n14387_), .ZN(new_n14388_));
  OR2_X2     g11952(.A1(new_n14379_), .A2(new_n12796_), .Z(new_n14389_));
  OAI22_X1   g11953(.A1(new_n14389_), .A2(new_n14371_), .B1(pi0789), .B2(new_n14368_), .ZN(new_n14390_));
  NAND2_X1   g11954(.A1(new_n14390_), .A2(new_n12804_), .ZN(new_n14391_));
  OAI21_X1   g11955(.A1(new_n12749_), .A2(new_n14282_), .B(new_n14391_), .ZN(new_n14392_));
  AND2_X2    g11956(.A1(new_n14392_), .A2(new_n12914_), .Z(new_n14393_));
  OAI21_X1   g11957(.A1(new_n14393_), .A2(new_n14388_), .B(pi0788), .ZN(new_n14394_));
  NAND2_X1   g11958(.A1(new_n14385_), .A2(new_n14394_), .ZN(new_n14395_));
  INV_X1     g11959(.I(new_n14395_), .ZN(new_n14396_));
  NOR2_X1    g11960(.A1(new_n14396_), .A2(new_n12920_), .ZN(new_n14397_));
  NAND2_X1   g11961(.A1(new_n14392_), .A2(pi0788), .ZN(new_n14398_));
  NAND2_X1   g11962(.A1(new_n14390_), .A2(new_n12808_), .ZN(new_n14399_));
  NAND2_X1   g11963(.A1(new_n14398_), .A2(new_n14399_), .ZN(new_n14400_));
  AOI21_X1   g11964(.A1(new_n12920_), .A2(new_n14400_), .B(new_n14397_), .ZN(new_n14401_));
  OAI21_X1   g11965(.A1(new_n14294_), .A2(pi0628), .B(new_n14282_), .ZN(new_n14402_));
  AOI21_X1   g11966(.A1(new_n14402_), .A2(new_n12742_), .B(new_n12919_), .ZN(new_n14403_));
  OAI21_X1   g11967(.A1(new_n14401_), .A2(new_n12742_), .B(new_n14403_), .ZN(new_n14404_));
  NAND2_X1   g11968(.A1(new_n14400_), .A2(pi0628), .ZN(new_n14405_));
  OAI21_X1   g11969(.A1(new_n14396_), .A2(pi0628), .B(new_n14405_), .ZN(new_n14406_));
  NAND2_X1   g11970(.A1(new_n14406_), .A2(new_n12742_), .ZN(new_n14407_));
  OAI21_X1   g11971(.A1(new_n14294_), .A2(new_n12920_), .B(new_n14282_), .ZN(new_n14408_));
  NAND2_X1   g11972(.A1(new_n14408_), .A2(pi1156), .ZN(new_n14409_));
  AND3_X2    g11973(.A1(new_n14407_), .A2(new_n12919_), .A3(new_n14409_), .Z(new_n14410_));
  NOR2_X1    g11974(.A1(new_n14410_), .A2(new_n12937_), .ZN(new_n14411_));
  AOI22_X1   g11975(.A1(new_n14411_), .A2(new_n14404_), .B1(new_n12937_), .B2(new_n14395_), .ZN(new_n14412_));
  NAND2_X1   g11976(.A1(new_n14412_), .A2(new_n12972_), .ZN(new_n14413_));
  NOR2_X1    g11977(.A1(new_n14400_), .A2(new_n12943_), .ZN(new_n14414_));
  AOI21_X1   g11978(.A1(new_n12943_), .A2(new_n14282_), .B(new_n14414_), .ZN(new_n14415_));
  NOR2_X1    g11979(.A1(new_n14415_), .A2(pi0647), .ZN(new_n14416_));
  AOI21_X1   g11980(.A1(new_n14412_), .A2(pi0647), .B(new_n14416_), .ZN(new_n14417_));
  OAI21_X1   g11981(.A1(new_n14296_), .A2(pi0647), .B(new_n12965_), .ZN(new_n14418_));
  OAI22_X1   g11982(.A1(new_n14417_), .A2(new_n12965_), .B1(new_n14281_), .B2(new_n14418_), .ZN(new_n14419_));
  NAND2_X1   g11983(.A1(new_n14412_), .A2(new_n12741_), .ZN(new_n14420_));
  INV_X1     g11984(.I(new_n14415_), .ZN(new_n14421_));
  NAND2_X1   g11985(.A1(new_n14421_), .A2(pi0647), .ZN(new_n14422_));
  AOI21_X1   g11986(.A1(new_n14420_), .A2(new_n14422_), .B(pi1157), .ZN(new_n14423_));
  OAI21_X1   g11987(.A1(new_n14296_), .A2(new_n12741_), .B(pi1157), .ZN(new_n14424_));
  OAI21_X1   g11988(.A1(new_n14424_), .A2(new_n14281_), .B(new_n12981_), .ZN(new_n14425_));
  OAI22_X1   g11989(.A1(new_n14419_), .A2(new_n12981_), .B1(new_n14423_), .B2(new_n14425_), .ZN(new_n14426_));
  OAI21_X1   g11990(.A1(new_n14426_), .A2(new_n12972_), .B(new_n14413_), .ZN(new_n14427_));
  AND2_X2    g11991(.A1(new_n14427_), .A2(new_n12975_), .Z(new_n14428_));
  OAI21_X1   g11992(.A1(new_n14428_), .A2(new_n14302_), .B(new_n12740_), .ZN(new_n14429_));
  NAND2_X1   g11993(.A1(new_n12984_), .A2(new_n14281_), .ZN(new_n14430_));
  OAI21_X1   g11994(.A1(new_n14421_), .A2(new_n12984_), .B(new_n14430_), .ZN(new_n14431_));
  NOR2_X1    g11995(.A1(new_n14431_), .A2(pi0644), .ZN(new_n14432_));
  NOR2_X1    g11996(.A1(new_n14281_), .A2(new_n12975_), .ZN(new_n14433_));
  OAI21_X1   g11997(.A1(new_n14432_), .A2(new_n14433_), .B(pi0715), .ZN(new_n14434_));
  NAND3_X1   g11998(.A1(new_n14429_), .A2(new_n12739_), .A3(new_n14434_), .ZN(new_n14435_));
  NOR2_X1    g11999(.A1(new_n14301_), .A2(pi0644), .ZN(new_n14436_));
  AOI21_X1   g12000(.A1(new_n14427_), .A2(pi0644), .B(new_n14436_), .ZN(new_n14437_));
  NAND2_X1   g12001(.A1(new_n14282_), .A2(new_n12975_), .ZN(new_n14438_));
  OAI21_X1   g12002(.A1(new_n14431_), .A2(new_n12975_), .B(new_n14438_), .ZN(new_n14439_));
  AOI21_X1   g12003(.A1(new_n14439_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n14440_));
  OAI21_X1   g12004(.A1(new_n14437_), .A2(new_n12740_), .B(new_n14440_), .ZN(new_n14441_));
  NAND3_X1   g12005(.A1(new_n14435_), .A2(pi0790), .A3(new_n14441_), .ZN(new_n14442_));
  NAND2_X1   g12006(.A1(new_n14427_), .A2(new_n13000_), .ZN(new_n14443_));
  AOI21_X1   g12007(.A1(new_n14442_), .A2(new_n14443_), .B(new_n12738_), .ZN(new_n14444_));
  AOI21_X1   g12008(.A1(pi0057), .A2(pi0142), .B(pi0832), .ZN(new_n14445_));
  NOR2_X1    g12009(.A1(new_n13179_), .A2(new_n2724_), .ZN(new_n14446_));
  NAND2_X1   g12010(.A1(new_n14446_), .A2(new_n5422_), .ZN(new_n14447_));
  NOR2_X1    g12011(.A1(new_n13175_), .A2(new_n2724_), .ZN(new_n14448_));
  NAND2_X1   g12012(.A1(new_n14448_), .A2(new_n6764_), .ZN(new_n14449_));
  AOI21_X1   g12013(.A1(new_n14447_), .A2(new_n14449_), .B(new_n2436_), .ZN(new_n14450_));
  NOR2_X1    g12014(.A1(new_n13126_), .A2(new_n6764_), .ZN(new_n14451_));
  INV_X1     g12015(.I(new_n13093_), .ZN(new_n14452_));
  NOR2_X1    g12016(.A1(new_n14452_), .A2(new_n5422_), .ZN(new_n14453_));
  NOR3_X1    g12017(.A1(new_n14451_), .A2(new_n3303_), .A3(new_n14453_), .ZN(new_n14454_));
  NOR4_X1    g12018(.A1(new_n14454_), .A2(new_n2724_), .A3(pi0215), .A4(new_n13639_), .ZN(new_n14455_));
  OAI21_X1   g12019(.A1(new_n14455_), .A2(new_n14450_), .B(pi0299), .ZN(new_n14456_));
  OAI21_X1   g12020(.A1(new_n2627_), .A2(new_n13188_), .B(new_n13336_), .ZN(new_n14457_));
  OAI22_X1   g12021(.A1(new_n14457_), .A2(new_n2724_), .B1(new_n2627_), .B2(new_n14456_), .ZN(new_n14458_));
  AND2_X2    g12022(.A1(new_n14458_), .A2(new_n11503_), .Z(new_n14459_));
  NOR2_X1    g12023(.A1(new_n13005_), .A2(new_n2610_), .ZN(new_n14460_));
  NOR2_X1    g12024(.A1(new_n14460_), .A2(new_n2724_), .ZN(new_n14461_));
  NOR2_X1    g12025(.A1(new_n14459_), .A2(new_n14461_), .ZN(new_n14462_));
  INV_X1     g12026(.I(new_n14462_), .ZN(new_n14463_));
  NOR2_X1    g12027(.A1(new_n2609_), .A2(new_n2724_), .ZN(new_n14464_));
  AOI21_X1   g12028(.A1(pi0039), .A2(pi0142), .B(new_n3265_), .ZN(new_n14465_));
  NOR2_X1    g12029(.A1(new_n2530_), .A2(new_n14332_), .ZN(new_n14466_));
  NOR2_X1    g12030(.A1(new_n13136_), .A2(new_n2724_), .ZN(new_n14467_));
  OAI21_X1   g12031(.A1(new_n14467_), .A2(new_n14466_), .B(new_n2627_), .ZN(new_n14468_));
  AOI21_X1   g12032(.A1(new_n14468_), .A2(new_n14465_), .B(new_n2610_), .ZN(new_n14469_));
  INV_X1     g12033(.I(new_n14469_), .ZN(new_n14470_));
  NAND2_X1   g12034(.A1(new_n13405_), .A2(pi0142), .ZN(new_n14471_));
  OAI21_X1   g12035(.A1(pi0142), .A2(new_n13416_), .B(new_n14471_), .ZN(new_n14472_));
  NOR2_X1    g12036(.A1(new_n2724_), .A2(pi0735), .ZN(new_n14473_));
  AOI22_X1   g12037(.A1(new_n14472_), .A2(pi0735), .B1(new_n13060_), .B2(new_n14473_), .ZN(new_n14474_));
  OAI21_X1   g12038(.A1(new_n14474_), .A2(pi0039), .B(new_n3265_), .ZN(new_n14475_));
  NAND2_X1   g12039(.A1(new_n13473_), .A2(pi0142), .ZN(new_n14476_));
  NOR4_X1    g12040(.A1(new_n13422_), .A2(new_n13423_), .A3(pi0142), .A4(new_n12821_), .ZN(new_n14477_));
  NOR2_X1    g12041(.A1(new_n14477_), .A2(new_n14283_), .ZN(new_n14478_));
  NAND2_X1   g12042(.A1(new_n14476_), .A2(new_n14478_), .ZN(new_n14479_));
  OAI21_X1   g12043(.A1(new_n14446_), .A2(pi0735), .B(new_n14479_), .ZN(new_n14480_));
  OR2_X2     g12044(.A1(new_n14480_), .A2(new_n6764_), .Z(new_n14481_));
  INV_X1     g12045(.I(new_n14448_), .ZN(new_n14482_));
  OAI21_X1   g12046(.A1(new_n13468_), .A2(new_n13461_), .B(pi0142), .ZN(new_n14483_));
  AOI21_X1   g12047(.A1(new_n14477_), .A2(new_n13578_), .B(new_n14283_), .ZN(new_n14484_));
  AOI22_X1   g12048(.A1(new_n14482_), .A2(new_n14283_), .B1(new_n14483_), .B2(new_n14484_), .ZN(new_n14485_));
  NAND2_X1   g12049(.A1(new_n14485_), .A2(new_n6764_), .ZN(new_n14486_));
  AOI21_X1   g12050(.A1(new_n14481_), .A2(new_n14486_), .B(new_n2436_), .ZN(new_n14487_));
  NOR2_X1    g12051(.A1(new_n13098_), .A2(new_n2724_), .ZN(new_n14488_));
  AOI21_X1   g12052(.A1(new_n13087_), .A2(new_n14284_), .B(new_n14488_), .ZN(new_n14489_));
  AOI21_X1   g12053(.A1(new_n14489_), .A2(new_n3303_), .B(pi0215), .ZN(new_n14490_));
  INV_X1     g12054(.I(new_n14490_), .ZN(new_n14491_));
  INV_X1     g12055(.I(new_n14473_), .ZN(new_n14492_));
  NOR2_X1    g12056(.A1(new_n13438_), .A2(new_n13435_), .ZN(new_n14493_));
  AND2_X2    g12057(.A1(new_n13494_), .A2(pi0142), .Z(new_n14494_));
  AOI22_X1   g12058(.A1(new_n14494_), .A2(new_n13497_), .B1(new_n2724_), .B2(new_n14493_), .ZN(new_n14495_));
  OAI22_X1   g12059(.A1(new_n14495_), .A2(new_n14283_), .B1(new_n13126_), .B2(new_n14492_), .ZN(new_n14496_));
  NAND2_X1   g12060(.A1(new_n13487_), .A2(pi0142), .ZN(new_n14497_));
  OR2_X2     g12061(.A1(new_n13431_), .A2(pi0142), .Z(new_n14498_));
  NAND2_X1   g12062(.A1(new_n14497_), .A2(new_n14498_), .ZN(new_n14499_));
  NOR2_X1    g12063(.A1(new_n14452_), .A2(new_n14492_), .ZN(new_n14500_));
  AOI21_X1   g12064(.A1(new_n14499_), .A2(pi0735), .B(new_n14500_), .ZN(new_n14501_));
  NAND2_X1   g12065(.A1(new_n14501_), .A2(new_n6764_), .ZN(new_n14502_));
  OAI21_X1   g12066(.A1(new_n14496_), .A2(new_n6764_), .B(new_n14502_), .ZN(new_n14503_));
  AOI21_X1   g12067(.A1(new_n14503_), .A2(new_n3304_), .B(new_n14491_), .ZN(new_n14504_));
  NOR3_X1    g12068(.A1(new_n14504_), .A2(new_n2628_), .A3(new_n14487_), .ZN(new_n14505_));
  OR2_X2     g12069(.A1(new_n14480_), .A2(new_n5445_), .Z(new_n14506_));
  NAND2_X1   g12070(.A1(new_n14485_), .A2(new_n5445_), .ZN(new_n14507_));
  AOI21_X1   g12071(.A1(new_n14506_), .A2(new_n14507_), .B(new_n2668_), .ZN(new_n14508_));
  NAND2_X1   g12072(.A1(new_n14501_), .A2(new_n5445_), .ZN(new_n14509_));
  OAI21_X1   g12073(.A1(new_n14496_), .A2(new_n5445_), .B(new_n14509_), .ZN(new_n14510_));
  AOI21_X1   g12074(.A1(new_n14489_), .A2(new_n2641_), .B(pi0223), .ZN(new_n14511_));
  INV_X1     g12075(.I(new_n14511_), .ZN(new_n14512_));
  AOI21_X1   g12076(.A1(new_n14510_), .A2(new_n2642_), .B(new_n14512_), .ZN(new_n14513_));
  NOR3_X1    g12077(.A1(new_n14513_), .A2(pi0299), .A3(new_n14508_), .ZN(new_n14514_));
  NOR3_X1    g12078(.A1(new_n14505_), .A2(new_n14514_), .A3(new_n2627_), .ZN(new_n14515_));
  NOR2_X1    g12079(.A1(new_n14515_), .A2(new_n14475_), .ZN(new_n14516_));
  NOR2_X1    g12080(.A1(new_n14516_), .A2(new_n14470_), .ZN(new_n14517_));
  NOR2_X1    g12081(.A1(new_n14517_), .A2(new_n14464_), .ZN(new_n14518_));
  AOI21_X1   g12082(.A1(new_n14462_), .A2(pi0625), .B(pi1153), .ZN(new_n14519_));
  NOR2_X1    g12083(.A1(new_n14464_), .A2(pi0625), .ZN(new_n14520_));
  INV_X1     g12084(.I(new_n14520_), .ZN(new_n14521_));
  OAI21_X1   g12085(.A1(new_n14517_), .A2(new_n14521_), .B(new_n14519_), .ZN(new_n14522_));
  AOI21_X1   g12086(.A1(new_n14462_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n14523_));
  NOR2_X1    g12087(.A1(new_n14464_), .A2(new_n13521_), .ZN(new_n14524_));
  OAI21_X1   g12088(.A1(new_n14516_), .A2(new_n14470_), .B(new_n14524_), .ZN(new_n14525_));
  AOI21_X1   g12089(.A1(new_n14525_), .A2(new_n14523_), .B(new_n12758_), .ZN(new_n14526_));
  AOI22_X1   g12090(.A1(new_n14526_), .A2(new_n14522_), .B1(new_n12758_), .B2(new_n14518_), .ZN(new_n14527_));
  NOR2_X1    g12091(.A1(new_n14462_), .A2(new_n12870_), .ZN(new_n14528_));
  AOI21_X1   g12092(.A1(new_n14527_), .A2(new_n12870_), .B(new_n14528_), .ZN(new_n14529_));
  NOR2_X1    g12093(.A1(new_n14463_), .A2(new_n12888_), .ZN(new_n14530_));
  AOI21_X1   g12094(.A1(new_n14529_), .A2(new_n12888_), .B(new_n14530_), .ZN(new_n14531_));
  NOR2_X1    g12095(.A1(new_n14462_), .A2(new_n12911_), .ZN(new_n14532_));
  AOI21_X1   g12096(.A1(new_n14531_), .A2(new_n12911_), .B(new_n14532_), .ZN(new_n14533_));
  NOR2_X1    g12097(.A1(new_n14533_), .A2(new_n12817_), .ZN(new_n14534_));
  AOI21_X1   g12098(.A1(new_n12817_), .A2(new_n14463_), .B(new_n14534_), .ZN(new_n14535_));
  INV_X1     g12099(.I(new_n14535_), .ZN(new_n14536_));
  NAND2_X1   g12100(.A1(new_n14536_), .A2(new_n12920_), .ZN(new_n14537_));
  NAND2_X1   g12101(.A1(new_n14463_), .A2(pi0628), .ZN(new_n14538_));
  AOI21_X1   g12102(.A1(new_n14537_), .A2(new_n14538_), .B(pi1156), .ZN(new_n14539_));
  OR2_X2     g12103(.A1(new_n14539_), .A2(new_n12919_), .Z(new_n14540_));
  INV_X1     g12104(.I(new_n14464_), .ZN(new_n14541_));
  AOI21_X1   g12105(.A1(new_n2531_), .A2(new_n14305_), .B(new_n14467_), .ZN(new_n14542_));
  OAI21_X1   g12106(.A1(new_n14542_), .A2(pi0039), .B(new_n14465_), .ZN(new_n14543_));
  NAND2_X1   g12107(.A1(new_n14543_), .A2(new_n2609_), .ZN(new_n14544_));
  INV_X1     g12108(.I(new_n14544_), .ZN(new_n14545_));
  NOR2_X1    g12109(.A1(new_n13206_), .A2(new_n12751_), .ZN(new_n14546_));
  NAND2_X1   g12110(.A1(new_n13251_), .A2(new_n13254_), .ZN(new_n14547_));
  NOR2_X1    g12111(.A1(new_n14547_), .A2(new_n2724_), .ZN(new_n14548_));
  AOI21_X1   g12112(.A1(new_n2724_), .A2(new_n14546_), .B(new_n14548_), .ZN(new_n14549_));
  NOR2_X1    g12113(.A1(new_n2724_), .A2(pi0743), .ZN(new_n14550_));
  AOI21_X1   g12114(.A1(new_n13058_), .A2(new_n14550_), .B(pi0299), .ZN(new_n14551_));
  OAI21_X1   g12115(.A1(new_n14549_), .A2(new_n14304_), .B(new_n14551_), .ZN(new_n14552_));
  NOR2_X1    g12116(.A1(new_n13201_), .A2(new_n12751_), .ZN(new_n14553_));
  INV_X1     g12117(.I(new_n14553_), .ZN(new_n14554_));
  NAND2_X1   g12118(.A1(new_n14554_), .A2(new_n2724_), .ZN(new_n14555_));
  AOI22_X1   g12119(.A1(new_n14555_), .A2(pi0743), .B1(pi0142), .B2(new_n13055_), .ZN(new_n14556_));
  INV_X1     g12120(.I(new_n13055_), .ZN(new_n14557_));
  INV_X1     g12121(.I(new_n13803_), .ZN(new_n14558_));
  OAI21_X1   g12122(.A1(new_n12751_), .A2(new_n14558_), .B(new_n14557_), .ZN(new_n14559_));
  NOR2_X1    g12123(.A1(new_n14559_), .A2(new_n2724_), .ZN(new_n14560_));
  OAI21_X1   g12124(.A1(new_n14556_), .A2(new_n14560_), .B(pi0299), .ZN(new_n14561_));
  NAND3_X1   g12125(.A1(new_n14561_), .A2(new_n2627_), .A3(new_n14552_), .ZN(new_n14562_));
  NAND2_X1   g12126(.A1(new_n14562_), .A2(new_n3265_), .ZN(new_n14563_));
  OAI21_X1   g12127(.A1(new_n13179_), .A2(new_n2724_), .B(new_n14304_), .ZN(new_n14564_));
  NOR2_X1    g12128(.A1(new_n13217_), .A2(new_n14304_), .ZN(new_n14565_));
  OAI21_X1   g12129(.A1(new_n2724_), .A2(new_n13272_), .B(new_n14565_), .ZN(new_n14566_));
  NAND2_X1   g12130(.A1(new_n14566_), .A2(new_n14564_), .ZN(new_n14567_));
  NOR2_X1    g12131(.A1(new_n14567_), .A2(new_n5445_), .ZN(new_n14568_));
  NOR2_X1    g12132(.A1(new_n14448_), .A2(pi0743), .ZN(new_n14569_));
  NOR2_X1    g12133(.A1(new_n13281_), .A2(new_n2724_), .ZN(new_n14570_));
  NOR3_X1    g12134(.A1(new_n14570_), .A2(new_n14304_), .A3(new_n13581_), .ZN(new_n14571_));
  NOR2_X1    g12135(.A1(new_n14569_), .A2(new_n14571_), .ZN(new_n14572_));
  AOI21_X1   g12136(.A1(new_n5445_), .A2(new_n14572_), .B(new_n14568_), .ZN(new_n14573_));
  NAND2_X1   g12137(.A1(new_n13231_), .A2(new_n2724_), .ZN(new_n14574_));
  OR3_X2     g12138(.A1(new_n13294_), .A2(new_n2724_), .A3(new_n13306_), .Z(new_n14575_));
  NAND3_X1   g12139(.A1(new_n14575_), .A2(pi0743), .A3(new_n14574_), .ZN(new_n14576_));
  INV_X1     g12140(.I(new_n13126_), .ZN(new_n14577_));
  NAND2_X1   g12141(.A1(new_n14577_), .A2(new_n14550_), .ZN(new_n14578_));
  NAND2_X1   g12142(.A1(new_n14578_), .A2(new_n14576_), .ZN(new_n14579_));
  NOR2_X1    g12143(.A1(new_n14579_), .A2(new_n5445_), .ZN(new_n14580_));
  OAI21_X1   g12144(.A1(new_n13318_), .A2(new_n13308_), .B(pi0142), .ZN(new_n14581_));
  AND3_X2    g12145(.A1(new_n14581_), .A2(pi0743), .A3(new_n13239_), .Z(new_n14582_));
  AOI21_X1   g12146(.A1(new_n13093_), .A2(pi0142), .B(pi0743), .ZN(new_n14583_));
  NOR2_X1    g12147(.A1(new_n14582_), .A2(new_n14583_), .ZN(new_n14584_));
  NOR2_X1    g12148(.A1(new_n14584_), .A2(new_n5446_), .ZN(new_n14585_));
  OAI21_X1   g12149(.A1(new_n14585_), .A2(new_n14580_), .B(new_n2642_), .ZN(new_n14586_));
  AOI21_X1   g12150(.A1(new_n13210_), .A2(pi0743), .B(new_n14488_), .ZN(new_n14587_));
  AOI21_X1   g12151(.A1(new_n14587_), .A2(new_n2641_), .B(pi0223), .ZN(new_n14588_));
  AOI21_X1   g12152(.A1(new_n14586_), .A2(new_n14588_), .B(pi0299), .ZN(new_n14589_));
  OAI21_X1   g12153(.A1(new_n2668_), .A2(new_n14573_), .B(new_n14589_), .ZN(new_n14590_));
  INV_X1     g12154(.I(new_n14587_), .ZN(new_n14591_));
  NOR2_X1    g12155(.A1(new_n14591_), .A2(new_n3304_), .ZN(new_n14592_));
  INV_X1     g12156(.I(new_n14592_), .ZN(new_n14593_));
  NOR2_X1    g12157(.A1(new_n14579_), .A2(new_n6764_), .ZN(new_n14594_));
  NOR2_X1    g12158(.A1(new_n14584_), .A2(new_n5422_), .ZN(new_n14595_));
  OAI21_X1   g12159(.A1(new_n14595_), .A2(new_n14594_), .B(new_n3304_), .ZN(new_n14596_));
  AOI21_X1   g12160(.A1(new_n14596_), .A2(new_n14593_), .B(pi0215), .ZN(new_n14597_));
  INV_X1     g12161(.I(new_n14572_), .ZN(new_n14598_));
  NAND2_X1   g12162(.A1(new_n14598_), .A2(new_n6764_), .ZN(new_n14599_));
  NAND2_X1   g12163(.A1(new_n14567_), .A2(new_n5422_), .ZN(new_n14600_));
  AOI21_X1   g12164(.A1(new_n14599_), .A2(new_n14600_), .B(new_n2436_), .ZN(new_n14601_));
  OAI21_X1   g12165(.A1(new_n14597_), .A2(new_n14601_), .B(pi0299), .ZN(new_n14602_));
  AND3_X2    g12166(.A1(new_n14590_), .A2(pi0039), .A3(new_n14602_), .Z(new_n14603_));
  OAI21_X1   g12167(.A1(new_n14603_), .A2(new_n14563_), .B(new_n14545_), .ZN(new_n14604_));
  AOI21_X1   g12168(.A1(new_n14604_), .A2(new_n14541_), .B(new_n12760_), .ZN(new_n14605_));
  NOR2_X1    g12169(.A1(new_n14462_), .A2(new_n12761_), .ZN(new_n14606_));
  NOR3_X1    g12170(.A1(new_n14605_), .A2(pi0785), .A3(new_n14606_), .ZN(new_n14607_));
  INV_X1     g12171(.I(new_n14607_), .ZN(new_n14608_));
  AOI22_X1   g12172(.A1(new_n14605_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n14463_), .ZN(new_n14609_));
  OR2_X2     g12173(.A1(new_n14609_), .A2(pi1155), .Z(new_n14610_));
  AOI22_X1   g12174(.A1(new_n14605_), .A2(pi0609), .B1(new_n13357_), .B2(new_n14463_), .ZN(new_n14611_));
  NOR2_X1    g12175(.A1(new_n14611_), .A2(new_n12770_), .ZN(new_n14612_));
  NOR2_X1    g12176(.A1(new_n14612_), .A2(new_n12764_), .ZN(new_n14613_));
  NAND2_X1   g12177(.A1(new_n14613_), .A2(new_n14610_), .ZN(new_n14614_));
  NAND2_X1   g12178(.A1(new_n14614_), .A2(new_n14608_), .ZN(new_n14615_));
  NAND2_X1   g12179(.A1(new_n14463_), .A2(pi0618), .ZN(new_n14616_));
  OAI21_X1   g12180(.A1(new_n14615_), .A2(pi0618), .B(new_n14616_), .ZN(new_n14617_));
  NAND2_X1   g12181(.A1(new_n14617_), .A2(new_n12785_), .ZN(new_n14618_));
  NAND2_X1   g12182(.A1(new_n14463_), .A2(new_n12781_), .ZN(new_n14619_));
  OAI21_X1   g12183(.A1(new_n14615_), .A2(new_n12781_), .B(new_n14619_), .ZN(new_n14620_));
  AOI21_X1   g12184(.A1(new_n14620_), .A2(pi1154), .B(new_n12779_), .ZN(new_n14621_));
  AOI22_X1   g12185(.A1(new_n14621_), .A2(new_n14618_), .B1(new_n12779_), .B2(new_n14615_), .ZN(new_n14622_));
  NOR2_X1    g12186(.A1(new_n14462_), .A2(new_n12793_), .ZN(new_n14623_));
  AOI21_X1   g12187(.A1(new_n14622_), .A2(new_n12793_), .B(new_n14623_), .ZN(new_n14624_));
  NOR2_X1    g12188(.A1(new_n14624_), .A2(pi1159), .ZN(new_n14625_));
  NOR2_X1    g12189(.A1(new_n14462_), .A2(pi0619), .ZN(new_n14626_));
  AOI21_X1   g12190(.A1(new_n14622_), .A2(pi0619), .B(new_n14626_), .ZN(new_n14627_));
  OAI21_X1   g12191(.A1(new_n14627_), .A2(new_n12791_), .B(pi0789), .ZN(new_n14628_));
  OAI22_X1   g12192(.A1(new_n14628_), .A2(new_n14625_), .B1(pi0789), .B2(new_n14622_), .ZN(new_n14629_));
  NAND2_X1   g12193(.A1(new_n14463_), .A2(new_n12747_), .ZN(new_n14630_));
  OAI21_X1   g12194(.A1(new_n14629_), .A2(new_n12747_), .B(new_n14630_), .ZN(new_n14631_));
  NAND2_X1   g12195(.A1(new_n14631_), .A2(pi1158), .ZN(new_n14632_));
  NOR2_X1    g12196(.A1(new_n14462_), .A2(new_n12747_), .ZN(new_n14633_));
  INV_X1     g12197(.I(new_n14633_), .ZN(new_n14634_));
  OAI21_X1   g12198(.A1(new_n14629_), .A2(pi0626), .B(new_n14634_), .ZN(new_n14635_));
  AOI21_X1   g12199(.A1(new_n14635_), .A2(new_n12745_), .B(new_n12808_), .ZN(new_n14636_));
  AOI22_X1   g12200(.A1(new_n14636_), .A2(new_n14632_), .B1(new_n12808_), .B2(new_n14629_), .ZN(new_n14637_));
  NOR2_X1    g12201(.A1(new_n14637_), .A2(pi0628), .ZN(new_n14638_));
  NOR2_X1    g12202(.A1(new_n14638_), .A2(new_n12742_), .ZN(new_n14639_));
  NAND2_X1   g12203(.A1(new_n14525_), .A2(new_n14523_), .ZN(new_n14640_));
  AOI21_X1   g12204(.A1(new_n14604_), .A2(new_n14524_), .B(pi1153), .ZN(new_n14641_));
  INV_X1     g12205(.I(new_n14542_), .ZN(new_n14642_));
  INV_X1     g12206(.I(new_n13573_), .ZN(new_n14643_));
  NOR2_X1    g12207(.A1(new_n14643_), .A2(new_n14283_), .ZN(new_n14644_));
  OAI21_X1   g12208(.A1(new_n14644_), .A2(new_n14642_), .B(new_n2627_), .ZN(new_n14645_));
  AOI21_X1   g12209(.A1(new_n14645_), .A2(new_n14465_), .B(new_n2610_), .ZN(new_n14646_));
  INV_X1     g12210(.I(new_n14646_), .ZN(new_n14647_));
  AOI21_X1   g12211(.A1(new_n14561_), .A2(new_n14552_), .B(pi0735), .ZN(new_n14648_));
  NOR2_X1    g12212(.A1(new_n13403_), .A2(new_n13055_), .ZN(new_n14649_));
  NAND2_X1   g12213(.A1(new_n14554_), .A2(pi0142), .ZN(new_n14650_));
  OAI21_X1   g12214(.A1(new_n14650_), .A2(new_n14649_), .B(new_n14304_), .ZN(new_n14651_));
  NAND2_X1   g12215(.A1(new_n13804_), .A2(pi0680), .ZN(new_n14652_));
  NOR2_X1    g12216(.A1(new_n14652_), .A2(pi0142), .ZN(new_n14653_));
  OAI21_X1   g12217(.A1(new_n14651_), .A2(new_n14653_), .B(pi0299), .ZN(new_n14654_));
  INV_X1     g12218(.I(new_n13411_), .ZN(new_n14655_));
  NAND2_X1   g12219(.A1(new_n14655_), .A2(pi0680), .ZN(new_n14656_));
  NAND3_X1   g12220(.A1(new_n14554_), .A2(new_n14656_), .A3(new_n2724_), .ZN(new_n14657_));
  OR3_X2     g12221(.A1(new_n14559_), .A2(new_n2724_), .A3(new_n13403_), .Z(new_n14658_));
  AOI21_X1   g12222(.A1(new_n14658_), .A2(new_n14657_), .B(new_n14304_), .ZN(new_n14659_));
  NOR2_X1    g12223(.A1(new_n14654_), .A2(new_n14659_), .ZN(new_n14660_));
  NOR2_X1    g12224(.A1(new_n13401_), .A2(new_n13058_), .ZN(new_n14661_));
  NOR3_X1    g12225(.A1(new_n14661_), .A2(new_n14546_), .A3(new_n2724_), .ZN(new_n14662_));
  NAND2_X1   g12226(.A1(new_n13806_), .A2(pi0680), .ZN(new_n14663_));
  NOR2_X1    g12227(.A1(new_n14663_), .A2(pi0142), .ZN(new_n14664_));
  NOR3_X1    g12228(.A1(new_n14664_), .A2(pi0743), .A3(new_n14662_), .ZN(new_n14665_));
  INV_X1     g12229(.I(new_n14546_), .ZN(new_n14666_));
  INV_X1     g12230(.I(new_n13414_), .ZN(new_n14667_));
  NAND2_X1   g12231(.A1(new_n14667_), .A2(pi0680), .ZN(new_n14668_));
  NAND3_X1   g12232(.A1(new_n14668_), .A2(new_n14666_), .A3(new_n2724_), .ZN(new_n14669_));
  NAND3_X1   g12233(.A1(new_n14547_), .A2(new_n14661_), .A3(pi0142), .ZN(new_n14670_));
  AOI21_X1   g12234(.A1(new_n14669_), .A2(new_n14670_), .B(new_n14304_), .ZN(new_n14671_));
  NOR3_X1    g12235(.A1(new_n14665_), .A2(new_n14671_), .A3(pi0299), .ZN(new_n14672_));
  NOR3_X1    g12236(.A1(new_n14660_), .A2(new_n14283_), .A3(new_n14672_), .ZN(new_n14673_));
  OAI21_X1   g12237(.A1(new_n14673_), .A2(new_n14648_), .B(new_n2627_), .ZN(new_n14674_));
  OR3_X2     g12238(.A1(new_n13717_), .A2(new_n13711_), .A3(new_n13718_), .Z(new_n14675_));
  AND2_X2    g12239(.A1(new_n13783_), .A2(new_n2724_), .Z(new_n14676_));
  AOI21_X1   g12240(.A1(pi0142), .A2(new_n14675_), .B(new_n14676_), .ZN(new_n14677_));
  OAI21_X1   g12241(.A1(new_n13655_), .A2(new_n13657_), .B(pi0142), .ZN(new_n14678_));
  OAI21_X1   g12242(.A1(new_n13582_), .A2(pi0142), .B(new_n14678_), .ZN(new_n14679_));
  AOI21_X1   g12243(.A1(new_n14679_), .A2(pi0743), .B(new_n14283_), .ZN(new_n14680_));
  OAI21_X1   g12244(.A1(new_n14677_), .A2(pi0743), .B(new_n14680_), .ZN(new_n14681_));
  NAND2_X1   g12245(.A1(new_n14598_), .A2(new_n14283_), .ZN(new_n14682_));
  NAND3_X1   g12246(.A1(new_n14681_), .A2(new_n14682_), .A3(new_n5445_), .ZN(new_n14683_));
  OR2_X2     g12247(.A1(new_n13709_), .A2(new_n13696_), .Z(new_n14684_));
  AOI21_X1   g12248(.A1(new_n13775_), .A2(new_n13776_), .B(pi0142), .ZN(new_n14685_));
  AOI21_X1   g12249(.A1(new_n14684_), .A2(pi0142), .B(new_n14685_), .ZN(new_n14686_));
  NAND3_X1   g12250(.A1(new_n13661_), .A2(pi0142), .A3(new_n13660_), .ZN(new_n14687_));
  OAI21_X1   g12251(.A1(new_n13593_), .A2(pi0142), .B(new_n14687_), .ZN(new_n14688_));
  AOI21_X1   g12252(.A1(new_n14688_), .A2(pi0743), .B(new_n14283_), .ZN(new_n14689_));
  OAI21_X1   g12253(.A1(new_n14686_), .A2(pi0743), .B(new_n14689_), .ZN(new_n14690_));
  NAND2_X1   g12254(.A1(new_n14567_), .A2(new_n14283_), .ZN(new_n14691_));
  NAND3_X1   g12255(.A1(new_n14690_), .A2(new_n5446_), .A3(new_n14691_), .ZN(new_n14692_));
  AOI21_X1   g12256(.A1(new_n14692_), .A2(new_n14683_), .B(new_n2668_), .ZN(new_n14693_));
  NOR2_X1    g12257(.A1(new_n14579_), .A2(pi0735), .ZN(new_n14694_));
  OR2_X2     g12258(.A1(new_n13668_), .A2(new_n13669_), .Z(new_n14695_));
  OAI21_X1   g12259(.A1(new_n14695_), .A2(new_n13664_), .B(pi0142), .ZN(new_n14696_));
  NAND4_X1   g12260(.A1(new_n13631_), .A2(new_n13624_), .A3(new_n13619_), .A4(new_n2724_), .ZN(new_n14697_));
  AOI21_X1   g12261(.A1(new_n14696_), .A2(new_n14697_), .B(new_n14304_), .ZN(new_n14698_));
  NOR2_X1    g12262(.A1(new_n13764_), .A2(pi0142), .ZN(new_n14699_));
  NOR2_X1    g12263(.A1(new_n14699_), .A2(pi0743), .ZN(new_n14700_));
  OR3_X2     g12264(.A1(new_n13734_), .A2(new_n2724_), .A3(new_n13739_), .Z(new_n14701_));
  AOI21_X1   g12265(.A1(new_n14701_), .A2(new_n14700_), .B(new_n14698_), .ZN(new_n14702_));
  AOI21_X1   g12266(.A1(new_n14702_), .A2(pi0735), .B(new_n14694_), .ZN(new_n14703_));
  NAND3_X1   g12267(.A1(new_n13771_), .A2(new_n2724_), .A3(new_n13767_), .ZN(new_n14704_));
  NAND2_X1   g12268(.A1(new_n13725_), .A2(pi0142), .ZN(new_n14705_));
  AOI21_X1   g12269(.A1(new_n14704_), .A2(new_n14705_), .B(pi0743), .ZN(new_n14706_));
  OAI21_X1   g12270(.A1(new_n13674_), .A2(new_n13675_), .B(pi0142), .ZN(new_n14707_));
  INV_X1     g12271(.I(new_n13429_), .ZN(new_n14708_));
  NAND3_X1   g12272(.A1(new_n13239_), .A2(new_n14708_), .A3(new_n13585_), .ZN(new_n14709_));
  NAND2_X1   g12273(.A1(new_n13291_), .A2(new_n12822_), .ZN(new_n14710_));
  NAND3_X1   g12274(.A1(new_n13311_), .A2(new_n14710_), .A3(pi0603), .ZN(new_n14711_));
  AOI21_X1   g12275(.A1(new_n13768_), .A2(new_n14711_), .B(new_n13264_), .ZN(new_n14712_));
  AOI21_X1   g12276(.A1(new_n13617_), .A2(new_n13603_), .B(new_n5408_), .ZN(new_n14713_));
  OAI21_X1   g12277(.A1(new_n14712_), .A2(new_n14713_), .B(new_n13584_), .ZN(new_n14714_));
  NAND3_X1   g12278(.A1(new_n14714_), .A2(new_n2724_), .A3(new_n14709_), .ZN(new_n14715_));
  AOI21_X1   g12279(.A1(new_n14715_), .A2(new_n14707_), .B(new_n14304_), .ZN(new_n14716_));
  NOR3_X1    g12280(.A1(new_n14706_), .A2(new_n14716_), .A3(new_n14283_), .ZN(new_n14717_));
  NOR2_X1    g12281(.A1(new_n14584_), .A2(pi0735), .ZN(new_n14718_));
  OAI21_X1   g12282(.A1(new_n14718_), .A2(new_n14717_), .B(new_n5445_), .ZN(new_n14719_));
  OAI21_X1   g12283(.A1(new_n14703_), .A2(new_n5445_), .B(new_n14719_), .ZN(new_n14720_));
  OAI21_X1   g12284(.A1(new_n14642_), .A2(new_n13573_), .B(new_n13679_), .ZN(new_n14721_));
  NAND2_X1   g12285(.A1(new_n14721_), .A2(pi0735), .ZN(new_n14722_));
  OAI22_X1   g12286(.A1(new_n14591_), .A2(pi0735), .B1(new_n14488_), .B2(new_n14722_), .ZN(new_n14723_));
  AOI21_X1   g12287(.A1(new_n14723_), .A2(new_n2641_), .B(pi0223), .ZN(new_n14724_));
  INV_X1     g12288(.I(new_n14724_), .ZN(new_n14725_));
  AOI21_X1   g12289(.A1(new_n14720_), .A2(new_n2642_), .B(new_n14725_), .ZN(new_n14726_));
  OAI21_X1   g12290(.A1(new_n14726_), .A2(new_n14693_), .B(new_n2628_), .ZN(new_n14727_));
  NAND3_X1   g12291(.A1(new_n14681_), .A2(new_n14682_), .A3(new_n6764_), .ZN(new_n14728_));
  NAND3_X1   g12292(.A1(new_n14690_), .A2(new_n5422_), .A3(new_n14691_), .ZN(new_n14729_));
  AOI21_X1   g12293(.A1(new_n14729_), .A2(new_n14728_), .B(new_n2436_), .ZN(new_n14730_));
  NAND2_X1   g12294(.A1(new_n14723_), .A2(new_n3303_), .ZN(new_n14731_));
  NAND2_X1   g12295(.A1(new_n14731_), .A2(new_n2436_), .ZN(new_n14732_));
  NOR3_X1    g12296(.A1(new_n14718_), .A2(new_n14717_), .A3(new_n5422_), .ZN(new_n14733_));
  NOR2_X1    g12297(.A1(new_n14733_), .A2(new_n3303_), .ZN(new_n14734_));
  NAND2_X1   g12298(.A1(new_n14703_), .A2(new_n5422_), .ZN(new_n14735_));
  AOI21_X1   g12299(.A1(new_n14735_), .A2(new_n14734_), .B(new_n14732_), .ZN(new_n14736_));
  OAI21_X1   g12300(.A1(new_n14736_), .A2(new_n14730_), .B(pi0299), .ZN(new_n14737_));
  NAND3_X1   g12301(.A1(new_n14727_), .A2(new_n14737_), .A3(pi0039), .ZN(new_n14738_));
  AOI21_X1   g12302(.A1(new_n14738_), .A2(new_n14674_), .B(pi0038), .ZN(new_n14739_));
  NOR2_X1    g12303(.A1(new_n14739_), .A2(new_n14647_), .ZN(new_n14740_));
  OAI21_X1   g12304(.A1(new_n14740_), .A2(new_n14521_), .B(new_n14641_), .ZN(new_n14741_));
  NAND3_X1   g12305(.A1(new_n14741_), .A2(new_n13560_), .A3(new_n14640_), .ZN(new_n14742_));
  AOI21_X1   g12306(.A1(new_n14604_), .A2(new_n14520_), .B(new_n12841_), .ZN(new_n14743_));
  OAI21_X1   g12307(.A1(new_n14739_), .A2(new_n14647_), .B(new_n14524_), .ZN(new_n14744_));
  AOI21_X1   g12308(.A1(new_n14744_), .A2(new_n14743_), .B(new_n13560_), .ZN(new_n14745_));
  AOI21_X1   g12309(.A1(new_n14745_), .A2(new_n14522_), .B(new_n12758_), .ZN(new_n14746_));
  NOR2_X1    g12310(.A1(new_n14740_), .A2(new_n14464_), .ZN(new_n14747_));
  NOR2_X1    g12311(.A1(new_n14747_), .A2(pi0778), .ZN(new_n14748_));
  AOI21_X1   g12312(.A1(new_n14746_), .A2(new_n14742_), .B(new_n14748_), .ZN(new_n14749_));
  NOR2_X1    g12313(.A1(new_n14749_), .A2(pi0785), .ZN(new_n14750_));
  INV_X1     g12314(.I(new_n14750_), .ZN(new_n14751_));
  NAND2_X1   g12315(.A1(new_n14610_), .A2(pi0660), .ZN(new_n14752_));
  NOR2_X1    g12316(.A1(new_n14527_), .A2(pi0609), .ZN(new_n14753_));
  NOR2_X1    g12317(.A1(new_n14753_), .A2(new_n12770_), .ZN(new_n14754_));
  NAND2_X1   g12318(.A1(new_n14749_), .A2(pi0609), .ZN(new_n14755_));
  AOI21_X1   g12319(.A1(new_n14755_), .A2(new_n14754_), .B(new_n14752_), .ZN(new_n14756_));
  OAI21_X1   g12320(.A1(new_n14611_), .A2(new_n12770_), .B(new_n13829_), .ZN(new_n14757_));
  OAI21_X1   g12321(.A1(new_n14527_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n14758_));
  AOI21_X1   g12322(.A1(new_n14749_), .A2(new_n12766_), .B(new_n14758_), .ZN(new_n14759_));
  OAI21_X1   g12323(.A1(new_n14759_), .A2(new_n14757_), .B(pi0785), .ZN(new_n14760_));
  OAI21_X1   g12324(.A1(new_n14760_), .A2(new_n14756_), .B(new_n14751_), .ZN(new_n14761_));
  INV_X1     g12325(.I(new_n14761_), .ZN(new_n14762_));
  NOR2_X1    g12326(.A1(new_n14762_), .A2(pi0781), .ZN(new_n14763_));
  AOI21_X1   g12327(.A1(new_n14617_), .A2(new_n12785_), .B(new_n12880_), .ZN(new_n14764_));
  AOI21_X1   g12328(.A1(new_n14529_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n14765_));
  OAI21_X1   g12329(.A1(new_n14761_), .A2(new_n12781_), .B(new_n14765_), .ZN(new_n14766_));
  NAND2_X1   g12330(.A1(new_n14766_), .A2(new_n14764_), .ZN(new_n14767_));
  AOI21_X1   g12331(.A1(new_n14620_), .A2(pi1154), .B(pi0627), .ZN(new_n14768_));
  AOI21_X1   g12332(.A1(new_n14529_), .A2(pi0618), .B(pi1154), .ZN(new_n14769_));
  OAI21_X1   g12333(.A1(new_n14761_), .A2(pi0618), .B(new_n14769_), .ZN(new_n14770_));
  AOI21_X1   g12334(.A1(new_n14770_), .A2(new_n14768_), .B(new_n12779_), .ZN(new_n14771_));
  AOI21_X1   g12335(.A1(new_n14771_), .A2(new_n14767_), .B(new_n14763_), .ZN(new_n14772_));
  OR2_X2     g12336(.A1(new_n14772_), .A2(pi0789), .Z(new_n14773_));
  OAI21_X1   g12337(.A1(new_n14624_), .A2(pi1159), .B(pi0648), .ZN(new_n14774_));
  INV_X1     g12338(.I(new_n14531_), .ZN(new_n14775_));
  AOI21_X1   g12339(.A1(new_n14775_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n14776_));
  NAND2_X1   g12340(.A1(new_n14772_), .A2(pi0619), .ZN(new_n14777_));
  AOI21_X1   g12341(.A1(new_n14777_), .A2(new_n14776_), .B(new_n14774_), .ZN(new_n14778_));
  OAI21_X1   g12342(.A1(new_n14627_), .A2(new_n12791_), .B(new_n12895_), .ZN(new_n14779_));
  AOI21_X1   g12343(.A1(new_n14775_), .A2(pi0619), .B(pi1159), .ZN(new_n14780_));
  INV_X1     g12344(.I(new_n14780_), .ZN(new_n14781_));
  AOI21_X1   g12345(.A1(new_n14772_), .A2(new_n12793_), .B(new_n14781_), .ZN(new_n14782_));
  OAI21_X1   g12346(.A1(new_n14782_), .A2(new_n14779_), .B(pi0789), .ZN(new_n14783_));
  OAI21_X1   g12347(.A1(new_n14783_), .A2(new_n14778_), .B(new_n14773_), .ZN(new_n14784_));
  NOR2_X1    g12348(.A1(new_n14533_), .A2(pi0626), .ZN(new_n14785_));
  NOR2_X1    g12349(.A1(new_n14785_), .A2(new_n12814_), .ZN(new_n14786_));
  NAND2_X1   g12350(.A1(new_n14784_), .A2(pi0626), .ZN(new_n14787_));
  AOI22_X1   g12351(.A1(new_n14787_), .A2(new_n14786_), .B1(new_n13557_), .B2(new_n14632_), .ZN(new_n14788_));
  OAI21_X1   g12352(.A1(new_n14635_), .A2(new_n12814_), .B(new_n12745_), .ZN(new_n14789_));
  OAI21_X1   g12353(.A1(new_n14533_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n14790_));
  AOI21_X1   g12354(.A1(new_n14784_), .A2(new_n12747_), .B(new_n14790_), .ZN(new_n14791_));
  OAI21_X1   g12355(.A1(new_n14791_), .A2(new_n14789_), .B(pi0788), .ZN(new_n14792_));
  OAI22_X1   g12356(.A1(new_n14788_), .A2(new_n14792_), .B1(pi0788), .B2(new_n14784_), .ZN(new_n14793_));
  NAND2_X1   g12357(.A1(new_n14793_), .A2(pi0628), .ZN(new_n14794_));
  AOI21_X1   g12358(.A1(new_n14794_), .A2(new_n14639_), .B(new_n14540_), .ZN(new_n14795_));
  NOR2_X1    g12359(.A1(new_n14462_), .A2(pi0628), .ZN(new_n14796_));
  AOI21_X1   g12360(.A1(new_n14536_), .A2(pi0628), .B(new_n14796_), .ZN(new_n14797_));
  OAI21_X1   g12361(.A1(new_n14797_), .A2(new_n12742_), .B(new_n12919_), .ZN(new_n14798_));
  OAI21_X1   g12362(.A1(new_n14637_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n14799_));
  AOI21_X1   g12363(.A1(new_n14793_), .A2(new_n12920_), .B(new_n14799_), .ZN(new_n14800_));
  OAI21_X1   g12364(.A1(new_n14800_), .A2(new_n14798_), .B(pi0792), .ZN(new_n14801_));
  OR2_X2     g12365(.A1(new_n14793_), .A2(pi0792), .Z(new_n14802_));
  OAI21_X1   g12366(.A1(new_n14801_), .A2(new_n14795_), .B(new_n14802_), .ZN(new_n14803_));
  AND2_X2    g12367(.A1(new_n14803_), .A2(new_n12972_), .Z(new_n14804_));
  OAI21_X1   g12368(.A1(new_n14797_), .A2(new_n12742_), .B(pi0792), .ZN(new_n14805_));
  NOR2_X1    g12369(.A1(new_n14805_), .A2(new_n14539_), .ZN(new_n14806_));
  NOR2_X1    g12370(.A1(new_n14536_), .A2(pi0792), .ZN(new_n14807_));
  NOR2_X1    g12371(.A1(new_n14806_), .A2(new_n14807_), .ZN(new_n14808_));
  NAND2_X1   g12372(.A1(new_n14808_), .A2(new_n12741_), .ZN(new_n14809_));
  NAND2_X1   g12373(.A1(new_n14463_), .A2(pi0647), .ZN(new_n14810_));
  AOI21_X1   g12374(.A1(new_n14809_), .A2(new_n14810_), .B(pi1157), .ZN(new_n14811_));
  INV_X1     g12375(.I(new_n14811_), .ZN(new_n14812_));
  NOR2_X1    g12376(.A1(new_n14462_), .A2(new_n13384_), .ZN(new_n14813_));
  AOI21_X1   g12377(.A1(new_n14637_), .A2(new_n13384_), .B(new_n14813_), .ZN(new_n14814_));
  AOI21_X1   g12378(.A1(new_n14814_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n14815_));
  OAI21_X1   g12379(.A1(new_n14803_), .A2(new_n12741_), .B(new_n14815_), .ZN(new_n14816_));
  NAND3_X1   g12380(.A1(new_n14816_), .A2(pi0630), .A3(new_n14812_), .ZN(new_n14817_));
  NOR2_X1    g12381(.A1(new_n14462_), .A2(pi0647), .ZN(new_n14818_));
  AOI21_X1   g12382(.A1(new_n14808_), .A2(pi0647), .B(new_n14818_), .ZN(new_n14819_));
  NOR2_X1    g12383(.A1(new_n14819_), .A2(new_n12965_), .ZN(new_n14820_));
  NOR2_X1    g12384(.A1(new_n14820_), .A2(pi0630), .ZN(new_n14821_));
  AOI21_X1   g12385(.A1(new_n14814_), .A2(pi0647), .B(pi1157), .ZN(new_n14822_));
  OAI21_X1   g12386(.A1(new_n14803_), .A2(pi0647), .B(new_n14822_), .ZN(new_n14823_));
  AOI21_X1   g12387(.A1(new_n14823_), .A2(new_n14821_), .B(new_n12972_), .ZN(new_n14824_));
  AOI21_X1   g12388(.A1(new_n14824_), .A2(new_n14817_), .B(new_n14804_), .ZN(new_n14825_));
  OAI21_X1   g12389(.A1(new_n14825_), .A2(pi0790), .B(new_n5477_), .ZN(new_n14826_));
  NOR2_X1    g12390(.A1(new_n14463_), .A2(new_n12985_), .ZN(new_n14827_));
  AOI21_X1   g12391(.A1(new_n14814_), .A2(new_n12985_), .B(new_n14827_), .ZN(new_n14828_));
  NOR2_X1    g12392(.A1(new_n14462_), .A2(new_n12975_), .ZN(new_n14829_));
  AOI21_X1   g12393(.A1(new_n14828_), .A2(new_n12975_), .B(new_n14829_), .ZN(new_n14830_));
  OAI21_X1   g12394(.A1(new_n14830_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n14831_));
  INV_X1     g12395(.I(new_n14808_), .ZN(new_n14832_));
  NOR2_X1    g12396(.A1(new_n14820_), .A2(new_n12972_), .ZN(new_n14833_));
  AOI22_X1   g12397(.A1(new_n14833_), .A2(new_n14812_), .B1(new_n12972_), .B2(new_n14832_), .ZN(new_n14834_));
  NOR2_X1    g12398(.A1(new_n14834_), .A2(new_n12975_), .ZN(new_n14835_));
  NOR2_X1    g12399(.A1(new_n14835_), .A2(pi0715), .ZN(new_n14836_));
  NAND2_X1   g12400(.A1(new_n14825_), .A2(new_n12975_), .ZN(new_n14837_));
  AOI21_X1   g12401(.A1(new_n14837_), .A2(new_n14836_), .B(new_n14831_), .ZN(new_n14838_));
  NOR2_X1    g12402(.A1(new_n14462_), .A2(pi0644), .ZN(new_n14839_));
  AOI21_X1   g12403(.A1(new_n14828_), .A2(pi0644), .B(new_n14839_), .ZN(new_n14840_));
  OAI21_X1   g12404(.A1(new_n14840_), .A2(pi0715), .B(pi1160), .ZN(new_n14841_));
  OAI21_X1   g12405(.A1(new_n14834_), .A2(pi0644), .B(pi0715), .ZN(new_n14842_));
  AOI21_X1   g12406(.A1(new_n14825_), .A2(pi0644), .B(new_n14842_), .ZN(new_n14843_));
  OAI21_X1   g12407(.A1(new_n14843_), .A2(new_n14841_), .B(pi0790), .ZN(new_n14844_));
  NOR2_X1    g12408(.A1(new_n14844_), .A2(new_n14838_), .ZN(new_n14845_));
  AOI21_X1   g12409(.A1(new_n6165_), .A2(new_n2724_), .B(pi0057), .ZN(new_n14846_));
  OAI21_X1   g12410(.A1(new_n14845_), .A2(new_n14826_), .B(new_n14846_), .ZN(new_n14847_));
  AOI21_X1   g12411(.A1(new_n14847_), .A2(new_n14445_), .B(new_n14444_), .ZN(po0299));
  NOR2_X1    g12412(.A1(new_n3042_), .A2(pi0143), .ZN(new_n14849_));
  INV_X1     g12413(.I(new_n14849_), .ZN(new_n14850_));
  INV_X1     g12414(.I(pi0774), .ZN(new_n14851_));
  AOI21_X1   g12415(.A1(new_n12756_), .A2(new_n14851_), .B(new_n14849_), .ZN(new_n14852_));
  NOR3_X1    g12416(.A1(new_n14852_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n14853_));
  NOR2_X1    g12417(.A1(new_n14852_), .A2(new_n12762_), .ZN(new_n14854_));
  AOI21_X1   g12418(.A1(new_n14854_), .A2(new_n12768_), .B(pi1155), .ZN(new_n14855_));
  INV_X1     g12419(.I(new_n14852_), .ZN(new_n14856_));
  AOI21_X1   g12420(.A1(new_n14856_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n14857_));
  NOR3_X1    g12421(.A1(new_n14855_), .A2(new_n14857_), .A3(new_n12764_), .ZN(new_n14858_));
  NOR2_X1    g12422(.A1(new_n14858_), .A2(new_n14853_), .ZN(new_n14859_));
  NOR2_X1    g12423(.A1(new_n14859_), .A2(pi0781), .ZN(new_n14860_));
  INV_X1     g12424(.I(new_n14859_), .ZN(new_n14861_));
  AOI21_X1   g12425(.A1(new_n14861_), .A2(new_n12783_), .B(pi1154), .ZN(new_n14862_));
  AOI21_X1   g12426(.A1(new_n14861_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n14863_));
  NOR3_X1    g12427(.A1(new_n14862_), .A2(new_n14863_), .A3(new_n12779_), .ZN(new_n14864_));
  NOR2_X1    g12428(.A1(new_n14864_), .A2(new_n14860_), .ZN(new_n14865_));
  NOR3_X1    g12429(.A1(new_n14864_), .A2(pi0619), .A3(new_n14860_), .ZN(new_n14866_));
  NOR2_X1    g12430(.A1(new_n14849_), .A2(new_n12793_), .ZN(new_n14867_));
  OAI21_X1   g12431(.A1(new_n14866_), .A2(new_n14867_), .B(new_n12791_), .ZN(new_n14868_));
  NAND2_X1   g12432(.A1(new_n14865_), .A2(pi0619), .ZN(new_n14869_));
  NAND2_X1   g12433(.A1(new_n14850_), .A2(new_n12793_), .ZN(new_n14870_));
  AOI21_X1   g12434(.A1(new_n14869_), .A2(new_n14870_), .B(new_n12791_), .ZN(new_n14871_));
  NOR2_X1    g12435(.A1(new_n14871_), .A2(new_n12796_), .ZN(new_n14872_));
  NAND2_X1   g12436(.A1(new_n14872_), .A2(new_n14868_), .ZN(new_n14873_));
  OAI21_X1   g12437(.A1(pi0789), .A2(new_n14865_), .B(new_n14873_), .ZN(new_n14874_));
  NAND2_X1   g12438(.A1(new_n14874_), .A2(new_n12804_), .ZN(new_n14875_));
  OAI21_X1   g12439(.A1(new_n12749_), .A2(new_n14850_), .B(new_n14875_), .ZN(new_n14876_));
  NAND2_X1   g12440(.A1(new_n14876_), .A2(pi0788), .ZN(new_n14877_));
  NAND2_X1   g12441(.A1(new_n14874_), .A2(new_n12808_), .ZN(new_n14878_));
  NAND2_X1   g12442(.A1(new_n14877_), .A2(new_n14878_), .ZN(new_n14879_));
  NOR2_X1    g12443(.A1(new_n14879_), .A2(pi0628), .ZN(new_n14880_));
  AOI21_X1   g12444(.A1(new_n12826_), .A2(pi0687), .B(new_n14849_), .ZN(new_n14881_));
  NOR2_X1    g12445(.A1(new_n14881_), .A2(new_n12754_), .ZN(new_n14882_));
  NOR2_X1    g12446(.A1(new_n14882_), .A2(new_n14856_), .ZN(new_n14883_));
  NAND2_X1   g12447(.A1(new_n14883_), .A2(new_n12758_), .ZN(new_n14884_));
  INV_X1     g12448(.I(pi0687), .ZN(new_n14885_));
  NOR2_X1    g12449(.A1(new_n12834_), .A2(new_n14885_), .ZN(new_n14886_));
  INV_X1     g12450(.I(new_n14886_), .ZN(new_n14887_));
  NOR2_X1    g12451(.A1(new_n14849_), .A2(pi1153), .ZN(new_n14888_));
  NAND2_X1   g12452(.A1(new_n14887_), .A2(new_n14888_), .ZN(new_n14889_));
  NAND2_X1   g12453(.A1(new_n14882_), .A2(pi0625), .ZN(new_n14890_));
  NAND3_X1   g12454(.A1(new_n14890_), .A2(pi1153), .A3(new_n14852_), .ZN(new_n14891_));
  AND3_X2    g12455(.A1(new_n14889_), .A2(pi0608), .A3(new_n14891_), .Z(new_n14892_));
  NOR2_X1    g12456(.A1(new_n14886_), .A2(new_n14881_), .ZN(new_n14893_));
  NOR2_X1    g12457(.A1(new_n14893_), .A2(new_n12841_), .ZN(new_n14894_));
  NOR2_X1    g12458(.A1(new_n14894_), .A2(pi0608), .ZN(new_n14895_));
  INV_X1     g12459(.I(new_n14890_), .ZN(new_n14896_));
  OAI21_X1   g12460(.A1(new_n14896_), .A2(new_n14883_), .B(new_n14888_), .ZN(new_n14897_));
  NAND2_X1   g12461(.A1(new_n14895_), .A2(new_n14897_), .ZN(new_n14898_));
  NAND2_X1   g12462(.A1(new_n14898_), .A2(pi0778), .ZN(new_n14899_));
  OAI21_X1   g12463(.A1(new_n14899_), .A2(new_n14892_), .B(new_n14884_), .ZN(new_n14900_));
  INV_X1     g12464(.I(new_n14900_), .ZN(new_n14901_));
  NOR2_X1    g12465(.A1(new_n14881_), .A2(pi0778), .ZN(new_n14902_));
  INV_X1     g12466(.I(new_n14889_), .ZN(new_n14903_));
  NOR3_X1    g12467(.A1(new_n14903_), .A2(new_n12758_), .A3(new_n14894_), .ZN(new_n14904_));
  NOR2_X1    g12468(.A1(new_n14904_), .A2(new_n14902_), .ZN(new_n14905_));
  INV_X1     g12469(.I(new_n14905_), .ZN(new_n14906_));
  NOR2_X1    g12470(.A1(new_n14906_), .A2(pi0609), .ZN(new_n14907_));
  AOI21_X1   g12471(.A1(new_n14900_), .A2(pi0609), .B(new_n14907_), .ZN(new_n14908_));
  NOR2_X1    g12472(.A1(new_n14908_), .A2(new_n12770_), .ZN(new_n14909_));
  NOR2_X1    g12473(.A1(new_n14909_), .A2(new_n14855_), .ZN(new_n14910_));
  NOR2_X1    g12474(.A1(new_n14901_), .A2(pi0609), .ZN(new_n14911_));
  NOR2_X1    g12475(.A1(new_n14906_), .A2(new_n12766_), .ZN(new_n14912_));
  OAI21_X1   g12476(.A1(new_n14911_), .A2(new_n14912_), .B(new_n12770_), .ZN(new_n14913_));
  NOR2_X1    g12477(.A1(new_n14857_), .A2(pi0660), .ZN(new_n14914_));
  AOI22_X1   g12478(.A1(new_n14910_), .A2(pi0660), .B1(new_n14913_), .B2(new_n14914_), .ZN(new_n14915_));
  NAND2_X1   g12479(.A1(new_n14915_), .A2(pi0785), .ZN(new_n14916_));
  OAI21_X1   g12480(.A1(pi0785), .A2(new_n14901_), .B(new_n14916_), .ZN(new_n14917_));
  INV_X1     g12481(.I(new_n14863_), .ZN(new_n14918_));
  NOR2_X1    g12482(.A1(new_n14905_), .A2(new_n12871_), .ZN(new_n14919_));
  NOR2_X1    g12483(.A1(new_n14919_), .A2(new_n12781_), .ZN(new_n14920_));
  AOI21_X1   g12484(.A1(new_n14917_), .A2(new_n12781_), .B(new_n14920_), .ZN(new_n14921_));
  OAI21_X1   g12485(.A1(new_n14921_), .A2(pi1154), .B(new_n14918_), .ZN(new_n14922_));
  INV_X1     g12486(.I(new_n14919_), .ZN(new_n14923_));
  NAND2_X1   g12487(.A1(new_n14923_), .A2(new_n12781_), .ZN(new_n14924_));
  NAND2_X1   g12488(.A1(new_n14917_), .A2(pi0618), .ZN(new_n14925_));
  AOI21_X1   g12489(.A1(new_n14925_), .A2(new_n14924_), .B(new_n12785_), .ZN(new_n14926_));
  OR2_X2     g12490(.A1(new_n14862_), .A2(new_n12880_), .Z(new_n14927_));
  OAI22_X1   g12491(.A1(new_n14922_), .A2(pi0627), .B1(new_n14926_), .B2(new_n14927_), .ZN(new_n14928_));
  NOR2_X1    g12492(.A1(new_n14928_), .A2(new_n12779_), .ZN(new_n14929_));
  AOI21_X1   g12493(.A1(new_n12779_), .A2(new_n14917_), .B(new_n14929_), .ZN(new_n14930_));
  OAI21_X1   g12494(.A1(new_n14930_), .A2(pi0789), .B(new_n12819_), .ZN(new_n14931_));
  NOR2_X1    g12495(.A1(new_n14923_), .A2(new_n12889_), .ZN(new_n14932_));
  NOR2_X1    g12496(.A1(new_n14932_), .A2(pi0619), .ZN(new_n14933_));
  NOR2_X1    g12497(.A1(new_n14930_), .A2(new_n12793_), .ZN(new_n14934_));
  OAI21_X1   g12498(.A1(new_n14934_), .A2(new_n14933_), .B(pi1159), .ZN(new_n14935_));
  NAND3_X1   g12499(.A1(new_n14935_), .A2(pi0648), .A3(new_n14868_), .ZN(new_n14936_));
  INV_X1     g12500(.I(new_n14932_), .ZN(new_n14937_));
  NAND2_X1   g12501(.A1(new_n14937_), .A2(pi0619), .ZN(new_n14938_));
  OAI21_X1   g12502(.A1(new_n14930_), .A2(pi0619), .B(new_n14938_), .ZN(new_n14939_));
  AOI21_X1   g12503(.A1(new_n14939_), .A2(new_n12791_), .B(new_n14871_), .ZN(new_n14940_));
  AOI21_X1   g12504(.A1(new_n14940_), .A2(new_n12895_), .B(new_n12796_), .ZN(new_n14941_));
  AOI21_X1   g12505(.A1(new_n14941_), .A2(new_n14936_), .B(new_n14931_), .ZN(new_n14942_));
  AOI22_X1   g12506(.A1(new_n14876_), .A2(new_n12914_), .B1(new_n12913_), .B2(new_n14932_), .ZN(new_n14943_));
  NOR2_X1    g12507(.A1(new_n14943_), .A2(new_n12808_), .ZN(new_n14944_));
  NOR2_X1    g12508(.A1(new_n14942_), .A2(new_n14944_), .ZN(new_n14945_));
  AOI21_X1   g12509(.A1(new_n14945_), .A2(pi0628), .B(new_n14880_), .ZN(new_n14946_));
  NOR2_X1    g12510(.A1(new_n14937_), .A2(new_n12924_), .ZN(new_n14947_));
  NAND2_X1   g12511(.A1(new_n14947_), .A2(new_n12922_), .ZN(new_n14948_));
  AOI21_X1   g12512(.A1(new_n14948_), .A2(new_n12742_), .B(new_n12919_), .ZN(new_n14949_));
  OAI21_X1   g12513(.A1(new_n14946_), .A2(new_n12742_), .B(new_n14949_), .ZN(new_n14950_));
  NOR2_X1    g12514(.A1(new_n14879_), .A2(new_n12920_), .ZN(new_n14951_));
  AOI21_X1   g12515(.A1(new_n14945_), .A2(new_n12920_), .B(new_n14951_), .ZN(new_n14952_));
  NAND2_X1   g12516(.A1(new_n14947_), .A2(new_n12932_), .ZN(new_n14953_));
  AOI21_X1   g12517(.A1(new_n14953_), .A2(pi1156), .B(pi0629), .ZN(new_n14954_));
  OAI21_X1   g12518(.A1(new_n14952_), .A2(pi1156), .B(new_n14954_), .ZN(new_n14955_));
  NAND3_X1   g12519(.A1(new_n14950_), .A2(new_n14955_), .A3(pi0792), .ZN(new_n14956_));
  NAND2_X1   g12520(.A1(new_n14945_), .A2(new_n12937_), .ZN(new_n14957_));
  AOI21_X1   g12521(.A1(new_n14956_), .A2(new_n14957_), .B(new_n12741_), .ZN(new_n14958_));
  NOR2_X1    g12522(.A1(new_n14879_), .A2(new_n12943_), .ZN(new_n14959_));
  AOI21_X1   g12523(.A1(new_n12943_), .A2(new_n14850_), .B(new_n14959_), .ZN(new_n14960_));
  NOR2_X1    g12524(.A1(new_n14960_), .A2(pi0647), .ZN(new_n14961_));
  OAI21_X1   g12525(.A1(new_n14958_), .A2(new_n14961_), .B(pi1157), .ZN(new_n14962_));
  NAND2_X1   g12526(.A1(new_n14947_), .A2(new_n12954_), .ZN(new_n14963_));
  NAND2_X1   g12527(.A1(new_n14963_), .A2(new_n12741_), .ZN(new_n14964_));
  NOR2_X1    g12528(.A1(new_n14849_), .A2(new_n12741_), .ZN(new_n14965_));
  INV_X1     g12529(.I(new_n14965_), .ZN(new_n14966_));
  AOI21_X1   g12530(.A1(new_n14964_), .A2(new_n14966_), .B(pi1157), .ZN(new_n14967_));
  INV_X1     g12531(.I(new_n14967_), .ZN(new_n14968_));
  NAND3_X1   g12532(.A1(new_n14962_), .A2(pi0630), .A3(new_n14968_), .ZN(new_n14969_));
  NAND2_X1   g12533(.A1(new_n14956_), .A2(new_n14957_), .ZN(new_n14970_));
  NOR2_X1    g12534(.A1(new_n14960_), .A2(new_n12741_), .ZN(new_n14971_));
  AOI21_X1   g12535(.A1(new_n14970_), .A2(new_n12741_), .B(new_n14971_), .ZN(new_n14972_));
  NAND2_X1   g12536(.A1(new_n14963_), .A2(pi0647), .ZN(new_n14973_));
  NAND2_X1   g12537(.A1(new_n14850_), .A2(new_n12741_), .ZN(new_n14974_));
  AOI21_X1   g12538(.A1(new_n14973_), .A2(new_n14974_), .B(new_n12965_), .ZN(new_n14975_));
  NOR2_X1    g12539(.A1(new_n14975_), .A2(pi0630), .ZN(new_n14976_));
  OAI21_X1   g12540(.A1(new_n14972_), .A2(pi1157), .B(new_n14976_), .ZN(new_n14977_));
  NAND3_X1   g12541(.A1(new_n14969_), .A2(new_n14977_), .A3(pi0787), .ZN(new_n14978_));
  NAND2_X1   g12542(.A1(new_n14970_), .A2(new_n12972_), .ZN(new_n14979_));
  AOI21_X1   g12543(.A1(new_n14978_), .A2(new_n14979_), .B(pi0644), .ZN(new_n14980_));
  OR2_X2     g12544(.A1(new_n14975_), .A2(new_n12972_), .Z(new_n14981_));
  OAI22_X1   g12545(.A1(new_n14981_), .A2(new_n14967_), .B1(pi0787), .B2(new_n14963_), .ZN(new_n14982_));
  NOR2_X1    g12546(.A1(new_n14982_), .A2(new_n12975_), .ZN(new_n14983_));
  OAI21_X1   g12547(.A1(new_n14980_), .A2(new_n14983_), .B(new_n12740_), .ZN(new_n14984_));
  NAND2_X1   g12548(.A1(new_n14960_), .A2(new_n12985_), .ZN(new_n14985_));
  OAI21_X1   g12549(.A1(new_n12985_), .A2(new_n14850_), .B(new_n14985_), .ZN(new_n14986_));
  NOR2_X1    g12550(.A1(new_n14986_), .A2(pi0644), .ZN(new_n14987_));
  NOR2_X1    g12551(.A1(new_n14849_), .A2(new_n12975_), .ZN(new_n14988_));
  OAI21_X1   g12552(.A1(new_n14987_), .A2(new_n14988_), .B(pi0715), .ZN(new_n14989_));
  NAND3_X1   g12553(.A1(new_n14984_), .A2(new_n12739_), .A3(new_n14989_), .ZN(new_n14990_));
  NAND2_X1   g12554(.A1(new_n14978_), .A2(new_n14979_), .ZN(new_n14991_));
  NOR2_X1    g12555(.A1(new_n14982_), .A2(pi0644), .ZN(new_n14992_));
  AOI21_X1   g12556(.A1(new_n14991_), .A2(pi0644), .B(new_n14992_), .ZN(new_n14993_));
  NAND2_X1   g12557(.A1(new_n14850_), .A2(new_n12975_), .ZN(new_n14994_));
  OAI21_X1   g12558(.A1(new_n14986_), .A2(new_n12975_), .B(new_n14994_), .ZN(new_n14995_));
  AOI21_X1   g12559(.A1(new_n14995_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n14996_));
  OAI21_X1   g12560(.A1(new_n14993_), .A2(new_n12740_), .B(new_n14996_), .ZN(new_n14997_));
  NAND3_X1   g12561(.A1(new_n14990_), .A2(new_n14997_), .A3(pi0790), .ZN(new_n14998_));
  NAND2_X1   g12562(.A1(new_n14991_), .A2(new_n13000_), .ZN(new_n14999_));
  AOI21_X1   g12563(.A1(new_n14998_), .A2(new_n14999_), .B(new_n12738_), .ZN(new_n15000_));
  AOI21_X1   g12564(.A1(po1038), .A2(new_n10695_), .B(pi0832), .ZN(new_n15001_));
  NOR2_X1    g12565(.A1(new_n13193_), .A2(pi0143), .ZN(new_n15002_));
  AOI21_X1   g12566(.A1(new_n15002_), .A2(pi0644), .B(new_n12740_), .ZN(new_n15003_));
  NOR2_X1    g12567(.A1(new_n2609_), .A2(new_n10695_), .ZN(new_n15004_));
  INV_X1     g12568(.I(new_n15004_), .ZN(new_n15005_));
  NOR2_X1    g12569(.A1(new_n5346_), .A2(new_n13340_), .ZN(new_n15006_));
  INV_X1     g12570(.I(new_n15006_), .ZN(new_n15007_));
  NOR2_X1    g12571(.A1(new_n15007_), .A2(new_n3265_), .ZN(new_n15008_));
  NAND2_X1   g12572(.A1(new_n13245_), .A2(new_n3265_), .ZN(new_n15009_));
  NAND2_X1   g12573(.A1(new_n15009_), .A2(pi0143), .ZN(new_n15010_));
  AOI21_X1   g12574(.A1(new_n5336_), .A2(new_n13275_), .B(new_n3265_), .ZN(new_n15011_));
  AOI21_X1   g12575(.A1(new_n13333_), .A2(new_n13257_), .B(pi0038), .ZN(new_n15012_));
  NOR2_X1    g12576(.A1(new_n15012_), .A2(new_n15011_), .ZN(new_n15013_));
  NOR2_X1    g12577(.A1(pi0143), .A2(pi0774), .ZN(new_n15014_));
  NAND2_X1   g12578(.A1(new_n15013_), .A2(new_n15014_), .ZN(new_n15015_));
  AOI21_X1   g12579(.A1(new_n15015_), .A2(new_n15010_), .B(new_n15008_), .ZN(new_n15016_));
  AOI21_X1   g12580(.A1(new_n13395_), .A2(new_n10695_), .B(new_n14851_), .ZN(new_n15017_));
  OAI21_X1   g12581(.A1(new_n15016_), .A2(new_n15017_), .B(new_n2609_), .ZN(new_n15018_));
  AOI21_X1   g12582(.A1(new_n15018_), .A2(new_n15005_), .B(new_n12760_), .ZN(new_n15019_));
  NOR2_X1    g12583(.A1(new_n15002_), .A2(new_n12761_), .ZN(new_n15020_));
  NOR2_X1    g12584(.A1(new_n15019_), .A2(new_n15020_), .ZN(new_n15021_));
  NAND2_X1   g12585(.A1(new_n15019_), .A2(new_n12766_), .ZN(new_n15022_));
  OAI21_X1   g12586(.A1(new_n13353_), .A2(new_n15002_), .B(new_n15022_), .ZN(new_n15023_));
  NAND2_X1   g12587(.A1(new_n15023_), .A2(new_n12770_), .ZN(new_n15024_));
  INV_X1     g12588(.I(new_n15002_), .ZN(new_n15025_));
  AOI22_X1   g12589(.A1(new_n15019_), .A2(pi0609), .B1(new_n13357_), .B2(new_n15025_), .ZN(new_n15026_));
  NOR2_X1    g12590(.A1(new_n15026_), .A2(new_n12770_), .ZN(new_n15027_));
  NOR2_X1    g12591(.A1(new_n15027_), .A2(new_n12764_), .ZN(new_n15028_));
  AOI22_X1   g12592(.A1(new_n15028_), .A2(new_n15024_), .B1(new_n12764_), .B2(new_n15021_), .ZN(new_n15029_));
  NOR2_X1    g12593(.A1(new_n15002_), .A2(new_n12781_), .ZN(new_n15030_));
  AOI21_X1   g12594(.A1(new_n15029_), .A2(new_n12781_), .B(new_n15030_), .ZN(new_n15031_));
  NOR2_X1    g12595(.A1(new_n15031_), .A2(pi1154), .ZN(new_n15032_));
  NOR2_X1    g12596(.A1(new_n15002_), .A2(pi0618), .ZN(new_n15033_));
  AOI21_X1   g12597(.A1(new_n15029_), .A2(pi0618), .B(new_n15033_), .ZN(new_n15034_));
  OAI21_X1   g12598(.A1(new_n15034_), .A2(new_n12785_), .B(pi0781), .ZN(new_n15035_));
  OAI22_X1   g12599(.A1(new_n15035_), .A2(new_n15032_), .B1(pi0781), .B2(new_n15029_), .ZN(new_n15036_));
  NAND2_X1   g12600(.A1(new_n15025_), .A2(pi0619), .ZN(new_n15037_));
  OAI21_X1   g12601(.A1(new_n15036_), .A2(pi0619), .B(new_n15037_), .ZN(new_n15038_));
  NAND2_X1   g12602(.A1(new_n15038_), .A2(new_n12791_), .ZN(new_n15039_));
  NAND2_X1   g12603(.A1(new_n15025_), .A2(new_n12793_), .ZN(new_n15040_));
  OAI21_X1   g12604(.A1(new_n15036_), .A2(new_n12793_), .B(new_n15040_), .ZN(new_n15041_));
  AOI21_X1   g12605(.A1(new_n15041_), .A2(pi1159), .B(new_n12796_), .ZN(new_n15042_));
  AOI22_X1   g12606(.A1(new_n15042_), .A2(new_n15039_), .B1(new_n12796_), .B2(new_n15036_), .ZN(new_n15043_));
  NOR2_X1    g12607(.A1(new_n15002_), .A2(pi0626), .ZN(new_n15044_));
  AOI21_X1   g12608(.A1(new_n15043_), .A2(pi0626), .B(new_n15044_), .ZN(new_n15045_));
  NOR2_X1    g12609(.A1(new_n15045_), .A2(new_n12745_), .ZN(new_n15046_));
  NOR2_X1    g12610(.A1(new_n15002_), .A2(new_n12747_), .ZN(new_n15047_));
  AOI21_X1   g12611(.A1(new_n15043_), .A2(new_n12747_), .B(new_n15047_), .ZN(new_n15048_));
  OAI21_X1   g12612(.A1(new_n15048_), .A2(pi1158), .B(pi0788), .ZN(new_n15049_));
  OAI22_X1   g12613(.A1(new_n15049_), .A2(new_n15046_), .B1(pi0788), .B2(new_n15043_), .ZN(new_n15050_));
  NOR2_X1    g12614(.A1(new_n15050_), .A2(new_n12943_), .ZN(new_n15051_));
  NOR2_X1    g12615(.A1(new_n15002_), .A2(new_n13384_), .ZN(new_n15052_));
  NOR2_X1    g12616(.A1(new_n15051_), .A2(new_n15052_), .ZN(new_n15053_));
  INV_X1     g12617(.I(new_n15053_), .ZN(new_n15054_));
  NAND2_X1   g12618(.A1(new_n15002_), .A2(new_n12984_), .ZN(new_n15055_));
  OAI21_X1   g12619(.A1(new_n15054_), .A2(new_n12984_), .B(new_n15055_), .ZN(new_n15056_));
  NAND2_X1   g12620(.A1(new_n15056_), .A2(new_n12975_), .ZN(new_n15057_));
  AOI21_X1   g12621(.A1(new_n15057_), .A2(new_n15003_), .B(pi1160), .ZN(new_n15058_));
  NOR2_X1    g12622(.A1(new_n15025_), .A2(new_n12870_), .ZN(new_n15059_));
  AOI21_X1   g12623(.A1(new_n14117_), .A2(new_n14116_), .B(pi0143), .ZN(new_n15060_));
  AOI21_X1   g12624(.A1(new_n14121_), .A2(new_n14120_), .B(new_n10695_), .ZN(new_n15061_));
  OAI21_X1   g12625(.A1(new_n15060_), .A2(new_n15061_), .B(new_n3265_), .ZN(new_n15062_));
  NAND2_X1   g12626(.A1(new_n13397_), .A2(new_n10695_), .ZN(new_n15063_));
  AOI21_X1   g12627(.A1(new_n13399_), .A2(new_n15063_), .B(new_n14885_), .ZN(new_n15064_));
  NAND2_X1   g12628(.A1(new_n15062_), .A2(new_n15064_), .ZN(new_n15065_));
  NAND3_X1   g12629(.A1(new_n13395_), .A2(new_n10695_), .A3(new_n14885_), .ZN(new_n15066_));
  NAND3_X1   g12630(.A1(new_n15065_), .A2(new_n15066_), .A3(new_n2609_), .ZN(new_n15067_));
  NAND2_X1   g12631(.A1(new_n15067_), .A2(new_n15005_), .ZN(new_n15068_));
  NAND2_X1   g12632(.A1(new_n15068_), .A2(new_n13521_), .ZN(new_n15069_));
  NAND2_X1   g12633(.A1(new_n15025_), .A2(pi0625), .ZN(new_n15070_));
  AOI21_X1   g12634(.A1(new_n15069_), .A2(new_n15070_), .B(pi1153), .ZN(new_n15071_));
  AOI21_X1   g12635(.A1(new_n15067_), .A2(new_n15005_), .B(new_n13521_), .ZN(new_n15072_));
  NOR2_X1    g12636(.A1(new_n15002_), .A2(pi0625), .ZN(new_n15073_));
  OAI21_X1   g12637(.A1(new_n15072_), .A2(new_n15073_), .B(pi1153), .ZN(new_n15074_));
  NAND2_X1   g12638(.A1(new_n15074_), .A2(pi0778), .ZN(new_n15075_));
  OAI22_X1   g12639(.A1(new_n15075_), .A2(new_n15071_), .B1(pi0778), .B2(new_n15068_), .ZN(new_n15076_));
  AOI21_X1   g12640(.A1(new_n15076_), .A2(new_n12870_), .B(new_n15059_), .ZN(new_n15077_));
  NOR2_X1    g12641(.A1(new_n15002_), .A2(new_n12888_), .ZN(new_n15078_));
  AOI21_X1   g12642(.A1(new_n15077_), .A2(new_n12888_), .B(new_n15078_), .ZN(new_n15079_));
  NOR2_X1    g12643(.A1(new_n15025_), .A2(new_n12911_), .ZN(new_n15080_));
  AOI21_X1   g12644(.A1(new_n15079_), .A2(new_n12911_), .B(new_n15080_), .ZN(new_n15081_));
  NAND2_X1   g12645(.A1(new_n15081_), .A2(new_n13392_), .ZN(new_n15082_));
  OAI21_X1   g12646(.A1(new_n13392_), .A2(new_n15002_), .B(new_n15082_), .ZN(new_n15083_));
  NAND2_X1   g12647(.A1(new_n15083_), .A2(new_n12920_), .ZN(new_n15084_));
  NAND2_X1   g12648(.A1(new_n15025_), .A2(pi0628), .ZN(new_n15085_));
  AOI21_X1   g12649(.A1(new_n15084_), .A2(new_n15085_), .B(pi1156), .ZN(new_n15086_));
  NAND2_X1   g12650(.A1(new_n15025_), .A2(new_n12920_), .ZN(new_n15087_));
  NAND2_X1   g12651(.A1(new_n15083_), .A2(pi0628), .ZN(new_n15088_));
  AOI21_X1   g12652(.A1(new_n15088_), .A2(new_n15087_), .B(new_n12742_), .ZN(new_n15089_));
  NOR3_X1    g12653(.A1(new_n15086_), .A2(new_n15089_), .A3(new_n12937_), .ZN(new_n15090_));
  NOR2_X1    g12654(.A1(new_n15083_), .A2(pi0792), .ZN(new_n15091_));
  NOR2_X1    g12655(.A1(new_n15090_), .A2(new_n15091_), .ZN(new_n15092_));
  NAND2_X1   g12656(.A1(new_n15092_), .A2(new_n12741_), .ZN(new_n15093_));
  NAND2_X1   g12657(.A1(new_n15025_), .A2(pi0647), .ZN(new_n15094_));
  AOI21_X1   g12658(.A1(new_n15093_), .A2(new_n15094_), .B(pi1157), .ZN(new_n15095_));
  NAND2_X1   g12659(.A1(new_n15092_), .A2(pi0647), .ZN(new_n15096_));
  OAI21_X1   g12660(.A1(pi0647), .A2(new_n15002_), .B(new_n15096_), .ZN(new_n15097_));
  NAND2_X1   g12661(.A1(new_n15097_), .A2(pi1157), .ZN(new_n15098_));
  NAND2_X1   g12662(.A1(new_n15098_), .A2(pi0787), .ZN(new_n15099_));
  OAI22_X1   g12663(.A1(new_n15099_), .A2(new_n15095_), .B1(pi0787), .B2(new_n15092_), .ZN(new_n15100_));
  AOI21_X1   g12664(.A1(new_n15100_), .A2(pi0644), .B(pi0715), .ZN(new_n15101_));
  NOR2_X1    g12665(.A1(new_n15086_), .A2(new_n12919_), .ZN(new_n15102_));
  AOI21_X1   g12666(.A1(new_n15050_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n15103_));
  OAI21_X1   g12667(.A1(new_n15045_), .A2(new_n12745_), .B(new_n13557_), .ZN(new_n15104_));
  AOI21_X1   g12668(.A1(new_n15081_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n15105_));
  NOR3_X1    g12669(.A1(new_n15016_), .A2(new_n15017_), .A3(pi0687), .ZN(new_n15106_));
  OAI21_X1   g12670(.A1(new_n13800_), .A2(pi0039), .B(new_n3265_), .ZN(new_n15107_));
  NOR3_X1    g12671(.A1(new_n13566_), .A2(new_n3265_), .A3(pi0039), .ZN(new_n15108_));
  INV_X1     g12672(.I(new_n15108_), .ZN(new_n15109_));
  NOR2_X1    g12673(.A1(new_n13692_), .A2(new_n2627_), .ZN(new_n15110_));
  AOI21_X1   g12674(.A1(new_n15107_), .A2(new_n15109_), .B(new_n15110_), .ZN(new_n15111_));
  OAI21_X1   g12675(.A1(new_n15111_), .A2(pi0143), .B(new_n14851_), .ZN(new_n15112_));
  AOI21_X1   g12676(.A1(new_n5336_), .A2(new_n13597_), .B(new_n3265_), .ZN(new_n15113_));
  NAND3_X1   g12677(.A1(new_n13416_), .A2(new_n13798_), .A3(new_n2627_), .ZN(new_n15114_));
  OAI21_X1   g12678(.A1(new_n13651_), .A2(new_n13634_), .B(pi0039), .ZN(new_n15115_));
  AOI21_X1   g12679(.A1(new_n15115_), .A2(new_n15114_), .B(pi0038), .ZN(new_n15116_));
  NOR3_X1    g12680(.A1(new_n15116_), .A2(new_n10695_), .A3(new_n15113_), .ZN(new_n15117_));
  OAI21_X1   g12681(.A1(new_n15117_), .A2(new_n15112_), .B(pi0687), .ZN(new_n15118_));
  NOR3_X1    g12682(.A1(new_n13794_), .A2(new_n13786_), .A3(new_n2627_), .ZN(new_n15119_));
  AOI21_X1   g12683(.A1(new_n13805_), .A2(new_n13807_), .B(pi0039), .ZN(new_n15120_));
  OAI21_X1   g12684(.A1(new_n15119_), .A2(new_n15120_), .B(new_n3265_), .ZN(new_n15121_));
  OAI21_X1   g12685(.A1(new_n15121_), .A2(new_n10695_), .B(pi0774), .ZN(new_n15122_));
  NOR3_X1    g12686(.A1(new_n14643_), .A2(new_n3265_), .A3(pi0039), .ZN(new_n15123_));
  NOR2_X1    g12687(.A1(new_n13397_), .A2(new_n13571_), .ZN(new_n15124_));
  NOR2_X1    g12688(.A1(new_n15124_), .A2(new_n3265_), .ZN(new_n15125_));
  INV_X1     g12689(.I(new_n15125_), .ZN(new_n15126_));
  OAI21_X1   g12690(.A1(new_n13809_), .A2(new_n13406_), .B(new_n2627_), .ZN(new_n15127_));
  OAI21_X1   g12691(.A1(new_n13745_), .A2(new_n13754_), .B(pi0039), .ZN(new_n15128_));
  NAND3_X1   g12692(.A1(new_n15128_), .A2(new_n15127_), .A3(new_n3265_), .ZN(new_n15129_));
  AOI21_X1   g12693(.A1(new_n15129_), .A2(new_n15126_), .B(pi0143), .ZN(new_n15130_));
  NOR3_X1    g12694(.A1(new_n15130_), .A2(new_n15122_), .A3(new_n15123_), .ZN(new_n15131_));
  OAI21_X1   g12695(.A1(new_n15118_), .A2(new_n15131_), .B(new_n2609_), .ZN(new_n15132_));
  OAI21_X1   g12696(.A1(new_n15132_), .A2(new_n15106_), .B(new_n15005_), .ZN(new_n15133_));
  NAND2_X1   g12697(.A1(new_n15133_), .A2(pi0625), .ZN(new_n15134_));
  NAND2_X1   g12698(.A1(new_n15018_), .A2(new_n15005_), .ZN(new_n15135_));
  NAND2_X1   g12699(.A1(new_n15135_), .A2(new_n13521_), .ZN(new_n15136_));
  AOI21_X1   g12700(.A1(new_n15134_), .A2(new_n15136_), .B(new_n12841_), .ZN(new_n15137_));
  NOR3_X1    g12701(.A1(new_n15137_), .A2(new_n13560_), .A3(new_n15071_), .ZN(new_n15138_));
  AOI21_X1   g12702(.A1(new_n15018_), .A2(new_n15005_), .B(new_n13521_), .ZN(new_n15139_));
  AOI21_X1   g12703(.A1(new_n15133_), .A2(new_n13521_), .B(new_n15139_), .ZN(new_n15140_));
  OAI21_X1   g12704(.A1(new_n15140_), .A2(pi1153), .B(new_n15074_), .ZN(new_n15141_));
  OAI21_X1   g12705(.A1(new_n15141_), .A2(pi0608), .B(pi0778), .ZN(new_n15142_));
  NAND2_X1   g12706(.A1(new_n15133_), .A2(new_n12758_), .ZN(new_n15143_));
  OAI21_X1   g12707(.A1(new_n15142_), .A2(new_n15138_), .B(new_n15143_), .ZN(new_n15144_));
  NAND2_X1   g12708(.A1(new_n15144_), .A2(new_n12764_), .ZN(new_n15145_));
  INV_X1     g12709(.I(new_n15145_), .ZN(new_n15146_));
  AOI21_X1   g12710(.A1(new_n15023_), .A2(new_n12770_), .B(new_n13829_), .ZN(new_n15147_));
  AOI21_X1   g12711(.A1(new_n15076_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n15148_));
  OAI21_X1   g12712(.A1(new_n15144_), .A2(new_n12766_), .B(new_n15148_), .ZN(new_n15149_));
  NAND2_X1   g12713(.A1(new_n15149_), .A2(new_n15147_), .ZN(new_n15150_));
  NOR2_X1    g12714(.A1(new_n15027_), .A2(pi0660), .ZN(new_n15151_));
  AOI21_X1   g12715(.A1(new_n15076_), .A2(pi0609), .B(pi1155), .ZN(new_n15152_));
  OAI21_X1   g12716(.A1(new_n15144_), .A2(pi0609), .B(new_n15152_), .ZN(new_n15153_));
  AOI21_X1   g12717(.A1(new_n15153_), .A2(new_n15151_), .B(new_n12764_), .ZN(new_n15154_));
  AOI21_X1   g12718(.A1(new_n15154_), .A2(new_n15150_), .B(new_n15146_), .ZN(new_n15155_));
  OR2_X2     g12719(.A1(new_n15155_), .A2(pi0781), .Z(new_n15156_));
  OAI21_X1   g12720(.A1(new_n15031_), .A2(pi1154), .B(pi0627), .ZN(new_n15157_));
  NOR2_X1    g12721(.A1(new_n15077_), .A2(pi0618), .ZN(new_n15158_));
  NOR2_X1    g12722(.A1(new_n15158_), .A2(new_n12785_), .ZN(new_n15159_));
  NAND2_X1   g12723(.A1(new_n15155_), .A2(pi0618), .ZN(new_n15160_));
  AOI21_X1   g12724(.A1(new_n15160_), .A2(new_n15159_), .B(new_n15157_), .ZN(new_n15161_));
  OAI21_X1   g12725(.A1(new_n15034_), .A2(new_n12785_), .B(new_n12880_), .ZN(new_n15162_));
  OAI21_X1   g12726(.A1(new_n15077_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n15163_));
  AOI21_X1   g12727(.A1(new_n15155_), .A2(new_n12781_), .B(new_n15163_), .ZN(new_n15164_));
  OAI21_X1   g12728(.A1(new_n15164_), .A2(new_n15162_), .B(pi0781), .ZN(new_n15165_));
  OAI21_X1   g12729(.A1(new_n15165_), .A2(new_n15161_), .B(new_n15156_), .ZN(new_n15166_));
  AND2_X2    g12730(.A1(new_n15166_), .A2(new_n12796_), .Z(new_n15167_));
  AOI21_X1   g12731(.A1(new_n15038_), .A2(new_n12791_), .B(new_n12895_), .ZN(new_n15168_));
  AOI21_X1   g12732(.A1(new_n15079_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n15169_));
  OAI21_X1   g12733(.A1(new_n15166_), .A2(new_n12793_), .B(new_n15169_), .ZN(new_n15170_));
  NAND2_X1   g12734(.A1(new_n15170_), .A2(new_n15168_), .ZN(new_n15171_));
  AOI21_X1   g12735(.A1(new_n15041_), .A2(pi1159), .B(pi0648), .ZN(new_n15172_));
  AOI21_X1   g12736(.A1(new_n15079_), .A2(pi0619), .B(pi1159), .ZN(new_n15173_));
  OAI21_X1   g12737(.A1(new_n15166_), .A2(pi0619), .B(new_n15173_), .ZN(new_n15174_));
  AOI21_X1   g12738(.A1(new_n15174_), .A2(new_n15172_), .B(new_n12796_), .ZN(new_n15175_));
  AOI21_X1   g12739(.A1(new_n15175_), .A2(new_n15171_), .B(new_n15167_), .ZN(new_n15176_));
  OAI21_X1   g12740(.A1(new_n15176_), .A2(new_n12747_), .B(new_n15105_), .ZN(new_n15177_));
  NAND2_X1   g12741(.A1(new_n15177_), .A2(new_n15104_), .ZN(new_n15178_));
  OAI21_X1   g12742(.A1(new_n15048_), .A2(pi1158), .B(new_n12904_), .ZN(new_n15179_));
  AOI21_X1   g12743(.A1(new_n15081_), .A2(pi0626), .B(pi0641), .ZN(new_n15180_));
  OAI21_X1   g12744(.A1(new_n15176_), .A2(pi0626), .B(new_n15180_), .ZN(new_n15181_));
  AOI21_X1   g12745(.A1(new_n15181_), .A2(new_n15179_), .B(new_n12808_), .ZN(new_n15182_));
  AND2_X2    g12746(.A1(new_n15176_), .A2(new_n12808_), .Z(new_n15183_));
  AOI21_X1   g12747(.A1(new_n15182_), .A2(new_n15178_), .B(new_n15183_), .ZN(new_n15184_));
  OAI21_X1   g12748(.A1(new_n15184_), .A2(new_n12920_), .B(new_n15103_), .ZN(new_n15185_));
  NAND2_X1   g12749(.A1(new_n15185_), .A2(new_n15102_), .ZN(new_n15186_));
  NOR2_X1    g12750(.A1(new_n15089_), .A2(pi0629), .ZN(new_n15187_));
  AOI21_X1   g12751(.A1(new_n15050_), .A2(pi0628), .B(pi1156), .ZN(new_n15188_));
  OAI21_X1   g12752(.A1(new_n15184_), .A2(pi0628), .B(new_n15188_), .ZN(new_n15189_));
  AOI21_X1   g12753(.A1(new_n15189_), .A2(new_n15187_), .B(new_n12937_), .ZN(new_n15190_));
  AND2_X2    g12754(.A1(new_n15184_), .A2(new_n12937_), .Z(new_n15191_));
  AOI21_X1   g12755(.A1(new_n15190_), .A2(new_n15186_), .B(new_n15191_), .ZN(new_n15192_));
  OR2_X2     g12756(.A1(new_n15192_), .A2(pi0787), .Z(new_n15193_));
  OR2_X2     g12757(.A1(new_n15095_), .A2(new_n12981_), .Z(new_n15194_));
  AOI21_X1   g12758(.A1(new_n15053_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n15195_));
  NAND2_X1   g12759(.A1(new_n15192_), .A2(pi0647), .ZN(new_n15196_));
  AOI21_X1   g12760(.A1(new_n15196_), .A2(new_n15195_), .B(new_n15194_), .ZN(new_n15197_));
  NAND2_X1   g12761(.A1(new_n15098_), .A2(new_n12981_), .ZN(new_n15198_));
  OAI21_X1   g12762(.A1(new_n15054_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n15199_));
  AOI21_X1   g12763(.A1(new_n15192_), .A2(new_n12741_), .B(new_n15199_), .ZN(new_n15200_));
  OAI21_X1   g12764(.A1(new_n15200_), .A2(new_n15198_), .B(pi0787), .ZN(new_n15201_));
  OAI21_X1   g12765(.A1(new_n15201_), .A2(new_n15197_), .B(new_n15193_), .ZN(new_n15202_));
  OAI21_X1   g12766(.A1(new_n15202_), .A2(pi0644), .B(new_n15101_), .ZN(new_n15203_));
  NAND2_X1   g12767(.A1(new_n15203_), .A2(new_n15058_), .ZN(new_n15204_));
  AOI21_X1   g12768(.A1(new_n15002_), .A2(new_n12975_), .B(pi0715), .ZN(new_n15205_));
  NAND2_X1   g12769(.A1(new_n15056_), .A2(pi0644), .ZN(new_n15206_));
  AOI21_X1   g12770(.A1(new_n15206_), .A2(new_n15205_), .B(new_n12739_), .ZN(new_n15207_));
  NOR2_X1    g12771(.A1(new_n15100_), .A2(pi0644), .ZN(new_n15208_));
  AOI21_X1   g12772(.A1(new_n15202_), .A2(pi0644), .B(new_n15208_), .ZN(new_n15209_));
  OAI21_X1   g12773(.A1(new_n15209_), .A2(new_n12740_), .B(new_n15207_), .ZN(new_n15210_));
  NAND3_X1   g12774(.A1(new_n15210_), .A2(new_n15204_), .A3(pi0790), .ZN(new_n15211_));
  AOI21_X1   g12775(.A1(new_n15202_), .A2(new_n13000_), .B(po1038), .ZN(new_n15212_));
  NAND2_X1   g12776(.A1(new_n15211_), .A2(new_n15212_), .ZN(new_n15213_));
  AOI21_X1   g12777(.A1(new_n15213_), .A2(new_n15001_), .B(new_n15000_), .ZN(po0300));
  NOR2_X1    g12778(.A1(new_n3042_), .A2(new_n8058_), .ZN(new_n15215_));
  INV_X1     g12779(.I(new_n15215_), .ZN(new_n15216_));
  NAND2_X1   g12780(.A1(new_n12826_), .A2(pi0736), .ZN(new_n15217_));
  NAND2_X1   g12781(.A1(new_n15217_), .A2(new_n15216_), .ZN(new_n15218_));
  INV_X1     g12782(.I(new_n15218_), .ZN(new_n15219_));
  NOR2_X1    g12783(.A1(new_n15217_), .A2(new_n13521_), .ZN(new_n15220_));
  NOR3_X1    g12784(.A1(new_n15220_), .A2(new_n12841_), .A3(new_n15215_), .ZN(new_n15221_));
  INV_X1     g12785(.I(new_n15221_), .ZN(new_n15222_));
  OAI21_X1   g12786(.A1(new_n15219_), .A2(new_n15220_), .B(new_n12841_), .ZN(new_n15223_));
  NAND3_X1   g12787(.A1(new_n15222_), .A2(new_n15223_), .A3(pi0778), .ZN(new_n15224_));
  OAI21_X1   g12788(.A1(pi0778), .A2(new_n15219_), .B(new_n15224_), .ZN(new_n15225_));
  AND2_X2    g12789(.A1(new_n15225_), .A2(new_n14291_), .Z(new_n15226_));
  NAND2_X1   g12790(.A1(new_n15226_), .A2(new_n12952_), .ZN(new_n15227_));
  NAND2_X1   g12791(.A1(new_n15227_), .A2(new_n12981_), .ZN(new_n15228_));
  NOR2_X1    g12792(.A1(new_n12770_), .A2(pi0609), .ZN(new_n15229_));
  NOR2_X1    g12793(.A1(new_n12766_), .A2(pi1155), .ZN(new_n15230_));
  OAI21_X1   g12794(.A1(new_n15229_), .A2(new_n15230_), .B(pi0785), .ZN(new_n15231_));
  INV_X1     g12795(.I(new_n15231_), .ZN(new_n15232_));
  INV_X1     g12796(.I(pi0758), .ZN(new_n15233_));
  NOR2_X1    g12797(.A1(new_n13340_), .A2(new_n15233_), .ZN(new_n15234_));
  INV_X1     g12798(.I(new_n15234_), .ZN(new_n15235_));
  NOR2_X1    g12799(.A1(new_n15235_), .A2(new_n15232_), .ZN(new_n15236_));
  INV_X1     g12800(.I(new_n15236_), .ZN(new_n15237_));
  XNOR2_X1   g12801(.A1(pi0618), .A2(pi1154), .ZN(new_n15238_));
  NOR2_X1    g12802(.A1(new_n15238_), .A2(new_n12779_), .ZN(new_n15239_));
  NOR2_X1    g12803(.A1(new_n12760_), .A2(new_n15239_), .ZN(new_n15240_));
  INV_X1     g12804(.I(new_n15240_), .ZN(new_n15241_));
  NOR2_X1    g12805(.A1(pi0619), .A2(pi1159), .ZN(new_n15242_));
  NOR2_X1    g12806(.A1(new_n12793_), .A2(new_n12791_), .ZN(new_n15243_));
  NOR3_X1    g12807(.A1(new_n15243_), .A2(new_n12796_), .A3(new_n15242_), .ZN(new_n15244_));
  NOR2_X1    g12808(.A1(new_n15241_), .A2(new_n15244_), .ZN(new_n15245_));
  INV_X1     g12809(.I(new_n15245_), .ZN(new_n15246_));
  NOR2_X1    g12810(.A1(new_n15237_), .A2(new_n15246_), .ZN(new_n15247_));
  INV_X1     g12811(.I(new_n15247_), .ZN(new_n15248_));
  NOR2_X1    g12812(.A1(new_n15248_), .A2(new_n12818_), .ZN(new_n15249_));
  NAND2_X1   g12813(.A1(new_n15249_), .A2(new_n13384_), .ZN(new_n15250_));
  OAI21_X1   g12814(.A1(new_n15250_), .A2(new_n12981_), .B(pi1157), .ZN(new_n15251_));
  AOI21_X1   g12815(.A1(new_n15228_), .A2(pi0647), .B(new_n15251_), .ZN(new_n15252_));
  NOR2_X1    g12816(.A1(new_n15227_), .A2(pi0647), .ZN(new_n15253_));
  AOI21_X1   g12817(.A1(new_n15250_), .A2(pi0647), .B(pi0630), .ZN(new_n15254_));
  NOR3_X1    g12818(.A1(new_n15253_), .A2(pi1157), .A3(new_n15254_), .ZN(new_n15255_));
  NOR2_X1    g12819(.A1(new_n15215_), .A2(new_n12972_), .ZN(new_n15256_));
  OAI21_X1   g12820(.A1(new_n15255_), .A2(new_n15252_), .B(new_n15256_), .ZN(new_n15257_));
  NAND2_X1   g12821(.A1(new_n15247_), .A2(new_n12747_), .ZN(new_n15258_));
  AOI21_X1   g12822(.A1(new_n15258_), .A2(new_n15216_), .B(pi1158), .ZN(new_n15259_));
  AOI21_X1   g12823(.A1(new_n15225_), .A2(new_n14289_), .B(new_n15215_), .ZN(new_n15260_));
  INV_X1     g12824(.I(new_n15260_), .ZN(new_n15261_));
  OAI21_X1   g12825(.A1(new_n12911_), .A2(new_n15215_), .B(new_n15261_), .ZN(new_n15262_));
  NOR3_X1    g12826(.A1(new_n15262_), .A2(pi0626), .A3(new_n12745_), .ZN(new_n15263_));
  NOR3_X1    g12827(.A1(new_n15263_), .A2(new_n12814_), .A3(new_n15259_), .ZN(new_n15264_));
  INV_X1     g12828(.I(new_n12748_), .ZN(new_n15265_));
  OAI21_X1   g12829(.A1(new_n15248_), .A2(new_n12747_), .B(new_n15216_), .ZN(new_n15266_));
  AOI21_X1   g12830(.A1(new_n15266_), .A2(pi1158), .B(pi0641), .ZN(new_n15267_));
  OAI21_X1   g12831(.A1(new_n15262_), .A2(new_n15265_), .B(new_n15267_), .ZN(new_n15268_));
  NAND2_X1   g12832(.A1(new_n15268_), .A2(pi0788), .ZN(new_n15269_));
  NOR2_X1    g12833(.A1(new_n15264_), .A2(new_n15269_), .ZN(new_n15270_));
  NOR2_X1    g12834(.A1(new_n15241_), .A2(pi0619), .ZN(new_n15271_));
  NAND2_X1   g12835(.A1(new_n15236_), .A2(new_n15271_), .ZN(new_n15272_));
  AND3_X2    g12836(.A1(new_n15272_), .A2(new_n12791_), .A3(new_n15216_), .Z(new_n15273_));
  NOR2_X1    g12837(.A1(new_n15225_), .A2(pi0609), .ZN(new_n15274_));
  INV_X1     g12838(.I(pi0736), .ZN(new_n15275_));
  NOR2_X1    g12839(.A1(new_n14328_), .A2(new_n15275_), .ZN(new_n15276_));
  NOR3_X1    g12840(.A1(new_n15276_), .A2(new_n15234_), .A3(new_n15215_), .ZN(new_n15277_));
  NAND2_X1   g12841(.A1(new_n15277_), .A2(new_n12758_), .ZN(new_n15278_));
  NOR2_X1    g12842(.A1(new_n14330_), .A2(new_n15275_), .ZN(new_n15279_));
  INV_X1     g12843(.I(new_n15279_), .ZN(new_n15280_));
  NAND4_X1   g12844(.A1(new_n15280_), .A2(pi1153), .A3(new_n15216_), .A4(new_n15235_), .ZN(new_n15281_));
  NAND3_X1   g12845(.A1(new_n15281_), .A2(pi0608), .A3(new_n15223_), .ZN(new_n15282_));
  OAI21_X1   g12846(.A1(new_n15279_), .A2(new_n15277_), .B(new_n12841_), .ZN(new_n15283_));
  NAND3_X1   g12847(.A1(new_n15283_), .A2(new_n13560_), .A3(new_n15222_), .ZN(new_n15284_));
  NAND3_X1   g12848(.A1(new_n15282_), .A2(pi0778), .A3(new_n15284_), .ZN(new_n15285_));
  AOI21_X1   g12849(.A1(new_n15285_), .A2(new_n15278_), .B(new_n12766_), .ZN(new_n15286_));
  OAI21_X1   g12850(.A1(new_n15286_), .A2(new_n15274_), .B(pi1155), .ZN(new_n15287_));
  NAND2_X1   g12851(.A1(new_n15234_), .A2(new_n13353_), .ZN(new_n15288_));
  NAND3_X1   g12852(.A1(new_n15288_), .A2(new_n12770_), .A3(new_n15216_), .ZN(new_n15289_));
  NAND3_X1   g12853(.A1(new_n15287_), .A2(pi0660), .A3(new_n15289_), .ZN(new_n15290_));
  NAND2_X1   g12854(.A1(new_n15285_), .A2(new_n15278_), .ZN(new_n15291_));
  NOR2_X1    g12855(.A1(new_n15225_), .A2(new_n12766_), .ZN(new_n15292_));
  AOI21_X1   g12856(.A1(new_n15291_), .A2(new_n12766_), .B(new_n15292_), .ZN(new_n15293_));
  AOI21_X1   g12857(.A1(new_n15234_), .A2(new_n12772_), .B(new_n12770_), .ZN(new_n15294_));
  AOI21_X1   g12858(.A1(new_n15294_), .A2(new_n15216_), .B(pi0660), .ZN(new_n15295_));
  OAI21_X1   g12859(.A1(new_n15293_), .A2(pi1155), .B(new_n15295_), .ZN(new_n15296_));
  NAND3_X1   g12860(.A1(new_n15290_), .A2(new_n15296_), .A3(pi0785), .ZN(new_n15297_));
  NAND2_X1   g12861(.A1(new_n15291_), .A2(new_n12764_), .ZN(new_n15298_));
  NAND2_X1   g12862(.A1(new_n15297_), .A2(new_n15298_), .ZN(new_n15299_));
  NAND2_X1   g12863(.A1(new_n15299_), .A2(pi0618), .ZN(new_n15300_));
  AOI21_X1   g12864(.A1(new_n15225_), .A2(new_n12870_), .B(new_n15215_), .ZN(new_n15301_));
  NAND2_X1   g12865(.A1(new_n15301_), .A2(new_n12781_), .ZN(new_n15302_));
  AOI21_X1   g12866(.A1(new_n15300_), .A2(new_n15302_), .B(new_n12785_), .ZN(new_n15303_));
  NAND2_X1   g12867(.A1(new_n12761_), .A2(new_n12781_), .ZN(new_n15304_));
  OAI21_X1   g12868(.A1(new_n15237_), .A2(new_n15304_), .B(new_n12785_), .ZN(new_n15305_));
  NOR2_X1    g12869(.A1(new_n15305_), .A2(new_n15215_), .ZN(new_n15306_));
  NOR3_X1    g12870(.A1(new_n15303_), .A2(new_n12880_), .A3(new_n15306_), .ZN(new_n15307_));
  NAND2_X1   g12871(.A1(new_n15301_), .A2(pi0618), .ZN(new_n15308_));
  NAND2_X1   g12872(.A1(new_n15299_), .A2(new_n12781_), .ZN(new_n15309_));
  NAND2_X1   g12873(.A1(new_n15309_), .A2(new_n15308_), .ZN(new_n15310_));
  NAND2_X1   g12874(.A1(new_n12761_), .A2(pi0618), .ZN(new_n15311_));
  OAI21_X1   g12875(.A1(new_n15237_), .A2(new_n15311_), .B(pi1154), .ZN(new_n15312_));
  OAI21_X1   g12876(.A1(new_n15312_), .A2(new_n15215_), .B(new_n12880_), .ZN(new_n15313_));
  AOI21_X1   g12877(.A1(new_n15310_), .A2(new_n12785_), .B(new_n15313_), .ZN(new_n15314_));
  OR3_X2     g12878(.A1(new_n15307_), .A2(new_n12779_), .A3(new_n15314_), .Z(new_n15315_));
  NAND2_X1   g12879(.A1(new_n15299_), .A2(new_n12779_), .ZN(new_n15316_));
  NAND2_X1   g12880(.A1(new_n15315_), .A2(new_n15316_), .ZN(new_n15317_));
  NAND2_X1   g12881(.A1(new_n15317_), .A2(pi0619), .ZN(new_n15318_));
  NAND2_X1   g12882(.A1(new_n15260_), .A2(new_n12793_), .ZN(new_n15319_));
  AOI21_X1   g12883(.A1(new_n15318_), .A2(new_n15319_), .B(new_n12791_), .ZN(new_n15320_));
  NOR3_X1    g12884(.A1(new_n15320_), .A2(new_n12895_), .A3(new_n15273_), .ZN(new_n15321_));
  NAND2_X1   g12885(.A1(new_n15317_), .A2(new_n12793_), .ZN(new_n15322_));
  OAI21_X1   g12886(.A1(new_n12793_), .A2(new_n15261_), .B(new_n15322_), .ZN(new_n15323_));
  NAND3_X1   g12887(.A1(new_n15236_), .A2(new_n15240_), .A3(pi0619), .ZN(new_n15324_));
  NAND3_X1   g12888(.A1(new_n15324_), .A2(pi1159), .A3(new_n15216_), .ZN(new_n15325_));
  NAND2_X1   g12889(.A1(new_n15325_), .A2(new_n12895_), .ZN(new_n15326_));
  AOI21_X1   g12890(.A1(new_n15323_), .A2(new_n12791_), .B(new_n15326_), .ZN(new_n15327_));
  OR3_X2     g12891(.A1(new_n15327_), .A2(new_n12796_), .A3(new_n15321_), .Z(new_n15328_));
  AOI21_X1   g12892(.A1(new_n15317_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n15329_));
  AOI21_X1   g12893(.A1(new_n15328_), .A2(new_n15329_), .B(new_n15270_), .ZN(new_n15330_));
  OAI21_X1   g12894(.A1(new_n15249_), .A2(pi0628), .B(pi0629), .ZN(new_n15331_));
  NAND2_X1   g12895(.A1(new_n15226_), .A2(pi0628), .ZN(new_n15332_));
  NAND3_X1   g12896(.A1(new_n15332_), .A2(pi1156), .A3(new_n15331_), .ZN(new_n15333_));
  INV_X1     g12897(.I(new_n15249_), .ZN(new_n15334_));
  NOR2_X1    g12898(.A1(new_n15226_), .A2(new_n12919_), .ZN(new_n15335_));
  OAI22_X1   g12899(.A1(new_n15335_), .A2(pi0628), .B1(pi0629), .B2(new_n15334_), .ZN(new_n15336_));
  OAI21_X1   g12900(.A1(new_n15336_), .A2(pi1156), .B(new_n15333_), .ZN(new_n15337_));
  NAND2_X1   g12901(.A1(new_n15337_), .A2(new_n15216_), .ZN(new_n15338_));
  NOR2_X1    g12902(.A1(new_n15338_), .A2(new_n12937_), .ZN(new_n15339_));
  AOI21_X1   g12903(.A1(new_n12942_), .A2(new_n12950_), .B(new_n12937_), .ZN(new_n15340_));
  AOI21_X1   g12904(.A1(new_n12983_), .A2(new_n14299_), .B(new_n12972_), .ZN(new_n15341_));
  AOI21_X1   g12905(.A1(new_n15338_), .A2(new_n15340_), .B(new_n15341_), .ZN(new_n15342_));
  OAI21_X1   g12906(.A1(new_n15330_), .A2(new_n15339_), .B(new_n15342_), .ZN(new_n15343_));
  NAND2_X1   g12907(.A1(new_n15343_), .A2(new_n15257_), .ZN(new_n15344_));
  NAND2_X1   g12908(.A1(new_n15344_), .A2(new_n13000_), .ZN(new_n15345_));
  AOI21_X1   g12909(.A1(new_n15343_), .A2(new_n15257_), .B(pi0644), .ZN(new_n15346_));
  OAI21_X1   g12910(.A1(new_n15227_), .A2(new_n14300_), .B(new_n15216_), .ZN(new_n15347_));
  NOR2_X1    g12911(.A1(new_n15347_), .A2(new_n12975_), .ZN(new_n15348_));
  OAI21_X1   g12912(.A1(new_n15346_), .A2(new_n15348_), .B(new_n12740_), .ZN(new_n15349_));
  NOR2_X1    g12913(.A1(new_n15250_), .A2(new_n12984_), .ZN(new_n15350_));
  NAND2_X1   g12914(.A1(new_n15350_), .A2(new_n12975_), .ZN(new_n15351_));
  NAND3_X1   g12915(.A1(new_n15351_), .A2(pi0715), .A3(new_n15216_), .ZN(new_n15352_));
  NAND3_X1   g12916(.A1(new_n15349_), .A2(new_n12739_), .A3(new_n15352_), .ZN(new_n15353_));
  NOR2_X1    g12917(.A1(new_n15347_), .A2(pi0644), .ZN(new_n15354_));
  AOI21_X1   g12918(.A1(new_n15344_), .A2(pi0644), .B(new_n15354_), .ZN(new_n15355_));
  AOI21_X1   g12919(.A1(new_n15350_), .A2(pi0644), .B(pi0715), .ZN(new_n15356_));
  AOI21_X1   g12920(.A1(new_n15356_), .A2(new_n15216_), .B(new_n12739_), .ZN(new_n15357_));
  OAI21_X1   g12921(.A1(new_n15355_), .A2(new_n12740_), .B(new_n15357_), .ZN(new_n15358_));
  NAND3_X1   g12922(.A1(new_n15353_), .A2(new_n15358_), .A3(pi0790), .ZN(new_n15359_));
  AOI21_X1   g12923(.A1(new_n15359_), .A2(new_n15345_), .B(new_n12738_), .ZN(new_n15360_));
  AOI21_X1   g12924(.A1(pi0057), .A2(pi0144), .B(pi0832), .ZN(new_n15361_));
  NAND2_X1   g12925(.A1(new_n13192_), .A2(pi0144), .ZN(new_n15362_));
  NOR2_X1    g12926(.A1(new_n15362_), .A2(new_n13521_), .ZN(new_n15363_));
  NOR2_X1    g12927(.A1(new_n2610_), .A2(new_n15275_), .ZN(new_n15364_));
  NOR2_X1    g12928(.A1(new_n14122_), .A2(pi0144), .ZN(new_n15365_));
  NOR2_X1    g12929(.A1(new_n14118_), .A2(new_n8058_), .ZN(new_n15366_));
  OAI21_X1   g12930(.A1(new_n15366_), .A2(new_n15365_), .B(new_n3265_), .ZN(new_n15367_));
  NOR2_X1    g12931(.A1(new_n13344_), .A2(new_n8058_), .ZN(new_n15368_));
  NOR2_X1    g12932(.A1(new_n13398_), .A2(new_n15368_), .ZN(new_n15369_));
  NOR2_X1    g12933(.A1(new_n15369_), .A2(new_n3265_), .ZN(new_n15370_));
  INV_X1     g12934(.I(new_n15370_), .ZN(new_n15371_));
  NAND3_X1   g12935(.A1(new_n15367_), .A2(new_n15364_), .A3(new_n15371_), .ZN(new_n15372_));
  INV_X1     g12936(.I(new_n15364_), .ZN(new_n15373_));
  NAND2_X1   g12937(.A1(new_n15362_), .A2(new_n15373_), .ZN(new_n15374_));
  AND3_X2    g12938(.A1(new_n15372_), .A2(new_n13521_), .A3(new_n15374_), .Z(new_n15375_));
  OAI21_X1   g12939(.A1(new_n15375_), .A2(new_n15363_), .B(new_n12841_), .ZN(new_n15376_));
  NAND3_X1   g12940(.A1(new_n15372_), .A2(new_n15374_), .A3(pi0625), .ZN(new_n15377_));
  INV_X1     g12941(.I(new_n15362_), .ZN(new_n15378_));
  NAND2_X1   g12942(.A1(new_n15378_), .A2(new_n13521_), .ZN(new_n15379_));
  AOI21_X1   g12943(.A1(new_n15377_), .A2(new_n15379_), .B(new_n12841_), .ZN(new_n15380_));
  NOR2_X1    g12944(.A1(new_n15380_), .A2(new_n12758_), .ZN(new_n15381_));
  AOI21_X1   g12945(.A1(new_n15372_), .A2(new_n15374_), .B(pi0778), .ZN(new_n15382_));
  AOI21_X1   g12946(.A1(new_n15381_), .A2(new_n15376_), .B(new_n15382_), .ZN(new_n15383_));
  NOR2_X1    g12947(.A1(new_n15362_), .A2(new_n12870_), .ZN(new_n15384_));
  AOI21_X1   g12948(.A1(new_n15383_), .A2(new_n12870_), .B(new_n15384_), .ZN(new_n15385_));
  NOR2_X1    g12949(.A1(new_n15378_), .A2(new_n12888_), .ZN(new_n15386_));
  AOI21_X1   g12950(.A1(new_n15385_), .A2(new_n12888_), .B(new_n15386_), .ZN(new_n15387_));
  NOR2_X1    g12951(.A1(new_n15362_), .A2(new_n12911_), .ZN(new_n15388_));
  AOI21_X1   g12952(.A1(new_n15387_), .A2(new_n12911_), .B(new_n15388_), .ZN(new_n15389_));
  NOR2_X1    g12953(.A1(new_n15378_), .A2(new_n13392_), .ZN(new_n15390_));
  AOI21_X1   g12954(.A1(new_n15389_), .A2(new_n13392_), .B(new_n15390_), .ZN(new_n15391_));
  NAND2_X1   g12955(.A1(new_n15391_), .A2(new_n12920_), .ZN(new_n15392_));
  NAND2_X1   g12956(.A1(new_n15378_), .A2(pi0628), .ZN(new_n15393_));
  AOI21_X1   g12957(.A1(new_n15392_), .A2(new_n15393_), .B(pi1156), .ZN(new_n15394_));
  OR2_X2     g12958(.A1(new_n15394_), .A2(new_n12919_), .Z(new_n15395_));
  NOR2_X1    g12959(.A1(new_n2609_), .A2(new_n8058_), .ZN(new_n15396_));
  INV_X1     g12960(.I(new_n15396_), .ZN(new_n15397_));
  NOR2_X1    g12961(.A1(new_n5337_), .A2(new_n15235_), .ZN(new_n15398_));
  OAI21_X1   g12962(.A1(new_n15368_), .A2(new_n15398_), .B(pi0038), .ZN(new_n15399_));
  INV_X1     g12963(.I(new_n15399_), .ZN(new_n15400_));
  NAND3_X1   g12964(.A1(new_n13245_), .A2(new_n8058_), .A3(pi0758), .ZN(new_n15401_));
  NAND2_X1   g12965(.A1(new_n13256_), .A2(pi0758), .ZN(new_n15402_));
  NAND2_X1   g12966(.A1(new_n13060_), .A2(new_n15233_), .ZN(new_n15403_));
  AOI21_X1   g12967(.A1(new_n15402_), .A2(new_n15403_), .B(pi0039), .ZN(new_n15404_));
  AOI21_X1   g12968(.A1(new_n13322_), .A2(new_n13332_), .B(new_n15233_), .ZN(new_n15405_));
  NOR3_X1    g12969(.A1(new_n13178_), .A2(new_n13188_), .A3(pi0758), .ZN(new_n15406_));
  NOR3_X1    g12970(.A1(new_n15405_), .A2(new_n15406_), .A3(new_n2627_), .ZN(new_n15407_));
  OAI21_X1   g12971(.A1(new_n15407_), .A2(new_n15404_), .B(pi0144), .ZN(new_n15408_));
  AOI21_X1   g12972(.A1(new_n15408_), .A2(new_n15401_), .B(pi0038), .ZN(new_n15409_));
  OAI21_X1   g12973(.A1(new_n15409_), .A2(new_n15400_), .B(new_n2609_), .ZN(new_n15410_));
  NAND2_X1   g12974(.A1(new_n15410_), .A2(new_n15397_), .ZN(new_n15411_));
  NAND2_X1   g12975(.A1(new_n15411_), .A2(new_n12761_), .ZN(new_n15412_));
  OAI21_X1   g12976(.A1(new_n12761_), .A2(new_n15362_), .B(new_n15412_), .ZN(new_n15413_));
  NOR2_X1    g12977(.A1(new_n15362_), .A2(new_n12766_), .ZN(new_n15414_));
  AOI21_X1   g12978(.A1(new_n15413_), .A2(new_n12766_), .B(new_n15414_), .ZN(new_n15415_));
  NOR2_X1    g12979(.A1(new_n15415_), .A2(pi1155), .ZN(new_n15416_));
  NOR2_X1    g12980(.A1(new_n15362_), .A2(pi0609), .ZN(new_n15417_));
  AOI21_X1   g12981(.A1(new_n15413_), .A2(pi0609), .B(new_n15417_), .ZN(new_n15418_));
  OAI21_X1   g12982(.A1(new_n15418_), .A2(new_n12770_), .B(pi0785), .ZN(new_n15419_));
  OAI22_X1   g12983(.A1(new_n15419_), .A2(new_n15416_), .B1(pi0785), .B2(new_n15413_), .ZN(new_n15420_));
  NAND2_X1   g12984(.A1(new_n15378_), .A2(pi0618), .ZN(new_n15421_));
  OAI21_X1   g12985(.A1(new_n15420_), .A2(pi0618), .B(new_n15421_), .ZN(new_n15422_));
  NAND2_X1   g12986(.A1(new_n15422_), .A2(new_n12785_), .ZN(new_n15423_));
  NAND2_X1   g12987(.A1(new_n15378_), .A2(new_n12781_), .ZN(new_n15424_));
  OAI21_X1   g12988(.A1(new_n15420_), .A2(new_n12781_), .B(new_n15424_), .ZN(new_n15425_));
  AOI21_X1   g12989(.A1(new_n15425_), .A2(pi1154), .B(new_n12779_), .ZN(new_n15426_));
  AOI22_X1   g12990(.A1(new_n15426_), .A2(new_n15423_), .B1(new_n12779_), .B2(new_n15420_), .ZN(new_n15427_));
  NOR2_X1    g12991(.A1(new_n15362_), .A2(new_n12793_), .ZN(new_n15428_));
  AOI21_X1   g12992(.A1(new_n15427_), .A2(new_n12793_), .B(new_n15428_), .ZN(new_n15429_));
  NOR2_X1    g12993(.A1(new_n15429_), .A2(pi1159), .ZN(new_n15430_));
  NOR2_X1    g12994(.A1(new_n15362_), .A2(pi0619), .ZN(new_n15431_));
  AOI21_X1   g12995(.A1(new_n15427_), .A2(pi0619), .B(new_n15431_), .ZN(new_n15432_));
  OAI21_X1   g12996(.A1(new_n15432_), .A2(new_n12791_), .B(pi0789), .ZN(new_n15433_));
  OAI22_X1   g12997(.A1(new_n15433_), .A2(new_n15430_), .B1(pi0789), .B2(new_n15427_), .ZN(new_n15434_));
  NOR2_X1    g12998(.A1(new_n15362_), .A2(pi0626), .ZN(new_n15435_));
  INV_X1     g12999(.I(new_n15435_), .ZN(new_n15436_));
  OAI21_X1   g13000(.A1(new_n15434_), .A2(new_n12747_), .B(new_n15436_), .ZN(new_n15437_));
  NAND2_X1   g13001(.A1(new_n15437_), .A2(pi1158), .ZN(new_n15438_));
  NOR2_X1    g13002(.A1(new_n15362_), .A2(new_n12747_), .ZN(new_n15439_));
  INV_X1     g13003(.I(new_n15439_), .ZN(new_n15440_));
  OAI21_X1   g13004(.A1(new_n15434_), .A2(pi0626), .B(new_n15440_), .ZN(new_n15441_));
  AOI21_X1   g13005(.A1(new_n15441_), .A2(new_n12745_), .B(new_n12808_), .ZN(new_n15442_));
  AOI22_X1   g13006(.A1(new_n15442_), .A2(new_n15438_), .B1(new_n12808_), .B2(new_n15434_), .ZN(new_n15443_));
  NOR2_X1    g13007(.A1(new_n15443_), .A2(pi0628), .ZN(new_n15444_));
  NOR2_X1    g13008(.A1(new_n15444_), .A2(new_n12742_), .ZN(new_n15445_));
  OAI21_X1   g13009(.A1(new_n15437_), .A2(pi0641), .B(pi1158), .ZN(new_n15446_));
  NOR2_X1    g13010(.A1(new_n15389_), .A2(pi0626), .ZN(new_n15447_));
  NOR2_X1    g13011(.A1(new_n15447_), .A2(new_n12814_), .ZN(new_n15448_));
  NOR3_X1    g13012(.A1(new_n15400_), .A2(new_n15275_), .A3(new_n15123_), .ZN(new_n15449_));
  AOI21_X1   g13013(.A1(new_n13692_), .A2(pi0144), .B(new_n15233_), .ZN(new_n15450_));
  OAI21_X1   g13014(.A1(new_n14187_), .A2(pi0144), .B(new_n15450_), .ZN(new_n15451_));
  OAI21_X1   g13015(.A1(new_n13794_), .A2(new_n13786_), .B(new_n8058_), .ZN(new_n15452_));
  OAI21_X1   g13016(.A1(new_n13745_), .A2(new_n13754_), .B(pi0144), .ZN(new_n15453_));
  NAND3_X1   g13017(.A1(new_n15453_), .A2(new_n15233_), .A3(new_n15452_), .ZN(new_n15454_));
  NAND3_X1   g13018(.A1(new_n15451_), .A2(new_n15454_), .A3(pi0039), .ZN(new_n15455_));
  AOI21_X1   g13019(.A1(new_n13416_), .A2(new_n13798_), .B(pi0144), .ZN(new_n15456_));
  NOR2_X1    g13020(.A1(new_n13800_), .A2(new_n8058_), .ZN(new_n15457_));
  OAI21_X1   g13021(.A1(new_n15457_), .A2(new_n15456_), .B(pi0758), .ZN(new_n15458_));
  NOR3_X1    g13022(.A1(new_n13809_), .A2(new_n13406_), .A3(new_n8058_), .ZN(new_n15459_));
  AOI21_X1   g13023(.A1(new_n13805_), .A2(new_n13807_), .B(pi0144), .ZN(new_n15460_));
  OAI21_X1   g13024(.A1(new_n15459_), .A2(new_n15460_), .B(new_n15233_), .ZN(new_n15461_));
  NAND3_X1   g13025(.A1(new_n15458_), .A2(new_n15461_), .A3(new_n2627_), .ZN(new_n15462_));
  NAND3_X1   g13026(.A1(new_n15455_), .A2(new_n15462_), .A3(new_n3265_), .ZN(new_n15463_));
  AOI21_X1   g13027(.A1(new_n15463_), .A2(new_n15449_), .B(new_n2610_), .ZN(new_n15464_));
  NOR2_X1    g13028(.A1(new_n15409_), .A2(new_n15400_), .ZN(new_n15465_));
  NAND2_X1   g13029(.A1(new_n15465_), .A2(new_n15275_), .ZN(new_n15466_));
  AOI21_X1   g13030(.A1(new_n15464_), .A2(new_n15466_), .B(new_n15396_), .ZN(new_n15467_));
  NOR2_X1    g13031(.A1(new_n15467_), .A2(new_n13521_), .ZN(new_n15468_));
  AOI21_X1   g13032(.A1(new_n15410_), .A2(new_n15397_), .B(pi0625), .ZN(new_n15469_));
  OAI21_X1   g13033(.A1(new_n15468_), .A2(new_n15469_), .B(pi1153), .ZN(new_n15470_));
  NAND3_X1   g13034(.A1(new_n15470_), .A2(pi0608), .A3(new_n15376_), .ZN(new_n15471_));
  NAND2_X1   g13035(.A1(new_n15411_), .A2(pi0625), .ZN(new_n15472_));
  OAI21_X1   g13036(.A1(new_n15467_), .A2(pi0625), .B(new_n15472_), .ZN(new_n15473_));
  AOI21_X1   g13037(.A1(new_n15473_), .A2(new_n12841_), .B(new_n15380_), .ZN(new_n15474_));
  AOI21_X1   g13038(.A1(new_n15474_), .A2(new_n13560_), .B(new_n12758_), .ZN(new_n15475_));
  NOR2_X1    g13039(.A1(new_n15467_), .A2(pi0778), .ZN(new_n15476_));
  AOI21_X1   g13040(.A1(new_n15475_), .A2(new_n15471_), .B(new_n15476_), .ZN(new_n15477_));
  NOR2_X1    g13041(.A1(new_n15477_), .A2(pi0785), .ZN(new_n15478_));
  INV_X1     g13042(.I(new_n15478_), .ZN(new_n15479_));
  OAI21_X1   g13043(.A1(new_n15415_), .A2(pi1155), .B(pi0660), .ZN(new_n15480_));
  NOR2_X1    g13044(.A1(new_n15383_), .A2(pi0609), .ZN(new_n15481_));
  NOR2_X1    g13045(.A1(new_n15481_), .A2(new_n12770_), .ZN(new_n15482_));
  NAND2_X1   g13046(.A1(new_n15477_), .A2(pi0609), .ZN(new_n15483_));
  AOI21_X1   g13047(.A1(new_n15483_), .A2(new_n15482_), .B(new_n15480_), .ZN(new_n15484_));
  OAI21_X1   g13048(.A1(new_n15418_), .A2(new_n12770_), .B(new_n13829_), .ZN(new_n15485_));
  OAI21_X1   g13049(.A1(new_n15383_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n15486_));
  AOI21_X1   g13050(.A1(new_n15477_), .A2(new_n12766_), .B(new_n15486_), .ZN(new_n15487_));
  OAI21_X1   g13051(.A1(new_n15487_), .A2(new_n15485_), .B(pi0785), .ZN(new_n15488_));
  OAI21_X1   g13052(.A1(new_n15488_), .A2(new_n15484_), .B(new_n15479_), .ZN(new_n15489_));
  NAND2_X1   g13053(.A1(new_n15489_), .A2(new_n12779_), .ZN(new_n15490_));
  INV_X1     g13054(.I(new_n15490_), .ZN(new_n15491_));
  AOI21_X1   g13055(.A1(new_n15422_), .A2(new_n12785_), .B(new_n12880_), .ZN(new_n15492_));
  AOI21_X1   g13056(.A1(new_n15385_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n15493_));
  OAI21_X1   g13057(.A1(new_n15489_), .A2(new_n12781_), .B(new_n15493_), .ZN(new_n15494_));
  NAND2_X1   g13058(.A1(new_n15494_), .A2(new_n15492_), .ZN(new_n15495_));
  AOI21_X1   g13059(.A1(new_n15425_), .A2(pi1154), .B(pi0627), .ZN(new_n15496_));
  AOI21_X1   g13060(.A1(new_n15385_), .A2(pi0618), .B(pi1154), .ZN(new_n15497_));
  OAI21_X1   g13061(.A1(new_n15489_), .A2(pi0618), .B(new_n15497_), .ZN(new_n15498_));
  AOI21_X1   g13062(.A1(new_n15498_), .A2(new_n15496_), .B(new_n12779_), .ZN(new_n15499_));
  AOI21_X1   g13063(.A1(new_n15499_), .A2(new_n15495_), .B(new_n15491_), .ZN(new_n15500_));
  OR2_X2     g13064(.A1(new_n15500_), .A2(pi0789), .Z(new_n15501_));
  OAI21_X1   g13065(.A1(new_n15429_), .A2(pi1159), .B(pi0648), .ZN(new_n15502_));
  INV_X1     g13066(.I(new_n15387_), .ZN(new_n15503_));
  AOI21_X1   g13067(.A1(new_n15503_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n15504_));
  NAND2_X1   g13068(.A1(new_n15500_), .A2(pi0619), .ZN(new_n15505_));
  AOI21_X1   g13069(.A1(new_n15505_), .A2(new_n15504_), .B(new_n15502_), .ZN(new_n15506_));
  OAI21_X1   g13070(.A1(new_n15432_), .A2(new_n12791_), .B(new_n12895_), .ZN(new_n15507_));
  AOI21_X1   g13071(.A1(new_n15503_), .A2(pi0619), .B(pi1159), .ZN(new_n15508_));
  INV_X1     g13072(.I(new_n15508_), .ZN(new_n15509_));
  AOI21_X1   g13073(.A1(new_n15500_), .A2(new_n12793_), .B(new_n15509_), .ZN(new_n15510_));
  OAI21_X1   g13074(.A1(new_n15510_), .A2(new_n15507_), .B(pi0789), .ZN(new_n15511_));
  OAI21_X1   g13075(.A1(new_n15511_), .A2(new_n15506_), .B(new_n15501_), .ZN(new_n15512_));
  NAND2_X1   g13076(.A1(new_n15512_), .A2(pi0626), .ZN(new_n15513_));
  AOI21_X1   g13077(.A1(new_n15513_), .A2(new_n15448_), .B(new_n15446_), .ZN(new_n15514_));
  OAI21_X1   g13078(.A1(new_n15441_), .A2(new_n12814_), .B(new_n12745_), .ZN(new_n15515_));
  OAI21_X1   g13079(.A1(new_n15389_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n15516_));
  AOI21_X1   g13080(.A1(new_n15512_), .A2(new_n12747_), .B(new_n15516_), .ZN(new_n15517_));
  OAI21_X1   g13081(.A1(new_n15517_), .A2(new_n15515_), .B(pi0788), .ZN(new_n15518_));
  OR2_X2     g13082(.A1(new_n15512_), .A2(pi0788), .Z(new_n15519_));
  OAI21_X1   g13083(.A1(new_n15518_), .A2(new_n15514_), .B(new_n15519_), .ZN(new_n15520_));
  NAND2_X1   g13084(.A1(new_n15520_), .A2(pi0628), .ZN(new_n15521_));
  AOI21_X1   g13085(.A1(new_n15521_), .A2(new_n15445_), .B(new_n15395_), .ZN(new_n15522_));
  NOR2_X1    g13086(.A1(new_n15362_), .A2(pi0628), .ZN(new_n15523_));
  AOI21_X1   g13087(.A1(new_n15391_), .A2(pi0628), .B(new_n15523_), .ZN(new_n15524_));
  OAI21_X1   g13088(.A1(new_n15524_), .A2(new_n12742_), .B(new_n12919_), .ZN(new_n15525_));
  OAI21_X1   g13089(.A1(new_n15443_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n15526_));
  AOI21_X1   g13090(.A1(new_n15520_), .A2(new_n12920_), .B(new_n15526_), .ZN(new_n15527_));
  OAI21_X1   g13091(.A1(new_n15527_), .A2(new_n15525_), .B(pi0792), .ZN(new_n15528_));
  OR2_X2     g13092(.A1(new_n15520_), .A2(pi0792), .Z(new_n15529_));
  OAI21_X1   g13093(.A1(new_n15528_), .A2(new_n15522_), .B(new_n15529_), .ZN(new_n15530_));
  AND2_X2    g13094(.A1(new_n15530_), .A2(new_n12972_), .Z(new_n15531_));
  NOR2_X1    g13095(.A1(new_n15391_), .A2(pi0792), .ZN(new_n15532_));
  OAI21_X1   g13096(.A1(new_n15524_), .A2(new_n12742_), .B(pi0792), .ZN(new_n15533_));
  NOR2_X1    g13097(.A1(new_n15533_), .A2(new_n15394_), .ZN(new_n15534_));
  NOR2_X1    g13098(.A1(new_n15534_), .A2(new_n15532_), .ZN(new_n15535_));
  NAND2_X1   g13099(.A1(new_n15535_), .A2(new_n12741_), .ZN(new_n15536_));
  NAND2_X1   g13100(.A1(new_n15378_), .A2(pi0647), .ZN(new_n15537_));
  AOI21_X1   g13101(.A1(new_n15536_), .A2(new_n15537_), .B(pi1157), .ZN(new_n15538_));
  NOR2_X1    g13102(.A1(new_n15538_), .A2(new_n12981_), .ZN(new_n15539_));
  NAND2_X1   g13103(.A1(new_n15362_), .A2(new_n12943_), .ZN(new_n15540_));
  OAI21_X1   g13104(.A1(new_n15443_), .A2(new_n12943_), .B(new_n15540_), .ZN(new_n15541_));
  AOI21_X1   g13105(.A1(new_n15541_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n15542_));
  OAI21_X1   g13106(.A1(new_n15530_), .A2(new_n12741_), .B(new_n15542_), .ZN(new_n15543_));
  NAND2_X1   g13107(.A1(new_n15543_), .A2(new_n15539_), .ZN(new_n15544_));
  NOR2_X1    g13108(.A1(new_n15362_), .A2(pi0647), .ZN(new_n15545_));
  AOI21_X1   g13109(.A1(new_n15535_), .A2(pi0647), .B(new_n15545_), .ZN(new_n15546_));
  NOR2_X1    g13110(.A1(new_n15546_), .A2(new_n12965_), .ZN(new_n15547_));
  NOR2_X1    g13111(.A1(new_n15547_), .A2(pi0630), .ZN(new_n15548_));
  AOI21_X1   g13112(.A1(new_n15541_), .A2(pi0647), .B(pi1157), .ZN(new_n15549_));
  OAI21_X1   g13113(.A1(new_n15530_), .A2(pi0647), .B(new_n15549_), .ZN(new_n15550_));
  AOI21_X1   g13114(.A1(new_n15550_), .A2(new_n15548_), .B(new_n12972_), .ZN(new_n15551_));
  AOI21_X1   g13115(.A1(new_n15551_), .A2(new_n15544_), .B(new_n15531_), .ZN(new_n15552_));
  OAI21_X1   g13116(.A1(new_n15552_), .A2(pi0790), .B(new_n5477_), .ZN(new_n15553_));
  OAI21_X1   g13117(.A1(new_n15378_), .A2(new_n12975_), .B(pi0715), .ZN(new_n15554_));
  NAND2_X1   g13118(.A1(new_n15378_), .A2(new_n12984_), .ZN(new_n15555_));
  OAI21_X1   g13119(.A1(new_n15541_), .A2(new_n12984_), .B(new_n15555_), .ZN(new_n15556_));
  NOR2_X1    g13120(.A1(new_n15556_), .A2(pi0644), .ZN(new_n15557_));
  OAI21_X1   g13121(.A1(new_n15557_), .A2(new_n15554_), .B(new_n12739_), .ZN(new_n15558_));
  NOR2_X1    g13122(.A1(new_n15547_), .A2(new_n12972_), .ZN(new_n15559_));
  INV_X1     g13123(.I(new_n15559_), .ZN(new_n15560_));
  OAI22_X1   g13124(.A1(new_n15560_), .A2(new_n15538_), .B1(pi0787), .B2(new_n15535_), .ZN(new_n15561_));
  AOI21_X1   g13125(.A1(new_n15561_), .A2(pi0644), .B(pi0715), .ZN(new_n15562_));
  NAND2_X1   g13126(.A1(new_n15552_), .A2(new_n12975_), .ZN(new_n15563_));
  AOI21_X1   g13127(.A1(new_n15563_), .A2(new_n15562_), .B(new_n15558_), .ZN(new_n15564_));
  OAI21_X1   g13128(.A1(new_n15378_), .A2(pi0644), .B(new_n12740_), .ZN(new_n15565_));
  NOR2_X1    g13129(.A1(new_n15556_), .A2(new_n12975_), .ZN(new_n15566_));
  OAI21_X1   g13130(.A1(new_n15566_), .A2(new_n15565_), .B(pi1160), .ZN(new_n15567_));
  NAND2_X1   g13131(.A1(new_n15561_), .A2(new_n12975_), .ZN(new_n15568_));
  NAND2_X1   g13132(.A1(new_n15568_), .A2(pi0715), .ZN(new_n15569_));
  AOI21_X1   g13133(.A1(new_n15552_), .A2(pi0644), .B(new_n15569_), .ZN(new_n15570_));
  OAI21_X1   g13134(.A1(new_n15570_), .A2(new_n15567_), .B(pi0790), .ZN(new_n15571_));
  NOR2_X1    g13135(.A1(new_n15571_), .A2(new_n15564_), .ZN(new_n15572_));
  AOI21_X1   g13136(.A1(new_n6165_), .A2(new_n8058_), .B(pi0057), .ZN(new_n15573_));
  OAI21_X1   g13137(.A1(new_n15572_), .A2(new_n15553_), .B(new_n15573_), .ZN(new_n15574_));
  AOI21_X1   g13138(.A1(new_n15574_), .A2(new_n15361_), .B(new_n15360_), .ZN(po0301));
  INV_X1     g13139(.I(new_n12980_), .ZN(new_n15576_));
  INV_X1     g13140(.I(pi0698), .ZN(new_n15577_));
  NOR2_X1    g13141(.A1(new_n3042_), .A2(pi0145), .ZN(new_n15578_));
  AOI21_X1   g13142(.A1(new_n12826_), .A2(new_n15577_), .B(new_n15578_), .ZN(new_n15579_));
  NOR2_X1    g13143(.A1(new_n15579_), .A2(pi0778), .ZN(new_n15580_));
  NOR2_X1    g13144(.A1(new_n15578_), .A2(pi1153), .ZN(new_n15581_));
  NOR2_X1    g13145(.A1(new_n12834_), .A2(pi0698), .ZN(new_n15582_));
  INV_X1     g13146(.I(new_n15582_), .ZN(new_n15583_));
  NAND2_X1   g13147(.A1(new_n15583_), .A2(new_n15581_), .ZN(new_n15584_));
  INV_X1     g13148(.I(new_n15584_), .ZN(new_n15585_));
  NOR2_X1    g13149(.A1(new_n15582_), .A2(new_n15579_), .ZN(new_n15586_));
  NOR2_X1    g13150(.A1(new_n15586_), .A2(new_n12841_), .ZN(new_n15587_));
  NOR3_X1    g13151(.A1(new_n15585_), .A2(new_n12758_), .A3(new_n15587_), .ZN(new_n15588_));
  NOR2_X1    g13152(.A1(new_n15588_), .A2(new_n15580_), .ZN(new_n15589_));
  NOR2_X1    g13153(.A1(new_n15589_), .A2(new_n12871_), .ZN(new_n15590_));
  INV_X1     g13154(.I(new_n15590_), .ZN(new_n15591_));
  NOR2_X1    g13155(.A1(new_n15591_), .A2(new_n12889_), .ZN(new_n15592_));
  INV_X1     g13156(.I(new_n15592_), .ZN(new_n15593_));
  NOR2_X1    g13157(.A1(new_n15593_), .A2(new_n12924_), .ZN(new_n15594_));
  INV_X1     g13158(.I(new_n15594_), .ZN(new_n15595_));
  NOR2_X1    g13159(.A1(new_n15595_), .A2(new_n12953_), .ZN(new_n15596_));
  INV_X1     g13160(.I(new_n15596_), .ZN(new_n15597_));
  NAND2_X1   g13161(.A1(new_n15597_), .A2(new_n12741_), .ZN(new_n15598_));
  INV_X1     g13162(.I(new_n15578_), .ZN(new_n15599_));
  NAND2_X1   g13163(.A1(new_n15599_), .A2(pi0647), .ZN(new_n15600_));
  AOI21_X1   g13164(.A1(new_n15598_), .A2(new_n15600_), .B(pi1157), .ZN(new_n15601_));
  INV_X1     g13165(.I(new_n15601_), .ZN(new_n15602_));
  NAND2_X1   g13166(.A1(new_n15578_), .A2(new_n12741_), .ZN(new_n15603_));
  OAI21_X1   g13167(.A1(new_n15597_), .A2(new_n12741_), .B(new_n15603_), .ZN(new_n15604_));
  OAI22_X1   g13168(.A1(new_n15602_), .A2(new_n12981_), .B1(new_n15576_), .B2(new_n15604_), .ZN(new_n15605_));
  INV_X1     g13169(.I(new_n14298_), .ZN(new_n15606_));
  NAND2_X1   g13170(.A1(new_n14297_), .A2(pi0630), .ZN(new_n15607_));
  OAI21_X1   g13171(.A1(pi0630), .A2(new_n15606_), .B(new_n15607_), .ZN(new_n15608_));
  INV_X1     g13172(.I(new_n12749_), .ZN(new_n15609_));
  NOR2_X1    g13173(.A1(new_n13340_), .A2(pi0767), .ZN(new_n15610_));
  NOR2_X1    g13174(.A1(new_n15610_), .A2(new_n15578_), .ZN(new_n15611_));
  NOR3_X1    g13175(.A1(new_n15611_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n15612_));
  NOR2_X1    g13176(.A1(new_n15611_), .A2(new_n12762_), .ZN(new_n15613_));
  AOI21_X1   g13177(.A1(new_n15613_), .A2(new_n12768_), .B(pi1155), .ZN(new_n15614_));
  INV_X1     g13178(.I(new_n15611_), .ZN(new_n15615_));
  AOI21_X1   g13179(.A1(new_n15615_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n15616_));
  NOR3_X1    g13180(.A1(new_n15614_), .A2(new_n15616_), .A3(new_n12764_), .ZN(new_n15617_));
  NOR2_X1    g13181(.A1(new_n15617_), .A2(new_n15612_), .ZN(new_n15618_));
  INV_X1     g13182(.I(new_n15618_), .ZN(new_n15619_));
  AOI21_X1   g13183(.A1(new_n15619_), .A2(new_n12783_), .B(pi1154), .ZN(new_n15620_));
  AOI21_X1   g13184(.A1(new_n15619_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n15621_));
  NOR3_X1    g13185(.A1(new_n15620_), .A2(new_n15621_), .A3(new_n12779_), .ZN(new_n15622_));
  AOI21_X1   g13186(.A1(new_n12779_), .A2(new_n15619_), .B(new_n15622_), .ZN(new_n15623_));
  NOR2_X1    g13187(.A1(new_n15623_), .A2(pi0789), .ZN(new_n15624_));
  NAND2_X1   g13188(.A1(new_n15623_), .A2(new_n12793_), .ZN(new_n15625_));
  NAND2_X1   g13189(.A1(new_n15599_), .A2(pi0619), .ZN(new_n15626_));
  AOI21_X1   g13190(.A1(new_n15625_), .A2(new_n15626_), .B(pi1159), .ZN(new_n15627_));
  NAND2_X1   g13191(.A1(new_n15623_), .A2(pi0619), .ZN(new_n15628_));
  NAND2_X1   g13192(.A1(new_n15599_), .A2(new_n12793_), .ZN(new_n15629_));
  AOI21_X1   g13193(.A1(new_n15628_), .A2(new_n15629_), .B(new_n12791_), .ZN(new_n15630_));
  NOR3_X1    g13194(.A1(new_n15627_), .A2(new_n15630_), .A3(new_n12796_), .ZN(new_n15631_));
  NOR2_X1    g13195(.A1(new_n15631_), .A2(new_n15624_), .ZN(new_n15632_));
  NOR2_X1    g13196(.A1(new_n15632_), .A2(new_n12803_), .ZN(new_n15633_));
  AOI21_X1   g13197(.A1(new_n15609_), .A2(new_n15578_), .B(new_n15633_), .ZN(new_n15634_));
  NOR2_X1    g13198(.A1(new_n15634_), .A2(new_n12808_), .ZN(new_n15635_));
  NOR2_X1    g13199(.A1(new_n15632_), .A2(pi0788), .ZN(new_n15636_));
  NOR2_X1    g13200(.A1(new_n15635_), .A2(new_n15636_), .ZN(new_n15637_));
  NAND2_X1   g13201(.A1(new_n15637_), .A2(new_n13384_), .ZN(new_n15638_));
  OAI21_X1   g13202(.A1(new_n13384_), .A2(new_n15578_), .B(new_n15638_), .ZN(new_n15639_));
  AOI21_X1   g13203(.A1(new_n15639_), .A2(new_n15608_), .B(new_n15605_), .ZN(new_n15640_));
  NOR2_X1    g13204(.A1(new_n15579_), .A2(new_n12754_), .ZN(new_n15641_));
  NOR2_X1    g13205(.A1(new_n15615_), .A2(new_n15641_), .ZN(new_n15642_));
  NAND2_X1   g13206(.A1(new_n15642_), .A2(new_n12758_), .ZN(new_n15643_));
  NAND2_X1   g13207(.A1(new_n15641_), .A2(pi0625), .ZN(new_n15644_));
  NAND3_X1   g13208(.A1(new_n15644_), .A2(pi1153), .A3(new_n15611_), .ZN(new_n15645_));
  AND3_X2    g13209(.A1(new_n15645_), .A2(pi0608), .A3(new_n15584_), .Z(new_n15646_));
  NOR2_X1    g13210(.A1(new_n15587_), .A2(pi0608), .ZN(new_n15647_));
  INV_X1     g13211(.I(new_n15644_), .ZN(new_n15648_));
  OAI21_X1   g13212(.A1(new_n15642_), .A2(new_n15648_), .B(new_n15581_), .ZN(new_n15649_));
  NAND2_X1   g13213(.A1(new_n15647_), .A2(new_n15649_), .ZN(new_n15650_));
  NAND2_X1   g13214(.A1(new_n15650_), .A2(pi0778), .ZN(new_n15651_));
  OAI21_X1   g13215(.A1(new_n15651_), .A2(new_n15646_), .B(new_n15643_), .ZN(new_n15652_));
  INV_X1     g13216(.I(new_n15652_), .ZN(new_n15653_));
  INV_X1     g13217(.I(new_n15589_), .ZN(new_n15654_));
  NOR2_X1    g13218(.A1(new_n15654_), .A2(pi0609), .ZN(new_n15655_));
  AOI21_X1   g13219(.A1(new_n15652_), .A2(pi0609), .B(new_n15655_), .ZN(new_n15656_));
  NOR2_X1    g13220(.A1(new_n15656_), .A2(new_n12770_), .ZN(new_n15657_));
  NOR2_X1    g13221(.A1(new_n15657_), .A2(new_n15614_), .ZN(new_n15658_));
  NOR2_X1    g13222(.A1(new_n15653_), .A2(pi0609), .ZN(new_n15659_));
  NOR2_X1    g13223(.A1(new_n15654_), .A2(new_n12766_), .ZN(new_n15660_));
  OAI21_X1   g13224(.A1(new_n15659_), .A2(new_n15660_), .B(new_n12770_), .ZN(new_n15661_));
  NOR2_X1    g13225(.A1(new_n15616_), .A2(pi0660), .ZN(new_n15662_));
  AOI22_X1   g13226(.A1(new_n15658_), .A2(pi0660), .B1(new_n15661_), .B2(new_n15662_), .ZN(new_n15663_));
  NAND2_X1   g13227(.A1(new_n15663_), .A2(pi0785), .ZN(new_n15664_));
  OAI21_X1   g13228(.A1(pi0785), .A2(new_n15653_), .B(new_n15664_), .ZN(new_n15665_));
  INV_X1     g13229(.I(new_n15665_), .ZN(new_n15666_));
  NAND2_X1   g13230(.A1(new_n15591_), .A2(pi0618), .ZN(new_n15667_));
  OAI21_X1   g13231(.A1(new_n15666_), .A2(pi0618), .B(new_n15667_), .ZN(new_n15668_));
  AOI21_X1   g13232(.A1(new_n15668_), .A2(new_n12785_), .B(new_n15621_), .ZN(new_n15669_));
  NOR2_X1    g13233(.A1(new_n15590_), .A2(pi0618), .ZN(new_n15670_));
  NOR2_X1    g13234(.A1(new_n15666_), .A2(new_n12781_), .ZN(new_n15671_));
  OAI21_X1   g13235(.A1(new_n15671_), .A2(new_n15670_), .B(pi1154), .ZN(new_n15672_));
  NOR2_X1    g13236(.A1(new_n15620_), .A2(new_n12880_), .ZN(new_n15673_));
  AOI22_X1   g13237(.A1(new_n15669_), .A2(new_n12880_), .B1(new_n15672_), .B2(new_n15673_), .ZN(new_n15674_));
  NAND2_X1   g13238(.A1(new_n15674_), .A2(pi0781), .ZN(new_n15675_));
  OAI21_X1   g13239(.A1(pi0781), .A2(new_n15666_), .B(new_n15675_), .ZN(new_n15676_));
  AOI21_X1   g13240(.A1(new_n15676_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n15677_));
  NAND2_X1   g13241(.A1(new_n15593_), .A2(new_n12793_), .ZN(new_n15678_));
  NAND2_X1   g13242(.A1(new_n15676_), .A2(pi0619), .ZN(new_n15679_));
  AOI21_X1   g13243(.A1(new_n15679_), .A2(new_n15678_), .B(new_n12791_), .ZN(new_n15680_));
  NOR3_X1    g13244(.A1(new_n15680_), .A2(new_n12895_), .A3(new_n15627_), .ZN(new_n15681_));
  INV_X1     g13245(.I(new_n15630_), .ZN(new_n15682_));
  NOR2_X1    g13246(.A1(new_n15592_), .A2(new_n12793_), .ZN(new_n15683_));
  AOI21_X1   g13247(.A1(new_n15676_), .A2(new_n12793_), .B(new_n15683_), .ZN(new_n15684_));
  OAI21_X1   g13248(.A1(new_n15684_), .A2(pi1159), .B(new_n15682_), .ZN(new_n15685_));
  OAI21_X1   g13249(.A1(new_n15685_), .A2(pi0648), .B(pi0789), .ZN(new_n15686_));
  OAI21_X1   g13250(.A1(new_n15686_), .A2(new_n15681_), .B(new_n15677_), .ZN(new_n15687_));
  INV_X1     g13251(.I(new_n12913_), .ZN(new_n15688_));
  INV_X1     g13252(.I(new_n12914_), .ZN(new_n15689_));
  OAI22_X1   g13253(.A1(new_n15634_), .A2(new_n15689_), .B1(new_n15688_), .B2(new_n15593_), .ZN(new_n15690_));
  NAND2_X1   g13254(.A1(new_n15690_), .A2(pi0788), .ZN(new_n15691_));
  AOI21_X1   g13255(.A1(new_n15687_), .A2(new_n15691_), .B(new_n15340_), .ZN(new_n15692_));
  INV_X1     g13256(.I(new_n15341_), .ZN(new_n15693_));
  INV_X1     g13257(.I(new_n12949_), .ZN(new_n15694_));
  NOR2_X1    g13258(.A1(new_n12931_), .A2(new_n12742_), .ZN(new_n15695_));
  INV_X1     g13259(.I(new_n15695_), .ZN(new_n15696_));
  OAI22_X1   g13260(.A1(new_n15637_), .A2(new_n15694_), .B1(new_n15595_), .B2(new_n15696_), .ZN(new_n15697_));
  NAND2_X1   g13261(.A1(new_n15697_), .A2(new_n12919_), .ZN(new_n15698_));
  INV_X1     g13262(.I(new_n12948_), .ZN(new_n15699_));
  NOR2_X1    g13263(.A1(new_n12921_), .A2(pi1156), .ZN(new_n15700_));
  INV_X1     g13264(.I(new_n15700_), .ZN(new_n15701_));
  OAI22_X1   g13265(.A1(new_n15637_), .A2(new_n15699_), .B1(new_n15595_), .B2(new_n15701_), .ZN(new_n15702_));
  NAND2_X1   g13266(.A1(new_n15702_), .A2(pi0629), .ZN(new_n15703_));
  NAND2_X1   g13267(.A1(new_n15698_), .A2(new_n15703_), .ZN(new_n15704_));
  NAND2_X1   g13268(.A1(new_n15704_), .A2(pi0792), .ZN(new_n15705_));
  NAND2_X1   g13269(.A1(new_n15705_), .A2(new_n15693_), .ZN(new_n15706_));
  OAI22_X1   g13270(.A1(new_n15692_), .A2(new_n15706_), .B1(new_n12972_), .B2(new_n15640_), .ZN(new_n15707_));
  NAND2_X1   g13271(.A1(new_n15707_), .A2(new_n13000_), .ZN(new_n15708_));
  AND2_X2    g13272(.A1(new_n15707_), .A2(new_n12975_), .Z(new_n15709_));
  OAI21_X1   g13273(.A1(new_n15604_), .A2(new_n12965_), .B(new_n15602_), .ZN(new_n15710_));
  NAND2_X1   g13274(.A1(new_n15596_), .A2(new_n12972_), .ZN(new_n15711_));
  OAI21_X1   g13275(.A1(new_n15710_), .A2(new_n12972_), .B(new_n15711_), .ZN(new_n15712_));
  NOR2_X1    g13276(.A1(new_n15712_), .A2(new_n12975_), .ZN(new_n15713_));
  OAI21_X1   g13277(.A1(new_n15709_), .A2(new_n15713_), .B(new_n12740_), .ZN(new_n15714_));
  NOR2_X1    g13278(.A1(new_n15578_), .A2(new_n12975_), .ZN(new_n15715_));
  NOR2_X1    g13279(.A1(new_n12985_), .A2(new_n15578_), .ZN(new_n15716_));
  AOI21_X1   g13280(.A1(new_n15639_), .A2(new_n12985_), .B(new_n15716_), .ZN(new_n15717_));
  NOR2_X1    g13281(.A1(new_n15717_), .A2(pi0644), .ZN(new_n15718_));
  OAI21_X1   g13282(.A1(new_n15718_), .A2(new_n15715_), .B(pi0715), .ZN(new_n15719_));
  NAND3_X1   g13283(.A1(new_n15714_), .A2(new_n12739_), .A3(new_n15719_), .ZN(new_n15720_));
  NOR2_X1    g13284(.A1(new_n15712_), .A2(pi0644), .ZN(new_n15721_));
  AOI21_X1   g13285(.A1(new_n15707_), .A2(pi0644), .B(new_n15721_), .ZN(new_n15722_));
  NAND2_X1   g13286(.A1(new_n15599_), .A2(new_n12975_), .ZN(new_n15723_));
  OAI21_X1   g13287(.A1(new_n15717_), .A2(new_n12975_), .B(new_n15723_), .ZN(new_n15724_));
  AOI21_X1   g13288(.A1(new_n15724_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n15725_));
  OAI21_X1   g13289(.A1(new_n15722_), .A2(new_n12740_), .B(new_n15725_), .ZN(new_n15726_));
  NAND3_X1   g13290(.A1(new_n15720_), .A2(pi0790), .A3(new_n15726_), .ZN(new_n15727_));
  NAND2_X1   g13291(.A1(new_n15727_), .A2(new_n15708_), .ZN(new_n15728_));
  AOI21_X1   g13292(.A1(po1038), .A2(new_n5656_), .B(pi0832), .ZN(new_n15729_));
  INV_X1     g13293(.I(new_n12982_), .ZN(new_n15730_));
  NAND2_X1   g13294(.A1(new_n13192_), .A2(new_n5656_), .ZN(new_n15731_));
  NOR2_X1    g13295(.A1(new_n15731_), .A2(new_n12870_), .ZN(new_n15732_));
  INV_X1     g13296(.I(new_n15732_), .ZN(new_n15733_));
  INV_X1     g13297(.I(new_n15731_), .ZN(new_n15734_));
  NOR2_X1    g13298(.A1(new_n13344_), .A2(pi0145), .ZN(new_n15735_));
  OAI21_X1   g13299(.A1(new_n14125_), .A2(new_n15735_), .B(new_n15577_), .ZN(new_n15736_));
  OAI21_X1   g13300(.A1(new_n14122_), .A2(new_n5656_), .B(new_n3265_), .ZN(new_n15737_));
  NAND2_X1   g13301(.A1(new_n15737_), .A2(new_n2609_), .ZN(new_n15738_));
  INV_X1     g13302(.I(new_n13501_), .ZN(new_n15739_));
  AOI21_X1   g13303(.A1(new_n15739_), .A2(new_n13476_), .B(pi0299), .ZN(new_n15740_));
  INV_X1     g13304(.I(new_n13513_), .ZN(new_n15741_));
  AOI21_X1   g13305(.A1(new_n15741_), .A2(new_n13506_), .B(new_n2628_), .ZN(new_n15742_));
  NOR2_X1    g13306(.A1(new_n15740_), .A2(new_n15742_), .ZN(new_n15743_));
  AOI21_X1   g13307(.A1(new_n15743_), .A2(pi0039), .B(new_n14115_), .ZN(new_n15744_));
  NAND2_X1   g13308(.A1(new_n15744_), .A2(new_n5656_), .ZN(new_n15745_));
  AOI21_X1   g13309(.A1(new_n15745_), .A2(new_n15738_), .B(new_n15736_), .ZN(new_n15746_));
  NAND2_X1   g13310(.A1(new_n2609_), .A2(new_n15577_), .ZN(new_n15747_));
  AOI21_X1   g13311(.A1(new_n15734_), .A2(new_n15747_), .B(new_n15746_), .ZN(new_n15748_));
  NAND2_X1   g13312(.A1(new_n15748_), .A2(new_n13521_), .ZN(new_n15749_));
  NOR2_X1    g13313(.A1(new_n15734_), .A2(new_n13521_), .ZN(new_n15750_));
  INV_X1     g13314(.I(new_n15750_), .ZN(new_n15751_));
  AOI21_X1   g13315(.A1(new_n15749_), .A2(new_n15751_), .B(pi1153), .ZN(new_n15752_));
  NAND2_X1   g13316(.A1(new_n15731_), .A2(new_n13521_), .ZN(new_n15753_));
  NAND2_X1   g13317(.A1(new_n15748_), .A2(pi0625), .ZN(new_n15754_));
  AOI21_X1   g13318(.A1(new_n15754_), .A2(new_n15753_), .B(new_n12841_), .ZN(new_n15755_));
  NOR3_X1    g13319(.A1(new_n15752_), .A2(new_n15755_), .A3(new_n12758_), .ZN(new_n15756_));
  NOR2_X1    g13320(.A1(new_n15748_), .A2(pi0778), .ZN(new_n15757_));
  NOR2_X1    g13321(.A1(new_n15756_), .A2(new_n15757_), .ZN(new_n15758_));
  OAI21_X1   g13322(.A1(new_n15758_), .A2(new_n12869_), .B(new_n15733_), .ZN(new_n15759_));
  INV_X1     g13323(.I(new_n15759_), .ZN(new_n15760_));
  NOR2_X1    g13324(.A1(new_n15734_), .A2(new_n12888_), .ZN(new_n15761_));
  AOI21_X1   g13325(.A1(new_n15760_), .A2(new_n12888_), .B(new_n15761_), .ZN(new_n15762_));
  NOR2_X1    g13326(.A1(new_n15762_), .A2(new_n14288_), .ZN(new_n15763_));
  AOI21_X1   g13327(.A1(new_n14288_), .A2(new_n15731_), .B(new_n15763_), .ZN(new_n15764_));
  NOR2_X1    g13328(.A1(new_n15764_), .A2(pi0628), .ZN(new_n15765_));
  NOR2_X1    g13329(.A1(new_n15734_), .A2(new_n12920_), .ZN(new_n15766_));
  OAI21_X1   g13330(.A1(new_n15765_), .A2(new_n15766_), .B(new_n12742_), .ZN(new_n15767_));
  NOR2_X1    g13331(.A1(new_n15734_), .A2(pi0628), .ZN(new_n15768_));
  NOR2_X1    g13332(.A1(new_n15764_), .A2(new_n12920_), .ZN(new_n15769_));
  OAI21_X1   g13333(.A1(new_n15769_), .A2(new_n15768_), .B(pi1156), .ZN(new_n15770_));
  NAND3_X1   g13334(.A1(new_n15767_), .A2(new_n15770_), .A3(pi0792), .ZN(new_n15771_));
  NAND2_X1   g13335(.A1(new_n15764_), .A2(new_n12937_), .ZN(new_n15772_));
  NAND2_X1   g13336(.A1(new_n15771_), .A2(new_n15772_), .ZN(new_n15773_));
  NAND2_X1   g13337(.A1(new_n15773_), .A2(pi0647), .ZN(new_n15774_));
  OAI21_X1   g13338(.A1(pi0647), .A2(new_n15731_), .B(new_n15774_), .ZN(new_n15775_));
  NAND2_X1   g13339(.A1(new_n15773_), .A2(new_n12741_), .ZN(new_n15776_));
  OAI21_X1   g13340(.A1(new_n12741_), .A2(new_n15731_), .B(new_n15776_), .ZN(new_n15777_));
  OAI22_X1   g13341(.A1(new_n15576_), .A2(new_n15775_), .B1(new_n15777_), .B2(new_n15730_), .ZN(new_n15778_));
  INV_X1     g13342(.I(new_n15244_), .ZN(new_n15779_));
  NOR2_X1    g13343(.A1(new_n2609_), .A2(new_n5656_), .ZN(new_n15780_));
  INV_X1     g13344(.I(new_n15735_), .ZN(new_n15781_));
  INV_X1     g13345(.I(pi0767), .ZN(new_n15782_));
  AOI21_X1   g13346(.A1(new_n13341_), .A2(new_n15782_), .B(new_n3265_), .ZN(new_n15783_));
  INV_X1     g13347(.I(new_n13245_), .ZN(new_n15784_));
  NOR2_X1    g13348(.A1(new_n13334_), .A2(pi0145), .ZN(new_n15785_));
  AOI22_X1   g13349(.A1(new_n15785_), .A2(new_n15782_), .B1(pi0145), .B2(new_n15784_), .ZN(new_n15786_));
  NAND2_X1   g13350(.A1(new_n13337_), .A2(new_n13336_), .ZN(new_n15787_));
  OAI21_X1   g13351(.A1(new_n15787_), .A2(pi0145), .B(pi0767), .ZN(new_n15788_));
  NAND2_X1   g13352(.A1(new_n15786_), .A2(new_n15788_), .ZN(new_n15789_));
  AOI22_X1   g13353(.A1(new_n15789_), .A2(new_n3265_), .B1(new_n15781_), .B2(new_n15783_), .ZN(new_n15790_));
  NOR2_X1    g13354(.A1(new_n15790_), .A2(new_n2610_), .ZN(new_n15791_));
  NOR2_X1    g13355(.A1(new_n15791_), .A2(new_n15780_), .ZN(new_n15792_));
  NOR2_X1    g13356(.A1(new_n15792_), .A2(new_n12760_), .ZN(new_n15793_));
  AOI21_X1   g13357(.A1(new_n12760_), .A2(new_n15731_), .B(new_n15793_), .ZN(new_n15794_));
  INV_X1     g13358(.I(new_n15793_), .ZN(new_n15795_));
  OAI22_X1   g13359(.A1(new_n15795_), .A2(pi0609), .B1(new_n13353_), .B2(new_n15734_), .ZN(new_n15796_));
  NAND2_X1   g13360(.A1(new_n15796_), .A2(new_n12770_), .ZN(new_n15797_));
  OAI22_X1   g13361(.A1(new_n15795_), .A2(new_n12766_), .B1(new_n12772_), .B2(new_n15734_), .ZN(new_n15798_));
  AOI21_X1   g13362(.A1(new_n15798_), .A2(pi1155), .B(new_n12764_), .ZN(new_n15799_));
  AOI22_X1   g13363(.A1(new_n15799_), .A2(new_n15797_), .B1(new_n12764_), .B2(new_n15794_), .ZN(new_n15800_));
  NOR2_X1    g13364(.A1(new_n12781_), .A2(new_n12785_), .ZN(new_n15801_));
  NOR2_X1    g13365(.A1(pi0618), .A2(pi1154), .ZN(new_n15802_));
  NOR3_X1    g13366(.A1(new_n15801_), .A2(new_n12779_), .A3(new_n15802_), .ZN(new_n15803_));
  INV_X1     g13367(.I(new_n15238_), .ZN(new_n15804_));
  NAND2_X1   g13368(.A1(new_n15734_), .A2(new_n15804_), .ZN(new_n15805_));
  OAI22_X1   g13369(.A1(new_n15800_), .A2(new_n15803_), .B1(new_n12779_), .B2(new_n15805_), .ZN(new_n15806_));
  XNOR2_X1   g13370(.A1(pi0619), .A2(pi1159), .ZN(new_n15807_));
  NOR2_X1    g13371(.A1(new_n15731_), .A2(new_n15807_), .ZN(new_n15808_));
  AOI22_X1   g13372(.A1(new_n15806_), .A2(new_n15779_), .B1(pi0789), .B2(new_n15808_), .ZN(new_n15809_));
  OAI22_X1   g13373(.A1(new_n15809_), .A2(new_n12803_), .B1(new_n12749_), .B2(new_n15731_), .ZN(new_n15810_));
  NAND2_X1   g13374(.A1(new_n15810_), .A2(pi0788), .ZN(new_n15811_));
  OAI21_X1   g13375(.A1(pi0788), .A2(new_n15809_), .B(new_n15811_), .ZN(new_n15812_));
  NOR2_X1    g13376(.A1(new_n15812_), .A2(new_n12943_), .ZN(new_n15813_));
  AOI21_X1   g13377(.A1(new_n12943_), .A2(new_n15731_), .B(new_n15813_), .ZN(new_n15814_));
  INV_X1     g13378(.I(new_n15814_), .ZN(new_n15815_));
  AOI21_X1   g13379(.A1(new_n15608_), .A2(new_n15815_), .B(new_n15778_), .ZN(new_n15816_));
  AND2_X2    g13380(.A1(new_n15770_), .A2(new_n12919_), .Z(new_n15817_));
  AOI21_X1   g13381(.A1(pi0629), .A2(new_n15767_), .B(new_n15817_), .ZN(new_n15818_));
  NOR3_X1    g13382(.A1(new_n12919_), .A2(new_n12742_), .A3(pi0628), .ZN(new_n15819_));
  NOR3_X1    g13383(.A1(new_n12920_), .A2(pi0629), .A3(pi1156), .ZN(new_n15820_));
  NOR2_X1    g13384(.A1(new_n15819_), .A2(new_n15820_), .ZN(new_n15821_));
  NOR2_X1    g13385(.A1(new_n15812_), .A2(new_n15821_), .ZN(new_n15822_));
  OAI21_X1   g13386(.A1(new_n15818_), .A2(new_n15822_), .B(pi0792), .ZN(new_n15823_));
  INV_X1     g13387(.I(new_n15340_), .ZN(new_n15824_));
  INV_X1     g13388(.I(new_n15780_), .ZN(new_n15825_));
  INV_X1     g13389(.I(new_n15124_), .ZN(new_n15826_));
  AOI21_X1   g13390(.A1(new_n15782_), .A2(new_n13566_), .B(new_n15826_), .ZN(new_n15827_));
  NOR2_X1    g13391(.A1(new_n13562_), .A2(new_n15610_), .ZN(new_n15828_));
  NOR2_X1    g13392(.A1(new_n15828_), .A2(new_n5656_), .ZN(new_n15829_));
  AOI21_X1   g13393(.A1(new_n15829_), .A2(new_n5336_), .B(new_n3265_), .ZN(new_n15830_));
  OAI21_X1   g13394(.A1(new_n15827_), .A2(pi0145), .B(new_n15830_), .ZN(new_n15831_));
  NAND2_X1   g13395(.A1(new_n14172_), .A2(pi0145), .ZN(new_n15832_));
  NAND2_X1   g13396(.A1(new_n14174_), .A2(new_n5656_), .ZN(new_n15833_));
  AOI21_X1   g13397(.A1(new_n15832_), .A2(new_n15833_), .B(pi0767), .ZN(new_n15834_));
  NAND2_X1   g13398(.A1(new_n13805_), .A2(new_n13807_), .ZN(new_n15835_));
  NAND2_X1   g13399(.A1(new_n15835_), .A2(pi0145), .ZN(new_n15836_));
  NAND2_X1   g13400(.A1(new_n14177_), .A2(new_n5656_), .ZN(new_n15837_));
  AOI21_X1   g13401(.A1(new_n15837_), .A2(new_n15836_), .B(new_n15782_), .ZN(new_n15838_));
  OAI21_X1   g13402(.A1(new_n15838_), .A2(new_n15834_), .B(new_n2627_), .ZN(new_n15839_));
  NOR2_X1    g13403(.A1(new_n14182_), .A2(pi0145), .ZN(new_n15840_));
  NOR2_X1    g13404(.A1(new_n14184_), .A2(new_n5656_), .ZN(new_n15841_));
  OAI21_X1   g13405(.A1(new_n15840_), .A2(new_n15841_), .B(pi0767), .ZN(new_n15842_));
  NOR2_X1    g13406(.A1(new_n14187_), .A2(new_n5656_), .ZN(new_n15843_));
  NOR2_X1    g13407(.A1(new_n14189_), .A2(pi0145), .ZN(new_n15844_));
  OAI21_X1   g13408(.A1(new_n15843_), .A2(new_n15844_), .B(new_n15782_), .ZN(new_n15845_));
  NAND3_X1   g13409(.A1(new_n15845_), .A2(new_n15842_), .A3(pi0039), .ZN(new_n15846_));
  NAND3_X1   g13410(.A1(new_n15846_), .A2(new_n3265_), .A3(new_n15839_), .ZN(new_n15847_));
  NAND3_X1   g13411(.A1(new_n15847_), .A2(new_n15577_), .A3(new_n15831_), .ZN(new_n15848_));
  NAND2_X1   g13412(.A1(new_n15790_), .A2(pi0698), .ZN(new_n15849_));
  NAND3_X1   g13413(.A1(new_n15849_), .A2(new_n15848_), .A3(new_n2609_), .ZN(new_n15850_));
  NAND2_X1   g13414(.A1(new_n15850_), .A2(new_n15825_), .ZN(new_n15851_));
  NAND2_X1   g13415(.A1(new_n15851_), .A2(new_n12758_), .ZN(new_n15852_));
  INV_X1     g13416(.I(new_n15755_), .ZN(new_n15853_));
  NOR2_X1    g13417(.A1(new_n15792_), .A2(new_n13521_), .ZN(new_n15854_));
  AOI21_X1   g13418(.A1(new_n15851_), .A2(new_n13521_), .B(new_n15854_), .ZN(new_n15855_));
  OAI21_X1   g13419(.A1(new_n15855_), .A2(pi1153), .B(new_n15853_), .ZN(new_n15856_));
  NOR2_X1    g13420(.A1(new_n15792_), .A2(pi0625), .ZN(new_n15857_));
  AOI21_X1   g13421(.A1(new_n15851_), .A2(pi0625), .B(new_n15857_), .ZN(new_n15858_));
  OAI21_X1   g13422(.A1(new_n15858_), .A2(new_n12841_), .B(pi0608), .ZN(new_n15859_));
  OAI22_X1   g13423(.A1(pi0608), .A2(new_n15856_), .B1(new_n15859_), .B2(new_n15752_), .ZN(new_n15860_));
  OAI21_X1   g13424(.A1(new_n15860_), .A2(new_n12758_), .B(new_n15852_), .ZN(new_n15861_));
  INV_X1     g13425(.I(new_n15861_), .ZN(new_n15862_));
  INV_X1     g13426(.I(new_n15758_), .ZN(new_n15863_));
  NOR2_X1    g13427(.A1(new_n15863_), .A2(pi0609), .ZN(new_n15864_));
  INV_X1     g13428(.I(new_n15864_), .ZN(new_n15865_));
  NAND2_X1   g13429(.A1(new_n15861_), .A2(pi0609), .ZN(new_n15866_));
  NAND2_X1   g13430(.A1(new_n15866_), .A2(new_n15865_), .ZN(new_n15867_));
  NAND2_X1   g13431(.A1(new_n15867_), .A2(pi1155), .ZN(new_n15868_));
  NAND3_X1   g13432(.A1(new_n15868_), .A2(pi0660), .A3(new_n15797_), .ZN(new_n15869_));
  NAND2_X1   g13433(.A1(new_n15798_), .A2(pi1155), .ZN(new_n15870_));
  NOR2_X1    g13434(.A1(new_n15862_), .A2(pi0609), .ZN(new_n15871_));
  NOR2_X1    g13435(.A1(new_n15863_), .A2(new_n12766_), .ZN(new_n15872_));
  OAI21_X1   g13436(.A1(new_n15871_), .A2(new_n15872_), .B(new_n12770_), .ZN(new_n15873_));
  NAND3_X1   g13437(.A1(new_n15873_), .A2(new_n13829_), .A3(new_n15870_), .ZN(new_n15874_));
  NAND3_X1   g13438(.A1(new_n15874_), .A2(new_n15869_), .A3(pi0785), .ZN(new_n15875_));
  OAI21_X1   g13439(.A1(pi0785), .A2(new_n15862_), .B(new_n15875_), .ZN(new_n15876_));
  AOI21_X1   g13440(.A1(new_n15734_), .A2(pi0618), .B(pi1154), .ZN(new_n15877_));
  OAI21_X1   g13441(.A1(new_n15800_), .A2(pi0618), .B(new_n15877_), .ZN(new_n15878_));
  AND2_X2    g13442(.A1(new_n15878_), .A2(pi0627), .Z(new_n15879_));
  OAI21_X1   g13443(.A1(new_n15760_), .A2(pi0618), .B(pi1154), .ZN(new_n15880_));
  NOR2_X1    g13444(.A1(new_n15876_), .A2(new_n12781_), .ZN(new_n15881_));
  OAI21_X1   g13445(.A1(new_n15881_), .A2(new_n15880_), .B(new_n15879_), .ZN(new_n15882_));
  AOI21_X1   g13446(.A1(new_n15734_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n15883_));
  OAI21_X1   g13447(.A1(new_n15800_), .A2(new_n12781_), .B(new_n15883_), .ZN(new_n15884_));
  AND2_X2    g13448(.A1(new_n15884_), .A2(new_n12880_), .Z(new_n15885_));
  AOI21_X1   g13449(.A1(new_n15759_), .A2(pi0618), .B(pi1154), .ZN(new_n15886_));
  OAI21_X1   g13450(.A1(new_n15876_), .A2(pi0618), .B(new_n15886_), .ZN(new_n15887_));
  AOI21_X1   g13451(.A1(new_n15887_), .A2(new_n15885_), .B(new_n12779_), .ZN(new_n15888_));
  AOI22_X1   g13452(.A1(new_n15888_), .A2(new_n15882_), .B1(new_n12779_), .B2(new_n15876_), .ZN(new_n15889_));
  NOR2_X1    g13453(.A1(new_n15889_), .A2(pi0789), .ZN(new_n15890_));
  NOR2_X1    g13454(.A1(new_n15890_), .A2(new_n14303_), .ZN(new_n15891_));
  OAI21_X1   g13455(.A1(new_n15731_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n15892_));
  AND2_X2    g13456(.A1(new_n15806_), .A2(new_n12793_), .Z(new_n15893_));
  OAI21_X1   g13457(.A1(new_n15893_), .A2(new_n15892_), .B(pi0648), .ZN(new_n15894_));
  AOI21_X1   g13458(.A1(new_n15762_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n15895_));
  NAND2_X1   g13459(.A1(new_n15889_), .A2(pi0619), .ZN(new_n15896_));
  AOI21_X1   g13460(.A1(new_n15896_), .A2(new_n15895_), .B(new_n15894_), .ZN(new_n15897_));
  OAI21_X1   g13461(.A1(new_n15731_), .A2(pi0619), .B(pi1159), .ZN(new_n15898_));
  AND2_X2    g13462(.A1(new_n15806_), .A2(pi0619), .Z(new_n15899_));
  OAI21_X1   g13463(.A1(new_n15899_), .A2(new_n15898_), .B(new_n12895_), .ZN(new_n15900_));
  NAND2_X1   g13464(.A1(new_n15762_), .A2(pi0619), .ZN(new_n15901_));
  NAND2_X1   g13465(.A1(new_n15901_), .A2(new_n12791_), .ZN(new_n15902_));
  AOI21_X1   g13466(.A1(new_n15889_), .A2(new_n12793_), .B(new_n15902_), .ZN(new_n15903_));
  OAI21_X1   g13467(.A1(new_n15903_), .A2(new_n15900_), .B(pi0789), .ZN(new_n15904_));
  OAI21_X1   g13468(.A1(new_n15904_), .A2(new_n15897_), .B(new_n15891_), .ZN(new_n15905_));
  NAND2_X1   g13469(.A1(new_n15762_), .A2(new_n12911_), .ZN(new_n15906_));
  NAND2_X1   g13470(.A1(new_n15734_), .A2(new_n12910_), .ZN(new_n15907_));
  AOI21_X1   g13471(.A1(new_n15906_), .A2(new_n15907_), .B(new_n12906_), .ZN(new_n15908_));
  AND2_X2    g13472(.A1(new_n15810_), .A2(new_n12914_), .Z(new_n15909_));
  OAI21_X1   g13473(.A1(new_n15909_), .A2(new_n15908_), .B(pi0788), .ZN(new_n15910_));
  NAND3_X1   g13474(.A1(new_n15905_), .A2(new_n15824_), .A3(new_n15910_), .ZN(new_n15911_));
  AND2_X2    g13475(.A1(new_n15911_), .A2(new_n15823_), .Z(new_n15912_));
  OAI22_X1   g13476(.A1(new_n15912_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n15816_), .ZN(new_n15913_));
  AOI21_X1   g13477(.A1(new_n15734_), .A2(new_n12975_), .B(pi0715), .ZN(new_n15914_));
  NOR2_X1    g13478(.A1(new_n15734_), .A2(new_n12985_), .ZN(new_n15915_));
  AOI21_X1   g13479(.A1(new_n15815_), .A2(new_n12985_), .B(new_n15915_), .ZN(new_n15916_));
  NAND2_X1   g13480(.A1(new_n15916_), .A2(pi0644), .ZN(new_n15917_));
  AOI21_X1   g13481(.A1(new_n15917_), .A2(new_n15914_), .B(new_n12739_), .ZN(new_n15918_));
  AOI21_X1   g13482(.A1(new_n15918_), .A2(pi0644), .B(new_n13000_), .ZN(new_n15919_));
  NOR2_X1    g13483(.A1(new_n15913_), .A2(new_n15919_), .ZN(new_n15920_));
  NOR2_X1    g13484(.A1(new_n15777_), .A2(pi1157), .ZN(new_n15921_));
  NOR2_X1    g13485(.A1(new_n15775_), .A2(new_n12965_), .ZN(new_n15922_));
  OAI21_X1   g13486(.A1(new_n15921_), .A2(new_n15922_), .B(pi0787), .ZN(new_n15923_));
  OAI21_X1   g13487(.A1(pi0787), .A2(new_n15773_), .B(new_n15923_), .ZN(new_n15924_));
  OAI21_X1   g13488(.A1(new_n15924_), .A2(pi0644), .B(pi0715), .ZN(new_n15925_));
  NAND2_X1   g13489(.A1(new_n15925_), .A2(new_n15918_), .ZN(new_n15926_));
  AND2_X2    g13490(.A1(new_n15924_), .A2(pi0644), .Z(new_n15927_));
  AOI21_X1   g13491(.A1(new_n15913_), .A2(new_n12975_), .B(new_n15927_), .ZN(new_n15928_));
  AOI21_X1   g13492(.A1(new_n15734_), .A2(pi0644), .B(new_n12740_), .ZN(new_n15929_));
  NAND2_X1   g13493(.A1(new_n15916_), .A2(new_n12975_), .ZN(new_n15930_));
  AOI21_X1   g13494(.A1(new_n15930_), .A2(new_n15929_), .B(pi1160), .ZN(new_n15931_));
  OAI21_X1   g13495(.A1(new_n15928_), .A2(pi0715), .B(new_n15931_), .ZN(new_n15932_));
  AOI21_X1   g13496(.A1(new_n15932_), .A2(new_n15926_), .B(new_n13000_), .ZN(new_n15933_));
  OAI21_X1   g13497(.A1(new_n15933_), .A2(new_n15920_), .B(new_n6643_), .ZN(new_n15934_));
  AOI22_X1   g13498(.A1(new_n15934_), .A2(new_n15729_), .B1(pi0832), .B2(new_n15728_), .ZN(po0302));
  NOR2_X1    g13499(.A1(new_n5473_), .A2(pi0947), .ZN(new_n15936_));
  AOI22_X1   g13500(.A1(new_n15936_), .A2(pi0735), .B1(pi0743), .B2(pi0947), .ZN(new_n15937_));
  INV_X1     g13501(.I(new_n15937_), .ZN(new_n15938_));
  NOR2_X1    g13502(.A1(new_n3042_), .A2(new_n3107_), .ZN(new_n15939_));
  AOI21_X1   g13503(.A1(new_n15938_), .A2(new_n3042_), .B(new_n15939_), .ZN(new_n15940_));
  OAI21_X1   g13504(.A1(new_n13397_), .A2(new_n15938_), .B(pi0038), .ZN(new_n15941_));
  NOR2_X1    g13505(.A1(new_n13344_), .A2(pi0146), .ZN(new_n15942_));
  OAI21_X1   g13506(.A1(new_n15941_), .A2(new_n15942_), .B(new_n8264_), .ZN(new_n15943_));
  NOR2_X1    g13507(.A1(new_n13058_), .A2(new_n15937_), .ZN(new_n15944_));
  INV_X1     g13508(.I(new_n13058_), .ZN(new_n15945_));
  NOR2_X1    g13509(.A1(new_n15945_), .A2(new_n3107_), .ZN(new_n15946_));
  OAI21_X1   g13510(.A1(new_n15946_), .A2(new_n15944_), .B(new_n2628_), .ZN(new_n15947_));
  NAND2_X1   g13511(.A1(new_n13055_), .A2(pi0146), .ZN(new_n15948_));
  OAI21_X1   g13512(.A1(new_n13055_), .A2(new_n15937_), .B(new_n15948_), .ZN(new_n15949_));
  AOI21_X1   g13513(.A1(new_n15949_), .A2(pi0299), .B(pi0039), .ZN(new_n15950_));
  AOI21_X1   g13514(.A1(new_n15950_), .A2(new_n15947_), .B(pi0038), .ZN(new_n15951_));
  NAND2_X1   g13515(.A1(new_n13179_), .A2(new_n15938_), .ZN(new_n15952_));
  INV_X1     g13516(.I(new_n13179_), .ZN(new_n15953_));
  NAND2_X1   g13517(.A1(new_n15953_), .A2(pi0146), .ZN(new_n15954_));
  AOI21_X1   g13518(.A1(new_n15954_), .A2(new_n15952_), .B(new_n5445_), .ZN(new_n15955_));
  INV_X1     g13519(.I(new_n13175_), .ZN(new_n15956_));
  NOR2_X1    g13520(.A1(new_n15956_), .A2(new_n15937_), .ZN(new_n15957_));
  AOI21_X1   g13521(.A1(pi0146), .A2(new_n15956_), .B(new_n15957_), .ZN(new_n15958_));
  NOR2_X1    g13522(.A1(new_n15958_), .A2(new_n5446_), .ZN(new_n15959_));
  OAI21_X1   g13523(.A1(new_n15959_), .A2(new_n15955_), .B(pi0223), .ZN(new_n15960_));
  NAND2_X1   g13524(.A1(new_n15960_), .A2(new_n2628_), .ZN(new_n15961_));
  NAND2_X1   g13525(.A1(new_n13093_), .A2(new_n3107_), .ZN(new_n15962_));
  NAND2_X1   g13526(.A1(new_n14452_), .A2(new_n15937_), .ZN(new_n15963_));
  AOI21_X1   g13527(.A1(new_n15963_), .A2(new_n15962_), .B(new_n5446_), .ZN(new_n15964_));
  NAND2_X1   g13528(.A1(new_n14577_), .A2(new_n3107_), .ZN(new_n15965_));
  NAND2_X1   g13529(.A1(new_n13126_), .A2(new_n15937_), .ZN(new_n15966_));
  AOI21_X1   g13530(.A1(new_n15965_), .A2(new_n15966_), .B(new_n5445_), .ZN(new_n15967_));
  OAI21_X1   g13531(.A1(new_n15967_), .A2(new_n15964_), .B(new_n2642_), .ZN(new_n15968_));
  NOR2_X1    g13532(.A1(new_n13098_), .A2(pi0146), .ZN(new_n15969_));
  AOI21_X1   g13533(.A1(new_n13098_), .A2(new_n15937_), .B(new_n15969_), .ZN(new_n15970_));
  NOR2_X1    g13534(.A1(new_n15970_), .A2(new_n2642_), .ZN(new_n15971_));
  NOR2_X1    g13535(.A1(new_n15971_), .A2(pi0223), .ZN(new_n15972_));
  AOI21_X1   g13536(.A1(new_n15968_), .A2(new_n15972_), .B(new_n15961_), .ZN(new_n15973_));
  INV_X1     g13537(.I(new_n13174_), .ZN(new_n15974_));
  NOR2_X1    g13538(.A1(new_n15956_), .A2(new_n5420_), .ZN(new_n15975_));
  NOR3_X1    g13539(.A1(new_n15974_), .A2(new_n3107_), .A3(new_n15975_), .ZN(new_n15976_));
  OR3_X2     g13540(.A1(new_n15976_), .A2(new_n2436_), .A3(new_n15957_), .Z(new_n15977_));
  NOR2_X1    g13541(.A1(new_n15970_), .A2(new_n3304_), .ZN(new_n15978_));
  NOR2_X1    g13542(.A1(new_n5419_), .A2(pi0907), .ZN(new_n15979_));
  NOR3_X1    g13543(.A1(new_n14452_), .A2(new_n3107_), .A3(new_n15979_), .ZN(new_n15980_));
  OAI21_X1   g13544(.A1(pi0743), .A2(new_n13093_), .B(new_n15962_), .ZN(new_n15981_));
  NAND3_X1   g13545(.A1(new_n14577_), .A2(pi0146), .A3(new_n15979_), .ZN(new_n15982_));
  NOR2_X1    g13546(.A1(new_n13093_), .A2(new_n5473_), .ZN(new_n15983_));
  AOI21_X1   g13547(.A1(new_n15983_), .A2(pi0735), .B(pi0947), .ZN(new_n15984_));
  AOI22_X1   g13548(.A1(new_n15982_), .A2(new_n15984_), .B1(pi0947), .B2(new_n15981_), .ZN(new_n15985_));
  NOR3_X1    g13549(.A1(new_n15985_), .A2(new_n3303_), .A3(new_n15980_), .ZN(new_n15986_));
  OAI21_X1   g13550(.A1(new_n15986_), .A2(new_n15978_), .B(new_n2436_), .ZN(new_n15987_));
  AOI21_X1   g13551(.A1(new_n15987_), .A2(new_n15977_), .B(new_n2628_), .ZN(new_n15988_));
  OAI21_X1   g13552(.A1(new_n15973_), .A2(new_n15988_), .B(pi0039), .ZN(new_n15989_));
  AOI21_X1   g13553(.A1(new_n15989_), .A2(new_n15951_), .B(new_n15943_), .ZN(new_n15990_));
  OAI21_X1   g13554(.A1(new_n8264_), .A2(pi0146), .B(new_n12738_), .ZN(new_n15991_));
  OAI22_X1   g13555(.A1(new_n15990_), .A2(new_n15991_), .B1(new_n12738_), .B2(new_n15940_), .ZN(po0303));
  INV_X1     g13556(.I(pi0726), .ZN(new_n15993_));
  INV_X1     g13557(.I(new_n15936_), .ZN(new_n15994_));
  OAI22_X1   g13558(.A1(new_n15994_), .A2(new_n15993_), .B1(pi0770), .B2(new_n5692_), .ZN(new_n15995_));
  NAND2_X1   g13559(.A1(new_n3043_), .A2(pi0147), .ZN(new_n15996_));
  OAI21_X1   g13560(.A1(new_n15995_), .A2(new_n3043_), .B(new_n15996_), .ZN(new_n15997_));
  AOI21_X1   g13561(.A1(new_n8265_), .A2(new_n9399_), .B(pi0832), .ZN(new_n15998_));
  AOI21_X1   g13562(.A1(new_n13344_), .A2(new_n15936_), .B(new_n3265_), .ZN(new_n15999_));
  OAI21_X1   g13563(.A1(pi0147), .A2(new_n13344_), .B(new_n15999_), .ZN(new_n16000_));
  NOR3_X1    g13564(.A1(new_n15956_), .A2(new_n2436_), .A3(new_n5692_), .ZN(new_n16001_));
  INV_X1     g13565(.I(new_n13127_), .ZN(new_n16002_));
  NOR2_X1    g13566(.A1(new_n13093_), .A2(new_n5692_), .ZN(new_n16003_));
  NOR2_X1    g13567(.A1(new_n16002_), .A2(new_n16003_), .ZN(new_n16004_));
  NOR2_X1    g13568(.A1(new_n16004_), .A2(new_n3303_), .ZN(new_n16005_));
  INV_X1     g13569(.I(new_n13639_), .ZN(new_n16006_));
  NOR2_X1    g13570(.A1(new_n16006_), .A2(new_n15936_), .ZN(new_n16007_));
  NOR3_X1    g13571(.A1(new_n16005_), .A2(pi0215), .A3(new_n16007_), .ZN(new_n16008_));
  AOI21_X1   g13572(.A1(pi0215), .A2(new_n13174_), .B(new_n16008_), .ZN(new_n16009_));
  NOR2_X1    g13573(.A1(new_n16009_), .A2(new_n16001_), .ZN(new_n16010_));
  NOR2_X1    g13574(.A1(new_n16010_), .A2(new_n2628_), .ZN(new_n16011_));
  INV_X1     g13575(.I(new_n13182_), .ZN(new_n16012_));
  INV_X1     g13576(.I(new_n13187_), .ZN(new_n16013_));
  NOR2_X1    g13577(.A1(new_n16013_), .A2(new_n16012_), .ZN(new_n16014_));
  INV_X1     g13578(.I(new_n16014_), .ZN(new_n16015_));
  NOR2_X1    g13579(.A1(new_n16015_), .A2(pi0299), .ZN(new_n16016_));
  INV_X1     g13580(.I(new_n16016_), .ZN(new_n16017_));
  NOR2_X1    g13581(.A1(new_n16017_), .A2(new_n15936_), .ZN(new_n16018_));
  NOR2_X1    g13582(.A1(new_n16011_), .A2(new_n16018_), .ZN(new_n16019_));
  INV_X1     g13583(.I(new_n16019_), .ZN(new_n16020_));
  AOI22_X1   g13584(.A1(new_n16020_), .A2(pi0039), .B1(new_n13061_), .B2(new_n15994_), .ZN(new_n16021_));
  NOR2_X1    g13585(.A1(new_n16021_), .A2(pi0147), .ZN(new_n16022_));
  NOR2_X1    g13586(.A1(new_n13060_), .A2(new_n15994_), .ZN(new_n16023_));
  NOR2_X1    g13587(.A1(new_n16023_), .A2(pi0039), .ZN(new_n16024_));
  AOI21_X1   g13588(.A1(new_n16014_), .A2(new_n15936_), .B(pi0299), .ZN(new_n16025_));
  NOR2_X1    g13589(.A1(new_n15956_), .A2(new_n15994_), .ZN(new_n16026_));
  INV_X1     g13590(.I(new_n16026_), .ZN(new_n16027_));
  NOR2_X1    g13591(.A1(new_n13093_), .A2(new_n15994_), .ZN(new_n16028_));
  NOR2_X1    g13592(.A1(new_n16028_), .A2(new_n3303_), .ZN(new_n16029_));
  NOR2_X1    g13593(.A1(new_n13088_), .A2(new_n15994_), .ZN(new_n16030_));
  OAI21_X1   g13594(.A1(new_n16030_), .A2(new_n3304_), .B(new_n2436_), .ZN(new_n16031_));
  OAI22_X1   g13595(.A1(new_n16027_), .A2(new_n2436_), .B1(new_n16029_), .B2(new_n16031_), .ZN(new_n16032_));
  NOR2_X1    g13596(.A1(new_n16032_), .A2(new_n2628_), .ZN(new_n16033_));
  NOR2_X1    g13597(.A1(new_n16025_), .A2(new_n16033_), .ZN(new_n16034_));
  INV_X1     g13598(.I(new_n16034_), .ZN(new_n16035_));
  AOI21_X1   g13599(.A1(new_n16035_), .A2(pi0039), .B(new_n16024_), .ZN(new_n16036_));
  NOR2_X1    g13600(.A1(new_n16036_), .A2(new_n9399_), .ZN(new_n16037_));
  OAI21_X1   g13601(.A1(new_n16022_), .A2(new_n16037_), .B(new_n3265_), .ZN(new_n16038_));
  NAND3_X1   g13602(.A1(new_n16038_), .A2(pi0770), .A3(new_n16000_), .ZN(new_n16039_));
  NAND2_X1   g13603(.A1(new_n13180_), .A2(new_n13181_), .ZN(new_n16040_));
  INV_X1     g13604(.I(new_n16040_), .ZN(new_n16041_));
  NOR2_X1    g13605(.A1(new_n16041_), .A2(pi0947), .ZN(new_n16042_));
  NOR2_X1    g13606(.A1(new_n16042_), .A2(new_n2668_), .ZN(new_n16043_));
  AOI21_X1   g13607(.A1(new_n16040_), .A2(new_n15994_), .B(new_n2668_), .ZN(new_n16044_));
  INV_X1     g13608(.I(new_n13185_), .ZN(new_n16045_));
  OAI22_X1   g13609(.A1(new_n13184_), .A2(new_n2641_), .B1(new_n2530_), .B2(new_n16045_), .ZN(new_n16046_));
  AOI21_X1   g13610(.A1(new_n16046_), .A2(new_n5420_), .B(pi0223), .ZN(new_n16047_));
  NOR3_X1    g13611(.A1(new_n16043_), .A2(new_n16044_), .A3(new_n16047_), .ZN(new_n16048_));
  NOR2_X1    g13612(.A1(new_n16048_), .A2(pi0299), .ZN(new_n16049_));
  AOI21_X1   g13613(.A1(new_n16009_), .A2(new_n5692_), .B(new_n2628_), .ZN(new_n16050_));
  NOR2_X1    g13614(.A1(new_n16050_), .A2(new_n16049_), .ZN(new_n16051_));
  INV_X1     g13615(.I(new_n16051_), .ZN(new_n16052_));
  OAI22_X1   g13616(.A1(new_n16052_), .A2(new_n2627_), .B1(new_n5421_), .B2(new_n13336_), .ZN(new_n16053_));
  NOR2_X1    g13617(.A1(new_n16015_), .A2(new_n5420_), .ZN(new_n16054_));
  INV_X1     g13618(.I(new_n16054_), .ZN(new_n16055_));
  INV_X1     g13619(.I(new_n13176_), .ZN(new_n16056_));
  INV_X1     g13620(.I(new_n13128_), .ZN(new_n16057_));
  NOR2_X1    g13621(.A1(new_n13088_), .A2(new_n5420_), .ZN(new_n16058_));
  NOR2_X1    g13622(.A1(new_n16058_), .A2(new_n3304_), .ZN(new_n16059_));
  OAI21_X1   g13623(.A1(new_n16057_), .A2(new_n16059_), .B(new_n2436_), .ZN(new_n16060_));
  NAND3_X1   g13624(.A1(new_n16060_), .A2(pi0299), .A3(new_n16056_), .ZN(new_n16061_));
  OAI21_X1   g13625(.A1(new_n16055_), .A2(pi0299), .B(new_n16061_), .ZN(new_n16062_));
  NOR2_X1    g13626(.A1(new_n13060_), .A2(new_n5420_), .ZN(new_n16063_));
  INV_X1     g13627(.I(new_n16063_), .ZN(new_n16064_));
  NOR2_X1    g13628(.A1(new_n16064_), .A2(pi0039), .ZN(new_n16065_));
  AOI21_X1   g13629(.A1(new_n16062_), .A2(pi0039), .B(new_n16065_), .ZN(new_n16066_));
  INV_X1     g13630(.I(new_n16066_), .ZN(new_n16067_));
  NOR2_X1    g13631(.A1(new_n16067_), .A2(new_n9399_), .ZN(new_n16068_));
  AOI21_X1   g13632(.A1(new_n16053_), .A2(new_n9399_), .B(new_n16068_), .ZN(new_n16069_));
  NAND2_X1   g13633(.A1(new_n13344_), .A2(new_n5421_), .ZN(new_n16070_));
  NAND2_X1   g13634(.A1(new_n16070_), .A2(pi0038), .ZN(new_n16071_));
  INV_X1     g13635(.I(new_n16071_), .ZN(new_n16072_));
  INV_X1     g13636(.I(new_n13004_), .ZN(new_n16073_));
  NOR2_X1    g13637(.A1(new_n16073_), .A2(new_n5421_), .ZN(new_n16074_));
  INV_X1     g13638(.I(new_n16074_), .ZN(new_n16075_));
  NAND2_X1   g13639(.A1(new_n16075_), .A2(new_n9399_), .ZN(new_n16076_));
  AOI21_X1   g13640(.A1(new_n16076_), .A2(new_n16072_), .B(pi0770), .ZN(new_n16077_));
  OAI21_X1   g13641(.A1(new_n16069_), .A2(pi0038), .B(new_n16077_), .ZN(new_n16078_));
  NAND3_X1   g13642(.A1(new_n16039_), .A2(pi0726), .A3(new_n16078_), .ZN(new_n16079_));
  INV_X1     g13643(.I(pi0770), .ZN(new_n16080_));
  AOI21_X1   g13644(.A1(new_n13004_), .A2(pi0947), .B(new_n3265_), .ZN(new_n16081_));
  NOR2_X1    g13645(.A1(new_n13060_), .A2(new_n5692_), .ZN(new_n16082_));
  NOR2_X1    g13646(.A1(new_n16082_), .A2(pi0039), .ZN(new_n16083_));
  NAND2_X1   g13647(.A1(new_n16014_), .A2(pi0947), .ZN(new_n16084_));
  NAND2_X1   g13648(.A1(new_n16084_), .A2(new_n2628_), .ZN(new_n16085_));
  INV_X1     g13649(.I(new_n16085_), .ZN(new_n16086_));
  NOR2_X1    g13650(.A1(new_n16003_), .A2(new_n3303_), .ZN(new_n16087_));
  NOR2_X1    g13651(.A1(new_n13088_), .A2(new_n5692_), .ZN(new_n16088_));
  NOR2_X1    g13652(.A1(new_n16088_), .A2(new_n3304_), .ZN(new_n16089_));
  NOR3_X1    g13653(.A1(new_n16087_), .A2(pi0215), .A3(new_n16089_), .ZN(new_n16090_));
  NOR2_X1    g13654(.A1(new_n16001_), .A2(new_n2628_), .ZN(new_n16091_));
  INV_X1     g13655(.I(new_n16091_), .ZN(new_n16092_));
  NOR2_X1    g13656(.A1(new_n16092_), .A2(new_n16090_), .ZN(new_n16093_));
  NOR2_X1    g13657(.A1(new_n16086_), .A2(new_n16093_), .ZN(new_n16094_));
  INV_X1     g13658(.I(new_n16094_), .ZN(new_n16095_));
  AOI21_X1   g13659(.A1(new_n16095_), .A2(pi0039), .B(new_n16083_), .ZN(new_n16096_));
  NOR2_X1    g13660(.A1(new_n16096_), .A2(pi0038), .ZN(new_n16097_));
  NOR2_X1    g13661(.A1(new_n16097_), .A2(new_n16081_), .ZN(new_n16098_));
  NAND3_X1   g13662(.A1(new_n16098_), .A2(pi0147), .A3(new_n16080_), .ZN(new_n16099_));
  NOR3_X1    g13663(.A1(new_n16073_), .A2(new_n3265_), .A3(pi0947), .ZN(new_n16100_));
  INV_X1     g13664(.I(new_n16100_), .ZN(new_n16101_));
  INV_X1     g13665(.I(new_n13060_), .ZN(new_n16102_));
  AOI21_X1   g13666(.A1(new_n16102_), .A2(new_n5692_), .B(pi0039), .ZN(new_n16103_));
  INV_X1     g13667(.I(new_n16103_), .ZN(new_n16104_));
  NOR2_X1    g13668(.A1(new_n15974_), .A2(new_n2436_), .ZN(new_n16105_));
  INV_X1     g13669(.I(new_n16105_), .ZN(new_n16106_));
  NOR2_X1    g13670(.A1(new_n16106_), .A2(new_n16026_), .ZN(new_n16107_));
  NOR2_X1    g13671(.A1(new_n16002_), .A2(new_n16028_), .ZN(new_n16108_));
  NOR2_X1    g13672(.A1(new_n16108_), .A2(new_n3303_), .ZN(new_n16109_));
  NOR2_X1    g13673(.A1(new_n16109_), .A2(pi0215), .ZN(new_n16110_));
  INV_X1     g13674(.I(new_n16110_), .ZN(new_n16111_));
  AOI21_X1   g13675(.A1(new_n5692_), .A2(new_n13639_), .B(new_n16111_), .ZN(new_n16112_));
  NOR2_X1    g13676(.A1(new_n16112_), .A2(new_n16107_), .ZN(new_n16113_));
  INV_X1     g13677(.I(new_n16113_), .ZN(new_n16114_));
  NOR2_X1    g13678(.A1(new_n16114_), .A2(new_n2628_), .ZN(new_n16115_));
  INV_X1     g13679(.I(new_n16115_), .ZN(new_n16116_));
  OAI21_X1   g13680(.A1(pi0947), .A2(new_n16017_), .B(new_n16116_), .ZN(new_n16117_));
  OAI21_X1   g13681(.A1(new_n16117_), .A2(new_n2627_), .B(new_n16104_), .ZN(new_n16118_));
  OAI21_X1   g13682(.A1(new_n16118_), .A2(pi0038), .B(new_n16101_), .ZN(new_n16119_));
  NOR2_X1    g13683(.A1(new_n16119_), .A2(pi0770), .ZN(new_n16120_));
  NOR2_X1    g13684(.A1(new_n13191_), .A2(new_n16080_), .ZN(new_n16121_));
  OAI21_X1   g13685(.A1(new_n16120_), .A2(new_n16121_), .B(new_n9399_), .ZN(new_n16122_));
  NAND3_X1   g13686(.A1(new_n16122_), .A2(new_n15993_), .A3(new_n16099_), .ZN(new_n16123_));
  NAND3_X1   g13687(.A1(new_n16123_), .A2(new_n8264_), .A3(new_n16079_), .ZN(new_n16124_));
  AOI22_X1   g13688(.A1(new_n16124_), .A2(new_n15998_), .B1(pi0832), .B2(new_n15997_), .ZN(po0304));
  NOR2_X1    g13689(.A1(new_n14059_), .A2(new_n5692_), .ZN(new_n16126_));
  NOR2_X1    g13690(.A1(new_n15994_), .A2(new_n13935_), .ZN(new_n16127_));
  NOR3_X1    g13691(.A1(new_n16127_), .A2(new_n3043_), .A3(new_n16126_), .ZN(new_n16128_));
  OAI21_X1   g13692(.A1(new_n3042_), .A2(new_n4257_), .B(pi0832), .ZN(new_n16129_));
  OAI21_X1   g13693(.A1(new_n2582_), .A2(new_n4257_), .B(new_n12738_), .ZN(new_n16130_));
  AOI21_X1   g13694(.A1(new_n13060_), .A2(new_n4257_), .B(pi0039), .ZN(new_n16131_));
  OAI21_X1   g13695(.A1(pi0749), .A2(new_n5692_), .B(new_n16063_), .ZN(new_n16132_));
  AOI21_X1   g13696(.A1(new_n16132_), .A2(new_n16131_), .B(pi0038), .ZN(new_n16133_));
  NAND2_X1   g13697(.A1(new_n16052_), .A2(new_n4257_), .ZN(new_n16134_));
  NAND2_X1   g13698(.A1(new_n16062_), .A2(pi0148), .ZN(new_n16135_));
  AOI21_X1   g13699(.A1(new_n16134_), .A2(new_n16135_), .B(new_n14059_), .ZN(new_n16136_));
  AOI21_X1   g13700(.A1(pi0299), .A2(new_n16032_), .B(new_n16016_), .ZN(new_n16137_));
  NAND2_X1   g13701(.A1(new_n16137_), .A2(pi0148), .ZN(new_n16138_));
  NAND2_X1   g13702(.A1(new_n16138_), .A2(new_n14059_), .ZN(new_n16139_));
  NOR2_X1    g13703(.A1(new_n16019_), .A2(new_n12662_), .ZN(new_n16140_));
  OAI21_X1   g13704(.A1(new_n16140_), .A2(new_n16139_), .B(pi0039), .ZN(new_n16141_));
  OAI21_X1   g13705(.A1(new_n16141_), .A2(new_n16136_), .B(new_n16133_), .ZN(new_n16142_));
  NOR2_X1    g13706(.A1(new_n5692_), .A2(pi0749), .ZN(new_n16143_));
  OAI22_X1   g13707(.A1(new_n16070_), .A2(new_n16143_), .B1(pi0148), .B2(new_n13344_), .ZN(new_n16144_));
  AOI21_X1   g13708(.A1(new_n16144_), .A2(pi0038), .B(new_n13935_), .ZN(new_n16145_));
  NAND2_X1   g13709(.A1(new_n16142_), .A2(new_n16145_), .ZN(new_n16146_));
  NOR2_X1    g13710(.A1(new_n2610_), .A2(new_n6165_), .ZN(new_n16147_));
  INV_X1     g13711(.I(new_n16147_), .ZN(new_n16148_));
  NOR2_X1    g13712(.A1(new_n13397_), .A2(new_n16126_), .ZN(new_n16149_));
  NOR2_X1    g13713(.A1(new_n16149_), .A2(new_n3265_), .ZN(new_n16150_));
  NAND2_X1   g13714(.A1(new_n16073_), .A2(pi0148), .ZN(new_n16151_));
  AOI21_X1   g13715(.A1(new_n16151_), .A2(new_n16150_), .B(pi0706), .ZN(new_n16152_));
  NAND2_X1   g13716(.A1(new_n16102_), .A2(new_n16126_), .ZN(new_n16153_));
  AOI21_X1   g13717(.A1(new_n16153_), .A2(new_n16131_), .B(pi0038), .ZN(new_n16154_));
  NAND2_X1   g13718(.A1(new_n4257_), .A2(new_n14059_), .ZN(new_n16155_));
  OAI21_X1   g13719(.A1(new_n14064_), .A2(new_n16155_), .B(pi0039), .ZN(new_n16156_));
  NOR2_X1    g13720(.A1(new_n16090_), .A2(new_n16001_), .ZN(new_n16157_));
  NAND2_X1   g13721(.A1(new_n16157_), .A2(pi0148), .ZN(new_n16158_));
  OAI21_X1   g13722(.A1(new_n16114_), .A2(pi0148), .B(new_n16158_), .ZN(new_n16159_));
  NOR2_X1    g13723(.A1(new_n16014_), .A2(pi0148), .ZN(new_n16160_));
  OAI21_X1   g13724(.A1(new_n16085_), .A2(new_n16160_), .B(pi0749), .ZN(new_n16161_));
  AOI21_X1   g13725(.A1(new_n16159_), .A2(pi0299), .B(new_n16161_), .ZN(new_n16162_));
  OAI21_X1   g13726(.A1(new_n16162_), .A2(new_n16156_), .B(new_n16154_), .ZN(new_n16163_));
  AOI21_X1   g13727(.A1(new_n16163_), .A2(new_n16152_), .B(new_n16148_), .ZN(new_n16164_));
  OAI21_X1   g13728(.A1(new_n16147_), .A2(pi0148), .B(new_n2582_), .ZN(new_n16165_));
  AOI21_X1   g13729(.A1(new_n16146_), .A2(new_n16164_), .B(new_n16165_), .ZN(new_n16166_));
  OAI22_X1   g13730(.A1(new_n16166_), .A2(new_n16130_), .B1(new_n16128_), .B2(new_n16129_), .ZN(po0305));
  INV_X1     g13731(.I(pi0725), .ZN(new_n16168_));
  INV_X1     g13732(.I(pi0755), .ZN(new_n16169_));
  NOR2_X1    g13733(.A1(new_n16018_), .A2(new_n16169_), .ZN(new_n16170_));
  NOR2_X1    g13734(.A1(new_n16011_), .A2(pi0149), .ZN(new_n16171_));
  NOR2_X1    g13735(.A1(new_n16137_), .A2(new_n7455_), .ZN(new_n16172_));
  OAI21_X1   g13736(.A1(new_n16171_), .A2(new_n16172_), .B(new_n16170_), .ZN(new_n16173_));
  NOR2_X1    g13737(.A1(new_n16051_), .A2(pi0149), .ZN(new_n16174_));
  INV_X1     g13738(.I(new_n16062_), .ZN(new_n16175_));
  NOR2_X1    g13739(.A1(new_n16175_), .A2(new_n7455_), .ZN(new_n16176_));
  OAI21_X1   g13740(.A1(new_n16174_), .A2(new_n16176_), .B(new_n16169_), .ZN(new_n16177_));
  NAND3_X1   g13741(.A1(new_n16177_), .A2(new_n16173_), .A3(pi0039), .ZN(new_n16178_));
  NOR2_X1    g13742(.A1(new_n5692_), .A2(pi0755), .ZN(new_n16179_));
  NOR2_X1    g13743(.A1(new_n13060_), .A2(new_n16179_), .ZN(new_n16180_));
  NOR2_X1    g13744(.A1(new_n16102_), .A2(new_n7455_), .ZN(new_n16181_));
  OAI21_X1   g13745(.A1(new_n16181_), .A2(new_n16180_), .B(new_n2627_), .ZN(new_n16182_));
  OR2_X2     g13746(.A1(new_n16182_), .A2(new_n16023_), .Z(new_n16183_));
  AOI21_X1   g13747(.A1(new_n16178_), .A2(new_n16183_), .B(pi0038), .ZN(new_n16184_));
  NOR2_X1    g13748(.A1(new_n13568_), .A2(new_n5420_), .ZN(new_n16185_));
  INV_X1     g13749(.I(new_n16185_), .ZN(new_n16186_));
  NOR2_X1    g13750(.A1(new_n16169_), .A2(new_n5692_), .ZN(new_n16187_));
  NOR3_X1    g13751(.A1(new_n16186_), .A2(pi0039), .A3(new_n16187_), .ZN(new_n16188_));
  OAI21_X1   g13752(.A1(new_n13344_), .A2(pi0149), .B(pi0038), .ZN(new_n16189_));
  OAI21_X1   g13753(.A1(new_n16188_), .A2(new_n16189_), .B(new_n16168_), .ZN(new_n16190_));
  INV_X1     g13754(.I(new_n16179_), .ZN(new_n16191_));
  AOI21_X1   g13755(.A1(new_n13344_), .A2(new_n16191_), .B(new_n3265_), .ZN(new_n16192_));
  NAND2_X1   g13756(.A1(new_n16073_), .A2(pi0149), .ZN(new_n16193_));
  NOR2_X1    g13757(.A1(new_n16169_), .A2(pi0149), .ZN(new_n16194_));
  AOI21_X1   g13758(.A1(new_n14065_), .A2(new_n16194_), .B(new_n2627_), .ZN(new_n16195_));
  OAI21_X1   g13759(.A1(pi0149), .A2(new_n16014_), .B(new_n16086_), .ZN(new_n16196_));
  OAI21_X1   g13760(.A1(new_n16113_), .A2(pi0149), .B(new_n16093_), .ZN(new_n16197_));
  NAND2_X1   g13761(.A1(new_n16115_), .A2(new_n7455_), .ZN(new_n16198_));
  NAND4_X1   g13762(.A1(new_n16198_), .A2(new_n16169_), .A3(new_n16196_), .A4(new_n16197_), .ZN(new_n16199_));
  AOI21_X1   g13763(.A1(new_n16199_), .A2(new_n16195_), .B(pi0038), .ZN(new_n16200_));
  AOI22_X1   g13764(.A1(new_n16200_), .A2(new_n16182_), .B1(new_n16192_), .B2(new_n16193_), .ZN(new_n16201_));
  OAI22_X1   g13765(.A1(new_n16201_), .A2(new_n16168_), .B1(new_n16184_), .B2(new_n16190_), .ZN(new_n16202_));
  NAND2_X1   g13766(.A1(new_n8265_), .A2(pi0149), .ZN(new_n16203_));
  OAI21_X1   g13767(.A1(new_n16202_), .A2(new_n8265_), .B(new_n16203_), .ZN(new_n16204_));
  NAND2_X1   g13768(.A1(new_n15936_), .A2(new_n16168_), .ZN(new_n16205_));
  NAND3_X1   g13769(.A1(new_n16205_), .A2(new_n16191_), .A3(new_n3042_), .ZN(new_n16206_));
  NAND2_X1   g13770(.A1(new_n3043_), .A2(pi0149), .ZN(new_n16207_));
  AOI21_X1   g13771(.A1(new_n16206_), .A2(new_n16207_), .B(new_n12738_), .ZN(new_n16208_));
  AOI21_X1   g13772(.A1(new_n16204_), .A2(new_n12738_), .B(new_n16208_), .ZN(po0306));
  INV_X1     g13773(.I(pi0751), .ZN(new_n16210_));
  NOR2_X1    g13774(.A1(new_n16102_), .A2(pi0150), .ZN(new_n16211_));
  AOI21_X1   g13775(.A1(new_n16210_), .A2(new_n16102_), .B(new_n16211_), .ZN(new_n16212_));
  NAND2_X1   g13776(.A1(new_n16094_), .A2(pi0150), .ZN(new_n16213_));
  OAI21_X1   g13777(.A1(new_n16117_), .A2(pi0150), .B(new_n16213_), .ZN(new_n16214_));
  NOR2_X1    g13778(.A1(new_n16210_), .A2(pi0150), .ZN(new_n16215_));
  AOI22_X1   g13779(.A1(new_n16214_), .A2(new_n16210_), .B1(new_n14065_), .B2(new_n16215_), .ZN(new_n16216_));
  OAI22_X1   g13780(.A1(new_n16216_), .A2(new_n2627_), .B1(new_n16104_), .B2(new_n16212_), .ZN(new_n16217_));
  INV_X1     g13781(.I(pi0701), .ZN(new_n16218_));
  NOR2_X1    g13782(.A1(new_n5692_), .A2(pi0751), .ZN(new_n16219_));
  OAI22_X1   g13783(.A1(new_n13004_), .A2(new_n10672_), .B1(new_n13397_), .B2(new_n16219_), .ZN(new_n16220_));
  AOI21_X1   g13784(.A1(new_n16220_), .A2(pi0038), .B(new_n16218_), .ZN(new_n16221_));
  OAI21_X1   g13785(.A1(new_n16217_), .A2(pi0038), .B(new_n16221_), .ZN(new_n16222_));
  NAND2_X1   g13786(.A1(new_n16052_), .A2(new_n10672_), .ZN(new_n16223_));
  NAND2_X1   g13787(.A1(new_n16062_), .A2(pi0150), .ZN(new_n16224_));
  AOI21_X1   g13788(.A1(new_n16223_), .A2(new_n16224_), .B(pi0751), .ZN(new_n16225_));
  NAND2_X1   g13789(.A1(new_n16034_), .A2(pi0150), .ZN(new_n16226_));
  NAND2_X1   g13790(.A1(new_n16019_), .A2(new_n10672_), .ZN(new_n16227_));
  AOI21_X1   g13791(.A1(new_n16227_), .A2(new_n16226_), .B(new_n16210_), .ZN(new_n16228_));
  OAI21_X1   g13792(.A1(new_n16228_), .A2(new_n16225_), .B(pi0039), .ZN(new_n16229_));
  NOR2_X1    g13793(.A1(new_n16210_), .A2(new_n5692_), .ZN(new_n16230_));
  NOR3_X1    g13794(.A1(new_n13060_), .A2(new_n5420_), .A3(new_n16230_), .ZN(new_n16231_));
  OAI21_X1   g13795(.A1(new_n16211_), .A2(new_n16231_), .B(new_n2627_), .ZN(new_n16232_));
  NAND3_X1   g13796(.A1(new_n16229_), .A2(new_n3265_), .A3(new_n16232_), .ZN(new_n16233_));
  OR3_X2     g13797(.A1(new_n16186_), .A2(pi0039), .A3(new_n16230_), .Z(new_n16234_));
  AOI21_X1   g13798(.A1(new_n13397_), .A2(new_n10672_), .B(new_n3265_), .ZN(new_n16235_));
  AOI21_X1   g13799(.A1(new_n16234_), .A2(new_n16235_), .B(pi0701), .ZN(new_n16236_));
  NAND2_X1   g13800(.A1(new_n16233_), .A2(new_n16236_), .ZN(new_n16237_));
  NAND3_X1   g13801(.A1(new_n16222_), .A2(new_n8264_), .A3(new_n16237_), .ZN(new_n16238_));
  OAI21_X1   g13802(.A1(new_n10672_), .A2(new_n8264_), .B(new_n16238_), .ZN(new_n16239_));
  AOI21_X1   g13803(.A1(new_n16218_), .A2(new_n15936_), .B(new_n16219_), .ZN(new_n16240_));
  NAND2_X1   g13804(.A1(new_n16240_), .A2(new_n3042_), .ZN(new_n16241_));
  NAND2_X1   g13805(.A1(new_n3043_), .A2(pi0150), .ZN(new_n16242_));
  AOI21_X1   g13806(.A1(new_n16241_), .A2(new_n16242_), .B(new_n12738_), .ZN(new_n16243_));
  AOI21_X1   g13807(.A1(new_n16239_), .A2(new_n12738_), .B(new_n16243_), .ZN(po0307));
  INV_X1     g13808(.I(pi0745), .ZN(new_n16245_));
  INV_X1     g13809(.I(new_n13178_), .ZN(new_n16246_));
  OAI22_X1   g13810(.A1(new_n16246_), .A2(new_n16245_), .B1(new_n16014_), .B2(pi0299), .ZN(new_n16247_));
  NOR2_X1    g13811(.A1(new_n13093_), .A2(new_n5420_), .ZN(new_n16248_));
  OAI21_X1   g13812(.A1(new_n3533_), .A2(new_n16248_), .B(new_n13127_), .ZN(new_n16249_));
  NAND2_X1   g13813(.A1(new_n13088_), .A2(new_n3533_), .ZN(new_n16250_));
  AOI22_X1   g13814(.A1(new_n16249_), .A2(new_n3304_), .B1(new_n16089_), .B2(new_n16250_), .ZN(new_n16251_));
  AOI21_X1   g13815(.A1(new_n16110_), .A2(new_n16251_), .B(new_n2628_), .ZN(new_n16252_));
  INV_X1     g13816(.I(new_n15975_), .ZN(new_n16253_));
  NOR2_X1    g13817(.A1(new_n15974_), .A2(new_n16026_), .ZN(new_n16254_));
  NAND2_X1   g13818(.A1(new_n16254_), .A2(new_n3533_), .ZN(new_n16255_));
  AOI21_X1   g13819(.A1(new_n16255_), .A2(new_n16253_), .B(new_n2436_), .ZN(new_n16256_));
  NAND2_X1   g13820(.A1(new_n16256_), .A2(new_n16027_), .ZN(new_n16257_));
  AOI21_X1   g13821(.A1(new_n16252_), .A2(new_n16257_), .B(pi0745), .ZN(new_n16258_));
  AOI22_X1   g13822(.A1(new_n16258_), .A2(new_n16085_), .B1(new_n3533_), .B2(new_n16247_), .ZN(new_n16259_));
  AOI22_X1   g13823(.A1(new_n16082_), .A2(new_n16245_), .B1(new_n3533_), .B2(new_n13060_), .ZN(new_n16260_));
  AND2_X2    g13824(.A1(new_n16260_), .A2(new_n2627_), .Z(new_n16261_));
  AOI21_X1   g13825(.A1(new_n16259_), .A2(pi0039), .B(new_n16261_), .ZN(new_n16262_));
  INV_X1     g13826(.I(pi0723), .ZN(new_n16263_));
  NOR2_X1    g13827(.A1(new_n5692_), .A2(pi0745), .ZN(new_n16264_));
  OAI22_X1   g13828(.A1(new_n13004_), .A2(new_n3533_), .B1(new_n13397_), .B2(new_n16264_), .ZN(new_n16265_));
  AOI21_X1   g13829(.A1(new_n16265_), .A2(pi0038), .B(new_n16263_), .ZN(new_n16266_));
  OAI21_X1   g13830(.A1(new_n16262_), .A2(pi0038), .B(new_n16266_), .ZN(new_n16267_));
  INV_X1     g13831(.I(new_n16049_), .ZN(new_n16268_));
  AOI21_X1   g13832(.A1(pi0151), .A2(new_n16055_), .B(new_n16268_), .ZN(new_n16269_));
  NOR2_X1    g13833(.A1(new_n16030_), .A2(new_n3304_), .ZN(new_n16270_));
  INV_X1     g13834(.I(new_n16058_), .ZN(new_n16271_));
  NAND3_X1   g13835(.A1(new_n16270_), .A2(new_n16271_), .A3(new_n16250_), .ZN(new_n16272_));
  AOI21_X1   g13836(.A1(new_n16249_), .A2(new_n3304_), .B(pi0215), .ZN(new_n16273_));
  AOI21_X1   g13837(.A1(new_n16272_), .A2(new_n16273_), .B(new_n16256_), .ZN(new_n16274_));
  NOR2_X1    g13838(.A1(new_n16274_), .A2(new_n2628_), .ZN(new_n16275_));
  OAI21_X1   g13839(.A1(new_n16269_), .A2(new_n16275_), .B(new_n16245_), .ZN(new_n16276_));
  NAND2_X1   g13840(.A1(new_n16015_), .A2(new_n3533_), .ZN(new_n16277_));
  AOI21_X1   g13841(.A1(new_n16277_), .A2(new_n16025_), .B(new_n16245_), .ZN(new_n16278_));
  AOI21_X1   g13842(.A1(new_n16270_), .A2(new_n16250_), .B(new_n16005_), .ZN(new_n16279_));
  AOI21_X1   g13843(.A1(new_n16279_), .A2(new_n16273_), .B(new_n16256_), .ZN(new_n16280_));
  OAI21_X1   g13844(.A1(new_n16280_), .A2(new_n16001_), .B(pi0299), .ZN(new_n16281_));
  AOI21_X1   g13845(.A1(new_n16281_), .A2(new_n16278_), .B(new_n2627_), .ZN(new_n16282_));
  AOI22_X1   g13846(.A1(new_n16276_), .A2(new_n16282_), .B1(new_n16024_), .B2(new_n16260_), .ZN(new_n16283_));
  NAND2_X1   g13847(.A1(pi0745), .A2(pi0947), .ZN(new_n16284_));
  NAND3_X1   g13848(.A1(new_n16185_), .A2(new_n2627_), .A3(new_n16284_), .ZN(new_n16285_));
  AOI21_X1   g13849(.A1(new_n13397_), .A2(new_n3533_), .B(new_n3265_), .ZN(new_n16286_));
  AOI21_X1   g13850(.A1(new_n16286_), .A2(new_n16285_), .B(pi0723), .ZN(new_n16287_));
  OAI21_X1   g13851(.A1(new_n16283_), .A2(pi0038), .B(new_n16287_), .ZN(new_n16288_));
  NAND3_X1   g13852(.A1(new_n16288_), .A2(new_n8264_), .A3(new_n16267_), .ZN(new_n16289_));
  OAI21_X1   g13853(.A1(new_n3533_), .A2(new_n8264_), .B(new_n16289_), .ZN(new_n16290_));
  AOI21_X1   g13854(.A1(new_n16263_), .A2(new_n15936_), .B(new_n16264_), .ZN(new_n16291_));
  NAND2_X1   g13855(.A1(new_n16291_), .A2(new_n3042_), .ZN(new_n16292_));
  NAND2_X1   g13856(.A1(new_n3043_), .A2(pi0151), .ZN(new_n16293_));
  AOI21_X1   g13857(.A1(new_n16292_), .A2(new_n16293_), .B(new_n12738_), .ZN(new_n16294_));
  AOI21_X1   g13858(.A1(new_n16290_), .A2(new_n12738_), .B(new_n16294_), .ZN(po0308));
  INV_X1     g13859(.I(pi0759), .ZN(new_n16296_));
  NOR2_X1    g13860(.A1(new_n16296_), .A2(new_n5692_), .ZN(new_n16297_));
  NOR2_X1    g13861(.A1(new_n13060_), .A2(new_n16297_), .ZN(new_n16298_));
  NOR2_X1    g13862(.A1(new_n16102_), .A2(pi0152), .ZN(new_n16299_));
  OAI21_X1   g13863(.A1(new_n16299_), .A2(new_n16298_), .B(new_n2627_), .ZN(new_n16300_));
  NOR2_X1    g13864(.A1(new_n3369_), .A2(pi0759), .ZN(new_n16301_));
  AOI21_X1   g13865(.A1(new_n14065_), .A2(new_n16301_), .B(new_n2627_), .ZN(new_n16302_));
  INV_X1     g13866(.I(new_n16109_), .ZN(new_n16303_));
  INV_X1     g13867(.I(new_n16004_), .ZN(new_n16304_));
  OAI21_X1   g13868(.A1(new_n16304_), .A2(new_n3369_), .B(new_n16029_), .ZN(new_n16305_));
  AOI21_X1   g13869(.A1(new_n16305_), .A2(new_n16303_), .B(new_n16003_), .ZN(new_n16306_));
  INV_X1     g13870(.I(new_n16088_), .ZN(new_n16307_));
  NAND2_X1   g13871(.A1(new_n13088_), .A2(pi0152), .ZN(new_n16308_));
  NAND2_X1   g13872(.A1(new_n16307_), .A2(new_n16308_), .ZN(new_n16309_));
  OAI21_X1   g13873(.A1(new_n16309_), .A2(new_n3304_), .B(new_n2436_), .ZN(new_n16310_));
  AOI21_X1   g13874(.A1(new_n16107_), .A2(pi0152), .B(new_n16092_), .ZN(new_n16311_));
  OAI21_X1   g13875(.A1(new_n16306_), .A2(new_n16310_), .B(new_n16311_), .ZN(new_n16312_));
  NOR2_X1    g13876(.A1(new_n13184_), .A2(new_n5692_), .ZN(new_n16313_));
  INV_X1     g13877(.I(new_n16313_), .ZN(new_n16314_));
  INV_X1     g13878(.I(new_n13184_), .ZN(new_n16315_));
  NOR2_X1    g13879(.A1(new_n16315_), .A2(new_n3369_), .ZN(new_n16316_));
  INV_X1     g13880(.I(new_n16316_), .ZN(new_n16317_));
  AOI21_X1   g13881(.A1(new_n16317_), .A2(new_n16314_), .B(new_n2641_), .ZN(new_n16318_));
  AOI21_X1   g13882(.A1(new_n2641_), .A2(new_n16309_), .B(new_n16318_), .ZN(new_n16319_));
  NAND2_X1   g13883(.A1(new_n16041_), .A2(new_n3369_), .ZN(new_n16320_));
  AOI21_X1   g13884(.A1(new_n16043_), .A2(new_n16320_), .B(pi0299), .ZN(new_n16321_));
  OAI21_X1   g13885(.A1(new_n16319_), .A2(pi0223), .B(new_n16321_), .ZN(new_n16322_));
  NAND3_X1   g13886(.A1(new_n16322_), .A2(new_n16312_), .A3(pi0759), .ZN(new_n16323_));
  AOI21_X1   g13887(.A1(new_n16323_), .A2(new_n16302_), .B(pi0038), .ZN(new_n16324_));
  INV_X1     g13888(.I(pi0696), .ZN(new_n16325_));
  OAI21_X1   g13889(.A1(new_n13397_), .A2(new_n16297_), .B(pi0038), .ZN(new_n16326_));
  NOR2_X1    g13890(.A1(new_n13004_), .A2(pi0152), .ZN(new_n16327_));
  OAI21_X1   g13891(.A1(new_n16327_), .A2(new_n16326_), .B(new_n16325_), .ZN(new_n16328_));
  AOI21_X1   g13892(.A1(new_n16324_), .A2(new_n16300_), .B(new_n16328_), .ZN(new_n16329_));
  AOI21_X1   g13893(.A1(new_n3369_), .A2(new_n16253_), .B(new_n16106_), .ZN(new_n16330_));
  NAND2_X1   g13894(.A1(new_n16056_), .A2(new_n15994_), .ZN(new_n16331_));
  NAND2_X1   g13895(.A1(new_n16330_), .A2(new_n16331_), .ZN(new_n16332_));
  INV_X1     g13896(.I(new_n16007_), .ZN(new_n16333_));
  AOI21_X1   g13897(.A1(new_n16059_), .A2(new_n16308_), .B(pi0215), .ZN(new_n16334_));
  NAND3_X1   g13898(.A1(new_n16305_), .A2(new_n16333_), .A3(new_n16334_), .ZN(new_n16335_));
  NAND3_X1   g13899(.A1(new_n16335_), .A2(new_n16332_), .A3(pi0299), .ZN(new_n16336_));
  NAND2_X1   g13900(.A1(new_n16315_), .A2(new_n15936_), .ZN(new_n16337_));
  NAND2_X1   g13901(.A1(new_n16317_), .A2(new_n16337_), .ZN(new_n16338_));
  INV_X1     g13902(.I(new_n16030_), .ZN(new_n16339_));
  AOI21_X1   g13903(.A1(new_n16339_), .A2(new_n16308_), .B(new_n2642_), .ZN(new_n16340_));
  AOI21_X1   g13904(.A1(new_n16338_), .A2(new_n2642_), .B(new_n16340_), .ZN(new_n16341_));
  AOI21_X1   g13905(.A1(new_n16320_), .A2(new_n16044_), .B(pi0299), .ZN(new_n16342_));
  OAI21_X1   g13906(.A1(new_n16341_), .A2(pi0223), .B(new_n16342_), .ZN(new_n16343_));
  NAND3_X1   g13907(.A1(new_n16336_), .A2(new_n16343_), .A3(new_n16296_), .ZN(new_n16344_));
  NAND2_X1   g13908(.A1(new_n16320_), .A2(new_n16044_), .ZN(new_n16345_));
  NAND3_X1   g13909(.A1(new_n16271_), .A2(new_n2641_), .A3(new_n16308_), .ZN(new_n16346_));
  AOI21_X1   g13910(.A1(new_n16315_), .A2(new_n5421_), .B(new_n2641_), .ZN(new_n16347_));
  INV_X1     g13911(.I(new_n16347_), .ZN(new_n16348_));
  OR2_X2     g13912(.A1(new_n16318_), .A2(new_n16348_), .Z(new_n16349_));
  NAND3_X1   g13913(.A1(new_n16349_), .A2(new_n2668_), .A3(new_n16346_), .ZN(new_n16350_));
  NAND3_X1   g13914(.A1(new_n16350_), .A2(new_n16321_), .A3(new_n16345_), .ZN(new_n16351_));
  INV_X1     g13915(.I(new_n16330_), .ZN(new_n16352_));
  OAI21_X1   g13916(.A1(new_n16305_), .A2(new_n16248_), .B(new_n16334_), .ZN(new_n16353_));
  NAND3_X1   g13917(.A1(new_n16353_), .A2(pi0299), .A3(new_n16352_), .ZN(new_n16354_));
  NAND3_X1   g13918(.A1(new_n16351_), .A2(pi0759), .A3(new_n16354_), .ZN(new_n16355_));
  NAND3_X1   g13919(.A1(new_n16355_), .A2(pi0039), .A3(new_n16344_), .ZN(new_n16356_));
  NOR2_X1    g13920(.A1(new_n16300_), .A2(new_n16023_), .ZN(new_n16357_));
  NOR2_X1    g13921(.A1(new_n16357_), .A2(pi0038), .ZN(new_n16358_));
  NAND2_X1   g13922(.A1(new_n16356_), .A2(new_n16358_), .ZN(new_n16359_));
  INV_X1     g13923(.I(new_n16297_), .ZN(new_n16360_));
  NOR3_X1    g13924(.A1(new_n13568_), .A2(pi0039), .A3(new_n15936_), .ZN(new_n16361_));
  AOI21_X1   g13925(.A1(new_n16361_), .A2(new_n16360_), .B(new_n3265_), .ZN(new_n16362_));
  NAND2_X1   g13926(.A1(new_n13397_), .A2(new_n3369_), .ZN(new_n16363_));
  AOI21_X1   g13927(.A1(new_n16363_), .A2(new_n16362_), .B(new_n16325_), .ZN(new_n16364_));
  AOI21_X1   g13928(.A1(new_n16359_), .A2(new_n16364_), .B(new_n16329_), .ZN(new_n16365_));
  NOR2_X1    g13929(.A1(new_n8264_), .A2(new_n3369_), .ZN(new_n16366_));
  AOI21_X1   g13930(.A1(new_n16365_), .A2(new_n8264_), .B(new_n16366_), .ZN(new_n16367_));
  NOR2_X1    g13931(.A1(new_n15994_), .A2(new_n16325_), .ZN(new_n16368_));
  NOR3_X1    g13932(.A1(new_n16368_), .A2(new_n3043_), .A3(new_n16297_), .ZN(new_n16369_));
  OAI21_X1   g13933(.A1(new_n3042_), .A2(pi0152), .B(pi0832), .ZN(new_n16370_));
  OAI22_X1   g13934(.A1(new_n16367_), .A2(pi0832), .B1(new_n16369_), .B2(new_n16370_), .ZN(po0309));
  OAI21_X1   g13935(.A1(new_n3042_), .A2(new_n2455_), .B(pi0832), .ZN(new_n16372_));
  AOI21_X1   g13936(.A1(pi0766), .A2(pi0947), .B(new_n3043_), .ZN(new_n16373_));
  INV_X1     g13937(.I(new_n16373_), .ZN(new_n16374_));
  AOI21_X1   g13938(.A1(pi0700), .A2(new_n15936_), .B(new_n16374_), .ZN(new_n16375_));
  OAI21_X1   g13939(.A1(new_n2582_), .A2(new_n2455_), .B(new_n12738_), .ZN(new_n16376_));
  NAND2_X1   g13940(.A1(new_n5336_), .A2(new_n16373_), .ZN(new_n16377_));
  NAND2_X1   g13941(.A1(new_n16073_), .A2(pi0153), .ZN(new_n16378_));
  NAND3_X1   g13942(.A1(new_n16378_), .A2(pi0038), .A3(new_n16377_), .ZN(new_n16379_));
  NOR2_X1    g13943(.A1(new_n13336_), .A2(pi0766), .ZN(new_n16380_));
  OAI22_X1   g13944(.A1(new_n16380_), .A2(new_n16083_), .B1(pi0153), .B2(new_n16102_), .ZN(new_n16381_));
  NOR2_X1    g13945(.A1(pi0153), .A2(pi0766), .ZN(new_n16382_));
  AOI21_X1   g13946(.A1(new_n14065_), .A2(new_n16382_), .B(new_n2627_), .ZN(new_n16383_));
  INV_X1     g13947(.I(pi0766), .ZN(new_n16384_));
  NAND2_X1   g13948(.A1(new_n16253_), .A2(pi0153), .ZN(new_n16385_));
  AOI21_X1   g13949(.A1(new_n16107_), .A2(new_n16385_), .B(new_n2628_), .ZN(new_n16386_));
  NOR2_X1    g13950(.A1(new_n16248_), .A2(new_n2455_), .ZN(new_n16387_));
  OAI21_X1   g13951(.A1(new_n16002_), .A2(new_n16387_), .B(new_n3304_), .ZN(new_n16388_));
  NAND2_X1   g13952(.A1(new_n13088_), .A2(new_n2455_), .ZN(new_n16389_));
  NAND2_X1   g13953(.A1(new_n16089_), .A2(new_n16389_), .ZN(new_n16390_));
  NAND3_X1   g13954(.A1(new_n16110_), .A2(new_n16388_), .A3(new_n16390_), .ZN(new_n16391_));
  AOI21_X1   g13955(.A1(new_n16391_), .A2(new_n16386_), .B(new_n16384_), .ZN(new_n16392_));
  NAND2_X1   g13956(.A1(new_n16015_), .A2(new_n2455_), .ZN(new_n16393_));
  NAND2_X1   g13957(.A1(new_n16086_), .A2(new_n16393_), .ZN(new_n16394_));
  NAND2_X1   g13958(.A1(new_n16394_), .A2(new_n16392_), .ZN(new_n16395_));
  AOI21_X1   g13959(.A1(new_n16395_), .A2(new_n16383_), .B(pi0038), .ZN(new_n16396_));
  AOI21_X1   g13960(.A1(new_n16396_), .A2(new_n16381_), .B(pi0700), .ZN(new_n16397_));
  AOI21_X1   g13961(.A1(new_n16397_), .A2(new_n16379_), .B(new_n16148_), .ZN(new_n16398_));
  AOI21_X1   g13962(.A1(new_n16384_), .A2(pi0947), .B(new_n16186_), .ZN(new_n16399_));
  OAI21_X1   g13963(.A1(new_n13344_), .A2(pi0153), .B(pi0038), .ZN(new_n16400_));
  AOI21_X1   g13964(.A1(new_n16399_), .A2(new_n2627_), .B(new_n16400_), .ZN(new_n16401_));
  NAND2_X1   g13965(.A1(new_n16393_), .A2(new_n16025_), .ZN(new_n16402_));
  INV_X1     g13966(.I(new_n16001_), .ZN(new_n16403_));
  NAND2_X1   g13967(.A1(new_n16105_), .A2(new_n16385_), .ZN(new_n16404_));
  NAND2_X1   g13968(.A1(new_n16404_), .A2(new_n13176_), .ZN(new_n16405_));
  NAND2_X1   g13969(.A1(new_n16405_), .A2(new_n16403_), .ZN(new_n16406_));
  AOI21_X1   g13970(.A1(new_n16270_), .A2(new_n16389_), .B(new_n16005_), .ZN(new_n16407_));
  AOI21_X1   g13971(.A1(new_n16407_), .A2(new_n16388_), .B(pi0215), .ZN(new_n16408_));
  OAI21_X1   g13972(.A1(new_n16408_), .A2(new_n16406_), .B(pi0299), .ZN(new_n16409_));
  NAND3_X1   g13973(.A1(new_n16409_), .A2(new_n16384_), .A3(new_n16402_), .ZN(new_n16410_));
  NOR2_X1    g13974(.A1(new_n13088_), .A2(new_n5473_), .ZN(new_n16411_));
  NOR2_X1    g13975(.A1(new_n16390_), .A2(new_n16411_), .ZN(new_n16412_));
  NOR2_X1    g13976(.A1(new_n16412_), .A2(pi0215), .ZN(new_n16413_));
  NAND2_X1   g13977(.A1(new_n16388_), .A2(new_n16413_), .ZN(new_n16414_));
  AOI21_X1   g13978(.A1(new_n16414_), .A2(new_n16404_), .B(new_n2628_), .ZN(new_n16415_));
  AOI21_X1   g13979(.A1(pi0153), .A2(new_n16055_), .B(new_n16268_), .ZN(new_n16416_));
  OAI21_X1   g13980(.A1(new_n16416_), .A2(new_n16415_), .B(pi0766), .ZN(new_n16417_));
  NAND3_X1   g13981(.A1(new_n16417_), .A2(pi0039), .A3(new_n16410_), .ZN(new_n16418_));
  OR2_X2     g13982(.A1(new_n16381_), .A2(new_n16023_), .Z(new_n16419_));
  AOI21_X1   g13983(.A1(new_n16418_), .A2(new_n16419_), .B(pi0038), .ZN(new_n16420_));
  OAI21_X1   g13984(.A1(new_n16420_), .A2(new_n16401_), .B(pi0700), .ZN(new_n16421_));
  OAI21_X1   g13985(.A1(new_n16147_), .A2(pi0153), .B(new_n2582_), .ZN(new_n16422_));
  AOI21_X1   g13986(.A1(new_n16421_), .A2(new_n16398_), .B(new_n16422_), .ZN(new_n16423_));
  OAI22_X1   g13987(.A1(new_n16423_), .A2(new_n16376_), .B1(new_n16372_), .B2(new_n16375_), .ZN(po0310));
  OAI22_X1   g13988(.A1(new_n15994_), .A2(pi0704), .B1(pi0742), .B2(new_n5692_), .ZN(new_n16425_));
  NAND2_X1   g13989(.A1(new_n3043_), .A2(pi0154), .ZN(new_n16426_));
  OAI21_X1   g13990(.A1(new_n16425_), .A2(new_n3043_), .B(new_n16426_), .ZN(new_n16427_));
  AOI21_X1   g13991(.A1(new_n8265_), .A2(new_n3321_), .B(pi0832), .ZN(new_n16428_));
  INV_X1     g13992(.I(pi0704), .ZN(new_n16429_));
  INV_X1     g13993(.I(pi0742), .ZN(new_n16430_));
  NAND2_X1   g13994(.A1(new_n13397_), .A2(new_n3321_), .ZN(new_n16431_));
  AOI21_X1   g13995(.A1(new_n16431_), .A2(new_n15999_), .B(new_n16430_), .ZN(new_n16432_));
  INV_X1     g13996(.I(new_n16024_), .ZN(new_n16433_));
  NOR2_X1    g13997(.A1(new_n16102_), .A2(pi0154), .ZN(new_n16434_));
  NOR2_X1    g13998(.A1(new_n16433_), .A2(new_n16434_), .ZN(new_n16435_));
  NAND2_X1   g13999(.A1(new_n16020_), .A2(new_n3321_), .ZN(new_n16436_));
  NAND2_X1   g14000(.A1(new_n16035_), .A2(pi0154), .ZN(new_n16437_));
  AOI21_X1   g14001(.A1(new_n16436_), .A2(new_n16437_), .B(new_n2627_), .ZN(new_n16438_));
  OAI21_X1   g14002(.A1(new_n16438_), .A2(new_n16435_), .B(new_n3265_), .ZN(new_n16439_));
  NAND2_X1   g14003(.A1(new_n16439_), .A2(new_n16432_), .ZN(new_n16440_));
  AOI21_X1   g14004(.A1(new_n16072_), .A2(new_n16431_), .B(pi0742), .ZN(new_n16441_));
  NAND2_X1   g14005(.A1(new_n16175_), .A2(pi0154), .ZN(new_n16442_));
  OAI21_X1   g14006(.A1(new_n16052_), .A2(pi0154), .B(new_n16442_), .ZN(new_n16443_));
  AOI22_X1   g14007(.A1(new_n16443_), .A2(pi0039), .B1(new_n16064_), .B2(new_n16435_), .ZN(new_n16444_));
  OAI21_X1   g14008(.A1(new_n16444_), .A2(pi0038), .B(new_n16441_), .ZN(new_n16445_));
  NAND3_X1   g14009(.A1(new_n16440_), .A2(new_n16429_), .A3(new_n16445_), .ZN(new_n16446_));
  NOR2_X1    g14010(.A1(new_n13191_), .A2(new_n16430_), .ZN(new_n16447_));
  AOI21_X1   g14011(.A1(new_n16447_), .A2(new_n3321_), .B(new_n16429_), .ZN(new_n16448_));
  OAI21_X1   g14012(.A1(pi0154), .A2(new_n13004_), .B(new_n16081_), .ZN(new_n16449_));
  NAND2_X1   g14013(.A1(new_n16095_), .A2(pi0154), .ZN(new_n16450_));
  NAND2_X1   g14014(.A1(new_n16117_), .A2(new_n3321_), .ZN(new_n16451_));
  AOI21_X1   g14015(.A1(new_n16451_), .A2(new_n16450_), .B(new_n2627_), .ZN(new_n16452_));
  NOR3_X1    g14016(.A1(new_n16434_), .A2(pi0039), .A3(new_n16082_), .ZN(new_n16453_));
  OAI21_X1   g14017(.A1(new_n16452_), .A2(new_n16453_), .B(new_n3265_), .ZN(new_n16454_));
  NAND3_X1   g14018(.A1(new_n16454_), .A2(new_n16430_), .A3(new_n16449_), .ZN(new_n16455_));
  NAND2_X1   g14019(.A1(new_n16455_), .A2(new_n16448_), .ZN(new_n16456_));
  NAND3_X1   g14020(.A1(new_n16456_), .A2(new_n8264_), .A3(new_n16446_), .ZN(new_n16457_));
  AOI22_X1   g14021(.A1(new_n16457_), .A2(new_n16428_), .B1(pi0832), .B2(new_n16427_), .ZN(po0311));
  INV_X1     g14022(.I(pi0686), .ZN(new_n16459_));
  INV_X1     g14023(.I(pi0757), .ZN(new_n16460_));
  AOI22_X1   g14024(.A1(new_n15936_), .A2(new_n16459_), .B1(new_n16460_), .B2(pi0947), .ZN(new_n16461_));
  NAND2_X1   g14025(.A1(new_n16461_), .A2(new_n3042_), .ZN(new_n16462_));
  NAND2_X1   g14026(.A1(new_n3043_), .A2(pi0155), .ZN(new_n16463_));
  AOI21_X1   g14027(.A1(new_n16462_), .A2(new_n16463_), .B(new_n12738_), .ZN(new_n16464_));
  OAI21_X1   g14028(.A1(new_n13190_), .A2(new_n13005_), .B(pi0757), .ZN(new_n16465_));
  OAI21_X1   g14029(.A1(new_n16119_), .A2(pi0757), .B(new_n16465_), .ZN(new_n16466_));
  NOR2_X1    g14030(.A1(new_n16466_), .A2(new_n16459_), .ZN(new_n16467_));
  NOR2_X1    g14031(.A1(new_n13397_), .A2(new_n3265_), .ZN(new_n16468_));
  INV_X1     g14032(.I(new_n16468_), .ZN(new_n16469_));
  OAI22_X1   g14033(.A1(new_n16021_), .A2(pi0038), .B1(new_n15936_), .B2(new_n16469_), .ZN(new_n16470_));
  NAND2_X1   g14034(.A1(new_n16470_), .A2(pi0757), .ZN(new_n16471_));
  NOR2_X1    g14035(.A1(new_n16053_), .A2(pi0038), .ZN(new_n16472_));
  AOI21_X1   g14036(.A1(pi0038), .A2(new_n16075_), .B(new_n16472_), .ZN(new_n16473_));
  NAND2_X1   g14037(.A1(new_n16473_), .A2(new_n16460_), .ZN(new_n16474_));
  AOI21_X1   g14038(.A1(new_n16474_), .A2(new_n16471_), .B(pi0686), .ZN(new_n16475_));
  OAI21_X1   g14039(.A1(new_n16467_), .A2(new_n16475_), .B(new_n8264_), .ZN(new_n16476_));
  OAI21_X1   g14040(.A1(new_n16067_), .A2(pi0038), .B(new_n16071_), .ZN(new_n16477_));
  NAND2_X1   g14041(.A1(new_n16477_), .A2(new_n16460_), .ZN(new_n16478_));
  INV_X1     g14042(.I(new_n16036_), .ZN(new_n16479_));
  AOI21_X1   g14043(.A1(new_n16479_), .A2(new_n3265_), .B(new_n15999_), .ZN(new_n16480_));
  INV_X1     g14044(.I(new_n16480_), .ZN(new_n16481_));
  NAND2_X1   g14045(.A1(new_n16481_), .A2(pi0757), .ZN(new_n16482_));
  AOI21_X1   g14046(.A1(new_n16482_), .A2(new_n16478_), .B(pi0686), .ZN(new_n16483_));
  INV_X1     g14047(.I(new_n16098_), .ZN(new_n16484_));
  OAI21_X1   g14048(.A1(new_n16484_), .A2(pi0757), .B(pi0686), .ZN(new_n16485_));
  NAND2_X1   g14049(.A1(new_n16485_), .A2(new_n8264_), .ZN(new_n16486_));
  OAI21_X1   g14050(.A1(new_n16486_), .A2(new_n16483_), .B(pi0155), .ZN(new_n16487_));
  OAI21_X1   g14051(.A1(new_n16476_), .A2(pi0155), .B(new_n16487_), .ZN(new_n16488_));
  AOI21_X1   g14052(.A1(new_n16488_), .A2(new_n12738_), .B(new_n16464_), .ZN(po0312));
  OAI22_X1   g14053(.A1(new_n15994_), .A2(pi0724), .B1(pi0741), .B2(new_n5692_), .ZN(new_n16490_));
  NAND2_X1   g14054(.A1(new_n3043_), .A2(pi0156), .ZN(new_n16491_));
  OAI21_X1   g14055(.A1(new_n16490_), .A2(new_n3043_), .B(new_n16491_), .ZN(new_n16492_));
  NOR2_X1    g14056(.A1(new_n16477_), .A2(pi0741), .ZN(new_n16493_));
  AOI21_X1   g14057(.A1(pi0741), .A2(new_n16480_), .B(new_n16493_), .ZN(new_n16494_));
  NAND2_X1   g14058(.A1(new_n16098_), .A2(pi0724), .ZN(new_n16495_));
  OAI22_X1   g14059(.A1(new_n16494_), .A2(pi0724), .B1(pi0741), .B2(new_n16495_), .ZN(new_n16496_));
  NOR2_X1    g14060(.A1(new_n8265_), .A2(new_n9471_), .ZN(new_n16497_));
  AOI21_X1   g14061(.A1(new_n16496_), .A2(new_n16497_), .B(pi0832), .ZN(new_n16498_));
  INV_X1     g14062(.I(pi0724), .ZN(new_n16499_));
  INV_X1     g14063(.I(pi0741), .ZN(new_n16500_));
  NOR2_X1    g14064(.A1(new_n16470_), .A2(new_n16500_), .ZN(new_n16501_));
  NOR2_X1    g14065(.A1(new_n16473_), .A2(pi0741), .ZN(new_n16502_));
  OAI21_X1   g14066(.A1(new_n16502_), .A2(new_n16501_), .B(new_n16499_), .ZN(new_n16503_));
  NOR3_X1    g14067(.A1(new_n13190_), .A2(new_n16500_), .A3(new_n13005_), .ZN(new_n16504_));
  AOI21_X1   g14068(.A1(new_n16119_), .A2(new_n16500_), .B(new_n16504_), .ZN(new_n16505_));
  NAND2_X1   g14069(.A1(new_n16505_), .A2(pi0724), .ZN(new_n16506_));
  NAND3_X1   g14070(.A1(new_n16506_), .A2(new_n8264_), .A3(new_n16503_), .ZN(new_n16507_));
  NAND2_X1   g14071(.A1(new_n16507_), .A2(new_n9471_), .ZN(new_n16508_));
  AOI22_X1   g14072(.A1(new_n16508_), .A2(new_n16498_), .B1(pi0832), .B2(new_n16492_), .ZN(po0313));
  INV_X1     g14073(.I(pi0688), .ZN(new_n16510_));
  NOR2_X1    g14074(.A1(new_n16051_), .A2(pi0760), .ZN(new_n16511_));
  INV_X1     g14075(.I(pi0760), .ZN(new_n16512_));
  NOR2_X1    g14076(.A1(new_n16020_), .A2(new_n16512_), .ZN(new_n16513_));
  OAI21_X1   g14077(.A1(new_n16513_), .A2(new_n16511_), .B(new_n10834_), .ZN(new_n16514_));
  NOR2_X1    g14078(.A1(new_n16175_), .A2(pi0760), .ZN(new_n16515_));
  NOR2_X1    g14079(.A1(new_n16035_), .A2(new_n16512_), .ZN(new_n16516_));
  OAI21_X1   g14080(.A1(new_n16515_), .A2(new_n16516_), .B(pi0157), .ZN(new_n16517_));
  NAND3_X1   g14081(.A1(new_n16514_), .A2(pi0039), .A3(new_n16517_), .ZN(new_n16518_));
  INV_X1     g14082(.I(new_n16023_), .ZN(new_n16519_));
  NOR2_X1    g14083(.A1(new_n5692_), .A2(pi0760), .ZN(new_n16520_));
  INV_X1     g14084(.I(new_n16520_), .ZN(new_n16521_));
  NAND2_X1   g14085(.A1(new_n16102_), .A2(new_n16521_), .ZN(new_n16522_));
  NAND2_X1   g14086(.A1(new_n13060_), .A2(pi0157), .ZN(new_n16523_));
  AOI21_X1   g14087(.A1(new_n16522_), .A2(new_n16523_), .B(pi0039), .ZN(new_n16524_));
  NAND2_X1   g14088(.A1(new_n16524_), .A2(new_n16519_), .ZN(new_n16525_));
  AOI21_X1   g14089(.A1(new_n16518_), .A2(new_n16525_), .B(pi0038), .ZN(new_n16526_));
  NOR2_X1    g14090(.A1(new_n16512_), .A2(new_n5692_), .ZN(new_n16527_));
  NOR3_X1    g14091(.A1(new_n16186_), .A2(pi0039), .A3(new_n16527_), .ZN(new_n16528_));
  OAI21_X1   g14092(.A1(new_n13344_), .A2(pi0157), .B(pi0038), .ZN(new_n16529_));
  OAI21_X1   g14093(.A1(new_n16528_), .A2(new_n16529_), .B(new_n16510_), .ZN(new_n16530_));
  OAI21_X1   g14094(.A1(new_n13397_), .A2(new_n16520_), .B(pi0038), .ZN(new_n16531_));
  AOI21_X1   g14095(.A1(new_n16073_), .A2(pi0157), .B(new_n16531_), .ZN(new_n16532_));
  NAND2_X1   g14096(.A1(new_n10834_), .A2(pi0760), .ZN(new_n16533_));
  OAI21_X1   g14097(.A1(new_n14064_), .A2(new_n16533_), .B(pi0039), .ZN(new_n16534_));
  OAI21_X1   g14098(.A1(pi0157), .A2(new_n16014_), .B(new_n16086_), .ZN(new_n16535_));
  NAND2_X1   g14099(.A1(new_n16114_), .A2(new_n10834_), .ZN(new_n16536_));
  OAI22_X1   g14100(.A1(new_n16092_), .A2(new_n16090_), .B1(pi0157), .B2(new_n2628_), .ZN(new_n16537_));
  AOI21_X1   g14101(.A1(new_n16536_), .A2(new_n16537_), .B(pi0760), .ZN(new_n16538_));
  AOI21_X1   g14102(.A1(new_n16538_), .A2(new_n16535_), .B(new_n16534_), .ZN(new_n16539_));
  NOR3_X1    g14103(.A1(new_n16539_), .A2(pi0038), .A3(new_n16524_), .ZN(new_n16540_));
  NOR2_X1    g14104(.A1(new_n16540_), .A2(new_n16532_), .ZN(new_n16541_));
  OAI22_X1   g14105(.A1(new_n16526_), .A2(new_n16530_), .B1(new_n16541_), .B2(new_n16510_), .ZN(new_n16542_));
  NAND2_X1   g14106(.A1(new_n8265_), .A2(pi0157), .ZN(new_n16543_));
  OAI21_X1   g14107(.A1(new_n16542_), .A2(new_n8265_), .B(new_n16543_), .ZN(new_n16544_));
  NAND2_X1   g14108(.A1(new_n15936_), .A2(new_n16510_), .ZN(new_n16545_));
  NAND3_X1   g14109(.A1(new_n16545_), .A2(new_n16521_), .A3(new_n3042_), .ZN(new_n16546_));
  NAND2_X1   g14110(.A1(new_n3043_), .A2(pi0157), .ZN(new_n16547_));
  AOI21_X1   g14111(.A1(new_n16546_), .A2(new_n16547_), .B(new_n12738_), .ZN(new_n16548_));
  AOI21_X1   g14112(.A1(new_n16544_), .A2(new_n12738_), .B(new_n16548_), .ZN(po0314));
  INV_X1     g14113(.I(pi0753), .ZN(new_n16550_));
  NOR2_X1    g14114(.A1(new_n16102_), .A2(pi0158), .ZN(new_n16551_));
  AOI21_X1   g14115(.A1(new_n16550_), .A2(new_n16102_), .B(new_n16551_), .ZN(new_n16552_));
  NAND2_X1   g14116(.A1(new_n16094_), .A2(pi0158), .ZN(new_n16553_));
  OAI21_X1   g14117(.A1(new_n16117_), .A2(pi0158), .B(new_n16553_), .ZN(new_n16554_));
  NOR2_X1    g14118(.A1(new_n16550_), .A2(pi0158), .ZN(new_n16555_));
  AOI22_X1   g14119(.A1(new_n16554_), .A2(new_n16550_), .B1(new_n14065_), .B2(new_n16555_), .ZN(new_n16556_));
  OAI22_X1   g14120(.A1(new_n16556_), .A2(new_n2627_), .B1(new_n16104_), .B2(new_n16552_), .ZN(new_n16557_));
  INV_X1     g14121(.I(pi0702), .ZN(new_n16558_));
  NOR2_X1    g14122(.A1(new_n5692_), .A2(pi0753), .ZN(new_n16559_));
  OAI22_X1   g14123(.A1(new_n13004_), .A2(new_n5631_), .B1(new_n13397_), .B2(new_n16559_), .ZN(new_n16560_));
  AOI21_X1   g14124(.A1(new_n16560_), .A2(pi0038), .B(new_n16558_), .ZN(new_n16561_));
  OAI21_X1   g14125(.A1(new_n16557_), .A2(pi0038), .B(new_n16561_), .ZN(new_n16562_));
  NAND2_X1   g14126(.A1(new_n16052_), .A2(new_n5631_), .ZN(new_n16563_));
  NAND2_X1   g14127(.A1(new_n16062_), .A2(pi0158), .ZN(new_n16564_));
  AOI21_X1   g14128(.A1(new_n16563_), .A2(new_n16564_), .B(pi0753), .ZN(new_n16565_));
  NAND2_X1   g14129(.A1(new_n16034_), .A2(pi0158), .ZN(new_n16566_));
  NAND2_X1   g14130(.A1(new_n16019_), .A2(new_n5631_), .ZN(new_n16567_));
  AOI21_X1   g14131(.A1(new_n16567_), .A2(new_n16566_), .B(new_n16550_), .ZN(new_n16568_));
  OAI21_X1   g14132(.A1(new_n16568_), .A2(new_n16565_), .B(pi0039), .ZN(new_n16569_));
  NOR2_X1    g14133(.A1(new_n16550_), .A2(new_n5692_), .ZN(new_n16570_));
  NOR3_X1    g14134(.A1(new_n13060_), .A2(new_n5420_), .A3(new_n16570_), .ZN(new_n16571_));
  OAI21_X1   g14135(.A1(new_n16551_), .A2(new_n16571_), .B(new_n2627_), .ZN(new_n16572_));
  NAND3_X1   g14136(.A1(new_n16569_), .A2(new_n3265_), .A3(new_n16572_), .ZN(new_n16573_));
  OR3_X2     g14137(.A1(new_n16186_), .A2(pi0039), .A3(new_n16570_), .Z(new_n16574_));
  AOI21_X1   g14138(.A1(new_n13397_), .A2(new_n5631_), .B(new_n3265_), .ZN(new_n16575_));
  AOI21_X1   g14139(.A1(new_n16574_), .A2(new_n16575_), .B(pi0702), .ZN(new_n16576_));
  NAND2_X1   g14140(.A1(new_n16573_), .A2(new_n16576_), .ZN(new_n16577_));
  NAND3_X1   g14141(.A1(new_n16562_), .A2(new_n8264_), .A3(new_n16577_), .ZN(new_n16578_));
  OAI21_X1   g14142(.A1(new_n5631_), .A2(new_n8264_), .B(new_n16578_), .ZN(new_n16579_));
  AOI21_X1   g14143(.A1(new_n16558_), .A2(new_n15936_), .B(new_n16559_), .ZN(new_n16580_));
  NAND2_X1   g14144(.A1(new_n16580_), .A2(new_n3042_), .ZN(new_n16581_));
  NAND2_X1   g14145(.A1(new_n3043_), .A2(pi0158), .ZN(new_n16582_));
  AOI21_X1   g14146(.A1(new_n16581_), .A2(new_n16582_), .B(new_n12738_), .ZN(new_n16583_));
  AOI21_X1   g14147(.A1(new_n16579_), .A2(new_n12738_), .B(new_n16583_), .ZN(po0315));
  INV_X1     g14148(.I(pi0754), .ZN(new_n16585_));
  NOR2_X1    g14149(.A1(new_n16102_), .A2(pi0159), .ZN(new_n16586_));
  AOI21_X1   g14150(.A1(new_n16585_), .A2(new_n16102_), .B(new_n16586_), .ZN(new_n16587_));
  NAND2_X1   g14151(.A1(new_n16094_), .A2(pi0159), .ZN(new_n16588_));
  OAI21_X1   g14152(.A1(new_n16117_), .A2(pi0159), .B(new_n16588_), .ZN(new_n16589_));
  NOR2_X1    g14153(.A1(new_n16585_), .A2(pi0159), .ZN(new_n16590_));
  AOI22_X1   g14154(.A1(new_n16589_), .A2(new_n16585_), .B1(new_n14065_), .B2(new_n16590_), .ZN(new_n16591_));
  OAI22_X1   g14155(.A1(new_n16591_), .A2(new_n2627_), .B1(new_n16104_), .B2(new_n16587_), .ZN(new_n16592_));
  INV_X1     g14156(.I(pi0709), .ZN(new_n16593_));
  NOR2_X1    g14157(.A1(new_n5692_), .A2(pi0754), .ZN(new_n16594_));
  OAI22_X1   g14158(.A1(new_n13004_), .A2(new_n5632_), .B1(new_n13397_), .B2(new_n16594_), .ZN(new_n16595_));
  AOI21_X1   g14159(.A1(new_n16595_), .A2(pi0038), .B(new_n16593_), .ZN(new_n16596_));
  OAI21_X1   g14160(.A1(new_n16592_), .A2(pi0038), .B(new_n16596_), .ZN(new_n16597_));
  NAND2_X1   g14161(.A1(new_n16052_), .A2(new_n5632_), .ZN(new_n16598_));
  NAND2_X1   g14162(.A1(new_n16062_), .A2(pi0159), .ZN(new_n16599_));
  AOI21_X1   g14163(.A1(new_n16598_), .A2(new_n16599_), .B(pi0754), .ZN(new_n16600_));
  NAND2_X1   g14164(.A1(new_n16034_), .A2(pi0159), .ZN(new_n16601_));
  NAND2_X1   g14165(.A1(new_n16019_), .A2(new_n5632_), .ZN(new_n16602_));
  AOI21_X1   g14166(.A1(new_n16602_), .A2(new_n16601_), .B(new_n16585_), .ZN(new_n16603_));
  OAI21_X1   g14167(.A1(new_n16603_), .A2(new_n16600_), .B(pi0039), .ZN(new_n16604_));
  NOR2_X1    g14168(.A1(new_n16585_), .A2(new_n5692_), .ZN(new_n16605_));
  NOR3_X1    g14169(.A1(new_n13060_), .A2(new_n5420_), .A3(new_n16605_), .ZN(new_n16606_));
  OAI21_X1   g14170(.A1(new_n16586_), .A2(new_n16606_), .B(new_n2627_), .ZN(new_n16607_));
  NAND3_X1   g14171(.A1(new_n16604_), .A2(new_n3265_), .A3(new_n16607_), .ZN(new_n16608_));
  OR3_X2     g14172(.A1(new_n16186_), .A2(pi0039), .A3(new_n16605_), .Z(new_n16609_));
  AOI21_X1   g14173(.A1(new_n13397_), .A2(new_n5632_), .B(new_n3265_), .ZN(new_n16610_));
  AOI21_X1   g14174(.A1(new_n16609_), .A2(new_n16610_), .B(pi0709), .ZN(new_n16611_));
  NAND2_X1   g14175(.A1(new_n16608_), .A2(new_n16611_), .ZN(new_n16612_));
  NAND3_X1   g14176(.A1(new_n16597_), .A2(new_n8264_), .A3(new_n16612_), .ZN(new_n16613_));
  OAI21_X1   g14177(.A1(new_n5632_), .A2(new_n8264_), .B(new_n16613_), .ZN(new_n16614_));
  AOI21_X1   g14178(.A1(new_n16593_), .A2(new_n15936_), .B(new_n16594_), .ZN(new_n16615_));
  NAND2_X1   g14179(.A1(new_n16615_), .A2(new_n3042_), .ZN(new_n16616_));
  NAND2_X1   g14180(.A1(new_n3043_), .A2(pi0159), .ZN(new_n16617_));
  AOI21_X1   g14181(.A1(new_n16616_), .A2(new_n16617_), .B(new_n12738_), .ZN(new_n16618_));
  AOI21_X1   g14182(.A1(new_n16614_), .A2(new_n12738_), .B(new_n16618_), .ZN(po0316));
  INV_X1     g14183(.I(pi0734), .ZN(new_n16620_));
  INV_X1     g14184(.I(pi0756), .ZN(new_n16621_));
  NOR2_X1    g14185(.A1(new_n16018_), .A2(new_n16621_), .ZN(new_n16622_));
  NOR2_X1    g14186(.A1(new_n16011_), .A2(pi0160), .ZN(new_n16623_));
  NOR2_X1    g14187(.A1(new_n16137_), .A2(new_n5635_), .ZN(new_n16624_));
  OAI21_X1   g14188(.A1(new_n16623_), .A2(new_n16624_), .B(new_n16622_), .ZN(new_n16625_));
  NOR2_X1    g14189(.A1(new_n16051_), .A2(pi0160), .ZN(new_n16626_));
  NOR2_X1    g14190(.A1(new_n16175_), .A2(new_n5635_), .ZN(new_n16627_));
  OAI21_X1   g14191(.A1(new_n16626_), .A2(new_n16627_), .B(new_n16621_), .ZN(new_n16628_));
  NAND3_X1   g14192(.A1(new_n16628_), .A2(new_n16625_), .A3(pi0039), .ZN(new_n16629_));
  NOR2_X1    g14193(.A1(new_n5692_), .A2(pi0756), .ZN(new_n16630_));
  NOR2_X1    g14194(.A1(new_n13060_), .A2(new_n16630_), .ZN(new_n16631_));
  NOR2_X1    g14195(.A1(new_n16102_), .A2(new_n5635_), .ZN(new_n16632_));
  OAI21_X1   g14196(.A1(new_n16632_), .A2(new_n16631_), .B(new_n2627_), .ZN(new_n16633_));
  OR2_X2     g14197(.A1(new_n16633_), .A2(new_n16023_), .Z(new_n16634_));
  AOI21_X1   g14198(.A1(new_n16629_), .A2(new_n16634_), .B(pi0038), .ZN(new_n16635_));
  NOR2_X1    g14199(.A1(new_n16621_), .A2(new_n5692_), .ZN(new_n16636_));
  NOR3_X1    g14200(.A1(new_n16186_), .A2(pi0039), .A3(new_n16636_), .ZN(new_n16637_));
  OAI21_X1   g14201(.A1(new_n13344_), .A2(pi0160), .B(pi0038), .ZN(new_n16638_));
  OAI21_X1   g14202(.A1(new_n16637_), .A2(new_n16638_), .B(new_n16620_), .ZN(new_n16639_));
  INV_X1     g14203(.I(new_n16630_), .ZN(new_n16640_));
  AOI21_X1   g14204(.A1(new_n13344_), .A2(new_n16640_), .B(new_n3265_), .ZN(new_n16641_));
  NAND2_X1   g14205(.A1(new_n16073_), .A2(pi0160), .ZN(new_n16642_));
  NOR2_X1    g14206(.A1(new_n16621_), .A2(pi0160), .ZN(new_n16643_));
  AOI21_X1   g14207(.A1(new_n14065_), .A2(new_n16643_), .B(new_n2627_), .ZN(new_n16644_));
  OAI21_X1   g14208(.A1(pi0160), .A2(new_n16014_), .B(new_n16086_), .ZN(new_n16645_));
  INV_X1     g14209(.I(new_n16157_), .ZN(new_n16646_));
  NOR2_X1    g14210(.A1(new_n16646_), .A2(new_n5635_), .ZN(new_n16647_));
  NOR2_X1    g14211(.A1(new_n16114_), .A2(pi0160), .ZN(new_n16648_));
  OAI21_X1   g14212(.A1(new_n16648_), .A2(new_n16647_), .B(pi0299), .ZN(new_n16649_));
  NAND3_X1   g14213(.A1(new_n16649_), .A2(new_n16621_), .A3(new_n16645_), .ZN(new_n16650_));
  AOI21_X1   g14214(.A1(new_n16650_), .A2(new_n16644_), .B(pi0038), .ZN(new_n16651_));
  AOI22_X1   g14215(.A1(new_n16651_), .A2(new_n16633_), .B1(new_n16641_), .B2(new_n16642_), .ZN(new_n16652_));
  OAI22_X1   g14216(.A1(new_n16652_), .A2(new_n16620_), .B1(new_n16635_), .B2(new_n16639_), .ZN(new_n16653_));
  NAND2_X1   g14217(.A1(new_n8265_), .A2(pi0160), .ZN(new_n16654_));
  OAI21_X1   g14218(.A1(new_n16653_), .A2(new_n8265_), .B(new_n16654_), .ZN(new_n16655_));
  NAND2_X1   g14219(.A1(new_n15936_), .A2(new_n16620_), .ZN(new_n16656_));
  NAND3_X1   g14220(.A1(new_n16656_), .A2(new_n16640_), .A3(new_n3042_), .ZN(new_n16657_));
  NAND2_X1   g14221(.A1(new_n3043_), .A2(pi0160), .ZN(new_n16658_));
  AOI21_X1   g14222(.A1(new_n16657_), .A2(new_n16658_), .B(new_n12738_), .ZN(new_n16659_));
  AOI21_X1   g14223(.A1(new_n16655_), .A2(new_n12738_), .B(new_n16659_), .ZN(po0317));
  NOR2_X1    g14224(.A1(new_n15233_), .A2(new_n5692_), .ZN(new_n16661_));
  NOR2_X1    g14225(.A1(new_n13060_), .A2(new_n16661_), .ZN(new_n16662_));
  NOR2_X1    g14226(.A1(new_n16102_), .A2(pi0161), .ZN(new_n16663_));
  OAI21_X1   g14227(.A1(new_n16663_), .A2(new_n16662_), .B(new_n2627_), .ZN(new_n16664_));
  NOR2_X1    g14228(.A1(new_n3360_), .A2(pi0758), .ZN(new_n16665_));
  AOI21_X1   g14229(.A1(new_n14065_), .A2(new_n16665_), .B(new_n2627_), .ZN(new_n16666_));
  OAI21_X1   g14230(.A1(new_n16304_), .A2(new_n3360_), .B(new_n16029_), .ZN(new_n16667_));
  AOI21_X1   g14231(.A1(new_n16667_), .A2(new_n16303_), .B(new_n16003_), .ZN(new_n16668_));
  NAND2_X1   g14232(.A1(new_n13088_), .A2(pi0161), .ZN(new_n16669_));
  NAND2_X1   g14233(.A1(new_n16307_), .A2(new_n16669_), .ZN(new_n16670_));
  OAI21_X1   g14234(.A1(new_n16670_), .A2(new_n3304_), .B(new_n2436_), .ZN(new_n16671_));
  AOI21_X1   g14235(.A1(new_n16107_), .A2(pi0161), .B(new_n16092_), .ZN(new_n16672_));
  OAI21_X1   g14236(.A1(new_n16668_), .A2(new_n16671_), .B(new_n16672_), .ZN(new_n16673_));
  NOR2_X1    g14237(.A1(new_n16315_), .A2(new_n3360_), .ZN(new_n16674_));
  INV_X1     g14238(.I(new_n16674_), .ZN(new_n16675_));
  AOI21_X1   g14239(.A1(new_n16675_), .A2(new_n16314_), .B(new_n2641_), .ZN(new_n16676_));
  AOI21_X1   g14240(.A1(new_n2641_), .A2(new_n16670_), .B(new_n16676_), .ZN(new_n16677_));
  NAND2_X1   g14241(.A1(new_n16041_), .A2(new_n3360_), .ZN(new_n16678_));
  AOI21_X1   g14242(.A1(new_n16043_), .A2(new_n16678_), .B(pi0299), .ZN(new_n16679_));
  OAI21_X1   g14243(.A1(new_n16677_), .A2(pi0223), .B(new_n16679_), .ZN(new_n16680_));
  NAND3_X1   g14244(.A1(new_n16680_), .A2(new_n16673_), .A3(pi0758), .ZN(new_n16681_));
  AOI21_X1   g14245(.A1(new_n16681_), .A2(new_n16666_), .B(pi0038), .ZN(new_n16682_));
  OAI21_X1   g14246(.A1(new_n13397_), .A2(new_n16661_), .B(pi0038), .ZN(new_n16683_));
  NOR2_X1    g14247(.A1(new_n13004_), .A2(pi0161), .ZN(new_n16684_));
  OAI21_X1   g14248(.A1(new_n16684_), .A2(new_n16683_), .B(new_n15275_), .ZN(new_n16685_));
  AOI21_X1   g14249(.A1(new_n16682_), .A2(new_n16664_), .B(new_n16685_), .ZN(new_n16686_));
  AOI21_X1   g14250(.A1(new_n3360_), .A2(new_n16253_), .B(new_n16106_), .ZN(new_n16687_));
  NAND2_X1   g14251(.A1(new_n16687_), .A2(new_n16331_), .ZN(new_n16688_));
  AOI21_X1   g14252(.A1(new_n16059_), .A2(new_n16669_), .B(pi0215), .ZN(new_n16689_));
  NAND3_X1   g14253(.A1(new_n16667_), .A2(new_n16333_), .A3(new_n16689_), .ZN(new_n16690_));
  NAND3_X1   g14254(.A1(new_n16690_), .A2(new_n16688_), .A3(pi0299), .ZN(new_n16691_));
  AOI21_X1   g14255(.A1(new_n16339_), .A2(new_n16669_), .B(new_n2642_), .ZN(new_n16692_));
  NAND2_X1   g14256(.A1(new_n16675_), .A2(new_n16337_), .ZN(new_n16693_));
  AOI21_X1   g14257(.A1(new_n16693_), .A2(new_n2642_), .B(new_n16692_), .ZN(new_n16694_));
  AOI21_X1   g14258(.A1(new_n16678_), .A2(new_n16044_), .B(pi0299), .ZN(new_n16695_));
  OAI21_X1   g14259(.A1(new_n16694_), .A2(pi0223), .B(new_n16695_), .ZN(new_n16696_));
  NAND3_X1   g14260(.A1(new_n16691_), .A2(new_n16696_), .A3(new_n15233_), .ZN(new_n16697_));
  NAND2_X1   g14261(.A1(new_n16678_), .A2(new_n16044_), .ZN(new_n16698_));
  NAND3_X1   g14262(.A1(new_n16271_), .A2(new_n2641_), .A3(new_n16669_), .ZN(new_n16699_));
  OR2_X2     g14263(.A1(new_n16676_), .A2(new_n16348_), .Z(new_n16700_));
  NAND3_X1   g14264(.A1(new_n16700_), .A2(new_n2668_), .A3(new_n16699_), .ZN(new_n16701_));
  NAND3_X1   g14265(.A1(new_n16701_), .A2(new_n16679_), .A3(new_n16698_), .ZN(new_n16702_));
  INV_X1     g14266(.I(new_n16687_), .ZN(new_n16703_));
  OAI21_X1   g14267(.A1(new_n16667_), .A2(new_n16248_), .B(new_n16689_), .ZN(new_n16704_));
  NAND3_X1   g14268(.A1(new_n16704_), .A2(pi0299), .A3(new_n16703_), .ZN(new_n16705_));
  NAND3_X1   g14269(.A1(new_n16702_), .A2(pi0758), .A3(new_n16705_), .ZN(new_n16706_));
  NAND3_X1   g14270(.A1(new_n16706_), .A2(pi0039), .A3(new_n16697_), .ZN(new_n16707_));
  NOR2_X1    g14271(.A1(new_n16664_), .A2(new_n16023_), .ZN(new_n16708_));
  NOR2_X1    g14272(.A1(new_n16708_), .A2(pi0038), .ZN(new_n16709_));
  NAND2_X1   g14273(.A1(new_n16707_), .A2(new_n16709_), .ZN(new_n16710_));
  INV_X1     g14274(.I(new_n16661_), .ZN(new_n16711_));
  AOI21_X1   g14275(.A1(new_n16361_), .A2(new_n16711_), .B(new_n3265_), .ZN(new_n16712_));
  NAND2_X1   g14276(.A1(new_n13397_), .A2(new_n3360_), .ZN(new_n16713_));
  AOI21_X1   g14277(.A1(new_n16713_), .A2(new_n16712_), .B(new_n15275_), .ZN(new_n16714_));
  AOI21_X1   g14278(.A1(new_n16710_), .A2(new_n16714_), .B(new_n16686_), .ZN(new_n16715_));
  NOR2_X1    g14279(.A1(new_n8264_), .A2(new_n3360_), .ZN(new_n16716_));
  AOI21_X1   g14280(.A1(new_n16715_), .A2(new_n8264_), .B(new_n16716_), .ZN(new_n16717_));
  NOR2_X1    g14281(.A1(new_n15994_), .A2(new_n15275_), .ZN(new_n16718_));
  NOR3_X1    g14282(.A1(new_n16718_), .A2(new_n3043_), .A3(new_n16661_), .ZN(new_n16719_));
  OAI21_X1   g14283(.A1(new_n3042_), .A2(pi0161), .B(pi0832), .ZN(new_n16720_));
  OAI22_X1   g14284(.A1(new_n16717_), .A2(pi0832), .B1(new_n16719_), .B2(new_n16720_), .ZN(po0318));
  AOI21_X1   g14285(.A1(new_n16137_), .A2(pi0162), .B(new_n12750_), .ZN(new_n16722_));
  INV_X1     g14286(.I(new_n11535_), .ZN(new_n16723_));
  NAND2_X1   g14287(.A1(new_n16020_), .A2(new_n16723_), .ZN(new_n16724_));
  NAND2_X1   g14288(.A1(new_n16062_), .A2(pi0162), .ZN(new_n16725_));
  OAI21_X1   g14289(.A1(pi0162), .A2(new_n16051_), .B(new_n16725_), .ZN(new_n16726_));
  AOI22_X1   g14290(.A1(new_n16724_), .A2(new_n16722_), .B1(new_n12750_), .B2(new_n16726_), .ZN(new_n16727_));
  NOR2_X1    g14291(.A1(new_n5692_), .A2(pi0761), .ZN(new_n16728_));
  INV_X1     g14292(.I(new_n16728_), .ZN(new_n16729_));
  NAND2_X1   g14293(.A1(new_n16102_), .A2(new_n16729_), .ZN(new_n16730_));
  NAND2_X1   g14294(.A1(new_n13060_), .A2(pi0162), .ZN(new_n16731_));
  AOI21_X1   g14295(.A1(new_n16730_), .A2(new_n16731_), .B(pi0039), .ZN(new_n16732_));
  AOI22_X1   g14296(.A1(new_n16727_), .A2(pi0039), .B1(new_n16519_), .B2(new_n16732_), .ZN(new_n16733_));
  NAND2_X1   g14297(.A1(pi0761), .A2(pi0947), .ZN(new_n16734_));
  NAND3_X1   g14298(.A1(new_n16185_), .A2(new_n2627_), .A3(new_n16734_), .ZN(new_n16735_));
  AOI21_X1   g14299(.A1(new_n13397_), .A2(new_n7985_), .B(new_n3265_), .ZN(new_n16736_));
  AOI21_X1   g14300(.A1(new_n16736_), .A2(new_n16735_), .B(pi0738), .ZN(new_n16737_));
  OAI21_X1   g14301(.A1(new_n16733_), .A2(pi0038), .B(new_n16737_), .ZN(new_n16738_));
  OAI21_X1   g14302(.A1(new_n13397_), .A2(new_n16728_), .B(pi0038), .ZN(new_n16739_));
  AOI21_X1   g14303(.A1(new_n16073_), .A2(pi0162), .B(new_n16739_), .ZN(new_n16740_));
  NAND3_X1   g14304(.A1(new_n16116_), .A2(new_n12750_), .A3(new_n16017_), .ZN(new_n16741_));
  OAI21_X1   g14305(.A1(new_n12750_), .A2(new_n14064_), .B(new_n16741_), .ZN(new_n16742_));
  OAI22_X1   g14306(.A1(new_n16084_), .A2(pi0299), .B1(new_n16723_), .B2(new_n16157_), .ZN(new_n16743_));
  NAND2_X1   g14307(.A1(new_n16743_), .A2(new_n12750_), .ZN(new_n16744_));
  NAND2_X1   g14308(.A1(new_n16744_), .A2(pi0039), .ZN(new_n16745_));
  AOI21_X1   g14309(.A1(new_n16742_), .A2(new_n7985_), .B(new_n16745_), .ZN(new_n16746_));
  NOR3_X1    g14310(.A1(new_n16746_), .A2(pi0038), .A3(new_n16732_), .ZN(new_n16747_));
  OAI21_X1   g14311(.A1(new_n16747_), .A2(new_n16740_), .B(pi0738), .ZN(new_n16748_));
  NAND3_X1   g14312(.A1(new_n16748_), .A2(new_n8264_), .A3(new_n16738_), .ZN(new_n16749_));
  OAI21_X1   g14313(.A1(new_n7985_), .A2(new_n8264_), .B(new_n16749_), .ZN(new_n16750_));
  NAND2_X1   g14314(.A1(new_n15936_), .A2(new_n12820_), .ZN(new_n16751_));
  NAND3_X1   g14315(.A1(new_n16751_), .A2(new_n16729_), .A3(new_n3042_), .ZN(new_n16752_));
  NAND2_X1   g14316(.A1(new_n3043_), .A2(pi0162), .ZN(new_n16753_));
  AOI21_X1   g14317(.A1(new_n16752_), .A2(new_n16753_), .B(new_n12738_), .ZN(new_n16754_));
  AOI21_X1   g14318(.A1(new_n16750_), .A2(new_n12738_), .B(new_n16754_), .ZN(po0319));
  INV_X1     g14319(.I(pi0737), .ZN(new_n16756_));
  INV_X1     g14320(.I(pi0777), .ZN(new_n16757_));
  NOR2_X1    g14321(.A1(new_n16018_), .A2(new_n16757_), .ZN(new_n16758_));
  NOR2_X1    g14322(.A1(new_n16011_), .A2(pi0163), .ZN(new_n16759_));
  NOR2_X1    g14323(.A1(new_n16137_), .A2(new_n9392_), .ZN(new_n16760_));
  OAI21_X1   g14324(.A1(new_n16759_), .A2(new_n16760_), .B(new_n16758_), .ZN(new_n16761_));
  NOR2_X1    g14325(.A1(new_n16051_), .A2(pi0163), .ZN(new_n16762_));
  NOR2_X1    g14326(.A1(new_n16175_), .A2(new_n9392_), .ZN(new_n16763_));
  OAI21_X1   g14327(.A1(new_n16762_), .A2(new_n16763_), .B(new_n16757_), .ZN(new_n16764_));
  NAND3_X1   g14328(.A1(new_n16764_), .A2(new_n16761_), .A3(pi0039), .ZN(new_n16765_));
  NOR2_X1    g14329(.A1(new_n5692_), .A2(pi0777), .ZN(new_n16766_));
  NOR2_X1    g14330(.A1(new_n13060_), .A2(new_n16766_), .ZN(new_n16767_));
  NOR2_X1    g14331(.A1(new_n16102_), .A2(new_n9392_), .ZN(new_n16768_));
  OAI21_X1   g14332(.A1(new_n16768_), .A2(new_n16767_), .B(new_n2627_), .ZN(new_n16769_));
  OR2_X2     g14333(.A1(new_n16769_), .A2(new_n16023_), .Z(new_n16770_));
  AOI21_X1   g14334(.A1(new_n16765_), .A2(new_n16770_), .B(pi0038), .ZN(new_n16771_));
  NOR2_X1    g14335(.A1(new_n16757_), .A2(new_n5692_), .ZN(new_n16772_));
  NOR3_X1    g14336(.A1(new_n16186_), .A2(pi0039), .A3(new_n16772_), .ZN(new_n16773_));
  OAI21_X1   g14337(.A1(new_n13344_), .A2(pi0163), .B(pi0038), .ZN(new_n16774_));
  OAI21_X1   g14338(.A1(new_n16773_), .A2(new_n16774_), .B(new_n16756_), .ZN(new_n16775_));
  INV_X1     g14339(.I(new_n16766_), .ZN(new_n16776_));
  AOI21_X1   g14340(.A1(new_n13344_), .A2(new_n16776_), .B(new_n3265_), .ZN(new_n16777_));
  NAND2_X1   g14341(.A1(new_n16073_), .A2(pi0163), .ZN(new_n16778_));
  NOR2_X1    g14342(.A1(new_n16757_), .A2(pi0163), .ZN(new_n16779_));
  AOI21_X1   g14343(.A1(new_n14065_), .A2(new_n16779_), .B(new_n2627_), .ZN(new_n16780_));
  OAI21_X1   g14344(.A1(pi0163), .A2(new_n16014_), .B(new_n16086_), .ZN(new_n16781_));
  OAI21_X1   g14345(.A1(new_n16113_), .A2(pi0163), .B(new_n16093_), .ZN(new_n16782_));
  NAND2_X1   g14346(.A1(new_n16115_), .A2(new_n9392_), .ZN(new_n16783_));
  NAND4_X1   g14347(.A1(new_n16783_), .A2(new_n16757_), .A3(new_n16781_), .A4(new_n16782_), .ZN(new_n16784_));
  AOI21_X1   g14348(.A1(new_n16784_), .A2(new_n16780_), .B(pi0038), .ZN(new_n16785_));
  AOI22_X1   g14349(.A1(new_n16785_), .A2(new_n16769_), .B1(new_n16777_), .B2(new_n16778_), .ZN(new_n16786_));
  OAI22_X1   g14350(.A1(new_n16786_), .A2(new_n16756_), .B1(new_n16771_), .B2(new_n16775_), .ZN(new_n16787_));
  NAND2_X1   g14351(.A1(new_n8265_), .A2(pi0163), .ZN(new_n16788_));
  OAI21_X1   g14352(.A1(new_n16787_), .A2(new_n8265_), .B(new_n16788_), .ZN(new_n16789_));
  NAND2_X1   g14353(.A1(new_n15936_), .A2(new_n16756_), .ZN(new_n16790_));
  NAND3_X1   g14354(.A1(new_n16790_), .A2(new_n16776_), .A3(new_n3042_), .ZN(new_n16791_));
  NAND2_X1   g14355(.A1(new_n3043_), .A2(pi0163), .ZN(new_n16792_));
  AOI21_X1   g14356(.A1(new_n16791_), .A2(new_n16792_), .B(new_n12738_), .ZN(new_n16793_));
  AOI21_X1   g14357(.A1(new_n16789_), .A2(new_n12738_), .B(new_n16793_), .ZN(po0320));
  INV_X1     g14358(.I(pi0703), .ZN(new_n16795_));
  AOI21_X1   g14359(.A1(new_n16101_), .A2(pi0164), .B(pi0752), .ZN(new_n16796_));
  NAND2_X1   g14360(.A1(new_n16119_), .A2(new_n16796_), .ZN(new_n16797_));
  NAND2_X1   g14361(.A1(new_n13191_), .A2(pi0752), .ZN(new_n16798_));
  OAI21_X1   g14362(.A1(new_n16484_), .A2(pi0752), .B(pi0164), .ZN(new_n16799_));
  NAND4_X1   g14363(.A1(new_n16797_), .A2(new_n16795_), .A3(new_n16798_), .A4(new_n16799_), .ZN(new_n16800_));
  NAND2_X1   g14364(.A1(new_n16053_), .A2(new_n7359_), .ZN(new_n16801_));
  OAI21_X1   g14365(.A1(new_n16067_), .A2(new_n7359_), .B(new_n16801_), .ZN(new_n16802_));
  INV_X1     g14366(.I(pi0752), .ZN(new_n16803_));
  OAI21_X1   g14367(.A1(new_n16074_), .A2(pi0164), .B(new_n16072_), .ZN(new_n16804_));
  NAND2_X1   g14368(.A1(new_n16804_), .A2(new_n16803_), .ZN(new_n16805_));
  AOI21_X1   g14369(.A1(new_n16802_), .A2(new_n3265_), .B(new_n16805_), .ZN(new_n16806_));
  NAND2_X1   g14370(.A1(new_n16479_), .A2(pi0164), .ZN(new_n16807_));
  OAI21_X1   g14371(.A1(new_n16021_), .A2(pi0164), .B(new_n16807_), .ZN(new_n16808_));
  INV_X1     g14372(.I(new_n15999_), .ZN(new_n16809_));
  NOR2_X1    g14373(.A1(new_n13344_), .A2(pi0164), .ZN(new_n16810_));
  OAI21_X1   g14374(.A1(new_n16809_), .A2(new_n16810_), .B(pi0752), .ZN(new_n16811_));
  AOI21_X1   g14375(.A1(new_n16808_), .A2(new_n3265_), .B(new_n16811_), .ZN(new_n16812_));
  OAI21_X1   g14376(.A1(new_n16806_), .A2(new_n16812_), .B(pi0703), .ZN(new_n16813_));
  NAND3_X1   g14377(.A1(new_n16800_), .A2(new_n8264_), .A3(new_n16813_), .ZN(new_n16814_));
  OAI21_X1   g14378(.A1(new_n7359_), .A2(new_n8264_), .B(new_n16814_), .ZN(new_n16815_));
  AOI22_X1   g14379(.A1(new_n15936_), .A2(pi0703), .B1(new_n16803_), .B2(pi0947), .ZN(new_n16816_));
  NAND2_X1   g14380(.A1(new_n16816_), .A2(new_n3042_), .ZN(new_n16817_));
  NAND2_X1   g14381(.A1(new_n3043_), .A2(pi0164), .ZN(new_n16818_));
  AOI21_X1   g14382(.A1(new_n16817_), .A2(new_n16818_), .B(new_n12738_), .ZN(new_n16819_));
  AOI21_X1   g14383(.A1(new_n16815_), .A2(new_n12738_), .B(new_n16819_), .ZN(po0321));
  AOI21_X1   g14384(.A1(new_n16101_), .A2(pi0165), .B(pi0774), .ZN(new_n16821_));
  NAND2_X1   g14385(.A1(new_n16119_), .A2(new_n16821_), .ZN(new_n16822_));
  NAND2_X1   g14386(.A1(new_n13191_), .A2(pi0774), .ZN(new_n16823_));
  OAI21_X1   g14387(.A1(new_n16484_), .A2(pi0774), .B(pi0165), .ZN(new_n16824_));
  NAND4_X1   g14388(.A1(new_n16822_), .A2(new_n14885_), .A3(new_n16823_), .A4(new_n16824_), .ZN(new_n16825_));
  NAND2_X1   g14389(.A1(new_n16053_), .A2(new_n10665_), .ZN(new_n16826_));
  OAI21_X1   g14390(.A1(new_n16067_), .A2(new_n10665_), .B(new_n16826_), .ZN(new_n16827_));
  OAI21_X1   g14391(.A1(new_n16074_), .A2(pi0165), .B(new_n16072_), .ZN(new_n16828_));
  NAND2_X1   g14392(.A1(new_n16828_), .A2(new_n14851_), .ZN(new_n16829_));
  AOI21_X1   g14393(.A1(new_n16827_), .A2(new_n3265_), .B(new_n16829_), .ZN(new_n16830_));
  NAND2_X1   g14394(.A1(new_n16479_), .A2(pi0165), .ZN(new_n16831_));
  OAI21_X1   g14395(.A1(new_n16021_), .A2(pi0165), .B(new_n16831_), .ZN(new_n16832_));
  NOR2_X1    g14396(.A1(new_n13344_), .A2(pi0165), .ZN(new_n16833_));
  OAI21_X1   g14397(.A1(new_n16809_), .A2(new_n16833_), .B(pi0774), .ZN(new_n16834_));
  AOI21_X1   g14398(.A1(new_n16832_), .A2(new_n3265_), .B(new_n16834_), .ZN(new_n16835_));
  OAI21_X1   g14399(.A1(new_n16830_), .A2(new_n16835_), .B(pi0687), .ZN(new_n16836_));
  NAND3_X1   g14400(.A1(new_n16825_), .A2(new_n8264_), .A3(new_n16836_), .ZN(new_n16837_));
  OAI21_X1   g14401(.A1(new_n10665_), .A2(new_n8264_), .B(new_n16837_), .ZN(new_n16838_));
  AOI22_X1   g14402(.A1(new_n15936_), .A2(pi0687), .B1(new_n14851_), .B2(pi0947), .ZN(new_n16839_));
  NAND2_X1   g14403(.A1(new_n16839_), .A2(new_n3042_), .ZN(new_n16840_));
  NAND2_X1   g14404(.A1(new_n3043_), .A2(pi0165), .ZN(new_n16841_));
  AOI21_X1   g14405(.A1(new_n16840_), .A2(new_n16841_), .B(new_n12738_), .ZN(new_n16842_));
  AOI21_X1   g14406(.A1(new_n16838_), .A2(new_n12738_), .B(new_n16842_), .ZN(po0322));
  INV_X1     g14407(.I(pi0727), .ZN(new_n16844_));
  INV_X1     g14408(.I(pi0772), .ZN(new_n16845_));
  NOR2_X1    g14409(.A1(new_n16845_), .A2(new_n5692_), .ZN(new_n16846_));
  OAI21_X1   g14410(.A1(new_n13397_), .A2(new_n16846_), .B(pi0038), .ZN(new_n16847_));
  NOR2_X1    g14411(.A1(new_n13004_), .A2(pi0166), .ZN(new_n16848_));
  OAI21_X1   g14412(.A1(new_n16848_), .A2(new_n16847_), .B(new_n16844_), .ZN(new_n16849_));
  NOR2_X1    g14413(.A1(new_n13060_), .A2(new_n16846_), .ZN(new_n16850_));
  NOR2_X1    g14414(.A1(new_n16102_), .A2(pi0166), .ZN(new_n16851_));
  OAI21_X1   g14415(.A1(new_n16851_), .A2(new_n16850_), .B(new_n2627_), .ZN(new_n16852_));
  NOR2_X1    g14416(.A1(new_n3361_), .A2(pi0772), .ZN(new_n16853_));
  AOI21_X1   g14417(.A1(new_n14065_), .A2(new_n16853_), .B(new_n2627_), .ZN(new_n16854_));
  NAND2_X1   g14418(.A1(new_n16041_), .A2(new_n3361_), .ZN(new_n16855_));
  AOI21_X1   g14419(.A1(new_n16043_), .A2(new_n16855_), .B(pi0299), .ZN(new_n16856_));
  NAND2_X1   g14420(.A1(new_n13184_), .A2(pi0166), .ZN(new_n16857_));
  AOI21_X1   g14421(.A1(new_n16314_), .A2(new_n16857_), .B(new_n2641_), .ZN(new_n16858_));
  NOR2_X1    g14422(.A1(new_n13098_), .A2(pi0166), .ZN(new_n16859_));
  AOI21_X1   g14423(.A1(new_n5692_), .A2(new_n13098_), .B(new_n16859_), .ZN(new_n16860_));
  AOI21_X1   g14424(.A1(new_n2641_), .A2(new_n16860_), .B(new_n16858_), .ZN(new_n16861_));
  OAI21_X1   g14425(.A1(new_n16861_), .A2(pi0223), .B(new_n16856_), .ZN(new_n16862_));
  OAI21_X1   g14426(.A1(new_n16304_), .A2(new_n3361_), .B(new_n16029_), .ZN(new_n16863_));
  AOI21_X1   g14427(.A1(new_n16863_), .A2(new_n16303_), .B(new_n16003_), .ZN(new_n16864_));
  OAI21_X1   g14428(.A1(new_n16860_), .A2(new_n3304_), .B(new_n2436_), .ZN(new_n16865_));
  AOI21_X1   g14429(.A1(new_n16107_), .A2(pi0166), .B(new_n16092_), .ZN(new_n16866_));
  OAI21_X1   g14430(.A1(new_n16864_), .A2(new_n16865_), .B(new_n16866_), .ZN(new_n16867_));
  NAND3_X1   g14431(.A1(new_n16867_), .A2(pi0772), .A3(new_n16862_), .ZN(new_n16868_));
  AOI21_X1   g14432(.A1(new_n16868_), .A2(new_n16854_), .B(pi0038), .ZN(new_n16869_));
  AOI21_X1   g14433(.A1(new_n16869_), .A2(new_n16852_), .B(new_n16849_), .ZN(new_n16870_));
  OAI21_X1   g14434(.A1(new_n16041_), .A2(new_n5420_), .B(new_n3361_), .ZN(new_n16871_));
  NAND2_X1   g14435(.A1(new_n16871_), .A2(new_n16044_), .ZN(new_n16872_));
  AOI21_X1   g14436(.A1(new_n5420_), .A2(new_n13098_), .B(new_n16859_), .ZN(new_n16873_));
  INV_X1     g14437(.I(new_n16873_), .ZN(new_n16874_));
  AOI21_X1   g14438(.A1(new_n16874_), .A2(new_n2641_), .B(pi0223), .ZN(new_n16875_));
  INV_X1     g14439(.I(new_n16875_), .ZN(new_n16876_));
  AOI21_X1   g14440(.A1(new_n2641_), .A2(new_n16088_), .B(new_n16876_), .ZN(new_n16877_));
  NAND2_X1   g14441(.A1(new_n16337_), .A2(new_n16857_), .ZN(new_n16878_));
  OAI21_X1   g14442(.A1(new_n16878_), .A2(new_n2641_), .B(new_n16877_), .ZN(new_n16879_));
  NAND3_X1   g14443(.A1(new_n16879_), .A2(new_n2628_), .A3(new_n16872_), .ZN(new_n16880_));
  AOI21_X1   g14444(.A1(new_n3361_), .A2(new_n16253_), .B(new_n16106_), .ZN(new_n16881_));
  NAND2_X1   g14445(.A1(new_n16881_), .A2(new_n16331_), .ZN(new_n16882_));
  AOI21_X1   g14446(.A1(new_n16874_), .A2(new_n3303_), .B(pi0215), .ZN(new_n16883_));
  NAND3_X1   g14447(.A1(new_n16863_), .A2(new_n16333_), .A3(new_n16883_), .ZN(new_n16884_));
  NAND3_X1   g14448(.A1(new_n16884_), .A2(new_n16882_), .A3(pi0299), .ZN(new_n16885_));
  NAND3_X1   g14449(.A1(new_n16885_), .A2(new_n16845_), .A3(new_n16880_), .ZN(new_n16886_));
  INV_X1     g14450(.I(new_n16881_), .ZN(new_n16887_));
  OAI21_X1   g14451(.A1(new_n16863_), .A2(new_n16248_), .B(new_n16883_), .ZN(new_n16888_));
  NAND3_X1   g14452(.A1(new_n16888_), .A2(pi0299), .A3(new_n16887_), .ZN(new_n16889_));
  OAI21_X1   g14453(.A1(new_n16348_), .A2(new_n16878_), .B(new_n16875_), .ZN(new_n16890_));
  NAND3_X1   g14454(.A1(new_n16856_), .A2(new_n16890_), .A3(new_n16872_), .ZN(new_n16891_));
  NAND3_X1   g14455(.A1(new_n16889_), .A2(pi0772), .A3(new_n16891_), .ZN(new_n16892_));
  NAND3_X1   g14456(.A1(new_n16892_), .A2(new_n16886_), .A3(pi0039), .ZN(new_n16893_));
  NOR2_X1    g14457(.A1(new_n16852_), .A2(new_n16023_), .ZN(new_n16894_));
  NOR2_X1    g14458(.A1(new_n16894_), .A2(pi0038), .ZN(new_n16895_));
  OAI21_X1   g14459(.A1(new_n13344_), .A2(pi0166), .B(pi0038), .ZN(new_n16896_));
  NOR4_X1    g14460(.A1(new_n13568_), .A2(pi0039), .A3(new_n15936_), .A4(new_n16846_), .ZN(new_n16897_));
  OAI21_X1   g14461(.A1(new_n16896_), .A2(new_n16897_), .B(pi0727), .ZN(new_n16898_));
  AOI21_X1   g14462(.A1(new_n16893_), .A2(new_n16895_), .B(new_n16898_), .ZN(new_n16899_));
  NOR3_X1    g14463(.A1(new_n16899_), .A2(new_n16870_), .A3(new_n8265_), .ZN(new_n16900_));
  AOI21_X1   g14464(.A1(pi0166), .A2(new_n8265_), .B(new_n16900_), .ZN(new_n16901_));
  OAI21_X1   g14465(.A1(new_n15994_), .A2(new_n16844_), .B(new_n3042_), .ZN(new_n16902_));
  NOR2_X1    g14466(.A1(new_n16902_), .A2(new_n16846_), .ZN(new_n16903_));
  OAI21_X1   g14467(.A1(new_n3042_), .A2(pi0166), .B(pi0832), .ZN(new_n16904_));
  OAI22_X1   g14468(.A1(new_n16901_), .A2(pi0832), .B1(new_n16903_), .B2(new_n16904_), .ZN(po0323));
  INV_X1     g14469(.I(pi0705), .ZN(new_n16906_));
  OAI22_X1   g14470(.A1(new_n15994_), .A2(new_n16906_), .B1(pi0768), .B2(new_n5692_), .ZN(new_n16907_));
  NAND2_X1   g14471(.A1(new_n3043_), .A2(pi0167), .ZN(new_n16908_));
  OAI21_X1   g14472(.A1(new_n16907_), .A2(new_n3043_), .B(new_n16908_), .ZN(new_n16909_));
  AOI21_X1   g14473(.A1(new_n8265_), .A2(new_n7925_), .B(pi0832), .ZN(new_n16910_));
  AOI21_X1   g14474(.A1(new_n16075_), .A2(new_n7925_), .B(new_n16071_), .ZN(new_n16911_));
  INV_X1     g14475(.I(pi0768), .ZN(new_n16912_));
  NOR2_X1    g14476(.A1(new_n16067_), .A2(new_n7925_), .ZN(new_n16913_));
  AOI21_X1   g14477(.A1(new_n16053_), .A2(new_n7925_), .B(new_n16913_), .ZN(new_n16914_));
  OAI21_X1   g14478(.A1(new_n16914_), .A2(pi0038), .B(new_n16912_), .ZN(new_n16915_));
  OAI21_X1   g14479(.A1(new_n16915_), .A2(new_n16911_), .B(pi0705), .ZN(new_n16916_));
  NAND2_X1   g14480(.A1(new_n16479_), .A2(pi0167), .ZN(new_n16917_));
  OAI21_X1   g14481(.A1(new_n16021_), .A2(pi0167), .B(new_n16917_), .ZN(new_n16918_));
  NOR2_X1    g14482(.A1(new_n13344_), .A2(pi0167), .ZN(new_n16919_));
  OAI21_X1   g14483(.A1(new_n16809_), .A2(new_n16919_), .B(pi0768), .ZN(new_n16920_));
  AOI21_X1   g14484(.A1(new_n16918_), .A2(new_n3265_), .B(new_n16920_), .ZN(new_n16921_));
  NOR2_X1    g14485(.A1(new_n13191_), .A2(new_n16912_), .ZN(new_n16922_));
  AOI21_X1   g14486(.A1(new_n16922_), .A2(new_n7925_), .B(pi0705), .ZN(new_n16923_));
  NOR2_X1    g14487(.A1(new_n16118_), .A2(pi0167), .ZN(new_n16924_));
  NOR2_X1    g14488(.A1(new_n16096_), .A2(new_n7925_), .ZN(new_n16925_));
  OAI21_X1   g14489(.A1(new_n16924_), .A2(new_n16925_), .B(new_n3265_), .ZN(new_n16926_));
  NAND2_X1   g14490(.A1(new_n16073_), .A2(new_n7925_), .ZN(new_n16927_));
  AOI21_X1   g14491(.A1(new_n16927_), .A2(new_n16081_), .B(pi0768), .ZN(new_n16928_));
  NAND2_X1   g14492(.A1(new_n16926_), .A2(new_n16928_), .ZN(new_n16929_));
  AOI21_X1   g14493(.A1(new_n16929_), .A2(new_n16923_), .B(new_n8265_), .ZN(new_n16930_));
  OAI21_X1   g14494(.A1(new_n16916_), .A2(new_n16921_), .B(new_n16930_), .ZN(new_n16931_));
  AOI22_X1   g14495(.A1(new_n16931_), .A2(new_n16910_), .B1(pi0832), .B2(new_n16909_), .ZN(po0324));
  OAI21_X1   g14496(.A1(new_n3042_), .A2(new_n4571_), .B(pi0832), .ZN(new_n16933_));
  AOI21_X1   g14497(.A1(pi0763), .A2(pi0947), .B(new_n3043_), .ZN(new_n16934_));
  INV_X1     g14498(.I(new_n16934_), .ZN(new_n16935_));
  AOI21_X1   g14499(.A1(pi0699), .A2(new_n15936_), .B(new_n16935_), .ZN(new_n16936_));
  OAI21_X1   g14500(.A1(new_n2582_), .A2(new_n4571_), .B(new_n12738_), .ZN(new_n16937_));
  NAND2_X1   g14501(.A1(new_n5336_), .A2(new_n16934_), .ZN(new_n16938_));
  NAND2_X1   g14502(.A1(new_n16073_), .A2(pi0168), .ZN(new_n16939_));
  NAND3_X1   g14503(.A1(new_n16939_), .A2(pi0038), .A3(new_n16938_), .ZN(new_n16940_));
  NOR2_X1    g14504(.A1(new_n13336_), .A2(pi0763), .ZN(new_n16941_));
  OAI22_X1   g14505(.A1(new_n16941_), .A2(new_n16083_), .B1(pi0168), .B2(new_n16102_), .ZN(new_n16942_));
  NOR2_X1    g14506(.A1(pi0168), .A2(pi0763), .ZN(new_n16943_));
  AOI21_X1   g14507(.A1(new_n14065_), .A2(new_n16943_), .B(new_n2627_), .ZN(new_n16944_));
  INV_X1     g14508(.I(pi0763), .ZN(new_n16945_));
  NAND2_X1   g14509(.A1(new_n16253_), .A2(pi0168), .ZN(new_n16946_));
  AOI21_X1   g14510(.A1(new_n16107_), .A2(new_n16946_), .B(new_n2628_), .ZN(new_n16947_));
  NOR2_X1    g14511(.A1(new_n16248_), .A2(new_n4571_), .ZN(new_n16948_));
  OAI21_X1   g14512(.A1(new_n16002_), .A2(new_n16948_), .B(new_n3304_), .ZN(new_n16949_));
  NAND2_X1   g14513(.A1(new_n13088_), .A2(new_n4571_), .ZN(new_n16950_));
  NAND2_X1   g14514(.A1(new_n16089_), .A2(new_n16950_), .ZN(new_n16951_));
  NAND3_X1   g14515(.A1(new_n16110_), .A2(new_n16949_), .A3(new_n16951_), .ZN(new_n16952_));
  AOI21_X1   g14516(.A1(new_n16952_), .A2(new_n16947_), .B(new_n16945_), .ZN(new_n16953_));
  NAND2_X1   g14517(.A1(new_n16015_), .A2(new_n4571_), .ZN(new_n16954_));
  NAND2_X1   g14518(.A1(new_n16086_), .A2(new_n16954_), .ZN(new_n16955_));
  NAND2_X1   g14519(.A1(new_n16955_), .A2(new_n16953_), .ZN(new_n16956_));
  AOI21_X1   g14520(.A1(new_n16956_), .A2(new_n16944_), .B(pi0038), .ZN(new_n16957_));
  AOI21_X1   g14521(.A1(new_n16957_), .A2(new_n16942_), .B(pi0699), .ZN(new_n16958_));
  AOI21_X1   g14522(.A1(new_n16958_), .A2(new_n16940_), .B(new_n16148_), .ZN(new_n16959_));
  AOI21_X1   g14523(.A1(new_n16945_), .A2(pi0947), .B(new_n16186_), .ZN(new_n16960_));
  OAI21_X1   g14524(.A1(new_n13344_), .A2(pi0168), .B(pi0038), .ZN(new_n16961_));
  AOI21_X1   g14525(.A1(new_n16960_), .A2(new_n2627_), .B(new_n16961_), .ZN(new_n16962_));
  NAND2_X1   g14526(.A1(new_n16954_), .A2(new_n16025_), .ZN(new_n16963_));
  NAND2_X1   g14527(.A1(new_n16105_), .A2(new_n16946_), .ZN(new_n16964_));
  NAND2_X1   g14528(.A1(new_n16964_), .A2(new_n13176_), .ZN(new_n16965_));
  NAND2_X1   g14529(.A1(new_n16965_), .A2(new_n16403_), .ZN(new_n16966_));
  AOI21_X1   g14530(.A1(new_n16270_), .A2(new_n16950_), .B(new_n16005_), .ZN(new_n16967_));
  AOI21_X1   g14531(.A1(new_n16967_), .A2(new_n16949_), .B(pi0215), .ZN(new_n16968_));
  OAI21_X1   g14532(.A1(new_n16968_), .A2(new_n16966_), .B(pi0299), .ZN(new_n16969_));
  NAND3_X1   g14533(.A1(new_n16969_), .A2(new_n16945_), .A3(new_n16963_), .ZN(new_n16970_));
  NOR2_X1    g14534(.A1(new_n16951_), .A2(new_n16411_), .ZN(new_n16971_));
  NOR2_X1    g14535(.A1(new_n16971_), .A2(pi0215), .ZN(new_n16972_));
  NAND2_X1   g14536(.A1(new_n16949_), .A2(new_n16972_), .ZN(new_n16973_));
  AOI21_X1   g14537(.A1(new_n16973_), .A2(new_n16964_), .B(new_n2628_), .ZN(new_n16974_));
  AOI21_X1   g14538(.A1(pi0168), .A2(new_n16055_), .B(new_n16268_), .ZN(new_n16975_));
  OAI21_X1   g14539(.A1(new_n16975_), .A2(new_n16974_), .B(pi0763), .ZN(new_n16976_));
  NAND3_X1   g14540(.A1(new_n16976_), .A2(pi0039), .A3(new_n16970_), .ZN(new_n16977_));
  OR2_X2     g14541(.A1(new_n16942_), .A2(new_n16023_), .Z(new_n16978_));
  AOI21_X1   g14542(.A1(new_n16977_), .A2(new_n16978_), .B(pi0038), .ZN(new_n16979_));
  OAI21_X1   g14543(.A1(new_n16979_), .A2(new_n16962_), .B(pi0699), .ZN(new_n16980_));
  OAI21_X1   g14544(.A1(new_n16147_), .A2(pi0168), .B(new_n2582_), .ZN(new_n16981_));
  AOI21_X1   g14545(.A1(new_n16980_), .A2(new_n16959_), .B(new_n16981_), .ZN(new_n16982_));
  OAI22_X1   g14546(.A1(new_n16982_), .A2(new_n16937_), .B1(new_n16933_), .B2(new_n16936_), .ZN(po0325));
  OAI21_X1   g14547(.A1(new_n3042_), .A2(new_n4414_), .B(pi0832), .ZN(new_n16984_));
  AOI21_X1   g14548(.A1(pi0746), .A2(pi0947), .B(new_n3043_), .ZN(new_n16985_));
  INV_X1     g14549(.I(new_n16985_), .ZN(new_n16986_));
  AOI21_X1   g14550(.A1(pi0729), .A2(new_n15936_), .B(new_n16986_), .ZN(new_n16987_));
  OAI21_X1   g14551(.A1(new_n2582_), .A2(new_n4414_), .B(new_n12738_), .ZN(new_n16988_));
  NAND2_X1   g14552(.A1(new_n5336_), .A2(new_n16985_), .ZN(new_n16989_));
  NAND2_X1   g14553(.A1(new_n16073_), .A2(pi0169), .ZN(new_n16990_));
  NAND3_X1   g14554(.A1(new_n16990_), .A2(pi0038), .A3(new_n16989_), .ZN(new_n16991_));
  NOR2_X1    g14555(.A1(new_n13336_), .A2(pi0746), .ZN(new_n16992_));
  OAI22_X1   g14556(.A1(new_n16992_), .A2(new_n16083_), .B1(pi0169), .B2(new_n16102_), .ZN(new_n16993_));
  NOR2_X1    g14557(.A1(pi0169), .A2(pi0746), .ZN(new_n16994_));
  AOI21_X1   g14558(.A1(new_n14065_), .A2(new_n16994_), .B(new_n2627_), .ZN(new_n16995_));
  INV_X1     g14559(.I(pi0746), .ZN(new_n16996_));
  NAND2_X1   g14560(.A1(new_n16253_), .A2(pi0169), .ZN(new_n16997_));
  AOI21_X1   g14561(.A1(new_n16107_), .A2(new_n16997_), .B(new_n2628_), .ZN(new_n16998_));
  NOR2_X1    g14562(.A1(new_n16248_), .A2(new_n4414_), .ZN(new_n16999_));
  OAI21_X1   g14563(.A1(new_n16002_), .A2(new_n16999_), .B(new_n3304_), .ZN(new_n17000_));
  NAND2_X1   g14564(.A1(new_n13088_), .A2(new_n4414_), .ZN(new_n17001_));
  NAND2_X1   g14565(.A1(new_n16089_), .A2(new_n17001_), .ZN(new_n17002_));
  NAND3_X1   g14566(.A1(new_n16110_), .A2(new_n17000_), .A3(new_n17002_), .ZN(new_n17003_));
  AOI21_X1   g14567(.A1(new_n17003_), .A2(new_n16998_), .B(new_n16996_), .ZN(new_n17004_));
  NAND2_X1   g14568(.A1(new_n16015_), .A2(new_n4414_), .ZN(new_n17005_));
  NAND2_X1   g14569(.A1(new_n16086_), .A2(new_n17005_), .ZN(new_n17006_));
  NAND2_X1   g14570(.A1(new_n17006_), .A2(new_n17004_), .ZN(new_n17007_));
  AOI21_X1   g14571(.A1(new_n17007_), .A2(new_n16995_), .B(pi0038), .ZN(new_n17008_));
  AOI21_X1   g14572(.A1(new_n17008_), .A2(new_n16993_), .B(pi0729), .ZN(new_n17009_));
  AOI21_X1   g14573(.A1(new_n17009_), .A2(new_n16991_), .B(new_n16148_), .ZN(new_n17010_));
  AOI21_X1   g14574(.A1(new_n16996_), .A2(pi0947), .B(new_n16186_), .ZN(new_n17011_));
  OAI21_X1   g14575(.A1(new_n13344_), .A2(pi0169), .B(pi0038), .ZN(new_n17012_));
  AOI21_X1   g14576(.A1(new_n17011_), .A2(new_n2627_), .B(new_n17012_), .ZN(new_n17013_));
  NAND2_X1   g14577(.A1(new_n17005_), .A2(new_n16025_), .ZN(new_n17014_));
  NAND2_X1   g14578(.A1(new_n16105_), .A2(new_n16997_), .ZN(new_n17015_));
  NAND2_X1   g14579(.A1(new_n17015_), .A2(new_n13176_), .ZN(new_n17016_));
  NAND2_X1   g14580(.A1(new_n17016_), .A2(new_n16403_), .ZN(new_n17017_));
  AOI21_X1   g14581(.A1(new_n16270_), .A2(new_n17001_), .B(new_n16005_), .ZN(new_n17018_));
  AOI21_X1   g14582(.A1(new_n17018_), .A2(new_n17000_), .B(pi0215), .ZN(new_n17019_));
  OAI21_X1   g14583(.A1(new_n17019_), .A2(new_n17017_), .B(pi0299), .ZN(new_n17020_));
  NAND3_X1   g14584(.A1(new_n17020_), .A2(new_n16996_), .A3(new_n17014_), .ZN(new_n17021_));
  NOR2_X1    g14585(.A1(new_n17002_), .A2(new_n16411_), .ZN(new_n17022_));
  NOR2_X1    g14586(.A1(new_n17022_), .A2(pi0215), .ZN(new_n17023_));
  NAND2_X1   g14587(.A1(new_n17000_), .A2(new_n17023_), .ZN(new_n17024_));
  AOI21_X1   g14588(.A1(new_n17024_), .A2(new_n17015_), .B(new_n2628_), .ZN(new_n17025_));
  AOI21_X1   g14589(.A1(pi0169), .A2(new_n16055_), .B(new_n16268_), .ZN(new_n17026_));
  OAI21_X1   g14590(.A1(new_n17026_), .A2(new_n17025_), .B(pi0746), .ZN(new_n17027_));
  NAND3_X1   g14591(.A1(new_n17027_), .A2(pi0039), .A3(new_n17021_), .ZN(new_n17028_));
  OR2_X2     g14592(.A1(new_n16993_), .A2(new_n16023_), .Z(new_n17029_));
  AOI21_X1   g14593(.A1(new_n17028_), .A2(new_n17029_), .B(pi0038), .ZN(new_n17030_));
  OAI21_X1   g14594(.A1(new_n17030_), .A2(new_n17013_), .B(pi0729), .ZN(new_n17031_));
  OAI21_X1   g14595(.A1(new_n16147_), .A2(pi0169), .B(new_n2582_), .ZN(new_n17032_));
  AOI21_X1   g14596(.A1(new_n17031_), .A2(new_n17010_), .B(new_n17032_), .ZN(new_n17033_));
  OAI22_X1   g14597(.A1(new_n17033_), .A2(new_n16988_), .B1(new_n16984_), .B2(new_n16987_), .ZN(po0326));
  OAI21_X1   g14598(.A1(new_n3042_), .A2(new_n4089_), .B(pi0832), .ZN(new_n17035_));
  INV_X1     g14599(.I(pi0748), .ZN(new_n17036_));
  OAI21_X1   g14600(.A1(new_n17036_), .A2(new_n5692_), .B(new_n3042_), .ZN(new_n17037_));
  AOI21_X1   g14601(.A1(pi0730), .A2(new_n15936_), .B(new_n17037_), .ZN(new_n17038_));
  OAI21_X1   g14602(.A1(new_n2582_), .A2(new_n4089_), .B(new_n12738_), .ZN(new_n17039_));
  NOR2_X1    g14603(.A1(new_n13191_), .A2(pi0748), .ZN(new_n17040_));
  AOI21_X1   g14604(.A1(new_n17040_), .A2(new_n4089_), .B(pi0730), .ZN(new_n17041_));
  OAI21_X1   g14605(.A1(new_n4089_), .A2(new_n15975_), .B(new_n16107_), .ZN(new_n17042_));
  NAND2_X1   g14606(.A1(new_n17042_), .A2(pi0299), .ZN(new_n17043_));
  NAND2_X1   g14607(.A1(new_n13088_), .A2(new_n4089_), .ZN(new_n17044_));
  NAND2_X1   g14608(.A1(new_n16089_), .A2(new_n17044_), .ZN(new_n17045_));
  OAI21_X1   g14609(.A1(new_n13093_), .A2(new_n5420_), .B(pi0170), .ZN(new_n17046_));
  AOI21_X1   g14610(.A1(new_n13127_), .A2(new_n17046_), .B(new_n3303_), .ZN(new_n17047_));
  INV_X1     g14611(.I(new_n17047_), .ZN(new_n17048_));
  AND3_X2    g14612(.A1(new_n16110_), .A2(new_n17045_), .A3(new_n17048_), .Z(new_n17049_));
  NOR2_X1    g14613(.A1(new_n16014_), .A2(pi0170), .ZN(new_n17050_));
  OAI22_X1   g14614(.A1(new_n17043_), .A2(new_n17049_), .B1(new_n16085_), .B2(new_n17050_), .ZN(new_n17051_));
  NOR2_X1    g14615(.A1(new_n16102_), .A2(pi0170), .ZN(new_n17052_));
  INV_X1     g14616(.I(new_n17052_), .ZN(new_n17053_));
  AOI22_X1   g14617(.A1(new_n17051_), .A2(pi0039), .B1(new_n16083_), .B2(new_n17053_), .ZN(new_n17054_));
  NAND2_X1   g14618(.A1(new_n16073_), .A2(new_n4089_), .ZN(new_n17055_));
  AOI21_X1   g14619(.A1(new_n17055_), .A2(new_n16081_), .B(new_n17036_), .ZN(new_n17056_));
  OAI21_X1   g14620(.A1(new_n17054_), .A2(pi0038), .B(new_n17056_), .ZN(new_n17057_));
  AOI21_X1   g14621(.A1(new_n17057_), .A2(new_n17041_), .B(new_n16148_), .ZN(new_n17058_));
  NAND2_X1   g14622(.A1(new_n13397_), .A2(new_n4089_), .ZN(new_n17059_));
  AOI21_X1   g14623(.A1(new_n16072_), .A2(new_n17059_), .B(new_n17036_), .ZN(new_n17060_));
  NOR2_X1    g14624(.A1(new_n17052_), .A2(new_n16063_), .ZN(new_n17061_));
  AOI21_X1   g14625(.A1(pi0170), .A2(new_n16253_), .B(new_n16106_), .ZN(new_n17062_));
  OAI21_X1   g14626(.A1(new_n17045_), .A2(new_n16411_), .B(new_n2436_), .ZN(new_n17063_));
  NOR2_X1    g14627(.A1(new_n17047_), .A2(new_n17063_), .ZN(new_n17064_));
  OAI21_X1   g14628(.A1(new_n17062_), .A2(new_n17064_), .B(pi0299), .ZN(new_n17065_));
  NAND2_X1   g14629(.A1(new_n16055_), .A2(pi0170), .ZN(new_n17066_));
  AOI21_X1   g14630(.A1(new_n17066_), .A2(new_n16049_), .B(new_n2627_), .ZN(new_n17067_));
  AOI22_X1   g14631(.A1(new_n17067_), .A2(new_n17065_), .B1(new_n2627_), .B2(new_n17061_), .ZN(new_n17068_));
  OAI21_X1   g14632(.A1(new_n17068_), .A2(pi0038), .B(new_n17060_), .ZN(new_n17069_));
  OAI21_X1   g14633(.A1(new_n17062_), .A2(new_n16056_), .B(new_n16403_), .ZN(new_n17070_));
  AOI21_X1   g14634(.A1(new_n16270_), .A2(new_n17044_), .B(new_n16005_), .ZN(new_n17071_));
  AOI21_X1   g14635(.A1(new_n17071_), .A2(new_n17048_), .B(pi0215), .ZN(new_n17072_));
  OAI21_X1   g14636(.A1(new_n17072_), .A2(new_n17070_), .B(pi0299), .ZN(new_n17073_));
  OAI21_X1   g14637(.A1(pi0170), .A2(new_n16014_), .B(new_n16025_), .ZN(new_n17074_));
  AOI21_X1   g14638(.A1(new_n17073_), .A2(new_n17074_), .B(new_n2627_), .ZN(new_n17075_));
  NOR2_X1    g14639(.A1(new_n16433_), .A2(new_n17052_), .ZN(new_n17076_));
  OAI21_X1   g14640(.A1(new_n17075_), .A2(new_n17076_), .B(new_n3265_), .ZN(new_n17077_));
  AOI21_X1   g14641(.A1(new_n17059_), .A2(new_n15999_), .B(pi0748), .ZN(new_n17078_));
  NAND2_X1   g14642(.A1(new_n17077_), .A2(new_n17078_), .ZN(new_n17079_));
  NAND3_X1   g14643(.A1(new_n17069_), .A2(new_n17079_), .A3(pi0730), .ZN(new_n17080_));
  OAI21_X1   g14644(.A1(new_n16147_), .A2(pi0170), .B(new_n2582_), .ZN(new_n17081_));
  AOI21_X1   g14645(.A1(new_n17080_), .A2(new_n17058_), .B(new_n17081_), .ZN(new_n17082_));
  OAI22_X1   g14646(.A1(new_n17082_), .A2(new_n17039_), .B1(new_n17035_), .B2(new_n17038_), .ZN(po0327));
  OAI21_X1   g14647(.A1(new_n3042_), .A2(new_n3932_), .B(pi0832), .ZN(new_n17084_));
  AOI21_X1   g14648(.A1(pi0764), .A2(pi0947), .B(new_n3043_), .ZN(new_n17085_));
  INV_X1     g14649(.I(new_n17085_), .ZN(new_n17086_));
  AOI21_X1   g14650(.A1(pi0691), .A2(new_n15936_), .B(new_n17086_), .ZN(new_n17087_));
  OAI21_X1   g14651(.A1(new_n2582_), .A2(new_n3932_), .B(new_n12738_), .ZN(new_n17088_));
  NAND2_X1   g14652(.A1(new_n5336_), .A2(new_n17085_), .ZN(new_n17089_));
  NAND2_X1   g14653(.A1(new_n16073_), .A2(pi0171), .ZN(new_n17090_));
  NAND3_X1   g14654(.A1(new_n17090_), .A2(pi0038), .A3(new_n17089_), .ZN(new_n17091_));
  NOR2_X1    g14655(.A1(new_n13336_), .A2(pi0764), .ZN(new_n17092_));
  OAI22_X1   g14656(.A1(new_n17092_), .A2(new_n16083_), .B1(pi0171), .B2(new_n16102_), .ZN(new_n17093_));
  NOR2_X1    g14657(.A1(pi0171), .A2(pi0764), .ZN(new_n17094_));
  AOI21_X1   g14658(.A1(new_n14065_), .A2(new_n17094_), .B(new_n2627_), .ZN(new_n17095_));
  INV_X1     g14659(.I(pi0764), .ZN(new_n17096_));
  NAND2_X1   g14660(.A1(new_n16253_), .A2(pi0171), .ZN(new_n17097_));
  AOI21_X1   g14661(.A1(new_n16107_), .A2(new_n17097_), .B(new_n2628_), .ZN(new_n17098_));
  NOR2_X1    g14662(.A1(new_n16248_), .A2(new_n3932_), .ZN(new_n17099_));
  OAI21_X1   g14663(.A1(new_n16002_), .A2(new_n17099_), .B(new_n3304_), .ZN(new_n17100_));
  NAND2_X1   g14664(.A1(new_n13088_), .A2(new_n3932_), .ZN(new_n17101_));
  NAND2_X1   g14665(.A1(new_n16089_), .A2(new_n17101_), .ZN(new_n17102_));
  NAND3_X1   g14666(.A1(new_n16110_), .A2(new_n17100_), .A3(new_n17102_), .ZN(new_n17103_));
  AOI21_X1   g14667(.A1(new_n17103_), .A2(new_n17098_), .B(new_n17096_), .ZN(new_n17104_));
  NAND2_X1   g14668(.A1(new_n16015_), .A2(new_n3932_), .ZN(new_n17105_));
  NAND2_X1   g14669(.A1(new_n16086_), .A2(new_n17105_), .ZN(new_n17106_));
  NAND2_X1   g14670(.A1(new_n17106_), .A2(new_n17104_), .ZN(new_n17107_));
  AOI21_X1   g14671(.A1(new_n17107_), .A2(new_n17095_), .B(pi0038), .ZN(new_n17108_));
  AOI21_X1   g14672(.A1(new_n17108_), .A2(new_n17093_), .B(pi0691), .ZN(new_n17109_));
  AOI21_X1   g14673(.A1(new_n17109_), .A2(new_n17091_), .B(new_n16148_), .ZN(new_n17110_));
  AOI21_X1   g14674(.A1(new_n17096_), .A2(pi0947), .B(new_n16186_), .ZN(new_n17111_));
  OAI21_X1   g14675(.A1(new_n13344_), .A2(pi0171), .B(pi0038), .ZN(new_n17112_));
  AOI21_X1   g14676(.A1(new_n17111_), .A2(new_n2627_), .B(new_n17112_), .ZN(new_n17113_));
  NAND2_X1   g14677(.A1(new_n17105_), .A2(new_n16025_), .ZN(new_n17114_));
  NAND2_X1   g14678(.A1(new_n16105_), .A2(new_n17097_), .ZN(new_n17115_));
  NAND2_X1   g14679(.A1(new_n17115_), .A2(new_n13176_), .ZN(new_n17116_));
  NAND2_X1   g14680(.A1(new_n17116_), .A2(new_n16403_), .ZN(new_n17117_));
  AOI21_X1   g14681(.A1(new_n16270_), .A2(new_n17101_), .B(new_n16005_), .ZN(new_n17118_));
  AOI21_X1   g14682(.A1(new_n17118_), .A2(new_n17100_), .B(pi0215), .ZN(new_n17119_));
  OAI21_X1   g14683(.A1(new_n17119_), .A2(new_n17117_), .B(pi0299), .ZN(new_n17120_));
  NAND3_X1   g14684(.A1(new_n17120_), .A2(new_n17096_), .A3(new_n17114_), .ZN(new_n17121_));
  NOR2_X1    g14685(.A1(new_n17102_), .A2(new_n16411_), .ZN(new_n17122_));
  NOR2_X1    g14686(.A1(new_n17122_), .A2(pi0215), .ZN(new_n17123_));
  NAND2_X1   g14687(.A1(new_n17100_), .A2(new_n17123_), .ZN(new_n17124_));
  AOI21_X1   g14688(.A1(new_n17124_), .A2(new_n17115_), .B(new_n2628_), .ZN(new_n17125_));
  AOI21_X1   g14689(.A1(pi0171), .A2(new_n16055_), .B(new_n16268_), .ZN(new_n17126_));
  OAI21_X1   g14690(.A1(new_n17126_), .A2(new_n17125_), .B(pi0764), .ZN(new_n17127_));
  NAND3_X1   g14691(.A1(new_n17127_), .A2(pi0039), .A3(new_n17121_), .ZN(new_n17128_));
  OR2_X2     g14692(.A1(new_n17093_), .A2(new_n16023_), .Z(new_n17129_));
  AOI21_X1   g14693(.A1(new_n17128_), .A2(new_n17129_), .B(pi0038), .ZN(new_n17130_));
  OAI21_X1   g14694(.A1(new_n17130_), .A2(new_n17113_), .B(pi0691), .ZN(new_n17131_));
  OAI21_X1   g14695(.A1(new_n16147_), .A2(pi0171), .B(new_n2582_), .ZN(new_n17132_));
  AOI21_X1   g14696(.A1(new_n17131_), .A2(new_n17110_), .B(new_n17132_), .ZN(new_n17133_));
  OAI22_X1   g14697(.A1(new_n17133_), .A2(new_n17088_), .B1(new_n17084_), .B2(new_n17087_), .ZN(po0328));
  INV_X1     g14698(.I(pi0739), .ZN(new_n17135_));
  NOR2_X1    g14699(.A1(new_n17135_), .A2(new_n5692_), .ZN(new_n17136_));
  INV_X1     g14700(.I(pi0690), .ZN(new_n17137_));
  NOR2_X1    g14701(.A1(new_n15994_), .A2(new_n17137_), .ZN(new_n17138_));
  NOR3_X1    g14702(.A1(new_n17138_), .A2(new_n3043_), .A3(new_n17136_), .ZN(new_n17139_));
  OAI21_X1   g14703(.A1(new_n3042_), .A2(new_n3778_), .B(pi0832), .ZN(new_n17140_));
  OAI21_X1   g14704(.A1(new_n2582_), .A2(new_n3778_), .B(new_n12738_), .ZN(new_n17141_));
  AOI21_X1   g14705(.A1(new_n16073_), .A2(pi0172), .B(new_n3265_), .ZN(new_n17142_));
  OAI21_X1   g14706(.A1(new_n13397_), .A2(new_n17136_), .B(new_n17142_), .ZN(new_n17143_));
  NOR2_X1    g14707(.A1(new_n13060_), .A2(new_n17136_), .ZN(new_n17144_));
  NOR2_X1    g14708(.A1(new_n16102_), .A2(new_n3778_), .ZN(new_n17145_));
  OAI21_X1   g14709(.A1(new_n17145_), .A2(new_n17144_), .B(new_n2627_), .ZN(new_n17146_));
  NOR2_X1    g14710(.A1(pi0172), .A2(pi0739), .ZN(new_n17147_));
  AOI21_X1   g14711(.A1(new_n14065_), .A2(new_n17147_), .B(new_n2627_), .ZN(new_n17148_));
  NAND2_X1   g14712(.A1(new_n16253_), .A2(pi0172), .ZN(new_n17149_));
  AOI21_X1   g14713(.A1(new_n16107_), .A2(new_n17149_), .B(new_n2628_), .ZN(new_n17150_));
  NOR2_X1    g14714(.A1(new_n16248_), .A2(new_n3778_), .ZN(new_n17151_));
  OAI21_X1   g14715(.A1(new_n16002_), .A2(new_n17151_), .B(new_n3304_), .ZN(new_n17152_));
  NAND2_X1   g14716(.A1(new_n13088_), .A2(new_n3778_), .ZN(new_n17153_));
  NAND2_X1   g14717(.A1(new_n16089_), .A2(new_n17153_), .ZN(new_n17154_));
  NAND3_X1   g14718(.A1(new_n16110_), .A2(new_n17152_), .A3(new_n17154_), .ZN(new_n17155_));
  AOI21_X1   g14719(.A1(new_n17155_), .A2(new_n17150_), .B(new_n17135_), .ZN(new_n17156_));
  NAND2_X1   g14720(.A1(new_n16015_), .A2(new_n3778_), .ZN(new_n17157_));
  NAND2_X1   g14721(.A1(new_n16086_), .A2(new_n17157_), .ZN(new_n17158_));
  NAND2_X1   g14722(.A1(new_n17158_), .A2(new_n17156_), .ZN(new_n17159_));
  AOI21_X1   g14723(.A1(new_n17159_), .A2(new_n17148_), .B(pi0038), .ZN(new_n17160_));
  AOI21_X1   g14724(.A1(new_n17160_), .A2(new_n17146_), .B(pi0690), .ZN(new_n17161_));
  AOI21_X1   g14725(.A1(new_n17161_), .A2(new_n17143_), .B(new_n16148_), .ZN(new_n17162_));
  AOI21_X1   g14726(.A1(new_n17135_), .A2(pi0947), .B(new_n16186_), .ZN(new_n17163_));
  OAI21_X1   g14727(.A1(new_n13344_), .A2(pi0172), .B(pi0038), .ZN(new_n17164_));
  AOI21_X1   g14728(.A1(new_n17163_), .A2(new_n2627_), .B(new_n17164_), .ZN(new_n17165_));
  NAND2_X1   g14729(.A1(new_n17157_), .A2(new_n16025_), .ZN(new_n17166_));
  NAND2_X1   g14730(.A1(new_n16105_), .A2(new_n17149_), .ZN(new_n17167_));
  NAND2_X1   g14731(.A1(new_n17167_), .A2(new_n13176_), .ZN(new_n17168_));
  NAND2_X1   g14732(.A1(new_n17168_), .A2(new_n16403_), .ZN(new_n17169_));
  AOI21_X1   g14733(.A1(new_n16270_), .A2(new_n17153_), .B(new_n16005_), .ZN(new_n17170_));
  AOI21_X1   g14734(.A1(new_n17170_), .A2(new_n17152_), .B(pi0215), .ZN(new_n17171_));
  OAI21_X1   g14735(.A1(new_n17171_), .A2(new_n17169_), .B(pi0299), .ZN(new_n17172_));
  NAND3_X1   g14736(.A1(new_n17172_), .A2(new_n17135_), .A3(new_n17166_), .ZN(new_n17173_));
  NOR2_X1    g14737(.A1(new_n17154_), .A2(new_n16411_), .ZN(new_n17174_));
  NOR2_X1    g14738(.A1(new_n17174_), .A2(pi0215), .ZN(new_n17175_));
  NAND2_X1   g14739(.A1(new_n17152_), .A2(new_n17175_), .ZN(new_n17176_));
  AOI21_X1   g14740(.A1(new_n17176_), .A2(new_n17167_), .B(new_n2628_), .ZN(new_n17177_));
  AOI21_X1   g14741(.A1(pi0172), .A2(new_n16055_), .B(new_n16268_), .ZN(new_n17178_));
  OAI21_X1   g14742(.A1(new_n17178_), .A2(new_n17177_), .B(pi0739), .ZN(new_n17179_));
  NAND3_X1   g14743(.A1(new_n17179_), .A2(pi0039), .A3(new_n17173_), .ZN(new_n17180_));
  OR2_X2     g14744(.A1(new_n17146_), .A2(new_n16023_), .Z(new_n17181_));
  AOI21_X1   g14745(.A1(new_n17180_), .A2(new_n17181_), .B(pi0038), .ZN(new_n17182_));
  OAI21_X1   g14746(.A1(new_n17182_), .A2(new_n17165_), .B(pi0690), .ZN(new_n17183_));
  OAI21_X1   g14747(.A1(new_n16147_), .A2(pi0172), .B(new_n2582_), .ZN(new_n17184_));
  AOI21_X1   g14748(.A1(new_n17183_), .A2(new_n17162_), .B(new_n17184_), .ZN(new_n17185_));
  OAI22_X1   g14749(.A1(new_n17185_), .A2(new_n17141_), .B1(new_n17139_), .B2(new_n17140_), .ZN(po0329));
  INV_X1     g14750(.I(new_n12871_), .ZN(new_n17187_));
  NOR2_X1    g14751(.A1(new_n3042_), .A2(pi0173), .ZN(new_n17188_));
  AOI21_X1   g14752(.A1(new_n12826_), .A2(new_n16263_), .B(new_n17188_), .ZN(new_n17189_));
  NOR2_X1    g14753(.A1(new_n17188_), .A2(pi1153), .ZN(new_n17190_));
  NOR2_X1    g14754(.A1(new_n12834_), .A2(pi0723), .ZN(new_n17191_));
  INV_X1     g14755(.I(new_n17191_), .ZN(new_n17192_));
  NAND2_X1   g14756(.A1(new_n17192_), .A2(new_n17190_), .ZN(new_n17193_));
  NOR2_X1    g14757(.A1(new_n17191_), .A2(new_n17189_), .ZN(new_n17194_));
  NOR2_X1    g14758(.A1(new_n17194_), .A2(new_n12841_), .ZN(new_n17195_));
  INV_X1     g14759(.I(new_n17195_), .ZN(new_n17196_));
  NAND3_X1   g14760(.A1(new_n17196_), .A2(pi0778), .A3(new_n17193_), .ZN(new_n17197_));
  OAI21_X1   g14761(.A1(pi0778), .A2(new_n17189_), .B(new_n17197_), .ZN(new_n17198_));
  NAND2_X1   g14762(.A1(new_n17198_), .A2(new_n17187_), .ZN(new_n17199_));
  NOR2_X1    g14763(.A1(new_n17199_), .A2(new_n12889_), .ZN(new_n17200_));
  INV_X1     g14764(.I(new_n17200_), .ZN(new_n17201_));
  NOR2_X1    g14765(.A1(new_n17201_), .A2(new_n12924_), .ZN(new_n17202_));
  NAND2_X1   g14766(.A1(new_n17202_), .A2(new_n12954_), .ZN(new_n17203_));
  NAND2_X1   g14767(.A1(new_n17203_), .A2(new_n12741_), .ZN(new_n17204_));
  INV_X1     g14768(.I(new_n17188_), .ZN(new_n17205_));
  NAND2_X1   g14769(.A1(new_n17205_), .A2(pi0647), .ZN(new_n17206_));
  AOI21_X1   g14770(.A1(new_n17204_), .A2(new_n17206_), .B(pi1157), .ZN(new_n17207_));
  INV_X1     g14771(.I(new_n17207_), .ZN(new_n17208_));
  NAND2_X1   g14772(.A1(new_n17188_), .A2(new_n12741_), .ZN(new_n17209_));
  OAI21_X1   g14773(.A1(new_n17203_), .A2(new_n12741_), .B(new_n17209_), .ZN(new_n17210_));
  OAI22_X1   g14774(.A1(new_n17208_), .A2(new_n12981_), .B1(new_n15576_), .B2(new_n17210_), .ZN(new_n17211_));
  INV_X1     g14775(.I(new_n15608_), .ZN(new_n17212_));
  NOR2_X1    g14776(.A1(new_n13340_), .A2(pi0745), .ZN(new_n17213_));
  NOR2_X1    g14777(.A1(new_n17213_), .A2(new_n17188_), .ZN(new_n17214_));
  NOR3_X1    g14778(.A1(new_n17214_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n17215_));
  INV_X1     g14779(.I(new_n17213_), .ZN(new_n17216_));
  NOR2_X1    g14780(.A1(new_n17216_), .A2(new_n13354_), .ZN(new_n17217_));
  NOR3_X1    g14781(.A1(new_n17217_), .A2(new_n12762_), .A3(new_n17214_), .ZN(new_n17218_));
  NOR2_X1    g14782(.A1(new_n17218_), .A2(new_n12770_), .ZN(new_n17219_));
  NOR3_X1    g14783(.A1(new_n17217_), .A2(pi1155), .A3(new_n17188_), .ZN(new_n17220_));
  NOR3_X1    g14784(.A1(new_n17219_), .A2(new_n12764_), .A3(new_n17220_), .ZN(new_n17221_));
  NOR2_X1    g14785(.A1(new_n17221_), .A2(new_n17215_), .ZN(new_n17222_));
  INV_X1     g14786(.I(new_n17222_), .ZN(new_n17223_));
  AOI21_X1   g14787(.A1(new_n17223_), .A2(new_n12783_), .B(pi1154), .ZN(new_n17224_));
  INV_X1     g14788(.I(new_n17224_), .ZN(new_n17225_));
  AOI21_X1   g14789(.A1(new_n17223_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n17226_));
  NOR2_X1    g14790(.A1(new_n17226_), .A2(new_n12779_), .ZN(new_n17227_));
  AOI22_X1   g14791(.A1(new_n17227_), .A2(new_n17225_), .B1(new_n12779_), .B2(new_n17223_), .ZN(new_n17228_));
  NOR2_X1    g14792(.A1(new_n3043_), .A2(new_n12793_), .ZN(new_n17229_));
  NOR2_X1    g14793(.A1(new_n17228_), .A2(new_n17229_), .ZN(new_n17230_));
  NOR2_X1    g14794(.A1(new_n17230_), .A2(pi1159), .ZN(new_n17231_));
  NOR2_X1    g14795(.A1(new_n3043_), .A2(pi0619), .ZN(new_n17232_));
  OAI21_X1   g14796(.A1(new_n17228_), .A2(new_n17232_), .B(pi1159), .ZN(new_n17233_));
  NAND2_X1   g14797(.A1(new_n17233_), .A2(pi0789), .ZN(new_n17234_));
  OAI22_X1   g14798(.A1(new_n17234_), .A2(new_n17231_), .B1(pi0789), .B2(new_n17228_), .ZN(new_n17235_));
  AOI22_X1   g14799(.A1(new_n17235_), .A2(new_n12804_), .B1(new_n15609_), .B2(new_n17188_), .ZN(new_n17236_));
  NAND2_X1   g14800(.A1(new_n17235_), .A2(new_n12808_), .ZN(new_n17237_));
  OAI21_X1   g14801(.A1(new_n17236_), .A2(new_n12808_), .B(new_n17237_), .ZN(new_n17238_));
  NOR2_X1    g14802(.A1(new_n17238_), .A2(new_n12943_), .ZN(new_n17239_));
  AOI21_X1   g14803(.A1(new_n12943_), .A2(new_n17205_), .B(new_n17239_), .ZN(new_n17240_));
  NOR2_X1    g14804(.A1(new_n17240_), .A2(new_n17212_), .ZN(new_n17241_));
  NOR2_X1    g14805(.A1(new_n17241_), .A2(new_n17211_), .ZN(new_n17242_));
  INV_X1     g14806(.I(new_n17220_), .ZN(new_n17243_));
  NOR2_X1    g14807(.A1(new_n17189_), .A2(new_n12754_), .ZN(new_n17244_));
  NOR3_X1    g14808(.A1(new_n17244_), .A2(new_n17188_), .A3(new_n17213_), .ZN(new_n17245_));
  NAND2_X1   g14809(.A1(new_n17245_), .A2(new_n12758_), .ZN(new_n17246_));
  NAND2_X1   g14810(.A1(new_n17244_), .A2(pi0625), .ZN(new_n17247_));
  NAND3_X1   g14811(.A1(new_n17247_), .A2(pi1153), .A3(new_n17214_), .ZN(new_n17248_));
  NAND3_X1   g14812(.A1(new_n17193_), .A2(pi0608), .A3(new_n17248_), .ZN(new_n17249_));
  INV_X1     g14813(.I(new_n17247_), .ZN(new_n17250_));
  OAI21_X1   g14814(.A1(new_n17250_), .A2(new_n17245_), .B(new_n17190_), .ZN(new_n17251_));
  NAND3_X1   g14815(.A1(new_n17196_), .A2(new_n13560_), .A3(new_n17251_), .ZN(new_n17252_));
  NAND3_X1   g14816(.A1(new_n17252_), .A2(pi0778), .A3(new_n17249_), .ZN(new_n17253_));
  AOI21_X1   g14817(.A1(new_n17253_), .A2(new_n17246_), .B(new_n12766_), .ZN(new_n17254_));
  NOR2_X1    g14818(.A1(new_n17198_), .A2(pi0609), .ZN(new_n17255_));
  OAI21_X1   g14819(.A1(new_n17255_), .A2(new_n17254_), .B(pi1155), .ZN(new_n17256_));
  NAND3_X1   g14820(.A1(new_n17256_), .A2(pi0660), .A3(new_n17243_), .ZN(new_n17257_));
  NAND2_X1   g14821(.A1(new_n17253_), .A2(new_n17246_), .ZN(new_n17258_));
  NOR2_X1    g14822(.A1(new_n17198_), .A2(new_n12766_), .ZN(new_n17259_));
  AOI21_X1   g14823(.A1(new_n17258_), .A2(new_n12766_), .B(new_n17259_), .ZN(new_n17260_));
  NOR2_X1    g14824(.A1(new_n17219_), .A2(pi0660), .ZN(new_n17261_));
  OAI21_X1   g14825(.A1(new_n17260_), .A2(pi1155), .B(new_n17261_), .ZN(new_n17262_));
  NAND3_X1   g14826(.A1(new_n17262_), .A2(new_n17257_), .A3(pi0785), .ZN(new_n17263_));
  NAND2_X1   g14827(.A1(new_n17258_), .A2(new_n12764_), .ZN(new_n17264_));
  NAND2_X1   g14828(.A1(new_n17263_), .A2(new_n17264_), .ZN(new_n17265_));
  NAND2_X1   g14829(.A1(new_n17265_), .A2(new_n12781_), .ZN(new_n17266_));
  NAND2_X1   g14830(.A1(new_n17199_), .A2(pi0618), .ZN(new_n17267_));
  AOI21_X1   g14831(.A1(new_n17266_), .A2(new_n17267_), .B(pi1154), .ZN(new_n17268_));
  NOR3_X1    g14832(.A1(new_n17268_), .A2(pi0627), .A3(new_n17226_), .ZN(new_n17269_));
  NAND2_X1   g14833(.A1(new_n17199_), .A2(new_n12781_), .ZN(new_n17270_));
  NAND2_X1   g14834(.A1(new_n17265_), .A2(pi0618), .ZN(new_n17271_));
  AOI21_X1   g14835(.A1(new_n17271_), .A2(new_n17270_), .B(new_n12785_), .ZN(new_n17272_));
  NOR3_X1    g14836(.A1(new_n17272_), .A2(new_n12880_), .A3(new_n17224_), .ZN(new_n17273_));
  OR3_X2     g14837(.A1(new_n17269_), .A2(new_n17273_), .A3(new_n12779_), .Z(new_n17274_));
  NAND2_X1   g14838(.A1(new_n17265_), .A2(new_n12779_), .ZN(new_n17275_));
  NAND2_X1   g14839(.A1(new_n17274_), .A2(new_n17275_), .ZN(new_n17276_));
  AOI21_X1   g14840(.A1(new_n17276_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n17277_));
  NAND2_X1   g14841(.A1(new_n17201_), .A2(new_n12793_), .ZN(new_n17278_));
  NAND2_X1   g14842(.A1(new_n17276_), .A2(pi0619), .ZN(new_n17279_));
  AOI21_X1   g14843(.A1(new_n17279_), .A2(new_n17278_), .B(new_n12791_), .ZN(new_n17280_));
  NOR3_X1    g14844(.A1(new_n17280_), .A2(new_n12895_), .A3(new_n17231_), .ZN(new_n17281_));
  AOI21_X1   g14845(.A1(new_n17274_), .A2(new_n17275_), .B(pi0619), .ZN(new_n17282_));
  NOR2_X1    g14846(.A1(new_n17200_), .A2(new_n12793_), .ZN(new_n17283_));
  OAI21_X1   g14847(.A1(new_n17282_), .A2(new_n17283_), .B(new_n12791_), .ZN(new_n17284_));
  NAND3_X1   g14848(.A1(new_n17284_), .A2(new_n12895_), .A3(new_n17233_), .ZN(new_n17285_));
  NAND2_X1   g14849(.A1(new_n17285_), .A2(pi0789), .ZN(new_n17286_));
  OAI21_X1   g14850(.A1(new_n17286_), .A2(new_n17281_), .B(new_n17277_), .ZN(new_n17287_));
  OAI22_X1   g14851(.A1(new_n17236_), .A2(new_n15689_), .B1(new_n15688_), .B2(new_n17201_), .ZN(new_n17288_));
  NAND2_X1   g14852(.A1(new_n17288_), .A2(pi0788), .ZN(new_n17289_));
  AOI21_X1   g14853(.A1(new_n17287_), .A2(new_n17289_), .B(new_n15340_), .ZN(new_n17290_));
  AOI22_X1   g14854(.A1(new_n17238_), .A2(new_n12949_), .B1(new_n15695_), .B2(new_n17202_), .ZN(new_n17291_));
  NOR2_X1    g14855(.A1(new_n17291_), .A2(pi0629), .ZN(new_n17292_));
  AOI22_X1   g14856(.A1(new_n17238_), .A2(new_n12948_), .B1(new_n15700_), .B2(new_n17202_), .ZN(new_n17293_));
  NOR2_X1    g14857(.A1(new_n17293_), .A2(new_n12919_), .ZN(new_n17294_));
  OAI21_X1   g14858(.A1(new_n17292_), .A2(new_n17294_), .B(pi0792), .ZN(new_n17295_));
  NAND2_X1   g14859(.A1(new_n17295_), .A2(new_n15693_), .ZN(new_n17296_));
  OAI22_X1   g14860(.A1(new_n17290_), .A2(new_n17296_), .B1(new_n12972_), .B2(new_n17242_), .ZN(new_n17297_));
  NAND2_X1   g14861(.A1(new_n17297_), .A2(new_n13000_), .ZN(new_n17298_));
  AND2_X2    g14862(.A1(new_n17297_), .A2(new_n12975_), .Z(new_n17299_));
  NOR2_X1    g14863(.A1(new_n17210_), .A2(new_n12965_), .ZN(new_n17300_));
  NOR3_X1    g14864(.A1(new_n17300_), .A2(new_n17207_), .A3(new_n12972_), .ZN(new_n17301_));
  NOR2_X1    g14865(.A1(new_n17203_), .A2(pi0787), .ZN(new_n17302_));
  NOR3_X1    g14866(.A1(new_n17301_), .A2(new_n12975_), .A3(new_n17302_), .ZN(new_n17303_));
  OAI21_X1   g14867(.A1(new_n17299_), .A2(new_n17303_), .B(new_n12740_), .ZN(new_n17304_));
  NOR2_X1    g14868(.A1(new_n17188_), .A2(new_n12975_), .ZN(new_n17305_));
  NOR2_X1    g14869(.A1(new_n17240_), .A2(new_n12984_), .ZN(new_n17306_));
  AOI21_X1   g14870(.A1(new_n12984_), .A2(new_n17205_), .B(new_n17306_), .ZN(new_n17307_));
  NOR2_X1    g14871(.A1(new_n17307_), .A2(pi0644), .ZN(new_n17308_));
  OAI21_X1   g14872(.A1(new_n17308_), .A2(new_n17305_), .B(pi0715), .ZN(new_n17309_));
  NAND3_X1   g14873(.A1(new_n17304_), .A2(new_n12739_), .A3(new_n17309_), .ZN(new_n17310_));
  NOR3_X1    g14874(.A1(new_n17301_), .A2(pi0644), .A3(new_n17302_), .ZN(new_n17311_));
  AOI21_X1   g14875(.A1(new_n17297_), .A2(pi0644), .B(new_n17311_), .ZN(new_n17312_));
  NAND2_X1   g14876(.A1(new_n17205_), .A2(new_n12975_), .ZN(new_n17313_));
  OAI21_X1   g14877(.A1(new_n17307_), .A2(new_n12975_), .B(new_n17313_), .ZN(new_n17314_));
  AOI21_X1   g14878(.A1(new_n17314_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n17315_));
  OAI21_X1   g14879(.A1(new_n17312_), .A2(new_n12740_), .B(new_n17315_), .ZN(new_n17316_));
  NAND3_X1   g14880(.A1(new_n17310_), .A2(pi0790), .A3(new_n17316_), .ZN(new_n17317_));
  NAND2_X1   g14881(.A1(new_n17317_), .A2(new_n17298_), .ZN(new_n17318_));
  AOI21_X1   g14882(.A1(po1038), .A2(new_n10736_), .B(pi0832), .ZN(new_n17319_));
  NAND2_X1   g14883(.A1(new_n13192_), .A2(new_n10736_), .ZN(new_n17320_));
  NOR2_X1    g14884(.A1(new_n17320_), .A2(new_n12870_), .ZN(new_n17321_));
  INV_X1     g14885(.I(new_n17321_), .ZN(new_n17322_));
  INV_X1     g14886(.I(new_n17320_), .ZN(new_n17323_));
  NOR2_X1    g14887(.A1(new_n13344_), .A2(pi0173), .ZN(new_n17324_));
  OAI21_X1   g14888(.A1(new_n14125_), .A2(new_n17324_), .B(new_n16263_), .ZN(new_n17325_));
  OAI21_X1   g14889(.A1(new_n14122_), .A2(new_n10736_), .B(new_n3265_), .ZN(new_n17326_));
  NAND2_X1   g14890(.A1(new_n17326_), .A2(new_n2609_), .ZN(new_n17327_));
  NAND2_X1   g14891(.A1(new_n15744_), .A2(new_n10736_), .ZN(new_n17328_));
  AOI21_X1   g14892(.A1(new_n17328_), .A2(new_n17327_), .B(new_n17325_), .ZN(new_n17329_));
  NAND2_X1   g14893(.A1(new_n2609_), .A2(new_n16263_), .ZN(new_n17330_));
  AOI21_X1   g14894(.A1(new_n17323_), .A2(new_n17330_), .B(new_n17329_), .ZN(new_n17331_));
  NAND2_X1   g14895(.A1(new_n17331_), .A2(new_n13521_), .ZN(new_n17332_));
  NOR2_X1    g14896(.A1(new_n17323_), .A2(new_n13521_), .ZN(new_n17333_));
  INV_X1     g14897(.I(new_n17333_), .ZN(new_n17334_));
  AOI21_X1   g14898(.A1(new_n17332_), .A2(new_n17334_), .B(pi1153), .ZN(new_n17335_));
  NAND2_X1   g14899(.A1(new_n17320_), .A2(new_n13521_), .ZN(new_n17336_));
  NAND2_X1   g14900(.A1(new_n17331_), .A2(pi0625), .ZN(new_n17337_));
  AOI21_X1   g14901(.A1(new_n17337_), .A2(new_n17336_), .B(new_n12841_), .ZN(new_n17338_));
  NOR3_X1    g14902(.A1(new_n17335_), .A2(new_n17338_), .A3(new_n12758_), .ZN(new_n17339_));
  NOR2_X1    g14903(.A1(new_n17331_), .A2(pi0778), .ZN(new_n17340_));
  NOR2_X1    g14904(.A1(new_n17339_), .A2(new_n17340_), .ZN(new_n17341_));
  OAI21_X1   g14905(.A1(new_n17341_), .A2(new_n12869_), .B(new_n17322_), .ZN(new_n17342_));
  INV_X1     g14906(.I(new_n17342_), .ZN(new_n17343_));
  NOR2_X1    g14907(.A1(new_n17323_), .A2(new_n12888_), .ZN(new_n17344_));
  AOI21_X1   g14908(.A1(new_n17343_), .A2(new_n12888_), .B(new_n17344_), .ZN(new_n17345_));
  NOR2_X1    g14909(.A1(new_n17345_), .A2(new_n14288_), .ZN(new_n17346_));
  AOI21_X1   g14910(.A1(new_n14288_), .A2(new_n17320_), .B(new_n17346_), .ZN(new_n17347_));
  NOR2_X1    g14911(.A1(new_n17347_), .A2(pi0628), .ZN(new_n17348_));
  NOR2_X1    g14912(.A1(new_n17323_), .A2(new_n12920_), .ZN(new_n17349_));
  OAI21_X1   g14913(.A1(new_n17348_), .A2(new_n17349_), .B(new_n12742_), .ZN(new_n17350_));
  NOR2_X1    g14914(.A1(new_n17323_), .A2(pi0628), .ZN(new_n17351_));
  NOR2_X1    g14915(.A1(new_n17347_), .A2(new_n12920_), .ZN(new_n17352_));
  OAI21_X1   g14916(.A1(new_n17352_), .A2(new_n17351_), .B(pi1156), .ZN(new_n17353_));
  NAND3_X1   g14917(.A1(new_n17350_), .A2(new_n17353_), .A3(pi0792), .ZN(new_n17354_));
  NAND2_X1   g14918(.A1(new_n17347_), .A2(new_n12937_), .ZN(new_n17355_));
  NAND2_X1   g14919(.A1(new_n17354_), .A2(new_n17355_), .ZN(new_n17356_));
  NAND2_X1   g14920(.A1(new_n17356_), .A2(pi0647), .ZN(new_n17357_));
  OAI21_X1   g14921(.A1(pi0647), .A2(new_n17320_), .B(new_n17357_), .ZN(new_n17358_));
  NAND2_X1   g14922(.A1(new_n17356_), .A2(new_n12741_), .ZN(new_n17359_));
  OAI21_X1   g14923(.A1(new_n12741_), .A2(new_n17320_), .B(new_n17359_), .ZN(new_n17360_));
  OAI22_X1   g14924(.A1(new_n15576_), .A2(new_n17358_), .B1(new_n17360_), .B2(new_n15730_), .ZN(new_n17361_));
  NOR2_X1    g14925(.A1(new_n2609_), .A2(new_n10736_), .ZN(new_n17362_));
  INV_X1     g14926(.I(new_n17324_), .ZN(new_n17363_));
  AOI21_X1   g14927(.A1(new_n13341_), .A2(new_n16245_), .B(new_n3265_), .ZN(new_n17364_));
  NOR2_X1    g14928(.A1(new_n13334_), .A2(pi0173), .ZN(new_n17365_));
  AOI22_X1   g14929(.A1(new_n17365_), .A2(new_n16245_), .B1(pi0173), .B2(new_n15784_), .ZN(new_n17366_));
  OAI21_X1   g14930(.A1(new_n15787_), .A2(pi0173), .B(pi0745), .ZN(new_n17367_));
  NAND2_X1   g14931(.A1(new_n17366_), .A2(new_n17367_), .ZN(new_n17368_));
  AOI22_X1   g14932(.A1(new_n17368_), .A2(new_n3265_), .B1(new_n17363_), .B2(new_n17364_), .ZN(new_n17369_));
  NOR2_X1    g14933(.A1(new_n17369_), .A2(new_n2610_), .ZN(new_n17370_));
  NOR2_X1    g14934(.A1(new_n17370_), .A2(new_n17362_), .ZN(new_n17371_));
  NOR2_X1    g14935(.A1(new_n17371_), .A2(new_n12760_), .ZN(new_n17372_));
  AOI21_X1   g14936(.A1(new_n12760_), .A2(new_n17320_), .B(new_n17372_), .ZN(new_n17373_));
  INV_X1     g14937(.I(new_n17372_), .ZN(new_n17374_));
  OAI22_X1   g14938(.A1(new_n17374_), .A2(pi0609), .B1(new_n13353_), .B2(new_n17323_), .ZN(new_n17375_));
  NAND2_X1   g14939(.A1(new_n17375_), .A2(new_n12770_), .ZN(new_n17376_));
  OAI22_X1   g14940(.A1(new_n17374_), .A2(new_n12766_), .B1(new_n12772_), .B2(new_n17323_), .ZN(new_n17377_));
  AOI21_X1   g14941(.A1(new_n17377_), .A2(pi1155), .B(new_n12764_), .ZN(new_n17378_));
  AOI22_X1   g14942(.A1(new_n17378_), .A2(new_n17376_), .B1(new_n12764_), .B2(new_n17373_), .ZN(new_n17379_));
  NAND2_X1   g14943(.A1(new_n17323_), .A2(new_n15804_), .ZN(new_n17380_));
  OAI22_X1   g14944(.A1(new_n17379_), .A2(new_n15803_), .B1(new_n12779_), .B2(new_n17380_), .ZN(new_n17381_));
  NOR2_X1    g14945(.A1(new_n17320_), .A2(new_n15807_), .ZN(new_n17382_));
  AOI22_X1   g14946(.A1(new_n17381_), .A2(new_n15779_), .B1(pi0789), .B2(new_n17382_), .ZN(new_n17383_));
  OAI22_X1   g14947(.A1(new_n17383_), .A2(new_n12803_), .B1(new_n12749_), .B2(new_n17320_), .ZN(new_n17384_));
  NAND2_X1   g14948(.A1(new_n17384_), .A2(pi0788), .ZN(new_n17385_));
  OAI21_X1   g14949(.A1(pi0788), .A2(new_n17383_), .B(new_n17385_), .ZN(new_n17386_));
  NOR2_X1    g14950(.A1(new_n17386_), .A2(new_n12943_), .ZN(new_n17387_));
  AOI21_X1   g14951(.A1(new_n12943_), .A2(new_n17320_), .B(new_n17387_), .ZN(new_n17388_));
  INV_X1     g14952(.I(new_n17388_), .ZN(new_n17389_));
  AOI21_X1   g14953(.A1(new_n15608_), .A2(new_n17389_), .B(new_n17361_), .ZN(new_n17390_));
  AND2_X2    g14954(.A1(new_n17353_), .A2(new_n12919_), .Z(new_n17391_));
  AOI21_X1   g14955(.A1(pi0629), .A2(new_n17350_), .B(new_n17391_), .ZN(new_n17392_));
  NOR2_X1    g14956(.A1(new_n17386_), .A2(new_n15821_), .ZN(new_n17393_));
  OAI21_X1   g14957(.A1(new_n17392_), .A2(new_n17393_), .B(pi0792), .ZN(new_n17394_));
  INV_X1     g14958(.I(new_n17362_), .ZN(new_n17395_));
  AOI21_X1   g14959(.A1(new_n16245_), .A2(new_n13566_), .B(new_n15826_), .ZN(new_n17396_));
  AOI21_X1   g14960(.A1(new_n14328_), .A2(new_n17216_), .B(new_n10736_), .ZN(new_n17397_));
  AOI21_X1   g14961(.A1(new_n17397_), .A2(new_n5336_), .B(new_n3265_), .ZN(new_n17398_));
  OAI21_X1   g14962(.A1(new_n17396_), .A2(pi0173), .B(new_n17398_), .ZN(new_n17399_));
  NAND2_X1   g14963(.A1(new_n14172_), .A2(pi0173), .ZN(new_n17400_));
  NAND2_X1   g14964(.A1(new_n14174_), .A2(new_n10736_), .ZN(new_n17401_));
  AOI21_X1   g14965(.A1(new_n17400_), .A2(new_n17401_), .B(pi0745), .ZN(new_n17402_));
  NAND2_X1   g14966(.A1(new_n15835_), .A2(pi0173), .ZN(new_n17403_));
  NAND2_X1   g14967(.A1(new_n14177_), .A2(new_n10736_), .ZN(new_n17404_));
  AOI21_X1   g14968(.A1(new_n17404_), .A2(new_n17403_), .B(new_n16245_), .ZN(new_n17405_));
  OAI21_X1   g14969(.A1(new_n17405_), .A2(new_n17402_), .B(new_n2627_), .ZN(new_n17406_));
  NOR2_X1    g14970(.A1(new_n14182_), .A2(pi0173), .ZN(new_n17407_));
  NOR2_X1    g14971(.A1(new_n14184_), .A2(new_n10736_), .ZN(new_n17408_));
  OAI21_X1   g14972(.A1(new_n17407_), .A2(new_n17408_), .B(pi0745), .ZN(new_n17409_));
  NOR2_X1    g14973(.A1(new_n14187_), .A2(new_n10736_), .ZN(new_n17410_));
  NOR2_X1    g14974(.A1(new_n14189_), .A2(pi0173), .ZN(new_n17411_));
  OAI21_X1   g14975(.A1(new_n17410_), .A2(new_n17411_), .B(new_n16245_), .ZN(new_n17412_));
  NAND3_X1   g14976(.A1(new_n17412_), .A2(new_n17409_), .A3(pi0039), .ZN(new_n17413_));
  NAND3_X1   g14977(.A1(new_n17413_), .A2(new_n3265_), .A3(new_n17406_), .ZN(new_n17414_));
  NAND3_X1   g14978(.A1(new_n17414_), .A2(new_n16263_), .A3(new_n17399_), .ZN(new_n17415_));
  NAND2_X1   g14979(.A1(new_n17369_), .A2(pi0723), .ZN(new_n17416_));
  NAND3_X1   g14980(.A1(new_n17416_), .A2(new_n17415_), .A3(new_n2609_), .ZN(new_n17417_));
  NAND2_X1   g14981(.A1(new_n17417_), .A2(new_n17395_), .ZN(new_n17418_));
  NAND2_X1   g14982(.A1(new_n17418_), .A2(new_n12758_), .ZN(new_n17419_));
  INV_X1     g14983(.I(new_n17338_), .ZN(new_n17420_));
  NOR2_X1    g14984(.A1(new_n17371_), .A2(new_n13521_), .ZN(new_n17421_));
  AOI21_X1   g14985(.A1(new_n17418_), .A2(new_n13521_), .B(new_n17421_), .ZN(new_n17422_));
  OAI21_X1   g14986(.A1(new_n17422_), .A2(pi1153), .B(new_n17420_), .ZN(new_n17423_));
  NOR2_X1    g14987(.A1(new_n17371_), .A2(pi0625), .ZN(new_n17424_));
  AOI21_X1   g14988(.A1(new_n17418_), .A2(pi0625), .B(new_n17424_), .ZN(new_n17425_));
  OAI21_X1   g14989(.A1(new_n17425_), .A2(new_n12841_), .B(pi0608), .ZN(new_n17426_));
  OAI22_X1   g14990(.A1(pi0608), .A2(new_n17423_), .B1(new_n17426_), .B2(new_n17335_), .ZN(new_n17427_));
  OAI21_X1   g14991(.A1(new_n17427_), .A2(new_n12758_), .B(new_n17419_), .ZN(new_n17428_));
  INV_X1     g14992(.I(new_n17428_), .ZN(new_n17429_));
  INV_X1     g14993(.I(new_n17341_), .ZN(new_n17430_));
  NOR2_X1    g14994(.A1(new_n17430_), .A2(pi0609), .ZN(new_n17431_));
  INV_X1     g14995(.I(new_n17431_), .ZN(new_n17432_));
  NAND2_X1   g14996(.A1(new_n17428_), .A2(pi0609), .ZN(new_n17433_));
  NAND2_X1   g14997(.A1(new_n17433_), .A2(new_n17432_), .ZN(new_n17434_));
  NAND2_X1   g14998(.A1(new_n17434_), .A2(pi1155), .ZN(new_n17435_));
  NAND3_X1   g14999(.A1(new_n17435_), .A2(pi0660), .A3(new_n17376_), .ZN(new_n17436_));
  NAND2_X1   g15000(.A1(new_n17377_), .A2(pi1155), .ZN(new_n17437_));
  NOR2_X1    g15001(.A1(new_n17429_), .A2(pi0609), .ZN(new_n17438_));
  NOR2_X1    g15002(.A1(new_n17430_), .A2(new_n12766_), .ZN(new_n17439_));
  OAI21_X1   g15003(.A1(new_n17438_), .A2(new_n17439_), .B(new_n12770_), .ZN(new_n17440_));
  NAND3_X1   g15004(.A1(new_n17440_), .A2(new_n13829_), .A3(new_n17437_), .ZN(new_n17441_));
  NAND3_X1   g15005(.A1(new_n17441_), .A2(new_n17436_), .A3(pi0785), .ZN(new_n17442_));
  OAI21_X1   g15006(.A1(pi0785), .A2(new_n17429_), .B(new_n17442_), .ZN(new_n17443_));
  AOI21_X1   g15007(.A1(new_n17323_), .A2(pi0618), .B(pi1154), .ZN(new_n17444_));
  OAI21_X1   g15008(.A1(new_n17379_), .A2(pi0618), .B(new_n17444_), .ZN(new_n17445_));
  AND2_X2    g15009(.A1(new_n17445_), .A2(pi0627), .Z(new_n17446_));
  OAI21_X1   g15010(.A1(new_n17343_), .A2(pi0618), .B(pi1154), .ZN(new_n17447_));
  NOR2_X1    g15011(.A1(new_n17443_), .A2(new_n12781_), .ZN(new_n17448_));
  OAI21_X1   g15012(.A1(new_n17448_), .A2(new_n17447_), .B(new_n17446_), .ZN(new_n17449_));
  AOI21_X1   g15013(.A1(new_n17323_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n17450_));
  OAI21_X1   g15014(.A1(new_n17379_), .A2(new_n12781_), .B(new_n17450_), .ZN(new_n17451_));
  AND2_X2    g15015(.A1(new_n17451_), .A2(new_n12880_), .Z(new_n17452_));
  AOI21_X1   g15016(.A1(new_n17342_), .A2(pi0618), .B(pi1154), .ZN(new_n17453_));
  OAI21_X1   g15017(.A1(new_n17443_), .A2(pi0618), .B(new_n17453_), .ZN(new_n17454_));
  AOI21_X1   g15018(.A1(new_n17454_), .A2(new_n17452_), .B(new_n12779_), .ZN(new_n17455_));
  AOI22_X1   g15019(.A1(new_n17455_), .A2(new_n17449_), .B1(new_n12779_), .B2(new_n17443_), .ZN(new_n17456_));
  NOR2_X1    g15020(.A1(new_n17456_), .A2(pi0789), .ZN(new_n17457_));
  NOR2_X1    g15021(.A1(new_n17457_), .A2(new_n14303_), .ZN(new_n17458_));
  OAI21_X1   g15022(.A1(new_n17320_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n17459_));
  AND2_X2    g15023(.A1(new_n17381_), .A2(new_n12793_), .Z(new_n17460_));
  OAI21_X1   g15024(.A1(new_n17460_), .A2(new_n17459_), .B(pi0648), .ZN(new_n17461_));
  AOI21_X1   g15025(.A1(new_n17345_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n17462_));
  NAND2_X1   g15026(.A1(new_n17456_), .A2(pi0619), .ZN(new_n17463_));
  AOI21_X1   g15027(.A1(new_n17463_), .A2(new_n17462_), .B(new_n17461_), .ZN(new_n17464_));
  OAI21_X1   g15028(.A1(new_n17320_), .A2(pi0619), .B(pi1159), .ZN(new_n17465_));
  AND2_X2    g15029(.A1(new_n17381_), .A2(pi0619), .Z(new_n17466_));
  OAI21_X1   g15030(.A1(new_n17466_), .A2(new_n17465_), .B(new_n12895_), .ZN(new_n17467_));
  NAND2_X1   g15031(.A1(new_n17345_), .A2(pi0619), .ZN(new_n17468_));
  NAND2_X1   g15032(.A1(new_n17468_), .A2(new_n12791_), .ZN(new_n17469_));
  AOI21_X1   g15033(.A1(new_n17456_), .A2(new_n12793_), .B(new_n17469_), .ZN(new_n17470_));
  OAI21_X1   g15034(.A1(new_n17470_), .A2(new_n17467_), .B(pi0789), .ZN(new_n17471_));
  OAI21_X1   g15035(.A1(new_n17471_), .A2(new_n17464_), .B(new_n17458_), .ZN(new_n17472_));
  NAND2_X1   g15036(.A1(new_n17345_), .A2(new_n12911_), .ZN(new_n17473_));
  NAND2_X1   g15037(.A1(new_n17323_), .A2(new_n12910_), .ZN(new_n17474_));
  AOI21_X1   g15038(.A1(new_n17473_), .A2(new_n17474_), .B(new_n12906_), .ZN(new_n17475_));
  AND2_X2    g15039(.A1(new_n17384_), .A2(new_n12914_), .Z(new_n17476_));
  OAI21_X1   g15040(.A1(new_n17476_), .A2(new_n17475_), .B(pi0788), .ZN(new_n17477_));
  NAND3_X1   g15041(.A1(new_n17472_), .A2(new_n15824_), .A3(new_n17477_), .ZN(new_n17478_));
  AND2_X2    g15042(.A1(new_n17478_), .A2(new_n17394_), .Z(new_n17479_));
  OAI22_X1   g15043(.A1(new_n17479_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n17390_), .ZN(new_n17480_));
  AOI21_X1   g15044(.A1(new_n17323_), .A2(new_n12975_), .B(pi0715), .ZN(new_n17481_));
  NOR2_X1    g15045(.A1(new_n17323_), .A2(new_n12985_), .ZN(new_n17482_));
  AOI21_X1   g15046(.A1(new_n17389_), .A2(new_n12985_), .B(new_n17482_), .ZN(new_n17483_));
  NAND2_X1   g15047(.A1(new_n17483_), .A2(pi0644), .ZN(new_n17484_));
  AOI21_X1   g15048(.A1(new_n17484_), .A2(new_n17481_), .B(new_n12739_), .ZN(new_n17485_));
  AOI21_X1   g15049(.A1(new_n17485_), .A2(pi0644), .B(new_n13000_), .ZN(new_n17486_));
  NOR2_X1    g15050(.A1(new_n17480_), .A2(new_n17486_), .ZN(new_n17487_));
  NOR2_X1    g15051(.A1(new_n17360_), .A2(pi1157), .ZN(new_n17488_));
  NOR2_X1    g15052(.A1(new_n17358_), .A2(new_n12965_), .ZN(new_n17489_));
  OAI21_X1   g15053(.A1(new_n17488_), .A2(new_n17489_), .B(pi0787), .ZN(new_n17490_));
  OAI21_X1   g15054(.A1(pi0787), .A2(new_n17356_), .B(new_n17490_), .ZN(new_n17491_));
  OAI21_X1   g15055(.A1(new_n17491_), .A2(pi0644), .B(pi0715), .ZN(new_n17492_));
  NAND2_X1   g15056(.A1(new_n17492_), .A2(new_n17485_), .ZN(new_n17493_));
  AND2_X2    g15057(.A1(new_n17491_), .A2(pi0644), .Z(new_n17494_));
  AOI21_X1   g15058(.A1(new_n17480_), .A2(new_n12975_), .B(new_n17494_), .ZN(new_n17495_));
  AOI21_X1   g15059(.A1(new_n17323_), .A2(pi0644), .B(new_n12740_), .ZN(new_n17496_));
  NAND2_X1   g15060(.A1(new_n17483_), .A2(new_n12975_), .ZN(new_n17497_));
  AOI21_X1   g15061(.A1(new_n17497_), .A2(new_n17496_), .B(pi1160), .ZN(new_n17498_));
  OAI21_X1   g15062(.A1(new_n17495_), .A2(pi0715), .B(new_n17498_), .ZN(new_n17499_));
  AOI21_X1   g15063(.A1(new_n17499_), .A2(new_n17493_), .B(new_n13000_), .ZN(new_n17500_));
  OAI21_X1   g15064(.A1(new_n17500_), .A2(new_n17487_), .B(new_n6643_), .ZN(new_n17501_));
  AOI22_X1   g15065(.A1(new_n17501_), .A2(new_n17319_), .B1(pi0832), .B2(new_n17318_), .ZN(po0330));
  NOR2_X1    g15066(.A1(new_n3042_), .A2(new_n7488_), .ZN(new_n17503_));
  INV_X1     g15067(.I(new_n12818_), .ZN(new_n17504_));
  NOR2_X1    g15068(.A1(new_n13340_), .A2(new_n16296_), .ZN(new_n17505_));
  INV_X1     g15069(.I(new_n17505_), .ZN(new_n17506_));
  NOR2_X1    g15070(.A1(new_n17506_), .A2(new_n15232_), .ZN(new_n17507_));
  INV_X1     g15071(.I(new_n17507_), .ZN(new_n17508_));
  NOR2_X1    g15072(.A1(new_n17508_), .A2(new_n15246_), .ZN(new_n17509_));
  NAND2_X1   g15073(.A1(new_n17509_), .A2(new_n17504_), .ZN(new_n17510_));
  NOR3_X1    g15074(.A1(new_n17510_), .A2(new_n12981_), .A3(new_n12943_), .ZN(new_n17511_));
  INV_X1     g15075(.I(new_n17503_), .ZN(new_n17512_));
  NAND2_X1   g15076(.A1(new_n12826_), .A2(pi0696), .ZN(new_n17513_));
  NAND2_X1   g15077(.A1(new_n17513_), .A2(new_n17512_), .ZN(new_n17514_));
  INV_X1     g15078(.I(new_n17514_), .ZN(new_n17515_));
  NOR2_X1    g15079(.A1(new_n17513_), .A2(new_n13521_), .ZN(new_n17516_));
  NOR3_X1    g15080(.A1(new_n17516_), .A2(new_n12841_), .A3(new_n17503_), .ZN(new_n17517_));
  INV_X1     g15081(.I(new_n17517_), .ZN(new_n17518_));
  OAI21_X1   g15082(.A1(new_n17515_), .A2(new_n17516_), .B(new_n12841_), .ZN(new_n17519_));
  NAND3_X1   g15083(.A1(new_n17518_), .A2(new_n17519_), .A3(pi0778), .ZN(new_n17520_));
  OAI21_X1   g15084(.A1(pi0778), .A2(new_n17515_), .B(new_n17520_), .ZN(new_n17521_));
  AND2_X2    g15085(.A1(new_n17521_), .A2(new_n14291_), .Z(new_n17522_));
  NAND2_X1   g15086(.A1(new_n17522_), .A2(new_n12952_), .ZN(new_n17523_));
  AOI21_X1   g15087(.A1(new_n17523_), .A2(new_n12981_), .B(new_n12741_), .ZN(new_n17524_));
  NOR3_X1    g15088(.A1(new_n17524_), .A2(new_n12965_), .A3(new_n17511_), .ZN(new_n17525_));
  NOR2_X1    g15089(.A1(new_n17510_), .A2(pi0630), .ZN(new_n17526_));
  AOI21_X1   g15090(.A1(new_n17526_), .A2(new_n13384_), .B(new_n12741_), .ZN(new_n17527_));
  AOI21_X1   g15091(.A1(new_n17522_), .A2(new_n12952_), .B(new_n12981_), .ZN(new_n17528_));
  NOR2_X1    g15092(.A1(new_n17528_), .A2(new_n17527_), .ZN(new_n17529_));
  NOR2_X1    g15093(.A1(new_n17529_), .A2(pi1157), .ZN(new_n17530_));
  OAI21_X1   g15094(.A1(new_n17530_), .A2(new_n17525_), .B(pi0787), .ZN(new_n17531_));
  NAND2_X1   g15095(.A1(new_n17522_), .A2(pi0628), .ZN(new_n17532_));
  NAND2_X1   g15096(.A1(new_n17510_), .A2(new_n12920_), .ZN(new_n17533_));
  AOI21_X1   g15097(.A1(new_n17533_), .A2(pi0629), .B(new_n12742_), .ZN(new_n17534_));
  NAND2_X1   g15098(.A1(new_n17510_), .A2(pi0628), .ZN(new_n17535_));
  AOI22_X1   g15099(.A1(new_n17522_), .A2(new_n12920_), .B1(new_n12919_), .B2(new_n17535_), .ZN(new_n17536_));
  AOI22_X1   g15100(.A1(new_n17536_), .A2(new_n12742_), .B1(new_n17532_), .B2(new_n17534_), .ZN(new_n17537_));
  NOR2_X1    g15101(.A1(new_n17537_), .A2(new_n17503_), .ZN(new_n17538_));
  AOI21_X1   g15102(.A1(new_n17509_), .A2(pi0626), .B(new_n17503_), .ZN(new_n17539_));
  NAND2_X1   g15103(.A1(new_n17521_), .A2(new_n14289_), .ZN(new_n17540_));
  OAI21_X1   g15104(.A1(new_n17540_), .A2(new_n12910_), .B(new_n17512_), .ZN(new_n17541_));
  AOI21_X1   g15105(.A1(new_n17541_), .A2(new_n12748_), .B(pi0641), .ZN(new_n17542_));
  OAI21_X1   g15106(.A1(new_n12745_), .A2(new_n17539_), .B(new_n17542_), .ZN(new_n17543_));
  AOI21_X1   g15107(.A1(new_n17509_), .A2(new_n12747_), .B(new_n17503_), .ZN(new_n17544_));
  OR2_X2     g15108(.A1(new_n17544_), .A2(pi1158), .Z(new_n17545_));
  AOI21_X1   g15109(.A1(new_n17541_), .A2(new_n12746_), .B(new_n12814_), .ZN(new_n17546_));
  AOI21_X1   g15110(.A1(new_n17546_), .A2(new_n17545_), .B(new_n12808_), .ZN(new_n17547_));
  AOI21_X1   g15111(.A1(new_n17543_), .A2(new_n17547_), .B(new_n15340_), .ZN(new_n17548_));
  NOR2_X1    g15112(.A1(new_n17521_), .A2(pi0609), .ZN(new_n17549_));
  NOR2_X1    g15113(.A1(new_n14328_), .A2(new_n16325_), .ZN(new_n17550_));
  NOR3_X1    g15114(.A1(new_n17550_), .A2(new_n17505_), .A3(new_n17503_), .ZN(new_n17551_));
  NAND2_X1   g15115(.A1(new_n17551_), .A2(new_n12758_), .ZN(new_n17552_));
  NOR2_X1    g15116(.A1(new_n14330_), .A2(new_n16325_), .ZN(new_n17553_));
  INV_X1     g15117(.I(new_n17553_), .ZN(new_n17554_));
  NAND4_X1   g15118(.A1(new_n17554_), .A2(pi1153), .A3(new_n17512_), .A4(new_n17506_), .ZN(new_n17555_));
  NAND3_X1   g15119(.A1(new_n17555_), .A2(pi0608), .A3(new_n17519_), .ZN(new_n17556_));
  OAI21_X1   g15120(.A1(new_n17553_), .A2(new_n17551_), .B(new_n12841_), .ZN(new_n17557_));
  NAND3_X1   g15121(.A1(new_n17557_), .A2(new_n13560_), .A3(new_n17518_), .ZN(new_n17558_));
  NAND3_X1   g15122(.A1(new_n17556_), .A2(pi0778), .A3(new_n17558_), .ZN(new_n17559_));
  AOI21_X1   g15123(.A1(new_n17559_), .A2(new_n17552_), .B(new_n12766_), .ZN(new_n17560_));
  OAI21_X1   g15124(.A1(new_n17560_), .A2(new_n17549_), .B(pi1155), .ZN(new_n17561_));
  NAND2_X1   g15125(.A1(new_n17505_), .A2(new_n13353_), .ZN(new_n17562_));
  NAND3_X1   g15126(.A1(new_n17562_), .A2(new_n12770_), .A3(new_n17512_), .ZN(new_n17563_));
  NAND3_X1   g15127(.A1(new_n17561_), .A2(pi0660), .A3(new_n17563_), .ZN(new_n17564_));
  NAND2_X1   g15128(.A1(new_n17559_), .A2(new_n17552_), .ZN(new_n17565_));
  NOR2_X1    g15129(.A1(new_n17521_), .A2(new_n12766_), .ZN(new_n17566_));
  AOI21_X1   g15130(.A1(new_n17565_), .A2(new_n12766_), .B(new_n17566_), .ZN(new_n17567_));
  AOI21_X1   g15131(.A1(new_n17505_), .A2(new_n12772_), .B(new_n12770_), .ZN(new_n17568_));
  AOI21_X1   g15132(.A1(new_n17568_), .A2(new_n17512_), .B(pi0660), .ZN(new_n17569_));
  OAI21_X1   g15133(.A1(new_n17567_), .A2(pi1155), .B(new_n17569_), .ZN(new_n17570_));
  NAND3_X1   g15134(.A1(new_n17564_), .A2(new_n17570_), .A3(pi0785), .ZN(new_n17571_));
  NAND2_X1   g15135(.A1(new_n17565_), .A2(new_n12764_), .ZN(new_n17572_));
  NAND2_X1   g15136(.A1(new_n17571_), .A2(new_n17572_), .ZN(new_n17573_));
  NAND2_X1   g15137(.A1(new_n17573_), .A2(pi0618), .ZN(new_n17574_));
  AOI21_X1   g15138(.A1(new_n17521_), .A2(new_n12870_), .B(new_n17503_), .ZN(new_n17575_));
  NAND2_X1   g15139(.A1(new_n17575_), .A2(new_n12781_), .ZN(new_n17576_));
  AOI21_X1   g15140(.A1(new_n17574_), .A2(new_n17576_), .B(new_n12785_), .ZN(new_n17577_));
  OAI21_X1   g15141(.A1(new_n17508_), .A2(new_n15304_), .B(new_n12785_), .ZN(new_n17578_));
  NOR2_X1    g15142(.A1(new_n17578_), .A2(new_n17503_), .ZN(new_n17579_));
  NOR3_X1    g15143(.A1(new_n17577_), .A2(new_n12880_), .A3(new_n17579_), .ZN(new_n17580_));
  NAND2_X1   g15144(.A1(new_n17575_), .A2(pi0618), .ZN(new_n17581_));
  NAND2_X1   g15145(.A1(new_n17573_), .A2(new_n12781_), .ZN(new_n17582_));
  NAND2_X1   g15146(.A1(new_n17582_), .A2(new_n17581_), .ZN(new_n17583_));
  OAI21_X1   g15147(.A1(new_n17508_), .A2(new_n15311_), .B(pi1154), .ZN(new_n17584_));
  OAI21_X1   g15148(.A1(new_n17584_), .A2(new_n17503_), .B(new_n12880_), .ZN(new_n17585_));
  AOI21_X1   g15149(.A1(new_n17583_), .A2(new_n12785_), .B(new_n17585_), .ZN(new_n17586_));
  NOR3_X1    g15150(.A1(new_n17580_), .A2(new_n17586_), .A3(new_n12779_), .ZN(new_n17587_));
  AOI21_X1   g15151(.A1(new_n17571_), .A2(new_n17572_), .B(pi0781), .ZN(new_n17588_));
  NAND2_X1   g15152(.A1(new_n12909_), .A2(new_n15807_), .ZN(new_n17589_));
  INV_X1     g15153(.I(new_n17589_), .ZN(new_n17590_));
  NOR2_X1    g15154(.A1(new_n17590_), .A2(new_n12796_), .ZN(new_n17591_));
  INV_X1     g15155(.I(new_n17591_), .ZN(new_n17592_));
  OAI21_X1   g15156(.A1(new_n17587_), .A2(new_n17588_), .B(new_n17592_), .ZN(new_n17593_));
  NAND3_X1   g15157(.A1(new_n17507_), .A2(new_n15240_), .A3(pi0619), .ZN(new_n17594_));
  NAND2_X1   g15158(.A1(new_n17507_), .A2(new_n15271_), .ZN(new_n17595_));
  AOI22_X1   g15159(.A1(new_n17594_), .A2(new_n12907_), .B1(new_n17595_), .B2(new_n12908_), .ZN(new_n17596_));
  NAND3_X1   g15160(.A1(new_n12793_), .A2(pi0648), .A3(pi1159), .ZN(new_n17597_));
  NAND3_X1   g15161(.A1(new_n12895_), .A2(new_n12791_), .A3(pi0619), .ZN(new_n17598_));
  NAND2_X1   g15162(.A1(new_n17598_), .A2(new_n17597_), .ZN(new_n17599_));
  NAND2_X1   g15163(.A1(new_n17540_), .A2(new_n17599_), .ZN(new_n17600_));
  AOI21_X1   g15164(.A1(new_n17600_), .A2(new_n17596_), .B(new_n12796_), .ZN(new_n17601_));
  AOI21_X1   g15165(.A1(new_n17601_), .A2(new_n17512_), .B(new_n14303_), .ZN(new_n17602_));
  NAND2_X1   g15166(.A1(new_n17593_), .A2(new_n17602_), .ZN(new_n17603_));
  AOI22_X1   g15167(.A1(new_n17603_), .A2(new_n17548_), .B1(pi0792), .B2(new_n17538_), .ZN(new_n17604_));
  OAI22_X1   g15168(.A1(new_n17604_), .A2(new_n15341_), .B1(new_n17503_), .B2(new_n17531_), .ZN(new_n17605_));
  NAND2_X1   g15169(.A1(new_n17605_), .A2(new_n13000_), .ZN(new_n17606_));
  AND2_X2    g15170(.A1(new_n17605_), .A2(new_n12975_), .Z(new_n17607_));
  OAI21_X1   g15171(.A1(new_n17523_), .A2(new_n14300_), .B(new_n17512_), .ZN(new_n17608_));
  NOR2_X1    g15172(.A1(new_n17608_), .A2(new_n12975_), .ZN(new_n17609_));
  OAI21_X1   g15173(.A1(new_n17607_), .A2(new_n17609_), .B(new_n12740_), .ZN(new_n17610_));
  NOR2_X1    g15174(.A1(new_n12943_), .A2(new_n12984_), .ZN(new_n17611_));
  INV_X1     g15175(.I(new_n17611_), .ZN(new_n17612_));
  NOR2_X1    g15176(.A1(new_n17510_), .A2(new_n17612_), .ZN(new_n17613_));
  NAND2_X1   g15177(.A1(new_n17613_), .A2(new_n12975_), .ZN(new_n17614_));
  NAND3_X1   g15178(.A1(new_n17614_), .A2(pi0715), .A3(new_n17512_), .ZN(new_n17615_));
  NAND3_X1   g15179(.A1(new_n17610_), .A2(new_n12739_), .A3(new_n17615_), .ZN(new_n17616_));
  NOR2_X1    g15180(.A1(new_n17608_), .A2(pi0644), .ZN(new_n17617_));
  AOI21_X1   g15181(.A1(new_n17605_), .A2(pi0644), .B(new_n17617_), .ZN(new_n17618_));
  AOI21_X1   g15182(.A1(new_n17613_), .A2(pi0644), .B(pi0715), .ZN(new_n17619_));
  AOI21_X1   g15183(.A1(new_n17619_), .A2(new_n17512_), .B(new_n12739_), .ZN(new_n17620_));
  OAI21_X1   g15184(.A1(new_n17618_), .A2(new_n12740_), .B(new_n17620_), .ZN(new_n17621_));
  NAND3_X1   g15185(.A1(new_n17616_), .A2(pi0790), .A3(new_n17621_), .ZN(new_n17622_));
  AOI21_X1   g15186(.A1(new_n17622_), .A2(new_n17606_), .B(new_n12738_), .ZN(new_n17623_));
  AOI21_X1   g15187(.A1(pi0057), .A2(pi0174), .B(pi0832), .ZN(new_n17624_));
  NAND2_X1   g15188(.A1(new_n13192_), .A2(pi0174), .ZN(new_n17625_));
  NOR2_X1    g15189(.A1(new_n17625_), .A2(new_n13521_), .ZN(new_n17626_));
  NOR2_X1    g15190(.A1(new_n2610_), .A2(new_n16325_), .ZN(new_n17627_));
  NOR2_X1    g15191(.A1(new_n14122_), .A2(pi0174), .ZN(new_n17628_));
  NOR2_X1    g15192(.A1(new_n14118_), .A2(new_n7488_), .ZN(new_n17629_));
  OAI21_X1   g15193(.A1(new_n17629_), .A2(new_n17628_), .B(new_n3265_), .ZN(new_n17630_));
  NOR2_X1    g15194(.A1(new_n13344_), .A2(new_n7488_), .ZN(new_n17631_));
  NOR2_X1    g15195(.A1(new_n13398_), .A2(new_n17631_), .ZN(new_n17632_));
  NOR2_X1    g15196(.A1(new_n17632_), .A2(new_n3265_), .ZN(new_n17633_));
  INV_X1     g15197(.I(new_n17633_), .ZN(new_n17634_));
  NAND3_X1   g15198(.A1(new_n17630_), .A2(new_n17627_), .A3(new_n17634_), .ZN(new_n17635_));
  INV_X1     g15199(.I(new_n17627_), .ZN(new_n17636_));
  NAND2_X1   g15200(.A1(new_n17625_), .A2(new_n17636_), .ZN(new_n17637_));
  AND3_X2    g15201(.A1(new_n17635_), .A2(new_n13521_), .A3(new_n17637_), .Z(new_n17638_));
  OAI21_X1   g15202(.A1(new_n17638_), .A2(new_n17626_), .B(new_n12841_), .ZN(new_n17639_));
  NAND3_X1   g15203(.A1(new_n17635_), .A2(new_n17637_), .A3(pi0625), .ZN(new_n17640_));
  INV_X1     g15204(.I(new_n17625_), .ZN(new_n17641_));
  NAND2_X1   g15205(.A1(new_n17641_), .A2(new_n13521_), .ZN(new_n17642_));
  AOI21_X1   g15206(.A1(new_n17640_), .A2(new_n17642_), .B(new_n12841_), .ZN(new_n17643_));
  NOR2_X1    g15207(.A1(new_n17643_), .A2(new_n12758_), .ZN(new_n17644_));
  AOI21_X1   g15208(.A1(new_n17635_), .A2(new_n17637_), .B(pi0778), .ZN(new_n17645_));
  AOI21_X1   g15209(.A1(new_n17644_), .A2(new_n17639_), .B(new_n17645_), .ZN(new_n17646_));
  NOR2_X1    g15210(.A1(new_n17625_), .A2(new_n12870_), .ZN(new_n17647_));
  AOI21_X1   g15211(.A1(new_n17646_), .A2(new_n12870_), .B(new_n17647_), .ZN(new_n17648_));
  NOR2_X1    g15212(.A1(new_n17641_), .A2(new_n12888_), .ZN(new_n17649_));
  AOI21_X1   g15213(.A1(new_n17648_), .A2(new_n12888_), .B(new_n17649_), .ZN(new_n17650_));
  NOR2_X1    g15214(.A1(new_n17625_), .A2(new_n12911_), .ZN(new_n17651_));
  AOI21_X1   g15215(.A1(new_n17650_), .A2(new_n12911_), .B(new_n17651_), .ZN(new_n17652_));
  NOR2_X1    g15216(.A1(new_n17641_), .A2(new_n13392_), .ZN(new_n17653_));
  AOI21_X1   g15217(.A1(new_n17652_), .A2(new_n13392_), .B(new_n17653_), .ZN(new_n17654_));
  NAND2_X1   g15218(.A1(new_n17654_), .A2(new_n12920_), .ZN(new_n17655_));
  NAND2_X1   g15219(.A1(new_n17641_), .A2(pi0628), .ZN(new_n17656_));
  AOI21_X1   g15220(.A1(new_n17655_), .A2(new_n17656_), .B(pi1156), .ZN(new_n17657_));
  OR2_X2     g15221(.A1(new_n17657_), .A2(new_n12919_), .Z(new_n17658_));
  NOR2_X1    g15222(.A1(new_n2609_), .A2(new_n7488_), .ZN(new_n17659_));
  INV_X1     g15223(.I(new_n17659_), .ZN(new_n17660_));
  NOR2_X1    g15224(.A1(new_n5337_), .A2(new_n17506_), .ZN(new_n17661_));
  OAI21_X1   g15225(.A1(new_n17631_), .A2(new_n17661_), .B(pi0038), .ZN(new_n17662_));
  INV_X1     g15226(.I(new_n17662_), .ZN(new_n17663_));
  NAND3_X1   g15227(.A1(new_n13245_), .A2(new_n7488_), .A3(pi0759), .ZN(new_n17664_));
  NAND2_X1   g15228(.A1(new_n13256_), .A2(pi0759), .ZN(new_n17665_));
  NAND2_X1   g15229(.A1(new_n13060_), .A2(new_n16296_), .ZN(new_n17666_));
  AOI21_X1   g15230(.A1(new_n17665_), .A2(new_n17666_), .B(pi0039), .ZN(new_n17667_));
  AOI21_X1   g15231(.A1(new_n13322_), .A2(new_n13332_), .B(new_n16296_), .ZN(new_n17668_));
  NOR3_X1    g15232(.A1(new_n13178_), .A2(new_n13188_), .A3(pi0759), .ZN(new_n17669_));
  NOR3_X1    g15233(.A1(new_n17668_), .A2(new_n17669_), .A3(new_n2627_), .ZN(new_n17670_));
  OAI21_X1   g15234(.A1(new_n17670_), .A2(new_n17667_), .B(pi0174), .ZN(new_n17671_));
  AOI21_X1   g15235(.A1(new_n17671_), .A2(new_n17664_), .B(pi0038), .ZN(new_n17672_));
  OAI21_X1   g15236(.A1(new_n17672_), .A2(new_n17663_), .B(new_n2609_), .ZN(new_n17673_));
  NAND2_X1   g15237(.A1(new_n17673_), .A2(new_n17660_), .ZN(new_n17674_));
  NAND2_X1   g15238(.A1(new_n17674_), .A2(new_n12761_), .ZN(new_n17675_));
  OAI21_X1   g15239(.A1(new_n12761_), .A2(new_n17625_), .B(new_n17675_), .ZN(new_n17676_));
  NOR2_X1    g15240(.A1(new_n17625_), .A2(new_n12766_), .ZN(new_n17677_));
  AOI21_X1   g15241(.A1(new_n17676_), .A2(new_n12766_), .B(new_n17677_), .ZN(new_n17678_));
  NOR2_X1    g15242(.A1(new_n17678_), .A2(pi1155), .ZN(new_n17679_));
  NOR2_X1    g15243(.A1(new_n17625_), .A2(pi0609), .ZN(new_n17680_));
  AOI21_X1   g15244(.A1(new_n17676_), .A2(pi0609), .B(new_n17680_), .ZN(new_n17681_));
  OAI21_X1   g15245(.A1(new_n17681_), .A2(new_n12770_), .B(pi0785), .ZN(new_n17682_));
  OAI22_X1   g15246(.A1(new_n17682_), .A2(new_n17679_), .B1(pi0785), .B2(new_n17676_), .ZN(new_n17683_));
  NAND2_X1   g15247(.A1(new_n17641_), .A2(pi0618), .ZN(new_n17684_));
  OAI21_X1   g15248(.A1(new_n17683_), .A2(pi0618), .B(new_n17684_), .ZN(new_n17685_));
  NAND2_X1   g15249(.A1(new_n17685_), .A2(new_n12785_), .ZN(new_n17686_));
  NAND2_X1   g15250(.A1(new_n17641_), .A2(new_n12781_), .ZN(new_n17687_));
  OAI21_X1   g15251(.A1(new_n17683_), .A2(new_n12781_), .B(new_n17687_), .ZN(new_n17688_));
  AOI21_X1   g15252(.A1(new_n17688_), .A2(pi1154), .B(new_n12779_), .ZN(new_n17689_));
  AOI22_X1   g15253(.A1(new_n17689_), .A2(new_n17686_), .B1(new_n12779_), .B2(new_n17683_), .ZN(new_n17690_));
  NOR2_X1    g15254(.A1(new_n17690_), .A2(pi0789), .ZN(new_n17691_));
  NOR2_X1    g15255(.A1(new_n17625_), .A2(new_n12793_), .ZN(new_n17692_));
  AOI21_X1   g15256(.A1(new_n17690_), .A2(new_n12793_), .B(new_n17692_), .ZN(new_n17693_));
  NOR2_X1    g15257(.A1(new_n17693_), .A2(pi1159), .ZN(new_n17694_));
  NOR2_X1    g15258(.A1(new_n17625_), .A2(pi0619), .ZN(new_n17695_));
  AOI21_X1   g15259(.A1(new_n17690_), .A2(pi0619), .B(new_n17695_), .ZN(new_n17696_));
  NOR2_X1    g15260(.A1(new_n17696_), .A2(new_n12791_), .ZN(new_n17697_));
  NOR3_X1    g15261(.A1(new_n17694_), .A2(new_n17697_), .A3(new_n12796_), .ZN(new_n17698_));
  NOR2_X1    g15262(.A1(new_n17698_), .A2(new_n17691_), .ZN(new_n17699_));
  NOR2_X1    g15263(.A1(new_n17699_), .A2(new_n12818_), .ZN(new_n17700_));
  AOI21_X1   g15264(.A1(new_n12818_), .A2(new_n17625_), .B(new_n17700_), .ZN(new_n17701_));
  NOR2_X1    g15265(.A1(new_n17701_), .A2(pi0628), .ZN(new_n17702_));
  NOR2_X1    g15266(.A1(new_n17702_), .A2(new_n12742_), .ZN(new_n17703_));
  AOI21_X1   g15267(.A1(new_n17641_), .A2(new_n12747_), .B(pi0641), .ZN(new_n17704_));
  INV_X1     g15268(.I(new_n17704_), .ZN(new_n17705_));
  NOR3_X1    g15269(.A1(new_n17698_), .A2(new_n12747_), .A3(new_n17691_), .ZN(new_n17706_));
  OAI21_X1   g15270(.A1(new_n17706_), .A2(new_n17705_), .B(pi1158), .ZN(new_n17707_));
  INV_X1     g15271(.I(new_n17652_), .ZN(new_n17708_));
  AOI21_X1   g15272(.A1(new_n17708_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n17709_));
  NOR3_X1    g15273(.A1(new_n17663_), .A2(new_n16325_), .A3(new_n15123_), .ZN(new_n17710_));
  AOI21_X1   g15274(.A1(new_n13692_), .A2(pi0174), .B(new_n16296_), .ZN(new_n17711_));
  OAI21_X1   g15275(.A1(new_n14187_), .A2(pi0174), .B(new_n17711_), .ZN(new_n17712_));
  OAI21_X1   g15276(.A1(new_n13794_), .A2(new_n13786_), .B(new_n7488_), .ZN(new_n17713_));
  OAI21_X1   g15277(.A1(new_n13745_), .A2(new_n13754_), .B(pi0174), .ZN(new_n17714_));
  NAND3_X1   g15278(.A1(new_n17714_), .A2(new_n16296_), .A3(new_n17713_), .ZN(new_n17715_));
  NAND3_X1   g15279(.A1(new_n17712_), .A2(new_n17715_), .A3(pi0039), .ZN(new_n17716_));
  AOI21_X1   g15280(.A1(new_n13416_), .A2(new_n13798_), .B(pi0174), .ZN(new_n17717_));
  NOR2_X1    g15281(.A1(new_n13800_), .A2(new_n7488_), .ZN(new_n17718_));
  OAI21_X1   g15282(.A1(new_n17718_), .A2(new_n17717_), .B(pi0759), .ZN(new_n17719_));
  NOR3_X1    g15283(.A1(new_n13809_), .A2(new_n13406_), .A3(new_n7488_), .ZN(new_n17720_));
  AOI21_X1   g15284(.A1(new_n13805_), .A2(new_n13807_), .B(pi0174), .ZN(new_n17721_));
  OAI21_X1   g15285(.A1(new_n17720_), .A2(new_n17721_), .B(new_n16296_), .ZN(new_n17722_));
  NAND3_X1   g15286(.A1(new_n17719_), .A2(new_n17722_), .A3(new_n2627_), .ZN(new_n17723_));
  NAND3_X1   g15287(.A1(new_n17716_), .A2(new_n17723_), .A3(new_n3265_), .ZN(new_n17724_));
  AOI21_X1   g15288(.A1(new_n17724_), .A2(new_n17710_), .B(new_n2610_), .ZN(new_n17725_));
  OR3_X2     g15289(.A1(new_n17672_), .A2(pi0696), .A3(new_n17663_), .Z(new_n17726_));
  AOI21_X1   g15290(.A1(new_n17725_), .A2(new_n17726_), .B(new_n17659_), .ZN(new_n17727_));
  NOR2_X1    g15291(.A1(new_n17727_), .A2(new_n13521_), .ZN(new_n17728_));
  AOI21_X1   g15292(.A1(new_n17673_), .A2(new_n17660_), .B(pi0625), .ZN(new_n17729_));
  OAI21_X1   g15293(.A1(new_n17728_), .A2(new_n17729_), .B(pi1153), .ZN(new_n17730_));
  NAND3_X1   g15294(.A1(new_n17730_), .A2(pi0608), .A3(new_n17639_), .ZN(new_n17731_));
  NAND2_X1   g15295(.A1(new_n17674_), .A2(pi0625), .ZN(new_n17732_));
  OAI21_X1   g15296(.A1(new_n17727_), .A2(pi0625), .B(new_n17732_), .ZN(new_n17733_));
  AOI21_X1   g15297(.A1(new_n17733_), .A2(new_n12841_), .B(new_n17643_), .ZN(new_n17734_));
  AOI21_X1   g15298(.A1(new_n17734_), .A2(new_n13560_), .B(new_n12758_), .ZN(new_n17735_));
  NOR2_X1    g15299(.A1(new_n17727_), .A2(pi0778), .ZN(new_n17736_));
  AOI21_X1   g15300(.A1(new_n17735_), .A2(new_n17731_), .B(new_n17736_), .ZN(new_n17737_));
  NOR2_X1    g15301(.A1(new_n17737_), .A2(pi0785), .ZN(new_n17738_));
  INV_X1     g15302(.I(new_n17738_), .ZN(new_n17739_));
  NOR2_X1    g15303(.A1(new_n17679_), .A2(new_n13829_), .ZN(new_n17740_));
  INV_X1     g15304(.I(new_n17740_), .ZN(new_n17741_));
  INV_X1     g15305(.I(new_n17646_), .ZN(new_n17742_));
  AOI21_X1   g15306(.A1(new_n17742_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n17743_));
  NAND2_X1   g15307(.A1(new_n17737_), .A2(pi0609), .ZN(new_n17744_));
  AOI21_X1   g15308(.A1(new_n17744_), .A2(new_n17743_), .B(new_n17741_), .ZN(new_n17745_));
  OAI21_X1   g15309(.A1(new_n17681_), .A2(new_n12770_), .B(new_n13829_), .ZN(new_n17746_));
  OAI21_X1   g15310(.A1(new_n17646_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n17747_));
  AOI21_X1   g15311(.A1(new_n17737_), .A2(new_n12766_), .B(new_n17747_), .ZN(new_n17748_));
  OAI21_X1   g15312(.A1(new_n17748_), .A2(new_n17746_), .B(pi0785), .ZN(new_n17749_));
  OAI21_X1   g15313(.A1(new_n17749_), .A2(new_n17745_), .B(new_n17739_), .ZN(new_n17750_));
  NAND2_X1   g15314(.A1(new_n17750_), .A2(new_n12779_), .ZN(new_n17751_));
  INV_X1     g15315(.I(new_n17751_), .ZN(new_n17752_));
  AOI21_X1   g15316(.A1(new_n17685_), .A2(new_n12785_), .B(new_n12880_), .ZN(new_n17753_));
  AOI21_X1   g15317(.A1(new_n17648_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n17754_));
  OAI21_X1   g15318(.A1(new_n17750_), .A2(new_n12781_), .B(new_n17754_), .ZN(new_n17755_));
  NAND2_X1   g15319(.A1(new_n17755_), .A2(new_n17753_), .ZN(new_n17756_));
  AOI21_X1   g15320(.A1(new_n17688_), .A2(pi1154), .B(pi0627), .ZN(new_n17757_));
  AOI21_X1   g15321(.A1(new_n17648_), .A2(pi0618), .B(pi1154), .ZN(new_n17758_));
  OAI21_X1   g15322(.A1(new_n17750_), .A2(pi0618), .B(new_n17758_), .ZN(new_n17759_));
  AOI21_X1   g15323(.A1(new_n17759_), .A2(new_n17757_), .B(new_n12779_), .ZN(new_n17760_));
  AOI21_X1   g15324(.A1(new_n17760_), .A2(new_n17756_), .B(new_n17752_), .ZN(new_n17761_));
  NOR2_X1    g15325(.A1(new_n17761_), .A2(pi0789), .ZN(new_n17762_));
  INV_X1     g15326(.I(new_n17762_), .ZN(new_n17763_));
  OAI21_X1   g15327(.A1(new_n17693_), .A2(pi1159), .B(pi0648), .ZN(new_n17764_));
  INV_X1     g15328(.I(new_n17650_), .ZN(new_n17765_));
  AOI21_X1   g15329(.A1(new_n17765_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n17766_));
  NAND2_X1   g15330(.A1(new_n17761_), .A2(pi0619), .ZN(new_n17767_));
  AOI21_X1   g15331(.A1(new_n17767_), .A2(new_n17766_), .B(new_n17764_), .ZN(new_n17768_));
  NOR2_X1    g15332(.A1(new_n17697_), .A2(pi0648), .ZN(new_n17769_));
  INV_X1     g15333(.I(new_n17769_), .ZN(new_n17770_));
  AOI21_X1   g15334(.A1(new_n17765_), .A2(pi0619), .B(pi1159), .ZN(new_n17771_));
  INV_X1     g15335(.I(new_n17771_), .ZN(new_n17772_));
  AOI21_X1   g15336(.A1(new_n17761_), .A2(new_n12793_), .B(new_n17772_), .ZN(new_n17773_));
  OAI21_X1   g15337(.A1(new_n17773_), .A2(new_n17770_), .B(pi0789), .ZN(new_n17774_));
  OAI21_X1   g15338(.A1(new_n17774_), .A2(new_n17768_), .B(new_n17763_), .ZN(new_n17775_));
  NAND2_X1   g15339(.A1(new_n17775_), .A2(pi0626), .ZN(new_n17776_));
  AOI21_X1   g15340(.A1(new_n17776_), .A2(new_n17709_), .B(new_n17707_), .ZN(new_n17777_));
  AOI21_X1   g15341(.A1(new_n17641_), .A2(pi0626), .B(new_n12814_), .ZN(new_n17778_));
  NAND2_X1   g15342(.A1(new_n17699_), .A2(new_n12747_), .ZN(new_n17779_));
  NAND2_X1   g15343(.A1(new_n17779_), .A2(new_n17778_), .ZN(new_n17780_));
  NAND2_X1   g15344(.A1(new_n17780_), .A2(new_n12745_), .ZN(new_n17781_));
  AOI21_X1   g15345(.A1(new_n17708_), .A2(pi0626), .B(pi0641), .ZN(new_n17782_));
  INV_X1     g15346(.I(new_n17782_), .ZN(new_n17783_));
  AOI21_X1   g15347(.A1(new_n17775_), .A2(new_n12747_), .B(new_n17783_), .ZN(new_n17784_));
  OAI21_X1   g15348(.A1(new_n17784_), .A2(new_n17781_), .B(pi0788), .ZN(new_n17785_));
  OR2_X2     g15349(.A1(new_n17775_), .A2(pi0788), .Z(new_n17786_));
  OAI21_X1   g15350(.A1(new_n17785_), .A2(new_n17777_), .B(new_n17786_), .ZN(new_n17787_));
  NAND2_X1   g15351(.A1(new_n17787_), .A2(pi0628), .ZN(new_n17788_));
  AOI21_X1   g15352(.A1(new_n17788_), .A2(new_n17703_), .B(new_n17658_), .ZN(new_n17789_));
  NOR2_X1    g15353(.A1(new_n17625_), .A2(pi0628), .ZN(new_n17790_));
  AOI21_X1   g15354(.A1(new_n17654_), .A2(pi0628), .B(new_n17790_), .ZN(new_n17791_));
  OAI21_X1   g15355(.A1(new_n17791_), .A2(new_n12742_), .B(new_n12919_), .ZN(new_n17792_));
  OAI21_X1   g15356(.A1(new_n17701_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n17793_));
  AOI21_X1   g15357(.A1(new_n17787_), .A2(new_n12920_), .B(new_n17793_), .ZN(new_n17794_));
  OAI21_X1   g15358(.A1(new_n17794_), .A2(new_n17792_), .B(pi0792), .ZN(new_n17795_));
  OR2_X2     g15359(.A1(new_n17787_), .A2(pi0792), .Z(new_n17796_));
  OAI21_X1   g15360(.A1(new_n17795_), .A2(new_n17789_), .B(new_n17796_), .ZN(new_n17797_));
  AND2_X2    g15361(.A1(new_n17797_), .A2(new_n12972_), .Z(new_n17798_));
  NOR2_X1    g15362(.A1(new_n17654_), .A2(pi0792), .ZN(new_n17799_));
  OAI21_X1   g15363(.A1(new_n17791_), .A2(new_n12742_), .B(pi0792), .ZN(new_n17800_));
  NOR2_X1    g15364(.A1(new_n17800_), .A2(new_n17657_), .ZN(new_n17801_));
  NOR2_X1    g15365(.A1(new_n17801_), .A2(new_n17799_), .ZN(new_n17802_));
  NAND2_X1   g15366(.A1(new_n17802_), .A2(new_n12741_), .ZN(new_n17803_));
  NAND2_X1   g15367(.A1(new_n17641_), .A2(pi0647), .ZN(new_n17804_));
  AOI21_X1   g15368(.A1(new_n17803_), .A2(new_n17804_), .B(pi1157), .ZN(new_n17805_));
  NOR2_X1    g15369(.A1(new_n17805_), .A2(new_n12981_), .ZN(new_n17806_));
  NAND2_X1   g15370(.A1(new_n17625_), .A2(new_n12943_), .ZN(new_n17807_));
  OAI21_X1   g15371(.A1(new_n17701_), .A2(new_n12943_), .B(new_n17807_), .ZN(new_n17808_));
  AOI21_X1   g15372(.A1(new_n17808_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n17809_));
  OAI21_X1   g15373(.A1(new_n17797_), .A2(new_n12741_), .B(new_n17809_), .ZN(new_n17810_));
  NAND2_X1   g15374(.A1(new_n17810_), .A2(new_n17806_), .ZN(new_n17811_));
  NOR2_X1    g15375(.A1(new_n17625_), .A2(pi0647), .ZN(new_n17812_));
  AOI21_X1   g15376(.A1(new_n17802_), .A2(pi0647), .B(new_n17812_), .ZN(new_n17813_));
  NOR2_X1    g15377(.A1(new_n17813_), .A2(new_n12965_), .ZN(new_n17814_));
  NOR2_X1    g15378(.A1(new_n17814_), .A2(pi0630), .ZN(new_n17815_));
  AOI21_X1   g15379(.A1(new_n17808_), .A2(pi0647), .B(pi1157), .ZN(new_n17816_));
  OAI21_X1   g15380(.A1(new_n17797_), .A2(pi0647), .B(new_n17816_), .ZN(new_n17817_));
  AOI21_X1   g15381(.A1(new_n17817_), .A2(new_n17815_), .B(new_n12972_), .ZN(new_n17818_));
  AOI21_X1   g15382(.A1(new_n17818_), .A2(new_n17811_), .B(new_n17798_), .ZN(new_n17819_));
  OAI21_X1   g15383(.A1(new_n17819_), .A2(pi0790), .B(new_n5477_), .ZN(new_n17820_));
  OAI21_X1   g15384(.A1(new_n17641_), .A2(new_n12975_), .B(pi0715), .ZN(new_n17821_));
  NAND2_X1   g15385(.A1(new_n17641_), .A2(new_n12984_), .ZN(new_n17822_));
  OAI21_X1   g15386(.A1(new_n17808_), .A2(new_n12984_), .B(new_n17822_), .ZN(new_n17823_));
  NOR2_X1    g15387(.A1(new_n17823_), .A2(pi0644), .ZN(new_n17824_));
  OAI21_X1   g15388(.A1(new_n17824_), .A2(new_n17821_), .B(new_n12739_), .ZN(new_n17825_));
  NOR2_X1    g15389(.A1(new_n17814_), .A2(new_n12972_), .ZN(new_n17826_));
  INV_X1     g15390(.I(new_n17826_), .ZN(new_n17827_));
  OAI22_X1   g15391(.A1(new_n17827_), .A2(new_n17805_), .B1(pi0787), .B2(new_n17802_), .ZN(new_n17828_));
  AOI21_X1   g15392(.A1(new_n17828_), .A2(pi0644), .B(pi0715), .ZN(new_n17829_));
  NAND2_X1   g15393(.A1(new_n17819_), .A2(new_n12975_), .ZN(new_n17830_));
  AOI21_X1   g15394(.A1(new_n17830_), .A2(new_n17829_), .B(new_n17825_), .ZN(new_n17831_));
  OAI21_X1   g15395(.A1(new_n17641_), .A2(pi0644), .B(new_n12740_), .ZN(new_n17832_));
  NOR2_X1    g15396(.A1(new_n17823_), .A2(new_n12975_), .ZN(new_n17833_));
  OAI21_X1   g15397(.A1(new_n17833_), .A2(new_n17832_), .B(pi1160), .ZN(new_n17834_));
  NAND2_X1   g15398(.A1(new_n17828_), .A2(new_n12975_), .ZN(new_n17835_));
  NAND2_X1   g15399(.A1(new_n17835_), .A2(pi0715), .ZN(new_n17836_));
  AOI21_X1   g15400(.A1(new_n17819_), .A2(pi0644), .B(new_n17836_), .ZN(new_n17837_));
  OAI21_X1   g15401(.A1(new_n17837_), .A2(new_n17834_), .B(pi0790), .ZN(new_n17838_));
  NOR2_X1    g15402(.A1(new_n17838_), .A2(new_n17831_), .ZN(new_n17839_));
  AOI21_X1   g15403(.A1(new_n6165_), .A2(new_n7488_), .B(pi0057), .ZN(new_n17840_));
  OAI21_X1   g15404(.A1(new_n17839_), .A2(new_n17820_), .B(new_n17840_), .ZN(new_n17841_));
  AOI21_X1   g15405(.A1(new_n17841_), .A2(new_n17624_), .B(new_n17623_), .ZN(po0331));
  NOR2_X1    g15406(.A1(new_n3042_), .A2(pi0175), .ZN(new_n17843_));
  NOR2_X1    g15407(.A1(new_n13340_), .A2(new_n16384_), .ZN(new_n17844_));
  NOR2_X1    g15408(.A1(new_n17844_), .A2(new_n17843_), .ZN(new_n17845_));
  NOR3_X1    g15409(.A1(new_n17845_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n17846_));
  INV_X1     g15410(.I(new_n17844_), .ZN(new_n17847_));
  NOR2_X1    g15411(.A1(new_n17847_), .A2(new_n13354_), .ZN(new_n17848_));
  NOR3_X1    g15412(.A1(new_n17848_), .A2(new_n12762_), .A3(new_n17845_), .ZN(new_n17849_));
  NOR2_X1    g15413(.A1(new_n17849_), .A2(new_n12770_), .ZN(new_n17850_));
  NOR3_X1    g15414(.A1(new_n17848_), .A2(pi1155), .A3(new_n17843_), .ZN(new_n17851_));
  NOR3_X1    g15415(.A1(new_n17850_), .A2(new_n12764_), .A3(new_n17851_), .ZN(new_n17852_));
  NOR2_X1    g15416(.A1(new_n17852_), .A2(new_n17846_), .ZN(new_n17853_));
  NOR2_X1    g15417(.A1(new_n17853_), .A2(pi0781), .ZN(new_n17854_));
  INV_X1     g15418(.I(new_n17853_), .ZN(new_n17855_));
  AOI21_X1   g15419(.A1(new_n17855_), .A2(new_n12783_), .B(pi1154), .ZN(new_n17856_));
  AOI21_X1   g15420(.A1(new_n17855_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n17857_));
  NOR3_X1    g15421(.A1(new_n17856_), .A2(new_n17857_), .A3(new_n12779_), .ZN(new_n17858_));
  NOR2_X1    g15422(.A1(new_n17858_), .A2(new_n17854_), .ZN(new_n17859_));
  NOR2_X1    g15423(.A1(new_n17859_), .A2(new_n17229_), .ZN(new_n17860_));
  NOR2_X1    g15424(.A1(new_n17860_), .A2(pi1159), .ZN(new_n17861_));
  OAI21_X1   g15425(.A1(new_n17859_), .A2(new_n17232_), .B(pi1159), .ZN(new_n17862_));
  NAND2_X1   g15426(.A1(new_n17862_), .A2(pi0789), .ZN(new_n17863_));
  OAI22_X1   g15427(.A1(new_n17863_), .A2(new_n17861_), .B1(pi0789), .B2(new_n17859_), .ZN(new_n17864_));
  INV_X1     g15428(.I(new_n17843_), .ZN(new_n17865_));
  NAND2_X1   g15429(.A1(new_n12818_), .A2(new_n17865_), .ZN(new_n17866_));
  OAI21_X1   g15430(.A1(new_n17864_), .A2(new_n12818_), .B(new_n17866_), .ZN(new_n17867_));
  AOI21_X1   g15431(.A1(new_n12826_), .A2(pi0700), .B(new_n17843_), .ZN(new_n17868_));
  INV_X1     g15432(.I(pi0700), .ZN(new_n17869_));
  NOR2_X1    g15433(.A1(new_n12834_), .A2(new_n17869_), .ZN(new_n17870_));
  INV_X1     g15434(.I(new_n17870_), .ZN(new_n17871_));
  NOR2_X1    g15435(.A1(new_n17843_), .A2(pi1153), .ZN(new_n17872_));
  NAND2_X1   g15436(.A1(new_n17871_), .A2(new_n17872_), .ZN(new_n17873_));
  NOR2_X1    g15437(.A1(new_n17870_), .A2(new_n17868_), .ZN(new_n17874_));
  NOR2_X1    g15438(.A1(new_n17874_), .A2(new_n12841_), .ZN(new_n17875_));
  INV_X1     g15439(.I(new_n17875_), .ZN(new_n17876_));
  NAND3_X1   g15440(.A1(new_n17876_), .A2(pi0778), .A3(new_n17873_), .ZN(new_n17877_));
  OAI21_X1   g15441(.A1(pi0778), .A2(new_n17868_), .B(new_n17877_), .ZN(new_n17878_));
  NAND2_X1   g15442(.A1(new_n17878_), .A2(new_n17187_), .ZN(new_n17879_));
  NOR2_X1    g15443(.A1(new_n17879_), .A2(new_n12889_), .ZN(new_n17880_));
  INV_X1     g15444(.I(new_n17880_), .ZN(new_n17881_));
  NOR2_X1    g15445(.A1(new_n17881_), .A2(new_n12912_), .ZN(new_n17882_));
  INV_X1     g15446(.I(new_n17882_), .ZN(new_n17883_));
  NOR2_X1    g15447(.A1(new_n13392_), .A2(new_n3043_), .ZN(new_n17884_));
  NOR2_X1    g15448(.A1(new_n17883_), .A2(new_n17884_), .ZN(new_n17885_));
  INV_X1     g15449(.I(new_n17885_), .ZN(new_n17886_));
  OAI22_X1   g15450(.A1(new_n17867_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n17886_), .ZN(new_n17887_));
  NAND2_X1   g15451(.A1(new_n17887_), .A2(new_n12919_), .ZN(new_n17888_));
  OAI22_X1   g15452(.A1(new_n17867_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n17886_), .ZN(new_n17889_));
  NAND2_X1   g15453(.A1(new_n17889_), .A2(pi0629), .ZN(new_n17890_));
  AOI21_X1   g15454(.A1(new_n17888_), .A2(new_n17890_), .B(new_n12937_), .ZN(new_n17891_));
  INV_X1     g15455(.I(new_n17851_), .ZN(new_n17892_));
  NOR2_X1    g15456(.A1(new_n17868_), .A2(new_n12754_), .ZN(new_n17893_));
  NOR3_X1    g15457(.A1(new_n17893_), .A2(new_n17843_), .A3(new_n17844_), .ZN(new_n17894_));
  NAND2_X1   g15458(.A1(new_n17894_), .A2(new_n12758_), .ZN(new_n17895_));
  NAND2_X1   g15459(.A1(new_n17893_), .A2(pi0625), .ZN(new_n17896_));
  NAND3_X1   g15460(.A1(new_n17896_), .A2(pi1153), .A3(new_n17845_), .ZN(new_n17897_));
  NAND3_X1   g15461(.A1(new_n17873_), .A2(pi0608), .A3(new_n17897_), .ZN(new_n17898_));
  INV_X1     g15462(.I(new_n17896_), .ZN(new_n17899_));
  OAI21_X1   g15463(.A1(new_n17899_), .A2(new_n17894_), .B(new_n17872_), .ZN(new_n17900_));
  NAND3_X1   g15464(.A1(new_n17876_), .A2(new_n13560_), .A3(new_n17900_), .ZN(new_n17901_));
  NAND3_X1   g15465(.A1(new_n17901_), .A2(pi0778), .A3(new_n17898_), .ZN(new_n17902_));
  AOI21_X1   g15466(.A1(new_n17902_), .A2(new_n17895_), .B(new_n12766_), .ZN(new_n17903_));
  NOR2_X1    g15467(.A1(new_n17878_), .A2(pi0609), .ZN(new_n17904_));
  OAI21_X1   g15468(.A1(new_n17904_), .A2(new_n17903_), .B(pi1155), .ZN(new_n17905_));
  NAND3_X1   g15469(.A1(new_n17905_), .A2(pi0660), .A3(new_n17892_), .ZN(new_n17906_));
  NAND2_X1   g15470(.A1(new_n17902_), .A2(new_n17895_), .ZN(new_n17907_));
  NOR2_X1    g15471(.A1(new_n17878_), .A2(new_n12766_), .ZN(new_n17908_));
  AOI21_X1   g15472(.A1(new_n17907_), .A2(new_n12766_), .B(new_n17908_), .ZN(new_n17909_));
  NOR2_X1    g15473(.A1(new_n17850_), .A2(pi0660), .ZN(new_n17910_));
  OAI21_X1   g15474(.A1(new_n17909_), .A2(pi1155), .B(new_n17910_), .ZN(new_n17911_));
  NAND3_X1   g15475(.A1(new_n17911_), .A2(new_n17906_), .A3(pi0785), .ZN(new_n17912_));
  NAND2_X1   g15476(.A1(new_n17907_), .A2(new_n12764_), .ZN(new_n17913_));
  NAND2_X1   g15477(.A1(new_n17912_), .A2(new_n17913_), .ZN(new_n17914_));
  NAND2_X1   g15478(.A1(new_n17914_), .A2(new_n12781_), .ZN(new_n17915_));
  NAND2_X1   g15479(.A1(new_n17879_), .A2(pi0618), .ZN(new_n17916_));
  AOI21_X1   g15480(.A1(new_n17915_), .A2(new_n17916_), .B(pi1154), .ZN(new_n17917_));
  NOR3_X1    g15481(.A1(new_n17917_), .A2(pi0627), .A3(new_n17857_), .ZN(new_n17918_));
  NAND2_X1   g15482(.A1(new_n17879_), .A2(new_n12781_), .ZN(new_n17919_));
  NAND2_X1   g15483(.A1(new_n17914_), .A2(pi0618), .ZN(new_n17920_));
  AOI21_X1   g15484(.A1(new_n17920_), .A2(new_n17919_), .B(new_n12785_), .ZN(new_n17921_));
  NOR3_X1    g15485(.A1(new_n17921_), .A2(new_n12880_), .A3(new_n17856_), .ZN(new_n17922_));
  OR3_X2     g15486(.A1(new_n17918_), .A2(new_n17922_), .A3(new_n12779_), .Z(new_n17923_));
  NAND2_X1   g15487(.A1(new_n17914_), .A2(new_n12779_), .ZN(new_n17924_));
  NAND2_X1   g15488(.A1(new_n17923_), .A2(new_n17924_), .ZN(new_n17925_));
  AOI21_X1   g15489(.A1(new_n17925_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n17926_));
  NAND2_X1   g15490(.A1(new_n17881_), .A2(new_n12793_), .ZN(new_n17927_));
  NAND2_X1   g15491(.A1(new_n17925_), .A2(pi0619), .ZN(new_n17928_));
  AOI21_X1   g15492(.A1(new_n17928_), .A2(new_n17927_), .B(new_n12791_), .ZN(new_n17929_));
  NOR3_X1    g15493(.A1(new_n17929_), .A2(new_n12895_), .A3(new_n17861_), .ZN(new_n17930_));
  AOI21_X1   g15494(.A1(new_n17923_), .A2(new_n17924_), .B(pi0619), .ZN(new_n17931_));
  NOR2_X1    g15495(.A1(new_n17880_), .A2(new_n12793_), .ZN(new_n17932_));
  OAI21_X1   g15496(.A1(new_n17931_), .A2(new_n17932_), .B(new_n12791_), .ZN(new_n17933_));
  NAND3_X1   g15497(.A1(new_n17933_), .A2(new_n12895_), .A3(new_n17862_), .ZN(new_n17934_));
  NAND2_X1   g15498(.A1(new_n17934_), .A2(pi0789), .ZN(new_n17935_));
  OAI21_X1   g15499(.A1(new_n17935_), .A2(new_n17930_), .B(new_n17926_), .ZN(new_n17936_));
  NAND2_X1   g15500(.A1(new_n17843_), .A2(pi0626), .ZN(new_n17937_));
  NAND2_X1   g15501(.A1(new_n17864_), .A2(new_n12747_), .ZN(new_n17938_));
  AOI21_X1   g15502(.A1(new_n17938_), .A2(new_n17937_), .B(new_n12816_), .ZN(new_n17939_));
  NOR2_X1    g15503(.A1(new_n17865_), .A2(pi0626), .ZN(new_n17940_));
  AOI21_X1   g15504(.A1(new_n17864_), .A2(pi0626), .B(new_n17940_), .ZN(new_n17941_));
  OAI22_X1   g15505(.A1(new_n17941_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n17883_), .ZN(new_n17942_));
  OAI21_X1   g15506(.A1(new_n17942_), .A2(new_n17939_), .B(pi0788), .ZN(new_n17943_));
  AOI21_X1   g15507(.A1(new_n17936_), .A2(new_n17943_), .B(new_n15340_), .ZN(new_n17944_));
  OR2_X2     g15508(.A1(new_n17944_), .A2(new_n17891_), .Z(new_n17945_));
  NAND2_X1   g15509(.A1(new_n17867_), .A2(new_n13384_), .ZN(new_n17946_));
  NAND2_X1   g15510(.A1(new_n12943_), .A2(new_n17865_), .ZN(new_n17947_));
  AOI21_X1   g15511(.A1(new_n17946_), .A2(new_n17947_), .B(new_n17212_), .ZN(new_n17948_));
  NOR2_X1    g15512(.A1(new_n17886_), .A2(new_n12953_), .ZN(new_n17949_));
  NOR2_X1    g15513(.A1(new_n17949_), .A2(pi0647), .ZN(new_n17950_));
  NOR2_X1    g15514(.A1(new_n17843_), .A2(new_n12741_), .ZN(new_n17951_));
  OAI21_X1   g15515(.A1(new_n17950_), .A2(new_n17951_), .B(new_n12965_), .ZN(new_n17952_));
  NOR2_X1    g15516(.A1(new_n17865_), .A2(pi0647), .ZN(new_n17953_));
  AOI21_X1   g15517(.A1(new_n17949_), .A2(pi0647), .B(new_n17953_), .ZN(new_n17954_));
  INV_X1     g15518(.I(new_n17954_), .ZN(new_n17955_));
  OAI22_X1   g15519(.A1(new_n17952_), .A2(new_n12981_), .B1(new_n17955_), .B2(new_n15576_), .ZN(new_n17956_));
  NOR2_X1    g15520(.A1(new_n17956_), .A2(new_n17948_), .ZN(new_n17957_));
  OAI22_X1   g15521(.A1(new_n17945_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n17957_), .ZN(new_n17958_));
  OAI21_X1   g15522(.A1(new_n12965_), .A2(new_n17955_), .B(new_n17952_), .ZN(new_n17959_));
  NOR2_X1    g15523(.A1(new_n17959_), .A2(new_n12972_), .ZN(new_n17960_));
  AOI21_X1   g15524(.A1(new_n12972_), .A2(new_n17949_), .B(new_n17960_), .ZN(new_n17961_));
  AND2_X2    g15525(.A1(new_n17961_), .A2(pi0644), .Z(new_n17962_));
  AOI21_X1   g15526(.A1(new_n17958_), .A2(new_n12975_), .B(new_n17962_), .ZN(new_n17963_));
  NAND2_X1   g15527(.A1(new_n17865_), .A2(pi0644), .ZN(new_n17964_));
  NOR2_X1    g15528(.A1(new_n17611_), .A2(new_n17843_), .ZN(new_n17965_));
  AOI21_X1   g15529(.A1(new_n17867_), .A2(new_n17611_), .B(new_n17965_), .ZN(new_n17966_));
  OAI21_X1   g15530(.A1(new_n17966_), .A2(pi0644), .B(new_n17964_), .ZN(new_n17967_));
  NAND2_X1   g15531(.A1(new_n17967_), .A2(pi0715), .ZN(new_n17968_));
  OAI21_X1   g15532(.A1(new_n17963_), .A2(pi0715), .B(new_n17968_), .ZN(new_n17969_));
  NAND2_X1   g15533(.A1(new_n17958_), .A2(pi0644), .ZN(new_n17970_));
  NAND2_X1   g15534(.A1(new_n17961_), .A2(new_n12975_), .ZN(new_n17971_));
  AOI21_X1   g15535(.A1(new_n17970_), .A2(new_n17971_), .B(new_n12740_), .ZN(new_n17972_));
  OAI21_X1   g15536(.A1(new_n17865_), .A2(pi0644), .B(new_n12740_), .ZN(new_n17973_));
  AND2_X2    g15537(.A1(new_n17966_), .A2(pi0644), .Z(new_n17974_));
  OAI21_X1   g15538(.A1(new_n17974_), .A2(new_n17973_), .B(pi1160), .ZN(new_n17975_));
  OAI22_X1   g15539(.A1(new_n17969_), .A2(pi1160), .B1(new_n17972_), .B2(new_n17975_), .ZN(new_n17976_));
  OAI21_X1   g15540(.A1(new_n17958_), .A2(pi0790), .B(pi0832), .ZN(new_n17977_));
  AOI21_X1   g15541(.A1(new_n17976_), .A2(pi0790), .B(new_n17977_), .ZN(new_n17978_));
  NOR2_X1    g15542(.A1(new_n13193_), .A2(pi0175), .ZN(new_n17979_));
  AOI21_X1   g15543(.A1(new_n17979_), .A2(pi0644), .B(new_n12740_), .ZN(new_n17980_));
  NOR2_X1    g15544(.A1(new_n17979_), .A2(new_n12985_), .ZN(new_n17981_));
  INV_X1     g15545(.I(new_n17979_), .ZN(new_n17982_));
  NAND2_X1   g15546(.A1(new_n17982_), .A2(new_n12943_), .ZN(new_n17983_));
  NOR2_X1    g15547(.A1(new_n2609_), .A2(new_n9541_), .ZN(new_n17984_));
  OAI22_X1   g15548(.A1(new_n16380_), .A2(pi0175), .B1(new_n16384_), .B2(new_n13208_), .ZN(new_n17985_));
  INV_X1     g15549(.I(new_n13334_), .ZN(new_n17986_));
  NAND3_X1   g15550(.A1(new_n17986_), .A2(new_n9541_), .A3(pi0766), .ZN(new_n17987_));
  NAND2_X1   g15551(.A1(new_n17987_), .A2(new_n17985_), .ZN(new_n17988_));
  OAI22_X1   g15552(.A1(new_n14065_), .A2(pi0766), .B1(new_n9541_), .B2(new_n14067_), .ZN(new_n17989_));
  AOI21_X1   g15553(.A1(pi0039), .A2(new_n17989_), .B(new_n17988_), .ZN(new_n17990_));
  NAND2_X1   g15554(.A1(new_n13397_), .A2(new_n9541_), .ZN(new_n17991_));
  NAND2_X1   g15555(.A1(new_n17991_), .A2(pi0038), .ZN(new_n17992_));
  NOR2_X1    g15556(.A1(new_n13342_), .A2(new_n16384_), .ZN(new_n17993_));
  OAI22_X1   g15557(.A1(new_n17990_), .A2(pi0038), .B1(new_n17992_), .B2(new_n17993_), .ZN(new_n17994_));
  AOI21_X1   g15558(.A1(new_n17994_), .A2(new_n2609_), .B(new_n17984_), .ZN(new_n17995_));
  NOR2_X1    g15559(.A1(new_n17995_), .A2(new_n12760_), .ZN(new_n17996_));
  NOR2_X1    g15560(.A1(new_n17979_), .A2(new_n12761_), .ZN(new_n17997_));
  NOR3_X1    g15561(.A1(new_n17996_), .A2(pi0785), .A3(new_n17997_), .ZN(new_n17998_));
  AOI22_X1   g15562(.A1(new_n17996_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n17982_), .ZN(new_n17999_));
  NOR2_X1    g15563(.A1(new_n17999_), .A2(pi1155), .ZN(new_n18000_));
  AOI22_X1   g15564(.A1(new_n17996_), .A2(pi0609), .B1(new_n13357_), .B2(new_n17982_), .ZN(new_n18001_));
  NOR2_X1    g15565(.A1(new_n18001_), .A2(new_n12770_), .ZN(new_n18002_));
  NOR3_X1    g15566(.A1(new_n18002_), .A2(new_n18000_), .A3(new_n12764_), .ZN(new_n18003_));
  NOR2_X1    g15567(.A1(new_n18003_), .A2(new_n17998_), .ZN(new_n18004_));
  NAND2_X1   g15568(.A1(new_n18004_), .A2(new_n12781_), .ZN(new_n18005_));
  NOR2_X1    g15569(.A1(new_n17979_), .A2(new_n12781_), .ZN(new_n18006_));
  INV_X1     g15570(.I(new_n18006_), .ZN(new_n18007_));
  AOI21_X1   g15571(.A1(new_n18005_), .A2(new_n18007_), .B(pi1154), .ZN(new_n18008_));
  NAND2_X1   g15572(.A1(new_n18004_), .A2(pi0618), .ZN(new_n18009_));
  NAND2_X1   g15573(.A1(new_n17982_), .A2(new_n12781_), .ZN(new_n18010_));
  AOI21_X1   g15574(.A1(new_n18009_), .A2(new_n18010_), .B(new_n12785_), .ZN(new_n18011_));
  OR2_X2     g15575(.A1(new_n18011_), .A2(new_n12779_), .Z(new_n18012_));
  OAI22_X1   g15576(.A1(new_n18012_), .A2(new_n18008_), .B1(pi0781), .B2(new_n18004_), .ZN(new_n18013_));
  NAND2_X1   g15577(.A1(new_n17982_), .A2(pi0619), .ZN(new_n18014_));
  OAI21_X1   g15578(.A1(new_n18013_), .A2(pi0619), .B(new_n18014_), .ZN(new_n18015_));
  NAND2_X1   g15579(.A1(new_n18015_), .A2(new_n12791_), .ZN(new_n18016_));
  NOR2_X1    g15580(.A1(new_n18013_), .A2(new_n12793_), .ZN(new_n18017_));
  AOI21_X1   g15581(.A1(new_n12793_), .A2(new_n17982_), .B(new_n18017_), .ZN(new_n18018_));
  NOR2_X1    g15582(.A1(new_n18018_), .A2(new_n12791_), .ZN(new_n18019_));
  NOR2_X1    g15583(.A1(new_n18019_), .A2(new_n12796_), .ZN(new_n18020_));
  AOI22_X1   g15584(.A1(new_n18020_), .A2(new_n18016_), .B1(new_n12796_), .B2(new_n18013_), .ZN(new_n18021_));
  NOR2_X1    g15585(.A1(new_n17979_), .A2(new_n17504_), .ZN(new_n18022_));
  AOI21_X1   g15586(.A1(new_n18021_), .A2(new_n17504_), .B(new_n18022_), .ZN(new_n18023_));
  OAI21_X1   g15587(.A1(new_n18023_), .A2(new_n12943_), .B(new_n17983_), .ZN(new_n18024_));
  AOI21_X1   g15588(.A1(new_n18024_), .A2(new_n12985_), .B(new_n17981_), .ZN(new_n18025_));
  NAND2_X1   g15589(.A1(new_n18025_), .A2(new_n12975_), .ZN(new_n18026_));
  AOI21_X1   g15590(.A1(new_n18026_), .A2(new_n17980_), .B(pi1160), .ZN(new_n18027_));
  NAND2_X1   g15591(.A1(new_n17982_), .A2(new_n12741_), .ZN(new_n18028_));
  NOR2_X1    g15592(.A1(new_n17979_), .A2(pi0628), .ZN(new_n18029_));
  NAND2_X1   g15593(.A1(new_n17979_), .A2(new_n12869_), .ZN(new_n18030_));
  INV_X1     g15594(.I(new_n17984_), .ZN(new_n18031_));
  NAND3_X1   g15595(.A1(new_n13395_), .A2(new_n9541_), .A3(new_n17869_), .ZN(new_n18032_));
  INV_X1     g15596(.I(new_n14122_), .ZN(new_n18033_));
  NOR2_X1    g15597(.A1(new_n18033_), .A2(new_n9541_), .ZN(new_n18034_));
  AOI21_X1   g15598(.A1(new_n9541_), .A2(new_n14118_), .B(new_n18034_), .ZN(new_n18035_));
  AOI21_X1   g15599(.A1(new_n13399_), .A2(new_n17991_), .B(new_n17869_), .ZN(new_n18036_));
  OAI21_X1   g15600(.A1(new_n18035_), .A2(pi0038), .B(new_n18036_), .ZN(new_n18037_));
  NAND3_X1   g15601(.A1(new_n18037_), .A2(new_n2609_), .A3(new_n18032_), .ZN(new_n18038_));
  NAND2_X1   g15602(.A1(new_n18038_), .A2(new_n18031_), .ZN(new_n18039_));
  NAND2_X1   g15603(.A1(new_n17982_), .A2(pi0625), .ZN(new_n18040_));
  NAND2_X1   g15604(.A1(new_n18039_), .A2(new_n13521_), .ZN(new_n18041_));
  AOI21_X1   g15605(.A1(new_n18041_), .A2(new_n18040_), .B(pi1153), .ZN(new_n18042_));
  NAND2_X1   g15606(.A1(new_n17982_), .A2(new_n13521_), .ZN(new_n18043_));
  NAND2_X1   g15607(.A1(new_n18039_), .A2(pi0625), .ZN(new_n18044_));
  AOI21_X1   g15608(.A1(new_n18044_), .A2(new_n18043_), .B(new_n12841_), .ZN(new_n18045_));
  OR2_X2     g15609(.A1(new_n18045_), .A2(new_n12758_), .Z(new_n18046_));
  OAI22_X1   g15610(.A1(new_n18046_), .A2(new_n18042_), .B1(pi0778), .B2(new_n18039_), .ZN(new_n18047_));
  NAND2_X1   g15611(.A1(new_n18047_), .A2(new_n12870_), .ZN(new_n18048_));
  NAND2_X1   g15612(.A1(new_n18048_), .A2(new_n18030_), .ZN(new_n18049_));
  NAND2_X1   g15613(.A1(new_n17982_), .A2(new_n12887_), .ZN(new_n18050_));
  OAI21_X1   g15614(.A1(new_n18049_), .A2(new_n12887_), .B(new_n18050_), .ZN(new_n18051_));
  NAND2_X1   g15615(.A1(new_n17979_), .A2(new_n12910_), .ZN(new_n18052_));
  OAI21_X1   g15616(.A1(new_n18051_), .A2(new_n12910_), .B(new_n18052_), .ZN(new_n18053_));
  NAND2_X1   g15617(.A1(new_n17982_), .A2(new_n12817_), .ZN(new_n18054_));
  OAI21_X1   g15618(.A1(new_n18053_), .A2(new_n12817_), .B(new_n18054_), .ZN(new_n18055_));
  AOI21_X1   g15619(.A1(new_n18055_), .A2(pi0628), .B(new_n18029_), .ZN(new_n18056_));
  NOR2_X1    g15620(.A1(new_n18056_), .A2(new_n12742_), .ZN(new_n18057_));
  NOR2_X1    g15621(.A1(new_n17979_), .A2(new_n12920_), .ZN(new_n18058_));
  AOI21_X1   g15622(.A1(new_n18055_), .A2(new_n12920_), .B(new_n18058_), .ZN(new_n18059_));
  NOR2_X1    g15623(.A1(new_n18059_), .A2(pi1156), .ZN(new_n18060_));
  OAI21_X1   g15624(.A1(new_n18057_), .A2(new_n18060_), .B(pi0792), .ZN(new_n18061_));
  NAND2_X1   g15625(.A1(new_n18055_), .A2(new_n12937_), .ZN(new_n18062_));
  NAND2_X1   g15626(.A1(new_n18061_), .A2(new_n18062_), .ZN(new_n18063_));
  NAND2_X1   g15627(.A1(new_n18063_), .A2(pi0647), .ZN(new_n18064_));
  AOI21_X1   g15628(.A1(new_n18064_), .A2(new_n18028_), .B(new_n12965_), .ZN(new_n18065_));
  NAND2_X1   g15629(.A1(new_n17982_), .A2(pi0647), .ZN(new_n18066_));
  NAND2_X1   g15630(.A1(new_n18063_), .A2(new_n12741_), .ZN(new_n18067_));
  AOI21_X1   g15631(.A1(new_n18067_), .A2(new_n18066_), .B(pi1157), .ZN(new_n18068_));
  OAI21_X1   g15632(.A1(new_n18065_), .A2(new_n18068_), .B(pi0787), .ZN(new_n18069_));
  NAND2_X1   g15633(.A1(new_n18063_), .A2(new_n12972_), .ZN(new_n18070_));
  NAND2_X1   g15634(.A1(new_n18069_), .A2(new_n18070_), .ZN(new_n18071_));
  OAI21_X1   g15635(.A1(new_n18071_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n18072_));
  AOI21_X1   g15636(.A1(new_n17979_), .A2(new_n12975_), .B(pi0715), .ZN(new_n18073_));
  NAND2_X1   g15637(.A1(new_n18025_), .A2(pi0644), .ZN(new_n18074_));
  AOI21_X1   g15638(.A1(new_n18074_), .A2(new_n18073_), .B(new_n12739_), .ZN(new_n18075_));
  OAI21_X1   g15639(.A1(new_n18071_), .A2(pi0644), .B(pi0715), .ZN(new_n18076_));
  AOI22_X1   g15640(.A1(new_n18027_), .A2(new_n18072_), .B1(new_n18075_), .B2(new_n18076_), .ZN(new_n18077_));
  NOR2_X1    g15641(.A1(new_n18077_), .A2(new_n13000_), .ZN(new_n18078_));
  OR2_X2     g15642(.A1(new_n18075_), .A2(new_n12975_), .Z(new_n18079_));
  OR2_X2     g15643(.A1(new_n18027_), .A2(pi0644), .Z(new_n18080_));
  AOI21_X1   g15644(.A1(new_n18079_), .A2(new_n18080_), .B(new_n13000_), .ZN(new_n18081_));
  NAND2_X1   g15645(.A1(new_n18064_), .A2(new_n18028_), .ZN(new_n18082_));
  NAND2_X1   g15646(.A1(new_n18067_), .A2(new_n18066_), .ZN(new_n18083_));
  AOI22_X1   g15647(.A1(new_n12980_), .A2(new_n18082_), .B1(new_n18083_), .B2(new_n12982_), .ZN(new_n18084_));
  NAND2_X1   g15648(.A1(new_n18024_), .A2(new_n15608_), .ZN(new_n18085_));
  AOI21_X1   g15649(.A1(new_n18085_), .A2(new_n18084_), .B(new_n12972_), .ZN(new_n18086_));
  INV_X1     g15650(.I(new_n12940_), .ZN(new_n18087_));
  INV_X1     g15651(.I(new_n12941_), .ZN(new_n18088_));
  OAI22_X1   g15652(.A1(new_n18087_), .A2(new_n18056_), .B1(new_n18059_), .B2(new_n18088_), .ZN(new_n18089_));
  NOR2_X1    g15653(.A1(new_n18023_), .A2(new_n15821_), .ZN(new_n18090_));
  OAI21_X1   g15654(.A1(new_n18090_), .A2(new_n18089_), .B(pi0792), .ZN(new_n18091_));
  NOR2_X1    g15655(.A1(new_n18021_), .A2(pi0626), .ZN(new_n18092_));
  AOI21_X1   g15656(.A1(pi0626), .A2(new_n17979_), .B(new_n18092_), .ZN(new_n18093_));
  NAND2_X1   g15657(.A1(new_n17979_), .A2(new_n12747_), .ZN(new_n18094_));
  OAI21_X1   g15658(.A1(new_n18021_), .A2(new_n12747_), .B(new_n18094_), .ZN(new_n18095_));
  AOI22_X1   g15659(.A1(new_n18095_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n18053_), .ZN(new_n18096_));
  OAI21_X1   g15660(.A1(new_n12816_), .A2(new_n18093_), .B(new_n18096_), .ZN(new_n18097_));
  AOI21_X1   g15661(.A1(new_n18097_), .A2(pi0788), .B(new_n15340_), .ZN(new_n18098_));
  OR2_X2     g15662(.A1(new_n18047_), .A2(pi0609), .Z(new_n18099_));
  OAI21_X1   g15663(.A1(new_n13562_), .A2(new_n17844_), .B(pi0175), .ZN(new_n18100_));
  NOR2_X1    g15664(.A1(new_n13568_), .A2(new_n13569_), .ZN(new_n18101_));
  INV_X1     g15665(.I(new_n18101_), .ZN(new_n18102_));
  OAI21_X1   g15666(.A1(new_n18102_), .A2(pi0766), .B(new_n13566_), .ZN(new_n18103_));
  NAND2_X1   g15667(.A1(new_n18103_), .A2(new_n2627_), .ZN(new_n18104_));
  AOI21_X1   g15668(.A1(new_n18104_), .A2(new_n9541_), .B(new_n3265_), .ZN(new_n18105_));
  OAI21_X1   g15669(.A1(new_n5337_), .A2(new_n18100_), .B(new_n18105_), .ZN(new_n18106_));
  NOR2_X1    g15670(.A1(new_n14172_), .A2(new_n9541_), .ZN(new_n18107_));
  NOR2_X1    g15671(.A1(new_n14174_), .A2(pi0175), .ZN(new_n18108_));
  OAI21_X1   g15672(.A1(new_n18107_), .A2(new_n18108_), .B(pi0766), .ZN(new_n18109_));
  OAI21_X1   g15673(.A1(new_n12821_), .A2(new_n13798_), .B(new_n13405_), .ZN(new_n18110_));
  NAND2_X1   g15674(.A1(new_n18110_), .A2(new_n9541_), .ZN(new_n18111_));
  OAI21_X1   g15675(.A1(new_n9541_), .A2(new_n15835_), .B(new_n18111_), .ZN(new_n18112_));
  NAND2_X1   g15676(.A1(new_n18112_), .A2(new_n16384_), .ZN(new_n18113_));
  NAND3_X1   g15677(.A1(new_n18113_), .A2(new_n2627_), .A3(new_n18109_), .ZN(new_n18114_));
  NOR2_X1    g15678(.A1(new_n14182_), .A2(pi0175), .ZN(new_n18115_));
  NOR2_X1    g15679(.A1(new_n14184_), .A2(new_n9541_), .ZN(new_n18116_));
  OAI21_X1   g15680(.A1(new_n18115_), .A2(new_n18116_), .B(new_n16384_), .ZN(new_n18117_));
  NOR2_X1    g15681(.A1(new_n14187_), .A2(new_n9541_), .ZN(new_n18118_));
  NOR2_X1    g15682(.A1(new_n14189_), .A2(pi0175), .ZN(new_n18119_));
  OAI21_X1   g15683(.A1(new_n18118_), .A2(new_n18119_), .B(pi0766), .ZN(new_n18120_));
  NAND3_X1   g15684(.A1(new_n18120_), .A2(new_n18117_), .A3(pi0039), .ZN(new_n18121_));
  NAND3_X1   g15685(.A1(new_n18114_), .A2(new_n18121_), .A3(new_n3265_), .ZN(new_n18122_));
  NAND3_X1   g15686(.A1(new_n18122_), .A2(pi0700), .A3(new_n18106_), .ZN(new_n18123_));
  NAND2_X1   g15687(.A1(new_n18123_), .A2(new_n2609_), .ZN(new_n18124_));
  NOR2_X1    g15688(.A1(new_n17994_), .A2(pi0700), .ZN(new_n18125_));
  OAI21_X1   g15689(.A1(new_n18124_), .A2(new_n18125_), .B(new_n18031_), .ZN(new_n18126_));
  OR2_X2     g15690(.A1(new_n17995_), .A2(new_n13521_), .Z(new_n18127_));
  NAND2_X1   g15691(.A1(new_n18126_), .A2(new_n13521_), .ZN(new_n18128_));
  AOI21_X1   g15692(.A1(new_n18128_), .A2(new_n18127_), .B(pi1153), .ZN(new_n18129_));
  NOR3_X1    g15693(.A1(new_n18129_), .A2(pi0608), .A3(new_n18045_), .ZN(new_n18130_));
  NOR2_X1    g15694(.A1(new_n17995_), .A2(pi0625), .ZN(new_n18131_));
  AOI21_X1   g15695(.A1(new_n18126_), .A2(pi0625), .B(new_n18131_), .ZN(new_n18132_));
  NOR2_X1    g15696(.A1(new_n18132_), .A2(new_n12841_), .ZN(new_n18133_));
  NOR3_X1    g15697(.A1(new_n18133_), .A2(new_n13560_), .A3(new_n18042_), .ZN(new_n18134_));
  NOR3_X1    g15698(.A1(new_n18134_), .A2(new_n18130_), .A3(new_n12758_), .ZN(new_n18135_));
  AOI21_X1   g15699(.A1(new_n12758_), .A2(new_n18126_), .B(new_n18135_), .ZN(new_n18136_));
  OAI21_X1   g15700(.A1(new_n18136_), .A2(new_n12766_), .B(new_n18099_), .ZN(new_n18137_));
  AOI21_X1   g15701(.A1(new_n18137_), .A2(pi1155), .B(new_n18000_), .ZN(new_n18138_));
  NOR2_X1    g15702(.A1(new_n18136_), .A2(pi0609), .ZN(new_n18139_));
  NOR2_X1    g15703(.A1(new_n18047_), .A2(new_n12766_), .ZN(new_n18140_));
  OAI21_X1   g15704(.A1(new_n18139_), .A2(new_n18140_), .B(new_n12770_), .ZN(new_n18141_));
  NOR2_X1    g15705(.A1(new_n18002_), .A2(pi0660), .ZN(new_n18142_));
  AOI22_X1   g15706(.A1(new_n18138_), .A2(pi0660), .B1(new_n18141_), .B2(new_n18142_), .ZN(new_n18143_));
  AND2_X2    g15707(.A1(new_n18143_), .A2(pi0785), .Z(new_n18144_));
  NOR2_X1    g15708(.A1(new_n18136_), .A2(pi0785), .ZN(new_n18145_));
  NOR2_X1    g15709(.A1(new_n18144_), .A2(new_n18145_), .ZN(new_n18146_));
  NOR2_X1    g15710(.A1(new_n18146_), .A2(pi0781), .ZN(new_n18147_));
  NOR2_X1    g15711(.A1(new_n18049_), .A2(pi0618), .ZN(new_n18148_));
  INV_X1     g15712(.I(new_n18148_), .ZN(new_n18149_));
  OAI21_X1   g15713(.A1(new_n18144_), .A2(new_n18145_), .B(pi0618), .ZN(new_n18150_));
  AOI21_X1   g15714(.A1(new_n18150_), .A2(new_n18149_), .B(new_n12785_), .ZN(new_n18151_));
  NOR3_X1    g15715(.A1(new_n18151_), .A2(new_n12880_), .A3(new_n18008_), .ZN(new_n18152_));
  OAI21_X1   g15716(.A1(new_n18144_), .A2(new_n18145_), .B(new_n12781_), .ZN(new_n18153_));
  NAND3_X1   g15717(.A1(new_n18048_), .A2(pi0618), .A3(new_n18030_), .ZN(new_n18154_));
  AOI21_X1   g15718(.A1(new_n18153_), .A2(new_n18154_), .B(pi1154), .ZN(new_n18155_));
  NOR3_X1    g15719(.A1(new_n18155_), .A2(pi0627), .A3(new_n18011_), .ZN(new_n18156_));
  NOR3_X1    g15720(.A1(new_n18152_), .A2(new_n18156_), .A3(new_n12779_), .ZN(new_n18157_));
  OAI21_X1   g15721(.A1(new_n18157_), .A2(new_n18147_), .B(new_n12796_), .ZN(new_n18158_));
  NAND2_X1   g15722(.A1(new_n18158_), .A2(new_n12819_), .ZN(new_n18159_));
  NAND2_X1   g15723(.A1(new_n18051_), .A2(pi0619), .ZN(new_n18160_));
  OAI21_X1   g15724(.A1(new_n18157_), .A2(new_n18147_), .B(new_n12793_), .ZN(new_n18161_));
  AOI21_X1   g15725(.A1(new_n18161_), .A2(new_n18160_), .B(pi1159), .ZN(new_n18162_));
  NOR3_X1    g15726(.A1(new_n18162_), .A2(pi0648), .A3(new_n18019_), .ZN(new_n18163_));
  INV_X1     g15727(.I(new_n18016_), .ZN(new_n18164_));
  OAI21_X1   g15728(.A1(new_n18157_), .A2(new_n18147_), .B(pi0619), .ZN(new_n18165_));
  NAND2_X1   g15729(.A1(new_n18051_), .A2(new_n12793_), .ZN(new_n18166_));
  AOI21_X1   g15730(.A1(new_n18165_), .A2(new_n18166_), .B(new_n12791_), .ZN(new_n18167_));
  NOR3_X1    g15731(.A1(new_n18167_), .A2(new_n12895_), .A3(new_n18164_), .ZN(new_n18168_));
  NOR3_X1    g15732(.A1(new_n18163_), .A2(new_n18168_), .A3(new_n12796_), .ZN(new_n18169_));
  OAI21_X1   g15733(.A1(new_n18169_), .A2(new_n18159_), .B(new_n18098_), .ZN(new_n18170_));
  AOI21_X1   g15734(.A1(new_n18170_), .A2(new_n18091_), .B(new_n15341_), .ZN(new_n18171_));
  NOR3_X1    g15735(.A1(new_n18081_), .A2(new_n18086_), .A3(new_n18171_), .ZN(new_n18172_));
  OAI21_X1   g15736(.A1(new_n18172_), .A2(new_n18078_), .B(new_n6643_), .ZN(new_n18173_));
  AOI21_X1   g15737(.A1(po1038), .A2(new_n9541_), .B(pi0832), .ZN(new_n18174_));
  AOI21_X1   g15738(.A1(new_n18173_), .A2(new_n18174_), .B(new_n17978_), .ZN(po0332));
  NOR2_X1    g15739(.A1(new_n3042_), .A2(pi0176), .ZN(new_n18176_));
  INV_X1     g15740(.I(new_n18176_), .ZN(new_n18177_));
  AOI21_X1   g15741(.A1(new_n12756_), .A2(new_n16430_), .B(new_n18176_), .ZN(new_n18178_));
  NOR3_X1    g15742(.A1(new_n18178_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n18179_));
  NOR2_X1    g15743(.A1(new_n18178_), .A2(new_n12762_), .ZN(new_n18180_));
  AOI21_X1   g15744(.A1(new_n18180_), .A2(new_n12768_), .B(pi1155), .ZN(new_n18181_));
  INV_X1     g15745(.I(new_n18178_), .ZN(new_n18182_));
  AOI21_X1   g15746(.A1(new_n18182_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n18183_));
  NOR3_X1    g15747(.A1(new_n18181_), .A2(new_n18183_), .A3(new_n12764_), .ZN(new_n18184_));
  NOR2_X1    g15748(.A1(new_n18184_), .A2(new_n18179_), .ZN(new_n18185_));
  NOR2_X1    g15749(.A1(new_n18185_), .A2(pi0781), .ZN(new_n18186_));
  INV_X1     g15750(.I(new_n18185_), .ZN(new_n18187_));
  AOI21_X1   g15751(.A1(new_n18187_), .A2(new_n12783_), .B(pi1154), .ZN(new_n18188_));
  AOI21_X1   g15752(.A1(new_n18187_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n18189_));
  NOR3_X1    g15753(.A1(new_n18188_), .A2(new_n18189_), .A3(new_n12779_), .ZN(new_n18190_));
  NOR2_X1    g15754(.A1(new_n18190_), .A2(new_n18186_), .ZN(new_n18191_));
  NOR3_X1    g15755(.A1(new_n18190_), .A2(pi0619), .A3(new_n18186_), .ZN(new_n18192_));
  NOR2_X1    g15756(.A1(new_n18176_), .A2(new_n12793_), .ZN(new_n18193_));
  OAI21_X1   g15757(.A1(new_n18192_), .A2(new_n18193_), .B(new_n12791_), .ZN(new_n18194_));
  NAND2_X1   g15758(.A1(new_n18191_), .A2(pi0619), .ZN(new_n18195_));
  NAND2_X1   g15759(.A1(new_n18177_), .A2(new_n12793_), .ZN(new_n18196_));
  AOI21_X1   g15760(.A1(new_n18195_), .A2(new_n18196_), .B(new_n12791_), .ZN(new_n18197_));
  INV_X1     g15761(.I(new_n18197_), .ZN(new_n18198_));
  NAND3_X1   g15762(.A1(new_n18198_), .A2(pi0789), .A3(new_n18194_), .ZN(new_n18199_));
  OAI21_X1   g15763(.A1(pi0789), .A2(new_n18191_), .B(new_n18199_), .ZN(new_n18200_));
  NOR2_X1    g15764(.A1(new_n18200_), .A2(new_n12818_), .ZN(new_n18201_));
  AOI21_X1   g15765(.A1(new_n12818_), .A2(new_n18177_), .B(new_n18201_), .ZN(new_n18202_));
  INV_X1     g15766(.I(new_n12912_), .ZN(new_n18203_));
  AOI21_X1   g15767(.A1(new_n12826_), .A2(new_n16429_), .B(new_n18176_), .ZN(new_n18204_));
  NOR2_X1    g15768(.A1(new_n18204_), .A2(pi0778), .ZN(new_n18205_));
  NOR2_X1    g15769(.A1(new_n18176_), .A2(pi1153), .ZN(new_n18206_));
  NOR2_X1    g15770(.A1(new_n12834_), .A2(pi0704), .ZN(new_n18207_));
  INV_X1     g15771(.I(new_n18207_), .ZN(new_n18208_));
  NAND2_X1   g15772(.A1(new_n18208_), .A2(new_n18206_), .ZN(new_n18209_));
  INV_X1     g15773(.I(new_n18209_), .ZN(new_n18210_));
  NOR2_X1    g15774(.A1(new_n18207_), .A2(new_n18204_), .ZN(new_n18211_));
  NOR2_X1    g15775(.A1(new_n18211_), .A2(new_n12841_), .ZN(new_n18212_));
  NOR2_X1    g15776(.A1(new_n18210_), .A2(new_n18212_), .ZN(new_n18213_));
  AOI21_X1   g15777(.A1(new_n18213_), .A2(pi0778), .B(new_n18205_), .ZN(new_n18214_));
  NOR2_X1    g15778(.A1(new_n18214_), .A2(new_n12871_), .ZN(new_n18215_));
  INV_X1     g15779(.I(new_n18215_), .ZN(new_n18216_));
  NOR2_X1    g15780(.A1(new_n18216_), .A2(new_n12889_), .ZN(new_n18217_));
  NAND2_X1   g15781(.A1(new_n18217_), .A2(new_n18203_), .ZN(new_n18218_));
  NOR2_X1    g15782(.A1(new_n18218_), .A2(new_n17884_), .ZN(new_n18219_));
  AOI22_X1   g15783(.A1(new_n18202_), .A2(new_n12949_), .B1(new_n15695_), .B2(new_n18219_), .ZN(new_n18220_));
  NOR2_X1    g15784(.A1(new_n18220_), .A2(pi0629), .ZN(new_n18221_));
  AOI22_X1   g15785(.A1(new_n18202_), .A2(new_n12948_), .B1(new_n15700_), .B2(new_n18219_), .ZN(new_n18222_));
  NOR2_X1    g15786(.A1(new_n18222_), .A2(new_n12919_), .ZN(new_n18223_));
  NOR2_X1    g15787(.A1(new_n18221_), .A2(new_n18223_), .ZN(new_n18224_));
  NOR2_X1    g15788(.A1(new_n18204_), .A2(new_n12754_), .ZN(new_n18225_));
  NOR2_X1    g15789(.A1(new_n18225_), .A2(new_n18182_), .ZN(new_n18226_));
  NAND2_X1   g15790(.A1(new_n18226_), .A2(new_n12758_), .ZN(new_n18227_));
  NAND2_X1   g15791(.A1(new_n18225_), .A2(pi0625), .ZN(new_n18228_));
  NAND3_X1   g15792(.A1(new_n18228_), .A2(pi1153), .A3(new_n18178_), .ZN(new_n18229_));
  AND3_X2    g15793(.A1(new_n18209_), .A2(pi0608), .A3(new_n18229_), .Z(new_n18230_));
  NOR2_X1    g15794(.A1(new_n18212_), .A2(pi0608), .ZN(new_n18231_));
  INV_X1     g15795(.I(new_n18228_), .ZN(new_n18232_));
  OAI21_X1   g15796(.A1(new_n18232_), .A2(new_n18226_), .B(new_n18206_), .ZN(new_n18233_));
  NAND2_X1   g15797(.A1(new_n18231_), .A2(new_n18233_), .ZN(new_n18234_));
  NAND2_X1   g15798(.A1(new_n18234_), .A2(pi0778), .ZN(new_n18235_));
  OAI21_X1   g15799(.A1(new_n18235_), .A2(new_n18230_), .B(new_n18227_), .ZN(new_n18236_));
  INV_X1     g15800(.I(new_n18236_), .ZN(new_n18237_));
  NAND2_X1   g15801(.A1(new_n18214_), .A2(new_n12766_), .ZN(new_n18238_));
  OAI21_X1   g15802(.A1(new_n18237_), .A2(new_n12766_), .B(new_n18238_), .ZN(new_n18239_));
  AOI21_X1   g15803(.A1(new_n18239_), .A2(pi1155), .B(new_n18181_), .ZN(new_n18240_));
  NAND2_X1   g15804(.A1(new_n18236_), .A2(new_n12766_), .ZN(new_n18241_));
  NAND2_X1   g15805(.A1(new_n18214_), .A2(pi0609), .ZN(new_n18242_));
  AOI21_X1   g15806(.A1(new_n18241_), .A2(new_n18242_), .B(pi1155), .ZN(new_n18243_));
  NOR3_X1    g15807(.A1(new_n18243_), .A2(pi0660), .A3(new_n18183_), .ZN(new_n18244_));
  AOI21_X1   g15808(.A1(pi0660), .A2(new_n18240_), .B(new_n18244_), .ZN(new_n18245_));
  NAND2_X1   g15809(.A1(new_n18245_), .A2(pi0785), .ZN(new_n18246_));
  OAI21_X1   g15810(.A1(pi0785), .A2(new_n18237_), .B(new_n18246_), .ZN(new_n18247_));
  INV_X1     g15811(.I(new_n18247_), .ZN(new_n18248_));
  NAND2_X1   g15812(.A1(new_n18216_), .A2(pi0618), .ZN(new_n18249_));
  OAI21_X1   g15813(.A1(new_n18248_), .A2(pi0618), .B(new_n18249_), .ZN(new_n18250_));
  AOI21_X1   g15814(.A1(new_n18250_), .A2(new_n12785_), .B(new_n18189_), .ZN(new_n18251_));
  NOR2_X1    g15815(.A1(new_n18215_), .A2(pi0618), .ZN(new_n18252_));
  NOR2_X1    g15816(.A1(new_n18248_), .A2(new_n12781_), .ZN(new_n18253_));
  OAI21_X1   g15817(.A1(new_n18253_), .A2(new_n18252_), .B(pi1154), .ZN(new_n18254_));
  NOR2_X1    g15818(.A1(new_n18188_), .A2(new_n12880_), .ZN(new_n18255_));
  AOI22_X1   g15819(.A1(new_n18251_), .A2(new_n12880_), .B1(new_n18254_), .B2(new_n18255_), .ZN(new_n18256_));
  NAND2_X1   g15820(.A1(new_n18256_), .A2(pi0781), .ZN(new_n18257_));
  NAND2_X1   g15821(.A1(new_n18247_), .A2(new_n12779_), .ZN(new_n18258_));
  NAND2_X1   g15822(.A1(new_n18257_), .A2(new_n18258_), .ZN(new_n18259_));
  AOI21_X1   g15823(.A1(new_n18259_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n18260_));
  NOR2_X1    g15824(.A1(new_n18217_), .A2(pi0619), .ZN(new_n18261_));
  INV_X1     g15825(.I(new_n18259_), .ZN(new_n18262_));
  NOR2_X1    g15826(.A1(new_n18262_), .A2(new_n12793_), .ZN(new_n18263_));
  OAI21_X1   g15827(.A1(new_n18263_), .A2(new_n18261_), .B(pi1159), .ZN(new_n18264_));
  NAND3_X1   g15828(.A1(new_n18264_), .A2(pi0648), .A3(new_n18194_), .ZN(new_n18265_));
  NOR2_X1    g15829(.A1(new_n18262_), .A2(pi0619), .ZN(new_n18266_));
  NOR2_X1    g15830(.A1(new_n18217_), .A2(new_n12793_), .ZN(new_n18267_));
  OAI21_X1   g15831(.A1(new_n18266_), .A2(new_n18267_), .B(new_n12791_), .ZN(new_n18268_));
  NAND3_X1   g15832(.A1(new_n18268_), .A2(new_n12895_), .A3(new_n18198_), .ZN(new_n18269_));
  NAND3_X1   g15833(.A1(new_n18265_), .A2(new_n18269_), .A3(pi0789), .ZN(new_n18270_));
  NOR2_X1    g15834(.A1(new_n18177_), .A2(new_n12747_), .ZN(new_n18271_));
  INV_X1     g15835(.I(new_n18200_), .ZN(new_n18272_));
  NOR2_X1    g15836(.A1(new_n18272_), .A2(pi0626), .ZN(new_n18273_));
  OAI21_X1   g15837(.A1(new_n18273_), .A2(new_n18271_), .B(new_n12815_), .ZN(new_n18274_));
  INV_X1     g15838(.I(new_n18218_), .ZN(new_n18275_));
  NAND2_X1   g15839(.A1(new_n18176_), .A2(new_n12747_), .ZN(new_n18276_));
  OAI21_X1   g15840(.A1(new_n18272_), .A2(new_n12747_), .B(new_n18276_), .ZN(new_n18277_));
  AOI22_X1   g15841(.A1(new_n18277_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n18275_), .ZN(new_n18278_));
  NAND2_X1   g15842(.A1(new_n18278_), .A2(new_n18274_), .ZN(new_n18279_));
  AOI22_X1   g15843(.A1(new_n18270_), .A2(new_n18260_), .B1(pi0788), .B2(new_n18279_), .ZN(new_n18280_));
  OAI22_X1   g15844(.A1(new_n18280_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n18224_), .ZN(new_n18281_));
  INV_X1     g15845(.I(new_n18202_), .ZN(new_n18282_));
  NAND2_X1   g15846(.A1(new_n18282_), .A2(new_n13384_), .ZN(new_n18283_));
  NAND2_X1   g15847(.A1(new_n12943_), .A2(new_n18177_), .ZN(new_n18284_));
  NAND2_X1   g15848(.A1(new_n18283_), .A2(new_n18284_), .ZN(new_n18285_));
  NAND2_X1   g15849(.A1(new_n18219_), .A2(new_n12954_), .ZN(new_n18286_));
  NAND2_X1   g15850(.A1(new_n18286_), .A2(new_n12741_), .ZN(new_n18287_));
  NOR2_X1    g15851(.A1(new_n18176_), .A2(new_n12741_), .ZN(new_n18288_));
  INV_X1     g15852(.I(new_n18288_), .ZN(new_n18289_));
  AOI21_X1   g15853(.A1(new_n18287_), .A2(new_n18289_), .B(pi1157), .ZN(new_n18290_));
  INV_X1     g15854(.I(new_n18290_), .ZN(new_n18291_));
  NAND2_X1   g15855(.A1(new_n18176_), .A2(new_n12741_), .ZN(new_n18292_));
  OAI21_X1   g15856(.A1(new_n18286_), .A2(new_n12741_), .B(new_n18292_), .ZN(new_n18293_));
  OAI22_X1   g15857(.A1(new_n18291_), .A2(new_n12981_), .B1(new_n18293_), .B2(new_n15576_), .ZN(new_n18294_));
  AOI21_X1   g15858(.A1(new_n18285_), .A2(new_n15608_), .B(new_n18294_), .ZN(new_n18295_));
  OAI22_X1   g15859(.A1(new_n18281_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n18295_), .ZN(new_n18296_));
  NAND2_X1   g15860(.A1(new_n18296_), .A2(new_n13000_), .ZN(new_n18297_));
  AND2_X2    g15861(.A1(new_n18296_), .A2(new_n12975_), .Z(new_n18298_));
  OAI21_X1   g15862(.A1(new_n12965_), .A2(new_n18293_), .B(new_n18291_), .ZN(new_n18299_));
  NAND3_X1   g15863(.A1(new_n18219_), .A2(new_n12972_), .A3(new_n12954_), .ZN(new_n18300_));
  OAI21_X1   g15864(.A1(new_n18299_), .A2(new_n12972_), .B(new_n18300_), .ZN(new_n18301_));
  NOR2_X1    g15865(.A1(new_n18301_), .A2(new_n12975_), .ZN(new_n18302_));
  OAI21_X1   g15866(.A1(new_n18298_), .A2(new_n18302_), .B(new_n12740_), .ZN(new_n18303_));
  NOR2_X1    g15867(.A1(new_n18176_), .A2(new_n12975_), .ZN(new_n18304_));
  NOR2_X1    g15868(.A1(new_n17611_), .A2(new_n18176_), .ZN(new_n18305_));
  AOI21_X1   g15869(.A1(new_n18282_), .A2(new_n17611_), .B(new_n18305_), .ZN(new_n18306_));
  NOR2_X1    g15870(.A1(new_n18306_), .A2(pi0644), .ZN(new_n18307_));
  OAI21_X1   g15871(.A1(new_n18307_), .A2(new_n18304_), .B(pi0715), .ZN(new_n18308_));
  NAND3_X1   g15872(.A1(new_n18303_), .A2(new_n12739_), .A3(new_n18308_), .ZN(new_n18309_));
  NOR2_X1    g15873(.A1(new_n18301_), .A2(pi0644), .ZN(new_n18310_));
  AOI21_X1   g15874(.A1(new_n18296_), .A2(pi0644), .B(new_n18310_), .ZN(new_n18311_));
  NAND2_X1   g15875(.A1(new_n18177_), .A2(new_n12975_), .ZN(new_n18312_));
  OAI21_X1   g15876(.A1(new_n18306_), .A2(new_n12975_), .B(new_n18312_), .ZN(new_n18313_));
  AOI21_X1   g15877(.A1(new_n18313_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n18314_));
  OAI21_X1   g15878(.A1(new_n18311_), .A2(new_n12740_), .B(new_n18314_), .ZN(new_n18315_));
  NAND3_X1   g15879(.A1(new_n18309_), .A2(pi0790), .A3(new_n18315_), .ZN(new_n18316_));
  NAND2_X1   g15880(.A1(new_n18316_), .A2(new_n18297_), .ZN(new_n18317_));
  AOI21_X1   g15881(.A1(po1038), .A2(new_n7518_), .B(pi0832), .ZN(new_n18318_));
  NOR2_X1    g15882(.A1(new_n13193_), .A2(pi0176), .ZN(new_n18319_));
  AOI21_X1   g15883(.A1(new_n18319_), .A2(pi0644), .B(new_n12740_), .ZN(new_n18320_));
  INV_X1     g15884(.I(new_n18319_), .ZN(new_n18321_));
  NAND2_X1   g15885(.A1(new_n18321_), .A2(new_n12984_), .ZN(new_n18322_));
  OAI21_X1   g15886(.A1(new_n15012_), .A2(new_n15011_), .B(new_n7518_), .ZN(new_n18323_));
  OAI21_X1   g15887(.A1(new_n13208_), .A2(new_n13244_), .B(new_n3265_), .ZN(new_n18324_));
  NOR2_X1    g15888(.A1(new_n15006_), .A2(new_n3265_), .ZN(new_n18325_));
  INV_X1     g15889(.I(new_n18325_), .ZN(new_n18326_));
  NAND2_X1   g15890(.A1(new_n18324_), .A2(new_n18326_), .ZN(new_n18327_));
  NOR2_X1    g15891(.A1(new_n18327_), .A2(new_n7518_), .ZN(new_n18328_));
  INV_X1     g15892(.I(new_n18328_), .ZN(new_n18329_));
  AOI21_X1   g15893(.A1(new_n18329_), .A2(new_n18323_), .B(pi0742), .ZN(new_n18330_));
  AOI21_X1   g15894(.A1(new_n7518_), .A2(new_n16447_), .B(new_n18330_), .ZN(new_n18331_));
  NOR2_X1    g15895(.A1(new_n18331_), .A2(new_n2610_), .ZN(new_n18332_));
  AOI21_X1   g15896(.A1(new_n7518_), .A2(new_n2610_), .B(new_n18332_), .ZN(new_n18333_));
  INV_X1     g15897(.I(new_n18333_), .ZN(new_n18334_));
  NOR2_X1    g15898(.A1(new_n18334_), .A2(new_n12760_), .ZN(new_n18335_));
  INV_X1     g15899(.I(new_n18335_), .ZN(new_n18336_));
  OAI21_X1   g15900(.A1(new_n12761_), .A2(new_n18319_), .B(new_n18336_), .ZN(new_n18337_));
  NOR2_X1    g15901(.A1(new_n18319_), .A2(new_n13353_), .ZN(new_n18338_));
  NOR2_X1    g15902(.A1(new_n18336_), .A2(pi0609), .ZN(new_n18339_));
  OAI21_X1   g15903(.A1(new_n18339_), .A2(new_n18338_), .B(new_n12770_), .ZN(new_n18340_));
  INV_X1     g15904(.I(new_n18340_), .ZN(new_n18341_));
  OAI22_X1   g15905(.A1(new_n18336_), .A2(new_n12766_), .B1(new_n12772_), .B2(new_n18319_), .ZN(new_n18342_));
  NAND2_X1   g15906(.A1(new_n18342_), .A2(pi1155), .ZN(new_n18343_));
  NAND2_X1   g15907(.A1(new_n18343_), .A2(pi0785), .ZN(new_n18344_));
  OAI22_X1   g15908(.A1(new_n18344_), .A2(new_n18341_), .B1(pi0785), .B2(new_n18337_), .ZN(new_n18345_));
  NAND2_X1   g15909(.A1(new_n18345_), .A2(new_n12779_), .ZN(new_n18346_));
  NOR2_X1    g15910(.A1(new_n18345_), .A2(pi0618), .ZN(new_n18347_));
  NOR2_X1    g15911(.A1(new_n18319_), .A2(new_n12781_), .ZN(new_n18348_));
  OAI21_X1   g15912(.A1(new_n18347_), .A2(new_n18348_), .B(new_n12785_), .ZN(new_n18349_));
  NOR2_X1    g15913(.A1(new_n18345_), .A2(new_n12781_), .ZN(new_n18350_));
  NOR2_X1    g15914(.A1(new_n18319_), .A2(pi0618), .ZN(new_n18351_));
  OAI21_X1   g15915(.A1(new_n18350_), .A2(new_n18351_), .B(pi1154), .ZN(new_n18352_));
  NAND3_X1   g15916(.A1(new_n18349_), .A2(new_n18352_), .A3(pi0781), .ZN(new_n18353_));
  NAND2_X1   g15917(.A1(new_n18353_), .A2(new_n18346_), .ZN(new_n18354_));
  NOR2_X1    g15918(.A1(new_n18321_), .A2(new_n15807_), .ZN(new_n18355_));
  AOI22_X1   g15919(.A1(new_n18354_), .A2(new_n15779_), .B1(pi0789), .B2(new_n18355_), .ZN(new_n18356_));
  NOR2_X1    g15920(.A1(new_n18319_), .A2(new_n17504_), .ZN(new_n18357_));
  AOI21_X1   g15921(.A1(new_n18356_), .A2(new_n17504_), .B(new_n18357_), .ZN(new_n18358_));
  NOR2_X1    g15922(.A1(new_n18358_), .A2(new_n12943_), .ZN(new_n18359_));
  AOI21_X1   g15923(.A1(new_n12943_), .A2(new_n18321_), .B(new_n18359_), .ZN(new_n18360_));
  OAI21_X1   g15924(.A1(new_n18360_), .A2(new_n12984_), .B(new_n18322_), .ZN(new_n18361_));
  OAI21_X1   g15925(.A1(new_n18361_), .A2(pi0644), .B(new_n18320_), .ZN(new_n18362_));
  AND2_X2    g15926(.A1(new_n18362_), .A2(new_n12739_), .Z(new_n18363_));
  NOR2_X1    g15927(.A1(new_n18319_), .A2(pi0647), .ZN(new_n18364_));
  NOR2_X1    g15928(.A1(new_n18321_), .A2(new_n12870_), .ZN(new_n18365_));
  NOR3_X1    g15929(.A1(new_n13191_), .A2(pi0176), .A3(new_n16429_), .ZN(new_n18366_));
  OAI22_X1   g15930(.A1(new_n15744_), .A2(pi0038), .B1(new_n12824_), .B2(new_n16469_), .ZN(new_n18367_));
  AOI21_X1   g15931(.A1(new_n18367_), .A2(new_n7518_), .B(pi0704), .ZN(new_n18368_));
  NOR3_X1    g15932(.A1(new_n18368_), .A2(new_n2610_), .A3(new_n18366_), .ZN(new_n18369_));
  NAND2_X1   g15933(.A1(new_n14122_), .A2(new_n3265_), .ZN(new_n18370_));
  NAND3_X1   g15934(.A1(new_n18370_), .A2(new_n2609_), .A3(new_n14125_), .ZN(new_n18371_));
  AND2_X2    g15935(.A1(new_n18371_), .A2(pi0176), .Z(new_n18372_));
  NOR2_X1    g15936(.A1(new_n18369_), .A2(new_n18372_), .ZN(new_n18373_));
  INV_X1     g15937(.I(new_n18373_), .ZN(new_n18374_));
  NOR2_X1    g15938(.A1(new_n18373_), .A2(pi0625), .ZN(new_n18375_));
  NOR2_X1    g15939(.A1(new_n18319_), .A2(new_n13521_), .ZN(new_n18376_));
  OAI21_X1   g15940(.A1(new_n18375_), .A2(new_n18376_), .B(new_n12841_), .ZN(new_n18377_));
  NOR2_X1    g15941(.A1(new_n18373_), .A2(new_n13521_), .ZN(new_n18378_));
  NOR2_X1    g15942(.A1(new_n18319_), .A2(pi0625), .ZN(new_n18379_));
  OAI21_X1   g15943(.A1(new_n18378_), .A2(new_n18379_), .B(pi1153), .ZN(new_n18380_));
  NAND3_X1   g15944(.A1(new_n18377_), .A2(new_n18380_), .A3(pi0778), .ZN(new_n18381_));
  OAI21_X1   g15945(.A1(pi0778), .A2(new_n18374_), .B(new_n18381_), .ZN(new_n18382_));
  AOI21_X1   g15946(.A1(new_n18382_), .A2(new_n12870_), .B(new_n18365_), .ZN(new_n18383_));
  NOR2_X1    g15947(.A1(new_n18319_), .A2(new_n12888_), .ZN(new_n18384_));
  AOI21_X1   g15948(.A1(new_n18383_), .A2(new_n12888_), .B(new_n18384_), .ZN(new_n18385_));
  INV_X1     g15949(.I(new_n18385_), .ZN(new_n18386_));
  NOR2_X1    g15950(.A1(new_n18319_), .A2(new_n12923_), .ZN(new_n18387_));
  AOI21_X1   g15951(.A1(new_n18386_), .A2(new_n12923_), .B(new_n18387_), .ZN(new_n18388_));
  XNOR2_X1   g15952(.A1(pi0628), .A2(pi1156), .ZN(new_n18389_));
  NOR2_X1    g15953(.A1(new_n18389_), .A2(new_n12937_), .ZN(new_n18390_));
  OAI21_X1   g15954(.A1(new_n12948_), .A2(new_n12949_), .B(new_n18321_), .ZN(new_n18391_));
  OAI22_X1   g15955(.A1(new_n18388_), .A2(new_n18390_), .B1(new_n12937_), .B2(new_n18391_), .ZN(new_n18392_));
  AOI21_X1   g15956(.A1(new_n18392_), .A2(pi0647), .B(new_n18364_), .ZN(new_n18393_));
  NOR2_X1    g15957(.A1(new_n18393_), .A2(new_n12965_), .ZN(new_n18394_));
  NOR2_X1    g15958(.A1(new_n18319_), .A2(new_n12741_), .ZN(new_n18395_));
  AOI21_X1   g15959(.A1(new_n18392_), .A2(new_n12741_), .B(new_n18395_), .ZN(new_n18396_));
  NOR2_X1    g15960(.A1(new_n18396_), .A2(pi1157), .ZN(new_n18397_));
  OAI21_X1   g15961(.A1(new_n18394_), .A2(new_n18397_), .B(pi0787), .ZN(new_n18398_));
  NAND2_X1   g15962(.A1(new_n18392_), .A2(new_n12972_), .ZN(new_n18399_));
  NAND2_X1   g15963(.A1(new_n18398_), .A2(new_n18399_), .ZN(new_n18400_));
  OAI21_X1   g15964(.A1(new_n18400_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n18401_));
  AOI21_X1   g15965(.A1(new_n18319_), .A2(new_n12975_), .B(pi0715), .ZN(new_n18402_));
  OAI21_X1   g15966(.A1(new_n18361_), .A2(new_n12975_), .B(new_n18402_), .ZN(new_n18403_));
  AND2_X2    g15967(.A1(new_n18403_), .A2(pi1160), .Z(new_n18404_));
  OAI21_X1   g15968(.A1(new_n18400_), .A2(pi0644), .B(pi0715), .ZN(new_n18405_));
  AOI22_X1   g15969(.A1(new_n18363_), .A2(new_n18401_), .B1(new_n18404_), .B2(new_n18405_), .ZN(new_n18406_));
  NOR2_X1    g15970(.A1(new_n18406_), .A2(new_n13000_), .ZN(new_n18407_));
  NAND2_X1   g15971(.A1(new_n18321_), .A2(pi0628), .ZN(new_n18408_));
  OR2_X2     g15972(.A1(new_n18388_), .A2(pi0628), .Z(new_n18409_));
  AOI21_X1   g15973(.A1(new_n18409_), .A2(new_n18408_), .B(new_n18088_), .ZN(new_n18410_));
  NOR2_X1    g15974(.A1(new_n18388_), .A2(new_n12920_), .ZN(new_n18411_));
  AOI21_X1   g15975(.A1(new_n12920_), .A2(new_n18321_), .B(new_n18411_), .ZN(new_n18412_));
  OAI22_X1   g15976(.A1(new_n18358_), .A2(new_n15821_), .B1(new_n18087_), .B2(new_n18412_), .ZN(new_n18413_));
  NOR2_X1    g15977(.A1(new_n18413_), .A2(new_n18410_), .ZN(new_n18414_));
  AOI21_X1   g15978(.A1(new_n18414_), .A2(new_n15340_), .B(new_n15341_), .ZN(new_n18415_));
  OR2_X2     g15979(.A1(new_n18382_), .A2(pi0609), .Z(new_n18416_));
  NOR2_X1    g15980(.A1(new_n18331_), .A2(new_n16429_), .ZN(new_n18417_));
  NAND2_X1   g15981(.A1(new_n15129_), .A2(new_n15126_), .ZN(new_n18418_));
  NOR2_X1    g15982(.A1(new_n18418_), .A2(pi0176), .ZN(new_n18419_));
  INV_X1     g15983(.I(new_n18419_), .ZN(new_n18420_));
  INV_X1     g15984(.I(new_n15123_), .ZN(new_n18421_));
  NAND3_X1   g15985(.A1(new_n15121_), .A2(pi0176), .A3(new_n18421_), .ZN(new_n18422_));
  AOI21_X1   g15986(.A1(new_n18420_), .A2(new_n18422_), .B(new_n16430_), .ZN(new_n18423_));
  INV_X1     g15987(.I(new_n15113_), .ZN(new_n18424_));
  INV_X1     g15988(.I(new_n15114_), .ZN(new_n18425_));
  INV_X1     g15989(.I(new_n13599_), .ZN(new_n18426_));
  NAND2_X1   g15990(.A1(new_n13632_), .A2(new_n2642_), .ZN(new_n18427_));
  AOI21_X1   g15991(.A1(new_n5445_), .A2(new_n13615_), .B(new_n18427_), .ZN(new_n18428_));
  OAI21_X1   g15992(.A1(new_n18428_), .A2(new_n18426_), .B(new_n13595_), .ZN(new_n18429_));
  INV_X1     g15993(.I(new_n13640_), .ZN(new_n18430_));
  NAND4_X1   g15994(.A1(new_n13631_), .A2(new_n13624_), .A3(new_n13619_), .A4(new_n5422_), .ZN(new_n18431_));
  NAND3_X1   g15995(.A1(new_n14714_), .A2(new_n6764_), .A3(new_n14709_), .ZN(new_n18432_));
  NAND2_X1   g15996(.A1(new_n18432_), .A2(new_n18431_), .ZN(new_n18433_));
  AOI21_X1   g15997(.A1(new_n18433_), .A2(new_n3304_), .B(new_n18430_), .ZN(new_n18434_));
  OAI21_X1   g15998(.A1(new_n18434_), .A2(new_n13637_), .B(pi0299), .ZN(new_n18435_));
  AOI21_X1   g15999(.A1(new_n18429_), .A2(new_n18435_), .B(new_n2627_), .ZN(new_n18436_));
  OAI21_X1   g16000(.A1(new_n18436_), .A2(new_n18425_), .B(new_n3265_), .ZN(new_n18437_));
  NAND2_X1   g16001(.A1(new_n18437_), .A2(new_n18424_), .ZN(new_n18438_));
  NAND2_X1   g16002(.A1(new_n18438_), .A2(pi0176), .ZN(new_n18439_));
  NAND2_X1   g16003(.A1(new_n15111_), .A2(new_n7518_), .ZN(new_n18440_));
  AOI21_X1   g16004(.A1(new_n18439_), .A2(new_n18440_), .B(pi0742), .ZN(new_n18441_));
  NOR3_X1    g16005(.A1(new_n18423_), .A2(pi0704), .A3(new_n18441_), .ZN(new_n18442_));
  OAI21_X1   g16006(.A1(new_n18442_), .A2(new_n18417_), .B(new_n2609_), .ZN(new_n18443_));
  OAI21_X1   g16007(.A1(pi0176), .A2(new_n2609_), .B(new_n18443_), .ZN(new_n18444_));
  NOR2_X1    g16008(.A1(new_n18444_), .A2(pi0625), .ZN(new_n18445_));
  NOR2_X1    g16009(.A1(new_n18334_), .A2(new_n13521_), .ZN(new_n18446_));
  OAI21_X1   g16010(.A1(new_n18445_), .A2(new_n18446_), .B(new_n12841_), .ZN(new_n18447_));
  NAND3_X1   g16011(.A1(new_n18447_), .A2(new_n13560_), .A3(new_n18380_), .ZN(new_n18448_));
  NOR2_X1    g16012(.A1(new_n18444_), .A2(new_n13521_), .ZN(new_n18449_));
  NOR2_X1    g16013(.A1(new_n18334_), .A2(pi0625), .ZN(new_n18450_));
  OAI21_X1   g16014(.A1(new_n18449_), .A2(new_n18450_), .B(pi1153), .ZN(new_n18451_));
  NAND3_X1   g16015(.A1(new_n18451_), .A2(pi0608), .A3(new_n18377_), .ZN(new_n18452_));
  NAND3_X1   g16016(.A1(new_n18448_), .A2(new_n18452_), .A3(pi0778), .ZN(new_n18453_));
  OAI21_X1   g16017(.A1(pi0778), .A2(new_n18444_), .B(new_n18453_), .ZN(new_n18454_));
  NAND2_X1   g16018(.A1(new_n18454_), .A2(pi0609), .ZN(new_n18455_));
  AOI21_X1   g16019(.A1(new_n18455_), .A2(new_n18416_), .B(new_n12770_), .ZN(new_n18456_));
  NOR3_X1    g16020(.A1(new_n18456_), .A2(new_n13829_), .A3(new_n18341_), .ZN(new_n18457_));
  NAND2_X1   g16021(.A1(new_n18454_), .A2(new_n12766_), .ZN(new_n18458_));
  OAI21_X1   g16022(.A1(new_n12766_), .A2(new_n18382_), .B(new_n18458_), .ZN(new_n18459_));
  NAND2_X1   g16023(.A1(new_n18343_), .A2(new_n13829_), .ZN(new_n18460_));
  AOI21_X1   g16024(.A1(new_n18459_), .A2(new_n12770_), .B(new_n18460_), .ZN(new_n18461_));
  NOR3_X1    g16025(.A1(new_n18461_), .A2(new_n18457_), .A3(new_n12764_), .ZN(new_n18462_));
  NAND2_X1   g16026(.A1(new_n18454_), .A2(new_n12764_), .ZN(new_n18463_));
  INV_X1     g16027(.I(new_n18463_), .ZN(new_n18464_));
  NOR2_X1    g16028(.A1(new_n18462_), .A2(new_n18464_), .ZN(new_n18465_));
  AND2_X2    g16029(.A1(new_n18383_), .A2(new_n12781_), .Z(new_n18466_));
  NOR2_X1    g16030(.A1(new_n18465_), .A2(new_n12781_), .ZN(new_n18467_));
  OAI21_X1   g16031(.A1(new_n18467_), .A2(new_n18466_), .B(pi1154), .ZN(new_n18468_));
  AND3_X2    g16032(.A1(new_n18468_), .A2(pi0627), .A3(new_n18349_), .Z(new_n18469_));
  INV_X1     g16033(.I(new_n18352_), .ZN(new_n18470_));
  OAI21_X1   g16034(.A1(new_n18462_), .A2(new_n18464_), .B(new_n12781_), .ZN(new_n18471_));
  NAND2_X1   g16035(.A1(new_n18383_), .A2(pi0618), .ZN(new_n18472_));
  AOI21_X1   g16036(.A1(new_n18471_), .A2(new_n18472_), .B(pi1154), .ZN(new_n18473_));
  NOR3_X1    g16037(.A1(new_n18473_), .A2(pi0627), .A3(new_n18470_), .ZN(new_n18474_));
  OR2_X2     g16038(.A1(new_n18474_), .A2(new_n12779_), .Z(new_n18475_));
  OAI22_X1   g16039(.A1(new_n18475_), .A2(new_n18469_), .B1(pi0781), .B2(new_n18465_), .ZN(new_n18476_));
  NAND2_X1   g16040(.A1(new_n18476_), .A2(new_n12796_), .ZN(new_n18477_));
  NAND2_X1   g16041(.A1(new_n18477_), .A2(new_n12819_), .ZN(new_n18478_));
  AOI21_X1   g16042(.A1(new_n18319_), .A2(pi0619), .B(pi1159), .ZN(new_n18479_));
  NAND2_X1   g16043(.A1(new_n18354_), .A2(new_n12793_), .ZN(new_n18480_));
  AOI21_X1   g16044(.A1(new_n18480_), .A2(new_n18479_), .B(new_n12895_), .ZN(new_n18481_));
  OAI21_X1   g16045(.A1(new_n18386_), .A2(pi0619), .B(pi1159), .ZN(new_n18482_));
  NOR2_X1    g16046(.A1(new_n18476_), .A2(new_n12793_), .ZN(new_n18483_));
  OAI21_X1   g16047(.A1(new_n18483_), .A2(new_n18482_), .B(new_n18481_), .ZN(new_n18484_));
  AOI21_X1   g16048(.A1(new_n18319_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n18485_));
  NAND2_X1   g16049(.A1(new_n18354_), .A2(pi0619), .ZN(new_n18486_));
  AOI21_X1   g16050(.A1(new_n18486_), .A2(new_n18485_), .B(pi0648), .ZN(new_n18487_));
  AOI21_X1   g16051(.A1(new_n18385_), .A2(pi0619), .B(pi1159), .ZN(new_n18488_));
  OAI21_X1   g16052(.A1(new_n18476_), .A2(pi0619), .B(new_n18488_), .ZN(new_n18489_));
  AOI21_X1   g16053(.A1(new_n18489_), .A2(new_n18487_), .B(new_n12796_), .ZN(new_n18490_));
  AOI21_X1   g16054(.A1(new_n18490_), .A2(new_n18484_), .B(new_n18478_), .ZN(new_n18491_));
  NAND2_X1   g16055(.A1(new_n18319_), .A2(new_n12747_), .ZN(new_n18492_));
  OAI21_X1   g16056(.A1(new_n18356_), .A2(new_n12747_), .B(new_n18492_), .ZN(new_n18493_));
  NAND2_X1   g16057(.A1(new_n18493_), .A2(new_n12812_), .ZN(new_n18494_));
  NAND2_X1   g16058(.A1(new_n18319_), .A2(new_n12910_), .ZN(new_n18495_));
  OAI21_X1   g16059(.A1(new_n18386_), .A2(new_n12910_), .B(new_n18495_), .ZN(new_n18496_));
  NAND2_X1   g16060(.A1(new_n18319_), .A2(pi0626), .ZN(new_n18497_));
  OAI21_X1   g16061(.A1(new_n18356_), .A2(pi0626), .B(new_n18497_), .ZN(new_n18498_));
  AOI22_X1   g16062(.A1(new_n18498_), .A2(new_n12815_), .B1(new_n14386_), .B2(new_n18496_), .ZN(new_n18499_));
  AOI21_X1   g16063(.A1(new_n18499_), .A2(new_n18494_), .B(new_n12808_), .ZN(new_n18500_));
  OAI22_X1   g16064(.A1(new_n18491_), .A2(new_n18500_), .B1(new_n12937_), .B2(new_n18414_), .ZN(new_n18501_));
  NOR2_X1    g16065(.A1(new_n18404_), .A2(new_n12975_), .ZN(new_n18502_));
  NOR2_X1    g16066(.A1(new_n18363_), .A2(pi0644), .ZN(new_n18503_));
  NOR2_X1    g16067(.A1(new_n18502_), .A2(new_n18503_), .ZN(new_n18504_));
  OAI22_X1   g16068(.A1(new_n15576_), .A2(new_n18393_), .B1(new_n18396_), .B2(new_n15730_), .ZN(new_n18505_));
  NOR2_X1    g16069(.A1(new_n18360_), .A2(new_n17212_), .ZN(new_n18506_));
  NOR2_X1    g16070(.A1(new_n18506_), .A2(new_n18505_), .ZN(new_n18507_));
  OAI22_X1   g16071(.A1(new_n18504_), .A2(new_n13000_), .B1(new_n12972_), .B2(new_n18507_), .ZN(new_n18508_));
  AOI21_X1   g16072(.A1(new_n18501_), .A2(new_n18415_), .B(new_n18508_), .ZN(new_n18509_));
  OAI21_X1   g16073(.A1(new_n18509_), .A2(new_n18407_), .B(new_n6643_), .ZN(new_n18510_));
  AOI22_X1   g16074(.A1(new_n18510_), .A2(new_n18318_), .B1(pi0832), .B2(new_n18317_), .ZN(po0333));
  NOR2_X1    g16075(.A1(new_n3042_), .A2(pi0177), .ZN(new_n18512_));
  INV_X1     g16076(.I(new_n18512_), .ZN(new_n18513_));
  AOI21_X1   g16077(.A1(new_n12756_), .A2(new_n16460_), .B(new_n18512_), .ZN(new_n18514_));
  NOR3_X1    g16078(.A1(new_n18514_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n18515_));
  NOR2_X1    g16079(.A1(new_n18514_), .A2(new_n12762_), .ZN(new_n18516_));
  AOI21_X1   g16080(.A1(new_n18516_), .A2(new_n12768_), .B(pi1155), .ZN(new_n18517_));
  INV_X1     g16081(.I(new_n18514_), .ZN(new_n18518_));
  AOI21_X1   g16082(.A1(new_n18518_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n18519_));
  NOR3_X1    g16083(.A1(new_n18517_), .A2(new_n18519_), .A3(new_n12764_), .ZN(new_n18520_));
  NOR2_X1    g16084(.A1(new_n18520_), .A2(new_n18515_), .ZN(new_n18521_));
  NOR2_X1    g16085(.A1(new_n18521_), .A2(pi0781), .ZN(new_n18522_));
  INV_X1     g16086(.I(new_n18521_), .ZN(new_n18523_));
  AOI21_X1   g16087(.A1(new_n18523_), .A2(new_n12783_), .B(pi1154), .ZN(new_n18524_));
  AOI21_X1   g16088(.A1(new_n18523_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n18525_));
  NOR3_X1    g16089(.A1(new_n18524_), .A2(new_n18525_), .A3(new_n12779_), .ZN(new_n18526_));
  NOR2_X1    g16090(.A1(new_n18526_), .A2(new_n18522_), .ZN(new_n18527_));
  NOR3_X1    g16091(.A1(new_n18526_), .A2(pi0619), .A3(new_n18522_), .ZN(new_n18528_));
  NOR2_X1    g16092(.A1(new_n18512_), .A2(new_n12793_), .ZN(new_n18529_));
  OAI21_X1   g16093(.A1(new_n18528_), .A2(new_n18529_), .B(new_n12791_), .ZN(new_n18530_));
  NAND2_X1   g16094(.A1(new_n18527_), .A2(pi0619), .ZN(new_n18531_));
  NAND2_X1   g16095(.A1(new_n18513_), .A2(new_n12793_), .ZN(new_n18532_));
  AOI21_X1   g16096(.A1(new_n18531_), .A2(new_n18532_), .B(new_n12791_), .ZN(new_n18533_));
  INV_X1     g16097(.I(new_n18533_), .ZN(new_n18534_));
  NAND3_X1   g16098(.A1(new_n18534_), .A2(pi0789), .A3(new_n18530_), .ZN(new_n18535_));
  OAI21_X1   g16099(.A1(pi0789), .A2(new_n18527_), .B(new_n18535_), .ZN(new_n18536_));
  NOR2_X1    g16100(.A1(new_n18536_), .A2(new_n12818_), .ZN(new_n18537_));
  AOI21_X1   g16101(.A1(new_n12818_), .A2(new_n18513_), .B(new_n18537_), .ZN(new_n18538_));
  AOI21_X1   g16102(.A1(new_n12826_), .A2(new_n16459_), .B(new_n18512_), .ZN(new_n18539_));
  NOR2_X1    g16103(.A1(new_n18539_), .A2(pi0778), .ZN(new_n18540_));
  NOR2_X1    g16104(.A1(new_n18512_), .A2(pi1153), .ZN(new_n18541_));
  NOR2_X1    g16105(.A1(new_n12834_), .A2(pi0686), .ZN(new_n18542_));
  INV_X1     g16106(.I(new_n18542_), .ZN(new_n18543_));
  NAND2_X1   g16107(.A1(new_n18543_), .A2(new_n18541_), .ZN(new_n18544_));
  INV_X1     g16108(.I(new_n18544_), .ZN(new_n18545_));
  NOR2_X1    g16109(.A1(new_n18542_), .A2(new_n18539_), .ZN(new_n18546_));
  NOR2_X1    g16110(.A1(new_n18546_), .A2(new_n12841_), .ZN(new_n18547_));
  NOR2_X1    g16111(.A1(new_n18545_), .A2(new_n18547_), .ZN(new_n18548_));
  AOI21_X1   g16112(.A1(new_n18548_), .A2(pi0778), .B(new_n18540_), .ZN(new_n18549_));
  NOR2_X1    g16113(.A1(new_n18549_), .A2(new_n12871_), .ZN(new_n18550_));
  INV_X1     g16114(.I(new_n18550_), .ZN(new_n18551_));
  NOR2_X1    g16115(.A1(new_n18551_), .A2(new_n12889_), .ZN(new_n18552_));
  NAND2_X1   g16116(.A1(new_n18552_), .A2(new_n18203_), .ZN(new_n18553_));
  NOR2_X1    g16117(.A1(new_n18553_), .A2(new_n17884_), .ZN(new_n18554_));
  AOI22_X1   g16118(.A1(new_n18538_), .A2(new_n12949_), .B1(new_n15695_), .B2(new_n18554_), .ZN(new_n18555_));
  NOR2_X1    g16119(.A1(new_n18555_), .A2(pi0629), .ZN(new_n18556_));
  AOI22_X1   g16120(.A1(new_n18538_), .A2(new_n12948_), .B1(new_n15700_), .B2(new_n18554_), .ZN(new_n18557_));
  NOR2_X1    g16121(.A1(new_n18557_), .A2(new_n12919_), .ZN(new_n18558_));
  NOR2_X1    g16122(.A1(new_n18556_), .A2(new_n18558_), .ZN(new_n18559_));
  NOR2_X1    g16123(.A1(new_n18539_), .A2(new_n12754_), .ZN(new_n18560_));
  NOR2_X1    g16124(.A1(new_n18560_), .A2(new_n18518_), .ZN(new_n18561_));
  NAND2_X1   g16125(.A1(new_n18561_), .A2(new_n12758_), .ZN(new_n18562_));
  NAND2_X1   g16126(.A1(new_n18560_), .A2(pi0625), .ZN(new_n18563_));
  NAND3_X1   g16127(.A1(new_n18563_), .A2(pi1153), .A3(new_n18514_), .ZN(new_n18564_));
  AND3_X2    g16128(.A1(new_n18544_), .A2(pi0608), .A3(new_n18564_), .Z(new_n18565_));
  NOR2_X1    g16129(.A1(new_n18547_), .A2(pi0608), .ZN(new_n18566_));
  INV_X1     g16130(.I(new_n18563_), .ZN(new_n18567_));
  OAI21_X1   g16131(.A1(new_n18567_), .A2(new_n18561_), .B(new_n18541_), .ZN(new_n18568_));
  NAND2_X1   g16132(.A1(new_n18566_), .A2(new_n18568_), .ZN(new_n18569_));
  NAND2_X1   g16133(.A1(new_n18569_), .A2(pi0778), .ZN(new_n18570_));
  OAI21_X1   g16134(.A1(new_n18570_), .A2(new_n18565_), .B(new_n18562_), .ZN(new_n18571_));
  INV_X1     g16135(.I(new_n18571_), .ZN(new_n18572_));
  NAND2_X1   g16136(.A1(new_n18549_), .A2(new_n12766_), .ZN(new_n18573_));
  OAI21_X1   g16137(.A1(new_n18572_), .A2(new_n12766_), .B(new_n18573_), .ZN(new_n18574_));
  AOI21_X1   g16138(.A1(new_n18574_), .A2(pi1155), .B(new_n18517_), .ZN(new_n18575_));
  NAND2_X1   g16139(.A1(new_n18571_), .A2(new_n12766_), .ZN(new_n18576_));
  NAND2_X1   g16140(.A1(new_n18549_), .A2(pi0609), .ZN(new_n18577_));
  AOI21_X1   g16141(.A1(new_n18576_), .A2(new_n18577_), .B(pi1155), .ZN(new_n18578_));
  NOR3_X1    g16142(.A1(new_n18578_), .A2(pi0660), .A3(new_n18519_), .ZN(new_n18579_));
  AOI21_X1   g16143(.A1(pi0660), .A2(new_n18575_), .B(new_n18579_), .ZN(new_n18580_));
  NAND2_X1   g16144(.A1(new_n18580_), .A2(pi0785), .ZN(new_n18581_));
  OAI21_X1   g16145(.A1(pi0785), .A2(new_n18572_), .B(new_n18581_), .ZN(new_n18582_));
  INV_X1     g16146(.I(new_n18582_), .ZN(new_n18583_));
  NAND2_X1   g16147(.A1(new_n18551_), .A2(pi0618), .ZN(new_n18584_));
  OAI21_X1   g16148(.A1(new_n18583_), .A2(pi0618), .B(new_n18584_), .ZN(new_n18585_));
  AOI21_X1   g16149(.A1(new_n18585_), .A2(new_n12785_), .B(new_n18525_), .ZN(new_n18586_));
  NOR2_X1    g16150(.A1(new_n18550_), .A2(pi0618), .ZN(new_n18587_));
  NOR2_X1    g16151(.A1(new_n18583_), .A2(new_n12781_), .ZN(new_n18588_));
  OAI21_X1   g16152(.A1(new_n18588_), .A2(new_n18587_), .B(pi1154), .ZN(new_n18589_));
  NOR2_X1    g16153(.A1(new_n18524_), .A2(new_n12880_), .ZN(new_n18590_));
  AOI22_X1   g16154(.A1(new_n18586_), .A2(new_n12880_), .B1(new_n18589_), .B2(new_n18590_), .ZN(new_n18591_));
  NAND2_X1   g16155(.A1(new_n18591_), .A2(pi0781), .ZN(new_n18592_));
  NAND2_X1   g16156(.A1(new_n18582_), .A2(new_n12779_), .ZN(new_n18593_));
  NAND2_X1   g16157(.A1(new_n18592_), .A2(new_n18593_), .ZN(new_n18594_));
  AOI21_X1   g16158(.A1(new_n18594_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n18595_));
  NOR2_X1    g16159(.A1(new_n18552_), .A2(pi0619), .ZN(new_n18596_));
  INV_X1     g16160(.I(new_n18594_), .ZN(new_n18597_));
  NOR2_X1    g16161(.A1(new_n18597_), .A2(new_n12793_), .ZN(new_n18598_));
  OAI21_X1   g16162(.A1(new_n18598_), .A2(new_n18596_), .B(pi1159), .ZN(new_n18599_));
  NAND3_X1   g16163(.A1(new_n18599_), .A2(pi0648), .A3(new_n18530_), .ZN(new_n18600_));
  NOR2_X1    g16164(.A1(new_n18597_), .A2(pi0619), .ZN(new_n18601_));
  NOR2_X1    g16165(.A1(new_n18552_), .A2(new_n12793_), .ZN(new_n18602_));
  OAI21_X1   g16166(.A1(new_n18601_), .A2(new_n18602_), .B(new_n12791_), .ZN(new_n18603_));
  NAND3_X1   g16167(.A1(new_n18603_), .A2(new_n12895_), .A3(new_n18534_), .ZN(new_n18604_));
  NAND3_X1   g16168(.A1(new_n18600_), .A2(new_n18604_), .A3(pi0789), .ZN(new_n18605_));
  NOR2_X1    g16169(.A1(new_n18513_), .A2(new_n12747_), .ZN(new_n18606_));
  INV_X1     g16170(.I(new_n18536_), .ZN(new_n18607_));
  NOR2_X1    g16171(.A1(new_n18607_), .A2(pi0626), .ZN(new_n18608_));
  OAI21_X1   g16172(.A1(new_n18608_), .A2(new_n18606_), .B(new_n12815_), .ZN(new_n18609_));
  INV_X1     g16173(.I(new_n18553_), .ZN(new_n18610_));
  NAND2_X1   g16174(.A1(new_n18512_), .A2(new_n12747_), .ZN(new_n18611_));
  OAI21_X1   g16175(.A1(new_n18607_), .A2(new_n12747_), .B(new_n18611_), .ZN(new_n18612_));
  AOI22_X1   g16176(.A1(new_n18612_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n18610_), .ZN(new_n18613_));
  NAND2_X1   g16177(.A1(new_n18613_), .A2(new_n18609_), .ZN(new_n18614_));
  AOI22_X1   g16178(.A1(new_n18605_), .A2(new_n18595_), .B1(pi0788), .B2(new_n18614_), .ZN(new_n18615_));
  OAI22_X1   g16179(.A1(new_n18615_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n18559_), .ZN(new_n18616_));
  INV_X1     g16180(.I(new_n18538_), .ZN(new_n18617_));
  NAND2_X1   g16181(.A1(new_n18617_), .A2(new_n13384_), .ZN(new_n18618_));
  NAND2_X1   g16182(.A1(new_n12943_), .A2(new_n18513_), .ZN(new_n18619_));
  NAND2_X1   g16183(.A1(new_n18618_), .A2(new_n18619_), .ZN(new_n18620_));
  NAND2_X1   g16184(.A1(new_n18554_), .A2(new_n12954_), .ZN(new_n18621_));
  NAND2_X1   g16185(.A1(new_n18621_), .A2(new_n12741_), .ZN(new_n18622_));
  NOR2_X1    g16186(.A1(new_n18512_), .A2(new_n12741_), .ZN(new_n18623_));
  INV_X1     g16187(.I(new_n18623_), .ZN(new_n18624_));
  AOI21_X1   g16188(.A1(new_n18622_), .A2(new_n18624_), .B(pi1157), .ZN(new_n18625_));
  INV_X1     g16189(.I(new_n18625_), .ZN(new_n18626_));
  NAND2_X1   g16190(.A1(new_n18512_), .A2(new_n12741_), .ZN(new_n18627_));
  OAI21_X1   g16191(.A1(new_n18621_), .A2(new_n12741_), .B(new_n18627_), .ZN(new_n18628_));
  OAI22_X1   g16192(.A1(new_n18626_), .A2(new_n12981_), .B1(new_n18628_), .B2(new_n15576_), .ZN(new_n18629_));
  AOI21_X1   g16193(.A1(new_n18620_), .A2(new_n15608_), .B(new_n18629_), .ZN(new_n18630_));
  OAI22_X1   g16194(.A1(new_n18616_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n18630_), .ZN(new_n18631_));
  NAND2_X1   g16195(.A1(new_n18631_), .A2(new_n13000_), .ZN(new_n18632_));
  AND2_X2    g16196(.A1(new_n18631_), .A2(new_n12975_), .Z(new_n18633_));
  OAI21_X1   g16197(.A1(new_n12965_), .A2(new_n18628_), .B(new_n18626_), .ZN(new_n18634_));
  NAND3_X1   g16198(.A1(new_n18554_), .A2(new_n12972_), .A3(new_n12954_), .ZN(new_n18635_));
  OAI21_X1   g16199(.A1(new_n18634_), .A2(new_n12972_), .B(new_n18635_), .ZN(new_n18636_));
  NOR2_X1    g16200(.A1(new_n18636_), .A2(new_n12975_), .ZN(new_n18637_));
  OAI21_X1   g16201(.A1(new_n18633_), .A2(new_n18637_), .B(new_n12740_), .ZN(new_n18638_));
  NOR2_X1    g16202(.A1(new_n18512_), .A2(new_n12975_), .ZN(new_n18639_));
  NOR2_X1    g16203(.A1(new_n17611_), .A2(new_n18512_), .ZN(new_n18640_));
  AOI21_X1   g16204(.A1(new_n18617_), .A2(new_n17611_), .B(new_n18640_), .ZN(new_n18641_));
  NOR2_X1    g16205(.A1(new_n18641_), .A2(pi0644), .ZN(new_n18642_));
  OAI21_X1   g16206(.A1(new_n18642_), .A2(new_n18639_), .B(pi0715), .ZN(new_n18643_));
  NAND3_X1   g16207(.A1(new_n18638_), .A2(new_n12739_), .A3(new_n18643_), .ZN(new_n18644_));
  NOR2_X1    g16208(.A1(new_n18636_), .A2(pi0644), .ZN(new_n18645_));
  AOI21_X1   g16209(.A1(new_n18631_), .A2(pi0644), .B(new_n18645_), .ZN(new_n18646_));
  NAND2_X1   g16210(.A1(new_n18513_), .A2(new_n12975_), .ZN(new_n18647_));
  OAI21_X1   g16211(.A1(new_n18641_), .A2(new_n12975_), .B(new_n18647_), .ZN(new_n18648_));
  AOI21_X1   g16212(.A1(new_n18648_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n18649_));
  OAI21_X1   g16213(.A1(new_n18646_), .A2(new_n12740_), .B(new_n18649_), .ZN(new_n18650_));
  NAND3_X1   g16214(.A1(new_n18644_), .A2(pi0790), .A3(new_n18650_), .ZN(new_n18651_));
  AOI21_X1   g16215(.A1(new_n18651_), .A2(new_n18632_), .B(new_n12738_), .ZN(new_n18652_));
  AOI21_X1   g16216(.A1(po1038), .A2(new_n8056_), .B(pi0832), .ZN(new_n18653_));
  NOR2_X1    g16217(.A1(new_n13193_), .A2(pi0177), .ZN(new_n18654_));
  INV_X1     g16218(.I(new_n18654_), .ZN(new_n18655_));
  OAI21_X1   g16219(.A1(new_n18655_), .A2(new_n12975_), .B(pi0715), .ZN(new_n18656_));
  NOR2_X1    g16220(.A1(new_n18654_), .A2(new_n13384_), .ZN(new_n18657_));
  NOR2_X1    g16221(.A1(new_n2609_), .A2(new_n8056_), .ZN(new_n18658_));
  INV_X1     g16222(.I(new_n15008_), .ZN(new_n18659_));
  NAND3_X1   g16223(.A1(new_n13245_), .A2(new_n3265_), .A3(pi0177), .ZN(new_n18660_));
  AOI21_X1   g16224(.A1(new_n18660_), .A2(new_n18659_), .B(pi0757), .ZN(new_n18661_));
  OAI21_X1   g16225(.A1(new_n15012_), .A2(new_n15011_), .B(new_n16460_), .ZN(new_n18662_));
  AOI21_X1   g16226(.A1(new_n18662_), .A2(new_n16465_), .B(pi0177), .ZN(new_n18663_));
  NOR2_X1    g16227(.A1(new_n18663_), .A2(new_n18661_), .ZN(new_n18664_));
  AOI21_X1   g16228(.A1(new_n18664_), .A2(new_n2609_), .B(new_n18658_), .ZN(new_n18665_));
  NOR2_X1    g16229(.A1(new_n18665_), .A2(new_n12760_), .ZN(new_n18666_));
  NOR2_X1    g16230(.A1(new_n18654_), .A2(new_n12761_), .ZN(new_n18667_));
  NOR3_X1    g16231(.A1(new_n18666_), .A2(pi0785), .A3(new_n18667_), .ZN(new_n18668_));
  AOI22_X1   g16232(.A1(new_n18666_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n18655_), .ZN(new_n18669_));
  OR2_X2     g16233(.A1(new_n18669_), .A2(pi1155), .Z(new_n18670_));
  AOI22_X1   g16234(.A1(new_n18666_), .A2(pi0609), .B1(new_n13357_), .B2(new_n18655_), .ZN(new_n18671_));
  NOR2_X1    g16235(.A1(new_n18671_), .A2(new_n12770_), .ZN(new_n18672_));
  NOR2_X1    g16236(.A1(new_n18672_), .A2(new_n12764_), .ZN(new_n18673_));
  AOI21_X1   g16237(.A1(new_n18673_), .A2(new_n18670_), .B(new_n18668_), .ZN(new_n18674_));
  NOR2_X1    g16238(.A1(new_n18654_), .A2(new_n12781_), .ZN(new_n18675_));
  AOI21_X1   g16239(.A1(new_n18674_), .A2(new_n12781_), .B(new_n18675_), .ZN(new_n18676_));
  NOR2_X1    g16240(.A1(new_n18676_), .A2(pi1154), .ZN(new_n18677_));
  NOR2_X1    g16241(.A1(new_n18654_), .A2(pi0618), .ZN(new_n18678_));
  AOI21_X1   g16242(.A1(new_n18674_), .A2(pi0618), .B(new_n18678_), .ZN(new_n18679_));
  OAI21_X1   g16243(.A1(new_n18679_), .A2(new_n12785_), .B(pi0781), .ZN(new_n18680_));
  OAI22_X1   g16244(.A1(new_n18680_), .A2(new_n18677_), .B1(pi0781), .B2(new_n18674_), .ZN(new_n18681_));
  NAND2_X1   g16245(.A1(new_n18681_), .A2(new_n12796_), .ZN(new_n18682_));
  NAND2_X1   g16246(.A1(new_n18655_), .A2(pi0619), .ZN(new_n18683_));
  OAI21_X1   g16247(.A1(new_n18681_), .A2(pi0619), .B(new_n18683_), .ZN(new_n18684_));
  NAND2_X1   g16248(.A1(new_n18684_), .A2(new_n12791_), .ZN(new_n18685_));
  NAND2_X1   g16249(.A1(new_n18655_), .A2(new_n12793_), .ZN(new_n18686_));
  OAI21_X1   g16250(.A1(new_n18681_), .A2(new_n12793_), .B(new_n18686_), .ZN(new_n18687_));
  AOI21_X1   g16251(.A1(new_n18687_), .A2(pi1159), .B(new_n12796_), .ZN(new_n18688_));
  NAND2_X1   g16252(.A1(new_n18688_), .A2(new_n18685_), .ZN(new_n18689_));
  NAND3_X1   g16253(.A1(new_n18689_), .A2(new_n17504_), .A3(new_n18682_), .ZN(new_n18690_));
  OAI21_X1   g16254(.A1(new_n17504_), .A2(new_n18654_), .B(new_n18690_), .ZN(new_n18691_));
  AOI21_X1   g16255(.A1(new_n18691_), .A2(new_n13384_), .B(new_n18657_), .ZN(new_n18692_));
  NOR2_X1    g16256(.A1(new_n18655_), .A2(new_n12985_), .ZN(new_n18693_));
  AOI21_X1   g16257(.A1(new_n18692_), .A2(new_n12985_), .B(new_n18693_), .ZN(new_n18694_));
  NOR2_X1    g16258(.A1(new_n18694_), .A2(pi0644), .ZN(new_n18695_));
  OAI21_X1   g16259(.A1(new_n18695_), .A2(new_n18656_), .B(new_n12739_), .ZN(new_n18696_));
  NOR2_X1    g16260(.A1(new_n18655_), .A2(new_n12870_), .ZN(new_n18697_));
  INV_X1     g16261(.I(new_n18658_), .ZN(new_n18698_));
  NOR2_X1    g16262(.A1(new_n16459_), .A2(pi0177), .ZN(new_n18699_));
  INV_X1     g16263(.I(new_n18699_), .ZN(new_n18700_));
  OAI21_X1   g16264(.A1(new_n13191_), .A2(new_n18700_), .B(new_n2609_), .ZN(new_n18701_));
  NAND2_X1   g16265(.A1(new_n14122_), .A2(pi0177), .ZN(new_n18702_));
  OAI21_X1   g16266(.A1(new_n15744_), .A2(pi0177), .B(new_n18702_), .ZN(new_n18703_));
  NOR2_X1    g16267(.A1(new_n13344_), .A2(pi0177), .ZN(new_n18704_));
  INV_X1     g16268(.I(new_n18704_), .ZN(new_n18705_));
  AOI21_X1   g16269(.A1(new_n13399_), .A2(new_n18705_), .B(pi0686), .ZN(new_n18706_));
  INV_X1     g16270(.I(new_n18706_), .ZN(new_n18707_));
  AOI21_X1   g16271(.A1(new_n18703_), .A2(new_n3265_), .B(new_n18707_), .ZN(new_n18708_));
  OAI21_X1   g16272(.A1(new_n18708_), .A2(new_n18701_), .B(new_n18698_), .ZN(new_n18709_));
  NOR2_X1    g16273(.A1(new_n18709_), .A2(new_n14131_), .ZN(new_n18710_));
  NOR3_X1    g16274(.A1(new_n18655_), .A2(new_n12758_), .A3(new_n14132_), .ZN(new_n18711_));
  NOR2_X1    g16275(.A1(new_n18710_), .A2(new_n18711_), .ZN(new_n18712_));
  INV_X1     g16276(.I(new_n18712_), .ZN(new_n18713_));
  AOI21_X1   g16277(.A1(new_n18713_), .A2(new_n12870_), .B(new_n18697_), .ZN(new_n18714_));
  NOR2_X1    g16278(.A1(new_n18654_), .A2(new_n12888_), .ZN(new_n18715_));
  AOI21_X1   g16279(.A1(new_n18714_), .A2(new_n12888_), .B(new_n18715_), .ZN(new_n18716_));
  NOR2_X1    g16280(.A1(new_n18655_), .A2(new_n12911_), .ZN(new_n18717_));
  AOI21_X1   g16281(.A1(new_n18716_), .A2(new_n12911_), .B(new_n18717_), .ZN(new_n18718_));
  INV_X1     g16282(.I(new_n18718_), .ZN(new_n18719_));
  NOR2_X1    g16283(.A1(new_n18719_), .A2(new_n12817_), .ZN(new_n18720_));
  AOI21_X1   g16284(.A1(new_n12817_), .A2(new_n18655_), .B(new_n18720_), .ZN(new_n18721_));
  INV_X1     g16285(.I(new_n18721_), .ZN(new_n18722_));
  NAND2_X1   g16286(.A1(new_n18722_), .A2(new_n12920_), .ZN(new_n18723_));
  NAND2_X1   g16287(.A1(new_n18655_), .A2(pi0628), .ZN(new_n18724_));
  AOI21_X1   g16288(.A1(new_n18723_), .A2(new_n18724_), .B(pi1156), .ZN(new_n18725_));
  INV_X1     g16289(.I(new_n18725_), .ZN(new_n18726_));
  NOR2_X1    g16290(.A1(new_n18654_), .A2(pi0628), .ZN(new_n18727_));
  AOI21_X1   g16291(.A1(new_n18722_), .A2(pi0628), .B(new_n18727_), .ZN(new_n18728_));
  NOR2_X1    g16292(.A1(new_n18728_), .A2(new_n12742_), .ZN(new_n18729_));
  NOR2_X1    g16293(.A1(new_n18729_), .A2(new_n12937_), .ZN(new_n18730_));
  AOI22_X1   g16294(.A1(new_n18730_), .A2(new_n18726_), .B1(new_n12937_), .B2(new_n18721_), .ZN(new_n18731_));
  NAND2_X1   g16295(.A1(new_n18731_), .A2(new_n12741_), .ZN(new_n18732_));
  OAI21_X1   g16296(.A1(new_n12741_), .A2(new_n18654_), .B(new_n18732_), .ZN(new_n18733_));
  NAND2_X1   g16297(.A1(new_n18733_), .A2(new_n12965_), .ZN(new_n18734_));
  NOR2_X1    g16298(.A1(new_n18654_), .A2(pi0647), .ZN(new_n18735_));
  AOI21_X1   g16299(.A1(new_n18731_), .A2(pi0647), .B(new_n18735_), .ZN(new_n18736_));
  NOR2_X1    g16300(.A1(new_n18736_), .A2(new_n12965_), .ZN(new_n18737_));
  NOR2_X1    g16301(.A1(new_n18737_), .A2(new_n12972_), .ZN(new_n18738_));
  NAND2_X1   g16302(.A1(new_n18738_), .A2(new_n18734_), .ZN(new_n18739_));
  OAI21_X1   g16303(.A1(pi0787), .A2(new_n18731_), .B(new_n18739_), .ZN(new_n18740_));
  AOI21_X1   g16304(.A1(new_n18740_), .A2(pi0644), .B(pi0715), .ZN(new_n18741_));
  NOR2_X1    g16305(.A1(new_n18725_), .A2(new_n12919_), .ZN(new_n18742_));
  OAI21_X1   g16306(.A1(new_n18691_), .A2(pi0628), .B(pi1156), .ZN(new_n18743_));
  AOI21_X1   g16307(.A1(new_n18655_), .A2(new_n12747_), .B(pi0641), .ZN(new_n18744_));
  NAND3_X1   g16308(.A1(new_n18689_), .A2(pi0626), .A3(new_n18682_), .ZN(new_n18745_));
  AOI21_X1   g16309(.A1(new_n18745_), .A2(new_n18744_), .B(new_n12745_), .ZN(new_n18746_));
  AOI21_X1   g16310(.A1(new_n18718_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n18747_));
  INV_X1     g16311(.I(new_n18747_), .ZN(new_n18748_));
  AOI21_X1   g16312(.A1(new_n14163_), .A2(new_n8056_), .B(pi1153), .ZN(new_n18749_));
  OAI21_X1   g16313(.A1(new_n18709_), .A2(pi0625), .B(new_n18749_), .ZN(new_n18750_));
  NAND2_X1   g16314(.A1(new_n18750_), .A2(pi0608), .ZN(new_n18751_));
  AOI21_X1   g16315(.A1(new_n18665_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n18752_));
  OAI21_X1   g16316(.A1(new_n18436_), .A2(new_n18425_), .B(pi0177), .ZN(new_n18753_));
  NAND2_X1   g16317(.A1(new_n14174_), .A2(new_n2627_), .ZN(new_n18754_));
  INV_X1     g16318(.I(new_n15110_), .ZN(new_n18755_));
  NAND3_X1   g16319(.A1(new_n18755_), .A2(new_n8056_), .A3(new_n18754_), .ZN(new_n18756_));
  AOI21_X1   g16320(.A1(new_n18756_), .A2(new_n18753_), .B(pi0038), .ZN(new_n18757_));
  AOI21_X1   g16321(.A1(new_n5336_), .A2(new_n13597_), .B(new_n8056_), .ZN(new_n18758_));
  NOR3_X1    g16322(.A1(new_n13566_), .A2(pi0039), .A3(pi0177), .ZN(new_n18759_));
  OAI21_X1   g16323(.A1(new_n18759_), .A2(new_n18758_), .B(pi0038), .ZN(new_n18760_));
  INV_X1     g16324(.I(new_n18760_), .ZN(new_n18761_));
  NOR3_X1    g16325(.A1(new_n18757_), .A2(pi0757), .A3(new_n18761_), .ZN(new_n18762_));
  AOI21_X1   g16326(.A1(new_n18705_), .A2(new_n14169_), .B(new_n16460_), .ZN(new_n18763_));
  INV_X1     g16327(.I(new_n18763_), .ZN(new_n18764_));
  OR2_X2     g16328(.A1(new_n15119_), .A2(new_n15120_), .Z(new_n18765_));
  AOI21_X1   g16329(.A1(new_n18765_), .A2(pi0177), .B(pi0038), .ZN(new_n18766_));
  NAND3_X1   g16330(.A1(new_n15128_), .A2(new_n15127_), .A3(new_n8056_), .ZN(new_n18767_));
  AOI21_X1   g16331(.A1(new_n18766_), .A2(new_n18767_), .B(new_n18764_), .ZN(new_n18768_));
  OAI21_X1   g16332(.A1(new_n18762_), .A2(new_n18768_), .B(new_n16459_), .ZN(new_n18769_));
  OAI21_X1   g16333(.A1(new_n18663_), .A2(new_n18661_), .B(pi0686), .ZN(new_n18770_));
  NAND3_X1   g16334(.A1(new_n18769_), .A2(new_n2609_), .A3(new_n18770_), .ZN(new_n18771_));
  NAND3_X1   g16335(.A1(new_n18771_), .A2(pi0625), .A3(new_n18698_), .ZN(new_n18772_));
  AOI21_X1   g16336(.A1(new_n18772_), .A2(new_n18752_), .B(new_n18751_), .ZN(new_n18773_));
  AOI21_X1   g16337(.A1(new_n14199_), .A2(new_n8056_), .B(new_n12841_), .ZN(new_n18774_));
  OAI21_X1   g16338(.A1(new_n18709_), .A2(new_n13521_), .B(new_n18774_), .ZN(new_n18775_));
  NAND2_X1   g16339(.A1(new_n18775_), .A2(new_n13560_), .ZN(new_n18776_));
  AOI21_X1   g16340(.A1(new_n18665_), .A2(pi0625), .B(pi1153), .ZN(new_n18777_));
  NAND3_X1   g16341(.A1(new_n18771_), .A2(new_n13521_), .A3(new_n18698_), .ZN(new_n18778_));
  AOI21_X1   g16342(.A1(new_n18778_), .A2(new_n18777_), .B(new_n18776_), .ZN(new_n18779_));
  NOR3_X1    g16343(.A1(new_n18773_), .A2(new_n18779_), .A3(new_n12758_), .ZN(new_n18780_));
  AOI21_X1   g16344(.A1(new_n18771_), .A2(new_n18698_), .B(pi0778), .ZN(new_n18781_));
  OAI21_X1   g16345(.A1(new_n18780_), .A2(new_n18781_), .B(new_n12764_), .ZN(new_n18782_));
  AND2_X2    g16346(.A1(new_n18670_), .A2(pi0660), .Z(new_n18783_));
  OAI21_X1   g16347(.A1(new_n18712_), .A2(pi0609), .B(pi1155), .ZN(new_n18784_));
  NOR3_X1    g16348(.A1(new_n18780_), .A2(new_n12766_), .A3(new_n18781_), .ZN(new_n18785_));
  OAI21_X1   g16349(.A1(new_n18785_), .A2(new_n18784_), .B(new_n18783_), .ZN(new_n18786_));
  NOR2_X1    g16350(.A1(new_n18672_), .A2(pi0660), .ZN(new_n18787_));
  OAI21_X1   g16351(.A1(new_n18712_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n18788_));
  NOR3_X1    g16352(.A1(new_n18780_), .A2(pi0609), .A3(new_n18781_), .ZN(new_n18789_));
  OAI21_X1   g16353(.A1(new_n18789_), .A2(new_n18788_), .B(new_n18787_), .ZN(new_n18790_));
  NAND3_X1   g16354(.A1(new_n18786_), .A2(new_n18790_), .A3(pi0785), .ZN(new_n18791_));
  AOI21_X1   g16355(.A1(new_n18791_), .A2(new_n18782_), .B(pi0781), .ZN(new_n18792_));
  OAI21_X1   g16356(.A1(new_n18676_), .A2(pi1154), .B(pi0627), .ZN(new_n18793_));
  INV_X1     g16357(.I(new_n18714_), .ZN(new_n18794_));
  AOI21_X1   g16358(.A1(new_n18794_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n18795_));
  NAND3_X1   g16359(.A1(new_n18791_), .A2(pi0618), .A3(new_n18782_), .ZN(new_n18796_));
  AOI21_X1   g16360(.A1(new_n18796_), .A2(new_n18795_), .B(new_n18793_), .ZN(new_n18797_));
  OAI21_X1   g16361(.A1(new_n18679_), .A2(new_n12785_), .B(new_n12880_), .ZN(new_n18798_));
  AOI21_X1   g16362(.A1(new_n18794_), .A2(pi0618), .B(pi1154), .ZN(new_n18799_));
  NAND3_X1   g16363(.A1(new_n18791_), .A2(new_n12781_), .A3(new_n18782_), .ZN(new_n18800_));
  AOI21_X1   g16364(.A1(new_n18800_), .A2(new_n18799_), .B(new_n18798_), .ZN(new_n18801_));
  NOR3_X1    g16365(.A1(new_n18797_), .A2(new_n18801_), .A3(new_n12779_), .ZN(new_n18802_));
  OAI21_X1   g16366(.A1(new_n18802_), .A2(new_n18792_), .B(new_n12796_), .ZN(new_n18803_));
  AOI21_X1   g16367(.A1(new_n18684_), .A2(new_n12791_), .B(new_n12895_), .ZN(new_n18804_));
  AOI21_X1   g16368(.A1(new_n18716_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n18805_));
  INV_X1     g16369(.I(new_n18805_), .ZN(new_n18806_));
  NOR3_X1    g16370(.A1(new_n18802_), .A2(new_n12793_), .A3(new_n18792_), .ZN(new_n18807_));
  OAI21_X1   g16371(.A1(new_n18807_), .A2(new_n18806_), .B(new_n18804_), .ZN(new_n18808_));
  AOI21_X1   g16372(.A1(new_n18687_), .A2(pi1159), .B(pi0648), .ZN(new_n18809_));
  NAND2_X1   g16373(.A1(new_n18716_), .A2(pi0619), .ZN(new_n18810_));
  NAND2_X1   g16374(.A1(new_n18810_), .A2(new_n12791_), .ZN(new_n18811_));
  NOR3_X1    g16375(.A1(new_n18802_), .A2(pi0619), .A3(new_n18792_), .ZN(new_n18812_));
  OAI21_X1   g16376(.A1(new_n18812_), .A2(new_n18811_), .B(new_n18809_), .ZN(new_n18813_));
  NAND3_X1   g16377(.A1(new_n18808_), .A2(new_n18813_), .A3(pi0789), .ZN(new_n18814_));
  AOI21_X1   g16378(.A1(new_n18814_), .A2(new_n18803_), .B(new_n12747_), .ZN(new_n18815_));
  OAI21_X1   g16379(.A1(new_n18815_), .A2(new_n18748_), .B(new_n18746_), .ZN(new_n18816_));
  AOI21_X1   g16380(.A1(new_n18655_), .A2(pi0626), .B(new_n12814_), .ZN(new_n18817_));
  NAND3_X1   g16381(.A1(new_n18689_), .A2(new_n12747_), .A3(new_n18682_), .ZN(new_n18818_));
  AOI21_X1   g16382(.A1(new_n18818_), .A2(new_n18817_), .B(pi1158), .ZN(new_n18819_));
  OAI21_X1   g16383(.A1(new_n18719_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n18820_));
  AOI21_X1   g16384(.A1(new_n18814_), .A2(new_n18803_), .B(pi0626), .ZN(new_n18821_));
  OAI21_X1   g16385(.A1(new_n18821_), .A2(new_n18820_), .B(new_n18819_), .ZN(new_n18822_));
  NAND3_X1   g16386(.A1(new_n18816_), .A2(new_n18822_), .A3(pi0788), .ZN(new_n18823_));
  NAND3_X1   g16387(.A1(new_n18814_), .A2(new_n12808_), .A3(new_n18803_), .ZN(new_n18824_));
  AOI21_X1   g16388(.A1(new_n18823_), .A2(new_n18824_), .B(new_n12920_), .ZN(new_n18825_));
  OAI21_X1   g16389(.A1(new_n18825_), .A2(new_n18743_), .B(new_n18742_), .ZN(new_n18826_));
  NOR2_X1    g16390(.A1(new_n18729_), .A2(pi0629), .ZN(new_n18827_));
  OAI21_X1   g16391(.A1(new_n18691_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n18828_));
  AOI21_X1   g16392(.A1(new_n18823_), .A2(new_n18824_), .B(pi0628), .ZN(new_n18829_));
  OAI21_X1   g16393(.A1(new_n18829_), .A2(new_n18828_), .B(new_n18827_), .ZN(new_n18830_));
  NAND3_X1   g16394(.A1(new_n18826_), .A2(new_n18830_), .A3(pi0792), .ZN(new_n18831_));
  NAND3_X1   g16395(.A1(new_n18823_), .A2(new_n12937_), .A3(new_n18824_), .ZN(new_n18832_));
  AOI21_X1   g16396(.A1(new_n18831_), .A2(new_n18832_), .B(pi0787), .ZN(new_n18833_));
  INV_X1     g16397(.I(new_n18833_), .ZN(new_n18834_));
  NAND2_X1   g16398(.A1(new_n18734_), .A2(pi0630), .ZN(new_n18835_));
  AOI21_X1   g16399(.A1(new_n18692_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n18836_));
  NAND3_X1   g16400(.A1(new_n18831_), .A2(pi0647), .A3(new_n18832_), .ZN(new_n18837_));
  AOI21_X1   g16401(.A1(new_n18837_), .A2(new_n18836_), .B(new_n18835_), .ZN(new_n18838_));
  NOR2_X1    g16402(.A1(new_n18737_), .A2(pi0630), .ZN(new_n18839_));
  INV_X1     g16403(.I(new_n18839_), .ZN(new_n18840_));
  AOI21_X1   g16404(.A1(new_n18692_), .A2(pi0647), .B(pi1157), .ZN(new_n18841_));
  NAND3_X1   g16405(.A1(new_n18831_), .A2(new_n12741_), .A3(new_n18832_), .ZN(new_n18842_));
  AOI21_X1   g16406(.A1(new_n18842_), .A2(new_n18841_), .B(new_n18840_), .ZN(new_n18843_));
  NOR3_X1    g16407(.A1(new_n18838_), .A2(new_n18843_), .A3(new_n12972_), .ZN(new_n18844_));
  INV_X1     g16408(.I(new_n18844_), .ZN(new_n18845_));
  NAND3_X1   g16409(.A1(new_n18845_), .A2(new_n12975_), .A3(new_n18834_), .ZN(new_n18846_));
  AOI21_X1   g16410(.A1(new_n18846_), .A2(new_n18741_), .B(new_n18696_), .ZN(new_n18847_));
  OAI21_X1   g16411(.A1(new_n18655_), .A2(pi0644), .B(new_n12740_), .ZN(new_n18848_));
  NOR2_X1    g16412(.A1(new_n18694_), .A2(new_n12975_), .ZN(new_n18849_));
  OAI21_X1   g16413(.A1(new_n18849_), .A2(new_n18848_), .B(pi1160), .ZN(new_n18850_));
  OR2_X2     g16414(.A1(new_n18740_), .A2(pi0644), .Z(new_n18851_));
  OAI21_X1   g16415(.A1(new_n18844_), .A2(new_n18833_), .B(pi0644), .ZN(new_n18852_));
  AOI21_X1   g16416(.A1(new_n18852_), .A2(new_n18851_), .B(new_n12740_), .ZN(new_n18853_));
  OAI21_X1   g16417(.A1(new_n18853_), .A2(new_n18850_), .B(pi0790), .ZN(new_n18854_));
  NAND2_X1   g16418(.A1(new_n18845_), .A2(new_n18834_), .ZN(new_n18855_));
  AOI21_X1   g16419(.A1(new_n18855_), .A2(new_n13000_), .B(po1038), .ZN(new_n18856_));
  OAI21_X1   g16420(.A1(new_n18854_), .A2(new_n18847_), .B(new_n18856_), .ZN(new_n18857_));
  AOI21_X1   g16421(.A1(new_n18857_), .A2(new_n18653_), .B(new_n18652_), .ZN(po0334));
  NOR2_X1    g16422(.A1(new_n13340_), .A2(pi0760), .ZN(new_n18859_));
  NOR2_X1    g16423(.A1(new_n3042_), .A2(pi0178), .ZN(new_n18860_));
  NOR2_X1    g16424(.A1(new_n18859_), .A2(new_n18860_), .ZN(new_n18861_));
  NOR3_X1    g16425(.A1(new_n18861_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n18862_));
  INV_X1     g16426(.I(new_n18859_), .ZN(new_n18863_));
  NOR2_X1    g16427(.A1(new_n18863_), .A2(new_n13354_), .ZN(new_n18864_));
  NOR3_X1    g16428(.A1(new_n18864_), .A2(new_n12762_), .A3(new_n18861_), .ZN(new_n18865_));
  NOR2_X1    g16429(.A1(new_n18865_), .A2(new_n12770_), .ZN(new_n18866_));
  NOR3_X1    g16430(.A1(new_n18864_), .A2(pi1155), .A3(new_n18860_), .ZN(new_n18867_));
  NOR3_X1    g16431(.A1(new_n18866_), .A2(new_n12764_), .A3(new_n18867_), .ZN(new_n18868_));
  NOR2_X1    g16432(.A1(new_n18868_), .A2(new_n18862_), .ZN(new_n18869_));
  INV_X1     g16433(.I(new_n18869_), .ZN(new_n18870_));
  AOI21_X1   g16434(.A1(new_n18870_), .A2(new_n12783_), .B(pi1154), .ZN(new_n18871_));
  AOI21_X1   g16435(.A1(new_n18870_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n18872_));
  NOR3_X1    g16436(.A1(new_n18871_), .A2(new_n18872_), .A3(new_n12779_), .ZN(new_n18873_));
  AOI21_X1   g16437(.A1(new_n12779_), .A2(new_n18870_), .B(new_n18873_), .ZN(new_n18874_));
  OAI21_X1   g16438(.A1(new_n18874_), .A2(new_n17229_), .B(new_n12791_), .ZN(new_n18875_));
  OAI21_X1   g16439(.A1(new_n18874_), .A2(new_n17232_), .B(pi1159), .ZN(new_n18876_));
  NAND3_X1   g16440(.A1(new_n18875_), .A2(new_n18876_), .A3(pi0789), .ZN(new_n18877_));
  OAI21_X1   g16441(.A1(pi0789), .A2(new_n18874_), .B(new_n18877_), .ZN(new_n18878_));
  INV_X1     g16442(.I(new_n18860_), .ZN(new_n18879_));
  NAND2_X1   g16443(.A1(new_n12818_), .A2(new_n18879_), .ZN(new_n18880_));
  OAI21_X1   g16444(.A1(new_n18878_), .A2(new_n12818_), .B(new_n18880_), .ZN(new_n18881_));
  AOI21_X1   g16445(.A1(new_n12826_), .A2(new_n16510_), .B(new_n18860_), .ZN(new_n18882_));
  NOR2_X1    g16446(.A1(new_n18860_), .A2(pi1153), .ZN(new_n18883_));
  NOR2_X1    g16447(.A1(new_n12834_), .A2(pi0688), .ZN(new_n18884_));
  INV_X1     g16448(.I(new_n18884_), .ZN(new_n18885_));
  NAND2_X1   g16449(.A1(new_n18885_), .A2(new_n18883_), .ZN(new_n18886_));
  NOR2_X1    g16450(.A1(new_n18884_), .A2(new_n18882_), .ZN(new_n18887_));
  NOR2_X1    g16451(.A1(new_n18887_), .A2(new_n12841_), .ZN(new_n18888_));
  INV_X1     g16452(.I(new_n18888_), .ZN(new_n18889_));
  NAND3_X1   g16453(.A1(new_n18889_), .A2(pi0778), .A3(new_n18886_), .ZN(new_n18890_));
  OAI21_X1   g16454(.A1(pi0778), .A2(new_n18882_), .B(new_n18890_), .ZN(new_n18891_));
  NAND2_X1   g16455(.A1(new_n18891_), .A2(new_n17187_), .ZN(new_n18892_));
  NOR2_X1    g16456(.A1(new_n18892_), .A2(new_n12889_), .ZN(new_n18893_));
  NAND2_X1   g16457(.A1(new_n18893_), .A2(new_n18203_), .ZN(new_n18894_));
  NOR2_X1    g16458(.A1(new_n18894_), .A2(new_n17884_), .ZN(new_n18895_));
  INV_X1     g16459(.I(new_n18895_), .ZN(new_n18896_));
  OAI22_X1   g16460(.A1(new_n18881_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n18896_), .ZN(new_n18897_));
  AND2_X2    g16461(.A1(new_n18897_), .A2(new_n12919_), .Z(new_n18898_));
  OAI22_X1   g16462(.A1(new_n18881_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n18896_), .ZN(new_n18899_));
  AOI21_X1   g16463(.A1(pi0629), .A2(new_n18899_), .B(new_n18898_), .ZN(new_n18900_));
  INV_X1     g16464(.I(new_n18867_), .ZN(new_n18901_));
  NOR2_X1    g16465(.A1(new_n18882_), .A2(new_n12754_), .ZN(new_n18902_));
  NOR3_X1    g16466(.A1(new_n18902_), .A2(new_n18859_), .A3(new_n18860_), .ZN(new_n18903_));
  NAND2_X1   g16467(.A1(new_n18903_), .A2(new_n12758_), .ZN(new_n18904_));
  NAND2_X1   g16468(.A1(new_n18902_), .A2(pi0625), .ZN(new_n18905_));
  NAND3_X1   g16469(.A1(new_n18905_), .A2(pi1153), .A3(new_n18861_), .ZN(new_n18906_));
  NAND3_X1   g16470(.A1(new_n18886_), .A2(pi0608), .A3(new_n18906_), .ZN(new_n18907_));
  INV_X1     g16471(.I(new_n18905_), .ZN(new_n18908_));
  OAI21_X1   g16472(.A1(new_n18908_), .A2(new_n18903_), .B(new_n18883_), .ZN(new_n18909_));
  NAND3_X1   g16473(.A1(new_n18889_), .A2(new_n13560_), .A3(new_n18909_), .ZN(new_n18910_));
  NAND3_X1   g16474(.A1(new_n18910_), .A2(pi0778), .A3(new_n18907_), .ZN(new_n18911_));
  AOI21_X1   g16475(.A1(new_n18911_), .A2(new_n18904_), .B(new_n12766_), .ZN(new_n18912_));
  NOR2_X1    g16476(.A1(new_n18891_), .A2(pi0609), .ZN(new_n18913_));
  OAI21_X1   g16477(.A1(new_n18913_), .A2(new_n18912_), .B(pi1155), .ZN(new_n18914_));
  NAND3_X1   g16478(.A1(new_n18914_), .A2(pi0660), .A3(new_n18901_), .ZN(new_n18915_));
  NAND2_X1   g16479(.A1(new_n18911_), .A2(new_n18904_), .ZN(new_n18916_));
  NOR2_X1    g16480(.A1(new_n18891_), .A2(new_n12766_), .ZN(new_n18917_));
  AOI21_X1   g16481(.A1(new_n18916_), .A2(new_n12766_), .B(new_n18917_), .ZN(new_n18918_));
  NOR2_X1    g16482(.A1(new_n18866_), .A2(pi0660), .ZN(new_n18919_));
  OAI21_X1   g16483(.A1(new_n18918_), .A2(pi1155), .B(new_n18919_), .ZN(new_n18920_));
  NAND3_X1   g16484(.A1(new_n18920_), .A2(new_n18915_), .A3(pi0785), .ZN(new_n18921_));
  NAND2_X1   g16485(.A1(new_n18916_), .A2(new_n12764_), .ZN(new_n18922_));
  NAND2_X1   g16486(.A1(new_n18921_), .A2(new_n18922_), .ZN(new_n18923_));
  NAND2_X1   g16487(.A1(new_n18923_), .A2(new_n12781_), .ZN(new_n18924_));
  NAND2_X1   g16488(.A1(new_n18892_), .A2(pi0618), .ZN(new_n18925_));
  AOI21_X1   g16489(.A1(new_n18924_), .A2(new_n18925_), .B(pi1154), .ZN(new_n18926_));
  NOR3_X1    g16490(.A1(new_n18926_), .A2(pi0627), .A3(new_n18872_), .ZN(new_n18927_));
  NAND2_X1   g16491(.A1(new_n18892_), .A2(new_n12781_), .ZN(new_n18928_));
  NAND2_X1   g16492(.A1(new_n18923_), .A2(pi0618), .ZN(new_n18929_));
  AOI21_X1   g16493(.A1(new_n18929_), .A2(new_n18928_), .B(new_n12785_), .ZN(new_n18930_));
  NOR3_X1    g16494(.A1(new_n18930_), .A2(new_n12880_), .A3(new_n18871_), .ZN(new_n18931_));
  OR3_X2     g16495(.A1(new_n18927_), .A2(new_n18931_), .A3(new_n12779_), .Z(new_n18932_));
  NAND2_X1   g16496(.A1(new_n18923_), .A2(new_n12779_), .ZN(new_n18933_));
  NAND2_X1   g16497(.A1(new_n18932_), .A2(new_n18933_), .ZN(new_n18934_));
  AOI21_X1   g16498(.A1(new_n18934_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n18935_));
  NOR2_X1    g16499(.A1(new_n18893_), .A2(pi0619), .ZN(new_n18936_));
  AOI21_X1   g16500(.A1(new_n18932_), .A2(new_n18933_), .B(new_n12793_), .ZN(new_n18937_));
  OAI21_X1   g16501(.A1(new_n18937_), .A2(new_n18936_), .B(pi1159), .ZN(new_n18938_));
  NAND3_X1   g16502(.A1(new_n18938_), .A2(pi0648), .A3(new_n18875_), .ZN(new_n18939_));
  NAND2_X1   g16503(.A1(new_n18934_), .A2(new_n12793_), .ZN(new_n18940_));
  OAI21_X1   g16504(.A1(new_n12793_), .A2(new_n18893_), .B(new_n18940_), .ZN(new_n18941_));
  NAND2_X1   g16505(.A1(new_n18941_), .A2(new_n12791_), .ZN(new_n18942_));
  NAND3_X1   g16506(.A1(new_n18942_), .A2(new_n12895_), .A3(new_n18876_), .ZN(new_n18943_));
  NAND3_X1   g16507(.A1(new_n18943_), .A2(pi0789), .A3(new_n18939_), .ZN(new_n18944_));
  NOR2_X1    g16508(.A1(new_n18879_), .A2(new_n12747_), .ZN(new_n18945_));
  AND2_X2    g16509(.A1(new_n18878_), .A2(new_n12747_), .Z(new_n18946_));
  OAI21_X1   g16510(.A1(new_n18946_), .A2(new_n18945_), .B(new_n12815_), .ZN(new_n18947_));
  INV_X1     g16511(.I(new_n18894_), .ZN(new_n18948_));
  NAND2_X1   g16512(.A1(new_n18878_), .A2(pi0626), .ZN(new_n18949_));
  OAI21_X1   g16513(.A1(pi0626), .A2(new_n18879_), .B(new_n18949_), .ZN(new_n18950_));
  AOI22_X1   g16514(.A1(new_n18950_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n18948_), .ZN(new_n18951_));
  NAND2_X1   g16515(.A1(new_n18951_), .A2(new_n18947_), .ZN(new_n18952_));
  AOI22_X1   g16516(.A1(new_n18944_), .A2(new_n18935_), .B1(pi0788), .B2(new_n18952_), .ZN(new_n18953_));
  OAI22_X1   g16517(.A1(new_n18953_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n18900_), .ZN(new_n18954_));
  NAND2_X1   g16518(.A1(new_n18881_), .A2(new_n13384_), .ZN(new_n18955_));
  NAND2_X1   g16519(.A1(new_n12943_), .A2(new_n18879_), .ZN(new_n18956_));
  NAND2_X1   g16520(.A1(new_n18955_), .A2(new_n18956_), .ZN(new_n18957_));
  NOR2_X1    g16521(.A1(new_n18896_), .A2(new_n12953_), .ZN(new_n18958_));
  NOR2_X1    g16522(.A1(new_n18958_), .A2(pi0647), .ZN(new_n18959_));
  NOR2_X1    g16523(.A1(new_n18860_), .A2(new_n12741_), .ZN(new_n18960_));
  OAI21_X1   g16524(.A1(new_n18959_), .A2(new_n18960_), .B(new_n12965_), .ZN(new_n18961_));
  NAND2_X1   g16525(.A1(new_n18958_), .A2(pi0647), .ZN(new_n18962_));
  OAI21_X1   g16526(.A1(pi0647), .A2(new_n18879_), .B(new_n18962_), .ZN(new_n18963_));
  OAI22_X1   g16527(.A1(new_n18963_), .A2(new_n15576_), .B1(new_n18961_), .B2(new_n12981_), .ZN(new_n18964_));
  AOI21_X1   g16528(.A1(new_n18957_), .A2(new_n15608_), .B(new_n18964_), .ZN(new_n18965_));
  OAI22_X1   g16529(.A1(new_n18954_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n18965_), .ZN(new_n18966_));
  NAND2_X1   g16530(.A1(new_n18966_), .A2(new_n13000_), .ZN(new_n18967_));
  AND2_X2    g16531(.A1(new_n18966_), .A2(new_n12975_), .Z(new_n18968_));
  OAI21_X1   g16532(.A1(new_n18963_), .A2(new_n12965_), .B(new_n18961_), .ZN(new_n18969_));
  NAND2_X1   g16533(.A1(new_n18958_), .A2(new_n12972_), .ZN(new_n18970_));
  OAI21_X1   g16534(.A1(new_n18969_), .A2(new_n12972_), .B(new_n18970_), .ZN(new_n18971_));
  NOR2_X1    g16535(.A1(new_n18971_), .A2(new_n12975_), .ZN(new_n18972_));
  OAI21_X1   g16536(.A1(new_n18968_), .A2(new_n18972_), .B(new_n12740_), .ZN(new_n18973_));
  NAND2_X1   g16537(.A1(new_n18879_), .A2(pi0644), .ZN(new_n18974_));
  NOR2_X1    g16538(.A1(new_n17611_), .A2(new_n18860_), .ZN(new_n18975_));
  AOI21_X1   g16539(.A1(new_n18881_), .A2(new_n17611_), .B(new_n18975_), .ZN(new_n18976_));
  OAI21_X1   g16540(.A1(new_n18976_), .A2(pi0644), .B(new_n18974_), .ZN(new_n18977_));
  NAND2_X1   g16541(.A1(new_n18977_), .A2(pi0715), .ZN(new_n18978_));
  NAND3_X1   g16542(.A1(new_n18973_), .A2(new_n12739_), .A3(new_n18978_), .ZN(new_n18979_));
  NOR2_X1    g16543(.A1(new_n18971_), .A2(pi0644), .ZN(new_n18980_));
  AOI21_X1   g16544(.A1(new_n18966_), .A2(pi0644), .B(new_n18980_), .ZN(new_n18981_));
  NAND2_X1   g16545(.A1(new_n18879_), .A2(new_n12975_), .ZN(new_n18982_));
  OAI21_X1   g16546(.A1(new_n18976_), .A2(new_n12975_), .B(new_n18982_), .ZN(new_n18983_));
  AOI21_X1   g16547(.A1(new_n18983_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n18984_));
  OAI21_X1   g16548(.A1(new_n18981_), .A2(new_n12740_), .B(new_n18984_), .ZN(new_n18985_));
  NAND3_X1   g16549(.A1(new_n18979_), .A2(pi0790), .A3(new_n18985_), .ZN(new_n18986_));
  NAND2_X1   g16550(.A1(new_n18986_), .A2(new_n18967_), .ZN(new_n18987_));
  AOI21_X1   g16551(.A1(po1038), .A2(new_n10724_), .B(pi0832), .ZN(new_n18988_));
  NAND2_X1   g16552(.A1(new_n13192_), .A2(new_n10724_), .ZN(new_n18989_));
  INV_X1     g16553(.I(new_n18989_), .ZN(new_n18990_));
  AOI21_X1   g16554(.A1(new_n18990_), .A2(pi0644), .B(new_n12740_), .ZN(new_n18991_));
  NAND2_X1   g16555(.A1(new_n18989_), .A2(new_n12984_), .ZN(new_n18992_));
  NOR2_X1    g16556(.A1(new_n18990_), .A2(new_n13384_), .ZN(new_n18993_));
  NOR2_X1    g16557(.A1(new_n2609_), .A2(new_n10724_), .ZN(new_n18994_));
  NOR2_X1    g16558(.A1(new_n13342_), .A2(pi0760), .ZN(new_n18995_));
  NOR2_X1    g16559(.A1(new_n13344_), .A2(pi0178), .ZN(new_n18996_));
  NOR3_X1    g16560(.A1(new_n18995_), .A2(new_n3265_), .A3(new_n18996_), .ZN(new_n18997_));
  NAND2_X1   g16561(.A1(new_n13334_), .A2(new_n10724_), .ZN(new_n18998_));
  NAND2_X1   g16562(.A1(new_n13245_), .A2(pi0178), .ZN(new_n18999_));
  AOI21_X1   g16563(.A1(new_n18998_), .A2(new_n18999_), .B(pi0760), .ZN(new_n19000_));
  NOR3_X1    g16564(.A1(new_n15787_), .A2(pi0178), .A3(new_n16512_), .ZN(new_n19001_));
  NOR2_X1    g16565(.A1(new_n19000_), .A2(new_n19001_), .ZN(new_n19002_));
  AOI21_X1   g16566(.A1(new_n19002_), .A2(new_n3265_), .B(new_n18997_), .ZN(new_n19003_));
  NOR2_X1    g16567(.A1(new_n19003_), .A2(new_n2610_), .ZN(new_n19004_));
  NOR2_X1    g16568(.A1(new_n19004_), .A2(new_n18994_), .ZN(new_n19005_));
  NOR2_X1    g16569(.A1(new_n19005_), .A2(new_n12760_), .ZN(new_n19006_));
  INV_X1     g16570(.I(new_n19006_), .ZN(new_n19007_));
  OAI21_X1   g16571(.A1(new_n12761_), .A2(new_n18990_), .B(new_n19007_), .ZN(new_n19008_));
  OAI22_X1   g16572(.A1(new_n19007_), .A2(pi0609), .B1(new_n13353_), .B2(new_n18990_), .ZN(new_n19009_));
  NAND2_X1   g16573(.A1(new_n19009_), .A2(new_n12770_), .ZN(new_n19010_));
  INV_X1     g16574(.I(new_n19010_), .ZN(new_n19011_));
  AOI22_X1   g16575(.A1(new_n19006_), .A2(pi0609), .B1(new_n13357_), .B2(new_n18989_), .ZN(new_n19012_));
  OAI21_X1   g16576(.A1(new_n19012_), .A2(new_n12770_), .B(pi0785), .ZN(new_n19013_));
  OAI22_X1   g16577(.A1(new_n19011_), .A2(new_n19013_), .B1(pi0785), .B2(new_n19008_), .ZN(new_n19014_));
  NAND2_X1   g16578(.A1(new_n19014_), .A2(new_n12779_), .ZN(new_n19015_));
  NAND2_X1   g16579(.A1(new_n18989_), .A2(pi0618), .ZN(new_n19016_));
  OAI21_X1   g16580(.A1(new_n19014_), .A2(pi0618), .B(new_n19016_), .ZN(new_n19017_));
  NAND2_X1   g16581(.A1(new_n19017_), .A2(new_n12785_), .ZN(new_n19018_));
  NAND2_X1   g16582(.A1(new_n18989_), .A2(new_n12781_), .ZN(new_n19019_));
  OAI21_X1   g16583(.A1(new_n19014_), .A2(new_n12781_), .B(new_n19019_), .ZN(new_n19020_));
  NAND2_X1   g16584(.A1(new_n19020_), .A2(pi1154), .ZN(new_n19021_));
  NAND3_X1   g16585(.A1(new_n19018_), .A2(new_n19021_), .A3(pi0781), .ZN(new_n19022_));
  NAND2_X1   g16586(.A1(new_n19022_), .A2(new_n19015_), .ZN(new_n19023_));
  NAND2_X1   g16587(.A1(new_n19023_), .A2(new_n12796_), .ZN(new_n19024_));
  NAND2_X1   g16588(.A1(new_n18989_), .A2(pi0619), .ZN(new_n19025_));
  OAI21_X1   g16589(.A1(new_n19023_), .A2(pi0619), .B(new_n19025_), .ZN(new_n19026_));
  NAND2_X1   g16590(.A1(new_n19026_), .A2(new_n12791_), .ZN(new_n19027_));
  NAND2_X1   g16591(.A1(new_n18989_), .A2(new_n12793_), .ZN(new_n19028_));
  OAI21_X1   g16592(.A1(new_n19023_), .A2(new_n12793_), .B(new_n19028_), .ZN(new_n19029_));
  NAND2_X1   g16593(.A1(new_n19029_), .A2(pi1159), .ZN(new_n19030_));
  NAND3_X1   g16594(.A1(new_n19027_), .A2(new_n19030_), .A3(pi0789), .ZN(new_n19031_));
  NAND2_X1   g16595(.A1(new_n19031_), .A2(new_n19024_), .ZN(new_n19032_));
  NAND2_X1   g16596(.A1(new_n18989_), .A2(new_n12818_), .ZN(new_n19033_));
  OAI21_X1   g16597(.A1(new_n19032_), .A2(new_n12818_), .B(new_n19033_), .ZN(new_n19034_));
  AOI21_X1   g16598(.A1(new_n19034_), .A2(new_n13384_), .B(new_n18993_), .ZN(new_n19035_));
  OAI21_X1   g16599(.A1(new_n19035_), .A2(new_n12984_), .B(new_n18992_), .ZN(new_n19036_));
  OAI21_X1   g16600(.A1(new_n19036_), .A2(pi0644), .B(new_n18991_), .ZN(new_n19037_));
  AND2_X2    g16601(.A1(new_n19037_), .A2(new_n12739_), .Z(new_n19038_));
  OAI21_X1   g16602(.A1(new_n14125_), .A2(new_n18996_), .B(new_n16510_), .ZN(new_n19039_));
  OAI21_X1   g16603(.A1(new_n14122_), .A2(new_n10724_), .B(new_n3265_), .ZN(new_n19040_));
  NAND2_X1   g16604(.A1(new_n19040_), .A2(new_n2609_), .ZN(new_n19041_));
  NAND2_X1   g16605(.A1(new_n15744_), .A2(new_n10724_), .ZN(new_n19042_));
  AOI21_X1   g16606(.A1(new_n19042_), .A2(new_n19041_), .B(new_n19039_), .ZN(new_n19043_));
  NAND2_X1   g16607(.A1(new_n2609_), .A2(new_n16510_), .ZN(new_n19044_));
  AOI21_X1   g16608(.A1(new_n18990_), .A2(new_n19044_), .B(new_n19043_), .ZN(new_n19045_));
  NAND2_X1   g16609(.A1(new_n19045_), .A2(new_n13521_), .ZN(new_n19046_));
  NAND2_X1   g16610(.A1(new_n18989_), .A2(pi0625), .ZN(new_n19047_));
  AOI21_X1   g16611(.A1(new_n19046_), .A2(new_n19047_), .B(pi1153), .ZN(new_n19048_));
  NAND2_X1   g16612(.A1(new_n18989_), .A2(new_n13521_), .ZN(new_n19049_));
  NAND2_X1   g16613(.A1(new_n19045_), .A2(pi0625), .ZN(new_n19050_));
  AOI21_X1   g16614(.A1(new_n19050_), .A2(new_n19049_), .B(new_n12841_), .ZN(new_n19051_));
  NOR3_X1    g16615(.A1(new_n19048_), .A2(new_n19051_), .A3(new_n12758_), .ZN(new_n19052_));
  NOR2_X1    g16616(.A1(new_n19045_), .A2(pi0778), .ZN(new_n19053_));
  NOR2_X1    g16617(.A1(new_n19052_), .A2(new_n19053_), .ZN(new_n19054_));
  NOR2_X1    g16618(.A1(new_n19054_), .A2(new_n12869_), .ZN(new_n19055_));
  AOI21_X1   g16619(.A1(new_n12869_), .A2(new_n18990_), .B(new_n19055_), .ZN(new_n19056_));
  NAND2_X1   g16620(.A1(new_n19056_), .A2(new_n12888_), .ZN(new_n19057_));
  OAI21_X1   g16621(.A1(new_n12888_), .A2(new_n18990_), .B(new_n19057_), .ZN(new_n19058_));
  INV_X1     g16622(.I(new_n19058_), .ZN(new_n19059_));
  NOR2_X1    g16623(.A1(new_n18989_), .A2(new_n12911_), .ZN(new_n19060_));
  AOI21_X1   g16624(.A1(new_n19059_), .A2(new_n12911_), .B(new_n19060_), .ZN(new_n19061_));
  NAND2_X1   g16625(.A1(new_n19061_), .A2(new_n13392_), .ZN(new_n19062_));
  OAI21_X1   g16626(.A1(new_n13392_), .A2(new_n18990_), .B(new_n19062_), .ZN(new_n19063_));
  NAND2_X1   g16627(.A1(new_n19063_), .A2(new_n12920_), .ZN(new_n19064_));
  NAND2_X1   g16628(.A1(new_n18989_), .A2(pi0628), .ZN(new_n19065_));
  AOI21_X1   g16629(.A1(new_n19064_), .A2(new_n19065_), .B(pi1156), .ZN(new_n19066_));
  NAND2_X1   g16630(.A1(new_n18989_), .A2(new_n12920_), .ZN(new_n19067_));
  NAND2_X1   g16631(.A1(new_n19063_), .A2(pi0628), .ZN(new_n19068_));
  AOI21_X1   g16632(.A1(new_n19068_), .A2(new_n19067_), .B(new_n12742_), .ZN(new_n19069_));
  OR2_X2     g16633(.A1(new_n19069_), .A2(new_n12937_), .Z(new_n19070_));
  OAI22_X1   g16634(.A1(new_n19070_), .A2(new_n19066_), .B1(pi0792), .B2(new_n19063_), .ZN(new_n19071_));
  NAND2_X1   g16635(.A1(new_n19071_), .A2(new_n12741_), .ZN(new_n19072_));
  OAI21_X1   g16636(.A1(new_n12741_), .A2(new_n18989_), .B(new_n19072_), .ZN(new_n19073_));
  NOR2_X1    g16637(.A1(new_n19073_), .A2(pi1157), .ZN(new_n19074_));
  NAND2_X1   g16638(.A1(new_n19071_), .A2(pi0647), .ZN(new_n19075_));
  OAI21_X1   g16639(.A1(pi0647), .A2(new_n18989_), .B(new_n19075_), .ZN(new_n19076_));
  NOR2_X1    g16640(.A1(new_n19076_), .A2(new_n12965_), .ZN(new_n19077_));
  OAI21_X1   g16641(.A1(new_n19074_), .A2(new_n19077_), .B(pi0787), .ZN(new_n19078_));
  OAI21_X1   g16642(.A1(pi0787), .A2(new_n19071_), .B(new_n19078_), .ZN(new_n19079_));
  OAI21_X1   g16643(.A1(new_n19079_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n19080_));
  AOI21_X1   g16644(.A1(new_n18990_), .A2(new_n12975_), .B(pi0715), .ZN(new_n19081_));
  OAI21_X1   g16645(.A1(new_n19036_), .A2(new_n12975_), .B(new_n19081_), .ZN(new_n19082_));
  AND2_X2    g16646(.A1(new_n19082_), .A2(pi1160), .Z(new_n19083_));
  OAI21_X1   g16647(.A1(new_n19079_), .A2(pi0644), .B(pi0715), .ZN(new_n19084_));
  AOI22_X1   g16648(.A1(new_n19038_), .A2(new_n19080_), .B1(new_n19084_), .B2(new_n19083_), .ZN(new_n19085_));
  NOR2_X1    g16649(.A1(new_n19085_), .A2(new_n13000_), .ZN(new_n19086_));
  NAND2_X1   g16650(.A1(new_n18990_), .A2(pi0626), .ZN(new_n19087_));
  NAND2_X1   g16651(.A1(new_n19032_), .A2(new_n12747_), .ZN(new_n19088_));
  AOI21_X1   g16652(.A1(new_n19088_), .A2(new_n19087_), .B(new_n12816_), .ZN(new_n19089_));
  NOR2_X1    g16653(.A1(new_n18989_), .A2(pi0626), .ZN(new_n19090_));
  AOI21_X1   g16654(.A1(new_n19032_), .A2(pi0626), .B(new_n19090_), .ZN(new_n19091_));
  OAI22_X1   g16655(.A1(new_n19091_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n19061_), .ZN(new_n19092_));
  OAI21_X1   g16656(.A1(new_n19092_), .A2(new_n19089_), .B(pi0788), .ZN(new_n19093_));
  NAND2_X1   g16657(.A1(new_n19093_), .A2(new_n15824_), .ZN(new_n19094_));
  NAND2_X1   g16658(.A1(new_n19054_), .A2(new_n12766_), .ZN(new_n19095_));
  AOI21_X1   g16659(.A1(new_n16512_), .A2(new_n13566_), .B(new_n15826_), .ZN(new_n19096_));
  AOI21_X1   g16660(.A1(new_n14328_), .A2(new_n18863_), .B(new_n10724_), .ZN(new_n19097_));
  AOI21_X1   g16661(.A1(new_n19097_), .A2(new_n5336_), .B(new_n3265_), .ZN(new_n19098_));
  OAI21_X1   g16662(.A1(new_n19096_), .A2(pi0178), .B(new_n19098_), .ZN(new_n19099_));
  NAND2_X1   g16663(.A1(new_n14172_), .A2(pi0178), .ZN(new_n19100_));
  NAND2_X1   g16664(.A1(new_n14174_), .A2(new_n10724_), .ZN(new_n19101_));
  AOI21_X1   g16665(.A1(new_n19100_), .A2(new_n19101_), .B(pi0760), .ZN(new_n19102_));
  NAND2_X1   g16666(.A1(new_n15835_), .A2(pi0178), .ZN(new_n19103_));
  NAND2_X1   g16667(.A1(new_n14177_), .A2(new_n10724_), .ZN(new_n19104_));
  AOI21_X1   g16668(.A1(new_n19104_), .A2(new_n19103_), .B(new_n16512_), .ZN(new_n19105_));
  OAI21_X1   g16669(.A1(new_n19105_), .A2(new_n19102_), .B(new_n2627_), .ZN(new_n19106_));
  NOR2_X1    g16670(.A1(new_n14182_), .A2(pi0178), .ZN(new_n19107_));
  NOR2_X1    g16671(.A1(new_n14184_), .A2(new_n10724_), .ZN(new_n19108_));
  OAI21_X1   g16672(.A1(new_n19107_), .A2(new_n19108_), .B(pi0760), .ZN(new_n19109_));
  NOR2_X1    g16673(.A1(new_n14187_), .A2(new_n10724_), .ZN(new_n19110_));
  NOR2_X1    g16674(.A1(new_n14189_), .A2(pi0178), .ZN(new_n19111_));
  OAI21_X1   g16675(.A1(new_n19110_), .A2(new_n19111_), .B(new_n16512_), .ZN(new_n19112_));
  NAND3_X1   g16676(.A1(new_n19112_), .A2(new_n19109_), .A3(pi0039), .ZN(new_n19113_));
  NAND3_X1   g16677(.A1(new_n19113_), .A2(new_n3265_), .A3(new_n19106_), .ZN(new_n19114_));
  NAND3_X1   g16678(.A1(new_n19114_), .A2(new_n16510_), .A3(new_n19099_), .ZN(new_n19115_));
  NAND2_X1   g16679(.A1(new_n19003_), .A2(pi0688), .ZN(new_n19116_));
  NAND3_X1   g16680(.A1(new_n19115_), .A2(new_n2609_), .A3(new_n19116_), .ZN(new_n19117_));
  OAI21_X1   g16681(.A1(new_n10724_), .A2(new_n2609_), .B(new_n19117_), .ZN(new_n19118_));
  INV_X1     g16682(.I(new_n19051_), .ZN(new_n19119_));
  NOR2_X1    g16683(.A1(new_n19005_), .A2(new_n13521_), .ZN(new_n19120_));
  AOI21_X1   g16684(.A1(new_n19118_), .A2(new_n13521_), .B(new_n19120_), .ZN(new_n19121_));
  OAI21_X1   g16685(.A1(new_n19121_), .A2(pi1153), .B(new_n19119_), .ZN(new_n19122_));
  NOR2_X1    g16686(.A1(new_n19005_), .A2(pi0625), .ZN(new_n19123_));
  AOI21_X1   g16687(.A1(new_n19118_), .A2(pi0625), .B(new_n19123_), .ZN(new_n19124_));
  OAI21_X1   g16688(.A1(new_n19124_), .A2(new_n12841_), .B(pi0608), .ZN(new_n19125_));
  OAI22_X1   g16689(.A1(pi0608), .A2(new_n19122_), .B1(new_n19125_), .B2(new_n19048_), .ZN(new_n19126_));
  NOR2_X1    g16690(.A1(new_n19126_), .A2(new_n12758_), .ZN(new_n19127_));
  AOI21_X1   g16691(.A1(new_n12758_), .A2(new_n19118_), .B(new_n19127_), .ZN(new_n19128_));
  OAI21_X1   g16692(.A1(new_n19128_), .A2(new_n12766_), .B(new_n19095_), .ZN(new_n19129_));
  AOI21_X1   g16693(.A1(new_n19129_), .A2(pi1155), .B(new_n19011_), .ZN(new_n19130_));
  NOR2_X1    g16694(.A1(new_n19128_), .A2(pi0609), .ZN(new_n19131_));
  NOR3_X1    g16695(.A1(new_n19052_), .A2(new_n12766_), .A3(new_n19053_), .ZN(new_n19132_));
  OAI21_X1   g16696(.A1(new_n19131_), .A2(new_n19132_), .B(new_n12770_), .ZN(new_n19133_));
  NOR2_X1    g16697(.A1(new_n19012_), .A2(new_n12770_), .ZN(new_n19134_));
  NOR2_X1    g16698(.A1(new_n19134_), .A2(pi0660), .ZN(new_n19135_));
  AOI22_X1   g16699(.A1(new_n19130_), .A2(pi0660), .B1(new_n19133_), .B2(new_n19135_), .ZN(new_n19136_));
  NOR2_X1    g16700(.A1(new_n19128_), .A2(pi0785), .ZN(new_n19137_));
  AOI21_X1   g16701(.A1(new_n19136_), .A2(pi0785), .B(new_n19137_), .ZN(new_n19138_));
  NOR2_X1    g16702(.A1(new_n19138_), .A2(pi0781), .ZN(new_n19139_));
  AND2_X2    g16703(.A1(new_n19056_), .A2(new_n12781_), .Z(new_n19140_));
  NOR2_X1    g16704(.A1(new_n19138_), .A2(new_n12781_), .ZN(new_n19141_));
  OAI21_X1   g16705(.A1(new_n19141_), .A2(new_n19140_), .B(pi1154), .ZN(new_n19142_));
  NAND3_X1   g16706(.A1(new_n19142_), .A2(pi0627), .A3(new_n19018_), .ZN(new_n19143_));
  INV_X1     g16707(.I(new_n19021_), .ZN(new_n19144_));
  NAND2_X1   g16708(.A1(new_n19056_), .A2(pi0618), .ZN(new_n19145_));
  OAI21_X1   g16709(.A1(new_n19138_), .A2(pi0618), .B(new_n19145_), .ZN(new_n19146_));
  AOI21_X1   g16710(.A1(new_n19146_), .A2(new_n12785_), .B(new_n19144_), .ZN(new_n19147_));
  AOI21_X1   g16711(.A1(new_n19147_), .A2(new_n12880_), .B(new_n12779_), .ZN(new_n19148_));
  AOI21_X1   g16712(.A1(new_n19148_), .A2(new_n19143_), .B(new_n19139_), .ZN(new_n19149_));
  OAI21_X1   g16713(.A1(new_n19149_), .A2(pi0789), .B(new_n12819_), .ZN(new_n19150_));
  NOR2_X1    g16714(.A1(new_n19059_), .A2(new_n12793_), .ZN(new_n19151_));
  NOR2_X1    g16715(.A1(new_n19149_), .A2(pi0619), .ZN(new_n19152_));
  OAI21_X1   g16716(.A1(new_n19152_), .A2(new_n19151_), .B(new_n12791_), .ZN(new_n19153_));
  NAND3_X1   g16717(.A1(new_n19153_), .A2(new_n12895_), .A3(new_n19030_), .ZN(new_n19154_));
  NAND2_X1   g16718(.A1(new_n19058_), .A2(new_n12793_), .ZN(new_n19155_));
  OAI21_X1   g16719(.A1(new_n19149_), .A2(new_n12793_), .B(new_n19155_), .ZN(new_n19156_));
  AOI21_X1   g16720(.A1(new_n19156_), .A2(pi1159), .B(new_n12895_), .ZN(new_n19157_));
  AOI21_X1   g16721(.A1(new_n19157_), .A2(new_n19027_), .B(new_n12796_), .ZN(new_n19158_));
  AOI21_X1   g16722(.A1(new_n19158_), .A2(new_n19154_), .B(new_n19150_), .ZN(new_n19159_));
  INV_X1     g16723(.I(new_n15821_), .ZN(new_n19160_));
  NOR2_X1    g16724(.A1(new_n19069_), .A2(pi0629), .ZN(new_n19161_));
  NOR2_X1    g16725(.A1(new_n19066_), .A2(new_n12919_), .ZN(new_n19162_));
  NOR2_X1    g16726(.A1(new_n19161_), .A2(new_n19162_), .ZN(new_n19163_));
  AOI21_X1   g16727(.A1(new_n19034_), .A2(new_n19160_), .B(new_n19163_), .ZN(new_n19164_));
  OAI22_X1   g16728(.A1(new_n19159_), .A2(new_n19094_), .B1(new_n12937_), .B2(new_n19164_), .ZN(new_n19165_));
  NOR2_X1    g16729(.A1(new_n19083_), .A2(new_n12975_), .ZN(new_n19166_));
  NOR2_X1    g16730(.A1(new_n19038_), .A2(pi0644), .ZN(new_n19167_));
  NOR2_X1    g16731(.A1(new_n19166_), .A2(new_n19167_), .ZN(new_n19168_));
  OAI22_X1   g16732(.A1(new_n15576_), .A2(new_n19076_), .B1(new_n19073_), .B2(new_n15730_), .ZN(new_n19169_));
  NOR2_X1    g16733(.A1(new_n19035_), .A2(new_n17212_), .ZN(new_n19170_));
  NOR2_X1    g16734(.A1(new_n19169_), .A2(new_n19170_), .ZN(new_n19171_));
  OAI22_X1   g16735(.A1(new_n19168_), .A2(new_n13000_), .B1(new_n19171_), .B2(new_n12972_), .ZN(new_n19172_));
  AOI21_X1   g16736(.A1(new_n15693_), .A2(new_n19165_), .B(new_n19172_), .ZN(new_n19173_));
  OAI21_X1   g16737(.A1(new_n19086_), .A2(new_n19173_), .B(new_n6643_), .ZN(new_n19174_));
  AOI22_X1   g16738(.A1(new_n19174_), .A2(new_n18988_), .B1(pi0832), .B2(new_n18987_), .ZN(po0335));
  NOR2_X1    g16739(.A1(new_n3042_), .A2(pi0179), .ZN(new_n19176_));
  INV_X1     g16740(.I(new_n19176_), .ZN(new_n19177_));
  AOI21_X1   g16741(.A1(new_n12756_), .A2(new_n16500_), .B(new_n19176_), .ZN(new_n19178_));
  NOR3_X1    g16742(.A1(new_n19178_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n19179_));
  NOR2_X1    g16743(.A1(new_n19178_), .A2(new_n12762_), .ZN(new_n19180_));
  AOI21_X1   g16744(.A1(new_n19180_), .A2(new_n12768_), .B(pi1155), .ZN(new_n19181_));
  INV_X1     g16745(.I(new_n19178_), .ZN(new_n19182_));
  AOI21_X1   g16746(.A1(new_n19182_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n19183_));
  NOR3_X1    g16747(.A1(new_n19181_), .A2(new_n19183_), .A3(new_n12764_), .ZN(new_n19184_));
  NOR2_X1    g16748(.A1(new_n19184_), .A2(new_n19179_), .ZN(new_n19185_));
  NOR2_X1    g16749(.A1(new_n19185_), .A2(pi0781), .ZN(new_n19186_));
  INV_X1     g16750(.I(new_n19185_), .ZN(new_n19187_));
  AOI21_X1   g16751(.A1(new_n19187_), .A2(new_n12783_), .B(pi1154), .ZN(new_n19188_));
  AOI21_X1   g16752(.A1(new_n19187_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n19189_));
  NOR3_X1    g16753(.A1(new_n19188_), .A2(new_n19189_), .A3(new_n12779_), .ZN(new_n19190_));
  NOR2_X1    g16754(.A1(new_n19190_), .A2(new_n19186_), .ZN(new_n19191_));
  NOR3_X1    g16755(.A1(new_n19190_), .A2(pi0619), .A3(new_n19186_), .ZN(new_n19192_));
  NOR2_X1    g16756(.A1(new_n19176_), .A2(new_n12793_), .ZN(new_n19193_));
  OAI21_X1   g16757(.A1(new_n19192_), .A2(new_n19193_), .B(new_n12791_), .ZN(new_n19194_));
  NAND2_X1   g16758(.A1(new_n19191_), .A2(pi0619), .ZN(new_n19195_));
  NAND2_X1   g16759(.A1(new_n19177_), .A2(new_n12793_), .ZN(new_n19196_));
  AOI21_X1   g16760(.A1(new_n19195_), .A2(new_n19196_), .B(new_n12791_), .ZN(new_n19197_));
  INV_X1     g16761(.I(new_n19197_), .ZN(new_n19198_));
  NAND3_X1   g16762(.A1(new_n19198_), .A2(pi0789), .A3(new_n19194_), .ZN(new_n19199_));
  OAI21_X1   g16763(.A1(pi0789), .A2(new_n19191_), .B(new_n19199_), .ZN(new_n19200_));
  NOR2_X1    g16764(.A1(new_n19200_), .A2(new_n12818_), .ZN(new_n19201_));
  AOI21_X1   g16765(.A1(new_n12818_), .A2(new_n19177_), .B(new_n19201_), .ZN(new_n19202_));
  AOI21_X1   g16766(.A1(new_n12826_), .A2(new_n16499_), .B(new_n19176_), .ZN(new_n19203_));
  NOR2_X1    g16767(.A1(new_n19203_), .A2(pi0778), .ZN(new_n19204_));
  NOR2_X1    g16768(.A1(new_n19176_), .A2(pi1153), .ZN(new_n19205_));
  NOR2_X1    g16769(.A1(new_n12834_), .A2(pi0724), .ZN(new_n19206_));
  INV_X1     g16770(.I(new_n19206_), .ZN(new_n19207_));
  NAND2_X1   g16771(.A1(new_n19207_), .A2(new_n19205_), .ZN(new_n19208_));
  INV_X1     g16772(.I(new_n19208_), .ZN(new_n19209_));
  NOR2_X1    g16773(.A1(new_n19206_), .A2(new_n19203_), .ZN(new_n19210_));
  NOR2_X1    g16774(.A1(new_n19210_), .A2(new_n12841_), .ZN(new_n19211_));
  NOR2_X1    g16775(.A1(new_n19209_), .A2(new_n19211_), .ZN(new_n19212_));
  AOI21_X1   g16776(.A1(new_n19212_), .A2(pi0778), .B(new_n19204_), .ZN(new_n19213_));
  NOR2_X1    g16777(.A1(new_n19213_), .A2(new_n12871_), .ZN(new_n19214_));
  INV_X1     g16778(.I(new_n19214_), .ZN(new_n19215_));
  NOR2_X1    g16779(.A1(new_n19215_), .A2(new_n12889_), .ZN(new_n19216_));
  NAND2_X1   g16780(.A1(new_n19216_), .A2(new_n18203_), .ZN(new_n19217_));
  NOR2_X1    g16781(.A1(new_n19217_), .A2(new_n17884_), .ZN(new_n19218_));
  AOI22_X1   g16782(.A1(new_n19202_), .A2(new_n12949_), .B1(new_n15695_), .B2(new_n19218_), .ZN(new_n19219_));
  NOR2_X1    g16783(.A1(new_n19219_), .A2(pi0629), .ZN(new_n19220_));
  AOI22_X1   g16784(.A1(new_n19202_), .A2(new_n12948_), .B1(new_n15700_), .B2(new_n19218_), .ZN(new_n19221_));
  NOR2_X1    g16785(.A1(new_n19221_), .A2(new_n12919_), .ZN(new_n19222_));
  NOR2_X1    g16786(.A1(new_n19220_), .A2(new_n19222_), .ZN(new_n19223_));
  NOR2_X1    g16787(.A1(new_n19203_), .A2(new_n12754_), .ZN(new_n19224_));
  NOR2_X1    g16788(.A1(new_n19224_), .A2(new_n19182_), .ZN(new_n19225_));
  NAND2_X1   g16789(.A1(new_n19225_), .A2(new_n12758_), .ZN(new_n19226_));
  NAND2_X1   g16790(.A1(new_n19224_), .A2(pi0625), .ZN(new_n19227_));
  NAND3_X1   g16791(.A1(new_n19227_), .A2(pi1153), .A3(new_n19178_), .ZN(new_n19228_));
  AND3_X2    g16792(.A1(new_n19208_), .A2(pi0608), .A3(new_n19228_), .Z(new_n19229_));
  NOR2_X1    g16793(.A1(new_n19211_), .A2(pi0608), .ZN(new_n19230_));
  INV_X1     g16794(.I(new_n19227_), .ZN(new_n19231_));
  OAI21_X1   g16795(.A1(new_n19231_), .A2(new_n19225_), .B(new_n19205_), .ZN(new_n19232_));
  NAND2_X1   g16796(.A1(new_n19230_), .A2(new_n19232_), .ZN(new_n19233_));
  NAND2_X1   g16797(.A1(new_n19233_), .A2(pi0778), .ZN(new_n19234_));
  OAI21_X1   g16798(.A1(new_n19234_), .A2(new_n19229_), .B(new_n19226_), .ZN(new_n19235_));
  INV_X1     g16799(.I(new_n19235_), .ZN(new_n19236_));
  NAND2_X1   g16800(.A1(new_n19213_), .A2(new_n12766_), .ZN(new_n19237_));
  OAI21_X1   g16801(.A1(new_n19236_), .A2(new_n12766_), .B(new_n19237_), .ZN(new_n19238_));
  AOI21_X1   g16802(.A1(new_n19238_), .A2(pi1155), .B(new_n19181_), .ZN(new_n19239_));
  NAND2_X1   g16803(.A1(new_n19235_), .A2(new_n12766_), .ZN(new_n19240_));
  NAND2_X1   g16804(.A1(new_n19213_), .A2(pi0609), .ZN(new_n19241_));
  AOI21_X1   g16805(.A1(new_n19240_), .A2(new_n19241_), .B(pi1155), .ZN(new_n19242_));
  NOR3_X1    g16806(.A1(new_n19242_), .A2(pi0660), .A3(new_n19183_), .ZN(new_n19243_));
  AOI21_X1   g16807(.A1(pi0660), .A2(new_n19239_), .B(new_n19243_), .ZN(new_n19244_));
  NAND2_X1   g16808(.A1(new_n19244_), .A2(pi0785), .ZN(new_n19245_));
  OAI21_X1   g16809(.A1(pi0785), .A2(new_n19236_), .B(new_n19245_), .ZN(new_n19246_));
  INV_X1     g16810(.I(new_n19246_), .ZN(new_n19247_));
  NAND2_X1   g16811(.A1(new_n19215_), .A2(pi0618), .ZN(new_n19248_));
  OAI21_X1   g16812(.A1(new_n19247_), .A2(pi0618), .B(new_n19248_), .ZN(new_n19249_));
  AOI21_X1   g16813(.A1(new_n19249_), .A2(new_n12785_), .B(new_n19189_), .ZN(new_n19250_));
  NOR2_X1    g16814(.A1(new_n19214_), .A2(pi0618), .ZN(new_n19251_));
  NOR2_X1    g16815(.A1(new_n19247_), .A2(new_n12781_), .ZN(new_n19252_));
  OAI21_X1   g16816(.A1(new_n19252_), .A2(new_n19251_), .B(pi1154), .ZN(new_n19253_));
  NOR2_X1    g16817(.A1(new_n19188_), .A2(new_n12880_), .ZN(new_n19254_));
  AOI22_X1   g16818(.A1(new_n19250_), .A2(new_n12880_), .B1(new_n19253_), .B2(new_n19254_), .ZN(new_n19255_));
  NAND2_X1   g16819(.A1(new_n19255_), .A2(pi0781), .ZN(new_n19256_));
  NAND2_X1   g16820(.A1(new_n19246_), .A2(new_n12779_), .ZN(new_n19257_));
  NAND2_X1   g16821(.A1(new_n19256_), .A2(new_n19257_), .ZN(new_n19258_));
  AOI21_X1   g16822(.A1(new_n19258_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n19259_));
  NOR2_X1    g16823(.A1(new_n19216_), .A2(pi0619), .ZN(new_n19260_));
  INV_X1     g16824(.I(new_n19258_), .ZN(new_n19261_));
  NOR2_X1    g16825(.A1(new_n19261_), .A2(new_n12793_), .ZN(new_n19262_));
  OAI21_X1   g16826(.A1(new_n19262_), .A2(new_n19260_), .B(pi1159), .ZN(new_n19263_));
  NAND3_X1   g16827(.A1(new_n19263_), .A2(pi0648), .A3(new_n19194_), .ZN(new_n19264_));
  NOR2_X1    g16828(.A1(new_n19261_), .A2(pi0619), .ZN(new_n19265_));
  NOR2_X1    g16829(.A1(new_n19216_), .A2(new_n12793_), .ZN(new_n19266_));
  OAI21_X1   g16830(.A1(new_n19265_), .A2(new_n19266_), .B(new_n12791_), .ZN(new_n19267_));
  NAND3_X1   g16831(.A1(new_n19267_), .A2(new_n12895_), .A3(new_n19198_), .ZN(new_n19268_));
  NAND3_X1   g16832(.A1(new_n19264_), .A2(new_n19268_), .A3(pi0789), .ZN(new_n19269_));
  NOR2_X1    g16833(.A1(new_n19177_), .A2(new_n12747_), .ZN(new_n19270_));
  INV_X1     g16834(.I(new_n19200_), .ZN(new_n19271_));
  NOR2_X1    g16835(.A1(new_n19271_), .A2(pi0626), .ZN(new_n19272_));
  OAI21_X1   g16836(.A1(new_n19272_), .A2(new_n19270_), .B(new_n12815_), .ZN(new_n19273_));
  INV_X1     g16837(.I(new_n19217_), .ZN(new_n19274_));
  NAND2_X1   g16838(.A1(new_n19176_), .A2(new_n12747_), .ZN(new_n19275_));
  OAI21_X1   g16839(.A1(new_n19271_), .A2(new_n12747_), .B(new_n19275_), .ZN(new_n19276_));
  AOI22_X1   g16840(.A1(new_n19276_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n19274_), .ZN(new_n19277_));
  NAND2_X1   g16841(.A1(new_n19277_), .A2(new_n19273_), .ZN(new_n19278_));
  AOI22_X1   g16842(.A1(new_n19269_), .A2(new_n19259_), .B1(pi0788), .B2(new_n19278_), .ZN(new_n19279_));
  OAI22_X1   g16843(.A1(new_n19279_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n19223_), .ZN(new_n19280_));
  INV_X1     g16844(.I(new_n19202_), .ZN(new_n19281_));
  NAND2_X1   g16845(.A1(new_n19281_), .A2(new_n13384_), .ZN(new_n19282_));
  NAND2_X1   g16846(.A1(new_n12943_), .A2(new_n19177_), .ZN(new_n19283_));
  NAND2_X1   g16847(.A1(new_n19282_), .A2(new_n19283_), .ZN(new_n19284_));
  NAND2_X1   g16848(.A1(new_n19218_), .A2(new_n12954_), .ZN(new_n19285_));
  NAND2_X1   g16849(.A1(new_n19285_), .A2(new_n12741_), .ZN(new_n19286_));
  NOR2_X1    g16850(.A1(new_n19176_), .A2(new_n12741_), .ZN(new_n19287_));
  INV_X1     g16851(.I(new_n19287_), .ZN(new_n19288_));
  AOI21_X1   g16852(.A1(new_n19286_), .A2(new_n19288_), .B(pi1157), .ZN(new_n19289_));
  INV_X1     g16853(.I(new_n19289_), .ZN(new_n19290_));
  NAND2_X1   g16854(.A1(new_n19176_), .A2(new_n12741_), .ZN(new_n19291_));
  OAI21_X1   g16855(.A1(new_n19285_), .A2(new_n12741_), .B(new_n19291_), .ZN(new_n19292_));
  OAI22_X1   g16856(.A1(new_n19290_), .A2(new_n12981_), .B1(new_n19292_), .B2(new_n15576_), .ZN(new_n19293_));
  AOI21_X1   g16857(.A1(new_n19284_), .A2(new_n15608_), .B(new_n19293_), .ZN(new_n19294_));
  OAI22_X1   g16858(.A1(new_n19280_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n19294_), .ZN(new_n19295_));
  NAND2_X1   g16859(.A1(new_n19295_), .A2(new_n13000_), .ZN(new_n19296_));
  AND2_X2    g16860(.A1(new_n19295_), .A2(new_n12975_), .Z(new_n19297_));
  OAI21_X1   g16861(.A1(new_n12965_), .A2(new_n19292_), .B(new_n19290_), .ZN(new_n19298_));
  NAND3_X1   g16862(.A1(new_n19218_), .A2(new_n12972_), .A3(new_n12954_), .ZN(new_n19299_));
  OAI21_X1   g16863(.A1(new_n19298_), .A2(new_n12972_), .B(new_n19299_), .ZN(new_n19300_));
  NOR2_X1    g16864(.A1(new_n19300_), .A2(new_n12975_), .ZN(new_n19301_));
  OAI21_X1   g16865(.A1(new_n19297_), .A2(new_n19301_), .B(new_n12740_), .ZN(new_n19302_));
  NOR2_X1    g16866(.A1(new_n19176_), .A2(new_n12975_), .ZN(new_n19303_));
  NOR2_X1    g16867(.A1(new_n17611_), .A2(new_n19176_), .ZN(new_n19304_));
  AOI21_X1   g16868(.A1(new_n19281_), .A2(new_n17611_), .B(new_n19304_), .ZN(new_n19305_));
  NOR2_X1    g16869(.A1(new_n19305_), .A2(pi0644), .ZN(new_n19306_));
  OAI21_X1   g16870(.A1(new_n19306_), .A2(new_n19303_), .B(pi0715), .ZN(new_n19307_));
  NAND3_X1   g16871(.A1(new_n19302_), .A2(new_n12739_), .A3(new_n19307_), .ZN(new_n19308_));
  NOR2_X1    g16872(.A1(new_n19300_), .A2(pi0644), .ZN(new_n19309_));
  AOI21_X1   g16873(.A1(new_n19295_), .A2(pi0644), .B(new_n19309_), .ZN(new_n19310_));
  NAND2_X1   g16874(.A1(new_n19177_), .A2(new_n12975_), .ZN(new_n19311_));
  OAI21_X1   g16875(.A1(new_n19305_), .A2(new_n12975_), .B(new_n19311_), .ZN(new_n19312_));
  AOI21_X1   g16876(.A1(new_n19312_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n19313_));
  OAI21_X1   g16877(.A1(new_n19310_), .A2(new_n12740_), .B(new_n19313_), .ZN(new_n19314_));
  NAND3_X1   g16878(.A1(new_n19308_), .A2(pi0790), .A3(new_n19314_), .ZN(new_n19315_));
  AOI21_X1   g16879(.A1(new_n19315_), .A2(new_n19296_), .B(new_n12738_), .ZN(new_n19316_));
  AOI21_X1   g16880(.A1(po1038), .A2(new_n9627_), .B(pi0832), .ZN(new_n19317_));
  NOR2_X1    g16881(.A1(new_n13193_), .A2(pi0179), .ZN(new_n19318_));
  AOI21_X1   g16882(.A1(new_n19318_), .A2(pi0644), .B(new_n12740_), .ZN(new_n19319_));
  NOR2_X1    g16883(.A1(new_n19318_), .A2(new_n13384_), .ZN(new_n19320_));
  NOR2_X1    g16884(.A1(new_n2609_), .A2(new_n9627_), .ZN(new_n19321_));
  INV_X1     g16885(.I(new_n19321_), .ZN(new_n19322_));
  NAND2_X1   g16886(.A1(new_n18659_), .A2(new_n9627_), .ZN(new_n19323_));
  NOR4_X1    g16887(.A1(new_n15012_), .A2(pi0741), .A3(new_n15011_), .A4(new_n19323_), .ZN(new_n19324_));
  NOR2_X1    g16888(.A1(new_n18327_), .A2(pi0741), .ZN(new_n19325_));
  NOR2_X1    g16889(.A1(new_n19325_), .A2(new_n9627_), .ZN(new_n19326_));
  NOR3_X1    g16890(.A1(new_n19326_), .A2(new_n16504_), .A3(new_n19324_), .ZN(new_n19327_));
  OAI21_X1   g16891(.A1(new_n19327_), .A2(new_n2610_), .B(new_n19322_), .ZN(new_n19328_));
  NAND2_X1   g16892(.A1(new_n19328_), .A2(new_n12761_), .ZN(new_n19329_));
  INV_X1     g16893(.I(new_n19318_), .ZN(new_n19330_));
  NAND2_X1   g16894(.A1(new_n19330_), .A2(new_n12760_), .ZN(new_n19331_));
  NAND2_X1   g16895(.A1(new_n19331_), .A2(new_n19329_), .ZN(new_n19332_));
  OAI22_X1   g16896(.A1(new_n19329_), .A2(pi0609), .B1(new_n13353_), .B2(new_n19318_), .ZN(new_n19333_));
  AND2_X2    g16897(.A1(new_n19333_), .A2(new_n12770_), .Z(new_n19334_));
  OAI22_X1   g16898(.A1(new_n19329_), .A2(new_n12766_), .B1(new_n12772_), .B2(new_n19318_), .ZN(new_n19335_));
  NAND2_X1   g16899(.A1(new_n19335_), .A2(pi1155), .ZN(new_n19336_));
  NAND2_X1   g16900(.A1(new_n19336_), .A2(pi0785), .ZN(new_n19337_));
  OAI22_X1   g16901(.A1(new_n19337_), .A2(new_n19334_), .B1(pi0785), .B2(new_n19332_), .ZN(new_n19338_));
  NAND2_X1   g16902(.A1(new_n19338_), .A2(new_n12779_), .ZN(new_n19339_));
  NAND2_X1   g16903(.A1(new_n19330_), .A2(pi0618), .ZN(new_n19340_));
  OAI21_X1   g16904(.A1(new_n19338_), .A2(pi0618), .B(new_n19340_), .ZN(new_n19341_));
  AND2_X2    g16905(.A1(new_n19341_), .A2(new_n12785_), .Z(new_n19342_));
  NOR2_X1    g16906(.A1(new_n19338_), .A2(new_n12781_), .ZN(new_n19343_));
  NOR2_X1    g16907(.A1(new_n19318_), .A2(pi0618), .ZN(new_n19344_));
  OAI21_X1   g16908(.A1(new_n19343_), .A2(new_n19344_), .B(pi1154), .ZN(new_n19345_));
  NAND2_X1   g16909(.A1(new_n19345_), .A2(pi0781), .ZN(new_n19346_));
  OAI21_X1   g16910(.A1(new_n19346_), .A2(new_n19342_), .B(new_n19339_), .ZN(new_n19347_));
  NAND2_X1   g16911(.A1(new_n19330_), .A2(pi0619), .ZN(new_n19348_));
  OAI21_X1   g16912(.A1(new_n19347_), .A2(pi0619), .B(new_n19348_), .ZN(new_n19349_));
  NAND2_X1   g16913(.A1(new_n19349_), .A2(new_n12791_), .ZN(new_n19350_));
  NAND2_X1   g16914(.A1(new_n19330_), .A2(new_n12793_), .ZN(new_n19351_));
  OAI21_X1   g16915(.A1(new_n19347_), .A2(new_n12793_), .B(new_n19351_), .ZN(new_n19352_));
  AOI21_X1   g16916(.A1(new_n19352_), .A2(pi1159), .B(new_n12796_), .ZN(new_n19353_));
  AOI22_X1   g16917(.A1(new_n19353_), .A2(new_n19350_), .B1(new_n12796_), .B2(new_n19347_), .ZN(new_n19354_));
  NOR2_X1    g16918(.A1(new_n19318_), .A2(new_n17504_), .ZN(new_n19355_));
  AOI21_X1   g16919(.A1(new_n19354_), .A2(new_n17504_), .B(new_n19355_), .ZN(new_n19356_));
  INV_X1     g16920(.I(new_n19356_), .ZN(new_n19357_));
  AOI21_X1   g16921(.A1(new_n19357_), .A2(new_n13384_), .B(new_n19320_), .ZN(new_n19358_));
  INV_X1     g16922(.I(new_n19358_), .ZN(new_n19359_));
  NAND2_X1   g16923(.A1(new_n19318_), .A2(new_n12984_), .ZN(new_n19360_));
  OAI21_X1   g16924(.A1(new_n19359_), .A2(new_n12984_), .B(new_n19360_), .ZN(new_n19361_));
  NAND2_X1   g16925(.A1(new_n19361_), .A2(new_n12975_), .ZN(new_n19362_));
  AOI21_X1   g16926(.A1(new_n19362_), .A2(new_n19319_), .B(pi1160), .ZN(new_n19363_));
  NOR2_X1    g16927(.A1(new_n19330_), .A2(new_n12870_), .ZN(new_n19364_));
  INV_X1     g16928(.I(new_n14131_), .ZN(new_n19365_));
  NOR2_X1    g16929(.A1(new_n13344_), .A2(pi0179), .ZN(new_n19366_));
  INV_X1     g16930(.I(new_n19366_), .ZN(new_n19367_));
  AOI21_X1   g16931(.A1(new_n13399_), .A2(new_n19367_), .B(pi0724), .ZN(new_n19368_));
  NAND2_X1   g16932(.A1(new_n18033_), .A2(pi0179), .ZN(new_n19369_));
  AOI21_X1   g16933(.A1(new_n19369_), .A2(new_n3265_), .B(new_n2610_), .ZN(new_n19370_));
  NOR2_X1    g16934(.A1(new_n14118_), .A2(pi0179), .ZN(new_n19371_));
  OAI21_X1   g16935(.A1(new_n19370_), .A2(new_n19371_), .B(new_n19368_), .ZN(new_n19372_));
  OAI21_X1   g16936(.A1(pi0724), .A2(new_n2610_), .B(new_n19318_), .ZN(new_n19373_));
  NAND2_X1   g16937(.A1(new_n19373_), .A2(new_n19372_), .ZN(new_n19374_));
  NOR3_X1    g16938(.A1(new_n19330_), .A2(new_n12758_), .A3(new_n14132_), .ZN(new_n19375_));
  AOI21_X1   g16939(.A1(new_n19374_), .A2(new_n19365_), .B(new_n19375_), .ZN(new_n19376_));
  INV_X1     g16940(.I(new_n19376_), .ZN(new_n19377_));
  AOI21_X1   g16941(.A1(new_n19377_), .A2(new_n12870_), .B(new_n19364_), .ZN(new_n19378_));
  NOR2_X1    g16942(.A1(new_n19318_), .A2(new_n12888_), .ZN(new_n19379_));
  AOI21_X1   g16943(.A1(new_n19378_), .A2(new_n12888_), .B(new_n19379_), .ZN(new_n19380_));
  NOR2_X1    g16944(.A1(new_n19330_), .A2(new_n12911_), .ZN(new_n19381_));
  AOI21_X1   g16945(.A1(new_n19380_), .A2(new_n12911_), .B(new_n19381_), .ZN(new_n19382_));
  AND2_X2    g16946(.A1(new_n19382_), .A2(new_n13392_), .Z(new_n19383_));
  AOI21_X1   g16947(.A1(new_n12817_), .A2(new_n19330_), .B(new_n19383_), .ZN(new_n19384_));
  INV_X1     g16948(.I(new_n19384_), .ZN(new_n19385_));
  NAND2_X1   g16949(.A1(new_n19385_), .A2(new_n12920_), .ZN(new_n19386_));
  NAND2_X1   g16950(.A1(new_n19330_), .A2(pi0628), .ZN(new_n19387_));
  AOI21_X1   g16951(.A1(new_n19386_), .A2(new_n19387_), .B(pi1156), .ZN(new_n19388_));
  NAND2_X1   g16952(.A1(new_n19330_), .A2(new_n12920_), .ZN(new_n19389_));
  NAND2_X1   g16953(.A1(new_n19385_), .A2(pi0628), .ZN(new_n19390_));
  AOI21_X1   g16954(.A1(new_n19390_), .A2(new_n19389_), .B(new_n12742_), .ZN(new_n19391_));
  NOR3_X1    g16955(.A1(new_n19388_), .A2(new_n19391_), .A3(new_n12937_), .ZN(new_n19392_));
  AOI21_X1   g16956(.A1(new_n12937_), .A2(new_n19384_), .B(new_n19392_), .ZN(new_n19393_));
  NAND2_X1   g16957(.A1(new_n19393_), .A2(new_n12741_), .ZN(new_n19394_));
  NAND2_X1   g16958(.A1(new_n19330_), .A2(pi0647), .ZN(new_n19395_));
  AOI21_X1   g16959(.A1(new_n19394_), .A2(new_n19395_), .B(pi1157), .ZN(new_n19396_));
  NAND2_X1   g16960(.A1(new_n19393_), .A2(pi0647), .ZN(new_n19397_));
  NAND2_X1   g16961(.A1(new_n19330_), .A2(new_n12741_), .ZN(new_n19398_));
  AOI21_X1   g16962(.A1(new_n19397_), .A2(new_n19398_), .B(new_n12965_), .ZN(new_n19399_));
  OR2_X2     g16963(.A1(new_n19399_), .A2(new_n12972_), .Z(new_n19400_));
  OAI22_X1   g16964(.A1(new_n19400_), .A2(new_n19396_), .B1(pi0787), .B2(new_n19393_), .ZN(new_n19401_));
  AOI21_X1   g16965(.A1(new_n19401_), .A2(pi0644), .B(pi0715), .ZN(new_n19402_));
  NOR2_X1    g16966(.A1(new_n19388_), .A2(new_n12919_), .ZN(new_n19403_));
  AOI21_X1   g16967(.A1(new_n19356_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n19404_));
  AOI21_X1   g16968(.A1(new_n19330_), .A2(new_n12747_), .B(pi0641), .ZN(new_n19405_));
  NAND2_X1   g16969(.A1(new_n19354_), .A2(pi0626), .ZN(new_n19406_));
  AOI21_X1   g16970(.A1(new_n19406_), .A2(new_n19405_), .B(new_n12745_), .ZN(new_n19407_));
  AOI21_X1   g16971(.A1(new_n19382_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n19408_));
  AOI21_X1   g16972(.A1(new_n19327_), .A2(pi0724), .B(new_n2610_), .ZN(new_n19409_));
  NAND2_X1   g16973(.A1(new_n19367_), .A2(new_n14169_), .ZN(new_n19410_));
  INV_X1     g16974(.I(new_n19410_), .ZN(new_n19411_));
  NOR2_X1    g16975(.A1(new_n14177_), .A2(pi0179), .ZN(new_n19412_));
  NOR2_X1    g16976(.A1(new_n15835_), .A2(new_n9627_), .ZN(new_n19413_));
  OAI21_X1   g16977(.A1(new_n19412_), .A2(new_n19413_), .B(new_n2627_), .ZN(new_n19414_));
  NOR2_X1    g16978(.A1(new_n14182_), .A2(pi0179), .ZN(new_n19415_));
  NOR2_X1    g16979(.A1(new_n14184_), .A2(new_n9627_), .ZN(new_n19416_));
  OAI21_X1   g16980(.A1(new_n19415_), .A2(new_n19416_), .B(pi0039), .ZN(new_n19417_));
  AOI21_X1   g16981(.A1(new_n19417_), .A2(new_n19414_), .B(pi0038), .ZN(new_n19418_));
  OAI21_X1   g16982(.A1(new_n19418_), .A2(new_n19411_), .B(pi0741), .ZN(new_n19419_));
  AOI21_X1   g16983(.A1(new_n18437_), .A2(new_n18424_), .B(new_n9627_), .ZN(new_n19420_));
  NAND2_X1   g16984(.A1(new_n15107_), .A2(new_n15109_), .ZN(new_n19421_));
  NAND2_X1   g16985(.A1(new_n19421_), .A2(new_n18755_), .ZN(new_n19422_));
  NOR2_X1    g16986(.A1(new_n19422_), .A2(pi0179), .ZN(new_n19423_));
  OAI21_X1   g16987(.A1(new_n19423_), .A2(new_n19420_), .B(new_n16500_), .ZN(new_n19424_));
  NAND3_X1   g16988(.A1(new_n19419_), .A2(new_n19424_), .A3(new_n16499_), .ZN(new_n19425_));
  AOI21_X1   g16989(.A1(new_n19425_), .A2(new_n19409_), .B(new_n19321_), .ZN(new_n19426_));
  INV_X1     g16990(.I(new_n14163_), .ZN(new_n19427_));
  OAI21_X1   g16991(.A1(new_n19427_), .A2(pi0179), .B(new_n12841_), .ZN(new_n19428_));
  AOI21_X1   g16992(.A1(new_n19373_), .A2(new_n19372_), .B(pi0625), .ZN(new_n19429_));
  OAI21_X1   g16993(.A1(new_n19429_), .A2(new_n19428_), .B(pi0608), .ZN(new_n19430_));
  NOR2_X1    g16994(.A1(new_n19328_), .A2(pi0625), .ZN(new_n19431_));
  NOR2_X1    g16995(.A1(new_n19431_), .A2(new_n12841_), .ZN(new_n19432_));
  NAND2_X1   g16996(.A1(new_n19426_), .A2(pi0625), .ZN(new_n19433_));
  AOI21_X1   g16997(.A1(new_n19433_), .A2(new_n19432_), .B(new_n19430_), .ZN(new_n19434_));
  INV_X1     g16998(.I(new_n14199_), .ZN(new_n19435_));
  OAI21_X1   g16999(.A1(new_n19435_), .A2(pi0179), .B(pi1153), .ZN(new_n19436_));
  AOI21_X1   g17000(.A1(new_n19373_), .A2(new_n19372_), .B(new_n13521_), .ZN(new_n19437_));
  OAI21_X1   g17001(.A1(new_n19437_), .A2(new_n19436_), .B(new_n13560_), .ZN(new_n19438_));
  OAI21_X1   g17002(.A1(new_n19328_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n19439_));
  AOI21_X1   g17003(.A1(new_n19426_), .A2(new_n13521_), .B(new_n19439_), .ZN(new_n19440_));
  OAI21_X1   g17004(.A1(new_n19440_), .A2(new_n19438_), .B(pi0778), .ZN(new_n19441_));
  OAI22_X1   g17005(.A1(new_n19434_), .A2(new_n19441_), .B1(pi0778), .B2(new_n19426_), .ZN(new_n19442_));
  NOR2_X1    g17006(.A1(new_n19334_), .A2(new_n13829_), .ZN(new_n19443_));
  OAI21_X1   g17007(.A1(new_n19376_), .A2(pi0609), .B(pi1155), .ZN(new_n19444_));
  NOR2_X1    g17008(.A1(new_n19442_), .A2(new_n12766_), .ZN(new_n19445_));
  OAI21_X1   g17009(.A1(new_n19445_), .A2(new_n19444_), .B(new_n19443_), .ZN(new_n19446_));
  AOI21_X1   g17010(.A1(new_n19335_), .A2(pi1155), .B(pi0660), .ZN(new_n19447_));
  AOI21_X1   g17011(.A1(new_n19377_), .A2(pi0609), .B(pi1155), .ZN(new_n19448_));
  OAI21_X1   g17012(.A1(new_n19442_), .A2(pi0609), .B(new_n19448_), .ZN(new_n19449_));
  AOI21_X1   g17013(.A1(new_n19449_), .A2(new_n19447_), .B(new_n12764_), .ZN(new_n19450_));
  AOI22_X1   g17014(.A1(new_n19450_), .A2(new_n19446_), .B1(new_n12764_), .B2(new_n19442_), .ZN(new_n19451_));
  NOR2_X1    g17015(.A1(new_n19451_), .A2(pi0781), .ZN(new_n19452_));
  INV_X1     g17016(.I(new_n19452_), .ZN(new_n19453_));
  OR2_X2     g17017(.A1(new_n19342_), .A2(new_n12880_), .Z(new_n19454_));
  INV_X1     g17018(.I(new_n19378_), .ZN(new_n19455_));
  AOI21_X1   g17019(.A1(new_n19455_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n19456_));
  NAND2_X1   g17020(.A1(new_n19451_), .A2(pi0618), .ZN(new_n19457_));
  AOI21_X1   g17021(.A1(new_n19457_), .A2(new_n19456_), .B(new_n19454_), .ZN(new_n19458_));
  NAND2_X1   g17022(.A1(new_n19345_), .A2(new_n12880_), .ZN(new_n19459_));
  AOI21_X1   g17023(.A1(new_n19455_), .A2(pi0618), .B(pi1154), .ZN(new_n19460_));
  INV_X1     g17024(.I(new_n19460_), .ZN(new_n19461_));
  AOI21_X1   g17025(.A1(new_n19451_), .A2(new_n12781_), .B(new_n19461_), .ZN(new_n19462_));
  OAI21_X1   g17026(.A1(new_n19462_), .A2(new_n19459_), .B(pi0781), .ZN(new_n19463_));
  OAI21_X1   g17027(.A1(new_n19463_), .A2(new_n19458_), .B(new_n19453_), .ZN(new_n19464_));
  AND2_X2    g17028(.A1(new_n19464_), .A2(new_n12796_), .Z(new_n19465_));
  AOI21_X1   g17029(.A1(new_n19349_), .A2(new_n12791_), .B(new_n12895_), .ZN(new_n19466_));
  AOI21_X1   g17030(.A1(new_n19380_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n19467_));
  OAI21_X1   g17031(.A1(new_n19464_), .A2(new_n12793_), .B(new_n19467_), .ZN(new_n19468_));
  NAND2_X1   g17032(.A1(new_n19468_), .A2(new_n19466_), .ZN(new_n19469_));
  AOI21_X1   g17033(.A1(new_n19352_), .A2(pi1159), .B(pi0648), .ZN(new_n19470_));
  AOI21_X1   g17034(.A1(new_n19380_), .A2(pi0619), .B(pi1159), .ZN(new_n19471_));
  OAI21_X1   g17035(.A1(new_n19464_), .A2(pi0619), .B(new_n19471_), .ZN(new_n19472_));
  AOI21_X1   g17036(.A1(new_n19472_), .A2(new_n19470_), .B(new_n12796_), .ZN(new_n19473_));
  AOI21_X1   g17037(.A1(new_n19473_), .A2(new_n19469_), .B(new_n19465_), .ZN(new_n19474_));
  OAI21_X1   g17038(.A1(new_n19474_), .A2(new_n12747_), .B(new_n19408_), .ZN(new_n19475_));
  NAND2_X1   g17039(.A1(new_n19475_), .A2(new_n19407_), .ZN(new_n19476_));
  AOI21_X1   g17040(.A1(new_n19330_), .A2(pi0626), .B(new_n12814_), .ZN(new_n19477_));
  NAND2_X1   g17041(.A1(new_n19354_), .A2(new_n12747_), .ZN(new_n19478_));
  AOI21_X1   g17042(.A1(new_n19478_), .A2(new_n19477_), .B(pi1158), .ZN(new_n19479_));
  AOI21_X1   g17043(.A1(new_n19382_), .A2(pi0626), .B(pi0641), .ZN(new_n19480_));
  OAI21_X1   g17044(.A1(new_n19474_), .A2(pi0626), .B(new_n19480_), .ZN(new_n19481_));
  AOI21_X1   g17045(.A1(new_n19481_), .A2(new_n19479_), .B(new_n12808_), .ZN(new_n19482_));
  AND2_X2    g17046(.A1(new_n19474_), .A2(new_n12808_), .Z(new_n19483_));
  AOI21_X1   g17047(.A1(new_n19482_), .A2(new_n19476_), .B(new_n19483_), .ZN(new_n19484_));
  OAI21_X1   g17048(.A1(new_n19484_), .A2(new_n12920_), .B(new_n19404_), .ZN(new_n19485_));
  NAND2_X1   g17049(.A1(new_n19485_), .A2(new_n19403_), .ZN(new_n19486_));
  NOR2_X1    g17050(.A1(new_n19391_), .A2(pi0629), .ZN(new_n19487_));
  AOI21_X1   g17051(.A1(new_n19356_), .A2(pi0628), .B(pi1156), .ZN(new_n19488_));
  OAI21_X1   g17052(.A1(new_n19484_), .A2(pi0628), .B(new_n19488_), .ZN(new_n19489_));
  AOI21_X1   g17053(.A1(new_n19489_), .A2(new_n19487_), .B(new_n12937_), .ZN(new_n19490_));
  AND2_X2    g17054(.A1(new_n19484_), .A2(new_n12937_), .Z(new_n19491_));
  AOI21_X1   g17055(.A1(new_n19490_), .A2(new_n19486_), .B(new_n19491_), .ZN(new_n19492_));
  OR2_X2     g17056(.A1(new_n19492_), .A2(pi0787), .Z(new_n19493_));
  OR2_X2     g17057(.A1(new_n19396_), .A2(new_n12981_), .Z(new_n19494_));
  AOI21_X1   g17058(.A1(new_n19358_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n19495_));
  NAND2_X1   g17059(.A1(new_n19492_), .A2(pi0647), .ZN(new_n19496_));
  AOI21_X1   g17060(.A1(new_n19496_), .A2(new_n19495_), .B(new_n19494_), .ZN(new_n19497_));
  OR2_X2     g17061(.A1(new_n19399_), .A2(pi0630), .Z(new_n19498_));
  OAI21_X1   g17062(.A1(new_n19359_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n19499_));
  AOI21_X1   g17063(.A1(new_n19492_), .A2(new_n12741_), .B(new_n19499_), .ZN(new_n19500_));
  OAI21_X1   g17064(.A1(new_n19500_), .A2(new_n19498_), .B(pi0787), .ZN(new_n19501_));
  OAI21_X1   g17065(.A1(new_n19501_), .A2(new_n19497_), .B(new_n19493_), .ZN(new_n19502_));
  OAI21_X1   g17066(.A1(new_n19502_), .A2(pi0644), .B(new_n19402_), .ZN(new_n19503_));
  NAND2_X1   g17067(.A1(new_n19503_), .A2(new_n19363_), .ZN(new_n19504_));
  AOI21_X1   g17068(.A1(new_n19318_), .A2(new_n12975_), .B(pi0715), .ZN(new_n19505_));
  NAND2_X1   g17069(.A1(new_n19361_), .A2(pi0644), .ZN(new_n19506_));
  AOI21_X1   g17070(.A1(new_n19506_), .A2(new_n19505_), .B(new_n12739_), .ZN(new_n19507_));
  NOR2_X1    g17071(.A1(new_n19401_), .A2(pi0644), .ZN(new_n19508_));
  AOI21_X1   g17072(.A1(new_n19502_), .A2(pi0644), .B(new_n19508_), .ZN(new_n19509_));
  OAI21_X1   g17073(.A1(new_n19509_), .A2(new_n12740_), .B(new_n19507_), .ZN(new_n19510_));
  NAND3_X1   g17074(.A1(new_n19510_), .A2(new_n19504_), .A3(pi0790), .ZN(new_n19511_));
  AOI21_X1   g17075(.A1(new_n19502_), .A2(new_n13000_), .B(po1038), .ZN(new_n19512_));
  NAND2_X1   g17076(.A1(new_n19511_), .A2(new_n19512_), .ZN(new_n19513_));
  AOI21_X1   g17077(.A1(new_n19513_), .A2(new_n19317_), .B(new_n19316_), .ZN(po0336));
  NOR2_X1    g17078(.A1(new_n13340_), .A2(pi0753), .ZN(new_n19515_));
  NOR2_X1    g17079(.A1(new_n3042_), .A2(pi0180), .ZN(new_n19516_));
  NOR2_X1    g17080(.A1(new_n19515_), .A2(new_n19516_), .ZN(new_n19517_));
  NOR3_X1    g17081(.A1(new_n19517_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n19518_));
  INV_X1     g17082(.I(new_n19515_), .ZN(new_n19519_));
  NOR2_X1    g17083(.A1(new_n19519_), .A2(new_n13354_), .ZN(new_n19520_));
  NOR3_X1    g17084(.A1(new_n19520_), .A2(new_n12762_), .A3(new_n19517_), .ZN(new_n19521_));
  NOR2_X1    g17085(.A1(new_n19521_), .A2(new_n12770_), .ZN(new_n19522_));
  NOR3_X1    g17086(.A1(new_n19520_), .A2(pi1155), .A3(new_n19516_), .ZN(new_n19523_));
  NOR3_X1    g17087(.A1(new_n19522_), .A2(new_n12764_), .A3(new_n19523_), .ZN(new_n19524_));
  NOR2_X1    g17088(.A1(new_n19524_), .A2(new_n19518_), .ZN(new_n19525_));
  INV_X1     g17089(.I(new_n19525_), .ZN(new_n19526_));
  AOI21_X1   g17090(.A1(new_n19526_), .A2(new_n12783_), .B(pi1154), .ZN(new_n19527_));
  AOI21_X1   g17091(.A1(new_n19526_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n19528_));
  NOR3_X1    g17092(.A1(new_n19527_), .A2(new_n19528_), .A3(new_n12779_), .ZN(new_n19529_));
  AOI21_X1   g17093(.A1(new_n12779_), .A2(new_n19526_), .B(new_n19529_), .ZN(new_n19530_));
  OAI21_X1   g17094(.A1(new_n19530_), .A2(new_n17229_), .B(new_n12791_), .ZN(new_n19531_));
  OAI21_X1   g17095(.A1(new_n19530_), .A2(new_n17232_), .B(pi1159), .ZN(new_n19532_));
  NAND3_X1   g17096(.A1(new_n19531_), .A2(new_n19532_), .A3(pi0789), .ZN(new_n19533_));
  OAI21_X1   g17097(.A1(pi0789), .A2(new_n19530_), .B(new_n19533_), .ZN(new_n19534_));
  INV_X1     g17098(.I(new_n19516_), .ZN(new_n19535_));
  NAND2_X1   g17099(.A1(new_n12818_), .A2(new_n19535_), .ZN(new_n19536_));
  OAI21_X1   g17100(.A1(new_n19534_), .A2(new_n12818_), .B(new_n19536_), .ZN(new_n19537_));
  AOI21_X1   g17101(.A1(new_n12826_), .A2(new_n16558_), .B(new_n19516_), .ZN(new_n19538_));
  NOR2_X1    g17102(.A1(new_n19516_), .A2(pi1153), .ZN(new_n19539_));
  NOR2_X1    g17103(.A1(new_n12834_), .A2(pi0702), .ZN(new_n19540_));
  INV_X1     g17104(.I(new_n19540_), .ZN(new_n19541_));
  NAND2_X1   g17105(.A1(new_n19541_), .A2(new_n19539_), .ZN(new_n19542_));
  NOR2_X1    g17106(.A1(new_n19540_), .A2(new_n19538_), .ZN(new_n19543_));
  NOR2_X1    g17107(.A1(new_n19543_), .A2(new_n12841_), .ZN(new_n19544_));
  INV_X1     g17108(.I(new_n19544_), .ZN(new_n19545_));
  NAND3_X1   g17109(.A1(new_n19545_), .A2(pi0778), .A3(new_n19542_), .ZN(new_n19546_));
  OAI21_X1   g17110(.A1(pi0778), .A2(new_n19538_), .B(new_n19546_), .ZN(new_n19547_));
  NAND2_X1   g17111(.A1(new_n19547_), .A2(new_n17187_), .ZN(new_n19548_));
  NOR2_X1    g17112(.A1(new_n19548_), .A2(new_n12889_), .ZN(new_n19549_));
  NAND2_X1   g17113(.A1(new_n19549_), .A2(new_n18203_), .ZN(new_n19550_));
  NOR2_X1    g17114(.A1(new_n19550_), .A2(new_n17884_), .ZN(new_n19551_));
  INV_X1     g17115(.I(new_n19551_), .ZN(new_n19552_));
  OAI22_X1   g17116(.A1(new_n19537_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n19552_), .ZN(new_n19553_));
  AND2_X2    g17117(.A1(new_n19553_), .A2(new_n12919_), .Z(new_n19554_));
  OAI22_X1   g17118(.A1(new_n19537_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n19552_), .ZN(new_n19555_));
  AOI21_X1   g17119(.A1(pi0629), .A2(new_n19555_), .B(new_n19554_), .ZN(new_n19556_));
  INV_X1     g17120(.I(new_n19523_), .ZN(new_n19557_));
  NOR2_X1    g17121(.A1(new_n19538_), .A2(new_n12754_), .ZN(new_n19558_));
  NOR3_X1    g17122(.A1(new_n19558_), .A2(new_n19515_), .A3(new_n19516_), .ZN(new_n19559_));
  NAND2_X1   g17123(.A1(new_n19559_), .A2(new_n12758_), .ZN(new_n19560_));
  NAND2_X1   g17124(.A1(new_n19558_), .A2(pi0625), .ZN(new_n19561_));
  NAND3_X1   g17125(.A1(new_n19561_), .A2(pi1153), .A3(new_n19517_), .ZN(new_n19562_));
  NAND3_X1   g17126(.A1(new_n19542_), .A2(pi0608), .A3(new_n19562_), .ZN(new_n19563_));
  INV_X1     g17127(.I(new_n19561_), .ZN(new_n19564_));
  OAI21_X1   g17128(.A1(new_n19564_), .A2(new_n19559_), .B(new_n19539_), .ZN(new_n19565_));
  NAND3_X1   g17129(.A1(new_n19545_), .A2(new_n13560_), .A3(new_n19565_), .ZN(new_n19566_));
  NAND3_X1   g17130(.A1(new_n19566_), .A2(pi0778), .A3(new_n19563_), .ZN(new_n19567_));
  AOI21_X1   g17131(.A1(new_n19567_), .A2(new_n19560_), .B(new_n12766_), .ZN(new_n19568_));
  NOR2_X1    g17132(.A1(new_n19547_), .A2(pi0609), .ZN(new_n19569_));
  OAI21_X1   g17133(.A1(new_n19569_), .A2(new_n19568_), .B(pi1155), .ZN(new_n19570_));
  NAND3_X1   g17134(.A1(new_n19570_), .A2(pi0660), .A3(new_n19557_), .ZN(new_n19571_));
  NAND2_X1   g17135(.A1(new_n19567_), .A2(new_n19560_), .ZN(new_n19572_));
  NOR2_X1    g17136(.A1(new_n19547_), .A2(new_n12766_), .ZN(new_n19573_));
  AOI21_X1   g17137(.A1(new_n19572_), .A2(new_n12766_), .B(new_n19573_), .ZN(new_n19574_));
  NOR2_X1    g17138(.A1(new_n19522_), .A2(pi0660), .ZN(new_n19575_));
  OAI21_X1   g17139(.A1(new_n19574_), .A2(pi1155), .B(new_n19575_), .ZN(new_n19576_));
  NAND3_X1   g17140(.A1(new_n19576_), .A2(new_n19571_), .A3(pi0785), .ZN(new_n19577_));
  NAND2_X1   g17141(.A1(new_n19572_), .A2(new_n12764_), .ZN(new_n19578_));
  NAND2_X1   g17142(.A1(new_n19577_), .A2(new_n19578_), .ZN(new_n19579_));
  NAND2_X1   g17143(.A1(new_n19579_), .A2(new_n12781_), .ZN(new_n19580_));
  NAND2_X1   g17144(.A1(new_n19548_), .A2(pi0618), .ZN(new_n19581_));
  AOI21_X1   g17145(.A1(new_n19580_), .A2(new_n19581_), .B(pi1154), .ZN(new_n19582_));
  NOR3_X1    g17146(.A1(new_n19582_), .A2(pi0627), .A3(new_n19528_), .ZN(new_n19583_));
  NAND2_X1   g17147(.A1(new_n19548_), .A2(new_n12781_), .ZN(new_n19584_));
  NAND2_X1   g17148(.A1(new_n19579_), .A2(pi0618), .ZN(new_n19585_));
  AOI21_X1   g17149(.A1(new_n19585_), .A2(new_n19584_), .B(new_n12785_), .ZN(new_n19586_));
  NOR3_X1    g17150(.A1(new_n19586_), .A2(new_n12880_), .A3(new_n19527_), .ZN(new_n19587_));
  OR3_X2     g17151(.A1(new_n19583_), .A2(new_n19587_), .A3(new_n12779_), .Z(new_n19588_));
  NAND2_X1   g17152(.A1(new_n19579_), .A2(new_n12779_), .ZN(new_n19589_));
  NAND2_X1   g17153(.A1(new_n19588_), .A2(new_n19589_), .ZN(new_n19590_));
  AOI21_X1   g17154(.A1(new_n19590_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n19591_));
  NOR2_X1    g17155(.A1(new_n19549_), .A2(pi0619), .ZN(new_n19592_));
  AOI21_X1   g17156(.A1(new_n19588_), .A2(new_n19589_), .B(new_n12793_), .ZN(new_n19593_));
  OAI21_X1   g17157(.A1(new_n19593_), .A2(new_n19592_), .B(pi1159), .ZN(new_n19594_));
  NAND3_X1   g17158(.A1(new_n19594_), .A2(pi0648), .A3(new_n19531_), .ZN(new_n19595_));
  NAND2_X1   g17159(.A1(new_n19590_), .A2(new_n12793_), .ZN(new_n19596_));
  OAI21_X1   g17160(.A1(new_n12793_), .A2(new_n19549_), .B(new_n19596_), .ZN(new_n19597_));
  NAND2_X1   g17161(.A1(new_n19597_), .A2(new_n12791_), .ZN(new_n19598_));
  NAND3_X1   g17162(.A1(new_n19598_), .A2(new_n12895_), .A3(new_n19532_), .ZN(new_n19599_));
  NAND3_X1   g17163(.A1(new_n19599_), .A2(pi0789), .A3(new_n19595_), .ZN(new_n19600_));
  NOR2_X1    g17164(.A1(new_n19535_), .A2(new_n12747_), .ZN(new_n19601_));
  AND2_X2    g17165(.A1(new_n19534_), .A2(new_n12747_), .Z(new_n19602_));
  OAI21_X1   g17166(.A1(new_n19602_), .A2(new_n19601_), .B(new_n12815_), .ZN(new_n19603_));
  INV_X1     g17167(.I(new_n19550_), .ZN(new_n19604_));
  NAND2_X1   g17168(.A1(new_n19534_), .A2(pi0626), .ZN(new_n19605_));
  OAI21_X1   g17169(.A1(pi0626), .A2(new_n19535_), .B(new_n19605_), .ZN(new_n19606_));
  AOI22_X1   g17170(.A1(new_n19606_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n19604_), .ZN(new_n19607_));
  NAND2_X1   g17171(.A1(new_n19607_), .A2(new_n19603_), .ZN(new_n19608_));
  AOI22_X1   g17172(.A1(new_n19600_), .A2(new_n19591_), .B1(pi0788), .B2(new_n19608_), .ZN(new_n19609_));
  OAI22_X1   g17173(.A1(new_n19609_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n19556_), .ZN(new_n19610_));
  NAND2_X1   g17174(.A1(new_n19537_), .A2(new_n13384_), .ZN(new_n19611_));
  NAND2_X1   g17175(.A1(new_n12943_), .A2(new_n19535_), .ZN(new_n19612_));
  NAND2_X1   g17176(.A1(new_n19611_), .A2(new_n19612_), .ZN(new_n19613_));
  NOR2_X1    g17177(.A1(new_n19552_), .A2(new_n12953_), .ZN(new_n19614_));
  NOR2_X1    g17178(.A1(new_n19614_), .A2(pi0647), .ZN(new_n19615_));
  NOR2_X1    g17179(.A1(new_n19516_), .A2(new_n12741_), .ZN(new_n19616_));
  OAI21_X1   g17180(.A1(new_n19615_), .A2(new_n19616_), .B(new_n12965_), .ZN(new_n19617_));
  NAND2_X1   g17181(.A1(new_n19614_), .A2(pi0647), .ZN(new_n19618_));
  OAI21_X1   g17182(.A1(pi0647), .A2(new_n19535_), .B(new_n19618_), .ZN(new_n19619_));
  OAI22_X1   g17183(.A1(new_n19619_), .A2(new_n15576_), .B1(new_n19617_), .B2(new_n12981_), .ZN(new_n19620_));
  AOI21_X1   g17184(.A1(new_n19613_), .A2(new_n15608_), .B(new_n19620_), .ZN(new_n19621_));
  OAI22_X1   g17185(.A1(new_n19610_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n19621_), .ZN(new_n19622_));
  NAND2_X1   g17186(.A1(new_n19622_), .A2(new_n13000_), .ZN(new_n19623_));
  AND2_X2    g17187(.A1(new_n19622_), .A2(new_n12975_), .Z(new_n19624_));
  OAI21_X1   g17188(.A1(new_n19619_), .A2(new_n12965_), .B(new_n19617_), .ZN(new_n19625_));
  NAND2_X1   g17189(.A1(new_n19614_), .A2(new_n12972_), .ZN(new_n19626_));
  OAI21_X1   g17190(.A1(new_n19625_), .A2(new_n12972_), .B(new_n19626_), .ZN(new_n19627_));
  NOR2_X1    g17191(.A1(new_n19627_), .A2(new_n12975_), .ZN(new_n19628_));
  OAI21_X1   g17192(.A1(new_n19624_), .A2(new_n19628_), .B(new_n12740_), .ZN(new_n19629_));
  NAND2_X1   g17193(.A1(new_n19535_), .A2(pi0644), .ZN(new_n19630_));
  NOR2_X1    g17194(.A1(new_n17611_), .A2(new_n19516_), .ZN(new_n19631_));
  AOI21_X1   g17195(.A1(new_n19537_), .A2(new_n17611_), .B(new_n19631_), .ZN(new_n19632_));
  OAI21_X1   g17196(.A1(new_n19632_), .A2(pi0644), .B(new_n19630_), .ZN(new_n19633_));
  NAND2_X1   g17197(.A1(new_n19633_), .A2(pi0715), .ZN(new_n19634_));
  NAND3_X1   g17198(.A1(new_n19629_), .A2(new_n12739_), .A3(new_n19634_), .ZN(new_n19635_));
  NOR2_X1    g17199(.A1(new_n19627_), .A2(pi0644), .ZN(new_n19636_));
  AOI21_X1   g17200(.A1(new_n19622_), .A2(pi0644), .B(new_n19636_), .ZN(new_n19637_));
  NAND2_X1   g17201(.A1(new_n19535_), .A2(new_n12975_), .ZN(new_n19638_));
  OAI21_X1   g17202(.A1(new_n19632_), .A2(new_n12975_), .B(new_n19638_), .ZN(new_n19639_));
  AOI21_X1   g17203(.A1(new_n19639_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n19640_));
  OAI21_X1   g17204(.A1(new_n19637_), .A2(new_n12740_), .B(new_n19640_), .ZN(new_n19641_));
  NAND3_X1   g17205(.A1(new_n19635_), .A2(pi0790), .A3(new_n19641_), .ZN(new_n19642_));
  NAND2_X1   g17206(.A1(new_n19642_), .A2(new_n19623_), .ZN(new_n19643_));
  AOI21_X1   g17207(.A1(po1038), .A2(new_n5657_), .B(pi0832), .ZN(new_n19644_));
  NAND2_X1   g17208(.A1(new_n13192_), .A2(new_n5657_), .ZN(new_n19645_));
  INV_X1     g17209(.I(new_n19645_), .ZN(new_n19646_));
  AOI21_X1   g17210(.A1(new_n19646_), .A2(pi0644), .B(new_n12740_), .ZN(new_n19647_));
  NAND2_X1   g17211(.A1(new_n19645_), .A2(new_n12984_), .ZN(new_n19648_));
  NOR2_X1    g17212(.A1(new_n19646_), .A2(new_n13384_), .ZN(new_n19649_));
  NAND2_X1   g17213(.A1(new_n2610_), .A2(pi0180), .ZN(new_n19650_));
  INV_X1     g17214(.I(new_n13798_), .ZN(new_n19651_));
  OAI22_X1   g17215(.A1(new_n19651_), .A2(new_n5657_), .B1(new_n16550_), .B2(new_n13060_), .ZN(new_n19652_));
  NAND2_X1   g17216(.A1(new_n5657_), .A2(pi0753), .ZN(new_n19653_));
  OAI21_X1   g17217(.A1(new_n13334_), .A2(pi0180), .B(new_n16550_), .ZN(new_n19654_));
  AOI22_X1   g17218(.A1(new_n19654_), .A2(new_n19653_), .B1(new_n2627_), .B2(new_n19652_), .ZN(new_n19655_));
  OAI22_X1   g17219(.A1(new_n14065_), .A2(new_n16550_), .B1(new_n5657_), .B2(new_n14067_), .ZN(new_n19656_));
  NAND2_X1   g17220(.A1(new_n19656_), .A2(pi0039), .ZN(new_n19657_));
  NAND2_X1   g17221(.A1(new_n19655_), .A2(new_n19657_), .ZN(new_n19658_));
  NOR2_X1    g17222(.A1(new_n13344_), .A2(pi0180), .ZN(new_n19659_));
  NOR2_X1    g17223(.A1(new_n19659_), .A2(new_n3265_), .ZN(new_n19660_));
  NAND2_X1   g17224(.A1(new_n13341_), .A2(new_n16550_), .ZN(new_n19661_));
  AOI22_X1   g17225(.A1(new_n19658_), .A2(new_n3265_), .B1(new_n19660_), .B2(new_n19661_), .ZN(new_n19662_));
  OAI21_X1   g17226(.A1(new_n19662_), .A2(new_n2610_), .B(new_n19650_), .ZN(new_n19663_));
  NAND2_X1   g17227(.A1(new_n19663_), .A2(new_n12761_), .ZN(new_n19664_));
  INV_X1     g17228(.I(new_n19664_), .ZN(new_n19665_));
  NOR2_X1    g17229(.A1(new_n19646_), .A2(new_n12761_), .ZN(new_n19666_));
  NOR3_X1    g17230(.A1(new_n19665_), .A2(pi0785), .A3(new_n19666_), .ZN(new_n19667_));
  AOI22_X1   g17231(.A1(new_n19665_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n19645_), .ZN(new_n19668_));
  NOR2_X1    g17232(.A1(new_n19668_), .A2(pi1155), .ZN(new_n19669_));
  AOI22_X1   g17233(.A1(new_n19665_), .A2(pi0609), .B1(new_n13357_), .B2(new_n19645_), .ZN(new_n19670_));
  NOR2_X1    g17234(.A1(new_n19670_), .A2(new_n12770_), .ZN(new_n19671_));
  NOR3_X1    g17235(.A1(new_n19671_), .A2(new_n19669_), .A3(new_n12764_), .ZN(new_n19672_));
  NOR2_X1    g17236(.A1(new_n19672_), .A2(new_n19667_), .ZN(new_n19673_));
  NOR2_X1    g17237(.A1(new_n19673_), .A2(pi0781), .ZN(new_n19674_));
  NOR3_X1    g17238(.A1(new_n19672_), .A2(pi0618), .A3(new_n19667_), .ZN(new_n19675_));
  NOR2_X1    g17239(.A1(new_n19646_), .A2(new_n12781_), .ZN(new_n19676_));
  OAI21_X1   g17240(.A1(new_n19675_), .A2(new_n19676_), .B(new_n12785_), .ZN(new_n19677_));
  NAND2_X1   g17241(.A1(new_n19673_), .A2(pi0618), .ZN(new_n19678_));
  NAND2_X1   g17242(.A1(new_n19645_), .A2(new_n12781_), .ZN(new_n19679_));
  AOI21_X1   g17243(.A1(new_n19678_), .A2(new_n19679_), .B(new_n12785_), .ZN(new_n19680_));
  NOR2_X1    g17244(.A1(new_n19680_), .A2(new_n12779_), .ZN(new_n19681_));
  AND2_X2    g17245(.A1(new_n19681_), .A2(new_n19677_), .Z(new_n19682_));
  NOR2_X1    g17246(.A1(new_n19682_), .A2(new_n19674_), .ZN(new_n19683_));
  NAND2_X1   g17247(.A1(new_n19683_), .A2(new_n12793_), .ZN(new_n19684_));
  NOR2_X1    g17248(.A1(new_n19646_), .A2(new_n12793_), .ZN(new_n19685_));
  INV_X1     g17249(.I(new_n19685_), .ZN(new_n19686_));
  AOI21_X1   g17250(.A1(new_n19684_), .A2(new_n19686_), .B(pi1159), .ZN(new_n19687_));
  NOR3_X1    g17251(.A1(new_n19682_), .A2(new_n12793_), .A3(new_n19674_), .ZN(new_n19688_));
  NOR2_X1    g17252(.A1(new_n19646_), .A2(pi0619), .ZN(new_n19689_));
  OAI21_X1   g17253(.A1(new_n19688_), .A2(new_n19689_), .B(pi1159), .ZN(new_n19690_));
  NAND2_X1   g17254(.A1(new_n19690_), .A2(pi0789), .ZN(new_n19691_));
  OAI22_X1   g17255(.A1(new_n19691_), .A2(new_n19687_), .B1(pi0789), .B2(new_n19683_), .ZN(new_n19692_));
  NAND2_X1   g17256(.A1(new_n19645_), .A2(new_n12818_), .ZN(new_n19693_));
  OAI21_X1   g17257(.A1(new_n19692_), .A2(new_n12818_), .B(new_n19693_), .ZN(new_n19694_));
  AOI21_X1   g17258(.A1(new_n19694_), .A2(new_n13384_), .B(new_n19649_), .ZN(new_n19695_));
  OAI21_X1   g17259(.A1(new_n19695_), .A2(new_n12984_), .B(new_n19648_), .ZN(new_n19696_));
  OAI21_X1   g17260(.A1(new_n19696_), .A2(pi0644), .B(new_n19647_), .ZN(new_n19697_));
  OAI21_X1   g17261(.A1(new_n14125_), .A2(new_n19659_), .B(new_n16558_), .ZN(new_n19698_));
  OAI21_X1   g17262(.A1(new_n14122_), .A2(new_n5657_), .B(new_n3265_), .ZN(new_n19699_));
  NAND2_X1   g17263(.A1(new_n19699_), .A2(new_n2609_), .ZN(new_n19700_));
  NAND2_X1   g17264(.A1(new_n15744_), .A2(new_n5657_), .ZN(new_n19701_));
  AOI21_X1   g17265(.A1(new_n19701_), .A2(new_n19700_), .B(new_n19698_), .ZN(new_n19702_));
  NAND2_X1   g17266(.A1(new_n2609_), .A2(new_n16558_), .ZN(new_n19703_));
  AOI21_X1   g17267(.A1(new_n19646_), .A2(new_n19703_), .B(new_n19702_), .ZN(new_n19704_));
  NAND2_X1   g17268(.A1(new_n19704_), .A2(new_n13521_), .ZN(new_n19705_));
  NAND2_X1   g17269(.A1(new_n19645_), .A2(pi0625), .ZN(new_n19706_));
  AOI21_X1   g17270(.A1(new_n19705_), .A2(new_n19706_), .B(pi1153), .ZN(new_n19707_));
  NAND2_X1   g17271(.A1(new_n19645_), .A2(new_n13521_), .ZN(new_n19708_));
  NAND2_X1   g17272(.A1(new_n19704_), .A2(pi0625), .ZN(new_n19709_));
  AOI21_X1   g17273(.A1(new_n19709_), .A2(new_n19708_), .B(new_n12841_), .ZN(new_n19710_));
  NOR3_X1    g17274(.A1(new_n19707_), .A2(new_n19710_), .A3(new_n12758_), .ZN(new_n19711_));
  NOR2_X1    g17275(.A1(new_n19704_), .A2(pi0778), .ZN(new_n19712_));
  NOR2_X1    g17276(.A1(new_n19711_), .A2(new_n19712_), .ZN(new_n19713_));
  NOR2_X1    g17277(.A1(new_n19713_), .A2(new_n12869_), .ZN(new_n19714_));
  AOI21_X1   g17278(.A1(new_n12869_), .A2(new_n19646_), .B(new_n19714_), .ZN(new_n19715_));
  NAND2_X1   g17279(.A1(new_n19715_), .A2(new_n12888_), .ZN(new_n19716_));
  OAI21_X1   g17280(.A1(new_n12888_), .A2(new_n19646_), .B(new_n19716_), .ZN(new_n19717_));
  INV_X1     g17281(.I(new_n19717_), .ZN(new_n19718_));
  NOR2_X1    g17282(.A1(new_n19645_), .A2(new_n12911_), .ZN(new_n19719_));
  AOI21_X1   g17283(.A1(new_n19718_), .A2(new_n12911_), .B(new_n19719_), .ZN(new_n19720_));
  NAND2_X1   g17284(.A1(new_n19720_), .A2(new_n13392_), .ZN(new_n19721_));
  OAI21_X1   g17285(.A1(new_n13392_), .A2(new_n19646_), .B(new_n19721_), .ZN(new_n19722_));
  NAND2_X1   g17286(.A1(new_n19722_), .A2(new_n12920_), .ZN(new_n19723_));
  NAND2_X1   g17287(.A1(new_n19645_), .A2(pi0628), .ZN(new_n19724_));
  AOI21_X1   g17288(.A1(new_n19723_), .A2(new_n19724_), .B(pi1156), .ZN(new_n19725_));
  NAND2_X1   g17289(.A1(new_n19645_), .A2(new_n12920_), .ZN(new_n19726_));
  NAND2_X1   g17290(.A1(new_n19722_), .A2(pi0628), .ZN(new_n19727_));
  AOI21_X1   g17291(.A1(new_n19727_), .A2(new_n19726_), .B(new_n12742_), .ZN(new_n19728_));
  OR2_X2     g17292(.A1(new_n19728_), .A2(new_n12937_), .Z(new_n19729_));
  OAI22_X1   g17293(.A1(new_n19729_), .A2(new_n19725_), .B1(pi0792), .B2(new_n19722_), .ZN(new_n19730_));
  NAND2_X1   g17294(.A1(new_n19730_), .A2(new_n12741_), .ZN(new_n19731_));
  OAI21_X1   g17295(.A1(new_n12741_), .A2(new_n19645_), .B(new_n19731_), .ZN(new_n19732_));
  NOR2_X1    g17296(.A1(new_n19732_), .A2(pi1157), .ZN(new_n19733_));
  NAND2_X1   g17297(.A1(new_n19730_), .A2(pi0647), .ZN(new_n19734_));
  OAI21_X1   g17298(.A1(pi0647), .A2(new_n19645_), .B(new_n19734_), .ZN(new_n19735_));
  NOR2_X1    g17299(.A1(new_n19735_), .A2(new_n12965_), .ZN(new_n19736_));
  OAI21_X1   g17300(.A1(new_n19733_), .A2(new_n19736_), .B(pi0787), .ZN(new_n19737_));
  OAI21_X1   g17301(.A1(pi0787), .A2(new_n19730_), .B(new_n19737_), .ZN(new_n19738_));
  OAI21_X1   g17302(.A1(new_n19738_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n19739_));
  NAND3_X1   g17303(.A1(new_n19739_), .A2(new_n12739_), .A3(new_n19697_), .ZN(new_n19740_));
  AOI21_X1   g17304(.A1(new_n19646_), .A2(new_n12975_), .B(pi0715), .ZN(new_n19741_));
  OAI21_X1   g17305(.A1(new_n19696_), .A2(new_n12975_), .B(new_n19741_), .ZN(new_n19742_));
  OAI21_X1   g17306(.A1(new_n19738_), .A2(pi0644), .B(pi0715), .ZN(new_n19743_));
  NAND3_X1   g17307(.A1(new_n19743_), .A2(pi1160), .A3(new_n19742_), .ZN(new_n19744_));
  AOI21_X1   g17308(.A1(new_n19740_), .A2(new_n19744_), .B(new_n13000_), .ZN(new_n19745_));
  NAND2_X1   g17309(.A1(new_n19646_), .A2(pi0626), .ZN(new_n19746_));
  NAND2_X1   g17310(.A1(new_n19692_), .A2(new_n12747_), .ZN(new_n19747_));
  AOI21_X1   g17311(.A1(new_n19747_), .A2(new_n19746_), .B(new_n12816_), .ZN(new_n19748_));
  NOR2_X1    g17312(.A1(new_n19645_), .A2(pi0626), .ZN(new_n19749_));
  AOI21_X1   g17313(.A1(new_n19692_), .A2(pi0626), .B(new_n19749_), .ZN(new_n19750_));
  OAI22_X1   g17314(.A1(new_n19750_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n19720_), .ZN(new_n19751_));
  OAI21_X1   g17315(.A1(new_n19751_), .A2(new_n19748_), .B(pi0788), .ZN(new_n19752_));
  NAND2_X1   g17316(.A1(new_n19752_), .A2(new_n15824_), .ZN(new_n19753_));
  NAND2_X1   g17317(.A1(new_n19713_), .A2(new_n12766_), .ZN(new_n19754_));
  AOI21_X1   g17318(.A1(new_n16550_), .A2(new_n13566_), .B(new_n15826_), .ZN(new_n19755_));
  AOI21_X1   g17319(.A1(new_n14328_), .A2(new_n19519_), .B(new_n5657_), .ZN(new_n19756_));
  AOI21_X1   g17320(.A1(new_n19756_), .A2(new_n5336_), .B(new_n3265_), .ZN(new_n19757_));
  OAI21_X1   g17321(.A1(new_n19755_), .A2(pi0180), .B(new_n19757_), .ZN(new_n19758_));
  NAND2_X1   g17322(.A1(new_n14172_), .A2(pi0180), .ZN(new_n19759_));
  NAND2_X1   g17323(.A1(new_n14174_), .A2(new_n5657_), .ZN(new_n19760_));
  AOI21_X1   g17324(.A1(new_n19759_), .A2(new_n19760_), .B(pi0753), .ZN(new_n19761_));
  NAND2_X1   g17325(.A1(new_n15835_), .A2(pi0180), .ZN(new_n19762_));
  NAND2_X1   g17326(.A1(new_n14177_), .A2(new_n5657_), .ZN(new_n19763_));
  AOI21_X1   g17327(.A1(new_n19763_), .A2(new_n19762_), .B(new_n16550_), .ZN(new_n19764_));
  OAI21_X1   g17328(.A1(new_n19764_), .A2(new_n19761_), .B(new_n2627_), .ZN(new_n19765_));
  NOR2_X1    g17329(.A1(new_n14182_), .A2(pi0180), .ZN(new_n19766_));
  NOR2_X1    g17330(.A1(new_n14184_), .A2(new_n5657_), .ZN(new_n19767_));
  OAI21_X1   g17331(.A1(new_n19766_), .A2(new_n19767_), .B(pi0753), .ZN(new_n19768_));
  NOR2_X1    g17332(.A1(new_n14187_), .A2(new_n5657_), .ZN(new_n19769_));
  NOR2_X1    g17333(.A1(new_n14189_), .A2(pi0180), .ZN(new_n19770_));
  OAI21_X1   g17334(.A1(new_n19769_), .A2(new_n19770_), .B(new_n16550_), .ZN(new_n19771_));
  NAND3_X1   g17335(.A1(new_n19771_), .A2(new_n19768_), .A3(pi0039), .ZN(new_n19772_));
  NAND3_X1   g17336(.A1(new_n19772_), .A2(new_n3265_), .A3(new_n19765_), .ZN(new_n19773_));
  NAND3_X1   g17337(.A1(new_n19773_), .A2(new_n16558_), .A3(new_n19758_), .ZN(new_n19774_));
  NAND2_X1   g17338(.A1(new_n19662_), .A2(pi0702), .ZN(new_n19775_));
  NAND3_X1   g17339(.A1(new_n19775_), .A2(new_n19774_), .A3(new_n2609_), .ZN(new_n19776_));
  AOI21_X1   g17340(.A1(new_n19776_), .A2(new_n19650_), .B(pi0778), .ZN(new_n19777_));
  INV_X1     g17341(.I(new_n19707_), .ZN(new_n19778_));
  NAND2_X1   g17342(.A1(new_n19663_), .A2(pi0625), .ZN(new_n19779_));
  NAND2_X1   g17343(.A1(new_n19776_), .A2(new_n19650_), .ZN(new_n19780_));
  NAND2_X1   g17344(.A1(new_n19780_), .A2(new_n13521_), .ZN(new_n19781_));
  NAND2_X1   g17345(.A1(new_n19781_), .A2(new_n19779_), .ZN(new_n19782_));
  AOI21_X1   g17346(.A1(new_n19782_), .A2(new_n12841_), .B(new_n19710_), .ZN(new_n19783_));
  NAND2_X1   g17347(.A1(new_n19663_), .A2(new_n13521_), .ZN(new_n19784_));
  NAND2_X1   g17348(.A1(new_n19780_), .A2(pi0625), .ZN(new_n19785_));
  NAND2_X1   g17349(.A1(new_n19785_), .A2(new_n19784_), .ZN(new_n19786_));
  AOI21_X1   g17350(.A1(new_n19786_), .A2(pi1153), .B(new_n13560_), .ZN(new_n19787_));
  AOI22_X1   g17351(.A1(new_n13560_), .A2(new_n19783_), .B1(new_n19787_), .B2(new_n19778_), .ZN(new_n19788_));
  AOI21_X1   g17352(.A1(new_n19788_), .A2(pi0778), .B(new_n19777_), .ZN(new_n19789_));
  OAI21_X1   g17353(.A1(new_n19789_), .A2(new_n12766_), .B(new_n19754_), .ZN(new_n19790_));
  AOI21_X1   g17354(.A1(new_n19790_), .A2(pi1155), .B(new_n19669_), .ZN(new_n19791_));
  NOR2_X1    g17355(.A1(new_n19789_), .A2(pi0609), .ZN(new_n19792_));
  NOR3_X1    g17356(.A1(new_n19711_), .A2(new_n12766_), .A3(new_n19712_), .ZN(new_n19793_));
  OAI21_X1   g17357(.A1(new_n19792_), .A2(new_n19793_), .B(new_n12770_), .ZN(new_n19794_));
  NOR2_X1    g17358(.A1(new_n19671_), .A2(pi0660), .ZN(new_n19795_));
  AOI22_X1   g17359(.A1(new_n19791_), .A2(pi0660), .B1(new_n19794_), .B2(new_n19795_), .ZN(new_n19796_));
  NOR2_X1    g17360(.A1(new_n19789_), .A2(pi0785), .ZN(new_n19797_));
  AOI21_X1   g17361(.A1(new_n19796_), .A2(pi0785), .B(new_n19797_), .ZN(new_n19798_));
  NOR2_X1    g17362(.A1(new_n19798_), .A2(pi0781), .ZN(new_n19799_));
  AND2_X2    g17363(.A1(new_n19715_), .A2(new_n12781_), .Z(new_n19800_));
  NOR2_X1    g17364(.A1(new_n19798_), .A2(new_n12781_), .ZN(new_n19801_));
  OAI21_X1   g17365(.A1(new_n19801_), .A2(new_n19800_), .B(pi1154), .ZN(new_n19802_));
  NAND3_X1   g17366(.A1(new_n19802_), .A2(pi0627), .A3(new_n19677_), .ZN(new_n19803_));
  NAND2_X1   g17367(.A1(new_n19715_), .A2(pi0618), .ZN(new_n19804_));
  OAI21_X1   g17368(.A1(new_n19798_), .A2(pi0618), .B(new_n19804_), .ZN(new_n19805_));
  AOI21_X1   g17369(.A1(new_n19805_), .A2(new_n12785_), .B(new_n19680_), .ZN(new_n19806_));
  AOI21_X1   g17370(.A1(new_n19806_), .A2(new_n12880_), .B(new_n12779_), .ZN(new_n19807_));
  AOI21_X1   g17371(.A1(new_n19807_), .A2(new_n19803_), .B(new_n19799_), .ZN(new_n19808_));
  OAI21_X1   g17372(.A1(new_n19808_), .A2(pi0789), .B(new_n12819_), .ZN(new_n19809_));
  NOR2_X1    g17373(.A1(new_n19718_), .A2(new_n12793_), .ZN(new_n19810_));
  NOR2_X1    g17374(.A1(new_n19808_), .A2(pi0619), .ZN(new_n19811_));
  OAI21_X1   g17375(.A1(new_n19811_), .A2(new_n19810_), .B(new_n12791_), .ZN(new_n19812_));
  NAND3_X1   g17376(.A1(new_n19812_), .A2(new_n12895_), .A3(new_n19690_), .ZN(new_n19813_));
  INV_X1     g17377(.I(new_n19687_), .ZN(new_n19814_));
  NAND2_X1   g17378(.A1(new_n19717_), .A2(new_n12793_), .ZN(new_n19815_));
  OAI21_X1   g17379(.A1(new_n19808_), .A2(new_n12793_), .B(new_n19815_), .ZN(new_n19816_));
  AOI21_X1   g17380(.A1(new_n19816_), .A2(pi1159), .B(new_n12895_), .ZN(new_n19817_));
  AOI21_X1   g17381(.A1(new_n19817_), .A2(new_n19814_), .B(new_n12796_), .ZN(new_n19818_));
  AOI21_X1   g17382(.A1(new_n19818_), .A2(new_n19813_), .B(new_n19809_), .ZN(new_n19819_));
  NOR2_X1    g17383(.A1(new_n19728_), .A2(pi0629), .ZN(new_n19820_));
  NOR2_X1    g17384(.A1(new_n19725_), .A2(new_n12919_), .ZN(new_n19821_));
  NOR2_X1    g17385(.A1(new_n19820_), .A2(new_n19821_), .ZN(new_n19822_));
  AOI21_X1   g17386(.A1(new_n19694_), .A2(new_n19160_), .B(new_n19822_), .ZN(new_n19823_));
  OAI22_X1   g17387(.A1(new_n19819_), .A2(new_n19753_), .B1(new_n12937_), .B2(new_n19823_), .ZN(new_n19824_));
  AOI21_X1   g17388(.A1(new_n19742_), .A2(pi1160), .B(new_n12975_), .ZN(new_n19825_));
  AOI21_X1   g17389(.A1(new_n19697_), .A2(new_n12739_), .B(pi0644), .ZN(new_n19826_));
  NOR2_X1    g17390(.A1(new_n19825_), .A2(new_n19826_), .ZN(new_n19827_));
  OAI22_X1   g17391(.A1(new_n15576_), .A2(new_n19735_), .B1(new_n19732_), .B2(new_n15730_), .ZN(new_n19828_));
  NOR2_X1    g17392(.A1(new_n19695_), .A2(new_n17212_), .ZN(new_n19829_));
  NOR2_X1    g17393(.A1(new_n19828_), .A2(new_n19829_), .ZN(new_n19830_));
  OAI22_X1   g17394(.A1(new_n19827_), .A2(new_n13000_), .B1(new_n19830_), .B2(new_n12972_), .ZN(new_n19831_));
  AOI21_X1   g17395(.A1(new_n19824_), .A2(new_n15693_), .B(new_n19831_), .ZN(new_n19832_));
  OAI21_X1   g17396(.A1(new_n19745_), .A2(new_n19832_), .B(new_n6643_), .ZN(new_n19833_));
  AOI22_X1   g17397(.A1(new_n19833_), .A2(new_n19644_), .B1(pi0832), .B2(new_n19643_), .ZN(po0337));
  NOR2_X1    g17398(.A1(new_n13340_), .A2(pi0754), .ZN(new_n19835_));
  NOR2_X1    g17399(.A1(new_n3042_), .A2(pi0181), .ZN(new_n19836_));
  NOR2_X1    g17400(.A1(new_n19835_), .A2(new_n19836_), .ZN(new_n19837_));
  NOR3_X1    g17401(.A1(new_n19837_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n19838_));
  INV_X1     g17402(.I(new_n19835_), .ZN(new_n19839_));
  NOR2_X1    g17403(.A1(new_n19839_), .A2(new_n13354_), .ZN(new_n19840_));
  NOR3_X1    g17404(.A1(new_n19840_), .A2(new_n12762_), .A3(new_n19837_), .ZN(new_n19841_));
  NOR2_X1    g17405(.A1(new_n19841_), .A2(new_n12770_), .ZN(new_n19842_));
  NOR3_X1    g17406(.A1(new_n19840_), .A2(pi1155), .A3(new_n19836_), .ZN(new_n19843_));
  NOR3_X1    g17407(.A1(new_n19842_), .A2(new_n12764_), .A3(new_n19843_), .ZN(new_n19844_));
  NOR2_X1    g17408(.A1(new_n19844_), .A2(new_n19838_), .ZN(new_n19845_));
  INV_X1     g17409(.I(new_n19845_), .ZN(new_n19846_));
  AOI21_X1   g17410(.A1(new_n19846_), .A2(new_n12783_), .B(pi1154), .ZN(new_n19847_));
  AOI21_X1   g17411(.A1(new_n19846_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n19848_));
  NOR3_X1    g17412(.A1(new_n19847_), .A2(new_n19848_), .A3(new_n12779_), .ZN(new_n19849_));
  AOI21_X1   g17413(.A1(new_n12779_), .A2(new_n19846_), .B(new_n19849_), .ZN(new_n19850_));
  OAI21_X1   g17414(.A1(new_n19850_), .A2(new_n17229_), .B(new_n12791_), .ZN(new_n19851_));
  OAI21_X1   g17415(.A1(new_n19850_), .A2(new_n17232_), .B(pi1159), .ZN(new_n19852_));
  NAND3_X1   g17416(.A1(new_n19851_), .A2(new_n19852_), .A3(pi0789), .ZN(new_n19853_));
  OAI21_X1   g17417(.A1(pi0789), .A2(new_n19850_), .B(new_n19853_), .ZN(new_n19854_));
  INV_X1     g17418(.I(new_n19836_), .ZN(new_n19855_));
  NAND2_X1   g17419(.A1(new_n12818_), .A2(new_n19855_), .ZN(new_n19856_));
  OAI21_X1   g17420(.A1(new_n19854_), .A2(new_n12818_), .B(new_n19856_), .ZN(new_n19857_));
  AOI21_X1   g17421(.A1(new_n12826_), .A2(new_n16593_), .B(new_n19836_), .ZN(new_n19858_));
  NOR2_X1    g17422(.A1(new_n19836_), .A2(pi1153), .ZN(new_n19859_));
  NOR2_X1    g17423(.A1(new_n12834_), .A2(pi0709), .ZN(new_n19860_));
  INV_X1     g17424(.I(new_n19860_), .ZN(new_n19861_));
  NAND2_X1   g17425(.A1(new_n19861_), .A2(new_n19859_), .ZN(new_n19862_));
  NOR2_X1    g17426(.A1(new_n19860_), .A2(new_n19858_), .ZN(new_n19863_));
  NOR2_X1    g17427(.A1(new_n19863_), .A2(new_n12841_), .ZN(new_n19864_));
  INV_X1     g17428(.I(new_n19864_), .ZN(new_n19865_));
  NAND3_X1   g17429(.A1(new_n19865_), .A2(pi0778), .A3(new_n19862_), .ZN(new_n19866_));
  OAI21_X1   g17430(.A1(pi0778), .A2(new_n19858_), .B(new_n19866_), .ZN(new_n19867_));
  NAND2_X1   g17431(.A1(new_n19867_), .A2(new_n17187_), .ZN(new_n19868_));
  NOR2_X1    g17432(.A1(new_n19868_), .A2(new_n12889_), .ZN(new_n19869_));
  NAND2_X1   g17433(.A1(new_n19869_), .A2(new_n18203_), .ZN(new_n19870_));
  NOR2_X1    g17434(.A1(new_n19870_), .A2(new_n17884_), .ZN(new_n19871_));
  INV_X1     g17435(.I(new_n19871_), .ZN(new_n19872_));
  OAI22_X1   g17436(.A1(new_n19857_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n19872_), .ZN(new_n19873_));
  AND2_X2    g17437(.A1(new_n19873_), .A2(new_n12919_), .Z(new_n19874_));
  OAI22_X1   g17438(.A1(new_n19857_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n19872_), .ZN(new_n19875_));
  AOI21_X1   g17439(.A1(pi0629), .A2(new_n19875_), .B(new_n19874_), .ZN(new_n19876_));
  INV_X1     g17440(.I(new_n19843_), .ZN(new_n19877_));
  NOR2_X1    g17441(.A1(new_n19858_), .A2(new_n12754_), .ZN(new_n19878_));
  NOR3_X1    g17442(.A1(new_n19878_), .A2(new_n19835_), .A3(new_n19836_), .ZN(new_n19879_));
  NAND2_X1   g17443(.A1(new_n19879_), .A2(new_n12758_), .ZN(new_n19880_));
  NAND2_X1   g17444(.A1(new_n19878_), .A2(pi0625), .ZN(new_n19881_));
  NAND3_X1   g17445(.A1(new_n19881_), .A2(pi1153), .A3(new_n19837_), .ZN(new_n19882_));
  NAND3_X1   g17446(.A1(new_n19862_), .A2(pi0608), .A3(new_n19882_), .ZN(new_n19883_));
  INV_X1     g17447(.I(new_n19881_), .ZN(new_n19884_));
  OAI21_X1   g17448(.A1(new_n19884_), .A2(new_n19879_), .B(new_n19859_), .ZN(new_n19885_));
  NAND3_X1   g17449(.A1(new_n19865_), .A2(new_n13560_), .A3(new_n19885_), .ZN(new_n19886_));
  NAND3_X1   g17450(.A1(new_n19886_), .A2(pi0778), .A3(new_n19883_), .ZN(new_n19887_));
  AOI21_X1   g17451(.A1(new_n19887_), .A2(new_n19880_), .B(new_n12766_), .ZN(new_n19888_));
  NOR2_X1    g17452(.A1(new_n19867_), .A2(pi0609), .ZN(new_n19889_));
  OAI21_X1   g17453(.A1(new_n19889_), .A2(new_n19888_), .B(pi1155), .ZN(new_n19890_));
  NAND3_X1   g17454(.A1(new_n19890_), .A2(pi0660), .A3(new_n19877_), .ZN(new_n19891_));
  NAND2_X1   g17455(.A1(new_n19887_), .A2(new_n19880_), .ZN(new_n19892_));
  NOR2_X1    g17456(.A1(new_n19867_), .A2(new_n12766_), .ZN(new_n19893_));
  AOI21_X1   g17457(.A1(new_n19892_), .A2(new_n12766_), .B(new_n19893_), .ZN(new_n19894_));
  NOR2_X1    g17458(.A1(new_n19842_), .A2(pi0660), .ZN(new_n19895_));
  OAI21_X1   g17459(.A1(new_n19894_), .A2(pi1155), .B(new_n19895_), .ZN(new_n19896_));
  NAND3_X1   g17460(.A1(new_n19896_), .A2(new_n19891_), .A3(pi0785), .ZN(new_n19897_));
  NAND2_X1   g17461(.A1(new_n19892_), .A2(new_n12764_), .ZN(new_n19898_));
  NAND2_X1   g17462(.A1(new_n19897_), .A2(new_n19898_), .ZN(new_n19899_));
  NAND2_X1   g17463(.A1(new_n19899_), .A2(new_n12781_), .ZN(new_n19900_));
  NAND2_X1   g17464(.A1(new_n19868_), .A2(pi0618), .ZN(new_n19901_));
  AOI21_X1   g17465(.A1(new_n19900_), .A2(new_n19901_), .B(pi1154), .ZN(new_n19902_));
  NOR3_X1    g17466(.A1(new_n19902_), .A2(pi0627), .A3(new_n19848_), .ZN(new_n19903_));
  NAND2_X1   g17467(.A1(new_n19868_), .A2(new_n12781_), .ZN(new_n19904_));
  NAND2_X1   g17468(.A1(new_n19899_), .A2(pi0618), .ZN(new_n19905_));
  AOI21_X1   g17469(.A1(new_n19905_), .A2(new_n19904_), .B(new_n12785_), .ZN(new_n19906_));
  NOR3_X1    g17470(.A1(new_n19906_), .A2(new_n12880_), .A3(new_n19847_), .ZN(new_n19907_));
  OR3_X2     g17471(.A1(new_n19903_), .A2(new_n19907_), .A3(new_n12779_), .Z(new_n19908_));
  NAND2_X1   g17472(.A1(new_n19899_), .A2(new_n12779_), .ZN(new_n19909_));
  NAND2_X1   g17473(.A1(new_n19908_), .A2(new_n19909_), .ZN(new_n19910_));
  AOI21_X1   g17474(.A1(new_n19910_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n19911_));
  NOR2_X1    g17475(.A1(new_n19869_), .A2(pi0619), .ZN(new_n19912_));
  AOI21_X1   g17476(.A1(new_n19908_), .A2(new_n19909_), .B(new_n12793_), .ZN(new_n19913_));
  OAI21_X1   g17477(.A1(new_n19913_), .A2(new_n19912_), .B(pi1159), .ZN(new_n19914_));
  NAND3_X1   g17478(.A1(new_n19914_), .A2(pi0648), .A3(new_n19851_), .ZN(new_n19915_));
  NAND2_X1   g17479(.A1(new_n19910_), .A2(new_n12793_), .ZN(new_n19916_));
  OAI21_X1   g17480(.A1(new_n12793_), .A2(new_n19869_), .B(new_n19916_), .ZN(new_n19917_));
  NAND2_X1   g17481(.A1(new_n19917_), .A2(new_n12791_), .ZN(new_n19918_));
  NAND3_X1   g17482(.A1(new_n19918_), .A2(new_n12895_), .A3(new_n19852_), .ZN(new_n19919_));
  NAND3_X1   g17483(.A1(new_n19919_), .A2(pi0789), .A3(new_n19915_), .ZN(new_n19920_));
  NOR2_X1    g17484(.A1(new_n19855_), .A2(new_n12747_), .ZN(new_n19921_));
  AND2_X2    g17485(.A1(new_n19854_), .A2(new_n12747_), .Z(new_n19922_));
  OAI21_X1   g17486(.A1(new_n19922_), .A2(new_n19921_), .B(new_n12815_), .ZN(new_n19923_));
  INV_X1     g17487(.I(new_n19870_), .ZN(new_n19924_));
  NAND2_X1   g17488(.A1(new_n19854_), .A2(pi0626), .ZN(new_n19925_));
  OAI21_X1   g17489(.A1(pi0626), .A2(new_n19855_), .B(new_n19925_), .ZN(new_n19926_));
  AOI22_X1   g17490(.A1(new_n19926_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n19924_), .ZN(new_n19927_));
  NAND2_X1   g17491(.A1(new_n19927_), .A2(new_n19923_), .ZN(new_n19928_));
  AOI22_X1   g17492(.A1(new_n19920_), .A2(new_n19911_), .B1(pi0788), .B2(new_n19928_), .ZN(new_n19929_));
  OAI22_X1   g17493(.A1(new_n19929_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n19876_), .ZN(new_n19930_));
  NAND2_X1   g17494(.A1(new_n19857_), .A2(new_n13384_), .ZN(new_n19931_));
  NAND2_X1   g17495(.A1(new_n12943_), .A2(new_n19855_), .ZN(new_n19932_));
  NAND2_X1   g17496(.A1(new_n19931_), .A2(new_n19932_), .ZN(new_n19933_));
  NOR2_X1    g17497(.A1(new_n19872_), .A2(new_n12953_), .ZN(new_n19934_));
  NOR2_X1    g17498(.A1(new_n19934_), .A2(pi0647), .ZN(new_n19935_));
  NOR2_X1    g17499(.A1(new_n19836_), .A2(new_n12741_), .ZN(new_n19936_));
  OAI21_X1   g17500(.A1(new_n19935_), .A2(new_n19936_), .B(new_n12965_), .ZN(new_n19937_));
  NAND2_X1   g17501(.A1(new_n19934_), .A2(pi0647), .ZN(new_n19938_));
  OAI21_X1   g17502(.A1(pi0647), .A2(new_n19855_), .B(new_n19938_), .ZN(new_n19939_));
  OAI22_X1   g17503(.A1(new_n19939_), .A2(new_n15576_), .B1(new_n19937_), .B2(new_n12981_), .ZN(new_n19940_));
  AOI21_X1   g17504(.A1(new_n19933_), .A2(new_n15608_), .B(new_n19940_), .ZN(new_n19941_));
  OAI22_X1   g17505(.A1(new_n19930_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n19941_), .ZN(new_n19942_));
  NAND2_X1   g17506(.A1(new_n19942_), .A2(new_n13000_), .ZN(new_n19943_));
  AND2_X2    g17507(.A1(new_n19942_), .A2(new_n12975_), .Z(new_n19944_));
  OAI21_X1   g17508(.A1(new_n19939_), .A2(new_n12965_), .B(new_n19937_), .ZN(new_n19945_));
  NAND2_X1   g17509(.A1(new_n19934_), .A2(new_n12972_), .ZN(new_n19946_));
  OAI21_X1   g17510(.A1(new_n19945_), .A2(new_n12972_), .B(new_n19946_), .ZN(new_n19947_));
  NOR2_X1    g17511(.A1(new_n19947_), .A2(new_n12975_), .ZN(new_n19948_));
  OAI21_X1   g17512(.A1(new_n19944_), .A2(new_n19948_), .B(new_n12740_), .ZN(new_n19949_));
  NAND2_X1   g17513(.A1(new_n19855_), .A2(pi0644), .ZN(new_n19950_));
  NOR2_X1    g17514(.A1(new_n17611_), .A2(new_n19836_), .ZN(new_n19951_));
  AOI21_X1   g17515(.A1(new_n19857_), .A2(new_n17611_), .B(new_n19951_), .ZN(new_n19952_));
  OAI21_X1   g17516(.A1(new_n19952_), .A2(pi0644), .B(new_n19950_), .ZN(new_n19953_));
  NAND2_X1   g17517(.A1(new_n19953_), .A2(pi0715), .ZN(new_n19954_));
  NAND3_X1   g17518(.A1(new_n19949_), .A2(new_n12739_), .A3(new_n19954_), .ZN(new_n19955_));
  NOR2_X1    g17519(.A1(new_n19947_), .A2(pi0644), .ZN(new_n19956_));
  AOI21_X1   g17520(.A1(new_n19942_), .A2(pi0644), .B(new_n19956_), .ZN(new_n19957_));
  NAND2_X1   g17521(.A1(new_n19855_), .A2(new_n12975_), .ZN(new_n19958_));
  OAI21_X1   g17522(.A1(new_n19952_), .A2(new_n12975_), .B(new_n19958_), .ZN(new_n19959_));
  AOI21_X1   g17523(.A1(new_n19959_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n19960_));
  OAI21_X1   g17524(.A1(new_n19957_), .A2(new_n12740_), .B(new_n19960_), .ZN(new_n19961_));
  NAND3_X1   g17525(.A1(new_n19955_), .A2(pi0790), .A3(new_n19961_), .ZN(new_n19962_));
  NAND2_X1   g17526(.A1(new_n19962_), .A2(new_n19943_), .ZN(new_n19963_));
  AOI21_X1   g17527(.A1(po1038), .A2(new_n5658_), .B(pi0832), .ZN(new_n19964_));
  NAND2_X1   g17528(.A1(new_n13192_), .A2(new_n5658_), .ZN(new_n19965_));
  INV_X1     g17529(.I(new_n19965_), .ZN(new_n19966_));
  AOI21_X1   g17530(.A1(new_n19966_), .A2(pi0644), .B(new_n12740_), .ZN(new_n19967_));
  NAND2_X1   g17531(.A1(new_n19965_), .A2(new_n12984_), .ZN(new_n19968_));
  NOR2_X1    g17532(.A1(new_n19966_), .A2(new_n13384_), .ZN(new_n19969_));
  NAND2_X1   g17533(.A1(new_n2610_), .A2(pi0181), .ZN(new_n19970_));
  OAI22_X1   g17534(.A1(new_n19651_), .A2(new_n5658_), .B1(new_n16585_), .B2(new_n13060_), .ZN(new_n19971_));
  NAND2_X1   g17535(.A1(new_n5658_), .A2(pi0754), .ZN(new_n19972_));
  OAI21_X1   g17536(.A1(new_n13334_), .A2(pi0181), .B(new_n16585_), .ZN(new_n19973_));
  AOI22_X1   g17537(.A1(new_n19973_), .A2(new_n19972_), .B1(new_n2627_), .B2(new_n19971_), .ZN(new_n19974_));
  OAI22_X1   g17538(.A1(new_n14065_), .A2(new_n16585_), .B1(new_n5658_), .B2(new_n14067_), .ZN(new_n19975_));
  NAND2_X1   g17539(.A1(new_n19975_), .A2(pi0039), .ZN(new_n19976_));
  NAND2_X1   g17540(.A1(new_n19974_), .A2(new_n19976_), .ZN(new_n19977_));
  NOR2_X1    g17541(.A1(new_n13344_), .A2(pi0181), .ZN(new_n19978_));
  NOR2_X1    g17542(.A1(new_n19978_), .A2(new_n3265_), .ZN(new_n19979_));
  NAND2_X1   g17543(.A1(new_n13341_), .A2(new_n16585_), .ZN(new_n19980_));
  AOI22_X1   g17544(.A1(new_n19977_), .A2(new_n3265_), .B1(new_n19979_), .B2(new_n19980_), .ZN(new_n19981_));
  OAI21_X1   g17545(.A1(new_n19981_), .A2(new_n2610_), .B(new_n19970_), .ZN(new_n19982_));
  NAND2_X1   g17546(.A1(new_n19982_), .A2(new_n12761_), .ZN(new_n19983_));
  INV_X1     g17547(.I(new_n19983_), .ZN(new_n19984_));
  NOR2_X1    g17548(.A1(new_n19966_), .A2(new_n12761_), .ZN(new_n19985_));
  NOR3_X1    g17549(.A1(new_n19984_), .A2(pi0785), .A3(new_n19985_), .ZN(new_n19986_));
  AOI22_X1   g17550(.A1(new_n19984_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n19965_), .ZN(new_n19987_));
  NOR2_X1    g17551(.A1(new_n19987_), .A2(pi1155), .ZN(new_n19988_));
  AOI22_X1   g17552(.A1(new_n19984_), .A2(pi0609), .B1(new_n13357_), .B2(new_n19965_), .ZN(new_n19989_));
  NOR2_X1    g17553(.A1(new_n19989_), .A2(new_n12770_), .ZN(new_n19990_));
  NOR3_X1    g17554(.A1(new_n19990_), .A2(new_n19988_), .A3(new_n12764_), .ZN(new_n19991_));
  NOR2_X1    g17555(.A1(new_n19991_), .A2(new_n19986_), .ZN(new_n19992_));
  NOR2_X1    g17556(.A1(new_n19992_), .A2(pi0781), .ZN(new_n19993_));
  NOR3_X1    g17557(.A1(new_n19991_), .A2(pi0618), .A3(new_n19986_), .ZN(new_n19994_));
  NOR2_X1    g17558(.A1(new_n19966_), .A2(new_n12781_), .ZN(new_n19995_));
  OAI21_X1   g17559(.A1(new_n19994_), .A2(new_n19995_), .B(new_n12785_), .ZN(new_n19996_));
  NAND2_X1   g17560(.A1(new_n19992_), .A2(pi0618), .ZN(new_n19997_));
  NAND2_X1   g17561(.A1(new_n19965_), .A2(new_n12781_), .ZN(new_n19998_));
  AOI21_X1   g17562(.A1(new_n19997_), .A2(new_n19998_), .B(new_n12785_), .ZN(new_n19999_));
  NOR2_X1    g17563(.A1(new_n19999_), .A2(new_n12779_), .ZN(new_n20000_));
  AND2_X2    g17564(.A1(new_n20000_), .A2(new_n19996_), .Z(new_n20001_));
  NOR2_X1    g17565(.A1(new_n20001_), .A2(new_n19993_), .ZN(new_n20002_));
  NAND2_X1   g17566(.A1(new_n20002_), .A2(new_n12793_), .ZN(new_n20003_));
  NOR2_X1    g17567(.A1(new_n19966_), .A2(new_n12793_), .ZN(new_n20004_));
  INV_X1     g17568(.I(new_n20004_), .ZN(new_n20005_));
  AOI21_X1   g17569(.A1(new_n20003_), .A2(new_n20005_), .B(pi1159), .ZN(new_n20006_));
  NOR3_X1    g17570(.A1(new_n20001_), .A2(new_n12793_), .A3(new_n19993_), .ZN(new_n20007_));
  NOR2_X1    g17571(.A1(new_n19966_), .A2(pi0619), .ZN(new_n20008_));
  OAI21_X1   g17572(.A1(new_n20007_), .A2(new_n20008_), .B(pi1159), .ZN(new_n20009_));
  NAND2_X1   g17573(.A1(new_n20009_), .A2(pi0789), .ZN(new_n20010_));
  OAI22_X1   g17574(.A1(new_n20010_), .A2(new_n20006_), .B1(pi0789), .B2(new_n20002_), .ZN(new_n20011_));
  NAND2_X1   g17575(.A1(new_n19965_), .A2(new_n12818_), .ZN(new_n20012_));
  OAI21_X1   g17576(.A1(new_n20011_), .A2(new_n12818_), .B(new_n20012_), .ZN(new_n20013_));
  AOI21_X1   g17577(.A1(new_n20013_), .A2(new_n13384_), .B(new_n19969_), .ZN(new_n20014_));
  OAI21_X1   g17578(.A1(new_n20014_), .A2(new_n12984_), .B(new_n19968_), .ZN(new_n20015_));
  OAI21_X1   g17579(.A1(new_n20015_), .A2(pi0644), .B(new_n19967_), .ZN(new_n20016_));
  OAI21_X1   g17580(.A1(new_n14125_), .A2(new_n19978_), .B(new_n16593_), .ZN(new_n20017_));
  OAI21_X1   g17581(.A1(new_n14122_), .A2(new_n5658_), .B(new_n3265_), .ZN(new_n20018_));
  NAND2_X1   g17582(.A1(new_n20018_), .A2(new_n2609_), .ZN(new_n20019_));
  NAND2_X1   g17583(.A1(new_n15744_), .A2(new_n5658_), .ZN(new_n20020_));
  AOI21_X1   g17584(.A1(new_n20020_), .A2(new_n20019_), .B(new_n20017_), .ZN(new_n20021_));
  NAND2_X1   g17585(.A1(new_n2609_), .A2(new_n16593_), .ZN(new_n20022_));
  AOI21_X1   g17586(.A1(new_n19966_), .A2(new_n20022_), .B(new_n20021_), .ZN(new_n20023_));
  NAND2_X1   g17587(.A1(new_n20023_), .A2(new_n13521_), .ZN(new_n20024_));
  NAND2_X1   g17588(.A1(new_n19965_), .A2(pi0625), .ZN(new_n20025_));
  AOI21_X1   g17589(.A1(new_n20024_), .A2(new_n20025_), .B(pi1153), .ZN(new_n20026_));
  NAND2_X1   g17590(.A1(new_n19965_), .A2(new_n13521_), .ZN(new_n20027_));
  NAND2_X1   g17591(.A1(new_n20023_), .A2(pi0625), .ZN(new_n20028_));
  AOI21_X1   g17592(.A1(new_n20028_), .A2(new_n20027_), .B(new_n12841_), .ZN(new_n20029_));
  NOR3_X1    g17593(.A1(new_n20026_), .A2(new_n20029_), .A3(new_n12758_), .ZN(new_n20030_));
  NOR2_X1    g17594(.A1(new_n20023_), .A2(pi0778), .ZN(new_n20031_));
  NOR2_X1    g17595(.A1(new_n20030_), .A2(new_n20031_), .ZN(new_n20032_));
  NOR2_X1    g17596(.A1(new_n20032_), .A2(new_n12869_), .ZN(new_n20033_));
  AOI21_X1   g17597(.A1(new_n12869_), .A2(new_n19966_), .B(new_n20033_), .ZN(new_n20034_));
  NAND2_X1   g17598(.A1(new_n20034_), .A2(new_n12888_), .ZN(new_n20035_));
  OAI21_X1   g17599(.A1(new_n12888_), .A2(new_n19966_), .B(new_n20035_), .ZN(new_n20036_));
  INV_X1     g17600(.I(new_n20036_), .ZN(new_n20037_));
  NOR2_X1    g17601(.A1(new_n19965_), .A2(new_n12911_), .ZN(new_n20038_));
  AOI21_X1   g17602(.A1(new_n20037_), .A2(new_n12911_), .B(new_n20038_), .ZN(new_n20039_));
  NAND2_X1   g17603(.A1(new_n20039_), .A2(new_n13392_), .ZN(new_n20040_));
  OAI21_X1   g17604(.A1(new_n13392_), .A2(new_n19966_), .B(new_n20040_), .ZN(new_n20041_));
  NAND2_X1   g17605(.A1(new_n20041_), .A2(new_n12920_), .ZN(new_n20042_));
  NAND2_X1   g17606(.A1(new_n19965_), .A2(pi0628), .ZN(new_n20043_));
  AOI21_X1   g17607(.A1(new_n20042_), .A2(new_n20043_), .B(pi1156), .ZN(new_n20044_));
  NAND2_X1   g17608(.A1(new_n19965_), .A2(new_n12920_), .ZN(new_n20045_));
  NAND2_X1   g17609(.A1(new_n20041_), .A2(pi0628), .ZN(new_n20046_));
  AOI21_X1   g17610(.A1(new_n20046_), .A2(new_n20045_), .B(new_n12742_), .ZN(new_n20047_));
  OR2_X2     g17611(.A1(new_n20047_), .A2(new_n12937_), .Z(new_n20048_));
  OAI22_X1   g17612(.A1(new_n20048_), .A2(new_n20044_), .B1(pi0792), .B2(new_n20041_), .ZN(new_n20049_));
  NAND2_X1   g17613(.A1(new_n20049_), .A2(new_n12741_), .ZN(new_n20050_));
  OAI21_X1   g17614(.A1(new_n12741_), .A2(new_n19965_), .B(new_n20050_), .ZN(new_n20051_));
  NOR2_X1    g17615(.A1(new_n20051_), .A2(pi1157), .ZN(new_n20052_));
  NAND2_X1   g17616(.A1(new_n20049_), .A2(pi0647), .ZN(new_n20053_));
  OAI21_X1   g17617(.A1(pi0647), .A2(new_n19965_), .B(new_n20053_), .ZN(new_n20054_));
  NOR2_X1    g17618(.A1(new_n20054_), .A2(new_n12965_), .ZN(new_n20055_));
  OAI21_X1   g17619(.A1(new_n20052_), .A2(new_n20055_), .B(pi0787), .ZN(new_n20056_));
  OAI21_X1   g17620(.A1(pi0787), .A2(new_n20049_), .B(new_n20056_), .ZN(new_n20057_));
  OAI21_X1   g17621(.A1(new_n20057_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n20058_));
  NAND3_X1   g17622(.A1(new_n20058_), .A2(new_n12739_), .A3(new_n20016_), .ZN(new_n20059_));
  AOI21_X1   g17623(.A1(new_n19966_), .A2(new_n12975_), .B(pi0715), .ZN(new_n20060_));
  OAI21_X1   g17624(.A1(new_n20015_), .A2(new_n12975_), .B(new_n20060_), .ZN(new_n20061_));
  OAI21_X1   g17625(.A1(new_n20057_), .A2(pi0644), .B(pi0715), .ZN(new_n20062_));
  NAND3_X1   g17626(.A1(new_n20062_), .A2(pi1160), .A3(new_n20061_), .ZN(new_n20063_));
  AOI21_X1   g17627(.A1(new_n20059_), .A2(new_n20063_), .B(new_n13000_), .ZN(new_n20064_));
  NAND2_X1   g17628(.A1(new_n19966_), .A2(pi0626), .ZN(new_n20065_));
  NAND2_X1   g17629(.A1(new_n20011_), .A2(new_n12747_), .ZN(new_n20066_));
  AOI21_X1   g17630(.A1(new_n20066_), .A2(new_n20065_), .B(new_n12816_), .ZN(new_n20067_));
  NOR2_X1    g17631(.A1(new_n19965_), .A2(pi0626), .ZN(new_n20068_));
  AOI21_X1   g17632(.A1(new_n20011_), .A2(pi0626), .B(new_n20068_), .ZN(new_n20069_));
  OAI22_X1   g17633(.A1(new_n20069_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n20039_), .ZN(new_n20070_));
  OAI21_X1   g17634(.A1(new_n20070_), .A2(new_n20067_), .B(pi0788), .ZN(new_n20071_));
  NAND2_X1   g17635(.A1(new_n20071_), .A2(new_n15824_), .ZN(new_n20072_));
  NAND2_X1   g17636(.A1(new_n20032_), .A2(new_n12766_), .ZN(new_n20073_));
  AOI21_X1   g17637(.A1(new_n16585_), .A2(new_n13566_), .B(new_n15826_), .ZN(new_n20074_));
  AOI21_X1   g17638(.A1(new_n14328_), .A2(new_n19839_), .B(new_n5658_), .ZN(new_n20075_));
  AOI21_X1   g17639(.A1(new_n20075_), .A2(new_n5336_), .B(new_n3265_), .ZN(new_n20076_));
  OAI21_X1   g17640(.A1(new_n20074_), .A2(pi0181), .B(new_n20076_), .ZN(new_n20077_));
  NAND2_X1   g17641(.A1(new_n14172_), .A2(pi0181), .ZN(new_n20078_));
  NAND2_X1   g17642(.A1(new_n14174_), .A2(new_n5658_), .ZN(new_n20079_));
  AOI21_X1   g17643(.A1(new_n20078_), .A2(new_n20079_), .B(pi0754), .ZN(new_n20080_));
  NAND2_X1   g17644(.A1(new_n15835_), .A2(pi0181), .ZN(new_n20081_));
  NAND2_X1   g17645(.A1(new_n14177_), .A2(new_n5658_), .ZN(new_n20082_));
  AOI21_X1   g17646(.A1(new_n20082_), .A2(new_n20081_), .B(new_n16585_), .ZN(new_n20083_));
  OAI21_X1   g17647(.A1(new_n20083_), .A2(new_n20080_), .B(new_n2627_), .ZN(new_n20084_));
  NOR2_X1    g17648(.A1(new_n14182_), .A2(pi0181), .ZN(new_n20085_));
  NOR2_X1    g17649(.A1(new_n14184_), .A2(new_n5658_), .ZN(new_n20086_));
  OAI21_X1   g17650(.A1(new_n20085_), .A2(new_n20086_), .B(pi0754), .ZN(new_n20087_));
  NOR2_X1    g17651(.A1(new_n14187_), .A2(new_n5658_), .ZN(new_n20088_));
  NOR2_X1    g17652(.A1(new_n14189_), .A2(pi0181), .ZN(new_n20089_));
  OAI21_X1   g17653(.A1(new_n20088_), .A2(new_n20089_), .B(new_n16585_), .ZN(new_n20090_));
  NAND3_X1   g17654(.A1(new_n20090_), .A2(new_n20087_), .A3(pi0039), .ZN(new_n20091_));
  NAND3_X1   g17655(.A1(new_n20091_), .A2(new_n3265_), .A3(new_n20084_), .ZN(new_n20092_));
  NAND3_X1   g17656(.A1(new_n20092_), .A2(new_n16593_), .A3(new_n20077_), .ZN(new_n20093_));
  NAND2_X1   g17657(.A1(new_n19981_), .A2(pi0709), .ZN(new_n20094_));
  NAND3_X1   g17658(.A1(new_n20094_), .A2(new_n20093_), .A3(new_n2609_), .ZN(new_n20095_));
  AOI21_X1   g17659(.A1(new_n20095_), .A2(new_n19970_), .B(pi0778), .ZN(new_n20096_));
  INV_X1     g17660(.I(new_n20026_), .ZN(new_n20097_));
  NAND2_X1   g17661(.A1(new_n19982_), .A2(pi0625), .ZN(new_n20098_));
  NAND2_X1   g17662(.A1(new_n20095_), .A2(new_n19970_), .ZN(new_n20099_));
  NAND2_X1   g17663(.A1(new_n20099_), .A2(new_n13521_), .ZN(new_n20100_));
  NAND2_X1   g17664(.A1(new_n20100_), .A2(new_n20098_), .ZN(new_n20101_));
  AOI21_X1   g17665(.A1(new_n20101_), .A2(new_n12841_), .B(new_n20029_), .ZN(new_n20102_));
  NAND2_X1   g17666(.A1(new_n19982_), .A2(new_n13521_), .ZN(new_n20103_));
  NAND2_X1   g17667(.A1(new_n20099_), .A2(pi0625), .ZN(new_n20104_));
  NAND2_X1   g17668(.A1(new_n20104_), .A2(new_n20103_), .ZN(new_n20105_));
  AOI21_X1   g17669(.A1(new_n20105_), .A2(pi1153), .B(new_n13560_), .ZN(new_n20106_));
  AOI22_X1   g17670(.A1(new_n13560_), .A2(new_n20102_), .B1(new_n20106_), .B2(new_n20097_), .ZN(new_n20107_));
  AOI21_X1   g17671(.A1(new_n20107_), .A2(pi0778), .B(new_n20096_), .ZN(new_n20108_));
  OAI21_X1   g17672(.A1(new_n20108_), .A2(new_n12766_), .B(new_n20073_), .ZN(new_n20109_));
  AOI21_X1   g17673(.A1(new_n20109_), .A2(pi1155), .B(new_n19988_), .ZN(new_n20110_));
  NOR2_X1    g17674(.A1(new_n20108_), .A2(pi0609), .ZN(new_n20111_));
  NOR3_X1    g17675(.A1(new_n20030_), .A2(new_n12766_), .A3(new_n20031_), .ZN(new_n20112_));
  OAI21_X1   g17676(.A1(new_n20111_), .A2(new_n20112_), .B(new_n12770_), .ZN(new_n20113_));
  NOR2_X1    g17677(.A1(new_n19990_), .A2(pi0660), .ZN(new_n20114_));
  AOI22_X1   g17678(.A1(new_n20110_), .A2(pi0660), .B1(new_n20113_), .B2(new_n20114_), .ZN(new_n20115_));
  NOR2_X1    g17679(.A1(new_n20108_), .A2(pi0785), .ZN(new_n20116_));
  AOI21_X1   g17680(.A1(new_n20115_), .A2(pi0785), .B(new_n20116_), .ZN(new_n20117_));
  NOR2_X1    g17681(.A1(new_n20117_), .A2(pi0781), .ZN(new_n20118_));
  AND2_X2    g17682(.A1(new_n20034_), .A2(new_n12781_), .Z(new_n20119_));
  NOR2_X1    g17683(.A1(new_n20117_), .A2(new_n12781_), .ZN(new_n20120_));
  OAI21_X1   g17684(.A1(new_n20120_), .A2(new_n20119_), .B(pi1154), .ZN(new_n20121_));
  NAND3_X1   g17685(.A1(new_n20121_), .A2(pi0627), .A3(new_n19996_), .ZN(new_n20122_));
  NAND2_X1   g17686(.A1(new_n20034_), .A2(pi0618), .ZN(new_n20123_));
  OAI21_X1   g17687(.A1(new_n20117_), .A2(pi0618), .B(new_n20123_), .ZN(new_n20124_));
  AOI21_X1   g17688(.A1(new_n20124_), .A2(new_n12785_), .B(new_n19999_), .ZN(new_n20125_));
  AOI21_X1   g17689(.A1(new_n20125_), .A2(new_n12880_), .B(new_n12779_), .ZN(new_n20126_));
  AOI21_X1   g17690(.A1(new_n20126_), .A2(new_n20122_), .B(new_n20118_), .ZN(new_n20127_));
  OAI21_X1   g17691(.A1(new_n20127_), .A2(pi0789), .B(new_n12819_), .ZN(new_n20128_));
  NOR2_X1    g17692(.A1(new_n20037_), .A2(new_n12793_), .ZN(new_n20129_));
  NOR2_X1    g17693(.A1(new_n20127_), .A2(pi0619), .ZN(new_n20130_));
  OAI21_X1   g17694(.A1(new_n20130_), .A2(new_n20129_), .B(new_n12791_), .ZN(new_n20131_));
  NAND3_X1   g17695(.A1(new_n20131_), .A2(new_n12895_), .A3(new_n20009_), .ZN(new_n20132_));
  INV_X1     g17696(.I(new_n20006_), .ZN(new_n20133_));
  NAND2_X1   g17697(.A1(new_n20036_), .A2(new_n12793_), .ZN(new_n20134_));
  OAI21_X1   g17698(.A1(new_n20127_), .A2(new_n12793_), .B(new_n20134_), .ZN(new_n20135_));
  AOI21_X1   g17699(.A1(new_n20135_), .A2(pi1159), .B(new_n12895_), .ZN(new_n20136_));
  AOI21_X1   g17700(.A1(new_n20136_), .A2(new_n20133_), .B(new_n12796_), .ZN(new_n20137_));
  AOI21_X1   g17701(.A1(new_n20137_), .A2(new_n20132_), .B(new_n20128_), .ZN(new_n20138_));
  NOR2_X1    g17702(.A1(new_n20047_), .A2(pi0629), .ZN(new_n20139_));
  NOR2_X1    g17703(.A1(new_n20044_), .A2(new_n12919_), .ZN(new_n20140_));
  NOR2_X1    g17704(.A1(new_n20139_), .A2(new_n20140_), .ZN(new_n20141_));
  AOI21_X1   g17705(.A1(new_n20013_), .A2(new_n19160_), .B(new_n20141_), .ZN(new_n20142_));
  OAI22_X1   g17706(.A1(new_n20138_), .A2(new_n20072_), .B1(new_n12937_), .B2(new_n20142_), .ZN(new_n20143_));
  AOI21_X1   g17707(.A1(new_n20061_), .A2(pi1160), .B(new_n12975_), .ZN(new_n20144_));
  AOI21_X1   g17708(.A1(new_n20016_), .A2(new_n12739_), .B(pi0644), .ZN(new_n20145_));
  NOR2_X1    g17709(.A1(new_n20144_), .A2(new_n20145_), .ZN(new_n20146_));
  OAI22_X1   g17710(.A1(new_n15576_), .A2(new_n20054_), .B1(new_n20051_), .B2(new_n15730_), .ZN(new_n20147_));
  NOR2_X1    g17711(.A1(new_n20014_), .A2(new_n17212_), .ZN(new_n20148_));
  NOR2_X1    g17712(.A1(new_n20147_), .A2(new_n20148_), .ZN(new_n20149_));
  OAI22_X1   g17713(.A1(new_n20146_), .A2(new_n13000_), .B1(new_n20149_), .B2(new_n12972_), .ZN(new_n20150_));
  AOI21_X1   g17714(.A1(new_n20143_), .A2(new_n15693_), .B(new_n20150_), .ZN(new_n20151_));
  OAI21_X1   g17715(.A1(new_n20064_), .A2(new_n20151_), .B(new_n6643_), .ZN(new_n20152_));
  AOI22_X1   g17716(.A1(new_n20152_), .A2(new_n19964_), .B1(pi0832), .B2(new_n19963_), .ZN(po0338));
  NOR2_X1    g17717(.A1(new_n13340_), .A2(pi0756), .ZN(new_n20154_));
  NOR2_X1    g17718(.A1(new_n3042_), .A2(pi0182), .ZN(new_n20155_));
  NOR2_X1    g17719(.A1(new_n20154_), .A2(new_n20155_), .ZN(new_n20156_));
  NOR3_X1    g17720(.A1(new_n20156_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n20157_));
  INV_X1     g17721(.I(new_n20154_), .ZN(new_n20158_));
  NOR2_X1    g17722(.A1(new_n20158_), .A2(new_n13354_), .ZN(new_n20159_));
  NOR3_X1    g17723(.A1(new_n20159_), .A2(new_n12762_), .A3(new_n20156_), .ZN(new_n20160_));
  NOR2_X1    g17724(.A1(new_n20160_), .A2(new_n12770_), .ZN(new_n20161_));
  NOR3_X1    g17725(.A1(new_n20159_), .A2(pi1155), .A3(new_n20155_), .ZN(new_n20162_));
  NOR3_X1    g17726(.A1(new_n20161_), .A2(new_n12764_), .A3(new_n20162_), .ZN(new_n20163_));
  NOR2_X1    g17727(.A1(new_n20163_), .A2(new_n20157_), .ZN(new_n20164_));
  INV_X1     g17728(.I(new_n20164_), .ZN(new_n20165_));
  AOI21_X1   g17729(.A1(new_n20165_), .A2(new_n12783_), .B(pi1154), .ZN(new_n20166_));
  AOI21_X1   g17730(.A1(new_n20165_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n20167_));
  NOR3_X1    g17731(.A1(new_n20166_), .A2(new_n20167_), .A3(new_n12779_), .ZN(new_n20168_));
  AOI21_X1   g17732(.A1(new_n12779_), .A2(new_n20165_), .B(new_n20168_), .ZN(new_n20169_));
  OAI21_X1   g17733(.A1(new_n20169_), .A2(new_n17229_), .B(new_n12791_), .ZN(new_n20170_));
  OAI21_X1   g17734(.A1(new_n20169_), .A2(new_n17232_), .B(pi1159), .ZN(new_n20171_));
  NAND3_X1   g17735(.A1(new_n20170_), .A2(new_n20171_), .A3(pi0789), .ZN(new_n20172_));
  OAI21_X1   g17736(.A1(pi0789), .A2(new_n20169_), .B(new_n20172_), .ZN(new_n20173_));
  INV_X1     g17737(.I(new_n20155_), .ZN(new_n20174_));
  NAND2_X1   g17738(.A1(new_n12818_), .A2(new_n20174_), .ZN(new_n20175_));
  OAI21_X1   g17739(.A1(new_n20173_), .A2(new_n12818_), .B(new_n20175_), .ZN(new_n20176_));
  AOI21_X1   g17740(.A1(new_n12826_), .A2(new_n16620_), .B(new_n20155_), .ZN(new_n20177_));
  NOR2_X1    g17741(.A1(new_n20155_), .A2(pi1153), .ZN(new_n20178_));
  NOR2_X1    g17742(.A1(new_n12834_), .A2(pi0734), .ZN(new_n20179_));
  INV_X1     g17743(.I(new_n20179_), .ZN(new_n20180_));
  NAND2_X1   g17744(.A1(new_n20180_), .A2(new_n20178_), .ZN(new_n20181_));
  NOR2_X1    g17745(.A1(new_n20179_), .A2(new_n20177_), .ZN(new_n20182_));
  NOR2_X1    g17746(.A1(new_n20182_), .A2(new_n12841_), .ZN(new_n20183_));
  INV_X1     g17747(.I(new_n20183_), .ZN(new_n20184_));
  NAND3_X1   g17748(.A1(new_n20184_), .A2(pi0778), .A3(new_n20181_), .ZN(new_n20185_));
  OAI21_X1   g17749(.A1(pi0778), .A2(new_n20177_), .B(new_n20185_), .ZN(new_n20186_));
  NAND2_X1   g17750(.A1(new_n20186_), .A2(new_n17187_), .ZN(new_n20187_));
  NOR2_X1    g17751(.A1(new_n20187_), .A2(new_n12889_), .ZN(new_n20188_));
  NAND2_X1   g17752(.A1(new_n20188_), .A2(new_n18203_), .ZN(new_n20189_));
  NOR2_X1    g17753(.A1(new_n20189_), .A2(new_n17884_), .ZN(new_n20190_));
  INV_X1     g17754(.I(new_n20190_), .ZN(new_n20191_));
  OAI22_X1   g17755(.A1(new_n20176_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n20191_), .ZN(new_n20192_));
  AND2_X2    g17756(.A1(new_n20192_), .A2(new_n12919_), .Z(new_n20193_));
  OAI22_X1   g17757(.A1(new_n20176_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n20191_), .ZN(new_n20194_));
  AOI21_X1   g17758(.A1(pi0629), .A2(new_n20194_), .B(new_n20193_), .ZN(new_n20195_));
  INV_X1     g17759(.I(new_n20162_), .ZN(new_n20196_));
  NOR2_X1    g17760(.A1(new_n20177_), .A2(new_n12754_), .ZN(new_n20197_));
  NOR3_X1    g17761(.A1(new_n20197_), .A2(new_n20154_), .A3(new_n20155_), .ZN(new_n20198_));
  NAND2_X1   g17762(.A1(new_n20198_), .A2(new_n12758_), .ZN(new_n20199_));
  NAND2_X1   g17763(.A1(new_n20197_), .A2(pi0625), .ZN(new_n20200_));
  NAND3_X1   g17764(.A1(new_n20200_), .A2(pi1153), .A3(new_n20156_), .ZN(new_n20201_));
  NAND3_X1   g17765(.A1(new_n20181_), .A2(pi0608), .A3(new_n20201_), .ZN(new_n20202_));
  INV_X1     g17766(.I(new_n20200_), .ZN(new_n20203_));
  OAI21_X1   g17767(.A1(new_n20203_), .A2(new_n20198_), .B(new_n20178_), .ZN(new_n20204_));
  NAND3_X1   g17768(.A1(new_n20184_), .A2(new_n13560_), .A3(new_n20204_), .ZN(new_n20205_));
  NAND3_X1   g17769(.A1(new_n20205_), .A2(pi0778), .A3(new_n20202_), .ZN(new_n20206_));
  AOI21_X1   g17770(.A1(new_n20206_), .A2(new_n20199_), .B(new_n12766_), .ZN(new_n20207_));
  NOR2_X1    g17771(.A1(new_n20186_), .A2(pi0609), .ZN(new_n20208_));
  OAI21_X1   g17772(.A1(new_n20208_), .A2(new_n20207_), .B(pi1155), .ZN(new_n20209_));
  NAND3_X1   g17773(.A1(new_n20209_), .A2(pi0660), .A3(new_n20196_), .ZN(new_n20210_));
  NAND2_X1   g17774(.A1(new_n20206_), .A2(new_n20199_), .ZN(new_n20211_));
  NOR2_X1    g17775(.A1(new_n20186_), .A2(new_n12766_), .ZN(new_n20212_));
  AOI21_X1   g17776(.A1(new_n20211_), .A2(new_n12766_), .B(new_n20212_), .ZN(new_n20213_));
  NOR2_X1    g17777(.A1(new_n20161_), .A2(pi0660), .ZN(new_n20214_));
  OAI21_X1   g17778(.A1(new_n20213_), .A2(pi1155), .B(new_n20214_), .ZN(new_n20215_));
  NAND3_X1   g17779(.A1(new_n20215_), .A2(new_n20210_), .A3(pi0785), .ZN(new_n20216_));
  NAND2_X1   g17780(.A1(new_n20211_), .A2(new_n12764_), .ZN(new_n20217_));
  NAND2_X1   g17781(.A1(new_n20216_), .A2(new_n20217_), .ZN(new_n20218_));
  NAND2_X1   g17782(.A1(new_n20218_), .A2(new_n12781_), .ZN(new_n20219_));
  NAND2_X1   g17783(.A1(new_n20187_), .A2(pi0618), .ZN(new_n20220_));
  AOI21_X1   g17784(.A1(new_n20219_), .A2(new_n20220_), .B(pi1154), .ZN(new_n20221_));
  NOR3_X1    g17785(.A1(new_n20221_), .A2(pi0627), .A3(new_n20167_), .ZN(new_n20222_));
  NAND2_X1   g17786(.A1(new_n20187_), .A2(new_n12781_), .ZN(new_n20223_));
  NAND2_X1   g17787(.A1(new_n20218_), .A2(pi0618), .ZN(new_n20224_));
  AOI21_X1   g17788(.A1(new_n20224_), .A2(new_n20223_), .B(new_n12785_), .ZN(new_n20225_));
  NOR3_X1    g17789(.A1(new_n20225_), .A2(new_n12880_), .A3(new_n20166_), .ZN(new_n20226_));
  OR3_X2     g17790(.A1(new_n20222_), .A2(new_n20226_), .A3(new_n12779_), .Z(new_n20227_));
  NAND2_X1   g17791(.A1(new_n20218_), .A2(new_n12779_), .ZN(new_n20228_));
  NAND2_X1   g17792(.A1(new_n20227_), .A2(new_n20228_), .ZN(new_n20229_));
  AOI21_X1   g17793(.A1(new_n20229_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n20230_));
  NOR2_X1    g17794(.A1(new_n20188_), .A2(pi0619), .ZN(new_n20231_));
  AOI21_X1   g17795(.A1(new_n20227_), .A2(new_n20228_), .B(new_n12793_), .ZN(new_n20232_));
  OAI21_X1   g17796(.A1(new_n20232_), .A2(new_n20231_), .B(pi1159), .ZN(new_n20233_));
  NAND3_X1   g17797(.A1(new_n20233_), .A2(pi0648), .A3(new_n20170_), .ZN(new_n20234_));
  NAND2_X1   g17798(.A1(new_n20229_), .A2(new_n12793_), .ZN(new_n20235_));
  OAI21_X1   g17799(.A1(new_n12793_), .A2(new_n20188_), .B(new_n20235_), .ZN(new_n20236_));
  NAND2_X1   g17800(.A1(new_n20236_), .A2(new_n12791_), .ZN(new_n20237_));
  NAND3_X1   g17801(.A1(new_n20237_), .A2(new_n12895_), .A3(new_n20171_), .ZN(new_n20238_));
  NAND3_X1   g17802(.A1(new_n20238_), .A2(pi0789), .A3(new_n20234_), .ZN(new_n20239_));
  NOR2_X1    g17803(.A1(new_n20174_), .A2(new_n12747_), .ZN(new_n20240_));
  AND2_X2    g17804(.A1(new_n20173_), .A2(new_n12747_), .Z(new_n20241_));
  OAI21_X1   g17805(.A1(new_n20241_), .A2(new_n20240_), .B(new_n12815_), .ZN(new_n20242_));
  INV_X1     g17806(.I(new_n20189_), .ZN(new_n20243_));
  NAND2_X1   g17807(.A1(new_n20173_), .A2(pi0626), .ZN(new_n20244_));
  OAI21_X1   g17808(.A1(pi0626), .A2(new_n20174_), .B(new_n20244_), .ZN(new_n20245_));
  AOI22_X1   g17809(.A1(new_n20245_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n20243_), .ZN(new_n20246_));
  NAND2_X1   g17810(.A1(new_n20246_), .A2(new_n20242_), .ZN(new_n20247_));
  AOI22_X1   g17811(.A1(new_n20239_), .A2(new_n20230_), .B1(pi0788), .B2(new_n20247_), .ZN(new_n20248_));
  OAI22_X1   g17812(.A1(new_n20248_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n20195_), .ZN(new_n20249_));
  NAND2_X1   g17813(.A1(new_n20176_), .A2(new_n13384_), .ZN(new_n20250_));
  NAND2_X1   g17814(.A1(new_n12943_), .A2(new_n20174_), .ZN(new_n20251_));
  NAND2_X1   g17815(.A1(new_n20250_), .A2(new_n20251_), .ZN(new_n20252_));
  NOR2_X1    g17816(.A1(new_n20191_), .A2(new_n12953_), .ZN(new_n20253_));
  NOR2_X1    g17817(.A1(new_n20253_), .A2(pi0647), .ZN(new_n20254_));
  NOR2_X1    g17818(.A1(new_n20155_), .A2(new_n12741_), .ZN(new_n20255_));
  OAI21_X1   g17819(.A1(new_n20254_), .A2(new_n20255_), .B(new_n12965_), .ZN(new_n20256_));
  NAND2_X1   g17820(.A1(new_n20253_), .A2(pi0647), .ZN(new_n20257_));
  OAI21_X1   g17821(.A1(pi0647), .A2(new_n20174_), .B(new_n20257_), .ZN(new_n20258_));
  OAI22_X1   g17822(.A1(new_n20258_), .A2(new_n15576_), .B1(new_n20256_), .B2(new_n12981_), .ZN(new_n20259_));
  AOI21_X1   g17823(.A1(new_n20252_), .A2(new_n15608_), .B(new_n20259_), .ZN(new_n20260_));
  OAI22_X1   g17824(.A1(new_n20249_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n20260_), .ZN(new_n20261_));
  NAND2_X1   g17825(.A1(new_n20261_), .A2(new_n13000_), .ZN(new_n20262_));
  AND2_X2    g17826(.A1(new_n20261_), .A2(new_n12975_), .Z(new_n20263_));
  OAI21_X1   g17827(.A1(new_n20258_), .A2(new_n12965_), .B(new_n20256_), .ZN(new_n20264_));
  NAND2_X1   g17828(.A1(new_n20253_), .A2(new_n12972_), .ZN(new_n20265_));
  OAI21_X1   g17829(.A1(new_n20264_), .A2(new_n12972_), .B(new_n20265_), .ZN(new_n20266_));
  NOR2_X1    g17830(.A1(new_n20266_), .A2(new_n12975_), .ZN(new_n20267_));
  OAI21_X1   g17831(.A1(new_n20263_), .A2(new_n20267_), .B(new_n12740_), .ZN(new_n20268_));
  NAND2_X1   g17832(.A1(new_n20174_), .A2(pi0644), .ZN(new_n20269_));
  NOR2_X1    g17833(.A1(new_n17611_), .A2(new_n20155_), .ZN(new_n20270_));
  AOI21_X1   g17834(.A1(new_n20176_), .A2(new_n17611_), .B(new_n20270_), .ZN(new_n20271_));
  OAI21_X1   g17835(.A1(new_n20271_), .A2(pi0644), .B(new_n20269_), .ZN(new_n20272_));
  NAND2_X1   g17836(.A1(new_n20272_), .A2(pi0715), .ZN(new_n20273_));
  NAND3_X1   g17837(.A1(new_n20268_), .A2(new_n12739_), .A3(new_n20273_), .ZN(new_n20274_));
  NOR2_X1    g17838(.A1(new_n20266_), .A2(pi0644), .ZN(new_n20275_));
  AOI21_X1   g17839(.A1(new_n20261_), .A2(pi0644), .B(new_n20275_), .ZN(new_n20276_));
  NAND2_X1   g17840(.A1(new_n20174_), .A2(new_n12975_), .ZN(new_n20277_));
  OAI21_X1   g17841(.A1(new_n20271_), .A2(new_n12975_), .B(new_n20277_), .ZN(new_n20278_));
  AOI21_X1   g17842(.A1(new_n20278_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n20279_));
  OAI21_X1   g17843(.A1(new_n20276_), .A2(new_n12740_), .B(new_n20279_), .ZN(new_n20280_));
  NAND3_X1   g17844(.A1(new_n20274_), .A2(pi0790), .A3(new_n20280_), .ZN(new_n20281_));
  NAND2_X1   g17845(.A1(new_n20281_), .A2(new_n20262_), .ZN(new_n20282_));
  AOI21_X1   g17846(.A1(po1038), .A2(new_n5659_), .B(pi0832), .ZN(new_n20283_));
  NAND2_X1   g17847(.A1(new_n13192_), .A2(new_n5659_), .ZN(new_n20284_));
  INV_X1     g17848(.I(new_n20284_), .ZN(new_n20285_));
  AOI21_X1   g17849(.A1(new_n20285_), .A2(pi0644), .B(new_n12740_), .ZN(new_n20286_));
  NAND2_X1   g17850(.A1(new_n20284_), .A2(new_n12984_), .ZN(new_n20287_));
  NOR2_X1    g17851(.A1(new_n20285_), .A2(new_n13384_), .ZN(new_n20288_));
  NOR2_X1    g17852(.A1(new_n2609_), .A2(new_n5659_), .ZN(new_n20289_));
  NOR2_X1    g17853(.A1(new_n13342_), .A2(pi0756), .ZN(new_n20290_));
  NOR2_X1    g17854(.A1(new_n13344_), .A2(pi0182), .ZN(new_n20291_));
  NOR3_X1    g17855(.A1(new_n20290_), .A2(new_n3265_), .A3(new_n20291_), .ZN(new_n20292_));
  NAND2_X1   g17856(.A1(new_n13334_), .A2(new_n5659_), .ZN(new_n20293_));
  NAND2_X1   g17857(.A1(new_n13245_), .A2(pi0182), .ZN(new_n20294_));
  AOI21_X1   g17858(.A1(new_n20293_), .A2(new_n20294_), .B(pi0756), .ZN(new_n20295_));
  NOR3_X1    g17859(.A1(new_n15787_), .A2(pi0182), .A3(new_n16621_), .ZN(new_n20296_));
  NOR2_X1    g17860(.A1(new_n20295_), .A2(new_n20296_), .ZN(new_n20297_));
  AOI21_X1   g17861(.A1(new_n20297_), .A2(new_n3265_), .B(new_n20292_), .ZN(new_n20298_));
  NOR2_X1    g17862(.A1(new_n20298_), .A2(new_n2610_), .ZN(new_n20299_));
  NOR2_X1    g17863(.A1(new_n20299_), .A2(new_n20289_), .ZN(new_n20300_));
  NOR2_X1    g17864(.A1(new_n20300_), .A2(new_n12760_), .ZN(new_n20301_));
  INV_X1     g17865(.I(new_n20301_), .ZN(new_n20302_));
  OAI21_X1   g17866(.A1(new_n12761_), .A2(new_n20285_), .B(new_n20302_), .ZN(new_n20303_));
  OAI22_X1   g17867(.A1(new_n20302_), .A2(pi0609), .B1(new_n13353_), .B2(new_n20285_), .ZN(new_n20304_));
  NAND2_X1   g17868(.A1(new_n20304_), .A2(new_n12770_), .ZN(new_n20305_));
  INV_X1     g17869(.I(new_n20305_), .ZN(new_n20306_));
  AOI22_X1   g17870(.A1(new_n20301_), .A2(pi0609), .B1(new_n13357_), .B2(new_n20284_), .ZN(new_n20307_));
  OAI21_X1   g17871(.A1(new_n20307_), .A2(new_n12770_), .B(pi0785), .ZN(new_n20308_));
  OAI22_X1   g17872(.A1(new_n20306_), .A2(new_n20308_), .B1(pi0785), .B2(new_n20303_), .ZN(new_n20309_));
  NAND2_X1   g17873(.A1(new_n20309_), .A2(new_n12779_), .ZN(new_n20310_));
  NAND2_X1   g17874(.A1(new_n20284_), .A2(pi0618), .ZN(new_n20311_));
  OAI21_X1   g17875(.A1(new_n20309_), .A2(pi0618), .B(new_n20311_), .ZN(new_n20312_));
  NAND2_X1   g17876(.A1(new_n20312_), .A2(new_n12785_), .ZN(new_n20313_));
  NAND2_X1   g17877(.A1(new_n20284_), .A2(new_n12781_), .ZN(new_n20314_));
  OAI21_X1   g17878(.A1(new_n20309_), .A2(new_n12781_), .B(new_n20314_), .ZN(new_n20315_));
  NAND2_X1   g17879(.A1(new_n20315_), .A2(pi1154), .ZN(new_n20316_));
  NAND3_X1   g17880(.A1(new_n20313_), .A2(new_n20316_), .A3(pi0781), .ZN(new_n20317_));
  NAND2_X1   g17881(.A1(new_n20317_), .A2(new_n20310_), .ZN(new_n20318_));
  NAND2_X1   g17882(.A1(new_n20318_), .A2(new_n12796_), .ZN(new_n20319_));
  NAND2_X1   g17883(.A1(new_n20284_), .A2(pi0619), .ZN(new_n20320_));
  OAI21_X1   g17884(.A1(new_n20318_), .A2(pi0619), .B(new_n20320_), .ZN(new_n20321_));
  NAND2_X1   g17885(.A1(new_n20321_), .A2(new_n12791_), .ZN(new_n20322_));
  NAND2_X1   g17886(.A1(new_n20284_), .A2(new_n12793_), .ZN(new_n20323_));
  OAI21_X1   g17887(.A1(new_n20318_), .A2(new_n12793_), .B(new_n20323_), .ZN(new_n20324_));
  NAND2_X1   g17888(.A1(new_n20324_), .A2(pi1159), .ZN(new_n20325_));
  NAND3_X1   g17889(.A1(new_n20322_), .A2(new_n20325_), .A3(pi0789), .ZN(new_n20326_));
  NAND2_X1   g17890(.A1(new_n20326_), .A2(new_n20319_), .ZN(new_n20327_));
  NAND2_X1   g17891(.A1(new_n20284_), .A2(new_n12818_), .ZN(new_n20328_));
  OAI21_X1   g17892(.A1(new_n20327_), .A2(new_n12818_), .B(new_n20328_), .ZN(new_n20329_));
  AOI21_X1   g17893(.A1(new_n20329_), .A2(new_n13384_), .B(new_n20288_), .ZN(new_n20330_));
  OAI21_X1   g17894(.A1(new_n20330_), .A2(new_n12984_), .B(new_n20287_), .ZN(new_n20331_));
  OAI21_X1   g17895(.A1(new_n20331_), .A2(pi0644), .B(new_n20286_), .ZN(new_n20332_));
  AND2_X2    g17896(.A1(new_n20332_), .A2(new_n12739_), .Z(new_n20333_));
  OAI21_X1   g17897(.A1(new_n14125_), .A2(new_n20291_), .B(new_n16620_), .ZN(new_n20334_));
  OAI21_X1   g17898(.A1(new_n14122_), .A2(new_n5659_), .B(new_n3265_), .ZN(new_n20335_));
  NAND2_X1   g17899(.A1(new_n20335_), .A2(new_n2609_), .ZN(new_n20336_));
  NAND2_X1   g17900(.A1(new_n15744_), .A2(new_n5659_), .ZN(new_n20337_));
  AOI21_X1   g17901(.A1(new_n20337_), .A2(new_n20336_), .B(new_n20334_), .ZN(new_n20338_));
  NAND2_X1   g17902(.A1(new_n2609_), .A2(new_n16620_), .ZN(new_n20339_));
  AOI21_X1   g17903(.A1(new_n20285_), .A2(new_n20339_), .B(new_n20338_), .ZN(new_n20340_));
  NAND2_X1   g17904(.A1(new_n20340_), .A2(new_n13521_), .ZN(new_n20341_));
  NAND2_X1   g17905(.A1(new_n20284_), .A2(pi0625), .ZN(new_n20342_));
  AOI21_X1   g17906(.A1(new_n20341_), .A2(new_n20342_), .B(pi1153), .ZN(new_n20343_));
  NAND2_X1   g17907(.A1(new_n20284_), .A2(new_n13521_), .ZN(new_n20344_));
  NAND2_X1   g17908(.A1(new_n20340_), .A2(pi0625), .ZN(new_n20345_));
  AOI21_X1   g17909(.A1(new_n20345_), .A2(new_n20344_), .B(new_n12841_), .ZN(new_n20346_));
  NOR3_X1    g17910(.A1(new_n20343_), .A2(new_n20346_), .A3(new_n12758_), .ZN(new_n20347_));
  NOR2_X1    g17911(.A1(new_n20340_), .A2(pi0778), .ZN(new_n20348_));
  NOR2_X1    g17912(.A1(new_n20347_), .A2(new_n20348_), .ZN(new_n20349_));
  NOR2_X1    g17913(.A1(new_n20349_), .A2(new_n12869_), .ZN(new_n20350_));
  AOI21_X1   g17914(.A1(new_n12869_), .A2(new_n20285_), .B(new_n20350_), .ZN(new_n20351_));
  NAND2_X1   g17915(.A1(new_n20351_), .A2(new_n12888_), .ZN(new_n20352_));
  OAI21_X1   g17916(.A1(new_n12888_), .A2(new_n20285_), .B(new_n20352_), .ZN(new_n20353_));
  INV_X1     g17917(.I(new_n20353_), .ZN(new_n20354_));
  NOR2_X1    g17918(.A1(new_n20284_), .A2(new_n12911_), .ZN(new_n20355_));
  AOI21_X1   g17919(.A1(new_n20354_), .A2(new_n12911_), .B(new_n20355_), .ZN(new_n20356_));
  NAND2_X1   g17920(.A1(new_n20356_), .A2(new_n13392_), .ZN(new_n20357_));
  OAI21_X1   g17921(.A1(new_n13392_), .A2(new_n20285_), .B(new_n20357_), .ZN(new_n20358_));
  NAND2_X1   g17922(.A1(new_n20358_), .A2(new_n12920_), .ZN(new_n20359_));
  NAND2_X1   g17923(.A1(new_n20284_), .A2(pi0628), .ZN(new_n20360_));
  AOI21_X1   g17924(.A1(new_n20359_), .A2(new_n20360_), .B(pi1156), .ZN(new_n20361_));
  NAND2_X1   g17925(.A1(new_n20284_), .A2(new_n12920_), .ZN(new_n20362_));
  NAND2_X1   g17926(.A1(new_n20358_), .A2(pi0628), .ZN(new_n20363_));
  AOI21_X1   g17927(.A1(new_n20363_), .A2(new_n20362_), .B(new_n12742_), .ZN(new_n20364_));
  OR2_X2     g17928(.A1(new_n20364_), .A2(new_n12937_), .Z(new_n20365_));
  OAI22_X1   g17929(.A1(new_n20365_), .A2(new_n20361_), .B1(pi0792), .B2(new_n20358_), .ZN(new_n20366_));
  NAND2_X1   g17930(.A1(new_n20366_), .A2(new_n12741_), .ZN(new_n20367_));
  OAI21_X1   g17931(.A1(new_n12741_), .A2(new_n20284_), .B(new_n20367_), .ZN(new_n20368_));
  NOR2_X1    g17932(.A1(new_n20368_), .A2(pi1157), .ZN(new_n20369_));
  NAND2_X1   g17933(.A1(new_n20366_), .A2(pi0647), .ZN(new_n20370_));
  OAI21_X1   g17934(.A1(pi0647), .A2(new_n20284_), .B(new_n20370_), .ZN(new_n20371_));
  NOR2_X1    g17935(.A1(new_n20371_), .A2(new_n12965_), .ZN(new_n20372_));
  OAI21_X1   g17936(.A1(new_n20369_), .A2(new_n20372_), .B(pi0787), .ZN(new_n20373_));
  OAI21_X1   g17937(.A1(pi0787), .A2(new_n20366_), .B(new_n20373_), .ZN(new_n20374_));
  OAI21_X1   g17938(.A1(new_n20374_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n20375_));
  AOI21_X1   g17939(.A1(new_n20285_), .A2(new_n12975_), .B(pi0715), .ZN(new_n20376_));
  OAI21_X1   g17940(.A1(new_n20331_), .A2(new_n12975_), .B(new_n20376_), .ZN(new_n20377_));
  AND2_X2    g17941(.A1(new_n20377_), .A2(pi1160), .Z(new_n20378_));
  OAI21_X1   g17942(.A1(new_n20374_), .A2(pi0644), .B(pi0715), .ZN(new_n20379_));
  AOI22_X1   g17943(.A1(new_n20333_), .A2(new_n20375_), .B1(new_n20379_), .B2(new_n20378_), .ZN(new_n20380_));
  NOR2_X1    g17944(.A1(new_n20380_), .A2(new_n13000_), .ZN(new_n20381_));
  NAND2_X1   g17945(.A1(new_n20285_), .A2(pi0626), .ZN(new_n20382_));
  NAND2_X1   g17946(.A1(new_n20327_), .A2(new_n12747_), .ZN(new_n20383_));
  AOI21_X1   g17947(.A1(new_n20383_), .A2(new_n20382_), .B(new_n12816_), .ZN(new_n20384_));
  NOR2_X1    g17948(.A1(new_n20284_), .A2(pi0626), .ZN(new_n20385_));
  AOI21_X1   g17949(.A1(new_n20327_), .A2(pi0626), .B(new_n20385_), .ZN(new_n20386_));
  OAI22_X1   g17950(.A1(new_n20386_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n20356_), .ZN(new_n20387_));
  OAI21_X1   g17951(.A1(new_n20387_), .A2(new_n20384_), .B(pi0788), .ZN(new_n20388_));
  NAND2_X1   g17952(.A1(new_n20388_), .A2(new_n15824_), .ZN(new_n20389_));
  NAND2_X1   g17953(.A1(new_n20349_), .A2(new_n12766_), .ZN(new_n20390_));
  AOI21_X1   g17954(.A1(new_n16621_), .A2(new_n13566_), .B(new_n15826_), .ZN(new_n20391_));
  AOI21_X1   g17955(.A1(new_n14328_), .A2(new_n20158_), .B(new_n5659_), .ZN(new_n20392_));
  AOI21_X1   g17956(.A1(new_n20392_), .A2(new_n5336_), .B(new_n3265_), .ZN(new_n20393_));
  OAI21_X1   g17957(.A1(new_n20391_), .A2(pi0182), .B(new_n20393_), .ZN(new_n20394_));
  NAND2_X1   g17958(.A1(new_n14172_), .A2(pi0182), .ZN(new_n20395_));
  NAND2_X1   g17959(.A1(new_n14174_), .A2(new_n5659_), .ZN(new_n20396_));
  AOI21_X1   g17960(.A1(new_n20395_), .A2(new_n20396_), .B(pi0756), .ZN(new_n20397_));
  NAND2_X1   g17961(.A1(new_n15835_), .A2(pi0182), .ZN(new_n20398_));
  NAND2_X1   g17962(.A1(new_n14177_), .A2(new_n5659_), .ZN(new_n20399_));
  AOI21_X1   g17963(.A1(new_n20399_), .A2(new_n20398_), .B(new_n16621_), .ZN(new_n20400_));
  OAI21_X1   g17964(.A1(new_n20400_), .A2(new_n20397_), .B(new_n2627_), .ZN(new_n20401_));
  NOR2_X1    g17965(.A1(new_n14182_), .A2(pi0182), .ZN(new_n20402_));
  NOR2_X1    g17966(.A1(new_n14184_), .A2(new_n5659_), .ZN(new_n20403_));
  OAI21_X1   g17967(.A1(new_n20402_), .A2(new_n20403_), .B(pi0756), .ZN(new_n20404_));
  NOR2_X1    g17968(.A1(new_n14187_), .A2(new_n5659_), .ZN(new_n20405_));
  NOR2_X1    g17969(.A1(new_n14189_), .A2(pi0182), .ZN(new_n20406_));
  OAI21_X1   g17970(.A1(new_n20405_), .A2(new_n20406_), .B(new_n16621_), .ZN(new_n20407_));
  NAND3_X1   g17971(.A1(new_n20407_), .A2(new_n20404_), .A3(pi0039), .ZN(new_n20408_));
  NAND3_X1   g17972(.A1(new_n20408_), .A2(new_n3265_), .A3(new_n20401_), .ZN(new_n20409_));
  NAND3_X1   g17973(.A1(new_n20409_), .A2(new_n16620_), .A3(new_n20394_), .ZN(new_n20410_));
  NAND2_X1   g17974(.A1(new_n20298_), .A2(pi0734), .ZN(new_n20411_));
  NAND3_X1   g17975(.A1(new_n20410_), .A2(new_n2609_), .A3(new_n20411_), .ZN(new_n20412_));
  OAI21_X1   g17976(.A1(new_n5659_), .A2(new_n2609_), .B(new_n20412_), .ZN(new_n20413_));
  INV_X1     g17977(.I(new_n20346_), .ZN(new_n20414_));
  NOR2_X1    g17978(.A1(new_n20300_), .A2(new_n13521_), .ZN(new_n20415_));
  AOI21_X1   g17979(.A1(new_n20413_), .A2(new_n13521_), .B(new_n20415_), .ZN(new_n20416_));
  OAI21_X1   g17980(.A1(new_n20416_), .A2(pi1153), .B(new_n20414_), .ZN(new_n20417_));
  NOR2_X1    g17981(.A1(new_n20300_), .A2(pi0625), .ZN(new_n20418_));
  AOI21_X1   g17982(.A1(new_n20413_), .A2(pi0625), .B(new_n20418_), .ZN(new_n20419_));
  OAI21_X1   g17983(.A1(new_n20419_), .A2(new_n12841_), .B(pi0608), .ZN(new_n20420_));
  OAI22_X1   g17984(.A1(pi0608), .A2(new_n20417_), .B1(new_n20420_), .B2(new_n20343_), .ZN(new_n20421_));
  NOR2_X1    g17985(.A1(new_n20421_), .A2(new_n12758_), .ZN(new_n20422_));
  AOI21_X1   g17986(.A1(new_n12758_), .A2(new_n20413_), .B(new_n20422_), .ZN(new_n20423_));
  OAI21_X1   g17987(.A1(new_n20423_), .A2(new_n12766_), .B(new_n20390_), .ZN(new_n20424_));
  AOI21_X1   g17988(.A1(new_n20424_), .A2(pi1155), .B(new_n20306_), .ZN(new_n20425_));
  NOR2_X1    g17989(.A1(new_n20423_), .A2(pi0609), .ZN(new_n20426_));
  NOR3_X1    g17990(.A1(new_n20347_), .A2(new_n12766_), .A3(new_n20348_), .ZN(new_n20427_));
  OAI21_X1   g17991(.A1(new_n20426_), .A2(new_n20427_), .B(new_n12770_), .ZN(new_n20428_));
  NOR2_X1    g17992(.A1(new_n20307_), .A2(new_n12770_), .ZN(new_n20429_));
  NOR2_X1    g17993(.A1(new_n20429_), .A2(pi0660), .ZN(new_n20430_));
  AOI22_X1   g17994(.A1(new_n20425_), .A2(pi0660), .B1(new_n20428_), .B2(new_n20430_), .ZN(new_n20431_));
  NOR2_X1    g17995(.A1(new_n20423_), .A2(pi0785), .ZN(new_n20432_));
  AOI21_X1   g17996(.A1(new_n20431_), .A2(pi0785), .B(new_n20432_), .ZN(new_n20433_));
  NOR2_X1    g17997(.A1(new_n20433_), .A2(pi0781), .ZN(new_n20434_));
  AND2_X2    g17998(.A1(new_n20351_), .A2(new_n12781_), .Z(new_n20435_));
  NOR2_X1    g17999(.A1(new_n20433_), .A2(new_n12781_), .ZN(new_n20436_));
  OAI21_X1   g18000(.A1(new_n20436_), .A2(new_n20435_), .B(pi1154), .ZN(new_n20437_));
  NAND3_X1   g18001(.A1(new_n20437_), .A2(pi0627), .A3(new_n20313_), .ZN(new_n20438_));
  INV_X1     g18002(.I(new_n20316_), .ZN(new_n20439_));
  NAND2_X1   g18003(.A1(new_n20351_), .A2(pi0618), .ZN(new_n20440_));
  OAI21_X1   g18004(.A1(new_n20433_), .A2(pi0618), .B(new_n20440_), .ZN(new_n20441_));
  AOI21_X1   g18005(.A1(new_n20441_), .A2(new_n12785_), .B(new_n20439_), .ZN(new_n20442_));
  AOI21_X1   g18006(.A1(new_n20442_), .A2(new_n12880_), .B(new_n12779_), .ZN(new_n20443_));
  AOI21_X1   g18007(.A1(new_n20443_), .A2(new_n20438_), .B(new_n20434_), .ZN(new_n20444_));
  OAI21_X1   g18008(.A1(new_n20444_), .A2(pi0789), .B(new_n12819_), .ZN(new_n20445_));
  NOR2_X1    g18009(.A1(new_n20354_), .A2(new_n12793_), .ZN(new_n20446_));
  NOR2_X1    g18010(.A1(new_n20444_), .A2(pi0619), .ZN(new_n20447_));
  OAI21_X1   g18011(.A1(new_n20447_), .A2(new_n20446_), .B(new_n12791_), .ZN(new_n20448_));
  NAND3_X1   g18012(.A1(new_n20448_), .A2(new_n12895_), .A3(new_n20325_), .ZN(new_n20449_));
  NAND2_X1   g18013(.A1(new_n20353_), .A2(new_n12793_), .ZN(new_n20450_));
  OAI21_X1   g18014(.A1(new_n20444_), .A2(new_n12793_), .B(new_n20450_), .ZN(new_n20451_));
  AOI21_X1   g18015(.A1(new_n20451_), .A2(pi1159), .B(new_n12895_), .ZN(new_n20452_));
  AOI21_X1   g18016(.A1(new_n20452_), .A2(new_n20322_), .B(new_n12796_), .ZN(new_n20453_));
  AOI21_X1   g18017(.A1(new_n20453_), .A2(new_n20449_), .B(new_n20445_), .ZN(new_n20454_));
  NOR2_X1    g18018(.A1(new_n20364_), .A2(pi0629), .ZN(new_n20455_));
  NOR2_X1    g18019(.A1(new_n20361_), .A2(new_n12919_), .ZN(new_n20456_));
  NOR2_X1    g18020(.A1(new_n20455_), .A2(new_n20456_), .ZN(new_n20457_));
  AOI21_X1   g18021(.A1(new_n20329_), .A2(new_n19160_), .B(new_n20457_), .ZN(new_n20458_));
  OAI22_X1   g18022(.A1(new_n20454_), .A2(new_n20389_), .B1(new_n12937_), .B2(new_n20458_), .ZN(new_n20459_));
  NOR2_X1    g18023(.A1(new_n20378_), .A2(new_n12975_), .ZN(new_n20460_));
  NOR2_X1    g18024(.A1(new_n20333_), .A2(pi0644), .ZN(new_n20461_));
  NOR2_X1    g18025(.A1(new_n20460_), .A2(new_n20461_), .ZN(new_n20462_));
  OAI22_X1   g18026(.A1(new_n15576_), .A2(new_n20371_), .B1(new_n20368_), .B2(new_n15730_), .ZN(new_n20463_));
  NOR2_X1    g18027(.A1(new_n20330_), .A2(new_n17212_), .ZN(new_n20464_));
  NOR2_X1    g18028(.A1(new_n20463_), .A2(new_n20464_), .ZN(new_n20465_));
  OAI22_X1   g18029(.A1(new_n20462_), .A2(new_n13000_), .B1(new_n20465_), .B2(new_n12972_), .ZN(new_n20466_));
  AOI21_X1   g18030(.A1(new_n15693_), .A2(new_n20459_), .B(new_n20466_), .ZN(new_n20467_));
  OAI21_X1   g18031(.A1(new_n20381_), .A2(new_n20467_), .B(new_n6643_), .ZN(new_n20468_));
  AOI22_X1   g18032(.A1(new_n20468_), .A2(new_n20283_), .B1(pi0832), .B2(new_n20282_), .ZN(po0339));
  NOR2_X1    g18033(.A1(new_n13340_), .A2(pi0755), .ZN(new_n20470_));
  NOR2_X1    g18034(.A1(new_n3042_), .A2(pi0183), .ZN(new_n20471_));
  NOR2_X1    g18035(.A1(new_n20470_), .A2(new_n20471_), .ZN(new_n20472_));
  NOR3_X1    g18036(.A1(new_n20472_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n20473_));
  INV_X1     g18037(.I(new_n20470_), .ZN(new_n20474_));
  NOR2_X1    g18038(.A1(new_n20474_), .A2(new_n13354_), .ZN(new_n20475_));
  NOR3_X1    g18039(.A1(new_n20475_), .A2(new_n12762_), .A3(new_n20472_), .ZN(new_n20476_));
  NOR2_X1    g18040(.A1(new_n20476_), .A2(new_n12770_), .ZN(new_n20477_));
  NOR3_X1    g18041(.A1(new_n20475_), .A2(pi1155), .A3(new_n20471_), .ZN(new_n20478_));
  NOR3_X1    g18042(.A1(new_n20477_), .A2(new_n12764_), .A3(new_n20478_), .ZN(new_n20479_));
  NOR2_X1    g18043(.A1(new_n20479_), .A2(new_n20473_), .ZN(new_n20480_));
  INV_X1     g18044(.I(new_n20480_), .ZN(new_n20481_));
  AOI21_X1   g18045(.A1(new_n20481_), .A2(new_n12783_), .B(pi1154), .ZN(new_n20482_));
  AOI21_X1   g18046(.A1(new_n20481_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n20483_));
  NOR3_X1    g18047(.A1(new_n20482_), .A2(new_n20483_), .A3(new_n12779_), .ZN(new_n20484_));
  AOI21_X1   g18048(.A1(new_n12779_), .A2(new_n20481_), .B(new_n20484_), .ZN(new_n20485_));
  OAI21_X1   g18049(.A1(new_n20485_), .A2(new_n17229_), .B(new_n12791_), .ZN(new_n20486_));
  OAI21_X1   g18050(.A1(new_n20485_), .A2(new_n17232_), .B(pi1159), .ZN(new_n20487_));
  NAND3_X1   g18051(.A1(new_n20486_), .A2(new_n20487_), .A3(pi0789), .ZN(new_n20488_));
  OAI21_X1   g18052(.A1(pi0789), .A2(new_n20485_), .B(new_n20488_), .ZN(new_n20489_));
  INV_X1     g18053(.I(new_n20471_), .ZN(new_n20490_));
  NAND2_X1   g18054(.A1(new_n12818_), .A2(new_n20490_), .ZN(new_n20491_));
  OAI21_X1   g18055(.A1(new_n20489_), .A2(new_n12818_), .B(new_n20491_), .ZN(new_n20492_));
  AOI21_X1   g18056(.A1(new_n12826_), .A2(new_n16168_), .B(new_n20471_), .ZN(new_n20493_));
  NOR2_X1    g18057(.A1(new_n20471_), .A2(pi1153), .ZN(new_n20494_));
  NOR2_X1    g18058(.A1(new_n12834_), .A2(pi0725), .ZN(new_n20495_));
  INV_X1     g18059(.I(new_n20495_), .ZN(new_n20496_));
  NAND2_X1   g18060(.A1(new_n20496_), .A2(new_n20494_), .ZN(new_n20497_));
  NOR2_X1    g18061(.A1(new_n20495_), .A2(new_n20493_), .ZN(new_n20498_));
  NOR2_X1    g18062(.A1(new_n20498_), .A2(new_n12841_), .ZN(new_n20499_));
  INV_X1     g18063(.I(new_n20499_), .ZN(new_n20500_));
  NAND3_X1   g18064(.A1(new_n20500_), .A2(pi0778), .A3(new_n20497_), .ZN(new_n20501_));
  OAI21_X1   g18065(.A1(pi0778), .A2(new_n20493_), .B(new_n20501_), .ZN(new_n20502_));
  NAND2_X1   g18066(.A1(new_n20502_), .A2(new_n17187_), .ZN(new_n20503_));
  NOR2_X1    g18067(.A1(new_n20503_), .A2(new_n12889_), .ZN(new_n20504_));
  NAND2_X1   g18068(.A1(new_n20504_), .A2(new_n18203_), .ZN(new_n20505_));
  NOR2_X1    g18069(.A1(new_n20505_), .A2(new_n17884_), .ZN(new_n20506_));
  INV_X1     g18070(.I(new_n20506_), .ZN(new_n20507_));
  OAI22_X1   g18071(.A1(new_n20492_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n20507_), .ZN(new_n20508_));
  AND2_X2    g18072(.A1(new_n20508_), .A2(new_n12919_), .Z(new_n20509_));
  OAI22_X1   g18073(.A1(new_n20492_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n20507_), .ZN(new_n20510_));
  AOI21_X1   g18074(.A1(pi0629), .A2(new_n20510_), .B(new_n20509_), .ZN(new_n20511_));
  INV_X1     g18075(.I(new_n20478_), .ZN(new_n20512_));
  NOR2_X1    g18076(.A1(new_n20493_), .A2(new_n12754_), .ZN(new_n20513_));
  NOR3_X1    g18077(.A1(new_n20513_), .A2(new_n20470_), .A3(new_n20471_), .ZN(new_n20514_));
  NAND2_X1   g18078(.A1(new_n20514_), .A2(new_n12758_), .ZN(new_n20515_));
  NAND2_X1   g18079(.A1(new_n20513_), .A2(pi0625), .ZN(new_n20516_));
  NAND3_X1   g18080(.A1(new_n20516_), .A2(pi1153), .A3(new_n20472_), .ZN(new_n20517_));
  NAND3_X1   g18081(.A1(new_n20497_), .A2(pi0608), .A3(new_n20517_), .ZN(new_n20518_));
  INV_X1     g18082(.I(new_n20516_), .ZN(new_n20519_));
  OAI21_X1   g18083(.A1(new_n20519_), .A2(new_n20514_), .B(new_n20494_), .ZN(new_n20520_));
  NAND3_X1   g18084(.A1(new_n20500_), .A2(new_n13560_), .A3(new_n20520_), .ZN(new_n20521_));
  NAND3_X1   g18085(.A1(new_n20521_), .A2(pi0778), .A3(new_n20518_), .ZN(new_n20522_));
  AOI21_X1   g18086(.A1(new_n20522_), .A2(new_n20515_), .B(new_n12766_), .ZN(new_n20523_));
  NOR2_X1    g18087(.A1(new_n20502_), .A2(pi0609), .ZN(new_n20524_));
  OAI21_X1   g18088(.A1(new_n20524_), .A2(new_n20523_), .B(pi1155), .ZN(new_n20525_));
  NAND3_X1   g18089(.A1(new_n20525_), .A2(pi0660), .A3(new_n20512_), .ZN(new_n20526_));
  NAND2_X1   g18090(.A1(new_n20522_), .A2(new_n20515_), .ZN(new_n20527_));
  NOR2_X1    g18091(.A1(new_n20502_), .A2(new_n12766_), .ZN(new_n20528_));
  AOI21_X1   g18092(.A1(new_n20527_), .A2(new_n12766_), .B(new_n20528_), .ZN(new_n20529_));
  NOR2_X1    g18093(.A1(new_n20477_), .A2(pi0660), .ZN(new_n20530_));
  OAI21_X1   g18094(.A1(new_n20529_), .A2(pi1155), .B(new_n20530_), .ZN(new_n20531_));
  NAND3_X1   g18095(.A1(new_n20531_), .A2(new_n20526_), .A3(pi0785), .ZN(new_n20532_));
  NAND2_X1   g18096(.A1(new_n20527_), .A2(new_n12764_), .ZN(new_n20533_));
  NAND2_X1   g18097(.A1(new_n20532_), .A2(new_n20533_), .ZN(new_n20534_));
  NAND2_X1   g18098(.A1(new_n20534_), .A2(new_n12781_), .ZN(new_n20535_));
  NAND2_X1   g18099(.A1(new_n20503_), .A2(pi0618), .ZN(new_n20536_));
  AOI21_X1   g18100(.A1(new_n20535_), .A2(new_n20536_), .B(pi1154), .ZN(new_n20537_));
  NOR3_X1    g18101(.A1(new_n20537_), .A2(pi0627), .A3(new_n20483_), .ZN(new_n20538_));
  NAND2_X1   g18102(.A1(new_n20503_), .A2(new_n12781_), .ZN(new_n20539_));
  NAND2_X1   g18103(.A1(new_n20534_), .A2(pi0618), .ZN(new_n20540_));
  AOI21_X1   g18104(.A1(new_n20540_), .A2(new_n20539_), .B(new_n12785_), .ZN(new_n20541_));
  NOR3_X1    g18105(.A1(new_n20541_), .A2(new_n12880_), .A3(new_n20482_), .ZN(new_n20542_));
  OR3_X2     g18106(.A1(new_n20538_), .A2(new_n20542_), .A3(new_n12779_), .Z(new_n20543_));
  NAND2_X1   g18107(.A1(new_n20534_), .A2(new_n12779_), .ZN(new_n20544_));
  NAND2_X1   g18108(.A1(new_n20543_), .A2(new_n20544_), .ZN(new_n20545_));
  AOI21_X1   g18109(.A1(new_n20545_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n20546_));
  NOR2_X1    g18110(.A1(new_n20504_), .A2(pi0619), .ZN(new_n20547_));
  AOI21_X1   g18111(.A1(new_n20543_), .A2(new_n20544_), .B(new_n12793_), .ZN(new_n20548_));
  OAI21_X1   g18112(.A1(new_n20548_), .A2(new_n20547_), .B(pi1159), .ZN(new_n20549_));
  NAND3_X1   g18113(.A1(new_n20549_), .A2(pi0648), .A3(new_n20486_), .ZN(new_n20550_));
  NAND2_X1   g18114(.A1(new_n20545_), .A2(new_n12793_), .ZN(new_n20551_));
  OAI21_X1   g18115(.A1(new_n12793_), .A2(new_n20504_), .B(new_n20551_), .ZN(new_n20552_));
  NAND2_X1   g18116(.A1(new_n20552_), .A2(new_n12791_), .ZN(new_n20553_));
  NAND3_X1   g18117(.A1(new_n20553_), .A2(new_n12895_), .A3(new_n20487_), .ZN(new_n20554_));
  NAND3_X1   g18118(.A1(new_n20554_), .A2(pi0789), .A3(new_n20550_), .ZN(new_n20555_));
  NOR2_X1    g18119(.A1(new_n20490_), .A2(new_n12747_), .ZN(new_n20556_));
  AND2_X2    g18120(.A1(new_n20489_), .A2(new_n12747_), .Z(new_n20557_));
  OAI21_X1   g18121(.A1(new_n20557_), .A2(new_n20556_), .B(new_n12815_), .ZN(new_n20558_));
  INV_X1     g18122(.I(new_n20505_), .ZN(new_n20559_));
  NAND2_X1   g18123(.A1(new_n20489_), .A2(pi0626), .ZN(new_n20560_));
  OAI21_X1   g18124(.A1(pi0626), .A2(new_n20490_), .B(new_n20560_), .ZN(new_n20561_));
  AOI22_X1   g18125(.A1(new_n20561_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n20559_), .ZN(new_n20562_));
  NAND2_X1   g18126(.A1(new_n20562_), .A2(new_n20558_), .ZN(new_n20563_));
  AOI22_X1   g18127(.A1(new_n20555_), .A2(new_n20546_), .B1(pi0788), .B2(new_n20563_), .ZN(new_n20564_));
  OAI22_X1   g18128(.A1(new_n20564_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n20511_), .ZN(new_n20565_));
  NAND2_X1   g18129(.A1(new_n20492_), .A2(new_n13384_), .ZN(new_n20566_));
  NAND2_X1   g18130(.A1(new_n12943_), .A2(new_n20490_), .ZN(new_n20567_));
  NAND2_X1   g18131(.A1(new_n20566_), .A2(new_n20567_), .ZN(new_n20568_));
  NOR2_X1    g18132(.A1(new_n20507_), .A2(new_n12953_), .ZN(new_n20569_));
  NOR2_X1    g18133(.A1(new_n20569_), .A2(pi0647), .ZN(new_n20570_));
  NOR2_X1    g18134(.A1(new_n20471_), .A2(new_n12741_), .ZN(new_n20571_));
  OAI21_X1   g18135(.A1(new_n20570_), .A2(new_n20571_), .B(new_n12965_), .ZN(new_n20572_));
  NAND2_X1   g18136(.A1(new_n20569_), .A2(pi0647), .ZN(new_n20573_));
  OAI21_X1   g18137(.A1(pi0647), .A2(new_n20490_), .B(new_n20573_), .ZN(new_n20574_));
  OAI22_X1   g18138(.A1(new_n20574_), .A2(new_n15576_), .B1(new_n20572_), .B2(new_n12981_), .ZN(new_n20575_));
  AOI21_X1   g18139(.A1(new_n20568_), .A2(new_n15608_), .B(new_n20575_), .ZN(new_n20576_));
  OAI22_X1   g18140(.A1(new_n20565_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n20576_), .ZN(new_n20577_));
  NAND2_X1   g18141(.A1(new_n20577_), .A2(new_n13000_), .ZN(new_n20578_));
  AND2_X2    g18142(.A1(new_n20577_), .A2(new_n12975_), .Z(new_n20579_));
  OAI21_X1   g18143(.A1(new_n20574_), .A2(new_n12965_), .B(new_n20572_), .ZN(new_n20580_));
  NAND2_X1   g18144(.A1(new_n20569_), .A2(new_n12972_), .ZN(new_n20581_));
  OAI21_X1   g18145(.A1(new_n20580_), .A2(new_n12972_), .B(new_n20581_), .ZN(new_n20582_));
  NOR2_X1    g18146(.A1(new_n20582_), .A2(new_n12975_), .ZN(new_n20583_));
  OAI21_X1   g18147(.A1(new_n20579_), .A2(new_n20583_), .B(new_n12740_), .ZN(new_n20584_));
  NAND2_X1   g18148(.A1(new_n20490_), .A2(pi0644), .ZN(new_n20585_));
  NOR2_X1    g18149(.A1(new_n17611_), .A2(new_n20471_), .ZN(new_n20586_));
  AOI21_X1   g18150(.A1(new_n20492_), .A2(new_n17611_), .B(new_n20586_), .ZN(new_n20587_));
  OAI21_X1   g18151(.A1(new_n20587_), .A2(pi0644), .B(new_n20585_), .ZN(new_n20588_));
  NAND2_X1   g18152(.A1(new_n20588_), .A2(pi0715), .ZN(new_n20589_));
  NAND3_X1   g18153(.A1(new_n20584_), .A2(new_n12739_), .A3(new_n20589_), .ZN(new_n20590_));
  NOR2_X1    g18154(.A1(new_n20582_), .A2(pi0644), .ZN(new_n20591_));
  AOI21_X1   g18155(.A1(new_n20577_), .A2(pi0644), .B(new_n20591_), .ZN(new_n20592_));
  NAND2_X1   g18156(.A1(new_n20490_), .A2(new_n12975_), .ZN(new_n20593_));
  OAI21_X1   g18157(.A1(new_n20587_), .A2(new_n12975_), .B(new_n20593_), .ZN(new_n20594_));
  AOI21_X1   g18158(.A1(new_n20594_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n20595_));
  OAI21_X1   g18159(.A1(new_n20592_), .A2(new_n12740_), .B(new_n20595_), .ZN(new_n20596_));
  NAND3_X1   g18160(.A1(new_n20590_), .A2(pi0790), .A3(new_n20596_), .ZN(new_n20597_));
  NAND2_X1   g18161(.A1(new_n20597_), .A2(new_n20578_), .ZN(new_n20598_));
  AOI21_X1   g18162(.A1(po1038), .A2(new_n7479_), .B(pi0832), .ZN(new_n20599_));
  NAND2_X1   g18163(.A1(new_n13192_), .A2(new_n7479_), .ZN(new_n20600_));
  INV_X1     g18164(.I(new_n20600_), .ZN(new_n20601_));
  AOI21_X1   g18165(.A1(new_n20601_), .A2(pi0644), .B(new_n12740_), .ZN(new_n20602_));
  NAND2_X1   g18166(.A1(new_n20600_), .A2(new_n12984_), .ZN(new_n20603_));
  NOR2_X1    g18167(.A1(new_n20601_), .A2(new_n13384_), .ZN(new_n20604_));
  NOR2_X1    g18168(.A1(new_n2609_), .A2(new_n7479_), .ZN(new_n20605_));
  NOR2_X1    g18169(.A1(new_n13342_), .A2(pi0755), .ZN(new_n20606_));
  NOR2_X1    g18170(.A1(new_n13344_), .A2(pi0183), .ZN(new_n20607_));
  NOR3_X1    g18171(.A1(new_n20606_), .A2(new_n3265_), .A3(new_n20607_), .ZN(new_n20608_));
  NAND2_X1   g18172(.A1(new_n13334_), .A2(new_n7479_), .ZN(new_n20609_));
  NAND2_X1   g18173(.A1(new_n13245_), .A2(pi0183), .ZN(new_n20610_));
  AOI21_X1   g18174(.A1(new_n20609_), .A2(new_n20610_), .B(pi0755), .ZN(new_n20611_));
  NOR3_X1    g18175(.A1(new_n15787_), .A2(pi0183), .A3(new_n16169_), .ZN(new_n20612_));
  NOR2_X1    g18176(.A1(new_n20611_), .A2(new_n20612_), .ZN(new_n20613_));
  AOI21_X1   g18177(.A1(new_n20613_), .A2(new_n3265_), .B(new_n20608_), .ZN(new_n20614_));
  NOR2_X1    g18178(.A1(new_n20614_), .A2(new_n2610_), .ZN(new_n20615_));
  NOR2_X1    g18179(.A1(new_n20615_), .A2(new_n20605_), .ZN(new_n20616_));
  NOR2_X1    g18180(.A1(new_n20616_), .A2(new_n12760_), .ZN(new_n20617_));
  INV_X1     g18181(.I(new_n20617_), .ZN(new_n20618_));
  OAI21_X1   g18182(.A1(new_n12761_), .A2(new_n20601_), .B(new_n20618_), .ZN(new_n20619_));
  OAI22_X1   g18183(.A1(new_n20618_), .A2(pi0609), .B1(new_n13353_), .B2(new_n20601_), .ZN(new_n20620_));
  NAND2_X1   g18184(.A1(new_n20620_), .A2(new_n12770_), .ZN(new_n20621_));
  INV_X1     g18185(.I(new_n20621_), .ZN(new_n20622_));
  AOI22_X1   g18186(.A1(new_n20617_), .A2(pi0609), .B1(new_n13357_), .B2(new_n20600_), .ZN(new_n20623_));
  OAI21_X1   g18187(.A1(new_n20623_), .A2(new_n12770_), .B(pi0785), .ZN(new_n20624_));
  OAI22_X1   g18188(.A1(new_n20622_), .A2(new_n20624_), .B1(pi0785), .B2(new_n20619_), .ZN(new_n20625_));
  NAND2_X1   g18189(.A1(new_n20625_), .A2(new_n12779_), .ZN(new_n20626_));
  NAND2_X1   g18190(.A1(new_n20600_), .A2(pi0618), .ZN(new_n20627_));
  OAI21_X1   g18191(.A1(new_n20625_), .A2(pi0618), .B(new_n20627_), .ZN(new_n20628_));
  NAND2_X1   g18192(.A1(new_n20628_), .A2(new_n12785_), .ZN(new_n20629_));
  NAND2_X1   g18193(.A1(new_n20600_), .A2(new_n12781_), .ZN(new_n20630_));
  OAI21_X1   g18194(.A1(new_n20625_), .A2(new_n12781_), .B(new_n20630_), .ZN(new_n20631_));
  NAND2_X1   g18195(.A1(new_n20631_), .A2(pi1154), .ZN(new_n20632_));
  NAND3_X1   g18196(.A1(new_n20629_), .A2(new_n20632_), .A3(pi0781), .ZN(new_n20633_));
  NAND2_X1   g18197(.A1(new_n20633_), .A2(new_n20626_), .ZN(new_n20634_));
  NAND2_X1   g18198(.A1(new_n20634_), .A2(new_n12796_), .ZN(new_n20635_));
  NAND2_X1   g18199(.A1(new_n20600_), .A2(pi0619), .ZN(new_n20636_));
  OAI21_X1   g18200(.A1(new_n20634_), .A2(pi0619), .B(new_n20636_), .ZN(new_n20637_));
  NAND2_X1   g18201(.A1(new_n20637_), .A2(new_n12791_), .ZN(new_n20638_));
  NAND2_X1   g18202(.A1(new_n20600_), .A2(new_n12793_), .ZN(new_n20639_));
  OAI21_X1   g18203(.A1(new_n20634_), .A2(new_n12793_), .B(new_n20639_), .ZN(new_n20640_));
  NAND2_X1   g18204(.A1(new_n20640_), .A2(pi1159), .ZN(new_n20641_));
  NAND3_X1   g18205(.A1(new_n20638_), .A2(new_n20641_), .A3(pi0789), .ZN(new_n20642_));
  NAND2_X1   g18206(.A1(new_n20642_), .A2(new_n20635_), .ZN(new_n20643_));
  NAND2_X1   g18207(.A1(new_n20600_), .A2(new_n12818_), .ZN(new_n20644_));
  OAI21_X1   g18208(.A1(new_n20643_), .A2(new_n12818_), .B(new_n20644_), .ZN(new_n20645_));
  AOI21_X1   g18209(.A1(new_n20645_), .A2(new_n13384_), .B(new_n20604_), .ZN(new_n20646_));
  OAI21_X1   g18210(.A1(new_n20646_), .A2(new_n12984_), .B(new_n20603_), .ZN(new_n20647_));
  OAI21_X1   g18211(.A1(new_n20647_), .A2(pi0644), .B(new_n20602_), .ZN(new_n20648_));
  AND2_X2    g18212(.A1(new_n20648_), .A2(new_n12739_), .Z(new_n20649_));
  OAI21_X1   g18213(.A1(new_n14125_), .A2(new_n20607_), .B(new_n16168_), .ZN(new_n20650_));
  OAI21_X1   g18214(.A1(new_n14122_), .A2(new_n7479_), .B(new_n3265_), .ZN(new_n20651_));
  NAND2_X1   g18215(.A1(new_n20651_), .A2(new_n2609_), .ZN(new_n20652_));
  NAND2_X1   g18216(.A1(new_n15744_), .A2(new_n7479_), .ZN(new_n20653_));
  AOI21_X1   g18217(.A1(new_n20653_), .A2(new_n20652_), .B(new_n20650_), .ZN(new_n20654_));
  NAND2_X1   g18218(.A1(new_n2609_), .A2(new_n16168_), .ZN(new_n20655_));
  AOI21_X1   g18219(.A1(new_n20601_), .A2(new_n20655_), .B(new_n20654_), .ZN(new_n20656_));
  NAND2_X1   g18220(.A1(new_n20656_), .A2(new_n13521_), .ZN(new_n20657_));
  NAND2_X1   g18221(.A1(new_n20600_), .A2(pi0625), .ZN(new_n20658_));
  AOI21_X1   g18222(.A1(new_n20657_), .A2(new_n20658_), .B(pi1153), .ZN(new_n20659_));
  NAND2_X1   g18223(.A1(new_n20600_), .A2(new_n13521_), .ZN(new_n20660_));
  NAND2_X1   g18224(.A1(new_n20656_), .A2(pi0625), .ZN(new_n20661_));
  AOI21_X1   g18225(.A1(new_n20661_), .A2(new_n20660_), .B(new_n12841_), .ZN(new_n20662_));
  NOR3_X1    g18226(.A1(new_n20659_), .A2(new_n20662_), .A3(new_n12758_), .ZN(new_n20663_));
  NOR2_X1    g18227(.A1(new_n20656_), .A2(pi0778), .ZN(new_n20664_));
  NOR2_X1    g18228(.A1(new_n20663_), .A2(new_n20664_), .ZN(new_n20665_));
  NOR2_X1    g18229(.A1(new_n20665_), .A2(new_n12869_), .ZN(new_n20666_));
  AOI21_X1   g18230(.A1(new_n12869_), .A2(new_n20601_), .B(new_n20666_), .ZN(new_n20667_));
  NAND2_X1   g18231(.A1(new_n20667_), .A2(new_n12888_), .ZN(new_n20668_));
  OAI21_X1   g18232(.A1(new_n12888_), .A2(new_n20601_), .B(new_n20668_), .ZN(new_n20669_));
  INV_X1     g18233(.I(new_n20669_), .ZN(new_n20670_));
  NOR2_X1    g18234(.A1(new_n20600_), .A2(new_n12911_), .ZN(new_n20671_));
  AOI21_X1   g18235(.A1(new_n20670_), .A2(new_n12911_), .B(new_n20671_), .ZN(new_n20672_));
  NAND2_X1   g18236(.A1(new_n20672_), .A2(new_n13392_), .ZN(new_n20673_));
  OAI21_X1   g18237(.A1(new_n13392_), .A2(new_n20601_), .B(new_n20673_), .ZN(new_n20674_));
  NAND2_X1   g18238(.A1(new_n20674_), .A2(new_n12920_), .ZN(new_n20675_));
  NAND2_X1   g18239(.A1(new_n20600_), .A2(pi0628), .ZN(new_n20676_));
  AOI21_X1   g18240(.A1(new_n20675_), .A2(new_n20676_), .B(pi1156), .ZN(new_n20677_));
  NAND2_X1   g18241(.A1(new_n20600_), .A2(new_n12920_), .ZN(new_n20678_));
  NAND2_X1   g18242(.A1(new_n20674_), .A2(pi0628), .ZN(new_n20679_));
  AOI21_X1   g18243(.A1(new_n20679_), .A2(new_n20678_), .B(new_n12742_), .ZN(new_n20680_));
  OR2_X2     g18244(.A1(new_n20680_), .A2(new_n12937_), .Z(new_n20681_));
  OAI22_X1   g18245(.A1(new_n20681_), .A2(new_n20677_), .B1(pi0792), .B2(new_n20674_), .ZN(new_n20682_));
  NAND2_X1   g18246(.A1(new_n20682_), .A2(new_n12741_), .ZN(new_n20683_));
  OAI21_X1   g18247(.A1(new_n12741_), .A2(new_n20600_), .B(new_n20683_), .ZN(new_n20684_));
  NOR2_X1    g18248(.A1(new_n20684_), .A2(pi1157), .ZN(new_n20685_));
  NAND2_X1   g18249(.A1(new_n20682_), .A2(pi0647), .ZN(new_n20686_));
  OAI21_X1   g18250(.A1(pi0647), .A2(new_n20600_), .B(new_n20686_), .ZN(new_n20687_));
  NOR2_X1    g18251(.A1(new_n20687_), .A2(new_n12965_), .ZN(new_n20688_));
  OAI21_X1   g18252(.A1(new_n20685_), .A2(new_n20688_), .B(pi0787), .ZN(new_n20689_));
  OAI21_X1   g18253(.A1(pi0787), .A2(new_n20682_), .B(new_n20689_), .ZN(new_n20690_));
  OAI21_X1   g18254(.A1(new_n20690_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n20691_));
  AOI21_X1   g18255(.A1(new_n20601_), .A2(new_n12975_), .B(pi0715), .ZN(new_n20692_));
  OAI21_X1   g18256(.A1(new_n20647_), .A2(new_n12975_), .B(new_n20692_), .ZN(new_n20693_));
  AND2_X2    g18257(.A1(new_n20693_), .A2(pi1160), .Z(new_n20694_));
  OAI21_X1   g18258(.A1(new_n20690_), .A2(pi0644), .B(pi0715), .ZN(new_n20695_));
  AOI22_X1   g18259(.A1(new_n20649_), .A2(new_n20691_), .B1(new_n20695_), .B2(new_n20694_), .ZN(new_n20696_));
  NOR2_X1    g18260(.A1(new_n20696_), .A2(new_n13000_), .ZN(new_n20697_));
  NAND2_X1   g18261(.A1(new_n20601_), .A2(pi0626), .ZN(new_n20698_));
  NAND2_X1   g18262(.A1(new_n20643_), .A2(new_n12747_), .ZN(new_n20699_));
  AOI21_X1   g18263(.A1(new_n20699_), .A2(new_n20698_), .B(new_n12816_), .ZN(new_n20700_));
  NOR2_X1    g18264(.A1(new_n20600_), .A2(pi0626), .ZN(new_n20701_));
  AOI21_X1   g18265(.A1(new_n20643_), .A2(pi0626), .B(new_n20701_), .ZN(new_n20702_));
  OAI22_X1   g18266(.A1(new_n20702_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n20672_), .ZN(new_n20703_));
  OAI21_X1   g18267(.A1(new_n20703_), .A2(new_n20700_), .B(pi0788), .ZN(new_n20704_));
  NAND2_X1   g18268(.A1(new_n20704_), .A2(new_n15824_), .ZN(new_n20705_));
  NAND2_X1   g18269(.A1(new_n20665_), .A2(new_n12766_), .ZN(new_n20706_));
  AOI21_X1   g18270(.A1(new_n16169_), .A2(new_n13566_), .B(new_n15826_), .ZN(new_n20707_));
  AOI21_X1   g18271(.A1(new_n14328_), .A2(new_n20474_), .B(new_n7479_), .ZN(new_n20708_));
  AOI21_X1   g18272(.A1(new_n20708_), .A2(new_n5336_), .B(new_n3265_), .ZN(new_n20709_));
  OAI21_X1   g18273(.A1(new_n20707_), .A2(pi0183), .B(new_n20709_), .ZN(new_n20710_));
  NAND2_X1   g18274(.A1(new_n14172_), .A2(pi0183), .ZN(new_n20711_));
  NAND2_X1   g18275(.A1(new_n14174_), .A2(new_n7479_), .ZN(new_n20712_));
  AOI21_X1   g18276(.A1(new_n20711_), .A2(new_n20712_), .B(pi0755), .ZN(new_n20713_));
  NAND2_X1   g18277(.A1(new_n15835_), .A2(pi0183), .ZN(new_n20714_));
  NAND2_X1   g18278(.A1(new_n14177_), .A2(new_n7479_), .ZN(new_n20715_));
  AOI21_X1   g18279(.A1(new_n20715_), .A2(new_n20714_), .B(new_n16169_), .ZN(new_n20716_));
  OAI21_X1   g18280(.A1(new_n20716_), .A2(new_n20713_), .B(new_n2627_), .ZN(new_n20717_));
  NOR2_X1    g18281(.A1(new_n14182_), .A2(pi0183), .ZN(new_n20718_));
  NOR2_X1    g18282(.A1(new_n14184_), .A2(new_n7479_), .ZN(new_n20719_));
  OAI21_X1   g18283(.A1(new_n20718_), .A2(new_n20719_), .B(pi0755), .ZN(new_n20720_));
  NOR2_X1    g18284(.A1(new_n14187_), .A2(new_n7479_), .ZN(new_n20721_));
  NOR2_X1    g18285(.A1(new_n14189_), .A2(pi0183), .ZN(new_n20722_));
  OAI21_X1   g18286(.A1(new_n20721_), .A2(new_n20722_), .B(new_n16169_), .ZN(new_n20723_));
  NAND3_X1   g18287(.A1(new_n20723_), .A2(new_n20720_), .A3(pi0039), .ZN(new_n20724_));
  NAND3_X1   g18288(.A1(new_n20724_), .A2(new_n3265_), .A3(new_n20717_), .ZN(new_n20725_));
  NAND3_X1   g18289(.A1(new_n20725_), .A2(new_n16168_), .A3(new_n20710_), .ZN(new_n20726_));
  NAND2_X1   g18290(.A1(new_n20614_), .A2(pi0725), .ZN(new_n20727_));
  NAND3_X1   g18291(.A1(new_n20726_), .A2(new_n2609_), .A3(new_n20727_), .ZN(new_n20728_));
  OAI21_X1   g18292(.A1(new_n7479_), .A2(new_n2609_), .B(new_n20728_), .ZN(new_n20729_));
  INV_X1     g18293(.I(new_n20662_), .ZN(new_n20730_));
  NOR2_X1    g18294(.A1(new_n20616_), .A2(new_n13521_), .ZN(new_n20731_));
  AOI21_X1   g18295(.A1(new_n20729_), .A2(new_n13521_), .B(new_n20731_), .ZN(new_n20732_));
  OAI21_X1   g18296(.A1(new_n20732_), .A2(pi1153), .B(new_n20730_), .ZN(new_n20733_));
  NOR2_X1    g18297(.A1(new_n20616_), .A2(pi0625), .ZN(new_n20734_));
  AOI21_X1   g18298(.A1(new_n20729_), .A2(pi0625), .B(new_n20734_), .ZN(new_n20735_));
  OAI21_X1   g18299(.A1(new_n20735_), .A2(new_n12841_), .B(pi0608), .ZN(new_n20736_));
  OAI22_X1   g18300(.A1(pi0608), .A2(new_n20733_), .B1(new_n20736_), .B2(new_n20659_), .ZN(new_n20737_));
  NOR2_X1    g18301(.A1(new_n20737_), .A2(new_n12758_), .ZN(new_n20738_));
  AOI21_X1   g18302(.A1(new_n12758_), .A2(new_n20729_), .B(new_n20738_), .ZN(new_n20739_));
  OAI21_X1   g18303(.A1(new_n20739_), .A2(new_n12766_), .B(new_n20706_), .ZN(new_n20740_));
  AOI21_X1   g18304(.A1(new_n20740_), .A2(pi1155), .B(new_n20622_), .ZN(new_n20741_));
  NOR2_X1    g18305(.A1(new_n20739_), .A2(pi0609), .ZN(new_n20742_));
  NOR3_X1    g18306(.A1(new_n20663_), .A2(new_n12766_), .A3(new_n20664_), .ZN(new_n20743_));
  OAI21_X1   g18307(.A1(new_n20742_), .A2(new_n20743_), .B(new_n12770_), .ZN(new_n20744_));
  NOR2_X1    g18308(.A1(new_n20623_), .A2(new_n12770_), .ZN(new_n20745_));
  NOR2_X1    g18309(.A1(new_n20745_), .A2(pi0660), .ZN(new_n20746_));
  AOI22_X1   g18310(.A1(new_n20741_), .A2(pi0660), .B1(new_n20744_), .B2(new_n20746_), .ZN(new_n20747_));
  NOR2_X1    g18311(.A1(new_n20739_), .A2(pi0785), .ZN(new_n20748_));
  AOI21_X1   g18312(.A1(new_n20747_), .A2(pi0785), .B(new_n20748_), .ZN(new_n20749_));
  NOR2_X1    g18313(.A1(new_n20749_), .A2(pi0781), .ZN(new_n20750_));
  AND2_X2    g18314(.A1(new_n20667_), .A2(new_n12781_), .Z(new_n20751_));
  NOR2_X1    g18315(.A1(new_n20749_), .A2(new_n12781_), .ZN(new_n20752_));
  OAI21_X1   g18316(.A1(new_n20752_), .A2(new_n20751_), .B(pi1154), .ZN(new_n20753_));
  NAND3_X1   g18317(.A1(new_n20753_), .A2(pi0627), .A3(new_n20629_), .ZN(new_n20754_));
  INV_X1     g18318(.I(new_n20632_), .ZN(new_n20755_));
  NAND2_X1   g18319(.A1(new_n20667_), .A2(pi0618), .ZN(new_n20756_));
  OAI21_X1   g18320(.A1(new_n20749_), .A2(pi0618), .B(new_n20756_), .ZN(new_n20757_));
  AOI21_X1   g18321(.A1(new_n20757_), .A2(new_n12785_), .B(new_n20755_), .ZN(new_n20758_));
  AOI21_X1   g18322(.A1(new_n20758_), .A2(new_n12880_), .B(new_n12779_), .ZN(new_n20759_));
  AOI21_X1   g18323(.A1(new_n20759_), .A2(new_n20754_), .B(new_n20750_), .ZN(new_n20760_));
  OAI21_X1   g18324(.A1(new_n20760_), .A2(pi0789), .B(new_n12819_), .ZN(new_n20761_));
  NOR2_X1    g18325(.A1(new_n20670_), .A2(new_n12793_), .ZN(new_n20762_));
  NOR2_X1    g18326(.A1(new_n20760_), .A2(pi0619), .ZN(new_n20763_));
  OAI21_X1   g18327(.A1(new_n20763_), .A2(new_n20762_), .B(new_n12791_), .ZN(new_n20764_));
  NAND3_X1   g18328(.A1(new_n20764_), .A2(new_n12895_), .A3(new_n20641_), .ZN(new_n20765_));
  NAND2_X1   g18329(.A1(new_n20669_), .A2(new_n12793_), .ZN(new_n20766_));
  OAI21_X1   g18330(.A1(new_n20760_), .A2(new_n12793_), .B(new_n20766_), .ZN(new_n20767_));
  AOI21_X1   g18331(.A1(new_n20767_), .A2(pi1159), .B(new_n12895_), .ZN(new_n20768_));
  AOI21_X1   g18332(.A1(new_n20768_), .A2(new_n20638_), .B(new_n12796_), .ZN(new_n20769_));
  AOI21_X1   g18333(.A1(new_n20769_), .A2(new_n20765_), .B(new_n20761_), .ZN(new_n20770_));
  NOR2_X1    g18334(.A1(new_n20680_), .A2(pi0629), .ZN(new_n20771_));
  NOR2_X1    g18335(.A1(new_n20677_), .A2(new_n12919_), .ZN(new_n20772_));
  NOR2_X1    g18336(.A1(new_n20771_), .A2(new_n20772_), .ZN(new_n20773_));
  AOI21_X1   g18337(.A1(new_n20645_), .A2(new_n19160_), .B(new_n20773_), .ZN(new_n20774_));
  OAI22_X1   g18338(.A1(new_n20770_), .A2(new_n20705_), .B1(new_n12937_), .B2(new_n20774_), .ZN(new_n20775_));
  NOR2_X1    g18339(.A1(new_n20694_), .A2(new_n12975_), .ZN(new_n20776_));
  NOR2_X1    g18340(.A1(new_n20649_), .A2(pi0644), .ZN(new_n20777_));
  NOR2_X1    g18341(.A1(new_n20776_), .A2(new_n20777_), .ZN(new_n20778_));
  OAI22_X1   g18342(.A1(new_n15576_), .A2(new_n20687_), .B1(new_n20684_), .B2(new_n15730_), .ZN(new_n20779_));
  NOR2_X1    g18343(.A1(new_n20646_), .A2(new_n17212_), .ZN(new_n20780_));
  NOR2_X1    g18344(.A1(new_n20779_), .A2(new_n20780_), .ZN(new_n20781_));
  OAI22_X1   g18345(.A1(new_n20778_), .A2(new_n13000_), .B1(new_n20781_), .B2(new_n12972_), .ZN(new_n20782_));
  AOI21_X1   g18346(.A1(new_n15693_), .A2(new_n20775_), .B(new_n20782_), .ZN(new_n20783_));
  OAI21_X1   g18347(.A1(new_n20697_), .A2(new_n20783_), .B(new_n6643_), .ZN(new_n20784_));
  AOI22_X1   g18348(.A1(new_n20784_), .A2(new_n20599_), .B1(pi0832), .B2(new_n20598_), .ZN(po0340));
  NOR2_X1    g18349(.A1(new_n13340_), .A2(pi0777), .ZN(new_n20786_));
  NOR2_X1    g18350(.A1(new_n3042_), .A2(pi0184), .ZN(new_n20787_));
  NOR2_X1    g18351(.A1(new_n20786_), .A2(new_n20787_), .ZN(new_n20788_));
  NOR3_X1    g18352(.A1(new_n20788_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n20789_));
  INV_X1     g18353(.I(new_n20786_), .ZN(new_n20790_));
  NOR2_X1    g18354(.A1(new_n20790_), .A2(new_n13354_), .ZN(new_n20791_));
  NOR3_X1    g18355(.A1(new_n20791_), .A2(new_n12762_), .A3(new_n20788_), .ZN(new_n20792_));
  NOR2_X1    g18356(.A1(new_n20792_), .A2(new_n12770_), .ZN(new_n20793_));
  NOR3_X1    g18357(.A1(new_n20791_), .A2(pi1155), .A3(new_n20787_), .ZN(new_n20794_));
  NOR3_X1    g18358(.A1(new_n20793_), .A2(new_n12764_), .A3(new_n20794_), .ZN(new_n20795_));
  NOR2_X1    g18359(.A1(new_n20795_), .A2(new_n20789_), .ZN(new_n20796_));
  INV_X1     g18360(.I(new_n20796_), .ZN(new_n20797_));
  AOI21_X1   g18361(.A1(new_n20797_), .A2(new_n12783_), .B(pi1154), .ZN(new_n20798_));
  AOI21_X1   g18362(.A1(new_n20797_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n20799_));
  NOR3_X1    g18363(.A1(new_n20798_), .A2(new_n20799_), .A3(new_n12779_), .ZN(new_n20800_));
  AOI21_X1   g18364(.A1(new_n12779_), .A2(new_n20797_), .B(new_n20800_), .ZN(new_n20801_));
  OAI21_X1   g18365(.A1(new_n20801_), .A2(new_n17229_), .B(new_n12791_), .ZN(new_n20802_));
  OAI21_X1   g18366(.A1(new_n20801_), .A2(new_n17232_), .B(pi1159), .ZN(new_n20803_));
  NAND3_X1   g18367(.A1(new_n20802_), .A2(new_n20803_), .A3(pi0789), .ZN(new_n20804_));
  OAI21_X1   g18368(.A1(pi0789), .A2(new_n20801_), .B(new_n20804_), .ZN(new_n20805_));
  INV_X1     g18369(.I(new_n20787_), .ZN(new_n20806_));
  NAND2_X1   g18370(.A1(new_n12818_), .A2(new_n20806_), .ZN(new_n20807_));
  OAI21_X1   g18371(.A1(new_n20805_), .A2(new_n12818_), .B(new_n20807_), .ZN(new_n20808_));
  AOI21_X1   g18372(.A1(new_n12826_), .A2(new_n16756_), .B(new_n20787_), .ZN(new_n20809_));
  NOR2_X1    g18373(.A1(new_n20787_), .A2(pi1153), .ZN(new_n20810_));
  NOR2_X1    g18374(.A1(new_n12834_), .A2(pi0737), .ZN(new_n20811_));
  INV_X1     g18375(.I(new_n20811_), .ZN(new_n20812_));
  NAND2_X1   g18376(.A1(new_n20812_), .A2(new_n20810_), .ZN(new_n20813_));
  NOR2_X1    g18377(.A1(new_n20811_), .A2(new_n20809_), .ZN(new_n20814_));
  NOR2_X1    g18378(.A1(new_n20814_), .A2(new_n12841_), .ZN(new_n20815_));
  INV_X1     g18379(.I(new_n20815_), .ZN(new_n20816_));
  NAND3_X1   g18380(.A1(new_n20816_), .A2(pi0778), .A3(new_n20813_), .ZN(new_n20817_));
  OAI21_X1   g18381(.A1(pi0778), .A2(new_n20809_), .B(new_n20817_), .ZN(new_n20818_));
  NAND2_X1   g18382(.A1(new_n20818_), .A2(new_n17187_), .ZN(new_n20819_));
  NOR2_X1    g18383(.A1(new_n20819_), .A2(new_n12889_), .ZN(new_n20820_));
  NAND2_X1   g18384(.A1(new_n20820_), .A2(new_n18203_), .ZN(new_n20821_));
  NOR2_X1    g18385(.A1(new_n20821_), .A2(new_n17884_), .ZN(new_n20822_));
  INV_X1     g18386(.I(new_n20822_), .ZN(new_n20823_));
  OAI22_X1   g18387(.A1(new_n20808_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n20823_), .ZN(new_n20824_));
  AND2_X2    g18388(.A1(new_n20824_), .A2(new_n12919_), .Z(new_n20825_));
  OAI22_X1   g18389(.A1(new_n20808_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n20823_), .ZN(new_n20826_));
  AOI21_X1   g18390(.A1(pi0629), .A2(new_n20826_), .B(new_n20825_), .ZN(new_n20827_));
  INV_X1     g18391(.I(new_n20794_), .ZN(new_n20828_));
  NOR2_X1    g18392(.A1(new_n20809_), .A2(new_n12754_), .ZN(new_n20829_));
  NOR3_X1    g18393(.A1(new_n20829_), .A2(new_n20786_), .A3(new_n20787_), .ZN(new_n20830_));
  NAND2_X1   g18394(.A1(new_n20830_), .A2(new_n12758_), .ZN(new_n20831_));
  NAND2_X1   g18395(.A1(new_n20829_), .A2(pi0625), .ZN(new_n20832_));
  NAND3_X1   g18396(.A1(new_n20832_), .A2(pi1153), .A3(new_n20788_), .ZN(new_n20833_));
  NAND3_X1   g18397(.A1(new_n20813_), .A2(pi0608), .A3(new_n20833_), .ZN(new_n20834_));
  INV_X1     g18398(.I(new_n20832_), .ZN(new_n20835_));
  OAI21_X1   g18399(.A1(new_n20835_), .A2(new_n20830_), .B(new_n20810_), .ZN(new_n20836_));
  NAND3_X1   g18400(.A1(new_n20816_), .A2(new_n13560_), .A3(new_n20836_), .ZN(new_n20837_));
  NAND3_X1   g18401(.A1(new_n20837_), .A2(pi0778), .A3(new_n20834_), .ZN(new_n20838_));
  AOI21_X1   g18402(.A1(new_n20838_), .A2(new_n20831_), .B(new_n12766_), .ZN(new_n20839_));
  NOR2_X1    g18403(.A1(new_n20818_), .A2(pi0609), .ZN(new_n20840_));
  OAI21_X1   g18404(.A1(new_n20840_), .A2(new_n20839_), .B(pi1155), .ZN(new_n20841_));
  NAND3_X1   g18405(.A1(new_n20841_), .A2(pi0660), .A3(new_n20828_), .ZN(new_n20842_));
  NAND2_X1   g18406(.A1(new_n20838_), .A2(new_n20831_), .ZN(new_n20843_));
  NOR2_X1    g18407(.A1(new_n20818_), .A2(new_n12766_), .ZN(new_n20844_));
  AOI21_X1   g18408(.A1(new_n20843_), .A2(new_n12766_), .B(new_n20844_), .ZN(new_n20845_));
  NOR2_X1    g18409(.A1(new_n20793_), .A2(pi0660), .ZN(new_n20846_));
  OAI21_X1   g18410(.A1(new_n20845_), .A2(pi1155), .B(new_n20846_), .ZN(new_n20847_));
  NAND3_X1   g18411(.A1(new_n20847_), .A2(new_n20842_), .A3(pi0785), .ZN(new_n20848_));
  NAND2_X1   g18412(.A1(new_n20843_), .A2(new_n12764_), .ZN(new_n20849_));
  NAND2_X1   g18413(.A1(new_n20848_), .A2(new_n20849_), .ZN(new_n20850_));
  NAND2_X1   g18414(.A1(new_n20850_), .A2(new_n12781_), .ZN(new_n20851_));
  NAND2_X1   g18415(.A1(new_n20819_), .A2(pi0618), .ZN(new_n20852_));
  AOI21_X1   g18416(.A1(new_n20851_), .A2(new_n20852_), .B(pi1154), .ZN(new_n20853_));
  NOR3_X1    g18417(.A1(new_n20853_), .A2(pi0627), .A3(new_n20799_), .ZN(new_n20854_));
  NAND2_X1   g18418(.A1(new_n20819_), .A2(new_n12781_), .ZN(new_n20855_));
  NAND2_X1   g18419(.A1(new_n20850_), .A2(pi0618), .ZN(new_n20856_));
  AOI21_X1   g18420(.A1(new_n20856_), .A2(new_n20855_), .B(new_n12785_), .ZN(new_n20857_));
  NOR3_X1    g18421(.A1(new_n20857_), .A2(new_n12880_), .A3(new_n20798_), .ZN(new_n20858_));
  OR3_X2     g18422(.A1(new_n20854_), .A2(new_n20858_), .A3(new_n12779_), .Z(new_n20859_));
  NAND2_X1   g18423(.A1(new_n20850_), .A2(new_n12779_), .ZN(new_n20860_));
  NAND2_X1   g18424(.A1(new_n20859_), .A2(new_n20860_), .ZN(new_n20861_));
  AOI21_X1   g18425(.A1(new_n20861_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n20862_));
  NOR2_X1    g18426(.A1(new_n20820_), .A2(pi0619), .ZN(new_n20863_));
  AOI21_X1   g18427(.A1(new_n20859_), .A2(new_n20860_), .B(new_n12793_), .ZN(new_n20864_));
  OAI21_X1   g18428(.A1(new_n20864_), .A2(new_n20863_), .B(pi1159), .ZN(new_n20865_));
  NAND3_X1   g18429(.A1(new_n20865_), .A2(pi0648), .A3(new_n20802_), .ZN(new_n20866_));
  NAND2_X1   g18430(.A1(new_n20861_), .A2(new_n12793_), .ZN(new_n20867_));
  OAI21_X1   g18431(.A1(new_n12793_), .A2(new_n20820_), .B(new_n20867_), .ZN(new_n20868_));
  NAND2_X1   g18432(.A1(new_n20868_), .A2(new_n12791_), .ZN(new_n20869_));
  NAND3_X1   g18433(.A1(new_n20869_), .A2(new_n12895_), .A3(new_n20803_), .ZN(new_n20870_));
  NAND3_X1   g18434(.A1(new_n20870_), .A2(pi0789), .A3(new_n20866_), .ZN(new_n20871_));
  NOR2_X1    g18435(.A1(new_n20806_), .A2(new_n12747_), .ZN(new_n20872_));
  AND2_X2    g18436(.A1(new_n20805_), .A2(new_n12747_), .Z(new_n20873_));
  OAI21_X1   g18437(.A1(new_n20873_), .A2(new_n20872_), .B(new_n12815_), .ZN(new_n20874_));
  INV_X1     g18438(.I(new_n20821_), .ZN(new_n20875_));
  NAND2_X1   g18439(.A1(new_n20805_), .A2(pi0626), .ZN(new_n20876_));
  OAI21_X1   g18440(.A1(pi0626), .A2(new_n20806_), .B(new_n20876_), .ZN(new_n20877_));
  AOI22_X1   g18441(.A1(new_n20877_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n20875_), .ZN(new_n20878_));
  NAND2_X1   g18442(.A1(new_n20878_), .A2(new_n20874_), .ZN(new_n20879_));
  AOI22_X1   g18443(.A1(new_n20871_), .A2(new_n20862_), .B1(pi0788), .B2(new_n20879_), .ZN(new_n20880_));
  OAI22_X1   g18444(.A1(new_n20880_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n20827_), .ZN(new_n20881_));
  NAND2_X1   g18445(.A1(new_n20808_), .A2(new_n13384_), .ZN(new_n20882_));
  NAND2_X1   g18446(.A1(new_n12943_), .A2(new_n20806_), .ZN(new_n20883_));
  NAND2_X1   g18447(.A1(new_n20882_), .A2(new_n20883_), .ZN(new_n20884_));
  NOR2_X1    g18448(.A1(new_n20823_), .A2(new_n12953_), .ZN(new_n20885_));
  NOR2_X1    g18449(.A1(new_n20885_), .A2(pi0647), .ZN(new_n20886_));
  NOR2_X1    g18450(.A1(new_n20787_), .A2(new_n12741_), .ZN(new_n20887_));
  OAI21_X1   g18451(.A1(new_n20886_), .A2(new_n20887_), .B(new_n12965_), .ZN(new_n20888_));
  NAND2_X1   g18452(.A1(new_n20885_), .A2(pi0647), .ZN(new_n20889_));
  OAI21_X1   g18453(.A1(pi0647), .A2(new_n20806_), .B(new_n20889_), .ZN(new_n20890_));
  OAI22_X1   g18454(.A1(new_n20890_), .A2(new_n15576_), .B1(new_n20888_), .B2(new_n12981_), .ZN(new_n20891_));
  AOI21_X1   g18455(.A1(new_n20884_), .A2(new_n15608_), .B(new_n20891_), .ZN(new_n20892_));
  OAI22_X1   g18456(.A1(new_n20881_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n20892_), .ZN(new_n20893_));
  NAND2_X1   g18457(.A1(new_n20893_), .A2(new_n13000_), .ZN(new_n20894_));
  AND2_X2    g18458(.A1(new_n20893_), .A2(new_n12975_), .Z(new_n20895_));
  OAI21_X1   g18459(.A1(new_n20890_), .A2(new_n12965_), .B(new_n20888_), .ZN(new_n20896_));
  NAND2_X1   g18460(.A1(new_n20885_), .A2(new_n12972_), .ZN(new_n20897_));
  OAI21_X1   g18461(.A1(new_n20896_), .A2(new_n12972_), .B(new_n20897_), .ZN(new_n20898_));
  NOR2_X1    g18462(.A1(new_n20898_), .A2(new_n12975_), .ZN(new_n20899_));
  OAI21_X1   g18463(.A1(new_n20895_), .A2(new_n20899_), .B(new_n12740_), .ZN(new_n20900_));
  NAND2_X1   g18464(.A1(new_n20806_), .A2(pi0644), .ZN(new_n20901_));
  NOR2_X1    g18465(.A1(new_n17611_), .A2(new_n20787_), .ZN(new_n20902_));
  AOI21_X1   g18466(.A1(new_n20808_), .A2(new_n17611_), .B(new_n20902_), .ZN(new_n20903_));
  OAI21_X1   g18467(.A1(new_n20903_), .A2(pi0644), .B(new_n20901_), .ZN(new_n20904_));
  NAND2_X1   g18468(.A1(new_n20904_), .A2(pi0715), .ZN(new_n20905_));
  NAND3_X1   g18469(.A1(new_n20900_), .A2(new_n12739_), .A3(new_n20905_), .ZN(new_n20906_));
  NOR2_X1    g18470(.A1(new_n20898_), .A2(pi0644), .ZN(new_n20907_));
  AOI21_X1   g18471(.A1(new_n20893_), .A2(pi0644), .B(new_n20907_), .ZN(new_n20908_));
  NAND2_X1   g18472(.A1(new_n20806_), .A2(new_n12975_), .ZN(new_n20909_));
  OAI21_X1   g18473(.A1(new_n20903_), .A2(new_n12975_), .B(new_n20909_), .ZN(new_n20910_));
  AOI21_X1   g18474(.A1(new_n20910_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n20911_));
  OAI21_X1   g18475(.A1(new_n20908_), .A2(new_n12740_), .B(new_n20911_), .ZN(new_n20912_));
  NAND3_X1   g18476(.A1(new_n20906_), .A2(pi0790), .A3(new_n20912_), .ZN(new_n20913_));
  NAND2_X1   g18477(.A1(new_n20913_), .A2(new_n20894_), .ZN(new_n20914_));
  AOI21_X1   g18478(.A1(po1038), .A2(new_n9517_), .B(pi0832), .ZN(new_n20915_));
  NAND2_X1   g18479(.A1(new_n13192_), .A2(new_n9517_), .ZN(new_n20916_));
  INV_X1     g18480(.I(new_n20916_), .ZN(new_n20917_));
  AOI21_X1   g18481(.A1(new_n20917_), .A2(pi0644), .B(new_n12740_), .ZN(new_n20918_));
  NAND2_X1   g18482(.A1(new_n20916_), .A2(new_n12984_), .ZN(new_n20919_));
  NOR2_X1    g18483(.A1(new_n20917_), .A2(new_n13384_), .ZN(new_n20920_));
  NOR2_X1    g18484(.A1(new_n2609_), .A2(new_n9517_), .ZN(new_n20921_));
  NOR2_X1    g18485(.A1(new_n13342_), .A2(pi0777), .ZN(new_n20922_));
  NOR2_X1    g18486(.A1(new_n13344_), .A2(pi0184), .ZN(new_n20923_));
  NOR3_X1    g18487(.A1(new_n20922_), .A2(new_n3265_), .A3(new_n20923_), .ZN(new_n20924_));
  NAND2_X1   g18488(.A1(new_n13334_), .A2(new_n9517_), .ZN(new_n20925_));
  NAND2_X1   g18489(.A1(new_n13245_), .A2(pi0184), .ZN(new_n20926_));
  AOI21_X1   g18490(.A1(new_n20925_), .A2(new_n20926_), .B(pi0777), .ZN(new_n20927_));
  NOR3_X1    g18491(.A1(new_n15787_), .A2(pi0184), .A3(new_n16757_), .ZN(new_n20928_));
  NOR2_X1    g18492(.A1(new_n20927_), .A2(new_n20928_), .ZN(new_n20929_));
  AOI21_X1   g18493(.A1(new_n20929_), .A2(new_n3265_), .B(new_n20924_), .ZN(new_n20930_));
  NOR2_X1    g18494(.A1(new_n20930_), .A2(new_n2610_), .ZN(new_n20931_));
  NOR2_X1    g18495(.A1(new_n20931_), .A2(new_n20921_), .ZN(new_n20932_));
  NOR2_X1    g18496(.A1(new_n20932_), .A2(new_n12760_), .ZN(new_n20933_));
  INV_X1     g18497(.I(new_n20933_), .ZN(new_n20934_));
  OAI21_X1   g18498(.A1(new_n12761_), .A2(new_n20917_), .B(new_n20934_), .ZN(new_n20935_));
  OAI22_X1   g18499(.A1(new_n20934_), .A2(pi0609), .B1(new_n13353_), .B2(new_n20917_), .ZN(new_n20936_));
  NAND2_X1   g18500(.A1(new_n20936_), .A2(new_n12770_), .ZN(new_n20937_));
  INV_X1     g18501(.I(new_n20937_), .ZN(new_n20938_));
  AOI22_X1   g18502(.A1(new_n20933_), .A2(pi0609), .B1(new_n13357_), .B2(new_n20916_), .ZN(new_n20939_));
  OAI21_X1   g18503(.A1(new_n20939_), .A2(new_n12770_), .B(pi0785), .ZN(new_n20940_));
  OAI22_X1   g18504(.A1(new_n20938_), .A2(new_n20940_), .B1(pi0785), .B2(new_n20935_), .ZN(new_n20941_));
  NAND2_X1   g18505(.A1(new_n20941_), .A2(new_n12779_), .ZN(new_n20942_));
  NAND2_X1   g18506(.A1(new_n20916_), .A2(pi0618), .ZN(new_n20943_));
  OAI21_X1   g18507(.A1(new_n20941_), .A2(pi0618), .B(new_n20943_), .ZN(new_n20944_));
  NAND2_X1   g18508(.A1(new_n20944_), .A2(new_n12785_), .ZN(new_n20945_));
  NAND2_X1   g18509(.A1(new_n20916_), .A2(new_n12781_), .ZN(new_n20946_));
  OAI21_X1   g18510(.A1(new_n20941_), .A2(new_n12781_), .B(new_n20946_), .ZN(new_n20947_));
  NAND2_X1   g18511(.A1(new_n20947_), .A2(pi1154), .ZN(new_n20948_));
  NAND3_X1   g18512(.A1(new_n20945_), .A2(new_n20948_), .A3(pi0781), .ZN(new_n20949_));
  NAND2_X1   g18513(.A1(new_n20949_), .A2(new_n20942_), .ZN(new_n20950_));
  NAND2_X1   g18514(.A1(new_n20950_), .A2(new_n12796_), .ZN(new_n20951_));
  NAND2_X1   g18515(.A1(new_n20916_), .A2(pi0619), .ZN(new_n20952_));
  OAI21_X1   g18516(.A1(new_n20950_), .A2(pi0619), .B(new_n20952_), .ZN(new_n20953_));
  NAND2_X1   g18517(.A1(new_n20953_), .A2(new_n12791_), .ZN(new_n20954_));
  NAND2_X1   g18518(.A1(new_n20916_), .A2(new_n12793_), .ZN(new_n20955_));
  OAI21_X1   g18519(.A1(new_n20950_), .A2(new_n12793_), .B(new_n20955_), .ZN(new_n20956_));
  NAND2_X1   g18520(.A1(new_n20956_), .A2(pi1159), .ZN(new_n20957_));
  NAND3_X1   g18521(.A1(new_n20954_), .A2(new_n20957_), .A3(pi0789), .ZN(new_n20958_));
  NAND2_X1   g18522(.A1(new_n20958_), .A2(new_n20951_), .ZN(new_n20959_));
  NAND2_X1   g18523(.A1(new_n20916_), .A2(new_n12818_), .ZN(new_n20960_));
  OAI21_X1   g18524(.A1(new_n20959_), .A2(new_n12818_), .B(new_n20960_), .ZN(new_n20961_));
  AOI21_X1   g18525(.A1(new_n20961_), .A2(new_n13384_), .B(new_n20920_), .ZN(new_n20962_));
  OAI21_X1   g18526(.A1(new_n20962_), .A2(new_n12984_), .B(new_n20919_), .ZN(new_n20963_));
  OAI21_X1   g18527(.A1(new_n20963_), .A2(pi0644), .B(new_n20918_), .ZN(new_n20964_));
  AND2_X2    g18528(.A1(new_n20964_), .A2(new_n12739_), .Z(new_n20965_));
  OAI21_X1   g18529(.A1(new_n14125_), .A2(new_n20923_), .B(new_n16756_), .ZN(new_n20966_));
  OAI21_X1   g18530(.A1(new_n14122_), .A2(new_n9517_), .B(new_n3265_), .ZN(new_n20967_));
  NAND2_X1   g18531(.A1(new_n20967_), .A2(new_n2609_), .ZN(new_n20968_));
  NAND2_X1   g18532(.A1(new_n15744_), .A2(new_n9517_), .ZN(new_n20969_));
  AOI21_X1   g18533(.A1(new_n20969_), .A2(new_n20968_), .B(new_n20966_), .ZN(new_n20970_));
  NAND2_X1   g18534(.A1(new_n2609_), .A2(new_n16756_), .ZN(new_n20971_));
  AOI21_X1   g18535(.A1(new_n20917_), .A2(new_n20971_), .B(new_n20970_), .ZN(new_n20972_));
  NAND2_X1   g18536(.A1(new_n20972_), .A2(new_n13521_), .ZN(new_n20973_));
  NAND2_X1   g18537(.A1(new_n20916_), .A2(pi0625), .ZN(new_n20974_));
  AOI21_X1   g18538(.A1(new_n20973_), .A2(new_n20974_), .B(pi1153), .ZN(new_n20975_));
  NAND2_X1   g18539(.A1(new_n20916_), .A2(new_n13521_), .ZN(new_n20976_));
  NAND2_X1   g18540(.A1(new_n20972_), .A2(pi0625), .ZN(new_n20977_));
  AOI21_X1   g18541(.A1(new_n20977_), .A2(new_n20976_), .B(new_n12841_), .ZN(new_n20978_));
  NOR3_X1    g18542(.A1(new_n20975_), .A2(new_n20978_), .A3(new_n12758_), .ZN(new_n20979_));
  NOR2_X1    g18543(.A1(new_n20972_), .A2(pi0778), .ZN(new_n20980_));
  NOR2_X1    g18544(.A1(new_n20979_), .A2(new_n20980_), .ZN(new_n20981_));
  NOR2_X1    g18545(.A1(new_n20981_), .A2(new_n12869_), .ZN(new_n20982_));
  AOI21_X1   g18546(.A1(new_n12869_), .A2(new_n20917_), .B(new_n20982_), .ZN(new_n20983_));
  NAND2_X1   g18547(.A1(new_n20983_), .A2(new_n12888_), .ZN(new_n20984_));
  OAI21_X1   g18548(.A1(new_n12888_), .A2(new_n20917_), .B(new_n20984_), .ZN(new_n20985_));
  INV_X1     g18549(.I(new_n20985_), .ZN(new_n20986_));
  NOR2_X1    g18550(.A1(new_n20916_), .A2(new_n12911_), .ZN(new_n20987_));
  AOI21_X1   g18551(.A1(new_n20986_), .A2(new_n12911_), .B(new_n20987_), .ZN(new_n20988_));
  NAND2_X1   g18552(.A1(new_n20988_), .A2(new_n13392_), .ZN(new_n20989_));
  OAI21_X1   g18553(.A1(new_n13392_), .A2(new_n20917_), .B(new_n20989_), .ZN(new_n20990_));
  NAND2_X1   g18554(.A1(new_n20990_), .A2(new_n12920_), .ZN(new_n20991_));
  NAND2_X1   g18555(.A1(new_n20916_), .A2(pi0628), .ZN(new_n20992_));
  AOI21_X1   g18556(.A1(new_n20991_), .A2(new_n20992_), .B(pi1156), .ZN(new_n20993_));
  NAND2_X1   g18557(.A1(new_n20916_), .A2(new_n12920_), .ZN(new_n20994_));
  NAND2_X1   g18558(.A1(new_n20990_), .A2(pi0628), .ZN(new_n20995_));
  AOI21_X1   g18559(.A1(new_n20995_), .A2(new_n20994_), .B(new_n12742_), .ZN(new_n20996_));
  OR2_X2     g18560(.A1(new_n20996_), .A2(new_n12937_), .Z(new_n20997_));
  OAI22_X1   g18561(.A1(new_n20997_), .A2(new_n20993_), .B1(pi0792), .B2(new_n20990_), .ZN(new_n20998_));
  NAND2_X1   g18562(.A1(new_n20998_), .A2(new_n12741_), .ZN(new_n20999_));
  OAI21_X1   g18563(.A1(new_n12741_), .A2(new_n20916_), .B(new_n20999_), .ZN(new_n21000_));
  NOR2_X1    g18564(.A1(new_n21000_), .A2(pi1157), .ZN(new_n21001_));
  NAND2_X1   g18565(.A1(new_n20998_), .A2(pi0647), .ZN(new_n21002_));
  OAI21_X1   g18566(.A1(pi0647), .A2(new_n20916_), .B(new_n21002_), .ZN(new_n21003_));
  NOR2_X1    g18567(.A1(new_n21003_), .A2(new_n12965_), .ZN(new_n21004_));
  OAI21_X1   g18568(.A1(new_n21001_), .A2(new_n21004_), .B(pi0787), .ZN(new_n21005_));
  OAI21_X1   g18569(.A1(pi0787), .A2(new_n20998_), .B(new_n21005_), .ZN(new_n21006_));
  OAI21_X1   g18570(.A1(new_n21006_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n21007_));
  AOI21_X1   g18571(.A1(new_n20917_), .A2(new_n12975_), .B(pi0715), .ZN(new_n21008_));
  OAI21_X1   g18572(.A1(new_n20963_), .A2(new_n12975_), .B(new_n21008_), .ZN(new_n21009_));
  AND2_X2    g18573(.A1(new_n21009_), .A2(pi1160), .Z(new_n21010_));
  OAI21_X1   g18574(.A1(new_n21006_), .A2(pi0644), .B(pi0715), .ZN(new_n21011_));
  AOI22_X1   g18575(.A1(new_n20965_), .A2(new_n21007_), .B1(new_n21011_), .B2(new_n21010_), .ZN(new_n21012_));
  NOR2_X1    g18576(.A1(new_n21012_), .A2(new_n13000_), .ZN(new_n21013_));
  NAND2_X1   g18577(.A1(new_n20917_), .A2(pi0626), .ZN(new_n21014_));
  NAND2_X1   g18578(.A1(new_n20959_), .A2(new_n12747_), .ZN(new_n21015_));
  AOI21_X1   g18579(.A1(new_n21015_), .A2(new_n21014_), .B(new_n12816_), .ZN(new_n21016_));
  NOR2_X1    g18580(.A1(new_n20916_), .A2(pi0626), .ZN(new_n21017_));
  AOI21_X1   g18581(.A1(new_n20959_), .A2(pi0626), .B(new_n21017_), .ZN(new_n21018_));
  OAI22_X1   g18582(.A1(new_n21018_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n20988_), .ZN(new_n21019_));
  OAI21_X1   g18583(.A1(new_n21019_), .A2(new_n21016_), .B(pi0788), .ZN(new_n21020_));
  NAND2_X1   g18584(.A1(new_n21020_), .A2(new_n15824_), .ZN(new_n21021_));
  NAND2_X1   g18585(.A1(new_n20981_), .A2(new_n12766_), .ZN(new_n21022_));
  AOI21_X1   g18586(.A1(new_n16757_), .A2(new_n13566_), .B(new_n15826_), .ZN(new_n21023_));
  AOI21_X1   g18587(.A1(new_n14328_), .A2(new_n20790_), .B(new_n9517_), .ZN(new_n21024_));
  AOI21_X1   g18588(.A1(new_n21024_), .A2(new_n5336_), .B(new_n3265_), .ZN(new_n21025_));
  OAI21_X1   g18589(.A1(new_n21023_), .A2(pi0184), .B(new_n21025_), .ZN(new_n21026_));
  NAND2_X1   g18590(.A1(new_n14172_), .A2(pi0184), .ZN(new_n21027_));
  NAND2_X1   g18591(.A1(new_n14174_), .A2(new_n9517_), .ZN(new_n21028_));
  AOI21_X1   g18592(.A1(new_n21027_), .A2(new_n21028_), .B(pi0777), .ZN(new_n21029_));
  NAND2_X1   g18593(.A1(new_n15835_), .A2(pi0184), .ZN(new_n21030_));
  NAND2_X1   g18594(.A1(new_n14177_), .A2(new_n9517_), .ZN(new_n21031_));
  AOI21_X1   g18595(.A1(new_n21031_), .A2(new_n21030_), .B(new_n16757_), .ZN(new_n21032_));
  OAI21_X1   g18596(.A1(new_n21032_), .A2(new_n21029_), .B(new_n2627_), .ZN(new_n21033_));
  NOR2_X1    g18597(.A1(new_n14182_), .A2(pi0184), .ZN(new_n21034_));
  NOR2_X1    g18598(.A1(new_n14184_), .A2(new_n9517_), .ZN(new_n21035_));
  OAI21_X1   g18599(.A1(new_n21034_), .A2(new_n21035_), .B(pi0777), .ZN(new_n21036_));
  NOR2_X1    g18600(.A1(new_n14187_), .A2(new_n9517_), .ZN(new_n21037_));
  NOR2_X1    g18601(.A1(new_n14189_), .A2(pi0184), .ZN(new_n21038_));
  OAI21_X1   g18602(.A1(new_n21037_), .A2(new_n21038_), .B(new_n16757_), .ZN(new_n21039_));
  NAND3_X1   g18603(.A1(new_n21039_), .A2(new_n21036_), .A3(pi0039), .ZN(new_n21040_));
  NAND3_X1   g18604(.A1(new_n21040_), .A2(new_n3265_), .A3(new_n21033_), .ZN(new_n21041_));
  NAND3_X1   g18605(.A1(new_n21041_), .A2(new_n16756_), .A3(new_n21026_), .ZN(new_n21042_));
  NAND2_X1   g18606(.A1(new_n20930_), .A2(pi0737), .ZN(new_n21043_));
  NAND3_X1   g18607(.A1(new_n21042_), .A2(new_n2609_), .A3(new_n21043_), .ZN(new_n21044_));
  OAI21_X1   g18608(.A1(new_n9517_), .A2(new_n2609_), .B(new_n21044_), .ZN(new_n21045_));
  INV_X1     g18609(.I(new_n20978_), .ZN(new_n21046_));
  NOR2_X1    g18610(.A1(new_n20932_), .A2(new_n13521_), .ZN(new_n21047_));
  AOI21_X1   g18611(.A1(new_n21045_), .A2(new_n13521_), .B(new_n21047_), .ZN(new_n21048_));
  OAI21_X1   g18612(.A1(new_n21048_), .A2(pi1153), .B(new_n21046_), .ZN(new_n21049_));
  NOR2_X1    g18613(.A1(new_n20932_), .A2(pi0625), .ZN(new_n21050_));
  AOI21_X1   g18614(.A1(new_n21045_), .A2(pi0625), .B(new_n21050_), .ZN(new_n21051_));
  OAI21_X1   g18615(.A1(new_n21051_), .A2(new_n12841_), .B(pi0608), .ZN(new_n21052_));
  OAI22_X1   g18616(.A1(pi0608), .A2(new_n21049_), .B1(new_n21052_), .B2(new_n20975_), .ZN(new_n21053_));
  NOR2_X1    g18617(.A1(new_n21053_), .A2(new_n12758_), .ZN(new_n21054_));
  AOI21_X1   g18618(.A1(new_n12758_), .A2(new_n21045_), .B(new_n21054_), .ZN(new_n21055_));
  OAI21_X1   g18619(.A1(new_n21055_), .A2(new_n12766_), .B(new_n21022_), .ZN(new_n21056_));
  AOI21_X1   g18620(.A1(new_n21056_), .A2(pi1155), .B(new_n20938_), .ZN(new_n21057_));
  NOR2_X1    g18621(.A1(new_n21055_), .A2(pi0609), .ZN(new_n21058_));
  NOR3_X1    g18622(.A1(new_n20979_), .A2(new_n12766_), .A3(new_n20980_), .ZN(new_n21059_));
  OAI21_X1   g18623(.A1(new_n21058_), .A2(new_n21059_), .B(new_n12770_), .ZN(new_n21060_));
  NOR2_X1    g18624(.A1(new_n20939_), .A2(new_n12770_), .ZN(new_n21061_));
  NOR2_X1    g18625(.A1(new_n21061_), .A2(pi0660), .ZN(new_n21062_));
  AOI22_X1   g18626(.A1(new_n21057_), .A2(pi0660), .B1(new_n21060_), .B2(new_n21062_), .ZN(new_n21063_));
  NOR2_X1    g18627(.A1(new_n21055_), .A2(pi0785), .ZN(new_n21064_));
  AOI21_X1   g18628(.A1(new_n21063_), .A2(pi0785), .B(new_n21064_), .ZN(new_n21065_));
  NOR2_X1    g18629(.A1(new_n21065_), .A2(pi0781), .ZN(new_n21066_));
  AND2_X2    g18630(.A1(new_n20983_), .A2(new_n12781_), .Z(new_n21067_));
  NOR2_X1    g18631(.A1(new_n21065_), .A2(new_n12781_), .ZN(new_n21068_));
  OAI21_X1   g18632(.A1(new_n21068_), .A2(new_n21067_), .B(pi1154), .ZN(new_n21069_));
  NAND3_X1   g18633(.A1(new_n21069_), .A2(pi0627), .A3(new_n20945_), .ZN(new_n21070_));
  INV_X1     g18634(.I(new_n20948_), .ZN(new_n21071_));
  NAND2_X1   g18635(.A1(new_n20983_), .A2(pi0618), .ZN(new_n21072_));
  OAI21_X1   g18636(.A1(new_n21065_), .A2(pi0618), .B(new_n21072_), .ZN(new_n21073_));
  AOI21_X1   g18637(.A1(new_n21073_), .A2(new_n12785_), .B(new_n21071_), .ZN(new_n21074_));
  AOI21_X1   g18638(.A1(new_n21074_), .A2(new_n12880_), .B(new_n12779_), .ZN(new_n21075_));
  AOI21_X1   g18639(.A1(new_n21075_), .A2(new_n21070_), .B(new_n21066_), .ZN(new_n21076_));
  OAI21_X1   g18640(.A1(new_n21076_), .A2(pi0789), .B(new_n12819_), .ZN(new_n21077_));
  NOR2_X1    g18641(.A1(new_n20986_), .A2(new_n12793_), .ZN(new_n21078_));
  NOR2_X1    g18642(.A1(new_n21076_), .A2(pi0619), .ZN(new_n21079_));
  OAI21_X1   g18643(.A1(new_n21079_), .A2(new_n21078_), .B(new_n12791_), .ZN(new_n21080_));
  NAND3_X1   g18644(.A1(new_n21080_), .A2(new_n12895_), .A3(new_n20957_), .ZN(new_n21081_));
  NAND2_X1   g18645(.A1(new_n20985_), .A2(new_n12793_), .ZN(new_n21082_));
  OAI21_X1   g18646(.A1(new_n21076_), .A2(new_n12793_), .B(new_n21082_), .ZN(new_n21083_));
  AOI21_X1   g18647(.A1(new_n21083_), .A2(pi1159), .B(new_n12895_), .ZN(new_n21084_));
  AOI21_X1   g18648(.A1(new_n21084_), .A2(new_n20954_), .B(new_n12796_), .ZN(new_n21085_));
  AOI21_X1   g18649(.A1(new_n21085_), .A2(new_n21081_), .B(new_n21077_), .ZN(new_n21086_));
  NOR2_X1    g18650(.A1(new_n20996_), .A2(pi0629), .ZN(new_n21087_));
  NOR2_X1    g18651(.A1(new_n20993_), .A2(new_n12919_), .ZN(new_n21088_));
  NOR2_X1    g18652(.A1(new_n21087_), .A2(new_n21088_), .ZN(new_n21089_));
  AOI21_X1   g18653(.A1(new_n20961_), .A2(new_n19160_), .B(new_n21089_), .ZN(new_n21090_));
  OAI22_X1   g18654(.A1(new_n21086_), .A2(new_n21021_), .B1(new_n12937_), .B2(new_n21090_), .ZN(new_n21091_));
  NOR2_X1    g18655(.A1(new_n21010_), .A2(new_n12975_), .ZN(new_n21092_));
  NOR2_X1    g18656(.A1(new_n20965_), .A2(pi0644), .ZN(new_n21093_));
  NOR2_X1    g18657(.A1(new_n21092_), .A2(new_n21093_), .ZN(new_n21094_));
  OAI22_X1   g18658(.A1(new_n15576_), .A2(new_n21003_), .B1(new_n21000_), .B2(new_n15730_), .ZN(new_n21095_));
  NOR2_X1    g18659(.A1(new_n20962_), .A2(new_n17212_), .ZN(new_n21096_));
  NOR2_X1    g18660(.A1(new_n21095_), .A2(new_n21096_), .ZN(new_n21097_));
  OAI22_X1   g18661(.A1(new_n21094_), .A2(new_n13000_), .B1(new_n21097_), .B2(new_n12972_), .ZN(new_n21098_));
  AOI21_X1   g18662(.A1(new_n15693_), .A2(new_n21091_), .B(new_n21098_), .ZN(new_n21099_));
  OAI21_X1   g18663(.A1(new_n21013_), .A2(new_n21099_), .B(new_n6643_), .ZN(new_n21100_));
  AOI22_X1   g18664(.A1(new_n21100_), .A2(new_n20915_), .B1(pi0832), .B2(new_n20914_), .ZN(po0341));
  NOR2_X1    g18665(.A1(new_n13340_), .A2(pi0751), .ZN(new_n21102_));
  NOR2_X1    g18666(.A1(new_n3042_), .A2(pi0185), .ZN(new_n21103_));
  NOR2_X1    g18667(.A1(new_n21102_), .A2(new_n21103_), .ZN(new_n21104_));
  NOR3_X1    g18668(.A1(new_n21104_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n21105_));
  INV_X1     g18669(.I(new_n21102_), .ZN(new_n21106_));
  NOR2_X1    g18670(.A1(new_n21106_), .A2(new_n13354_), .ZN(new_n21107_));
  NOR3_X1    g18671(.A1(new_n21107_), .A2(new_n12762_), .A3(new_n21104_), .ZN(new_n21108_));
  NOR2_X1    g18672(.A1(new_n21108_), .A2(new_n12770_), .ZN(new_n21109_));
  NOR3_X1    g18673(.A1(new_n21107_), .A2(pi1155), .A3(new_n21103_), .ZN(new_n21110_));
  NOR3_X1    g18674(.A1(new_n21109_), .A2(new_n12764_), .A3(new_n21110_), .ZN(new_n21111_));
  NOR2_X1    g18675(.A1(new_n21111_), .A2(new_n21105_), .ZN(new_n21112_));
  INV_X1     g18676(.I(new_n21112_), .ZN(new_n21113_));
  AOI21_X1   g18677(.A1(new_n21113_), .A2(new_n12783_), .B(pi1154), .ZN(new_n21114_));
  AOI21_X1   g18678(.A1(new_n21113_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n21115_));
  NOR3_X1    g18679(.A1(new_n21114_), .A2(new_n21115_), .A3(new_n12779_), .ZN(new_n21116_));
  AOI21_X1   g18680(.A1(new_n12779_), .A2(new_n21113_), .B(new_n21116_), .ZN(new_n21117_));
  OAI21_X1   g18681(.A1(new_n21117_), .A2(new_n17229_), .B(new_n12791_), .ZN(new_n21118_));
  OAI21_X1   g18682(.A1(new_n21117_), .A2(new_n17232_), .B(pi1159), .ZN(new_n21119_));
  NAND3_X1   g18683(.A1(new_n21118_), .A2(new_n21119_), .A3(pi0789), .ZN(new_n21120_));
  OAI21_X1   g18684(.A1(pi0789), .A2(new_n21117_), .B(new_n21120_), .ZN(new_n21121_));
  INV_X1     g18685(.I(new_n21103_), .ZN(new_n21122_));
  NAND2_X1   g18686(.A1(new_n12818_), .A2(new_n21122_), .ZN(new_n21123_));
  OAI21_X1   g18687(.A1(new_n21121_), .A2(new_n12818_), .B(new_n21123_), .ZN(new_n21124_));
  AOI21_X1   g18688(.A1(new_n12826_), .A2(new_n16218_), .B(new_n21103_), .ZN(new_n21125_));
  NOR2_X1    g18689(.A1(new_n21103_), .A2(pi1153), .ZN(new_n21126_));
  NOR2_X1    g18690(.A1(new_n12834_), .A2(pi0701), .ZN(new_n21127_));
  INV_X1     g18691(.I(new_n21127_), .ZN(new_n21128_));
  NAND2_X1   g18692(.A1(new_n21128_), .A2(new_n21126_), .ZN(new_n21129_));
  NOR2_X1    g18693(.A1(new_n21127_), .A2(new_n21125_), .ZN(new_n21130_));
  NOR2_X1    g18694(.A1(new_n21130_), .A2(new_n12841_), .ZN(new_n21131_));
  INV_X1     g18695(.I(new_n21131_), .ZN(new_n21132_));
  NAND3_X1   g18696(.A1(new_n21132_), .A2(pi0778), .A3(new_n21129_), .ZN(new_n21133_));
  OAI21_X1   g18697(.A1(pi0778), .A2(new_n21125_), .B(new_n21133_), .ZN(new_n21134_));
  NAND2_X1   g18698(.A1(new_n21134_), .A2(new_n17187_), .ZN(new_n21135_));
  NOR2_X1    g18699(.A1(new_n21135_), .A2(new_n12889_), .ZN(new_n21136_));
  NAND2_X1   g18700(.A1(new_n21136_), .A2(new_n18203_), .ZN(new_n21137_));
  NOR2_X1    g18701(.A1(new_n21137_), .A2(new_n17884_), .ZN(new_n21138_));
  INV_X1     g18702(.I(new_n21138_), .ZN(new_n21139_));
  OAI22_X1   g18703(.A1(new_n21124_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n21139_), .ZN(new_n21140_));
  AND2_X2    g18704(.A1(new_n21140_), .A2(new_n12919_), .Z(new_n21141_));
  OAI22_X1   g18705(.A1(new_n21124_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n21139_), .ZN(new_n21142_));
  AOI21_X1   g18706(.A1(pi0629), .A2(new_n21142_), .B(new_n21141_), .ZN(new_n21143_));
  INV_X1     g18707(.I(new_n21110_), .ZN(new_n21144_));
  NOR2_X1    g18708(.A1(new_n21125_), .A2(new_n12754_), .ZN(new_n21145_));
  NOR3_X1    g18709(.A1(new_n21145_), .A2(new_n21102_), .A3(new_n21103_), .ZN(new_n21146_));
  NAND2_X1   g18710(.A1(new_n21146_), .A2(new_n12758_), .ZN(new_n21147_));
  NAND2_X1   g18711(.A1(new_n21145_), .A2(pi0625), .ZN(new_n21148_));
  NAND3_X1   g18712(.A1(new_n21148_), .A2(pi1153), .A3(new_n21104_), .ZN(new_n21149_));
  NAND3_X1   g18713(.A1(new_n21129_), .A2(pi0608), .A3(new_n21149_), .ZN(new_n21150_));
  INV_X1     g18714(.I(new_n21148_), .ZN(new_n21151_));
  OAI21_X1   g18715(.A1(new_n21151_), .A2(new_n21146_), .B(new_n21126_), .ZN(new_n21152_));
  NAND3_X1   g18716(.A1(new_n21132_), .A2(new_n13560_), .A3(new_n21152_), .ZN(new_n21153_));
  NAND3_X1   g18717(.A1(new_n21153_), .A2(pi0778), .A3(new_n21150_), .ZN(new_n21154_));
  AOI21_X1   g18718(.A1(new_n21154_), .A2(new_n21147_), .B(new_n12766_), .ZN(new_n21155_));
  NOR2_X1    g18719(.A1(new_n21134_), .A2(pi0609), .ZN(new_n21156_));
  OAI21_X1   g18720(.A1(new_n21156_), .A2(new_n21155_), .B(pi1155), .ZN(new_n21157_));
  NAND3_X1   g18721(.A1(new_n21157_), .A2(pi0660), .A3(new_n21144_), .ZN(new_n21158_));
  NAND2_X1   g18722(.A1(new_n21154_), .A2(new_n21147_), .ZN(new_n21159_));
  NOR2_X1    g18723(.A1(new_n21134_), .A2(new_n12766_), .ZN(new_n21160_));
  AOI21_X1   g18724(.A1(new_n21159_), .A2(new_n12766_), .B(new_n21160_), .ZN(new_n21161_));
  NOR2_X1    g18725(.A1(new_n21109_), .A2(pi0660), .ZN(new_n21162_));
  OAI21_X1   g18726(.A1(new_n21161_), .A2(pi1155), .B(new_n21162_), .ZN(new_n21163_));
  NAND3_X1   g18727(.A1(new_n21163_), .A2(new_n21158_), .A3(pi0785), .ZN(new_n21164_));
  NAND2_X1   g18728(.A1(new_n21159_), .A2(new_n12764_), .ZN(new_n21165_));
  NAND2_X1   g18729(.A1(new_n21164_), .A2(new_n21165_), .ZN(new_n21166_));
  NAND2_X1   g18730(.A1(new_n21166_), .A2(new_n12781_), .ZN(new_n21167_));
  NAND2_X1   g18731(.A1(new_n21135_), .A2(pi0618), .ZN(new_n21168_));
  AOI21_X1   g18732(.A1(new_n21167_), .A2(new_n21168_), .B(pi1154), .ZN(new_n21169_));
  NOR3_X1    g18733(.A1(new_n21169_), .A2(pi0627), .A3(new_n21115_), .ZN(new_n21170_));
  NAND2_X1   g18734(.A1(new_n21135_), .A2(new_n12781_), .ZN(new_n21171_));
  NAND2_X1   g18735(.A1(new_n21166_), .A2(pi0618), .ZN(new_n21172_));
  AOI21_X1   g18736(.A1(new_n21172_), .A2(new_n21171_), .B(new_n12785_), .ZN(new_n21173_));
  NOR3_X1    g18737(.A1(new_n21173_), .A2(new_n12880_), .A3(new_n21114_), .ZN(new_n21174_));
  OR3_X2     g18738(.A1(new_n21170_), .A2(new_n21174_), .A3(new_n12779_), .Z(new_n21175_));
  NAND2_X1   g18739(.A1(new_n21166_), .A2(new_n12779_), .ZN(new_n21176_));
  NAND2_X1   g18740(.A1(new_n21175_), .A2(new_n21176_), .ZN(new_n21177_));
  AOI21_X1   g18741(.A1(new_n21177_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n21178_));
  NOR2_X1    g18742(.A1(new_n21136_), .A2(pi0619), .ZN(new_n21179_));
  AOI21_X1   g18743(.A1(new_n21175_), .A2(new_n21176_), .B(new_n12793_), .ZN(new_n21180_));
  OAI21_X1   g18744(.A1(new_n21180_), .A2(new_n21179_), .B(pi1159), .ZN(new_n21181_));
  NAND3_X1   g18745(.A1(new_n21181_), .A2(pi0648), .A3(new_n21118_), .ZN(new_n21182_));
  NAND2_X1   g18746(.A1(new_n21177_), .A2(new_n12793_), .ZN(new_n21183_));
  OAI21_X1   g18747(.A1(new_n12793_), .A2(new_n21136_), .B(new_n21183_), .ZN(new_n21184_));
  NAND2_X1   g18748(.A1(new_n21184_), .A2(new_n12791_), .ZN(new_n21185_));
  NAND3_X1   g18749(.A1(new_n21185_), .A2(new_n12895_), .A3(new_n21119_), .ZN(new_n21186_));
  NAND3_X1   g18750(.A1(new_n21186_), .A2(pi0789), .A3(new_n21182_), .ZN(new_n21187_));
  NOR2_X1    g18751(.A1(new_n21122_), .A2(new_n12747_), .ZN(new_n21188_));
  AND2_X2    g18752(.A1(new_n21121_), .A2(new_n12747_), .Z(new_n21189_));
  OAI21_X1   g18753(.A1(new_n21189_), .A2(new_n21188_), .B(new_n12815_), .ZN(new_n21190_));
  INV_X1     g18754(.I(new_n21137_), .ZN(new_n21191_));
  NAND2_X1   g18755(.A1(new_n21121_), .A2(pi0626), .ZN(new_n21192_));
  OAI21_X1   g18756(.A1(pi0626), .A2(new_n21122_), .B(new_n21192_), .ZN(new_n21193_));
  AOI22_X1   g18757(.A1(new_n21193_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n21191_), .ZN(new_n21194_));
  NAND2_X1   g18758(.A1(new_n21194_), .A2(new_n21190_), .ZN(new_n21195_));
  AOI22_X1   g18759(.A1(new_n21187_), .A2(new_n21178_), .B1(pi0788), .B2(new_n21195_), .ZN(new_n21196_));
  OAI22_X1   g18760(.A1(new_n21196_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n21143_), .ZN(new_n21197_));
  NAND2_X1   g18761(.A1(new_n21124_), .A2(new_n13384_), .ZN(new_n21198_));
  NAND2_X1   g18762(.A1(new_n12943_), .A2(new_n21122_), .ZN(new_n21199_));
  NAND2_X1   g18763(.A1(new_n21198_), .A2(new_n21199_), .ZN(new_n21200_));
  NOR2_X1    g18764(.A1(new_n21139_), .A2(new_n12953_), .ZN(new_n21201_));
  NOR2_X1    g18765(.A1(new_n21201_), .A2(pi0647), .ZN(new_n21202_));
  NOR2_X1    g18766(.A1(new_n21103_), .A2(new_n12741_), .ZN(new_n21203_));
  OAI21_X1   g18767(.A1(new_n21202_), .A2(new_n21203_), .B(new_n12965_), .ZN(new_n21204_));
  NAND2_X1   g18768(.A1(new_n21201_), .A2(pi0647), .ZN(new_n21205_));
  OAI21_X1   g18769(.A1(pi0647), .A2(new_n21122_), .B(new_n21205_), .ZN(new_n21206_));
  OAI22_X1   g18770(.A1(new_n21206_), .A2(new_n15576_), .B1(new_n21204_), .B2(new_n12981_), .ZN(new_n21207_));
  AOI21_X1   g18771(.A1(new_n21200_), .A2(new_n15608_), .B(new_n21207_), .ZN(new_n21208_));
  OAI22_X1   g18772(.A1(new_n21197_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n21208_), .ZN(new_n21209_));
  NAND2_X1   g18773(.A1(new_n21209_), .A2(new_n13000_), .ZN(new_n21210_));
  AND2_X2    g18774(.A1(new_n21209_), .A2(new_n12975_), .Z(new_n21211_));
  OAI21_X1   g18775(.A1(new_n21206_), .A2(new_n12965_), .B(new_n21204_), .ZN(new_n21212_));
  NAND2_X1   g18776(.A1(new_n21201_), .A2(new_n12972_), .ZN(new_n21213_));
  OAI21_X1   g18777(.A1(new_n21212_), .A2(new_n12972_), .B(new_n21213_), .ZN(new_n21214_));
  NOR2_X1    g18778(.A1(new_n21214_), .A2(new_n12975_), .ZN(new_n21215_));
  OAI21_X1   g18779(.A1(new_n21211_), .A2(new_n21215_), .B(new_n12740_), .ZN(new_n21216_));
  NAND2_X1   g18780(.A1(new_n21122_), .A2(pi0644), .ZN(new_n21217_));
  NOR2_X1    g18781(.A1(new_n17611_), .A2(new_n21103_), .ZN(new_n21218_));
  AOI21_X1   g18782(.A1(new_n21124_), .A2(new_n17611_), .B(new_n21218_), .ZN(new_n21219_));
  OAI21_X1   g18783(.A1(new_n21219_), .A2(pi0644), .B(new_n21217_), .ZN(new_n21220_));
  NAND2_X1   g18784(.A1(new_n21220_), .A2(pi0715), .ZN(new_n21221_));
  NAND3_X1   g18785(.A1(new_n21216_), .A2(new_n12739_), .A3(new_n21221_), .ZN(new_n21222_));
  NOR2_X1    g18786(.A1(new_n21214_), .A2(pi0644), .ZN(new_n21223_));
  AOI21_X1   g18787(.A1(new_n21209_), .A2(pi0644), .B(new_n21223_), .ZN(new_n21224_));
  NAND2_X1   g18788(.A1(new_n21122_), .A2(new_n12975_), .ZN(new_n21225_));
  OAI21_X1   g18789(.A1(new_n21219_), .A2(new_n12975_), .B(new_n21225_), .ZN(new_n21226_));
  AOI21_X1   g18790(.A1(new_n21226_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n21227_));
  OAI21_X1   g18791(.A1(new_n21224_), .A2(new_n12740_), .B(new_n21227_), .ZN(new_n21228_));
  NAND3_X1   g18792(.A1(new_n21222_), .A2(pi0790), .A3(new_n21228_), .ZN(new_n21229_));
  NAND2_X1   g18793(.A1(new_n21229_), .A2(new_n21210_), .ZN(new_n21230_));
  AOI21_X1   g18794(.A1(po1038), .A2(new_n10688_), .B(pi0832), .ZN(new_n21231_));
  NAND2_X1   g18795(.A1(new_n13192_), .A2(new_n10688_), .ZN(new_n21232_));
  INV_X1     g18796(.I(new_n21232_), .ZN(new_n21233_));
  AOI21_X1   g18797(.A1(new_n21233_), .A2(pi0644), .B(new_n12740_), .ZN(new_n21234_));
  NAND2_X1   g18798(.A1(new_n21232_), .A2(new_n12984_), .ZN(new_n21235_));
  NOR2_X1    g18799(.A1(new_n21233_), .A2(new_n13384_), .ZN(new_n21236_));
  NAND2_X1   g18800(.A1(new_n2610_), .A2(pi0185), .ZN(new_n21237_));
  OAI22_X1   g18801(.A1(new_n19651_), .A2(new_n10688_), .B1(new_n16210_), .B2(new_n13060_), .ZN(new_n21238_));
  NAND2_X1   g18802(.A1(new_n10688_), .A2(pi0751), .ZN(new_n21239_));
  OAI21_X1   g18803(.A1(new_n13334_), .A2(pi0185), .B(new_n16210_), .ZN(new_n21240_));
  AOI22_X1   g18804(.A1(new_n21240_), .A2(new_n21239_), .B1(new_n2627_), .B2(new_n21238_), .ZN(new_n21241_));
  OAI22_X1   g18805(.A1(new_n14065_), .A2(new_n16210_), .B1(new_n10688_), .B2(new_n14067_), .ZN(new_n21242_));
  NAND2_X1   g18806(.A1(new_n21242_), .A2(pi0039), .ZN(new_n21243_));
  NAND2_X1   g18807(.A1(new_n21241_), .A2(new_n21243_), .ZN(new_n21244_));
  NOR2_X1    g18808(.A1(new_n13344_), .A2(pi0185), .ZN(new_n21245_));
  NOR2_X1    g18809(.A1(new_n21245_), .A2(new_n3265_), .ZN(new_n21246_));
  NAND2_X1   g18810(.A1(new_n13341_), .A2(new_n16210_), .ZN(new_n21247_));
  AOI22_X1   g18811(.A1(new_n21244_), .A2(new_n3265_), .B1(new_n21246_), .B2(new_n21247_), .ZN(new_n21248_));
  OAI21_X1   g18812(.A1(new_n21248_), .A2(new_n2610_), .B(new_n21237_), .ZN(new_n21249_));
  NAND2_X1   g18813(.A1(new_n21249_), .A2(new_n12761_), .ZN(new_n21250_));
  INV_X1     g18814(.I(new_n21250_), .ZN(new_n21251_));
  NOR2_X1    g18815(.A1(new_n21233_), .A2(new_n12761_), .ZN(new_n21252_));
  NOR3_X1    g18816(.A1(new_n21251_), .A2(pi0785), .A3(new_n21252_), .ZN(new_n21253_));
  AOI22_X1   g18817(.A1(new_n21251_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n21232_), .ZN(new_n21254_));
  NOR2_X1    g18818(.A1(new_n21254_), .A2(pi1155), .ZN(new_n21255_));
  AOI22_X1   g18819(.A1(new_n21251_), .A2(pi0609), .B1(new_n13357_), .B2(new_n21232_), .ZN(new_n21256_));
  NOR2_X1    g18820(.A1(new_n21256_), .A2(new_n12770_), .ZN(new_n21257_));
  NOR3_X1    g18821(.A1(new_n21257_), .A2(new_n21255_), .A3(new_n12764_), .ZN(new_n21258_));
  NOR2_X1    g18822(.A1(new_n21258_), .A2(new_n21253_), .ZN(new_n21259_));
  NOR2_X1    g18823(.A1(new_n21259_), .A2(pi0781), .ZN(new_n21260_));
  NOR3_X1    g18824(.A1(new_n21258_), .A2(pi0618), .A3(new_n21253_), .ZN(new_n21261_));
  NOR2_X1    g18825(.A1(new_n21233_), .A2(new_n12781_), .ZN(new_n21262_));
  OAI21_X1   g18826(.A1(new_n21261_), .A2(new_n21262_), .B(new_n12785_), .ZN(new_n21263_));
  NAND2_X1   g18827(.A1(new_n21259_), .A2(pi0618), .ZN(new_n21264_));
  NAND2_X1   g18828(.A1(new_n21232_), .A2(new_n12781_), .ZN(new_n21265_));
  AOI21_X1   g18829(.A1(new_n21264_), .A2(new_n21265_), .B(new_n12785_), .ZN(new_n21266_));
  NOR2_X1    g18830(.A1(new_n21266_), .A2(new_n12779_), .ZN(new_n21267_));
  AND2_X2    g18831(.A1(new_n21267_), .A2(new_n21263_), .Z(new_n21268_));
  NOR2_X1    g18832(.A1(new_n21268_), .A2(new_n21260_), .ZN(new_n21269_));
  NAND2_X1   g18833(.A1(new_n21269_), .A2(new_n12793_), .ZN(new_n21270_));
  NOR2_X1    g18834(.A1(new_n21233_), .A2(new_n12793_), .ZN(new_n21271_));
  INV_X1     g18835(.I(new_n21271_), .ZN(new_n21272_));
  AOI21_X1   g18836(.A1(new_n21270_), .A2(new_n21272_), .B(pi1159), .ZN(new_n21273_));
  NOR3_X1    g18837(.A1(new_n21268_), .A2(new_n12793_), .A3(new_n21260_), .ZN(new_n21274_));
  NOR2_X1    g18838(.A1(new_n21233_), .A2(pi0619), .ZN(new_n21275_));
  OAI21_X1   g18839(.A1(new_n21274_), .A2(new_n21275_), .B(pi1159), .ZN(new_n21276_));
  NAND2_X1   g18840(.A1(new_n21276_), .A2(pi0789), .ZN(new_n21277_));
  OAI22_X1   g18841(.A1(new_n21277_), .A2(new_n21273_), .B1(pi0789), .B2(new_n21269_), .ZN(new_n21278_));
  NAND2_X1   g18842(.A1(new_n21232_), .A2(new_n12818_), .ZN(new_n21279_));
  OAI21_X1   g18843(.A1(new_n21278_), .A2(new_n12818_), .B(new_n21279_), .ZN(new_n21280_));
  AOI21_X1   g18844(.A1(new_n21280_), .A2(new_n13384_), .B(new_n21236_), .ZN(new_n21281_));
  OAI21_X1   g18845(.A1(new_n21281_), .A2(new_n12984_), .B(new_n21235_), .ZN(new_n21282_));
  OAI21_X1   g18846(.A1(new_n21282_), .A2(pi0644), .B(new_n21234_), .ZN(new_n21283_));
  OAI21_X1   g18847(.A1(new_n14125_), .A2(new_n21245_), .B(new_n16218_), .ZN(new_n21284_));
  OAI21_X1   g18848(.A1(new_n14122_), .A2(new_n10688_), .B(new_n3265_), .ZN(new_n21285_));
  NAND2_X1   g18849(.A1(new_n21285_), .A2(new_n2609_), .ZN(new_n21286_));
  NAND2_X1   g18850(.A1(new_n15744_), .A2(new_n10688_), .ZN(new_n21287_));
  AOI21_X1   g18851(.A1(new_n21287_), .A2(new_n21286_), .B(new_n21284_), .ZN(new_n21288_));
  NAND2_X1   g18852(.A1(new_n2609_), .A2(new_n16218_), .ZN(new_n21289_));
  AOI21_X1   g18853(.A1(new_n21233_), .A2(new_n21289_), .B(new_n21288_), .ZN(new_n21290_));
  NAND2_X1   g18854(.A1(new_n21290_), .A2(new_n13521_), .ZN(new_n21291_));
  NAND2_X1   g18855(.A1(new_n21232_), .A2(pi0625), .ZN(new_n21292_));
  AOI21_X1   g18856(.A1(new_n21291_), .A2(new_n21292_), .B(pi1153), .ZN(new_n21293_));
  NAND2_X1   g18857(.A1(new_n21232_), .A2(new_n13521_), .ZN(new_n21294_));
  NAND2_X1   g18858(.A1(new_n21290_), .A2(pi0625), .ZN(new_n21295_));
  AOI21_X1   g18859(.A1(new_n21295_), .A2(new_n21294_), .B(new_n12841_), .ZN(new_n21296_));
  NOR3_X1    g18860(.A1(new_n21293_), .A2(new_n21296_), .A3(new_n12758_), .ZN(new_n21297_));
  NOR2_X1    g18861(.A1(new_n21290_), .A2(pi0778), .ZN(new_n21298_));
  NOR2_X1    g18862(.A1(new_n21297_), .A2(new_n21298_), .ZN(new_n21299_));
  NOR2_X1    g18863(.A1(new_n21299_), .A2(new_n12869_), .ZN(new_n21300_));
  AOI21_X1   g18864(.A1(new_n12869_), .A2(new_n21233_), .B(new_n21300_), .ZN(new_n21301_));
  NAND2_X1   g18865(.A1(new_n21301_), .A2(new_n12888_), .ZN(new_n21302_));
  OAI21_X1   g18866(.A1(new_n12888_), .A2(new_n21233_), .B(new_n21302_), .ZN(new_n21303_));
  INV_X1     g18867(.I(new_n21303_), .ZN(new_n21304_));
  NOR2_X1    g18868(.A1(new_n21232_), .A2(new_n12911_), .ZN(new_n21305_));
  AOI21_X1   g18869(.A1(new_n21304_), .A2(new_n12911_), .B(new_n21305_), .ZN(new_n21306_));
  NAND2_X1   g18870(.A1(new_n21306_), .A2(new_n13392_), .ZN(new_n21307_));
  OAI21_X1   g18871(.A1(new_n13392_), .A2(new_n21233_), .B(new_n21307_), .ZN(new_n21308_));
  NAND2_X1   g18872(.A1(new_n21308_), .A2(new_n12920_), .ZN(new_n21309_));
  NAND2_X1   g18873(.A1(new_n21232_), .A2(pi0628), .ZN(new_n21310_));
  AOI21_X1   g18874(.A1(new_n21309_), .A2(new_n21310_), .B(pi1156), .ZN(new_n21311_));
  NAND2_X1   g18875(.A1(new_n21232_), .A2(new_n12920_), .ZN(new_n21312_));
  NAND2_X1   g18876(.A1(new_n21308_), .A2(pi0628), .ZN(new_n21313_));
  AOI21_X1   g18877(.A1(new_n21313_), .A2(new_n21312_), .B(new_n12742_), .ZN(new_n21314_));
  OR2_X2     g18878(.A1(new_n21314_), .A2(new_n12937_), .Z(new_n21315_));
  OAI22_X1   g18879(.A1(new_n21315_), .A2(new_n21311_), .B1(pi0792), .B2(new_n21308_), .ZN(new_n21316_));
  NAND2_X1   g18880(.A1(new_n21316_), .A2(new_n12741_), .ZN(new_n21317_));
  OAI21_X1   g18881(.A1(new_n12741_), .A2(new_n21232_), .B(new_n21317_), .ZN(new_n21318_));
  NOR2_X1    g18882(.A1(new_n21318_), .A2(pi1157), .ZN(new_n21319_));
  NAND2_X1   g18883(.A1(new_n21316_), .A2(pi0647), .ZN(new_n21320_));
  OAI21_X1   g18884(.A1(pi0647), .A2(new_n21232_), .B(new_n21320_), .ZN(new_n21321_));
  NOR2_X1    g18885(.A1(new_n21321_), .A2(new_n12965_), .ZN(new_n21322_));
  OAI21_X1   g18886(.A1(new_n21319_), .A2(new_n21322_), .B(pi0787), .ZN(new_n21323_));
  OAI21_X1   g18887(.A1(pi0787), .A2(new_n21316_), .B(new_n21323_), .ZN(new_n21324_));
  OAI21_X1   g18888(.A1(new_n21324_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n21325_));
  NAND3_X1   g18889(.A1(new_n21325_), .A2(new_n12739_), .A3(new_n21283_), .ZN(new_n21326_));
  AOI21_X1   g18890(.A1(new_n21233_), .A2(new_n12975_), .B(pi0715), .ZN(new_n21327_));
  OAI21_X1   g18891(.A1(new_n21282_), .A2(new_n12975_), .B(new_n21327_), .ZN(new_n21328_));
  OAI21_X1   g18892(.A1(new_n21324_), .A2(pi0644), .B(pi0715), .ZN(new_n21329_));
  NAND3_X1   g18893(.A1(new_n21329_), .A2(pi1160), .A3(new_n21328_), .ZN(new_n21330_));
  AOI21_X1   g18894(.A1(new_n21326_), .A2(new_n21330_), .B(new_n13000_), .ZN(new_n21331_));
  NAND2_X1   g18895(.A1(new_n21233_), .A2(pi0626), .ZN(new_n21332_));
  NAND2_X1   g18896(.A1(new_n21278_), .A2(new_n12747_), .ZN(new_n21333_));
  AOI21_X1   g18897(.A1(new_n21333_), .A2(new_n21332_), .B(new_n12816_), .ZN(new_n21334_));
  NOR2_X1    g18898(.A1(new_n21232_), .A2(pi0626), .ZN(new_n21335_));
  AOI21_X1   g18899(.A1(new_n21278_), .A2(pi0626), .B(new_n21335_), .ZN(new_n21336_));
  OAI22_X1   g18900(.A1(new_n21336_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n21306_), .ZN(new_n21337_));
  OAI21_X1   g18901(.A1(new_n21337_), .A2(new_n21334_), .B(pi0788), .ZN(new_n21338_));
  NAND2_X1   g18902(.A1(new_n21338_), .A2(new_n15824_), .ZN(new_n21339_));
  NAND2_X1   g18903(.A1(new_n21299_), .A2(new_n12766_), .ZN(new_n21340_));
  AOI21_X1   g18904(.A1(new_n16210_), .A2(new_n13566_), .B(new_n15826_), .ZN(new_n21341_));
  AOI21_X1   g18905(.A1(new_n14328_), .A2(new_n21106_), .B(new_n10688_), .ZN(new_n21342_));
  AOI21_X1   g18906(.A1(new_n21342_), .A2(new_n5336_), .B(new_n3265_), .ZN(new_n21343_));
  OAI21_X1   g18907(.A1(new_n21341_), .A2(pi0185), .B(new_n21343_), .ZN(new_n21344_));
  NAND2_X1   g18908(.A1(new_n14172_), .A2(pi0185), .ZN(new_n21345_));
  NAND2_X1   g18909(.A1(new_n14174_), .A2(new_n10688_), .ZN(new_n21346_));
  AOI21_X1   g18910(.A1(new_n21345_), .A2(new_n21346_), .B(pi0751), .ZN(new_n21347_));
  NAND2_X1   g18911(.A1(new_n15835_), .A2(pi0185), .ZN(new_n21348_));
  NAND2_X1   g18912(.A1(new_n14177_), .A2(new_n10688_), .ZN(new_n21349_));
  AOI21_X1   g18913(.A1(new_n21349_), .A2(new_n21348_), .B(new_n16210_), .ZN(new_n21350_));
  OAI21_X1   g18914(.A1(new_n21350_), .A2(new_n21347_), .B(new_n2627_), .ZN(new_n21351_));
  NOR2_X1    g18915(.A1(new_n14182_), .A2(pi0185), .ZN(new_n21352_));
  NOR2_X1    g18916(.A1(new_n14184_), .A2(new_n10688_), .ZN(new_n21353_));
  OAI21_X1   g18917(.A1(new_n21352_), .A2(new_n21353_), .B(pi0751), .ZN(new_n21354_));
  NOR2_X1    g18918(.A1(new_n14187_), .A2(new_n10688_), .ZN(new_n21355_));
  NOR2_X1    g18919(.A1(new_n14189_), .A2(pi0185), .ZN(new_n21356_));
  OAI21_X1   g18920(.A1(new_n21355_), .A2(new_n21356_), .B(new_n16210_), .ZN(new_n21357_));
  NAND3_X1   g18921(.A1(new_n21357_), .A2(new_n21354_), .A3(pi0039), .ZN(new_n21358_));
  NAND3_X1   g18922(.A1(new_n21358_), .A2(new_n3265_), .A3(new_n21351_), .ZN(new_n21359_));
  NAND3_X1   g18923(.A1(new_n21359_), .A2(new_n16218_), .A3(new_n21344_), .ZN(new_n21360_));
  NAND2_X1   g18924(.A1(new_n21248_), .A2(pi0701), .ZN(new_n21361_));
  NAND3_X1   g18925(.A1(new_n21361_), .A2(new_n21360_), .A3(new_n2609_), .ZN(new_n21362_));
  AOI21_X1   g18926(.A1(new_n21362_), .A2(new_n21237_), .B(pi0778), .ZN(new_n21363_));
  INV_X1     g18927(.I(new_n21293_), .ZN(new_n21364_));
  NAND2_X1   g18928(.A1(new_n21249_), .A2(pi0625), .ZN(new_n21365_));
  NAND2_X1   g18929(.A1(new_n21362_), .A2(new_n21237_), .ZN(new_n21366_));
  NAND2_X1   g18930(.A1(new_n21366_), .A2(new_n13521_), .ZN(new_n21367_));
  NAND2_X1   g18931(.A1(new_n21367_), .A2(new_n21365_), .ZN(new_n21368_));
  AOI21_X1   g18932(.A1(new_n21368_), .A2(new_n12841_), .B(new_n21296_), .ZN(new_n21369_));
  NAND2_X1   g18933(.A1(new_n21249_), .A2(new_n13521_), .ZN(new_n21370_));
  NAND2_X1   g18934(.A1(new_n21366_), .A2(pi0625), .ZN(new_n21371_));
  NAND2_X1   g18935(.A1(new_n21371_), .A2(new_n21370_), .ZN(new_n21372_));
  AOI21_X1   g18936(.A1(new_n21372_), .A2(pi1153), .B(new_n13560_), .ZN(new_n21373_));
  AOI22_X1   g18937(.A1(new_n13560_), .A2(new_n21369_), .B1(new_n21373_), .B2(new_n21364_), .ZN(new_n21374_));
  AOI21_X1   g18938(.A1(new_n21374_), .A2(pi0778), .B(new_n21363_), .ZN(new_n21375_));
  OAI21_X1   g18939(.A1(new_n21375_), .A2(new_n12766_), .B(new_n21340_), .ZN(new_n21376_));
  AOI21_X1   g18940(.A1(new_n21376_), .A2(pi1155), .B(new_n21255_), .ZN(new_n21377_));
  NOR2_X1    g18941(.A1(new_n21375_), .A2(pi0609), .ZN(new_n21378_));
  NOR3_X1    g18942(.A1(new_n21297_), .A2(new_n12766_), .A3(new_n21298_), .ZN(new_n21379_));
  OAI21_X1   g18943(.A1(new_n21378_), .A2(new_n21379_), .B(new_n12770_), .ZN(new_n21380_));
  NOR2_X1    g18944(.A1(new_n21257_), .A2(pi0660), .ZN(new_n21381_));
  AOI22_X1   g18945(.A1(new_n21377_), .A2(pi0660), .B1(new_n21380_), .B2(new_n21381_), .ZN(new_n21382_));
  NOR2_X1    g18946(.A1(new_n21375_), .A2(pi0785), .ZN(new_n21383_));
  AOI21_X1   g18947(.A1(new_n21382_), .A2(pi0785), .B(new_n21383_), .ZN(new_n21384_));
  NOR2_X1    g18948(.A1(new_n21384_), .A2(pi0781), .ZN(new_n21385_));
  AND2_X2    g18949(.A1(new_n21301_), .A2(new_n12781_), .Z(new_n21386_));
  NOR2_X1    g18950(.A1(new_n21384_), .A2(new_n12781_), .ZN(new_n21387_));
  OAI21_X1   g18951(.A1(new_n21387_), .A2(new_n21386_), .B(pi1154), .ZN(new_n21388_));
  NAND3_X1   g18952(.A1(new_n21388_), .A2(pi0627), .A3(new_n21263_), .ZN(new_n21389_));
  NAND2_X1   g18953(.A1(new_n21301_), .A2(pi0618), .ZN(new_n21390_));
  OAI21_X1   g18954(.A1(new_n21384_), .A2(pi0618), .B(new_n21390_), .ZN(new_n21391_));
  AOI21_X1   g18955(.A1(new_n21391_), .A2(new_n12785_), .B(new_n21266_), .ZN(new_n21392_));
  AOI21_X1   g18956(.A1(new_n21392_), .A2(new_n12880_), .B(new_n12779_), .ZN(new_n21393_));
  AOI21_X1   g18957(.A1(new_n21393_), .A2(new_n21389_), .B(new_n21385_), .ZN(new_n21394_));
  OAI21_X1   g18958(.A1(new_n21394_), .A2(pi0789), .B(new_n12819_), .ZN(new_n21395_));
  NOR2_X1    g18959(.A1(new_n21304_), .A2(new_n12793_), .ZN(new_n21396_));
  NOR2_X1    g18960(.A1(new_n21394_), .A2(pi0619), .ZN(new_n21397_));
  OAI21_X1   g18961(.A1(new_n21397_), .A2(new_n21396_), .B(new_n12791_), .ZN(new_n21398_));
  NAND3_X1   g18962(.A1(new_n21398_), .A2(new_n12895_), .A3(new_n21276_), .ZN(new_n21399_));
  INV_X1     g18963(.I(new_n21273_), .ZN(new_n21400_));
  NAND2_X1   g18964(.A1(new_n21303_), .A2(new_n12793_), .ZN(new_n21401_));
  OAI21_X1   g18965(.A1(new_n21394_), .A2(new_n12793_), .B(new_n21401_), .ZN(new_n21402_));
  AOI21_X1   g18966(.A1(new_n21402_), .A2(pi1159), .B(new_n12895_), .ZN(new_n21403_));
  AOI21_X1   g18967(.A1(new_n21403_), .A2(new_n21400_), .B(new_n12796_), .ZN(new_n21404_));
  AOI21_X1   g18968(.A1(new_n21404_), .A2(new_n21399_), .B(new_n21395_), .ZN(new_n21405_));
  NOR2_X1    g18969(.A1(new_n21314_), .A2(pi0629), .ZN(new_n21406_));
  NOR2_X1    g18970(.A1(new_n21311_), .A2(new_n12919_), .ZN(new_n21407_));
  NOR2_X1    g18971(.A1(new_n21406_), .A2(new_n21407_), .ZN(new_n21408_));
  AOI21_X1   g18972(.A1(new_n21280_), .A2(new_n19160_), .B(new_n21408_), .ZN(new_n21409_));
  OAI22_X1   g18973(.A1(new_n21405_), .A2(new_n21339_), .B1(new_n12937_), .B2(new_n21409_), .ZN(new_n21410_));
  AOI21_X1   g18974(.A1(new_n21328_), .A2(pi1160), .B(new_n12975_), .ZN(new_n21411_));
  AOI21_X1   g18975(.A1(new_n21283_), .A2(new_n12739_), .B(pi0644), .ZN(new_n21412_));
  NOR2_X1    g18976(.A1(new_n21411_), .A2(new_n21412_), .ZN(new_n21413_));
  OAI22_X1   g18977(.A1(new_n15576_), .A2(new_n21321_), .B1(new_n21318_), .B2(new_n15730_), .ZN(new_n21414_));
  NOR2_X1    g18978(.A1(new_n21281_), .A2(new_n17212_), .ZN(new_n21415_));
  NOR2_X1    g18979(.A1(new_n21414_), .A2(new_n21415_), .ZN(new_n21416_));
  OAI22_X1   g18980(.A1(new_n21413_), .A2(new_n13000_), .B1(new_n21416_), .B2(new_n12972_), .ZN(new_n21417_));
  AOI21_X1   g18981(.A1(new_n21410_), .A2(new_n15693_), .B(new_n21417_), .ZN(new_n21418_));
  OAI21_X1   g18982(.A1(new_n21331_), .A2(new_n21418_), .B(new_n6643_), .ZN(new_n21419_));
  AOI22_X1   g18983(.A1(new_n21419_), .A2(new_n21231_), .B1(pi0832), .B2(new_n21230_), .ZN(po0342));
  NOR2_X1    g18984(.A1(new_n3042_), .A2(pi0186), .ZN(new_n21421_));
  INV_X1     g18985(.I(new_n21421_), .ZN(new_n21422_));
  AOI21_X1   g18986(.A1(new_n12756_), .A2(new_n16803_), .B(new_n21421_), .ZN(new_n21423_));
  NOR3_X1    g18987(.A1(new_n21423_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n21424_));
  NOR2_X1    g18988(.A1(new_n21423_), .A2(new_n12762_), .ZN(new_n21425_));
  AOI21_X1   g18989(.A1(new_n21425_), .A2(new_n12768_), .B(pi1155), .ZN(new_n21426_));
  INV_X1     g18990(.I(new_n21423_), .ZN(new_n21427_));
  AOI21_X1   g18991(.A1(new_n21427_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n21428_));
  NOR3_X1    g18992(.A1(new_n21426_), .A2(new_n21428_), .A3(new_n12764_), .ZN(new_n21429_));
  NOR2_X1    g18993(.A1(new_n21429_), .A2(new_n21424_), .ZN(new_n21430_));
  NOR2_X1    g18994(.A1(new_n21430_), .A2(pi0781), .ZN(new_n21431_));
  INV_X1     g18995(.I(new_n21430_), .ZN(new_n21432_));
  AOI21_X1   g18996(.A1(new_n21432_), .A2(new_n12783_), .B(pi1154), .ZN(new_n21433_));
  AOI21_X1   g18997(.A1(new_n21432_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n21434_));
  NOR3_X1    g18998(.A1(new_n21433_), .A2(new_n21434_), .A3(new_n12779_), .ZN(new_n21435_));
  NOR2_X1    g18999(.A1(new_n21435_), .A2(new_n21431_), .ZN(new_n21436_));
  NOR3_X1    g19000(.A1(new_n21435_), .A2(pi0619), .A3(new_n21431_), .ZN(new_n21437_));
  NOR2_X1    g19001(.A1(new_n21421_), .A2(new_n12793_), .ZN(new_n21438_));
  OAI21_X1   g19002(.A1(new_n21437_), .A2(new_n21438_), .B(new_n12791_), .ZN(new_n21439_));
  NAND2_X1   g19003(.A1(new_n21436_), .A2(pi0619), .ZN(new_n21440_));
  NAND2_X1   g19004(.A1(new_n21422_), .A2(new_n12793_), .ZN(new_n21441_));
  AOI21_X1   g19005(.A1(new_n21440_), .A2(new_n21441_), .B(new_n12791_), .ZN(new_n21442_));
  INV_X1     g19006(.I(new_n21442_), .ZN(new_n21443_));
  NAND3_X1   g19007(.A1(new_n21443_), .A2(pi0789), .A3(new_n21439_), .ZN(new_n21444_));
  OAI21_X1   g19008(.A1(pi0789), .A2(new_n21436_), .B(new_n21444_), .ZN(new_n21445_));
  NOR2_X1    g19009(.A1(new_n21445_), .A2(new_n12818_), .ZN(new_n21446_));
  AOI21_X1   g19010(.A1(new_n12818_), .A2(new_n21422_), .B(new_n21446_), .ZN(new_n21447_));
  AOI21_X1   g19011(.A1(new_n12826_), .A2(pi0703), .B(new_n21421_), .ZN(new_n21448_));
  NOR2_X1    g19012(.A1(new_n21448_), .A2(pi0778), .ZN(new_n21449_));
  NOR2_X1    g19013(.A1(new_n12834_), .A2(new_n16795_), .ZN(new_n21450_));
  INV_X1     g19014(.I(new_n21450_), .ZN(new_n21451_));
  NOR2_X1    g19015(.A1(new_n21421_), .A2(pi1153), .ZN(new_n21452_));
  NAND2_X1   g19016(.A1(new_n21451_), .A2(new_n21452_), .ZN(new_n21453_));
  INV_X1     g19017(.I(new_n21453_), .ZN(new_n21454_));
  NOR2_X1    g19018(.A1(new_n21450_), .A2(new_n21448_), .ZN(new_n21455_));
  NOR2_X1    g19019(.A1(new_n21455_), .A2(new_n12841_), .ZN(new_n21456_));
  NOR2_X1    g19020(.A1(new_n21454_), .A2(new_n21456_), .ZN(new_n21457_));
  AOI21_X1   g19021(.A1(new_n21457_), .A2(pi0778), .B(new_n21449_), .ZN(new_n21458_));
  NOR2_X1    g19022(.A1(new_n21458_), .A2(new_n12871_), .ZN(new_n21459_));
  INV_X1     g19023(.I(new_n21459_), .ZN(new_n21460_));
  NOR2_X1    g19024(.A1(new_n21460_), .A2(new_n12889_), .ZN(new_n21461_));
  NAND2_X1   g19025(.A1(new_n21461_), .A2(new_n18203_), .ZN(new_n21462_));
  NOR2_X1    g19026(.A1(new_n21462_), .A2(new_n17884_), .ZN(new_n21463_));
  AOI22_X1   g19027(.A1(new_n21447_), .A2(new_n12949_), .B1(new_n15695_), .B2(new_n21463_), .ZN(new_n21464_));
  NOR2_X1    g19028(.A1(new_n21464_), .A2(pi0629), .ZN(new_n21465_));
  AOI22_X1   g19029(.A1(new_n21447_), .A2(new_n12948_), .B1(new_n15700_), .B2(new_n21463_), .ZN(new_n21466_));
  NOR2_X1    g19030(.A1(new_n21466_), .A2(new_n12919_), .ZN(new_n21467_));
  NOR2_X1    g19031(.A1(new_n21465_), .A2(new_n21467_), .ZN(new_n21468_));
  NOR2_X1    g19032(.A1(new_n21448_), .A2(new_n12754_), .ZN(new_n21469_));
  NOR2_X1    g19033(.A1(new_n21469_), .A2(new_n21427_), .ZN(new_n21470_));
  NAND2_X1   g19034(.A1(new_n21470_), .A2(new_n12758_), .ZN(new_n21471_));
  NAND2_X1   g19035(.A1(new_n21469_), .A2(pi0625), .ZN(new_n21472_));
  NAND3_X1   g19036(.A1(new_n21472_), .A2(pi1153), .A3(new_n21423_), .ZN(new_n21473_));
  AND3_X2    g19037(.A1(new_n21453_), .A2(pi0608), .A3(new_n21473_), .Z(new_n21474_));
  NOR2_X1    g19038(.A1(new_n21456_), .A2(pi0608), .ZN(new_n21475_));
  INV_X1     g19039(.I(new_n21472_), .ZN(new_n21476_));
  OAI21_X1   g19040(.A1(new_n21476_), .A2(new_n21470_), .B(new_n21452_), .ZN(new_n21477_));
  NAND2_X1   g19041(.A1(new_n21475_), .A2(new_n21477_), .ZN(new_n21478_));
  NAND2_X1   g19042(.A1(new_n21478_), .A2(pi0778), .ZN(new_n21479_));
  OAI21_X1   g19043(.A1(new_n21479_), .A2(new_n21474_), .B(new_n21471_), .ZN(new_n21480_));
  INV_X1     g19044(.I(new_n21480_), .ZN(new_n21481_));
  NAND2_X1   g19045(.A1(new_n21458_), .A2(new_n12766_), .ZN(new_n21482_));
  OAI21_X1   g19046(.A1(new_n21481_), .A2(new_n12766_), .B(new_n21482_), .ZN(new_n21483_));
  AOI21_X1   g19047(.A1(new_n21483_), .A2(pi1155), .B(new_n21426_), .ZN(new_n21484_));
  NAND2_X1   g19048(.A1(new_n21480_), .A2(new_n12766_), .ZN(new_n21485_));
  NAND2_X1   g19049(.A1(new_n21458_), .A2(pi0609), .ZN(new_n21486_));
  AOI21_X1   g19050(.A1(new_n21485_), .A2(new_n21486_), .B(pi1155), .ZN(new_n21487_));
  NOR3_X1    g19051(.A1(new_n21487_), .A2(pi0660), .A3(new_n21428_), .ZN(new_n21488_));
  AOI21_X1   g19052(.A1(pi0660), .A2(new_n21484_), .B(new_n21488_), .ZN(new_n21489_));
  NAND2_X1   g19053(.A1(new_n21489_), .A2(pi0785), .ZN(new_n21490_));
  OAI21_X1   g19054(.A1(pi0785), .A2(new_n21481_), .B(new_n21490_), .ZN(new_n21491_));
  INV_X1     g19055(.I(new_n21491_), .ZN(new_n21492_));
  NAND2_X1   g19056(.A1(new_n21460_), .A2(pi0618), .ZN(new_n21493_));
  OAI21_X1   g19057(.A1(new_n21492_), .A2(pi0618), .B(new_n21493_), .ZN(new_n21494_));
  AOI21_X1   g19058(.A1(new_n21494_), .A2(new_n12785_), .B(new_n21434_), .ZN(new_n21495_));
  NOR2_X1    g19059(.A1(new_n21459_), .A2(pi0618), .ZN(new_n21496_));
  NOR2_X1    g19060(.A1(new_n21492_), .A2(new_n12781_), .ZN(new_n21497_));
  OAI21_X1   g19061(.A1(new_n21497_), .A2(new_n21496_), .B(pi1154), .ZN(new_n21498_));
  NOR2_X1    g19062(.A1(new_n21433_), .A2(new_n12880_), .ZN(new_n21499_));
  AOI22_X1   g19063(.A1(new_n21495_), .A2(new_n12880_), .B1(new_n21498_), .B2(new_n21499_), .ZN(new_n21500_));
  NAND2_X1   g19064(.A1(new_n21500_), .A2(pi0781), .ZN(new_n21501_));
  NAND2_X1   g19065(.A1(new_n21491_), .A2(new_n12779_), .ZN(new_n21502_));
  NAND2_X1   g19066(.A1(new_n21501_), .A2(new_n21502_), .ZN(new_n21503_));
  AOI21_X1   g19067(.A1(new_n21503_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n21504_));
  NOR2_X1    g19068(.A1(new_n21461_), .A2(pi0619), .ZN(new_n21505_));
  INV_X1     g19069(.I(new_n21503_), .ZN(new_n21506_));
  NOR2_X1    g19070(.A1(new_n21506_), .A2(new_n12793_), .ZN(new_n21507_));
  OAI21_X1   g19071(.A1(new_n21507_), .A2(new_n21505_), .B(pi1159), .ZN(new_n21508_));
  NAND3_X1   g19072(.A1(new_n21508_), .A2(pi0648), .A3(new_n21439_), .ZN(new_n21509_));
  NOR2_X1    g19073(.A1(new_n21506_), .A2(pi0619), .ZN(new_n21510_));
  NOR2_X1    g19074(.A1(new_n21461_), .A2(new_n12793_), .ZN(new_n21511_));
  OAI21_X1   g19075(.A1(new_n21510_), .A2(new_n21511_), .B(new_n12791_), .ZN(new_n21512_));
  NAND3_X1   g19076(.A1(new_n21512_), .A2(new_n12895_), .A3(new_n21443_), .ZN(new_n21513_));
  NAND3_X1   g19077(.A1(new_n21509_), .A2(new_n21513_), .A3(pi0789), .ZN(new_n21514_));
  NOR2_X1    g19078(.A1(new_n21422_), .A2(new_n12747_), .ZN(new_n21515_));
  INV_X1     g19079(.I(new_n21445_), .ZN(new_n21516_));
  NOR2_X1    g19080(.A1(new_n21516_), .A2(pi0626), .ZN(new_n21517_));
  OAI21_X1   g19081(.A1(new_n21517_), .A2(new_n21515_), .B(new_n12815_), .ZN(new_n21518_));
  INV_X1     g19082(.I(new_n21462_), .ZN(new_n21519_));
  NAND2_X1   g19083(.A1(new_n21421_), .A2(new_n12747_), .ZN(new_n21520_));
  OAI21_X1   g19084(.A1(new_n21516_), .A2(new_n12747_), .B(new_n21520_), .ZN(new_n21521_));
  AOI22_X1   g19085(.A1(new_n21521_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n21519_), .ZN(new_n21522_));
  NAND2_X1   g19086(.A1(new_n21522_), .A2(new_n21518_), .ZN(new_n21523_));
  AOI22_X1   g19087(.A1(new_n21514_), .A2(new_n21504_), .B1(pi0788), .B2(new_n21523_), .ZN(new_n21524_));
  OAI22_X1   g19088(.A1(new_n21524_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n21468_), .ZN(new_n21525_));
  INV_X1     g19089(.I(new_n21447_), .ZN(new_n21526_));
  NAND2_X1   g19090(.A1(new_n21526_), .A2(new_n13384_), .ZN(new_n21527_));
  NAND2_X1   g19091(.A1(new_n12943_), .A2(new_n21422_), .ZN(new_n21528_));
  NAND2_X1   g19092(.A1(new_n21527_), .A2(new_n21528_), .ZN(new_n21529_));
  NAND2_X1   g19093(.A1(new_n21463_), .A2(new_n12954_), .ZN(new_n21530_));
  NAND2_X1   g19094(.A1(new_n21530_), .A2(new_n12741_), .ZN(new_n21531_));
  NOR2_X1    g19095(.A1(new_n21421_), .A2(new_n12741_), .ZN(new_n21532_));
  INV_X1     g19096(.I(new_n21532_), .ZN(new_n21533_));
  AOI21_X1   g19097(.A1(new_n21531_), .A2(new_n21533_), .B(pi1157), .ZN(new_n21534_));
  INV_X1     g19098(.I(new_n21534_), .ZN(new_n21535_));
  NAND2_X1   g19099(.A1(new_n21421_), .A2(new_n12741_), .ZN(new_n21536_));
  OAI21_X1   g19100(.A1(new_n21530_), .A2(new_n12741_), .B(new_n21536_), .ZN(new_n21537_));
  OAI22_X1   g19101(.A1(new_n21535_), .A2(new_n12981_), .B1(new_n21537_), .B2(new_n15576_), .ZN(new_n21538_));
  AOI21_X1   g19102(.A1(new_n21529_), .A2(new_n15608_), .B(new_n21538_), .ZN(new_n21539_));
  OAI22_X1   g19103(.A1(new_n21525_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n21539_), .ZN(new_n21540_));
  NAND2_X1   g19104(.A1(new_n21540_), .A2(new_n13000_), .ZN(new_n21541_));
  AND2_X2    g19105(.A1(new_n21540_), .A2(new_n12975_), .Z(new_n21542_));
  OAI21_X1   g19106(.A1(new_n12965_), .A2(new_n21537_), .B(new_n21535_), .ZN(new_n21543_));
  NAND3_X1   g19107(.A1(new_n21463_), .A2(new_n12972_), .A3(new_n12954_), .ZN(new_n21544_));
  OAI21_X1   g19108(.A1(new_n21543_), .A2(new_n12972_), .B(new_n21544_), .ZN(new_n21545_));
  NOR2_X1    g19109(.A1(new_n21545_), .A2(new_n12975_), .ZN(new_n21546_));
  OAI21_X1   g19110(.A1(new_n21542_), .A2(new_n21546_), .B(new_n12740_), .ZN(new_n21547_));
  NOR2_X1    g19111(.A1(new_n21421_), .A2(new_n12975_), .ZN(new_n21548_));
  NOR2_X1    g19112(.A1(new_n17611_), .A2(new_n21421_), .ZN(new_n21549_));
  AOI21_X1   g19113(.A1(new_n21526_), .A2(new_n17611_), .B(new_n21549_), .ZN(new_n21550_));
  NOR2_X1    g19114(.A1(new_n21550_), .A2(pi0644), .ZN(new_n21551_));
  OAI21_X1   g19115(.A1(new_n21551_), .A2(new_n21548_), .B(pi0715), .ZN(new_n21552_));
  NAND3_X1   g19116(.A1(new_n21547_), .A2(new_n12739_), .A3(new_n21552_), .ZN(new_n21553_));
  NOR2_X1    g19117(.A1(new_n21545_), .A2(pi0644), .ZN(new_n21554_));
  AOI21_X1   g19118(.A1(new_n21540_), .A2(pi0644), .B(new_n21554_), .ZN(new_n21555_));
  NAND2_X1   g19119(.A1(new_n21422_), .A2(new_n12975_), .ZN(new_n21556_));
  OAI21_X1   g19120(.A1(new_n21550_), .A2(new_n12975_), .B(new_n21556_), .ZN(new_n21557_));
  AOI21_X1   g19121(.A1(new_n21557_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n21558_));
  OAI21_X1   g19122(.A1(new_n21555_), .A2(new_n12740_), .B(new_n21558_), .ZN(new_n21559_));
  NAND3_X1   g19123(.A1(new_n21553_), .A2(pi0790), .A3(new_n21559_), .ZN(new_n21560_));
  AOI21_X1   g19124(.A1(new_n21560_), .A2(new_n21541_), .B(new_n12738_), .ZN(new_n21561_));
  AOI21_X1   g19125(.A1(po1038), .A2(new_n7381_), .B(pi0832), .ZN(new_n21562_));
  NOR2_X1    g19126(.A1(new_n13193_), .A2(pi0186), .ZN(new_n21563_));
  AOI21_X1   g19127(.A1(new_n21563_), .A2(pi0644), .B(new_n12740_), .ZN(new_n21564_));
  NOR2_X1    g19128(.A1(new_n21563_), .A2(new_n13384_), .ZN(new_n21565_));
  INV_X1     g19129(.I(new_n21565_), .ZN(new_n21566_));
  INV_X1     g19130(.I(new_n21563_), .ZN(new_n21567_));
  NOR2_X1    g19131(.A1(new_n2609_), .A2(new_n7381_), .ZN(new_n21568_));
  INV_X1     g19132(.I(new_n21568_), .ZN(new_n21569_));
  NAND2_X1   g19133(.A1(new_n15009_), .A2(pi0186), .ZN(new_n21570_));
  NOR2_X1    g19134(.A1(pi0186), .A2(pi0752), .ZN(new_n21571_));
  NAND2_X1   g19135(.A1(new_n15013_), .A2(new_n21571_), .ZN(new_n21572_));
  AOI21_X1   g19136(.A1(new_n21572_), .A2(new_n21570_), .B(new_n15008_), .ZN(new_n21573_));
  AOI21_X1   g19137(.A1(new_n13395_), .A2(new_n7381_), .B(new_n16803_), .ZN(new_n21574_));
  OAI21_X1   g19138(.A1(new_n21573_), .A2(new_n21574_), .B(new_n2609_), .ZN(new_n21575_));
  AOI21_X1   g19139(.A1(new_n21575_), .A2(new_n21569_), .B(new_n12760_), .ZN(new_n21576_));
  NOR2_X1    g19140(.A1(new_n21563_), .A2(new_n12761_), .ZN(new_n21577_));
  NOR2_X1    g19141(.A1(new_n21576_), .A2(new_n21577_), .ZN(new_n21578_));
  AOI22_X1   g19142(.A1(new_n21576_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n21567_), .ZN(new_n21579_));
  OR2_X2     g19143(.A1(new_n21579_), .A2(pi1155), .Z(new_n21580_));
  AOI22_X1   g19144(.A1(new_n21576_), .A2(pi0609), .B1(new_n13357_), .B2(new_n21567_), .ZN(new_n21581_));
  NOR2_X1    g19145(.A1(new_n21581_), .A2(new_n12770_), .ZN(new_n21582_));
  NOR2_X1    g19146(.A1(new_n21582_), .A2(new_n12764_), .ZN(new_n21583_));
  AOI22_X1   g19147(.A1(new_n21583_), .A2(new_n21580_), .B1(new_n12764_), .B2(new_n21578_), .ZN(new_n21584_));
  NOR2_X1    g19148(.A1(new_n21563_), .A2(new_n12781_), .ZN(new_n21585_));
  AOI21_X1   g19149(.A1(new_n21584_), .A2(new_n12781_), .B(new_n21585_), .ZN(new_n21586_));
  NOR2_X1    g19150(.A1(new_n21586_), .A2(pi1154), .ZN(new_n21587_));
  NAND2_X1   g19151(.A1(new_n21584_), .A2(pi0618), .ZN(new_n21588_));
  OAI21_X1   g19152(.A1(pi0618), .A2(new_n21563_), .B(new_n21588_), .ZN(new_n21589_));
  NAND2_X1   g19153(.A1(new_n21589_), .A2(pi1154), .ZN(new_n21590_));
  NAND2_X1   g19154(.A1(new_n21590_), .A2(pi0781), .ZN(new_n21591_));
  OAI22_X1   g19155(.A1(new_n21591_), .A2(new_n21587_), .B1(pi0781), .B2(new_n21584_), .ZN(new_n21592_));
  NAND2_X1   g19156(.A1(new_n21592_), .A2(new_n12796_), .ZN(new_n21593_));
  NAND2_X1   g19157(.A1(new_n21567_), .A2(pi0619), .ZN(new_n21594_));
  OAI21_X1   g19158(.A1(new_n21592_), .A2(pi0619), .B(new_n21594_), .ZN(new_n21595_));
  NAND2_X1   g19159(.A1(new_n21595_), .A2(new_n12791_), .ZN(new_n21596_));
  NAND2_X1   g19160(.A1(new_n21567_), .A2(new_n12793_), .ZN(new_n21597_));
  OAI21_X1   g19161(.A1(new_n21592_), .A2(new_n12793_), .B(new_n21597_), .ZN(new_n21598_));
  AOI21_X1   g19162(.A1(new_n21598_), .A2(pi1159), .B(new_n12796_), .ZN(new_n21599_));
  NAND2_X1   g19163(.A1(new_n21599_), .A2(new_n21596_), .ZN(new_n21600_));
  AND3_X2    g19164(.A1(new_n21600_), .A2(new_n17504_), .A3(new_n21593_), .Z(new_n21601_));
  AOI21_X1   g19165(.A1(new_n12818_), .A2(new_n21567_), .B(new_n21601_), .ZN(new_n21602_));
  OAI21_X1   g19166(.A1(new_n21602_), .A2(new_n12943_), .B(new_n21566_), .ZN(new_n21603_));
  NAND2_X1   g19167(.A1(new_n21563_), .A2(new_n12984_), .ZN(new_n21604_));
  OAI21_X1   g19168(.A1(new_n21603_), .A2(new_n12984_), .B(new_n21604_), .ZN(new_n21605_));
  NAND2_X1   g19169(.A1(new_n21605_), .A2(new_n12975_), .ZN(new_n21606_));
  AOI21_X1   g19170(.A1(new_n21606_), .A2(new_n21564_), .B(pi1160), .ZN(new_n21607_));
  NOR2_X1    g19171(.A1(new_n21567_), .A2(new_n12870_), .ZN(new_n21608_));
  AOI21_X1   g19172(.A1(new_n14117_), .A2(new_n14116_), .B(pi0186), .ZN(new_n21609_));
  AOI21_X1   g19173(.A1(new_n14121_), .A2(new_n14120_), .B(new_n7381_), .ZN(new_n21610_));
  OAI21_X1   g19174(.A1(new_n21609_), .A2(new_n21610_), .B(new_n3265_), .ZN(new_n21611_));
  NAND2_X1   g19175(.A1(new_n13397_), .A2(new_n7381_), .ZN(new_n21612_));
  AOI21_X1   g19176(.A1(new_n13399_), .A2(new_n21612_), .B(new_n16795_), .ZN(new_n21613_));
  NAND2_X1   g19177(.A1(new_n21611_), .A2(new_n21613_), .ZN(new_n21614_));
  NAND3_X1   g19178(.A1(new_n13395_), .A2(new_n7381_), .A3(new_n16795_), .ZN(new_n21615_));
  NAND3_X1   g19179(.A1(new_n21614_), .A2(new_n21615_), .A3(new_n2609_), .ZN(new_n21616_));
  NAND2_X1   g19180(.A1(new_n21616_), .A2(new_n21569_), .ZN(new_n21617_));
  NAND2_X1   g19181(.A1(new_n21617_), .A2(new_n13521_), .ZN(new_n21618_));
  NAND2_X1   g19182(.A1(new_n21567_), .A2(pi0625), .ZN(new_n21619_));
  AOI21_X1   g19183(.A1(new_n21618_), .A2(new_n21619_), .B(pi1153), .ZN(new_n21620_));
  AOI21_X1   g19184(.A1(new_n21616_), .A2(new_n21569_), .B(new_n13521_), .ZN(new_n21621_));
  NOR2_X1    g19185(.A1(new_n21563_), .A2(pi0625), .ZN(new_n21622_));
  OAI21_X1   g19186(.A1(new_n21621_), .A2(new_n21622_), .B(pi1153), .ZN(new_n21623_));
  NAND2_X1   g19187(.A1(new_n21623_), .A2(pi0778), .ZN(new_n21624_));
  OAI22_X1   g19188(.A1(new_n21624_), .A2(new_n21620_), .B1(pi0778), .B2(new_n21617_), .ZN(new_n21625_));
  AOI21_X1   g19189(.A1(new_n21625_), .A2(new_n12870_), .B(new_n21608_), .ZN(new_n21626_));
  NOR2_X1    g19190(.A1(new_n21563_), .A2(new_n12888_), .ZN(new_n21627_));
  AOI21_X1   g19191(.A1(new_n21626_), .A2(new_n12888_), .B(new_n21627_), .ZN(new_n21628_));
  NOR2_X1    g19192(.A1(new_n21567_), .A2(new_n12911_), .ZN(new_n21629_));
  AOI21_X1   g19193(.A1(new_n21628_), .A2(new_n12911_), .B(new_n21629_), .ZN(new_n21630_));
  NAND2_X1   g19194(.A1(new_n21630_), .A2(new_n13392_), .ZN(new_n21631_));
  OAI21_X1   g19195(.A1(new_n13392_), .A2(new_n21563_), .B(new_n21631_), .ZN(new_n21632_));
  NAND2_X1   g19196(.A1(new_n21632_), .A2(new_n12920_), .ZN(new_n21633_));
  NAND2_X1   g19197(.A1(new_n21567_), .A2(pi0628), .ZN(new_n21634_));
  AOI21_X1   g19198(.A1(new_n21633_), .A2(new_n21634_), .B(pi1156), .ZN(new_n21635_));
  NAND2_X1   g19199(.A1(new_n21567_), .A2(new_n12920_), .ZN(new_n21636_));
  NAND2_X1   g19200(.A1(new_n21632_), .A2(pi0628), .ZN(new_n21637_));
  AOI21_X1   g19201(.A1(new_n21637_), .A2(new_n21636_), .B(new_n12742_), .ZN(new_n21638_));
  NOR3_X1    g19202(.A1(new_n21638_), .A2(new_n21635_), .A3(new_n12937_), .ZN(new_n21639_));
  NOR2_X1    g19203(.A1(new_n21632_), .A2(pi0792), .ZN(new_n21640_));
  NOR2_X1    g19204(.A1(new_n21639_), .A2(new_n21640_), .ZN(new_n21641_));
  NAND2_X1   g19205(.A1(new_n21641_), .A2(new_n12741_), .ZN(new_n21642_));
  NAND2_X1   g19206(.A1(new_n21567_), .A2(pi0647), .ZN(new_n21643_));
  AOI21_X1   g19207(.A1(new_n21642_), .A2(new_n21643_), .B(pi1157), .ZN(new_n21644_));
  NAND2_X1   g19208(.A1(new_n21641_), .A2(pi0647), .ZN(new_n21645_));
  OAI21_X1   g19209(.A1(pi0647), .A2(new_n21563_), .B(new_n21645_), .ZN(new_n21646_));
  NAND2_X1   g19210(.A1(new_n21646_), .A2(pi1157), .ZN(new_n21647_));
  NAND2_X1   g19211(.A1(new_n21647_), .A2(pi0787), .ZN(new_n21648_));
  OAI22_X1   g19212(.A1(new_n21648_), .A2(new_n21644_), .B1(pi0787), .B2(new_n21641_), .ZN(new_n21649_));
  AOI21_X1   g19213(.A1(new_n21649_), .A2(pi0644), .B(pi0715), .ZN(new_n21650_));
  NOR2_X1    g19214(.A1(new_n21635_), .A2(new_n12919_), .ZN(new_n21651_));
  AOI21_X1   g19215(.A1(new_n21602_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n21652_));
  AOI21_X1   g19216(.A1(new_n21567_), .A2(new_n12747_), .B(pi0641), .ZN(new_n21653_));
  NAND3_X1   g19217(.A1(new_n21600_), .A2(pi0626), .A3(new_n21593_), .ZN(new_n21654_));
  AOI21_X1   g19218(.A1(new_n21654_), .A2(new_n21653_), .B(new_n12745_), .ZN(new_n21655_));
  AOI21_X1   g19219(.A1(new_n21630_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n21656_));
  NOR3_X1    g19220(.A1(new_n21573_), .A2(new_n21574_), .A3(pi0703), .ZN(new_n21657_));
  OAI21_X1   g19221(.A1(new_n15111_), .A2(pi0186), .B(new_n16803_), .ZN(new_n21658_));
  NOR3_X1    g19222(.A1(new_n15116_), .A2(new_n7381_), .A3(new_n15113_), .ZN(new_n21659_));
  OAI21_X1   g19223(.A1(new_n21659_), .A2(new_n21658_), .B(pi0703), .ZN(new_n21660_));
  OAI21_X1   g19224(.A1(new_n15121_), .A2(new_n7381_), .B(pi0752), .ZN(new_n21661_));
  AOI21_X1   g19225(.A1(new_n15129_), .A2(new_n15126_), .B(pi0186), .ZN(new_n21662_));
  NOR3_X1    g19226(.A1(new_n21662_), .A2(new_n15123_), .A3(new_n21661_), .ZN(new_n21663_));
  OAI21_X1   g19227(.A1(new_n21660_), .A2(new_n21663_), .B(new_n2609_), .ZN(new_n21664_));
  OAI21_X1   g19228(.A1(new_n21664_), .A2(new_n21657_), .B(new_n21569_), .ZN(new_n21665_));
  NAND2_X1   g19229(.A1(new_n21665_), .A2(pi0625), .ZN(new_n21666_));
  NAND2_X1   g19230(.A1(new_n21575_), .A2(new_n21569_), .ZN(new_n21667_));
  NAND2_X1   g19231(.A1(new_n21667_), .A2(new_n13521_), .ZN(new_n21668_));
  AOI21_X1   g19232(.A1(new_n21666_), .A2(new_n21668_), .B(new_n12841_), .ZN(new_n21669_));
  NOR3_X1    g19233(.A1(new_n21669_), .A2(new_n13560_), .A3(new_n21620_), .ZN(new_n21670_));
  AOI21_X1   g19234(.A1(new_n21575_), .A2(new_n21569_), .B(new_n13521_), .ZN(new_n21671_));
  AOI21_X1   g19235(.A1(new_n21665_), .A2(new_n13521_), .B(new_n21671_), .ZN(new_n21672_));
  OAI21_X1   g19236(.A1(new_n21672_), .A2(pi1153), .B(new_n21623_), .ZN(new_n21673_));
  OAI21_X1   g19237(.A1(new_n21673_), .A2(pi0608), .B(pi0778), .ZN(new_n21674_));
  NAND2_X1   g19238(.A1(new_n21665_), .A2(new_n12758_), .ZN(new_n21675_));
  OAI21_X1   g19239(.A1(new_n21674_), .A2(new_n21670_), .B(new_n21675_), .ZN(new_n21676_));
  NAND2_X1   g19240(.A1(new_n21676_), .A2(new_n12764_), .ZN(new_n21677_));
  INV_X1     g19241(.I(new_n21677_), .ZN(new_n21678_));
  AND2_X2    g19242(.A1(new_n21580_), .A2(pi0660), .Z(new_n21679_));
  AOI21_X1   g19243(.A1(new_n21625_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n21680_));
  OAI21_X1   g19244(.A1(new_n21676_), .A2(new_n12766_), .B(new_n21680_), .ZN(new_n21681_));
  NAND2_X1   g19245(.A1(new_n21681_), .A2(new_n21679_), .ZN(new_n21682_));
  NOR2_X1    g19246(.A1(new_n21582_), .A2(pi0660), .ZN(new_n21683_));
  AOI21_X1   g19247(.A1(new_n21625_), .A2(pi0609), .B(pi1155), .ZN(new_n21684_));
  OAI21_X1   g19248(.A1(new_n21676_), .A2(pi0609), .B(new_n21684_), .ZN(new_n21685_));
  AOI21_X1   g19249(.A1(new_n21685_), .A2(new_n21683_), .B(new_n12764_), .ZN(new_n21686_));
  AOI21_X1   g19250(.A1(new_n21686_), .A2(new_n21682_), .B(new_n21678_), .ZN(new_n21687_));
  OR2_X2     g19251(.A1(new_n21687_), .A2(pi0781), .Z(new_n21688_));
  OAI21_X1   g19252(.A1(new_n21586_), .A2(pi1154), .B(pi0627), .ZN(new_n21689_));
  NOR2_X1    g19253(.A1(new_n21626_), .A2(pi0618), .ZN(new_n21690_));
  NOR2_X1    g19254(.A1(new_n21690_), .A2(new_n12785_), .ZN(new_n21691_));
  NAND2_X1   g19255(.A1(new_n21687_), .A2(pi0618), .ZN(new_n21692_));
  AOI21_X1   g19256(.A1(new_n21692_), .A2(new_n21691_), .B(new_n21689_), .ZN(new_n21693_));
  NAND2_X1   g19257(.A1(new_n21590_), .A2(new_n12880_), .ZN(new_n21694_));
  OAI21_X1   g19258(.A1(new_n21626_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n21695_));
  AOI21_X1   g19259(.A1(new_n21687_), .A2(new_n12781_), .B(new_n21695_), .ZN(new_n21696_));
  OAI21_X1   g19260(.A1(new_n21696_), .A2(new_n21694_), .B(pi0781), .ZN(new_n21697_));
  OAI21_X1   g19261(.A1(new_n21697_), .A2(new_n21693_), .B(new_n21688_), .ZN(new_n21698_));
  AND2_X2    g19262(.A1(new_n21698_), .A2(new_n12796_), .Z(new_n21699_));
  AOI21_X1   g19263(.A1(new_n21595_), .A2(new_n12791_), .B(new_n12895_), .ZN(new_n21700_));
  AOI21_X1   g19264(.A1(new_n21628_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n21701_));
  OAI21_X1   g19265(.A1(new_n21698_), .A2(new_n12793_), .B(new_n21701_), .ZN(new_n21702_));
  NAND2_X1   g19266(.A1(new_n21702_), .A2(new_n21700_), .ZN(new_n21703_));
  AOI21_X1   g19267(.A1(new_n21598_), .A2(pi1159), .B(pi0648), .ZN(new_n21704_));
  AOI21_X1   g19268(.A1(new_n21628_), .A2(pi0619), .B(pi1159), .ZN(new_n21705_));
  OAI21_X1   g19269(.A1(new_n21698_), .A2(pi0619), .B(new_n21705_), .ZN(new_n21706_));
  AOI21_X1   g19270(.A1(new_n21706_), .A2(new_n21704_), .B(new_n12796_), .ZN(new_n21707_));
  AOI21_X1   g19271(.A1(new_n21707_), .A2(new_n21703_), .B(new_n21699_), .ZN(new_n21708_));
  OAI21_X1   g19272(.A1(new_n21708_), .A2(new_n12747_), .B(new_n21656_), .ZN(new_n21709_));
  NAND2_X1   g19273(.A1(new_n21709_), .A2(new_n21655_), .ZN(new_n21710_));
  AOI21_X1   g19274(.A1(new_n21567_), .A2(pi0626), .B(new_n12814_), .ZN(new_n21711_));
  NAND3_X1   g19275(.A1(new_n21600_), .A2(new_n12747_), .A3(new_n21593_), .ZN(new_n21712_));
  AOI21_X1   g19276(.A1(new_n21712_), .A2(new_n21711_), .B(pi1158), .ZN(new_n21713_));
  AOI21_X1   g19277(.A1(new_n21630_), .A2(pi0626), .B(pi0641), .ZN(new_n21714_));
  OAI21_X1   g19278(.A1(new_n21708_), .A2(pi0626), .B(new_n21714_), .ZN(new_n21715_));
  AOI21_X1   g19279(.A1(new_n21715_), .A2(new_n21713_), .B(new_n12808_), .ZN(new_n21716_));
  AND2_X2    g19280(.A1(new_n21708_), .A2(new_n12808_), .Z(new_n21717_));
  AOI21_X1   g19281(.A1(new_n21716_), .A2(new_n21710_), .B(new_n21717_), .ZN(new_n21718_));
  OAI21_X1   g19282(.A1(new_n21718_), .A2(new_n12920_), .B(new_n21652_), .ZN(new_n21719_));
  NAND2_X1   g19283(.A1(new_n21719_), .A2(new_n21651_), .ZN(new_n21720_));
  NOR2_X1    g19284(.A1(new_n21638_), .A2(pi0629), .ZN(new_n21721_));
  AOI21_X1   g19285(.A1(new_n21602_), .A2(pi0628), .B(pi1156), .ZN(new_n21722_));
  OAI21_X1   g19286(.A1(new_n21718_), .A2(pi0628), .B(new_n21722_), .ZN(new_n21723_));
  AOI21_X1   g19287(.A1(new_n21723_), .A2(new_n21721_), .B(new_n12937_), .ZN(new_n21724_));
  AND2_X2    g19288(.A1(new_n21718_), .A2(new_n12937_), .Z(new_n21725_));
  AOI21_X1   g19289(.A1(new_n21724_), .A2(new_n21720_), .B(new_n21725_), .ZN(new_n21726_));
  OR2_X2     g19290(.A1(new_n21726_), .A2(pi0787), .Z(new_n21727_));
  OR2_X2     g19291(.A1(new_n21644_), .A2(new_n12981_), .Z(new_n21728_));
  NOR2_X1    g19292(.A1(new_n21603_), .A2(pi0647), .ZN(new_n21729_));
  NOR2_X1    g19293(.A1(new_n21729_), .A2(new_n12965_), .ZN(new_n21730_));
  NAND2_X1   g19294(.A1(new_n21726_), .A2(pi0647), .ZN(new_n21731_));
  AOI21_X1   g19295(.A1(new_n21731_), .A2(new_n21730_), .B(new_n21728_), .ZN(new_n21732_));
  NAND2_X1   g19296(.A1(new_n21647_), .A2(new_n12981_), .ZN(new_n21733_));
  OAI21_X1   g19297(.A1(new_n21603_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n21734_));
  AOI21_X1   g19298(.A1(new_n21726_), .A2(new_n12741_), .B(new_n21734_), .ZN(new_n21735_));
  OAI21_X1   g19299(.A1(new_n21735_), .A2(new_n21733_), .B(pi0787), .ZN(new_n21736_));
  OAI21_X1   g19300(.A1(new_n21736_), .A2(new_n21732_), .B(new_n21727_), .ZN(new_n21737_));
  OAI21_X1   g19301(.A1(new_n21737_), .A2(pi0644), .B(new_n21650_), .ZN(new_n21738_));
  NAND2_X1   g19302(.A1(new_n21738_), .A2(new_n21607_), .ZN(new_n21739_));
  AOI21_X1   g19303(.A1(new_n21563_), .A2(new_n12975_), .B(pi0715), .ZN(new_n21740_));
  NAND2_X1   g19304(.A1(new_n21605_), .A2(pi0644), .ZN(new_n21741_));
  AOI21_X1   g19305(.A1(new_n21741_), .A2(new_n21740_), .B(new_n12739_), .ZN(new_n21742_));
  NOR2_X1    g19306(.A1(new_n21649_), .A2(pi0644), .ZN(new_n21743_));
  AOI21_X1   g19307(.A1(new_n21737_), .A2(pi0644), .B(new_n21743_), .ZN(new_n21744_));
  OAI21_X1   g19308(.A1(new_n21744_), .A2(new_n12740_), .B(new_n21742_), .ZN(new_n21745_));
  NAND3_X1   g19309(.A1(new_n21745_), .A2(new_n21739_), .A3(pi0790), .ZN(new_n21746_));
  AOI21_X1   g19310(.A1(new_n21737_), .A2(new_n13000_), .B(po1038), .ZN(new_n21747_));
  NAND2_X1   g19311(.A1(new_n21746_), .A2(new_n21747_), .ZN(new_n21748_));
  AOI21_X1   g19312(.A1(new_n21748_), .A2(new_n21562_), .B(new_n21561_), .ZN(po0343));
  NOR2_X1    g19313(.A1(new_n3042_), .A2(pi0187), .ZN(new_n21750_));
  INV_X1     g19314(.I(new_n21750_), .ZN(new_n21751_));
  AOI21_X1   g19315(.A1(new_n12756_), .A2(new_n16080_), .B(new_n21750_), .ZN(new_n21752_));
  NOR3_X1    g19316(.A1(new_n21752_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n21753_));
  NOR2_X1    g19317(.A1(new_n21752_), .A2(new_n12762_), .ZN(new_n21754_));
  AOI21_X1   g19318(.A1(new_n21754_), .A2(new_n12768_), .B(pi1155), .ZN(new_n21755_));
  INV_X1     g19319(.I(new_n21752_), .ZN(new_n21756_));
  AOI21_X1   g19320(.A1(new_n21756_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n21757_));
  NOR3_X1    g19321(.A1(new_n21755_), .A2(new_n21757_), .A3(new_n12764_), .ZN(new_n21758_));
  NOR2_X1    g19322(.A1(new_n21758_), .A2(new_n21753_), .ZN(new_n21759_));
  NOR2_X1    g19323(.A1(new_n21759_), .A2(pi0781), .ZN(new_n21760_));
  INV_X1     g19324(.I(new_n21759_), .ZN(new_n21761_));
  AOI21_X1   g19325(.A1(new_n21761_), .A2(new_n12783_), .B(pi1154), .ZN(new_n21762_));
  AOI21_X1   g19326(.A1(new_n21761_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n21763_));
  NOR3_X1    g19327(.A1(new_n21762_), .A2(new_n21763_), .A3(new_n12779_), .ZN(new_n21764_));
  NOR2_X1    g19328(.A1(new_n21764_), .A2(new_n21760_), .ZN(new_n21765_));
  NOR3_X1    g19329(.A1(new_n21764_), .A2(pi0619), .A3(new_n21760_), .ZN(new_n21766_));
  NOR2_X1    g19330(.A1(new_n21750_), .A2(new_n12793_), .ZN(new_n21767_));
  OAI21_X1   g19331(.A1(new_n21766_), .A2(new_n21767_), .B(new_n12791_), .ZN(new_n21768_));
  NAND2_X1   g19332(.A1(new_n21765_), .A2(pi0619), .ZN(new_n21769_));
  NAND2_X1   g19333(.A1(new_n21751_), .A2(new_n12793_), .ZN(new_n21770_));
  AOI21_X1   g19334(.A1(new_n21769_), .A2(new_n21770_), .B(new_n12791_), .ZN(new_n21771_));
  INV_X1     g19335(.I(new_n21771_), .ZN(new_n21772_));
  NAND3_X1   g19336(.A1(new_n21772_), .A2(pi0789), .A3(new_n21768_), .ZN(new_n21773_));
  OAI21_X1   g19337(.A1(pi0789), .A2(new_n21765_), .B(new_n21773_), .ZN(new_n21774_));
  NOR2_X1    g19338(.A1(new_n21774_), .A2(new_n12818_), .ZN(new_n21775_));
  AOI21_X1   g19339(.A1(new_n12818_), .A2(new_n21751_), .B(new_n21775_), .ZN(new_n21776_));
  AOI21_X1   g19340(.A1(new_n12826_), .A2(pi0726), .B(new_n21750_), .ZN(new_n21777_));
  NOR2_X1    g19341(.A1(new_n21777_), .A2(pi0778), .ZN(new_n21778_));
  NOR2_X1    g19342(.A1(new_n12834_), .A2(new_n15993_), .ZN(new_n21779_));
  INV_X1     g19343(.I(new_n21779_), .ZN(new_n21780_));
  NOR2_X1    g19344(.A1(new_n21750_), .A2(pi1153), .ZN(new_n21781_));
  NAND2_X1   g19345(.A1(new_n21780_), .A2(new_n21781_), .ZN(new_n21782_));
  INV_X1     g19346(.I(new_n21782_), .ZN(new_n21783_));
  NOR2_X1    g19347(.A1(new_n21779_), .A2(new_n21777_), .ZN(new_n21784_));
  NOR2_X1    g19348(.A1(new_n21784_), .A2(new_n12841_), .ZN(new_n21785_));
  NOR2_X1    g19349(.A1(new_n21783_), .A2(new_n21785_), .ZN(new_n21786_));
  AOI21_X1   g19350(.A1(new_n21786_), .A2(pi0778), .B(new_n21778_), .ZN(new_n21787_));
  NOR2_X1    g19351(.A1(new_n21787_), .A2(new_n12871_), .ZN(new_n21788_));
  INV_X1     g19352(.I(new_n21788_), .ZN(new_n21789_));
  NOR2_X1    g19353(.A1(new_n21789_), .A2(new_n12889_), .ZN(new_n21790_));
  NAND2_X1   g19354(.A1(new_n21790_), .A2(new_n18203_), .ZN(new_n21791_));
  NOR2_X1    g19355(.A1(new_n21791_), .A2(new_n17884_), .ZN(new_n21792_));
  AOI22_X1   g19356(.A1(new_n21776_), .A2(new_n12949_), .B1(new_n15695_), .B2(new_n21792_), .ZN(new_n21793_));
  NOR2_X1    g19357(.A1(new_n21793_), .A2(pi0629), .ZN(new_n21794_));
  AOI22_X1   g19358(.A1(new_n21776_), .A2(new_n12948_), .B1(new_n15700_), .B2(new_n21792_), .ZN(new_n21795_));
  NOR2_X1    g19359(.A1(new_n21795_), .A2(new_n12919_), .ZN(new_n21796_));
  NOR2_X1    g19360(.A1(new_n21794_), .A2(new_n21796_), .ZN(new_n21797_));
  NOR2_X1    g19361(.A1(new_n21777_), .A2(new_n12754_), .ZN(new_n21798_));
  NOR2_X1    g19362(.A1(new_n21798_), .A2(new_n21756_), .ZN(new_n21799_));
  NAND2_X1   g19363(.A1(new_n21799_), .A2(new_n12758_), .ZN(new_n21800_));
  NAND2_X1   g19364(.A1(new_n21798_), .A2(pi0625), .ZN(new_n21801_));
  NAND3_X1   g19365(.A1(new_n21801_), .A2(pi1153), .A3(new_n21752_), .ZN(new_n21802_));
  AND3_X2    g19366(.A1(new_n21782_), .A2(pi0608), .A3(new_n21802_), .Z(new_n21803_));
  NOR2_X1    g19367(.A1(new_n21785_), .A2(pi0608), .ZN(new_n21804_));
  INV_X1     g19368(.I(new_n21801_), .ZN(new_n21805_));
  OAI21_X1   g19369(.A1(new_n21805_), .A2(new_n21799_), .B(new_n21781_), .ZN(new_n21806_));
  NAND2_X1   g19370(.A1(new_n21804_), .A2(new_n21806_), .ZN(new_n21807_));
  NAND2_X1   g19371(.A1(new_n21807_), .A2(pi0778), .ZN(new_n21808_));
  OAI21_X1   g19372(.A1(new_n21808_), .A2(new_n21803_), .B(new_n21800_), .ZN(new_n21809_));
  INV_X1     g19373(.I(new_n21809_), .ZN(new_n21810_));
  NAND2_X1   g19374(.A1(new_n21787_), .A2(new_n12766_), .ZN(new_n21811_));
  OAI21_X1   g19375(.A1(new_n21810_), .A2(new_n12766_), .B(new_n21811_), .ZN(new_n21812_));
  AOI21_X1   g19376(.A1(new_n21812_), .A2(pi1155), .B(new_n21755_), .ZN(new_n21813_));
  NAND2_X1   g19377(.A1(new_n21809_), .A2(new_n12766_), .ZN(new_n21814_));
  NAND2_X1   g19378(.A1(new_n21787_), .A2(pi0609), .ZN(new_n21815_));
  AOI21_X1   g19379(.A1(new_n21814_), .A2(new_n21815_), .B(pi1155), .ZN(new_n21816_));
  NOR3_X1    g19380(.A1(new_n21816_), .A2(pi0660), .A3(new_n21757_), .ZN(new_n21817_));
  AOI21_X1   g19381(.A1(pi0660), .A2(new_n21813_), .B(new_n21817_), .ZN(new_n21818_));
  NAND2_X1   g19382(.A1(new_n21818_), .A2(pi0785), .ZN(new_n21819_));
  OAI21_X1   g19383(.A1(pi0785), .A2(new_n21810_), .B(new_n21819_), .ZN(new_n21820_));
  INV_X1     g19384(.I(new_n21820_), .ZN(new_n21821_));
  NAND2_X1   g19385(.A1(new_n21789_), .A2(pi0618), .ZN(new_n21822_));
  OAI21_X1   g19386(.A1(new_n21821_), .A2(pi0618), .B(new_n21822_), .ZN(new_n21823_));
  AOI21_X1   g19387(.A1(new_n21823_), .A2(new_n12785_), .B(new_n21763_), .ZN(new_n21824_));
  NOR2_X1    g19388(.A1(new_n21788_), .A2(pi0618), .ZN(new_n21825_));
  NOR2_X1    g19389(.A1(new_n21821_), .A2(new_n12781_), .ZN(new_n21826_));
  OAI21_X1   g19390(.A1(new_n21826_), .A2(new_n21825_), .B(pi1154), .ZN(new_n21827_));
  NOR2_X1    g19391(.A1(new_n21762_), .A2(new_n12880_), .ZN(new_n21828_));
  AOI22_X1   g19392(.A1(new_n21824_), .A2(new_n12880_), .B1(new_n21827_), .B2(new_n21828_), .ZN(new_n21829_));
  NAND2_X1   g19393(.A1(new_n21829_), .A2(pi0781), .ZN(new_n21830_));
  NAND2_X1   g19394(.A1(new_n21820_), .A2(new_n12779_), .ZN(new_n21831_));
  NAND2_X1   g19395(.A1(new_n21830_), .A2(new_n21831_), .ZN(new_n21832_));
  AOI21_X1   g19396(.A1(new_n21832_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n21833_));
  NOR2_X1    g19397(.A1(new_n21790_), .A2(pi0619), .ZN(new_n21834_));
  INV_X1     g19398(.I(new_n21832_), .ZN(new_n21835_));
  NOR2_X1    g19399(.A1(new_n21835_), .A2(new_n12793_), .ZN(new_n21836_));
  OAI21_X1   g19400(.A1(new_n21836_), .A2(new_n21834_), .B(pi1159), .ZN(new_n21837_));
  NAND3_X1   g19401(.A1(new_n21837_), .A2(pi0648), .A3(new_n21768_), .ZN(new_n21838_));
  NOR2_X1    g19402(.A1(new_n21835_), .A2(pi0619), .ZN(new_n21839_));
  NOR2_X1    g19403(.A1(new_n21790_), .A2(new_n12793_), .ZN(new_n21840_));
  OAI21_X1   g19404(.A1(new_n21839_), .A2(new_n21840_), .B(new_n12791_), .ZN(new_n21841_));
  NAND3_X1   g19405(.A1(new_n21841_), .A2(new_n12895_), .A3(new_n21772_), .ZN(new_n21842_));
  NAND3_X1   g19406(.A1(new_n21838_), .A2(new_n21842_), .A3(pi0789), .ZN(new_n21843_));
  NOR2_X1    g19407(.A1(new_n21751_), .A2(new_n12747_), .ZN(new_n21844_));
  INV_X1     g19408(.I(new_n21774_), .ZN(new_n21845_));
  NOR2_X1    g19409(.A1(new_n21845_), .A2(pi0626), .ZN(new_n21846_));
  OAI21_X1   g19410(.A1(new_n21846_), .A2(new_n21844_), .B(new_n12815_), .ZN(new_n21847_));
  INV_X1     g19411(.I(new_n21791_), .ZN(new_n21848_));
  NAND2_X1   g19412(.A1(new_n21750_), .A2(new_n12747_), .ZN(new_n21849_));
  OAI21_X1   g19413(.A1(new_n21845_), .A2(new_n12747_), .B(new_n21849_), .ZN(new_n21850_));
  AOI22_X1   g19414(.A1(new_n21850_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n21848_), .ZN(new_n21851_));
  NAND2_X1   g19415(.A1(new_n21851_), .A2(new_n21847_), .ZN(new_n21852_));
  AOI22_X1   g19416(.A1(new_n21843_), .A2(new_n21833_), .B1(pi0788), .B2(new_n21852_), .ZN(new_n21853_));
  OAI22_X1   g19417(.A1(new_n21853_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n21797_), .ZN(new_n21854_));
  INV_X1     g19418(.I(new_n21776_), .ZN(new_n21855_));
  NAND2_X1   g19419(.A1(new_n21855_), .A2(new_n13384_), .ZN(new_n21856_));
  NAND2_X1   g19420(.A1(new_n12943_), .A2(new_n21751_), .ZN(new_n21857_));
  NAND2_X1   g19421(.A1(new_n21856_), .A2(new_n21857_), .ZN(new_n21858_));
  NAND2_X1   g19422(.A1(new_n21792_), .A2(new_n12954_), .ZN(new_n21859_));
  NAND2_X1   g19423(.A1(new_n21859_), .A2(new_n12741_), .ZN(new_n21860_));
  NOR2_X1    g19424(.A1(new_n21750_), .A2(new_n12741_), .ZN(new_n21861_));
  INV_X1     g19425(.I(new_n21861_), .ZN(new_n21862_));
  AOI21_X1   g19426(.A1(new_n21860_), .A2(new_n21862_), .B(pi1157), .ZN(new_n21863_));
  INV_X1     g19427(.I(new_n21863_), .ZN(new_n21864_));
  NAND2_X1   g19428(.A1(new_n21750_), .A2(new_n12741_), .ZN(new_n21865_));
  OAI21_X1   g19429(.A1(new_n21859_), .A2(new_n12741_), .B(new_n21865_), .ZN(new_n21866_));
  OAI22_X1   g19430(.A1(new_n21864_), .A2(new_n12981_), .B1(new_n21866_), .B2(new_n15576_), .ZN(new_n21867_));
  AOI21_X1   g19431(.A1(new_n21858_), .A2(new_n15608_), .B(new_n21867_), .ZN(new_n21868_));
  OAI22_X1   g19432(.A1(new_n21854_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n21868_), .ZN(new_n21869_));
  NAND2_X1   g19433(.A1(new_n21869_), .A2(new_n13000_), .ZN(new_n21870_));
  AND2_X2    g19434(.A1(new_n21869_), .A2(new_n12975_), .Z(new_n21871_));
  OAI21_X1   g19435(.A1(new_n12965_), .A2(new_n21866_), .B(new_n21864_), .ZN(new_n21872_));
  NAND3_X1   g19436(.A1(new_n21792_), .A2(new_n12972_), .A3(new_n12954_), .ZN(new_n21873_));
  OAI21_X1   g19437(.A1(new_n21872_), .A2(new_n12972_), .B(new_n21873_), .ZN(new_n21874_));
  NOR2_X1    g19438(.A1(new_n21874_), .A2(new_n12975_), .ZN(new_n21875_));
  OAI21_X1   g19439(.A1(new_n21871_), .A2(new_n21875_), .B(new_n12740_), .ZN(new_n21876_));
  NOR2_X1    g19440(.A1(new_n21750_), .A2(new_n12975_), .ZN(new_n21877_));
  NOR2_X1    g19441(.A1(new_n17611_), .A2(new_n21750_), .ZN(new_n21878_));
  AOI21_X1   g19442(.A1(new_n21855_), .A2(new_n17611_), .B(new_n21878_), .ZN(new_n21879_));
  NOR2_X1    g19443(.A1(new_n21879_), .A2(pi0644), .ZN(new_n21880_));
  OAI21_X1   g19444(.A1(new_n21880_), .A2(new_n21877_), .B(pi0715), .ZN(new_n21881_));
  NAND3_X1   g19445(.A1(new_n21876_), .A2(new_n12739_), .A3(new_n21881_), .ZN(new_n21882_));
  NOR2_X1    g19446(.A1(new_n21874_), .A2(pi0644), .ZN(new_n21883_));
  AOI21_X1   g19447(.A1(new_n21869_), .A2(pi0644), .B(new_n21883_), .ZN(new_n21884_));
  NAND2_X1   g19448(.A1(new_n21751_), .A2(new_n12975_), .ZN(new_n21885_));
  OAI21_X1   g19449(.A1(new_n21879_), .A2(new_n12975_), .B(new_n21885_), .ZN(new_n21886_));
  AOI21_X1   g19450(.A1(new_n21886_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n21887_));
  OAI21_X1   g19451(.A1(new_n21884_), .A2(new_n12740_), .B(new_n21887_), .ZN(new_n21888_));
  NAND3_X1   g19452(.A1(new_n21882_), .A2(pi0790), .A3(new_n21888_), .ZN(new_n21889_));
  AOI21_X1   g19453(.A1(new_n21889_), .A2(new_n21870_), .B(new_n12738_), .ZN(new_n21890_));
  AOI21_X1   g19454(.A1(po1038), .A2(new_n9440_), .B(pi0832), .ZN(new_n21891_));
  NOR2_X1    g19455(.A1(new_n13193_), .A2(pi0187), .ZN(new_n21892_));
  AOI21_X1   g19456(.A1(new_n21892_), .A2(pi0644), .B(new_n12740_), .ZN(new_n21893_));
  NOR2_X1    g19457(.A1(new_n21892_), .A2(new_n13384_), .ZN(new_n21894_));
  INV_X1     g19458(.I(new_n21894_), .ZN(new_n21895_));
  INV_X1     g19459(.I(new_n21892_), .ZN(new_n21896_));
  NOR2_X1    g19460(.A1(new_n2609_), .A2(new_n9440_), .ZN(new_n21897_));
  INV_X1     g19461(.I(new_n21897_), .ZN(new_n21898_));
  OAI21_X1   g19462(.A1(new_n15009_), .A2(new_n9440_), .B(new_n18659_), .ZN(new_n21899_));
  NAND2_X1   g19463(.A1(new_n21899_), .A2(new_n16080_), .ZN(new_n21900_));
  NOR2_X1    g19464(.A1(new_n15013_), .A2(pi0770), .ZN(new_n21901_));
  OAI21_X1   g19465(.A1(new_n21901_), .A2(new_n16121_), .B(new_n9440_), .ZN(new_n21902_));
  NAND2_X1   g19466(.A1(new_n21902_), .A2(new_n21900_), .ZN(new_n21903_));
  OAI21_X1   g19467(.A1(new_n21903_), .A2(new_n2610_), .B(new_n21898_), .ZN(new_n21904_));
  INV_X1     g19468(.I(new_n21904_), .ZN(new_n21905_));
  NOR2_X1    g19469(.A1(new_n21905_), .A2(new_n12760_), .ZN(new_n21906_));
  NOR2_X1    g19470(.A1(new_n21892_), .A2(new_n12761_), .ZN(new_n21907_));
  NOR3_X1    g19471(.A1(new_n21906_), .A2(pi0785), .A3(new_n21907_), .ZN(new_n21908_));
  AOI22_X1   g19472(.A1(new_n21906_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n21896_), .ZN(new_n21909_));
  NOR2_X1    g19473(.A1(new_n21909_), .A2(pi1155), .ZN(new_n21910_));
  AOI22_X1   g19474(.A1(new_n21906_), .A2(pi0609), .B1(new_n13357_), .B2(new_n21896_), .ZN(new_n21911_));
  NOR2_X1    g19475(.A1(new_n21911_), .A2(new_n12770_), .ZN(new_n21912_));
  NOR3_X1    g19476(.A1(new_n21910_), .A2(new_n21912_), .A3(new_n12764_), .ZN(new_n21913_));
  NOR2_X1    g19477(.A1(new_n21913_), .A2(new_n21908_), .ZN(new_n21914_));
  NOR2_X1    g19478(.A1(new_n21892_), .A2(new_n12781_), .ZN(new_n21915_));
  AOI21_X1   g19479(.A1(new_n21914_), .A2(new_n12781_), .B(new_n21915_), .ZN(new_n21916_));
  NOR2_X1    g19480(.A1(new_n21916_), .A2(pi1154), .ZN(new_n21917_));
  NOR2_X1    g19481(.A1(new_n21892_), .A2(pi0618), .ZN(new_n21918_));
  AOI21_X1   g19482(.A1(new_n21914_), .A2(pi0618), .B(new_n21918_), .ZN(new_n21919_));
  OAI21_X1   g19483(.A1(new_n21919_), .A2(new_n12785_), .B(pi0781), .ZN(new_n21920_));
  OAI22_X1   g19484(.A1(new_n21920_), .A2(new_n21917_), .B1(pi0781), .B2(new_n21914_), .ZN(new_n21921_));
  NAND2_X1   g19485(.A1(new_n21921_), .A2(new_n12796_), .ZN(new_n21922_));
  NAND2_X1   g19486(.A1(new_n21896_), .A2(pi0619), .ZN(new_n21923_));
  OAI21_X1   g19487(.A1(new_n21921_), .A2(pi0619), .B(new_n21923_), .ZN(new_n21924_));
  NAND2_X1   g19488(.A1(new_n21924_), .A2(new_n12791_), .ZN(new_n21925_));
  NAND2_X1   g19489(.A1(new_n21896_), .A2(new_n12793_), .ZN(new_n21926_));
  OAI21_X1   g19490(.A1(new_n21921_), .A2(new_n12793_), .B(new_n21926_), .ZN(new_n21927_));
  AOI21_X1   g19491(.A1(new_n21927_), .A2(pi1159), .B(new_n12796_), .ZN(new_n21928_));
  NAND2_X1   g19492(.A1(new_n21928_), .A2(new_n21925_), .ZN(new_n21929_));
  AND3_X2    g19493(.A1(new_n21929_), .A2(new_n17504_), .A3(new_n21922_), .Z(new_n21930_));
  AOI21_X1   g19494(.A1(new_n12818_), .A2(new_n21896_), .B(new_n21930_), .ZN(new_n21931_));
  OAI21_X1   g19495(.A1(new_n21931_), .A2(new_n12943_), .B(new_n21895_), .ZN(new_n21932_));
  NAND2_X1   g19496(.A1(new_n21892_), .A2(new_n12984_), .ZN(new_n21933_));
  OAI21_X1   g19497(.A1(new_n21932_), .A2(new_n12984_), .B(new_n21933_), .ZN(new_n21934_));
  NAND2_X1   g19498(.A1(new_n21934_), .A2(new_n12975_), .ZN(new_n21935_));
  AOI21_X1   g19499(.A1(new_n21935_), .A2(new_n21893_), .B(pi1160), .ZN(new_n21936_));
  NOR2_X1    g19500(.A1(new_n21896_), .A2(new_n12870_), .ZN(new_n21937_));
  NAND2_X1   g19501(.A1(new_n9440_), .A2(new_n15993_), .ZN(new_n21938_));
  OAI21_X1   g19502(.A1(new_n13191_), .A2(new_n21938_), .B(new_n2609_), .ZN(new_n21939_));
  NAND2_X1   g19503(.A1(new_n14122_), .A2(pi0187), .ZN(new_n21940_));
  OAI21_X1   g19504(.A1(new_n15744_), .A2(pi0187), .B(new_n21940_), .ZN(new_n21941_));
  NOR2_X1    g19505(.A1(new_n13344_), .A2(pi0187), .ZN(new_n21942_));
  OAI21_X1   g19506(.A1(new_n14125_), .A2(new_n21942_), .B(pi0726), .ZN(new_n21943_));
  AOI21_X1   g19507(.A1(new_n21941_), .A2(new_n3265_), .B(new_n21943_), .ZN(new_n21944_));
  OAI21_X1   g19508(.A1(new_n21944_), .A2(new_n21939_), .B(new_n21898_), .ZN(new_n21945_));
  NAND2_X1   g19509(.A1(new_n21892_), .A2(new_n14133_), .ZN(new_n21946_));
  OAI22_X1   g19510(.A1(new_n14131_), .A2(new_n21945_), .B1(new_n21946_), .B2(new_n12758_), .ZN(new_n21947_));
  AOI21_X1   g19511(.A1(new_n21947_), .A2(new_n12870_), .B(new_n21937_), .ZN(new_n21948_));
  NOR2_X1    g19512(.A1(new_n21892_), .A2(new_n12888_), .ZN(new_n21949_));
  AOI21_X1   g19513(.A1(new_n21948_), .A2(new_n12888_), .B(new_n21949_), .ZN(new_n21950_));
  NOR2_X1    g19514(.A1(new_n21896_), .A2(new_n12911_), .ZN(new_n21951_));
  AOI21_X1   g19515(.A1(new_n21950_), .A2(new_n12911_), .B(new_n21951_), .ZN(new_n21952_));
  NOR2_X1    g19516(.A1(new_n21892_), .A2(new_n13392_), .ZN(new_n21953_));
  AOI21_X1   g19517(.A1(new_n21952_), .A2(new_n13392_), .B(new_n21953_), .ZN(new_n21954_));
  INV_X1     g19518(.I(new_n21954_), .ZN(new_n21955_));
  NAND2_X1   g19519(.A1(new_n21955_), .A2(new_n12920_), .ZN(new_n21956_));
  NAND2_X1   g19520(.A1(new_n21896_), .A2(pi0628), .ZN(new_n21957_));
  AOI21_X1   g19521(.A1(new_n21956_), .A2(new_n21957_), .B(pi1156), .ZN(new_n21958_));
  NAND2_X1   g19522(.A1(new_n21896_), .A2(new_n12920_), .ZN(new_n21959_));
  NAND2_X1   g19523(.A1(new_n21955_), .A2(pi0628), .ZN(new_n21960_));
  AOI21_X1   g19524(.A1(new_n21960_), .A2(new_n21959_), .B(new_n12742_), .ZN(new_n21961_));
  NOR3_X1    g19525(.A1(new_n21961_), .A2(new_n21958_), .A3(new_n12937_), .ZN(new_n21962_));
  AOI21_X1   g19526(.A1(new_n12937_), .A2(new_n21954_), .B(new_n21962_), .ZN(new_n21963_));
  NAND2_X1   g19527(.A1(new_n21963_), .A2(new_n12741_), .ZN(new_n21964_));
  NAND2_X1   g19528(.A1(new_n21896_), .A2(pi0647), .ZN(new_n21965_));
  AOI21_X1   g19529(.A1(new_n21964_), .A2(new_n21965_), .B(pi1157), .ZN(new_n21966_));
  NAND2_X1   g19530(.A1(new_n21963_), .A2(pi0647), .ZN(new_n21967_));
  OAI21_X1   g19531(.A1(pi0647), .A2(new_n21892_), .B(new_n21967_), .ZN(new_n21968_));
  NAND2_X1   g19532(.A1(new_n21968_), .A2(pi1157), .ZN(new_n21969_));
  NAND2_X1   g19533(.A1(new_n21969_), .A2(pi0787), .ZN(new_n21970_));
  OAI22_X1   g19534(.A1(new_n21970_), .A2(new_n21966_), .B1(pi0787), .B2(new_n21963_), .ZN(new_n21971_));
  AOI21_X1   g19535(.A1(new_n21971_), .A2(pi0644), .B(pi0715), .ZN(new_n21972_));
  NOR2_X1    g19536(.A1(new_n21958_), .A2(new_n12919_), .ZN(new_n21973_));
  AOI21_X1   g19537(.A1(new_n21931_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n21974_));
  AOI21_X1   g19538(.A1(new_n21896_), .A2(new_n12747_), .B(pi0641), .ZN(new_n21975_));
  NAND3_X1   g19539(.A1(new_n21929_), .A2(pi0626), .A3(new_n21922_), .ZN(new_n21976_));
  AOI21_X1   g19540(.A1(new_n21976_), .A2(new_n21975_), .B(new_n12745_), .ZN(new_n21977_));
  AOI21_X1   g19541(.A1(new_n21952_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n21978_));
  AOI21_X1   g19542(.A1(new_n14163_), .A2(new_n9440_), .B(pi1153), .ZN(new_n21979_));
  OAI21_X1   g19543(.A1(new_n21945_), .A2(pi0625), .B(new_n21979_), .ZN(new_n21980_));
  NAND2_X1   g19544(.A1(new_n21980_), .A2(pi0608), .ZN(new_n21981_));
  AOI21_X1   g19545(.A1(new_n21905_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n21982_));
  AOI21_X1   g19546(.A1(new_n18437_), .A2(new_n18424_), .B(new_n9440_), .ZN(new_n21983_));
  NOR2_X1    g19547(.A1(new_n19422_), .A2(pi0187), .ZN(new_n21984_));
  OAI21_X1   g19548(.A1(new_n21984_), .A2(new_n21983_), .B(new_n16080_), .ZN(new_n21985_));
  INV_X1     g19549(.I(new_n15121_), .ZN(new_n21986_));
  NAND2_X1   g19550(.A1(new_n21986_), .A2(pi0187), .ZN(new_n21987_));
  NAND2_X1   g19551(.A1(new_n18418_), .A2(new_n9440_), .ZN(new_n21988_));
  NAND4_X1   g19552(.A1(new_n21988_), .A2(pi0770), .A3(new_n18421_), .A4(new_n21987_), .ZN(new_n21989_));
  NAND3_X1   g19553(.A1(new_n21989_), .A2(new_n21985_), .A3(pi0726), .ZN(new_n21990_));
  AOI21_X1   g19554(.A1(new_n21903_), .A2(new_n15993_), .B(new_n2610_), .ZN(new_n21991_));
  AOI21_X1   g19555(.A1(new_n21991_), .A2(new_n21990_), .B(new_n21897_), .ZN(new_n21992_));
  NAND2_X1   g19556(.A1(new_n21992_), .A2(pi0625), .ZN(new_n21993_));
  AOI21_X1   g19557(.A1(new_n21993_), .A2(new_n21982_), .B(new_n21981_), .ZN(new_n21994_));
  AOI21_X1   g19558(.A1(new_n14199_), .A2(new_n9440_), .B(new_n12841_), .ZN(new_n21995_));
  OAI21_X1   g19559(.A1(new_n21945_), .A2(new_n13521_), .B(new_n21995_), .ZN(new_n21996_));
  NAND2_X1   g19560(.A1(new_n21996_), .A2(new_n13560_), .ZN(new_n21997_));
  OAI21_X1   g19561(.A1(new_n21904_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n21998_));
  AOI21_X1   g19562(.A1(new_n21992_), .A2(new_n13521_), .B(new_n21998_), .ZN(new_n21999_));
  OAI21_X1   g19563(.A1(new_n21999_), .A2(new_n21997_), .B(pi0778), .ZN(new_n22000_));
  OR2_X2     g19564(.A1(new_n21992_), .A2(pi0778), .Z(new_n22001_));
  OAI21_X1   g19565(.A1(new_n22000_), .A2(new_n21994_), .B(new_n22001_), .ZN(new_n22002_));
  NAND2_X1   g19566(.A1(new_n22002_), .A2(new_n12764_), .ZN(new_n22003_));
  INV_X1     g19567(.I(new_n22003_), .ZN(new_n22004_));
  NOR2_X1    g19568(.A1(new_n21910_), .A2(new_n13829_), .ZN(new_n22005_));
  NAND2_X1   g19569(.A1(new_n21947_), .A2(new_n12766_), .ZN(new_n22006_));
  NAND2_X1   g19570(.A1(new_n22006_), .A2(pi1155), .ZN(new_n22007_));
  NOR2_X1    g19571(.A1(new_n22002_), .A2(new_n12766_), .ZN(new_n22008_));
  OAI21_X1   g19572(.A1(new_n22008_), .A2(new_n22007_), .B(new_n22005_), .ZN(new_n22009_));
  NOR2_X1    g19573(.A1(new_n21912_), .A2(pi0660), .ZN(new_n22010_));
  AOI21_X1   g19574(.A1(new_n21947_), .A2(pi0609), .B(pi1155), .ZN(new_n22011_));
  OAI21_X1   g19575(.A1(new_n22002_), .A2(pi0609), .B(new_n22011_), .ZN(new_n22012_));
  AOI21_X1   g19576(.A1(new_n22012_), .A2(new_n22010_), .B(new_n12764_), .ZN(new_n22013_));
  AOI21_X1   g19577(.A1(new_n22013_), .A2(new_n22009_), .B(new_n22004_), .ZN(new_n22014_));
  OR2_X2     g19578(.A1(new_n22014_), .A2(pi0781), .Z(new_n22015_));
  OAI21_X1   g19579(.A1(new_n21916_), .A2(pi1154), .B(pi0627), .ZN(new_n22016_));
  INV_X1     g19580(.I(new_n21948_), .ZN(new_n22017_));
  AOI21_X1   g19581(.A1(new_n22017_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n22018_));
  NAND2_X1   g19582(.A1(new_n22014_), .A2(pi0618), .ZN(new_n22019_));
  AOI21_X1   g19583(.A1(new_n22019_), .A2(new_n22018_), .B(new_n22016_), .ZN(new_n22020_));
  OAI21_X1   g19584(.A1(new_n21919_), .A2(new_n12785_), .B(new_n12880_), .ZN(new_n22021_));
  AOI21_X1   g19585(.A1(new_n22017_), .A2(pi0618), .B(pi1154), .ZN(new_n22022_));
  INV_X1     g19586(.I(new_n22022_), .ZN(new_n22023_));
  AOI21_X1   g19587(.A1(new_n22014_), .A2(new_n12781_), .B(new_n22023_), .ZN(new_n22024_));
  OAI21_X1   g19588(.A1(new_n22024_), .A2(new_n22021_), .B(pi0781), .ZN(new_n22025_));
  OAI21_X1   g19589(.A1(new_n22025_), .A2(new_n22020_), .B(new_n22015_), .ZN(new_n22026_));
  AND2_X2    g19590(.A1(new_n22026_), .A2(new_n12796_), .Z(new_n22027_));
  AOI21_X1   g19591(.A1(new_n21950_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n22028_));
  OAI21_X1   g19592(.A1(new_n22026_), .A2(new_n12793_), .B(new_n22028_), .ZN(new_n22029_));
  NAND3_X1   g19593(.A1(new_n22029_), .A2(pi0648), .A3(new_n21925_), .ZN(new_n22030_));
  AOI21_X1   g19594(.A1(new_n21927_), .A2(pi1159), .B(pi0648), .ZN(new_n22031_));
  AOI21_X1   g19595(.A1(new_n21950_), .A2(pi0619), .B(pi1159), .ZN(new_n22032_));
  OAI21_X1   g19596(.A1(new_n22026_), .A2(pi0619), .B(new_n22032_), .ZN(new_n22033_));
  AOI21_X1   g19597(.A1(new_n22033_), .A2(new_n22031_), .B(new_n12796_), .ZN(new_n22034_));
  AOI21_X1   g19598(.A1(new_n22034_), .A2(new_n22030_), .B(new_n22027_), .ZN(new_n22035_));
  OAI21_X1   g19599(.A1(new_n22035_), .A2(new_n12747_), .B(new_n21978_), .ZN(new_n22036_));
  NAND2_X1   g19600(.A1(new_n22036_), .A2(new_n21977_), .ZN(new_n22037_));
  AOI21_X1   g19601(.A1(new_n21896_), .A2(pi0626), .B(new_n12814_), .ZN(new_n22038_));
  NAND3_X1   g19602(.A1(new_n21929_), .A2(new_n12747_), .A3(new_n21922_), .ZN(new_n22039_));
  AOI21_X1   g19603(.A1(new_n22039_), .A2(new_n22038_), .B(pi1158), .ZN(new_n22040_));
  AOI21_X1   g19604(.A1(new_n21952_), .A2(pi0626), .B(pi0641), .ZN(new_n22041_));
  OAI21_X1   g19605(.A1(new_n22035_), .A2(pi0626), .B(new_n22041_), .ZN(new_n22042_));
  AOI21_X1   g19606(.A1(new_n22042_), .A2(new_n22040_), .B(new_n12808_), .ZN(new_n22043_));
  AND2_X2    g19607(.A1(new_n22035_), .A2(new_n12808_), .Z(new_n22044_));
  AOI21_X1   g19608(.A1(new_n22043_), .A2(new_n22037_), .B(new_n22044_), .ZN(new_n22045_));
  OAI21_X1   g19609(.A1(new_n22045_), .A2(new_n12920_), .B(new_n21974_), .ZN(new_n22046_));
  NAND2_X1   g19610(.A1(new_n22046_), .A2(new_n21973_), .ZN(new_n22047_));
  NOR2_X1    g19611(.A1(new_n21961_), .A2(pi0629), .ZN(new_n22048_));
  AOI21_X1   g19612(.A1(new_n21931_), .A2(pi0628), .B(pi1156), .ZN(new_n22049_));
  OAI21_X1   g19613(.A1(new_n22045_), .A2(pi0628), .B(new_n22049_), .ZN(new_n22050_));
  AOI21_X1   g19614(.A1(new_n22050_), .A2(new_n22048_), .B(new_n12937_), .ZN(new_n22051_));
  AND2_X2    g19615(.A1(new_n22045_), .A2(new_n12937_), .Z(new_n22052_));
  AOI21_X1   g19616(.A1(new_n22051_), .A2(new_n22047_), .B(new_n22052_), .ZN(new_n22053_));
  OR2_X2     g19617(.A1(new_n22053_), .A2(pi0787), .Z(new_n22054_));
  OR2_X2     g19618(.A1(new_n21966_), .A2(new_n12981_), .Z(new_n22055_));
  NOR2_X1    g19619(.A1(new_n21932_), .A2(pi0647), .ZN(new_n22056_));
  NOR2_X1    g19620(.A1(new_n22056_), .A2(new_n12965_), .ZN(new_n22057_));
  NAND2_X1   g19621(.A1(new_n22053_), .A2(pi0647), .ZN(new_n22058_));
  AOI21_X1   g19622(.A1(new_n22058_), .A2(new_n22057_), .B(new_n22055_), .ZN(new_n22059_));
  NAND2_X1   g19623(.A1(new_n21969_), .A2(new_n12981_), .ZN(new_n22060_));
  OAI21_X1   g19624(.A1(new_n21932_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n22061_));
  AOI21_X1   g19625(.A1(new_n22053_), .A2(new_n12741_), .B(new_n22061_), .ZN(new_n22062_));
  OAI21_X1   g19626(.A1(new_n22062_), .A2(new_n22060_), .B(pi0787), .ZN(new_n22063_));
  OAI21_X1   g19627(.A1(new_n22063_), .A2(new_n22059_), .B(new_n22054_), .ZN(new_n22064_));
  OAI21_X1   g19628(.A1(new_n22064_), .A2(pi0644), .B(new_n21972_), .ZN(new_n22065_));
  NAND2_X1   g19629(.A1(new_n22065_), .A2(new_n21936_), .ZN(new_n22066_));
  AOI21_X1   g19630(.A1(new_n21892_), .A2(new_n12975_), .B(pi0715), .ZN(new_n22067_));
  NAND2_X1   g19631(.A1(new_n21934_), .A2(pi0644), .ZN(new_n22068_));
  AOI21_X1   g19632(.A1(new_n22068_), .A2(new_n22067_), .B(new_n12739_), .ZN(new_n22069_));
  NOR2_X1    g19633(.A1(new_n21971_), .A2(pi0644), .ZN(new_n22070_));
  AOI21_X1   g19634(.A1(new_n22064_), .A2(pi0644), .B(new_n22070_), .ZN(new_n22071_));
  OAI21_X1   g19635(.A1(new_n22071_), .A2(new_n12740_), .B(new_n22069_), .ZN(new_n22072_));
  NAND3_X1   g19636(.A1(new_n22072_), .A2(new_n22066_), .A3(pi0790), .ZN(new_n22073_));
  AOI21_X1   g19637(.A1(new_n22064_), .A2(new_n13000_), .B(po1038), .ZN(new_n22074_));
  NAND2_X1   g19638(.A1(new_n22073_), .A2(new_n22074_), .ZN(new_n22075_));
  AOI21_X1   g19639(.A1(new_n22075_), .A2(new_n21891_), .B(new_n21890_), .ZN(po0344));
  NOR2_X1    g19640(.A1(new_n3042_), .A2(pi0188), .ZN(new_n22077_));
  INV_X1     g19641(.I(new_n22077_), .ZN(new_n22078_));
  AOI21_X1   g19642(.A1(new_n12756_), .A2(new_n16912_), .B(new_n22077_), .ZN(new_n22079_));
  NOR3_X1    g19643(.A1(new_n22079_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n22080_));
  NOR2_X1    g19644(.A1(new_n22079_), .A2(new_n12762_), .ZN(new_n22081_));
  AOI21_X1   g19645(.A1(new_n22081_), .A2(new_n12768_), .B(pi1155), .ZN(new_n22082_));
  INV_X1     g19646(.I(new_n22079_), .ZN(new_n22083_));
  AOI21_X1   g19647(.A1(new_n22083_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n22084_));
  NOR3_X1    g19648(.A1(new_n22082_), .A2(new_n22084_), .A3(new_n12764_), .ZN(new_n22085_));
  NOR2_X1    g19649(.A1(new_n22085_), .A2(new_n22080_), .ZN(new_n22086_));
  NOR2_X1    g19650(.A1(new_n22086_), .A2(pi0781), .ZN(new_n22087_));
  INV_X1     g19651(.I(new_n22086_), .ZN(new_n22088_));
  AOI21_X1   g19652(.A1(new_n22088_), .A2(new_n12783_), .B(pi1154), .ZN(new_n22089_));
  AOI21_X1   g19653(.A1(new_n22088_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n22090_));
  NOR3_X1    g19654(.A1(new_n22089_), .A2(new_n22090_), .A3(new_n12779_), .ZN(new_n22091_));
  NOR2_X1    g19655(.A1(new_n22091_), .A2(new_n22087_), .ZN(new_n22092_));
  NOR3_X1    g19656(.A1(new_n22091_), .A2(pi0619), .A3(new_n22087_), .ZN(new_n22093_));
  NOR2_X1    g19657(.A1(new_n22077_), .A2(new_n12793_), .ZN(new_n22094_));
  OAI21_X1   g19658(.A1(new_n22093_), .A2(new_n22094_), .B(new_n12791_), .ZN(new_n22095_));
  NAND2_X1   g19659(.A1(new_n22092_), .A2(pi0619), .ZN(new_n22096_));
  NAND2_X1   g19660(.A1(new_n22078_), .A2(new_n12793_), .ZN(new_n22097_));
  AOI21_X1   g19661(.A1(new_n22096_), .A2(new_n22097_), .B(new_n12791_), .ZN(new_n22098_));
  INV_X1     g19662(.I(new_n22098_), .ZN(new_n22099_));
  NAND3_X1   g19663(.A1(new_n22099_), .A2(pi0789), .A3(new_n22095_), .ZN(new_n22100_));
  OAI21_X1   g19664(.A1(pi0789), .A2(new_n22092_), .B(new_n22100_), .ZN(new_n22101_));
  NOR2_X1    g19665(.A1(new_n22101_), .A2(new_n12818_), .ZN(new_n22102_));
  AOI21_X1   g19666(.A1(new_n12818_), .A2(new_n22078_), .B(new_n22102_), .ZN(new_n22103_));
  AOI21_X1   g19667(.A1(new_n12826_), .A2(pi0705), .B(new_n22077_), .ZN(new_n22104_));
  NOR2_X1    g19668(.A1(new_n22104_), .A2(pi0778), .ZN(new_n22105_));
  NOR2_X1    g19669(.A1(new_n12834_), .A2(new_n16906_), .ZN(new_n22106_));
  INV_X1     g19670(.I(new_n22106_), .ZN(new_n22107_));
  NOR2_X1    g19671(.A1(new_n22077_), .A2(pi1153), .ZN(new_n22108_));
  NAND2_X1   g19672(.A1(new_n22107_), .A2(new_n22108_), .ZN(new_n22109_));
  INV_X1     g19673(.I(new_n22109_), .ZN(new_n22110_));
  NOR2_X1    g19674(.A1(new_n22106_), .A2(new_n22104_), .ZN(new_n22111_));
  NOR2_X1    g19675(.A1(new_n22111_), .A2(new_n12841_), .ZN(new_n22112_));
  NOR2_X1    g19676(.A1(new_n22110_), .A2(new_n22112_), .ZN(new_n22113_));
  AOI21_X1   g19677(.A1(new_n22113_), .A2(pi0778), .B(new_n22105_), .ZN(new_n22114_));
  NOR2_X1    g19678(.A1(new_n22114_), .A2(new_n12871_), .ZN(new_n22115_));
  INV_X1     g19679(.I(new_n22115_), .ZN(new_n22116_));
  NOR2_X1    g19680(.A1(new_n22116_), .A2(new_n12889_), .ZN(new_n22117_));
  NAND2_X1   g19681(.A1(new_n22117_), .A2(new_n18203_), .ZN(new_n22118_));
  NOR2_X1    g19682(.A1(new_n22118_), .A2(new_n17884_), .ZN(new_n22119_));
  AOI22_X1   g19683(.A1(new_n22103_), .A2(new_n12949_), .B1(new_n15695_), .B2(new_n22119_), .ZN(new_n22120_));
  NOR2_X1    g19684(.A1(new_n22120_), .A2(pi0629), .ZN(new_n22121_));
  AOI22_X1   g19685(.A1(new_n22103_), .A2(new_n12948_), .B1(new_n15700_), .B2(new_n22119_), .ZN(new_n22122_));
  NOR2_X1    g19686(.A1(new_n22122_), .A2(new_n12919_), .ZN(new_n22123_));
  NOR2_X1    g19687(.A1(new_n22121_), .A2(new_n22123_), .ZN(new_n22124_));
  NOR2_X1    g19688(.A1(new_n22104_), .A2(new_n12754_), .ZN(new_n22125_));
  NOR2_X1    g19689(.A1(new_n22125_), .A2(new_n22083_), .ZN(new_n22126_));
  NAND2_X1   g19690(.A1(new_n22126_), .A2(new_n12758_), .ZN(new_n22127_));
  NAND2_X1   g19691(.A1(new_n22125_), .A2(pi0625), .ZN(new_n22128_));
  NAND3_X1   g19692(.A1(new_n22128_), .A2(pi1153), .A3(new_n22079_), .ZN(new_n22129_));
  AND3_X2    g19693(.A1(new_n22109_), .A2(pi0608), .A3(new_n22129_), .Z(new_n22130_));
  NOR2_X1    g19694(.A1(new_n22112_), .A2(pi0608), .ZN(new_n22131_));
  INV_X1     g19695(.I(new_n22128_), .ZN(new_n22132_));
  OAI21_X1   g19696(.A1(new_n22132_), .A2(new_n22126_), .B(new_n22108_), .ZN(new_n22133_));
  NAND2_X1   g19697(.A1(new_n22131_), .A2(new_n22133_), .ZN(new_n22134_));
  NAND2_X1   g19698(.A1(new_n22134_), .A2(pi0778), .ZN(new_n22135_));
  OAI21_X1   g19699(.A1(new_n22135_), .A2(new_n22130_), .B(new_n22127_), .ZN(new_n22136_));
  INV_X1     g19700(.I(new_n22136_), .ZN(new_n22137_));
  NAND2_X1   g19701(.A1(new_n22114_), .A2(new_n12766_), .ZN(new_n22138_));
  OAI21_X1   g19702(.A1(new_n22137_), .A2(new_n12766_), .B(new_n22138_), .ZN(new_n22139_));
  AOI21_X1   g19703(.A1(new_n22139_), .A2(pi1155), .B(new_n22082_), .ZN(new_n22140_));
  NAND2_X1   g19704(.A1(new_n22136_), .A2(new_n12766_), .ZN(new_n22141_));
  NAND2_X1   g19705(.A1(new_n22114_), .A2(pi0609), .ZN(new_n22142_));
  AOI21_X1   g19706(.A1(new_n22141_), .A2(new_n22142_), .B(pi1155), .ZN(new_n22143_));
  NOR3_X1    g19707(.A1(new_n22143_), .A2(pi0660), .A3(new_n22084_), .ZN(new_n22144_));
  AOI21_X1   g19708(.A1(pi0660), .A2(new_n22140_), .B(new_n22144_), .ZN(new_n22145_));
  NAND2_X1   g19709(.A1(new_n22145_), .A2(pi0785), .ZN(new_n22146_));
  OAI21_X1   g19710(.A1(pi0785), .A2(new_n22137_), .B(new_n22146_), .ZN(new_n22147_));
  INV_X1     g19711(.I(new_n22147_), .ZN(new_n22148_));
  NAND2_X1   g19712(.A1(new_n22116_), .A2(pi0618), .ZN(new_n22149_));
  OAI21_X1   g19713(.A1(new_n22148_), .A2(pi0618), .B(new_n22149_), .ZN(new_n22150_));
  AOI21_X1   g19714(.A1(new_n22150_), .A2(new_n12785_), .B(new_n22090_), .ZN(new_n22151_));
  NOR2_X1    g19715(.A1(new_n22115_), .A2(pi0618), .ZN(new_n22152_));
  NOR2_X1    g19716(.A1(new_n22148_), .A2(new_n12781_), .ZN(new_n22153_));
  OAI21_X1   g19717(.A1(new_n22153_), .A2(new_n22152_), .B(pi1154), .ZN(new_n22154_));
  NOR2_X1    g19718(.A1(new_n22089_), .A2(new_n12880_), .ZN(new_n22155_));
  AOI22_X1   g19719(.A1(new_n22151_), .A2(new_n12880_), .B1(new_n22154_), .B2(new_n22155_), .ZN(new_n22156_));
  NAND2_X1   g19720(.A1(new_n22156_), .A2(pi0781), .ZN(new_n22157_));
  NAND2_X1   g19721(.A1(new_n22147_), .A2(new_n12779_), .ZN(new_n22158_));
  NAND2_X1   g19722(.A1(new_n22157_), .A2(new_n22158_), .ZN(new_n22159_));
  AOI21_X1   g19723(.A1(new_n22159_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n22160_));
  NOR2_X1    g19724(.A1(new_n22117_), .A2(pi0619), .ZN(new_n22161_));
  INV_X1     g19725(.I(new_n22159_), .ZN(new_n22162_));
  NOR2_X1    g19726(.A1(new_n22162_), .A2(new_n12793_), .ZN(new_n22163_));
  OAI21_X1   g19727(.A1(new_n22163_), .A2(new_n22161_), .B(pi1159), .ZN(new_n22164_));
  NAND3_X1   g19728(.A1(new_n22164_), .A2(pi0648), .A3(new_n22095_), .ZN(new_n22165_));
  NOR2_X1    g19729(.A1(new_n22162_), .A2(pi0619), .ZN(new_n22166_));
  NOR2_X1    g19730(.A1(new_n22117_), .A2(new_n12793_), .ZN(new_n22167_));
  OAI21_X1   g19731(.A1(new_n22166_), .A2(new_n22167_), .B(new_n12791_), .ZN(new_n22168_));
  NAND3_X1   g19732(.A1(new_n22168_), .A2(new_n12895_), .A3(new_n22099_), .ZN(new_n22169_));
  NAND3_X1   g19733(.A1(new_n22165_), .A2(new_n22169_), .A3(pi0789), .ZN(new_n22170_));
  NOR2_X1    g19734(.A1(new_n22078_), .A2(new_n12747_), .ZN(new_n22171_));
  INV_X1     g19735(.I(new_n22101_), .ZN(new_n22172_));
  NOR2_X1    g19736(.A1(new_n22172_), .A2(pi0626), .ZN(new_n22173_));
  OAI21_X1   g19737(.A1(new_n22173_), .A2(new_n22171_), .B(new_n12815_), .ZN(new_n22174_));
  INV_X1     g19738(.I(new_n22118_), .ZN(new_n22175_));
  NAND2_X1   g19739(.A1(new_n22077_), .A2(new_n12747_), .ZN(new_n22176_));
  OAI21_X1   g19740(.A1(new_n22172_), .A2(new_n12747_), .B(new_n22176_), .ZN(new_n22177_));
  AOI22_X1   g19741(.A1(new_n22177_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n22175_), .ZN(new_n22178_));
  NAND2_X1   g19742(.A1(new_n22178_), .A2(new_n22174_), .ZN(new_n22179_));
  AOI22_X1   g19743(.A1(new_n22170_), .A2(new_n22160_), .B1(pi0788), .B2(new_n22179_), .ZN(new_n22180_));
  OAI22_X1   g19744(.A1(new_n22180_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n22124_), .ZN(new_n22181_));
  INV_X1     g19745(.I(new_n22103_), .ZN(new_n22182_));
  NAND2_X1   g19746(.A1(new_n22182_), .A2(new_n13384_), .ZN(new_n22183_));
  NAND2_X1   g19747(.A1(new_n12943_), .A2(new_n22078_), .ZN(new_n22184_));
  NAND2_X1   g19748(.A1(new_n22183_), .A2(new_n22184_), .ZN(new_n22185_));
  NAND2_X1   g19749(.A1(new_n22119_), .A2(new_n12954_), .ZN(new_n22186_));
  NAND2_X1   g19750(.A1(new_n22186_), .A2(new_n12741_), .ZN(new_n22187_));
  NOR2_X1    g19751(.A1(new_n22077_), .A2(new_n12741_), .ZN(new_n22188_));
  INV_X1     g19752(.I(new_n22188_), .ZN(new_n22189_));
  AOI21_X1   g19753(.A1(new_n22187_), .A2(new_n22189_), .B(pi1157), .ZN(new_n22190_));
  INV_X1     g19754(.I(new_n22190_), .ZN(new_n22191_));
  NAND2_X1   g19755(.A1(new_n22077_), .A2(new_n12741_), .ZN(new_n22192_));
  OAI21_X1   g19756(.A1(new_n22186_), .A2(new_n12741_), .B(new_n22192_), .ZN(new_n22193_));
  OAI22_X1   g19757(.A1(new_n22191_), .A2(new_n12981_), .B1(new_n22193_), .B2(new_n15576_), .ZN(new_n22194_));
  AOI21_X1   g19758(.A1(new_n22185_), .A2(new_n15608_), .B(new_n22194_), .ZN(new_n22195_));
  OAI22_X1   g19759(.A1(new_n22181_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n22195_), .ZN(new_n22196_));
  NAND2_X1   g19760(.A1(new_n22196_), .A2(new_n13000_), .ZN(new_n22197_));
  AND2_X2    g19761(.A1(new_n22196_), .A2(new_n12975_), .Z(new_n22198_));
  OAI21_X1   g19762(.A1(new_n12965_), .A2(new_n22193_), .B(new_n22191_), .ZN(new_n22199_));
  NAND3_X1   g19763(.A1(new_n22119_), .A2(new_n12972_), .A3(new_n12954_), .ZN(new_n22200_));
  OAI21_X1   g19764(.A1(new_n22199_), .A2(new_n12972_), .B(new_n22200_), .ZN(new_n22201_));
  NOR2_X1    g19765(.A1(new_n22201_), .A2(new_n12975_), .ZN(new_n22202_));
  OAI21_X1   g19766(.A1(new_n22198_), .A2(new_n22202_), .B(new_n12740_), .ZN(new_n22203_));
  NOR2_X1    g19767(.A1(new_n22077_), .A2(new_n12975_), .ZN(new_n22204_));
  NOR2_X1    g19768(.A1(new_n17611_), .A2(new_n22077_), .ZN(new_n22205_));
  AOI21_X1   g19769(.A1(new_n22182_), .A2(new_n17611_), .B(new_n22205_), .ZN(new_n22206_));
  NOR2_X1    g19770(.A1(new_n22206_), .A2(pi0644), .ZN(new_n22207_));
  OAI21_X1   g19771(.A1(new_n22207_), .A2(new_n22204_), .B(pi0715), .ZN(new_n22208_));
  NAND3_X1   g19772(.A1(new_n22203_), .A2(new_n12739_), .A3(new_n22208_), .ZN(new_n22209_));
  NOR2_X1    g19773(.A1(new_n22201_), .A2(pi0644), .ZN(new_n22210_));
  AOI21_X1   g19774(.A1(new_n22196_), .A2(pi0644), .B(new_n22210_), .ZN(new_n22211_));
  NAND2_X1   g19775(.A1(new_n22078_), .A2(new_n12975_), .ZN(new_n22212_));
  OAI21_X1   g19776(.A1(new_n22206_), .A2(new_n12975_), .B(new_n22212_), .ZN(new_n22213_));
  AOI21_X1   g19777(.A1(new_n22213_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n22214_));
  OAI21_X1   g19778(.A1(new_n22211_), .A2(new_n12740_), .B(new_n22214_), .ZN(new_n22215_));
  NAND3_X1   g19779(.A1(new_n22209_), .A2(pi0790), .A3(new_n22215_), .ZN(new_n22216_));
  AOI21_X1   g19780(.A1(new_n22216_), .A2(new_n22197_), .B(new_n12738_), .ZN(new_n22217_));
  AOI21_X1   g19781(.A1(po1038), .A2(new_n7958_), .B(pi0832), .ZN(new_n22218_));
  NOR2_X1    g19782(.A1(new_n13193_), .A2(pi0188), .ZN(new_n22219_));
  AOI21_X1   g19783(.A1(new_n22219_), .A2(pi0644), .B(new_n12740_), .ZN(new_n22220_));
  NOR2_X1    g19784(.A1(new_n22219_), .A2(new_n13384_), .ZN(new_n22221_));
  INV_X1     g19785(.I(new_n22221_), .ZN(new_n22222_));
  INV_X1     g19786(.I(new_n22219_), .ZN(new_n22223_));
  NOR2_X1    g19787(.A1(new_n2609_), .A2(new_n7958_), .ZN(new_n22224_));
  INV_X1     g19788(.I(new_n22224_), .ZN(new_n22225_));
  OAI21_X1   g19789(.A1(new_n15009_), .A2(new_n7958_), .B(new_n18659_), .ZN(new_n22226_));
  NAND2_X1   g19790(.A1(new_n22226_), .A2(new_n16912_), .ZN(new_n22227_));
  NOR2_X1    g19791(.A1(new_n15013_), .A2(pi0768), .ZN(new_n22228_));
  OAI21_X1   g19792(.A1(new_n22228_), .A2(new_n16922_), .B(new_n7958_), .ZN(new_n22229_));
  NAND2_X1   g19793(.A1(new_n22229_), .A2(new_n22227_), .ZN(new_n22230_));
  OAI21_X1   g19794(.A1(new_n22230_), .A2(new_n2610_), .B(new_n22225_), .ZN(new_n22231_));
  INV_X1     g19795(.I(new_n22231_), .ZN(new_n22232_));
  NOR2_X1    g19796(.A1(new_n22232_), .A2(new_n12760_), .ZN(new_n22233_));
  NOR2_X1    g19797(.A1(new_n22219_), .A2(new_n12761_), .ZN(new_n22234_));
  NOR3_X1    g19798(.A1(new_n22233_), .A2(pi0785), .A3(new_n22234_), .ZN(new_n22235_));
  AOI22_X1   g19799(.A1(new_n22233_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n22223_), .ZN(new_n22236_));
  NOR2_X1    g19800(.A1(new_n22236_), .A2(pi1155), .ZN(new_n22237_));
  AOI22_X1   g19801(.A1(new_n22233_), .A2(pi0609), .B1(new_n13357_), .B2(new_n22223_), .ZN(new_n22238_));
  NOR2_X1    g19802(.A1(new_n22238_), .A2(new_n12770_), .ZN(new_n22239_));
  NOR3_X1    g19803(.A1(new_n22237_), .A2(new_n22239_), .A3(new_n12764_), .ZN(new_n22240_));
  NOR2_X1    g19804(.A1(new_n22240_), .A2(new_n22235_), .ZN(new_n22241_));
  NOR2_X1    g19805(.A1(new_n22219_), .A2(new_n12781_), .ZN(new_n22242_));
  AOI21_X1   g19806(.A1(new_n22241_), .A2(new_n12781_), .B(new_n22242_), .ZN(new_n22243_));
  NOR2_X1    g19807(.A1(new_n22243_), .A2(pi1154), .ZN(new_n22244_));
  NOR2_X1    g19808(.A1(new_n22219_), .A2(pi0618), .ZN(new_n22245_));
  AOI21_X1   g19809(.A1(new_n22241_), .A2(pi0618), .B(new_n22245_), .ZN(new_n22246_));
  OAI21_X1   g19810(.A1(new_n22246_), .A2(new_n12785_), .B(pi0781), .ZN(new_n22247_));
  OAI22_X1   g19811(.A1(new_n22247_), .A2(new_n22244_), .B1(pi0781), .B2(new_n22241_), .ZN(new_n22248_));
  NAND2_X1   g19812(.A1(new_n22248_), .A2(new_n12796_), .ZN(new_n22249_));
  NAND2_X1   g19813(.A1(new_n22223_), .A2(pi0619), .ZN(new_n22250_));
  OAI21_X1   g19814(.A1(new_n22248_), .A2(pi0619), .B(new_n22250_), .ZN(new_n22251_));
  NAND2_X1   g19815(.A1(new_n22251_), .A2(new_n12791_), .ZN(new_n22252_));
  NAND2_X1   g19816(.A1(new_n22223_), .A2(new_n12793_), .ZN(new_n22253_));
  OAI21_X1   g19817(.A1(new_n22248_), .A2(new_n12793_), .B(new_n22253_), .ZN(new_n22254_));
  AOI21_X1   g19818(.A1(new_n22254_), .A2(pi1159), .B(new_n12796_), .ZN(new_n22255_));
  NAND2_X1   g19819(.A1(new_n22255_), .A2(new_n22252_), .ZN(new_n22256_));
  AND3_X2    g19820(.A1(new_n22256_), .A2(new_n17504_), .A3(new_n22249_), .Z(new_n22257_));
  AOI21_X1   g19821(.A1(new_n12818_), .A2(new_n22223_), .B(new_n22257_), .ZN(new_n22258_));
  OAI21_X1   g19822(.A1(new_n22258_), .A2(new_n12943_), .B(new_n22222_), .ZN(new_n22259_));
  NAND2_X1   g19823(.A1(new_n22219_), .A2(new_n12984_), .ZN(new_n22260_));
  OAI21_X1   g19824(.A1(new_n22259_), .A2(new_n12984_), .B(new_n22260_), .ZN(new_n22261_));
  NAND2_X1   g19825(.A1(new_n22261_), .A2(new_n12975_), .ZN(new_n22262_));
  AOI21_X1   g19826(.A1(new_n22262_), .A2(new_n22220_), .B(pi1160), .ZN(new_n22263_));
  NOR2_X1    g19827(.A1(new_n22223_), .A2(new_n12870_), .ZN(new_n22264_));
  NAND2_X1   g19828(.A1(new_n7958_), .A2(new_n16906_), .ZN(new_n22265_));
  OAI21_X1   g19829(.A1(new_n13191_), .A2(new_n22265_), .B(new_n2609_), .ZN(new_n22266_));
  NAND2_X1   g19830(.A1(new_n14122_), .A2(pi0188), .ZN(new_n22267_));
  OAI21_X1   g19831(.A1(new_n15744_), .A2(pi0188), .B(new_n22267_), .ZN(new_n22268_));
  NOR2_X1    g19832(.A1(new_n13344_), .A2(pi0188), .ZN(new_n22269_));
  OAI21_X1   g19833(.A1(new_n14125_), .A2(new_n22269_), .B(pi0705), .ZN(new_n22270_));
  AOI21_X1   g19834(.A1(new_n22268_), .A2(new_n3265_), .B(new_n22270_), .ZN(new_n22271_));
  OAI21_X1   g19835(.A1(new_n22271_), .A2(new_n22266_), .B(new_n22225_), .ZN(new_n22272_));
  NAND2_X1   g19836(.A1(new_n22219_), .A2(new_n14133_), .ZN(new_n22273_));
  OAI22_X1   g19837(.A1(new_n14131_), .A2(new_n22272_), .B1(new_n22273_), .B2(new_n12758_), .ZN(new_n22274_));
  AOI21_X1   g19838(.A1(new_n22274_), .A2(new_n12870_), .B(new_n22264_), .ZN(new_n22275_));
  NOR2_X1    g19839(.A1(new_n22219_), .A2(new_n12888_), .ZN(new_n22276_));
  AOI21_X1   g19840(.A1(new_n22275_), .A2(new_n12888_), .B(new_n22276_), .ZN(new_n22277_));
  NOR2_X1    g19841(.A1(new_n22223_), .A2(new_n12911_), .ZN(new_n22278_));
  AOI21_X1   g19842(.A1(new_n22277_), .A2(new_n12911_), .B(new_n22278_), .ZN(new_n22279_));
  NOR2_X1    g19843(.A1(new_n22219_), .A2(new_n13392_), .ZN(new_n22280_));
  AOI21_X1   g19844(.A1(new_n22279_), .A2(new_n13392_), .B(new_n22280_), .ZN(new_n22281_));
  INV_X1     g19845(.I(new_n22281_), .ZN(new_n22282_));
  NAND2_X1   g19846(.A1(new_n22282_), .A2(new_n12920_), .ZN(new_n22283_));
  NAND2_X1   g19847(.A1(new_n22223_), .A2(pi0628), .ZN(new_n22284_));
  AOI21_X1   g19848(.A1(new_n22283_), .A2(new_n22284_), .B(pi1156), .ZN(new_n22285_));
  NAND2_X1   g19849(.A1(new_n22223_), .A2(new_n12920_), .ZN(new_n22286_));
  NAND2_X1   g19850(.A1(new_n22282_), .A2(pi0628), .ZN(new_n22287_));
  AOI21_X1   g19851(.A1(new_n22287_), .A2(new_n22286_), .B(new_n12742_), .ZN(new_n22288_));
  NOR3_X1    g19852(.A1(new_n22288_), .A2(new_n22285_), .A3(new_n12937_), .ZN(new_n22289_));
  AOI21_X1   g19853(.A1(new_n12937_), .A2(new_n22281_), .B(new_n22289_), .ZN(new_n22290_));
  NAND2_X1   g19854(.A1(new_n22290_), .A2(new_n12741_), .ZN(new_n22291_));
  NAND2_X1   g19855(.A1(new_n22223_), .A2(pi0647), .ZN(new_n22292_));
  AOI21_X1   g19856(.A1(new_n22291_), .A2(new_n22292_), .B(pi1157), .ZN(new_n22293_));
  NAND2_X1   g19857(.A1(new_n22290_), .A2(pi0647), .ZN(new_n22294_));
  OAI21_X1   g19858(.A1(pi0647), .A2(new_n22219_), .B(new_n22294_), .ZN(new_n22295_));
  NAND2_X1   g19859(.A1(new_n22295_), .A2(pi1157), .ZN(new_n22296_));
  NAND2_X1   g19860(.A1(new_n22296_), .A2(pi0787), .ZN(new_n22297_));
  OAI22_X1   g19861(.A1(new_n22297_), .A2(new_n22293_), .B1(pi0787), .B2(new_n22290_), .ZN(new_n22298_));
  AOI21_X1   g19862(.A1(new_n22298_), .A2(pi0644), .B(pi0715), .ZN(new_n22299_));
  NOR2_X1    g19863(.A1(new_n22285_), .A2(new_n12919_), .ZN(new_n22300_));
  AOI21_X1   g19864(.A1(new_n22258_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n22301_));
  AOI21_X1   g19865(.A1(new_n22223_), .A2(new_n12747_), .B(pi0641), .ZN(new_n22302_));
  NAND3_X1   g19866(.A1(new_n22256_), .A2(pi0626), .A3(new_n22249_), .ZN(new_n22303_));
  AOI21_X1   g19867(.A1(new_n22303_), .A2(new_n22302_), .B(new_n12745_), .ZN(new_n22304_));
  AOI21_X1   g19868(.A1(new_n22279_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n22305_));
  AOI21_X1   g19869(.A1(new_n14163_), .A2(new_n7958_), .B(pi1153), .ZN(new_n22306_));
  OAI21_X1   g19870(.A1(new_n22272_), .A2(pi0625), .B(new_n22306_), .ZN(new_n22307_));
  NAND2_X1   g19871(.A1(new_n22307_), .A2(pi0608), .ZN(new_n22308_));
  AOI21_X1   g19872(.A1(new_n22232_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n22309_));
  AOI21_X1   g19873(.A1(new_n18437_), .A2(new_n18424_), .B(new_n7958_), .ZN(new_n22310_));
  NOR2_X1    g19874(.A1(new_n19422_), .A2(pi0188), .ZN(new_n22311_));
  OAI21_X1   g19875(.A1(new_n22311_), .A2(new_n22310_), .B(new_n16912_), .ZN(new_n22312_));
  NAND2_X1   g19876(.A1(new_n21986_), .A2(pi0188), .ZN(new_n22313_));
  NAND2_X1   g19877(.A1(new_n18418_), .A2(new_n7958_), .ZN(new_n22314_));
  NAND4_X1   g19878(.A1(new_n22314_), .A2(pi0768), .A3(new_n18421_), .A4(new_n22313_), .ZN(new_n22315_));
  NAND3_X1   g19879(.A1(new_n22315_), .A2(new_n22312_), .A3(pi0705), .ZN(new_n22316_));
  AOI21_X1   g19880(.A1(new_n22230_), .A2(new_n16906_), .B(new_n2610_), .ZN(new_n22317_));
  AOI21_X1   g19881(.A1(new_n22317_), .A2(new_n22316_), .B(new_n22224_), .ZN(new_n22318_));
  NAND2_X1   g19882(.A1(new_n22318_), .A2(pi0625), .ZN(new_n22319_));
  AOI21_X1   g19883(.A1(new_n22319_), .A2(new_n22309_), .B(new_n22308_), .ZN(new_n22320_));
  AOI21_X1   g19884(.A1(new_n14199_), .A2(new_n7958_), .B(new_n12841_), .ZN(new_n22321_));
  OAI21_X1   g19885(.A1(new_n22272_), .A2(new_n13521_), .B(new_n22321_), .ZN(new_n22322_));
  NAND2_X1   g19886(.A1(new_n22322_), .A2(new_n13560_), .ZN(new_n22323_));
  OAI21_X1   g19887(.A1(new_n22231_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n22324_));
  AOI21_X1   g19888(.A1(new_n22318_), .A2(new_n13521_), .B(new_n22324_), .ZN(new_n22325_));
  OAI21_X1   g19889(.A1(new_n22325_), .A2(new_n22323_), .B(pi0778), .ZN(new_n22326_));
  OR2_X2     g19890(.A1(new_n22318_), .A2(pi0778), .Z(new_n22327_));
  OAI21_X1   g19891(.A1(new_n22326_), .A2(new_n22320_), .B(new_n22327_), .ZN(new_n22328_));
  NAND2_X1   g19892(.A1(new_n22328_), .A2(new_n12764_), .ZN(new_n22329_));
  INV_X1     g19893(.I(new_n22329_), .ZN(new_n22330_));
  NOR2_X1    g19894(.A1(new_n22237_), .A2(new_n13829_), .ZN(new_n22331_));
  NAND2_X1   g19895(.A1(new_n22274_), .A2(new_n12766_), .ZN(new_n22332_));
  NAND2_X1   g19896(.A1(new_n22332_), .A2(pi1155), .ZN(new_n22333_));
  NOR2_X1    g19897(.A1(new_n22328_), .A2(new_n12766_), .ZN(new_n22334_));
  OAI21_X1   g19898(.A1(new_n22334_), .A2(new_n22333_), .B(new_n22331_), .ZN(new_n22335_));
  NOR2_X1    g19899(.A1(new_n22239_), .A2(pi0660), .ZN(new_n22336_));
  AOI21_X1   g19900(.A1(new_n22274_), .A2(pi0609), .B(pi1155), .ZN(new_n22337_));
  OAI21_X1   g19901(.A1(new_n22328_), .A2(pi0609), .B(new_n22337_), .ZN(new_n22338_));
  AOI21_X1   g19902(.A1(new_n22338_), .A2(new_n22336_), .B(new_n12764_), .ZN(new_n22339_));
  AOI21_X1   g19903(.A1(new_n22339_), .A2(new_n22335_), .B(new_n22330_), .ZN(new_n22340_));
  OR2_X2     g19904(.A1(new_n22340_), .A2(pi0781), .Z(new_n22341_));
  OAI21_X1   g19905(.A1(new_n22243_), .A2(pi1154), .B(pi0627), .ZN(new_n22342_));
  INV_X1     g19906(.I(new_n22275_), .ZN(new_n22343_));
  AOI21_X1   g19907(.A1(new_n22343_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n22344_));
  NAND2_X1   g19908(.A1(new_n22340_), .A2(pi0618), .ZN(new_n22345_));
  AOI21_X1   g19909(.A1(new_n22345_), .A2(new_n22344_), .B(new_n22342_), .ZN(new_n22346_));
  OAI21_X1   g19910(.A1(new_n22246_), .A2(new_n12785_), .B(new_n12880_), .ZN(new_n22347_));
  AOI21_X1   g19911(.A1(new_n22343_), .A2(pi0618), .B(pi1154), .ZN(new_n22348_));
  INV_X1     g19912(.I(new_n22348_), .ZN(new_n22349_));
  AOI21_X1   g19913(.A1(new_n22340_), .A2(new_n12781_), .B(new_n22349_), .ZN(new_n22350_));
  OAI21_X1   g19914(.A1(new_n22350_), .A2(new_n22347_), .B(pi0781), .ZN(new_n22351_));
  OAI21_X1   g19915(.A1(new_n22351_), .A2(new_n22346_), .B(new_n22341_), .ZN(new_n22352_));
  AND2_X2    g19916(.A1(new_n22352_), .A2(new_n12796_), .Z(new_n22353_));
  AOI21_X1   g19917(.A1(new_n22277_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n22354_));
  OAI21_X1   g19918(.A1(new_n22352_), .A2(new_n12793_), .B(new_n22354_), .ZN(new_n22355_));
  NAND3_X1   g19919(.A1(new_n22355_), .A2(pi0648), .A3(new_n22252_), .ZN(new_n22356_));
  AOI21_X1   g19920(.A1(new_n22254_), .A2(pi1159), .B(pi0648), .ZN(new_n22357_));
  AOI21_X1   g19921(.A1(new_n22277_), .A2(pi0619), .B(pi1159), .ZN(new_n22358_));
  OAI21_X1   g19922(.A1(new_n22352_), .A2(pi0619), .B(new_n22358_), .ZN(new_n22359_));
  AOI21_X1   g19923(.A1(new_n22359_), .A2(new_n22357_), .B(new_n12796_), .ZN(new_n22360_));
  AOI21_X1   g19924(.A1(new_n22360_), .A2(new_n22356_), .B(new_n22353_), .ZN(new_n22361_));
  OAI21_X1   g19925(.A1(new_n22361_), .A2(new_n12747_), .B(new_n22305_), .ZN(new_n22362_));
  NAND2_X1   g19926(.A1(new_n22362_), .A2(new_n22304_), .ZN(new_n22363_));
  AOI21_X1   g19927(.A1(new_n22223_), .A2(pi0626), .B(new_n12814_), .ZN(new_n22364_));
  NAND3_X1   g19928(.A1(new_n22256_), .A2(new_n12747_), .A3(new_n22249_), .ZN(new_n22365_));
  AOI21_X1   g19929(.A1(new_n22365_), .A2(new_n22364_), .B(pi1158), .ZN(new_n22366_));
  AOI21_X1   g19930(.A1(new_n22279_), .A2(pi0626), .B(pi0641), .ZN(new_n22367_));
  OAI21_X1   g19931(.A1(new_n22361_), .A2(pi0626), .B(new_n22367_), .ZN(new_n22368_));
  AOI21_X1   g19932(.A1(new_n22368_), .A2(new_n22366_), .B(new_n12808_), .ZN(new_n22369_));
  AND2_X2    g19933(.A1(new_n22361_), .A2(new_n12808_), .Z(new_n22370_));
  AOI21_X1   g19934(.A1(new_n22369_), .A2(new_n22363_), .B(new_n22370_), .ZN(new_n22371_));
  OAI21_X1   g19935(.A1(new_n22371_), .A2(new_n12920_), .B(new_n22301_), .ZN(new_n22372_));
  NAND2_X1   g19936(.A1(new_n22372_), .A2(new_n22300_), .ZN(new_n22373_));
  NOR2_X1    g19937(.A1(new_n22288_), .A2(pi0629), .ZN(new_n22374_));
  AOI21_X1   g19938(.A1(new_n22258_), .A2(pi0628), .B(pi1156), .ZN(new_n22375_));
  OAI21_X1   g19939(.A1(new_n22371_), .A2(pi0628), .B(new_n22375_), .ZN(new_n22376_));
  AOI21_X1   g19940(.A1(new_n22376_), .A2(new_n22374_), .B(new_n12937_), .ZN(new_n22377_));
  AND2_X2    g19941(.A1(new_n22371_), .A2(new_n12937_), .Z(new_n22378_));
  AOI21_X1   g19942(.A1(new_n22377_), .A2(new_n22373_), .B(new_n22378_), .ZN(new_n22379_));
  OR2_X2     g19943(.A1(new_n22379_), .A2(pi0787), .Z(new_n22380_));
  OR2_X2     g19944(.A1(new_n22293_), .A2(new_n12981_), .Z(new_n22381_));
  NOR2_X1    g19945(.A1(new_n22259_), .A2(pi0647), .ZN(new_n22382_));
  NOR2_X1    g19946(.A1(new_n22382_), .A2(new_n12965_), .ZN(new_n22383_));
  NAND2_X1   g19947(.A1(new_n22379_), .A2(pi0647), .ZN(new_n22384_));
  AOI21_X1   g19948(.A1(new_n22384_), .A2(new_n22383_), .B(new_n22381_), .ZN(new_n22385_));
  NAND2_X1   g19949(.A1(new_n22296_), .A2(new_n12981_), .ZN(new_n22386_));
  OAI21_X1   g19950(.A1(new_n22259_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n22387_));
  AOI21_X1   g19951(.A1(new_n22379_), .A2(new_n12741_), .B(new_n22387_), .ZN(new_n22388_));
  OAI21_X1   g19952(.A1(new_n22388_), .A2(new_n22386_), .B(pi0787), .ZN(new_n22389_));
  OAI21_X1   g19953(.A1(new_n22389_), .A2(new_n22385_), .B(new_n22380_), .ZN(new_n22390_));
  OAI21_X1   g19954(.A1(new_n22390_), .A2(pi0644), .B(new_n22299_), .ZN(new_n22391_));
  NAND2_X1   g19955(.A1(new_n22391_), .A2(new_n22263_), .ZN(new_n22392_));
  AOI21_X1   g19956(.A1(new_n22219_), .A2(new_n12975_), .B(pi0715), .ZN(new_n22393_));
  NAND2_X1   g19957(.A1(new_n22261_), .A2(pi0644), .ZN(new_n22394_));
  AOI21_X1   g19958(.A1(new_n22394_), .A2(new_n22393_), .B(new_n12739_), .ZN(new_n22395_));
  NOR2_X1    g19959(.A1(new_n22298_), .A2(pi0644), .ZN(new_n22396_));
  AOI21_X1   g19960(.A1(new_n22390_), .A2(pi0644), .B(new_n22396_), .ZN(new_n22397_));
  OAI21_X1   g19961(.A1(new_n22397_), .A2(new_n12740_), .B(new_n22395_), .ZN(new_n22398_));
  NAND3_X1   g19962(.A1(new_n22398_), .A2(new_n22392_), .A3(pi0790), .ZN(new_n22399_));
  AOI21_X1   g19963(.A1(new_n22390_), .A2(new_n13000_), .B(po1038), .ZN(new_n22400_));
  NAND2_X1   g19964(.A1(new_n22399_), .A2(new_n22400_), .ZN(new_n22401_));
  AOI21_X1   g19965(.A1(new_n22401_), .A2(new_n22218_), .B(new_n22217_), .ZN(po0345));
  NOR2_X1    g19966(.A1(new_n3042_), .A2(new_n9484_), .ZN(new_n22403_));
  NOR2_X1    g19967(.A1(new_n13340_), .A2(new_n16845_), .ZN(new_n22404_));
  INV_X1     g19968(.I(new_n22404_), .ZN(new_n22405_));
  NOR2_X1    g19969(.A1(new_n22405_), .A2(new_n15232_), .ZN(new_n22406_));
  INV_X1     g19970(.I(new_n22406_), .ZN(new_n22407_));
  NOR2_X1    g19971(.A1(new_n22407_), .A2(new_n15246_), .ZN(new_n22408_));
  INV_X1     g19972(.I(new_n22408_), .ZN(new_n22409_));
  NOR2_X1    g19973(.A1(new_n22409_), .A2(new_n12818_), .ZN(new_n22410_));
  INV_X1     g19974(.I(new_n22410_), .ZN(new_n22411_));
  NOR3_X1    g19975(.A1(new_n22411_), .A2(new_n12981_), .A3(new_n12943_), .ZN(new_n22412_));
  INV_X1     g19976(.I(new_n22403_), .ZN(new_n22413_));
  NAND2_X1   g19977(.A1(new_n12826_), .A2(pi0727), .ZN(new_n22414_));
  NAND2_X1   g19978(.A1(new_n22414_), .A2(new_n22413_), .ZN(new_n22415_));
  INV_X1     g19979(.I(new_n22415_), .ZN(new_n22416_));
  NOR2_X1    g19980(.A1(new_n22414_), .A2(new_n13521_), .ZN(new_n22417_));
  NOR3_X1    g19981(.A1(new_n22417_), .A2(new_n12841_), .A3(new_n22403_), .ZN(new_n22418_));
  INV_X1     g19982(.I(new_n22418_), .ZN(new_n22419_));
  OAI21_X1   g19983(.A1(new_n22416_), .A2(new_n22417_), .B(new_n12841_), .ZN(new_n22420_));
  NAND3_X1   g19984(.A1(new_n22419_), .A2(new_n22420_), .A3(pi0778), .ZN(new_n22421_));
  OAI21_X1   g19985(.A1(pi0778), .A2(new_n22416_), .B(new_n22421_), .ZN(new_n22422_));
  AND2_X2    g19986(.A1(new_n22422_), .A2(new_n14291_), .Z(new_n22423_));
  NAND2_X1   g19987(.A1(new_n22423_), .A2(new_n12952_), .ZN(new_n22424_));
  AOI21_X1   g19988(.A1(new_n22424_), .A2(new_n12981_), .B(new_n12741_), .ZN(new_n22425_));
  NOR3_X1    g19989(.A1(new_n22425_), .A2(new_n12965_), .A3(new_n22412_), .ZN(new_n22426_));
  NOR2_X1    g19990(.A1(new_n22411_), .A2(pi0630), .ZN(new_n22427_));
  AOI21_X1   g19991(.A1(new_n22427_), .A2(new_n13384_), .B(new_n12741_), .ZN(new_n22428_));
  AOI21_X1   g19992(.A1(new_n22423_), .A2(new_n12952_), .B(new_n12981_), .ZN(new_n22429_));
  NOR2_X1    g19993(.A1(new_n22428_), .A2(new_n22429_), .ZN(new_n22430_));
  NOR2_X1    g19994(.A1(new_n22430_), .A2(pi1157), .ZN(new_n22431_));
  OAI21_X1   g19995(.A1(new_n22431_), .A2(new_n22426_), .B(pi0787), .ZN(new_n22432_));
  OAI21_X1   g19996(.A1(new_n22410_), .A2(pi0628), .B(pi0629), .ZN(new_n22433_));
  AOI21_X1   g19997(.A1(new_n22423_), .A2(pi0628), .B(new_n12742_), .ZN(new_n22434_));
  NOR2_X1    g19998(.A1(new_n22411_), .A2(pi0629), .ZN(new_n22435_));
  OAI22_X1   g19999(.A1(new_n22435_), .A2(new_n12920_), .B1(new_n12919_), .B2(new_n22423_), .ZN(new_n22436_));
  AOI22_X1   g20000(.A1(new_n22436_), .A2(new_n12742_), .B1(new_n22433_), .B2(new_n22434_), .ZN(new_n22437_));
  NOR2_X1    g20001(.A1(new_n22437_), .A2(new_n12937_), .ZN(new_n22438_));
  AOI21_X1   g20002(.A1(new_n22408_), .A2(pi0626), .B(new_n22403_), .ZN(new_n22439_));
  NAND2_X1   g20003(.A1(new_n22422_), .A2(new_n14289_), .ZN(new_n22440_));
  OAI21_X1   g20004(.A1(new_n22440_), .A2(new_n12910_), .B(new_n22413_), .ZN(new_n22441_));
  AOI21_X1   g20005(.A1(new_n22441_), .A2(new_n12748_), .B(pi0641), .ZN(new_n22442_));
  OAI21_X1   g20006(.A1(new_n12745_), .A2(new_n22439_), .B(new_n22442_), .ZN(new_n22443_));
  OAI21_X1   g20007(.A1(new_n22409_), .A2(pi0626), .B(new_n22413_), .ZN(new_n22444_));
  NAND2_X1   g20008(.A1(new_n22444_), .A2(new_n12745_), .ZN(new_n22445_));
  AOI21_X1   g20009(.A1(new_n22441_), .A2(new_n12746_), .B(new_n12814_), .ZN(new_n22446_));
  AOI21_X1   g20010(.A1(new_n22446_), .A2(new_n22445_), .B(new_n12808_), .ZN(new_n22447_));
  AOI21_X1   g20011(.A1(new_n22443_), .A2(new_n22447_), .B(new_n15340_), .ZN(new_n22448_));
  AOI21_X1   g20012(.A1(new_n22422_), .A2(new_n12870_), .B(new_n22403_), .ZN(new_n22449_));
  NAND2_X1   g20013(.A1(new_n22449_), .A2(pi0618), .ZN(new_n22450_));
  NOR2_X1    g20014(.A1(new_n22422_), .A2(pi0609), .ZN(new_n22451_));
  NOR2_X1    g20015(.A1(new_n14328_), .A2(new_n16844_), .ZN(new_n22452_));
  NOR3_X1    g20016(.A1(new_n22452_), .A2(new_n22404_), .A3(new_n22403_), .ZN(new_n22453_));
  NAND2_X1   g20017(.A1(new_n22453_), .A2(new_n12758_), .ZN(new_n22454_));
  NOR2_X1    g20018(.A1(new_n14330_), .A2(new_n16844_), .ZN(new_n22455_));
  INV_X1     g20019(.I(new_n22455_), .ZN(new_n22456_));
  NAND4_X1   g20020(.A1(new_n22456_), .A2(pi1153), .A3(new_n22413_), .A4(new_n22405_), .ZN(new_n22457_));
  NAND3_X1   g20021(.A1(new_n22457_), .A2(pi0608), .A3(new_n22420_), .ZN(new_n22458_));
  OAI21_X1   g20022(.A1(new_n22455_), .A2(new_n22453_), .B(new_n12841_), .ZN(new_n22459_));
  NAND3_X1   g20023(.A1(new_n22459_), .A2(new_n13560_), .A3(new_n22419_), .ZN(new_n22460_));
  NAND3_X1   g20024(.A1(new_n22458_), .A2(pi0778), .A3(new_n22460_), .ZN(new_n22461_));
  AOI21_X1   g20025(.A1(new_n22461_), .A2(new_n22454_), .B(new_n12766_), .ZN(new_n22462_));
  OAI21_X1   g20026(.A1(new_n22462_), .A2(new_n22451_), .B(pi1155), .ZN(new_n22463_));
  NAND2_X1   g20027(.A1(new_n22404_), .A2(new_n13353_), .ZN(new_n22464_));
  NAND3_X1   g20028(.A1(new_n22464_), .A2(new_n12770_), .A3(new_n22413_), .ZN(new_n22465_));
  NAND3_X1   g20029(.A1(new_n22463_), .A2(pi0660), .A3(new_n22465_), .ZN(new_n22466_));
  NAND2_X1   g20030(.A1(new_n22461_), .A2(new_n22454_), .ZN(new_n22467_));
  NOR2_X1    g20031(.A1(new_n22422_), .A2(new_n12766_), .ZN(new_n22468_));
  AOI21_X1   g20032(.A1(new_n22467_), .A2(new_n12766_), .B(new_n22468_), .ZN(new_n22469_));
  AOI21_X1   g20033(.A1(new_n22404_), .A2(new_n12772_), .B(new_n12770_), .ZN(new_n22470_));
  AOI21_X1   g20034(.A1(new_n22470_), .A2(new_n22413_), .B(pi0660), .ZN(new_n22471_));
  OAI21_X1   g20035(.A1(new_n22469_), .A2(pi1155), .B(new_n22471_), .ZN(new_n22472_));
  NAND3_X1   g20036(.A1(new_n22466_), .A2(new_n22472_), .A3(pi0785), .ZN(new_n22473_));
  NAND2_X1   g20037(.A1(new_n22467_), .A2(new_n12764_), .ZN(new_n22474_));
  NAND2_X1   g20038(.A1(new_n22473_), .A2(new_n22474_), .ZN(new_n22475_));
  NAND2_X1   g20039(.A1(new_n22475_), .A2(new_n12781_), .ZN(new_n22476_));
  AOI21_X1   g20040(.A1(new_n22476_), .A2(new_n22450_), .B(pi1154), .ZN(new_n22477_));
  OAI21_X1   g20041(.A1(new_n22407_), .A2(new_n15311_), .B(pi1154), .ZN(new_n22478_));
  NOR2_X1    g20042(.A1(new_n22478_), .A2(new_n22403_), .ZN(new_n22479_));
  NOR3_X1    g20043(.A1(new_n22477_), .A2(pi0627), .A3(new_n22479_), .ZN(new_n22480_));
  NAND2_X1   g20044(.A1(new_n22475_), .A2(pi0618), .ZN(new_n22481_));
  NAND2_X1   g20045(.A1(new_n22449_), .A2(new_n12781_), .ZN(new_n22482_));
  NAND2_X1   g20046(.A1(new_n22481_), .A2(new_n22482_), .ZN(new_n22483_));
  OAI21_X1   g20047(.A1(new_n22407_), .A2(new_n15304_), .B(new_n12785_), .ZN(new_n22484_));
  OAI21_X1   g20048(.A1(new_n22484_), .A2(new_n22403_), .B(pi0627), .ZN(new_n22485_));
  AOI21_X1   g20049(.A1(new_n22483_), .A2(pi1154), .B(new_n22485_), .ZN(new_n22486_));
  NOR3_X1    g20050(.A1(new_n22480_), .A2(new_n22486_), .A3(new_n12779_), .ZN(new_n22487_));
  AOI21_X1   g20051(.A1(new_n22473_), .A2(new_n22474_), .B(pi0781), .ZN(new_n22488_));
  OAI21_X1   g20052(.A1(new_n22487_), .A2(new_n22488_), .B(new_n17592_), .ZN(new_n22489_));
  NAND3_X1   g20053(.A1(new_n22406_), .A2(new_n15240_), .A3(pi0619), .ZN(new_n22490_));
  NAND2_X1   g20054(.A1(new_n22406_), .A2(new_n15271_), .ZN(new_n22491_));
  AOI22_X1   g20055(.A1(new_n22490_), .A2(new_n12907_), .B1(new_n22491_), .B2(new_n12908_), .ZN(new_n22492_));
  NAND2_X1   g20056(.A1(new_n22440_), .A2(new_n17599_), .ZN(new_n22493_));
  AOI21_X1   g20057(.A1(new_n22493_), .A2(new_n22492_), .B(new_n12796_), .ZN(new_n22494_));
  AOI21_X1   g20058(.A1(new_n22494_), .A2(new_n22413_), .B(new_n14303_), .ZN(new_n22495_));
  NAND2_X1   g20059(.A1(new_n22489_), .A2(new_n22495_), .ZN(new_n22496_));
  AOI22_X1   g20060(.A1(new_n22496_), .A2(new_n22448_), .B1(new_n22413_), .B2(new_n22438_), .ZN(new_n22497_));
  OAI22_X1   g20061(.A1(new_n22497_), .A2(new_n15341_), .B1(new_n22403_), .B2(new_n22432_), .ZN(new_n22498_));
  NAND2_X1   g20062(.A1(new_n22498_), .A2(new_n13000_), .ZN(new_n22499_));
  AND2_X2    g20063(.A1(new_n22498_), .A2(new_n12975_), .Z(new_n22500_));
  OAI21_X1   g20064(.A1(new_n22424_), .A2(new_n14300_), .B(new_n22413_), .ZN(new_n22501_));
  NOR2_X1    g20065(.A1(new_n22501_), .A2(new_n12975_), .ZN(new_n22502_));
  OAI21_X1   g20066(.A1(new_n22500_), .A2(new_n22502_), .B(new_n12740_), .ZN(new_n22503_));
  NAND2_X1   g20067(.A1(new_n17611_), .A2(new_n17504_), .ZN(new_n22504_));
  NOR2_X1    g20068(.A1(new_n22409_), .A2(new_n22504_), .ZN(new_n22505_));
  NAND2_X1   g20069(.A1(new_n22505_), .A2(new_n12975_), .ZN(new_n22506_));
  NAND3_X1   g20070(.A1(new_n22506_), .A2(pi0715), .A3(new_n22413_), .ZN(new_n22507_));
  NAND3_X1   g20071(.A1(new_n22503_), .A2(new_n12739_), .A3(new_n22507_), .ZN(new_n22508_));
  NOR2_X1    g20072(.A1(new_n22501_), .A2(pi0644), .ZN(new_n22509_));
  AOI21_X1   g20073(.A1(new_n22498_), .A2(pi0644), .B(new_n22509_), .ZN(new_n22510_));
  AOI21_X1   g20074(.A1(new_n22505_), .A2(pi0644), .B(pi0715), .ZN(new_n22511_));
  AOI21_X1   g20075(.A1(new_n22511_), .A2(new_n22413_), .B(new_n12739_), .ZN(new_n22512_));
  OAI21_X1   g20076(.A1(new_n22510_), .A2(new_n12740_), .B(new_n22512_), .ZN(new_n22513_));
  NAND3_X1   g20077(.A1(new_n22508_), .A2(pi0790), .A3(new_n22513_), .ZN(new_n22514_));
  AOI21_X1   g20078(.A1(new_n22514_), .A2(new_n22499_), .B(new_n12738_), .ZN(new_n22515_));
  AOI21_X1   g20079(.A1(pi0057), .A2(pi0189), .B(pi0832), .ZN(new_n22516_));
  NAND2_X1   g20080(.A1(new_n13192_), .A2(pi0189), .ZN(new_n22517_));
  NOR2_X1    g20081(.A1(new_n22517_), .A2(new_n13521_), .ZN(new_n22518_));
  NOR2_X1    g20082(.A1(new_n2610_), .A2(new_n16844_), .ZN(new_n22519_));
  NOR2_X1    g20083(.A1(new_n14122_), .A2(pi0189), .ZN(new_n22520_));
  NOR2_X1    g20084(.A1(new_n14118_), .A2(new_n9484_), .ZN(new_n22521_));
  OAI21_X1   g20085(.A1(new_n22521_), .A2(new_n22520_), .B(new_n3265_), .ZN(new_n22522_));
  NOR2_X1    g20086(.A1(new_n13344_), .A2(new_n9484_), .ZN(new_n22523_));
  NOR2_X1    g20087(.A1(new_n13398_), .A2(new_n22523_), .ZN(new_n22524_));
  NOR2_X1    g20088(.A1(new_n22524_), .A2(new_n3265_), .ZN(new_n22525_));
  INV_X1     g20089(.I(new_n22525_), .ZN(new_n22526_));
  NAND3_X1   g20090(.A1(new_n22522_), .A2(new_n22519_), .A3(new_n22526_), .ZN(new_n22527_));
  INV_X1     g20091(.I(new_n22519_), .ZN(new_n22528_));
  NAND2_X1   g20092(.A1(new_n22517_), .A2(new_n22528_), .ZN(new_n22529_));
  AND3_X2    g20093(.A1(new_n22527_), .A2(new_n13521_), .A3(new_n22529_), .Z(new_n22530_));
  OAI21_X1   g20094(.A1(new_n22530_), .A2(new_n22518_), .B(new_n12841_), .ZN(new_n22531_));
  NAND3_X1   g20095(.A1(new_n22527_), .A2(new_n22529_), .A3(pi0625), .ZN(new_n22532_));
  INV_X1     g20096(.I(new_n22517_), .ZN(new_n22533_));
  NAND2_X1   g20097(.A1(new_n22533_), .A2(new_n13521_), .ZN(new_n22534_));
  AOI21_X1   g20098(.A1(new_n22532_), .A2(new_n22534_), .B(new_n12841_), .ZN(new_n22535_));
  NOR2_X1    g20099(.A1(new_n22535_), .A2(new_n12758_), .ZN(new_n22536_));
  AOI21_X1   g20100(.A1(new_n22527_), .A2(new_n22529_), .B(pi0778), .ZN(new_n22537_));
  AOI21_X1   g20101(.A1(new_n22536_), .A2(new_n22531_), .B(new_n22537_), .ZN(new_n22538_));
  NOR2_X1    g20102(.A1(new_n22517_), .A2(new_n12870_), .ZN(new_n22539_));
  AOI21_X1   g20103(.A1(new_n22538_), .A2(new_n12870_), .B(new_n22539_), .ZN(new_n22540_));
  NOR2_X1    g20104(.A1(new_n22533_), .A2(new_n12888_), .ZN(new_n22541_));
  AOI21_X1   g20105(.A1(new_n22540_), .A2(new_n12888_), .B(new_n22541_), .ZN(new_n22542_));
  NOR2_X1    g20106(.A1(new_n22517_), .A2(new_n12911_), .ZN(new_n22543_));
  AOI21_X1   g20107(.A1(new_n22542_), .A2(new_n12911_), .B(new_n22543_), .ZN(new_n22544_));
  NOR2_X1    g20108(.A1(new_n22533_), .A2(new_n13392_), .ZN(new_n22545_));
  AOI21_X1   g20109(.A1(new_n22544_), .A2(new_n13392_), .B(new_n22545_), .ZN(new_n22546_));
  NAND2_X1   g20110(.A1(new_n22546_), .A2(new_n12920_), .ZN(new_n22547_));
  NAND2_X1   g20111(.A1(new_n22533_), .A2(pi0628), .ZN(new_n22548_));
  AOI21_X1   g20112(.A1(new_n22547_), .A2(new_n22548_), .B(pi1156), .ZN(new_n22549_));
  OR2_X2     g20113(.A1(new_n22549_), .A2(new_n12919_), .Z(new_n22550_));
  NOR2_X1    g20114(.A1(new_n2609_), .A2(new_n9484_), .ZN(new_n22551_));
  INV_X1     g20115(.I(new_n22551_), .ZN(new_n22552_));
  NOR2_X1    g20116(.A1(new_n5337_), .A2(new_n22405_), .ZN(new_n22553_));
  OAI21_X1   g20117(.A1(new_n22523_), .A2(new_n22553_), .B(pi0038), .ZN(new_n22554_));
  INV_X1     g20118(.I(new_n22554_), .ZN(new_n22555_));
  NAND3_X1   g20119(.A1(new_n13245_), .A2(new_n9484_), .A3(pi0772), .ZN(new_n22556_));
  NAND2_X1   g20120(.A1(new_n13256_), .A2(pi0772), .ZN(new_n22557_));
  NAND2_X1   g20121(.A1(new_n13060_), .A2(new_n16845_), .ZN(new_n22558_));
  AOI21_X1   g20122(.A1(new_n22557_), .A2(new_n22558_), .B(pi0039), .ZN(new_n22559_));
  AOI21_X1   g20123(.A1(new_n13322_), .A2(new_n13332_), .B(new_n16845_), .ZN(new_n22560_));
  NOR3_X1    g20124(.A1(new_n13178_), .A2(new_n13188_), .A3(pi0772), .ZN(new_n22561_));
  NOR3_X1    g20125(.A1(new_n22560_), .A2(new_n22561_), .A3(new_n2627_), .ZN(new_n22562_));
  OAI21_X1   g20126(.A1(new_n22562_), .A2(new_n22559_), .B(pi0189), .ZN(new_n22563_));
  AOI21_X1   g20127(.A1(new_n22563_), .A2(new_n22556_), .B(pi0038), .ZN(new_n22564_));
  OAI21_X1   g20128(.A1(new_n22564_), .A2(new_n22555_), .B(new_n2609_), .ZN(new_n22565_));
  NAND2_X1   g20129(.A1(new_n22565_), .A2(new_n22552_), .ZN(new_n22566_));
  NAND2_X1   g20130(.A1(new_n22566_), .A2(new_n12761_), .ZN(new_n22567_));
  OAI21_X1   g20131(.A1(new_n12761_), .A2(new_n22517_), .B(new_n22567_), .ZN(new_n22568_));
  NOR2_X1    g20132(.A1(new_n22517_), .A2(new_n12766_), .ZN(new_n22569_));
  AOI21_X1   g20133(.A1(new_n22568_), .A2(new_n12766_), .B(new_n22569_), .ZN(new_n22570_));
  NOR2_X1    g20134(.A1(new_n22570_), .A2(pi1155), .ZN(new_n22571_));
  NOR2_X1    g20135(.A1(new_n22517_), .A2(pi0609), .ZN(new_n22572_));
  AOI21_X1   g20136(.A1(new_n22568_), .A2(pi0609), .B(new_n22572_), .ZN(new_n22573_));
  OAI21_X1   g20137(.A1(new_n22573_), .A2(new_n12770_), .B(pi0785), .ZN(new_n22574_));
  OAI22_X1   g20138(.A1(new_n22574_), .A2(new_n22571_), .B1(pi0785), .B2(new_n22568_), .ZN(new_n22575_));
  NAND2_X1   g20139(.A1(new_n22533_), .A2(pi0618), .ZN(new_n22576_));
  OAI21_X1   g20140(.A1(new_n22575_), .A2(pi0618), .B(new_n22576_), .ZN(new_n22577_));
  NAND2_X1   g20141(.A1(new_n22577_), .A2(new_n12785_), .ZN(new_n22578_));
  NAND2_X1   g20142(.A1(new_n22533_), .A2(new_n12781_), .ZN(new_n22579_));
  OAI21_X1   g20143(.A1(new_n22575_), .A2(new_n12781_), .B(new_n22579_), .ZN(new_n22580_));
  AOI21_X1   g20144(.A1(new_n22580_), .A2(pi1154), .B(new_n12779_), .ZN(new_n22581_));
  AOI22_X1   g20145(.A1(new_n22581_), .A2(new_n22578_), .B1(new_n12779_), .B2(new_n22575_), .ZN(new_n22582_));
  NOR2_X1    g20146(.A1(new_n22582_), .A2(pi0789), .ZN(new_n22583_));
  NOR2_X1    g20147(.A1(new_n22517_), .A2(new_n12793_), .ZN(new_n22584_));
  AOI21_X1   g20148(.A1(new_n22582_), .A2(new_n12793_), .B(new_n22584_), .ZN(new_n22585_));
  NOR2_X1    g20149(.A1(new_n22585_), .A2(pi1159), .ZN(new_n22586_));
  NOR2_X1    g20150(.A1(new_n22517_), .A2(pi0619), .ZN(new_n22587_));
  AOI21_X1   g20151(.A1(new_n22582_), .A2(pi0619), .B(new_n22587_), .ZN(new_n22588_));
  NOR2_X1    g20152(.A1(new_n22588_), .A2(new_n12791_), .ZN(new_n22589_));
  NOR3_X1    g20153(.A1(new_n22586_), .A2(new_n22589_), .A3(new_n12796_), .ZN(new_n22590_));
  NOR2_X1    g20154(.A1(new_n22590_), .A2(new_n22583_), .ZN(new_n22591_));
  NOR2_X1    g20155(.A1(new_n22591_), .A2(new_n12818_), .ZN(new_n22592_));
  AOI21_X1   g20156(.A1(new_n12818_), .A2(new_n22517_), .B(new_n22592_), .ZN(new_n22593_));
  NOR2_X1    g20157(.A1(new_n22593_), .A2(pi0628), .ZN(new_n22594_));
  NOR2_X1    g20158(.A1(new_n22594_), .A2(new_n12742_), .ZN(new_n22595_));
  AOI21_X1   g20159(.A1(new_n22533_), .A2(new_n12747_), .B(pi0641), .ZN(new_n22596_));
  INV_X1     g20160(.I(new_n22596_), .ZN(new_n22597_));
  NOR3_X1    g20161(.A1(new_n22590_), .A2(new_n12747_), .A3(new_n22583_), .ZN(new_n22598_));
  OAI21_X1   g20162(.A1(new_n22598_), .A2(new_n22597_), .B(pi1158), .ZN(new_n22599_));
  INV_X1     g20163(.I(new_n22544_), .ZN(new_n22600_));
  AOI21_X1   g20164(.A1(new_n22600_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n22601_));
  NOR3_X1    g20165(.A1(new_n22555_), .A2(new_n16844_), .A3(new_n15123_), .ZN(new_n22602_));
  AOI21_X1   g20166(.A1(new_n13692_), .A2(pi0189), .B(new_n16845_), .ZN(new_n22603_));
  OAI21_X1   g20167(.A1(new_n14187_), .A2(pi0189), .B(new_n22603_), .ZN(new_n22604_));
  OAI21_X1   g20168(.A1(new_n13794_), .A2(new_n13786_), .B(new_n9484_), .ZN(new_n22605_));
  OAI21_X1   g20169(.A1(new_n13745_), .A2(new_n13754_), .B(pi0189), .ZN(new_n22606_));
  NAND3_X1   g20170(.A1(new_n22606_), .A2(new_n16845_), .A3(new_n22605_), .ZN(new_n22607_));
  NAND3_X1   g20171(.A1(new_n22604_), .A2(new_n22607_), .A3(pi0039), .ZN(new_n22608_));
  AOI21_X1   g20172(.A1(new_n13416_), .A2(new_n13798_), .B(pi0189), .ZN(new_n22609_));
  NOR2_X1    g20173(.A1(new_n13800_), .A2(new_n9484_), .ZN(new_n22610_));
  OAI21_X1   g20174(.A1(new_n22610_), .A2(new_n22609_), .B(pi0772), .ZN(new_n22611_));
  NOR3_X1    g20175(.A1(new_n13809_), .A2(new_n13406_), .A3(new_n9484_), .ZN(new_n22612_));
  AOI21_X1   g20176(.A1(new_n13805_), .A2(new_n13807_), .B(pi0189), .ZN(new_n22613_));
  OAI21_X1   g20177(.A1(new_n22612_), .A2(new_n22613_), .B(new_n16845_), .ZN(new_n22614_));
  NAND3_X1   g20178(.A1(new_n22611_), .A2(new_n22614_), .A3(new_n2627_), .ZN(new_n22615_));
  NAND3_X1   g20179(.A1(new_n22608_), .A2(new_n22615_), .A3(new_n3265_), .ZN(new_n22616_));
  AOI21_X1   g20180(.A1(new_n22616_), .A2(new_n22602_), .B(new_n2610_), .ZN(new_n22617_));
  OR3_X2     g20181(.A1(new_n22564_), .A2(pi0727), .A3(new_n22555_), .Z(new_n22618_));
  AOI21_X1   g20182(.A1(new_n22617_), .A2(new_n22618_), .B(new_n22551_), .ZN(new_n22619_));
  NOR2_X1    g20183(.A1(new_n22619_), .A2(new_n13521_), .ZN(new_n22620_));
  AOI21_X1   g20184(.A1(new_n22565_), .A2(new_n22552_), .B(pi0625), .ZN(new_n22621_));
  OAI21_X1   g20185(.A1(new_n22620_), .A2(new_n22621_), .B(pi1153), .ZN(new_n22622_));
  NAND3_X1   g20186(.A1(new_n22622_), .A2(pi0608), .A3(new_n22531_), .ZN(new_n22623_));
  NAND2_X1   g20187(.A1(new_n22566_), .A2(pi0625), .ZN(new_n22624_));
  OAI21_X1   g20188(.A1(new_n22619_), .A2(pi0625), .B(new_n22624_), .ZN(new_n22625_));
  AOI21_X1   g20189(.A1(new_n22625_), .A2(new_n12841_), .B(new_n22535_), .ZN(new_n22626_));
  AOI21_X1   g20190(.A1(new_n22626_), .A2(new_n13560_), .B(new_n12758_), .ZN(new_n22627_));
  NOR2_X1    g20191(.A1(new_n22619_), .A2(pi0778), .ZN(new_n22628_));
  AOI21_X1   g20192(.A1(new_n22627_), .A2(new_n22623_), .B(new_n22628_), .ZN(new_n22629_));
  NOR2_X1    g20193(.A1(new_n22629_), .A2(pi0785), .ZN(new_n22630_));
  INV_X1     g20194(.I(new_n22630_), .ZN(new_n22631_));
  NOR2_X1    g20195(.A1(new_n22571_), .A2(new_n13829_), .ZN(new_n22632_));
  INV_X1     g20196(.I(new_n22632_), .ZN(new_n22633_));
  INV_X1     g20197(.I(new_n22538_), .ZN(new_n22634_));
  AOI21_X1   g20198(.A1(new_n22634_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n22635_));
  NAND2_X1   g20199(.A1(new_n22629_), .A2(pi0609), .ZN(new_n22636_));
  AOI21_X1   g20200(.A1(new_n22636_), .A2(new_n22635_), .B(new_n22633_), .ZN(new_n22637_));
  OAI21_X1   g20201(.A1(new_n22573_), .A2(new_n12770_), .B(new_n13829_), .ZN(new_n22638_));
  OAI21_X1   g20202(.A1(new_n22538_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n22639_));
  AOI21_X1   g20203(.A1(new_n22629_), .A2(new_n12766_), .B(new_n22639_), .ZN(new_n22640_));
  OAI21_X1   g20204(.A1(new_n22640_), .A2(new_n22638_), .B(pi0785), .ZN(new_n22641_));
  OAI21_X1   g20205(.A1(new_n22641_), .A2(new_n22637_), .B(new_n22631_), .ZN(new_n22642_));
  NAND2_X1   g20206(.A1(new_n22642_), .A2(new_n12779_), .ZN(new_n22643_));
  INV_X1     g20207(.I(new_n22643_), .ZN(new_n22644_));
  AOI21_X1   g20208(.A1(new_n22577_), .A2(new_n12785_), .B(new_n12880_), .ZN(new_n22645_));
  AOI21_X1   g20209(.A1(new_n22540_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n22646_));
  OAI21_X1   g20210(.A1(new_n22642_), .A2(new_n12781_), .B(new_n22646_), .ZN(new_n22647_));
  NAND2_X1   g20211(.A1(new_n22647_), .A2(new_n22645_), .ZN(new_n22648_));
  AOI21_X1   g20212(.A1(new_n22580_), .A2(pi1154), .B(pi0627), .ZN(new_n22649_));
  AOI21_X1   g20213(.A1(new_n22540_), .A2(pi0618), .B(pi1154), .ZN(new_n22650_));
  OAI21_X1   g20214(.A1(new_n22642_), .A2(pi0618), .B(new_n22650_), .ZN(new_n22651_));
  AOI21_X1   g20215(.A1(new_n22651_), .A2(new_n22649_), .B(new_n12779_), .ZN(new_n22652_));
  AOI21_X1   g20216(.A1(new_n22652_), .A2(new_n22648_), .B(new_n22644_), .ZN(new_n22653_));
  NOR2_X1    g20217(.A1(new_n22653_), .A2(pi0789), .ZN(new_n22654_));
  INV_X1     g20218(.I(new_n22654_), .ZN(new_n22655_));
  OAI21_X1   g20219(.A1(new_n22585_), .A2(pi1159), .B(pi0648), .ZN(new_n22656_));
  INV_X1     g20220(.I(new_n22542_), .ZN(new_n22657_));
  AOI21_X1   g20221(.A1(new_n22657_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n22658_));
  NAND2_X1   g20222(.A1(new_n22653_), .A2(pi0619), .ZN(new_n22659_));
  AOI21_X1   g20223(.A1(new_n22659_), .A2(new_n22658_), .B(new_n22656_), .ZN(new_n22660_));
  NOR2_X1    g20224(.A1(new_n22589_), .A2(pi0648), .ZN(new_n22661_));
  INV_X1     g20225(.I(new_n22661_), .ZN(new_n22662_));
  AOI21_X1   g20226(.A1(new_n22657_), .A2(pi0619), .B(pi1159), .ZN(new_n22663_));
  INV_X1     g20227(.I(new_n22663_), .ZN(new_n22664_));
  AOI21_X1   g20228(.A1(new_n22653_), .A2(new_n12793_), .B(new_n22664_), .ZN(new_n22665_));
  OAI21_X1   g20229(.A1(new_n22665_), .A2(new_n22662_), .B(pi0789), .ZN(new_n22666_));
  OAI21_X1   g20230(.A1(new_n22666_), .A2(new_n22660_), .B(new_n22655_), .ZN(new_n22667_));
  NAND2_X1   g20231(.A1(new_n22667_), .A2(pi0626), .ZN(new_n22668_));
  AOI21_X1   g20232(.A1(new_n22668_), .A2(new_n22601_), .B(new_n22599_), .ZN(new_n22669_));
  AOI21_X1   g20233(.A1(new_n22533_), .A2(pi0626), .B(new_n12814_), .ZN(new_n22670_));
  NAND2_X1   g20234(.A1(new_n22591_), .A2(new_n12747_), .ZN(new_n22671_));
  NAND2_X1   g20235(.A1(new_n22671_), .A2(new_n22670_), .ZN(new_n22672_));
  NAND2_X1   g20236(.A1(new_n22672_), .A2(new_n12745_), .ZN(new_n22673_));
  AOI21_X1   g20237(.A1(new_n22600_), .A2(pi0626), .B(pi0641), .ZN(new_n22674_));
  INV_X1     g20238(.I(new_n22674_), .ZN(new_n22675_));
  AOI21_X1   g20239(.A1(new_n22667_), .A2(new_n12747_), .B(new_n22675_), .ZN(new_n22676_));
  OAI21_X1   g20240(.A1(new_n22676_), .A2(new_n22673_), .B(pi0788), .ZN(new_n22677_));
  OR2_X2     g20241(.A1(new_n22667_), .A2(pi0788), .Z(new_n22678_));
  OAI21_X1   g20242(.A1(new_n22677_), .A2(new_n22669_), .B(new_n22678_), .ZN(new_n22679_));
  NAND2_X1   g20243(.A1(new_n22679_), .A2(pi0628), .ZN(new_n22680_));
  AOI21_X1   g20244(.A1(new_n22680_), .A2(new_n22595_), .B(new_n22550_), .ZN(new_n22681_));
  NOR2_X1    g20245(.A1(new_n22517_), .A2(pi0628), .ZN(new_n22682_));
  AOI21_X1   g20246(.A1(new_n22546_), .A2(pi0628), .B(new_n22682_), .ZN(new_n22683_));
  OAI21_X1   g20247(.A1(new_n22683_), .A2(new_n12742_), .B(new_n12919_), .ZN(new_n22684_));
  OAI21_X1   g20248(.A1(new_n22593_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n22685_));
  AOI21_X1   g20249(.A1(new_n22679_), .A2(new_n12920_), .B(new_n22685_), .ZN(new_n22686_));
  OAI21_X1   g20250(.A1(new_n22686_), .A2(new_n22684_), .B(pi0792), .ZN(new_n22687_));
  OR2_X2     g20251(.A1(new_n22679_), .A2(pi0792), .Z(new_n22688_));
  OAI21_X1   g20252(.A1(new_n22687_), .A2(new_n22681_), .B(new_n22688_), .ZN(new_n22689_));
  AND2_X2    g20253(.A1(new_n22689_), .A2(new_n12972_), .Z(new_n22690_));
  NOR2_X1    g20254(.A1(new_n22546_), .A2(pi0792), .ZN(new_n22691_));
  OAI21_X1   g20255(.A1(new_n22683_), .A2(new_n12742_), .B(pi0792), .ZN(new_n22692_));
  NOR2_X1    g20256(.A1(new_n22692_), .A2(new_n22549_), .ZN(new_n22693_));
  NOR2_X1    g20257(.A1(new_n22693_), .A2(new_n22691_), .ZN(new_n22694_));
  NAND2_X1   g20258(.A1(new_n22694_), .A2(new_n12741_), .ZN(new_n22695_));
  NAND2_X1   g20259(.A1(new_n22533_), .A2(pi0647), .ZN(new_n22696_));
  AOI21_X1   g20260(.A1(new_n22695_), .A2(new_n22696_), .B(pi1157), .ZN(new_n22697_));
  NOR2_X1    g20261(.A1(new_n22697_), .A2(new_n12981_), .ZN(new_n22698_));
  NAND2_X1   g20262(.A1(new_n22517_), .A2(new_n12943_), .ZN(new_n22699_));
  OAI21_X1   g20263(.A1(new_n22593_), .A2(new_n12943_), .B(new_n22699_), .ZN(new_n22700_));
  AOI21_X1   g20264(.A1(new_n22700_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n22701_));
  OAI21_X1   g20265(.A1(new_n22689_), .A2(new_n12741_), .B(new_n22701_), .ZN(new_n22702_));
  NAND2_X1   g20266(.A1(new_n22702_), .A2(new_n22698_), .ZN(new_n22703_));
  NOR2_X1    g20267(.A1(new_n22517_), .A2(pi0647), .ZN(new_n22704_));
  AOI21_X1   g20268(.A1(new_n22694_), .A2(pi0647), .B(new_n22704_), .ZN(new_n22705_));
  NOR2_X1    g20269(.A1(new_n22705_), .A2(new_n12965_), .ZN(new_n22706_));
  NOR2_X1    g20270(.A1(new_n22706_), .A2(pi0630), .ZN(new_n22707_));
  AOI21_X1   g20271(.A1(new_n22700_), .A2(pi0647), .B(pi1157), .ZN(new_n22708_));
  OAI21_X1   g20272(.A1(new_n22689_), .A2(pi0647), .B(new_n22708_), .ZN(new_n22709_));
  AOI21_X1   g20273(.A1(new_n22709_), .A2(new_n22707_), .B(new_n12972_), .ZN(new_n22710_));
  AOI21_X1   g20274(.A1(new_n22710_), .A2(new_n22703_), .B(new_n22690_), .ZN(new_n22711_));
  OAI21_X1   g20275(.A1(new_n22711_), .A2(pi0790), .B(new_n5477_), .ZN(new_n22712_));
  OAI21_X1   g20276(.A1(new_n22533_), .A2(new_n12975_), .B(pi0715), .ZN(new_n22713_));
  NAND2_X1   g20277(.A1(new_n22533_), .A2(new_n12984_), .ZN(new_n22714_));
  OAI21_X1   g20278(.A1(new_n22700_), .A2(new_n12984_), .B(new_n22714_), .ZN(new_n22715_));
  NOR2_X1    g20279(.A1(new_n22715_), .A2(pi0644), .ZN(new_n22716_));
  OAI21_X1   g20280(.A1(new_n22716_), .A2(new_n22713_), .B(new_n12739_), .ZN(new_n22717_));
  NOR2_X1    g20281(.A1(new_n22706_), .A2(new_n12972_), .ZN(new_n22718_));
  INV_X1     g20282(.I(new_n22718_), .ZN(new_n22719_));
  OAI22_X1   g20283(.A1(new_n22719_), .A2(new_n22697_), .B1(pi0787), .B2(new_n22694_), .ZN(new_n22720_));
  AOI21_X1   g20284(.A1(new_n22720_), .A2(pi0644), .B(pi0715), .ZN(new_n22721_));
  NAND2_X1   g20285(.A1(new_n22711_), .A2(new_n12975_), .ZN(new_n22722_));
  AOI21_X1   g20286(.A1(new_n22722_), .A2(new_n22721_), .B(new_n22717_), .ZN(new_n22723_));
  OAI21_X1   g20287(.A1(new_n22533_), .A2(pi0644), .B(new_n12740_), .ZN(new_n22724_));
  NOR2_X1    g20288(.A1(new_n22715_), .A2(new_n12975_), .ZN(new_n22725_));
  OAI21_X1   g20289(.A1(new_n22725_), .A2(new_n22724_), .B(pi1160), .ZN(new_n22726_));
  NAND2_X1   g20290(.A1(new_n22720_), .A2(new_n12975_), .ZN(new_n22727_));
  NAND2_X1   g20291(.A1(new_n22727_), .A2(pi0715), .ZN(new_n22728_));
  AOI21_X1   g20292(.A1(new_n22711_), .A2(pi0644), .B(new_n22728_), .ZN(new_n22729_));
  OAI21_X1   g20293(.A1(new_n22729_), .A2(new_n22726_), .B(pi0790), .ZN(new_n22730_));
  NOR2_X1    g20294(.A1(new_n22730_), .A2(new_n22723_), .ZN(new_n22731_));
  AOI21_X1   g20295(.A1(new_n6165_), .A2(new_n9484_), .B(pi0057), .ZN(new_n22732_));
  OAI21_X1   g20296(.A1(new_n22731_), .A2(new_n22712_), .B(new_n22732_), .ZN(new_n22733_));
  AOI21_X1   g20297(.A1(new_n22733_), .A2(new_n22516_), .B(new_n22515_), .ZN(po0346));
  NOR2_X1    g20298(.A1(new_n3042_), .A2(pi0190), .ZN(new_n22735_));
  NOR2_X1    g20299(.A1(new_n13340_), .A2(new_n16945_), .ZN(new_n22736_));
  NOR2_X1    g20300(.A1(new_n22736_), .A2(new_n22735_), .ZN(new_n22737_));
  NOR3_X1    g20301(.A1(new_n22737_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n22738_));
  INV_X1     g20302(.I(new_n22736_), .ZN(new_n22739_));
  NOR2_X1    g20303(.A1(new_n22739_), .A2(new_n13354_), .ZN(new_n22740_));
  NOR3_X1    g20304(.A1(new_n22740_), .A2(new_n12762_), .A3(new_n22737_), .ZN(new_n22741_));
  NOR2_X1    g20305(.A1(new_n22741_), .A2(new_n12770_), .ZN(new_n22742_));
  NOR3_X1    g20306(.A1(new_n22740_), .A2(pi1155), .A3(new_n22735_), .ZN(new_n22743_));
  NOR3_X1    g20307(.A1(new_n22742_), .A2(new_n12764_), .A3(new_n22743_), .ZN(new_n22744_));
  NOR2_X1    g20308(.A1(new_n22744_), .A2(new_n22738_), .ZN(new_n22745_));
  NOR2_X1    g20309(.A1(new_n22745_), .A2(pi0781), .ZN(new_n22746_));
  INV_X1     g20310(.I(new_n22745_), .ZN(new_n22747_));
  AOI21_X1   g20311(.A1(new_n22747_), .A2(new_n12783_), .B(pi1154), .ZN(new_n22748_));
  AOI21_X1   g20312(.A1(new_n22747_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n22749_));
  NOR3_X1    g20313(.A1(new_n22748_), .A2(new_n22749_), .A3(new_n12779_), .ZN(new_n22750_));
  NOR2_X1    g20314(.A1(new_n22750_), .A2(new_n22746_), .ZN(new_n22751_));
  NOR2_X1    g20315(.A1(new_n22751_), .A2(new_n17229_), .ZN(new_n22752_));
  NOR2_X1    g20316(.A1(new_n22752_), .A2(pi1159), .ZN(new_n22753_));
  OAI21_X1   g20317(.A1(new_n22751_), .A2(new_n17232_), .B(pi1159), .ZN(new_n22754_));
  NAND2_X1   g20318(.A1(new_n22754_), .A2(pi0789), .ZN(new_n22755_));
  OAI22_X1   g20319(.A1(new_n22755_), .A2(new_n22753_), .B1(pi0789), .B2(new_n22751_), .ZN(new_n22756_));
  INV_X1     g20320(.I(new_n22735_), .ZN(new_n22757_));
  NAND2_X1   g20321(.A1(new_n12818_), .A2(new_n22757_), .ZN(new_n22758_));
  OAI21_X1   g20322(.A1(new_n22756_), .A2(new_n12818_), .B(new_n22758_), .ZN(new_n22759_));
  AOI21_X1   g20323(.A1(new_n12826_), .A2(pi0699), .B(new_n22735_), .ZN(new_n22760_));
  INV_X1     g20324(.I(pi0699), .ZN(new_n22761_));
  NOR2_X1    g20325(.A1(new_n12834_), .A2(new_n22761_), .ZN(new_n22762_));
  INV_X1     g20326(.I(new_n22762_), .ZN(new_n22763_));
  NOR2_X1    g20327(.A1(new_n22735_), .A2(pi1153), .ZN(new_n22764_));
  NAND2_X1   g20328(.A1(new_n22763_), .A2(new_n22764_), .ZN(new_n22765_));
  NOR2_X1    g20329(.A1(new_n22762_), .A2(new_n22760_), .ZN(new_n22766_));
  NOR2_X1    g20330(.A1(new_n22766_), .A2(new_n12841_), .ZN(new_n22767_));
  INV_X1     g20331(.I(new_n22767_), .ZN(new_n22768_));
  NAND3_X1   g20332(.A1(new_n22768_), .A2(pi0778), .A3(new_n22765_), .ZN(new_n22769_));
  OAI21_X1   g20333(.A1(pi0778), .A2(new_n22760_), .B(new_n22769_), .ZN(new_n22770_));
  NAND2_X1   g20334(.A1(new_n22770_), .A2(new_n17187_), .ZN(new_n22771_));
  NOR2_X1    g20335(.A1(new_n22771_), .A2(new_n12889_), .ZN(new_n22772_));
  INV_X1     g20336(.I(new_n22772_), .ZN(new_n22773_));
  NOR2_X1    g20337(.A1(new_n22773_), .A2(new_n12912_), .ZN(new_n22774_));
  INV_X1     g20338(.I(new_n22774_), .ZN(new_n22775_));
  NOR2_X1    g20339(.A1(new_n22775_), .A2(new_n17884_), .ZN(new_n22776_));
  INV_X1     g20340(.I(new_n22776_), .ZN(new_n22777_));
  OAI22_X1   g20341(.A1(new_n22759_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n22777_), .ZN(new_n22778_));
  NAND2_X1   g20342(.A1(new_n22778_), .A2(new_n12919_), .ZN(new_n22779_));
  OAI22_X1   g20343(.A1(new_n22759_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n22777_), .ZN(new_n22780_));
  NAND2_X1   g20344(.A1(new_n22780_), .A2(pi0629), .ZN(new_n22781_));
  AOI21_X1   g20345(.A1(new_n22779_), .A2(new_n22781_), .B(new_n12937_), .ZN(new_n22782_));
  INV_X1     g20346(.I(new_n22743_), .ZN(new_n22783_));
  NOR2_X1    g20347(.A1(new_n22760_), .A2(new_n12754_), .ZN(new_n22784_));
  NOR3_X1    g20348(.A1(new_n22784_), .A2(new_n22735_), .A3(new_n22736_), .ZN(new_n22785_));
  NAND2_X1   g20349(.A1(new_n22785_), .A2(new_n12758_), .ZN(new_n22786_));
  NAND2_X1   g20350(.A1(new_n22784_), .A2(pi0625), .ZN(new_n22787_));
  NAND3_X1   g20351(.A1(new_n22787_), .A2(pi1153), .A3(new_n22737_), .ZN(new_n22788_));
  NAND3_X1   g20352(.A1(new_n22765_), .A2(pi0608), .A3(new_n22788_), .ZN(new_n22789_));
  INV_X1     g20353(.I(new_n22787_), .ZN(new_n22790_));
  OAI21_X1   g20354(.A1(new_n22790_), .A2(new_n22785_), .B(new_n22764_), .ZN(new_n22791_));
  NAND3_X1   g20355(.A1(new_n22768_), .A2(new_n13560_), .A3(new_n22791_), .ZN(new_n22792_));
  NAND3_X1   g20356(.A1(new_n22792_), .A2(pi0778), .A3(new_n22789_), .ZN(new_n22793_));
  AOI21_X1   g20357(.A1(new_n22793_), .A2(new_n22786_), .B(new_n12766_), .ZN(new_n22794_));
  NOR2_X1    g20358(.A1(new_n22770_), .A2(pi0609), .ZN(new_n22795_));
  OAI21_X1   g20359(.A1(new_n22795_), .A2(new_n22794_), .B(pi1155), .ZN(new_n22796_));
  NAND3_X1   g20360(.A1(new_n22796_), .A2(pi0660), .A3(new_n22783_), .ZN(new_n22797_));
  NAND2_X1   g20361(.A1(new_n22793_), .A2(new_n22786_), .ZN(new_n22798_));
  NOR2_X1    g20362(.A1(new_n22770_), .A2(new_n12766_), .ZN(new_n22799_));
  AOI21_X1   g20363(.A1(new_n22798_), .A2(new_n12766_), .B(new_n22799_), .ZN(new_n22800_));
  NOR2_X1    g20364(.A1(new_n22742_), .A2(pi0660), .ZN(new_n22801_));
  OAI21_X1   g20365(.A1(new_n22800_), .A2(pi1155), .B(new_n22801_), .ZN(new_n22802_));
  NAND3_X1   g20366(.A1(new_n22802_), .A2(new_n22797_), .A3(pi0785), .ZN(new_n22803_));
  NAND2_X1   g20367(.A1(new_n22798_), .A2(new_n12764_), .ZN(new_n22804_));
  NAND2_X1   g20368(.A1(new_n22803_), .A2(new_n22804_), .ZN(new_n22805_));
  NAND2_X1   g20369(.A1(new_n22805_), .A2(new_n12781_), .ZN(new_n22806_));
  NAND2_X1   g20370(.A1(new_n22771_), .A2(pi0618), .ZN(new_n22807_));
  AOI21_X1   g20371(.A1(new_n22806_), .A2(new_n22807_), .B(pi1154), .ZN(new_n22808_));
  NOR3_X1    g20372(.A1(new_n22808_), .A2(pi0627), .A3(new_n22749_), .ZN(new_n22809_));
  NAND2_X1   g20373(.A1(new_n22771_), .A2(new_n12781_), .ZN(new_n22810_));
  NAND2_X1   g20374(.A1(new_n22805_), .A2(pi0618), .ZN(new_n22811_));
  AOI21_X1   g20375(.A1(new_n22811_), .A2(new_n22810_), .B(new_n12785_), .ZN(new_n22812_));
  NOR3_X1    g20376(.A1(new_n22812_), .A2(new_n12880_), .A3(new_n22748_), .ZN(new_n22813_));
  OR3_X2     g20377(.A1(new_n22809_), .A2(new_n22813_), .A3(new_n12779_), .Z(new_n22814_));
  NAND2_X1   g20378(.A1(new_n22805_), .A2(new_n12779_), .ZN(new_n22815_));
  NAND2_X1   g20379(.A1(new_n22814_), .A2(new_n22815_), .ZN(new_n22816_));
  AOI21_X1   g20380(.A1(new_n22816_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n22817_));
  NAND2_X1   g20381(.A1(new_n22773_), .A2(new_n12793_), .ZN(new_n22818_));
  NAND2_X1   g20382(.A1(new_n22816_), .A2(pi0619), .ZN(new_n22819_));
  AOI21_X1   g20383(.A1(new_n22819_), .A2(new_n22818_), .B(new_n12791_), .ZN(new_n22820_));
  NOR3_X1    g20384(.A1(new_n22820_), .A2(new_n12895_), .A3(new_n22753_), .ZN(new_n22821_));
  AOI21_X1   g20385(.A1(new_n22814_), .A2(new_n22815_), .B(pi0619), .ZN(new_n22822_));
  NOR2_X1    g20386(.A1(new_n22772_), .A2(new_n12793_), .ZN(new_n22823_));
  OAI21_X1   g20387(.A1(new_n22822_), .A2(new_n22823_), .B(new_n12791_), .ZN(new_n22824_));
  NAND3_X1   g20388(.A1(new_n22824_), .A2(new_n12895_), .A3(new_n22754_), .ZN(new_n22825_));
  NAND2_X1   g20389(.A1(new_n22825_), .A2(pi0789), .ZN(new_n22826_));
  OAI21_X1   g20390(.A1(new_n22826_), .A2(new_n22821_), .B(new_n22817_), .ZN(new_n22827_));
  NAND2_X1   g20391(.A1(new_n22735_), .A2(pi0626), .ZN(new_n22828_));
  NAND2_X1   g20392(.A1(new_n22756_), .A2(new_n12747_), .ZN(new_n22829_));
  AOI21_X1   g20393(.A1(new_n22829_), .A2(new_n22828_), .B(new_n12816_), .ZN(new_n22830_));
  NOR2_X1    g20394(.A1(new_n22757_), .A2(pi0626), .ZN(new_n22831_));
  AOI21_X1   g20395(.A1(new_n22756_), .A2(pi0626), .B(new_n22831_), .ZN(new_n22832_));
  OAI22_X1   g20396(.A1(new_n22832_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n22775_), .ZN(new_n22833_));
  OAI21_X1   g20397(.A1(new_n22833_), .A2(new_n22830_), .B(pi0788), .ZN(new_n22834_));
  AOI21_X1   g20398(.A1(new_n22827_), .A2(new_n22834_), .B(new_n15340_), .ZN(new_n22835_));
  OR2_X2     g20399(.A1(new_n22835_), .A2(new_n22782_), .Z(new_n22836_));
  NAND2_X1   g20400(.A1(new_n22759_), .A2(new_n13384_), .ZN(new_n22837_));
  NAND2_X1   g20401(.A1(new_n12943_), .A2(new_n22757_), .ZN(new_n22838_));
  AOI21_X1   g20402(.A1(new_n22837_), .A2(new_n22838_), .B(new_n17212_), .ZN(new_n22839_));
  NOR2_X1    g20403(.A1(new_n22777_), .A2(new_n12953_), .ZN(new_n22840_));
  NOR2_X1    g20404(.A1(new_n22840_), .A2(pi0647), .ZN(new_n22841_));
  NOR2_X1    g20405(.A1(new_n22735_), .A2(new_n12741_), .ZN(new_n22842_));
  OAI21_X1   g20406(.A1(new_n22841_), .A2(new_n22842_), .B(new_n12965_), .ZN(new_n22843_));
  NOR2_X1    g20407(.A1(new_n22757_), .A2(pi0647), .ZN(new_n22844_));
  AOI21_X1   g20408(.A1(new_n22840_), .A2(pi0647), .B(new_n22844_), .ZN(new_n22845_));
  INV_X1     g20409(.I(new_n22845_), .ZN(new_n22846_));
  OAI22_X1   g20410(.A1(new_n22843_), .A2(new_n12981_), .B1(new_n22846_), .B2(new_n15576_), .ZN(new_n22847_));
  NOR2_X1    g20411(.A1(new_n22847_), .A2(new_n22839_), .ZN(new_n22848_));
  OAI22_X1   g20412(.A1(new_n22836_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n22848_), .ZN(new_n22849_));
  OAI21_X1   g20413(.A1(new_n12965_), .A2(new_n22846_), .B(new_n22843_), .ZN(new_n22850_));
  NOR2_X1    g20414(.A1(new_n22850_), .A2(new_n12972_), .ZN(new_n22851_));
  AOI21_X1   g20415(.A1(new_n12972_), .A2(new_n22840_), .B(new_n22851_), .ZN(new_n22852_));
  AND2_X2    g20416(.A1(new_n22852_), .A2(pi0644), .Z(new_n22853_));
  AOI21_X1   g20417(.A1(new_n22849_), .A2(new_n12975_), .B(new_n22853_), .ZN(new_n22854_));
  NAND2_X1   g20418(.A1(new_n22757_), .A2(pi0644), .ZN(new_n22855_));
  NOR2_X1    g20419(.A1(new_n17611_), .A2(new_n22735_), .ZN(new_n22856_));
  AOI21_X1   g20420(.A1(new_n22759_), .A2(new_n17611_), .B(new_n22856_), .ZN(new_n22857_));
  OAI21_X1   g20421(.A1(new_n22857_), .A2(pi0644), .B(new_n22855_), .ZN(new_n22858_));
  NAND2_X1   g20422(.A1(new_n22858_), .A2(pi0715), .ZN(new_n22859_));
  OAI21_X1   g20423(.A1(new_n22854_), .A2(pi0715), .B(new_n22859_), .ZN(new_n22860_));
  NAND2_X1   g20424(.A1(new_n22849_), .A2(pi0644), .ZN(new_n22861_));
  NAND2_X1   g20425(.A1(new_n22852_), .A2(new_n12975_), .ZN(new_n22862_));
  AOI21_X1   g20426(.A1(new_n22861_), .A2(new_n22862_), .B(new_n12740_), .ZN(new_n22863_));
  OAI21_X1   g20427(.A1(new_n22757_), .A2(pi0644), .B(new_n12740_), .ZN(new_n22864_));
  AND2_X2    g20428(.A1(new_n22857_), .A2(pi0644), .Z(new_n22865_));
  OAI21_X1   g20429(.A1(new_n22865_), .A2(new_n22864_), .B(pi1160), .ZN(new_n22866_));
  OAI22_X1   g20430(.A1(new_n22860_), .A2(pi1160), .B1(new_n22863_), .B2(new_n22866_), .ZN(new_n22867_));
  OAI21_X1   g20431(.A1(new_n22849_), .A2(pi0790), .B(pi0832), .ZN(new_n22868_));
  AOI21_X1   g20432(.A1(new_n22867_), .A2(pi0790), .B(new_n22868_), .ZN(new_n22869_));
  NOR2_X1    g20433(.A1(new_n13193_), .A2(pi0190), .ZN(new_n22870_));
  AOI21_X1   g20434(.A1(new_n22870_), .A2(pi0644), .B(new_n12740_), .ZN(new_n22871_));
  NOR2_X1    g20435(.A1(new_n22870_), .A2(new_n12985_), .ZN(new_n22872_));
  INV_X1     g20436(.I(new_n22870_), .ZN(new_n22873_));
  NAND2_X1   g20437(.A1(new_n22873_), .A2(new_n12943_), .ZN(new_n22874_));
  NOR2_X1    g20438(.A1(new_n2609_), .A2(new_n10721_), .ZN(new_n22875_));
  OAI22_X1   g20439(.A1(new_n16941_), .A2(pi0190), .B1(new_n16945_), .B2(new_n13208_), .ZN(new_n22876_));
  NAND3_X1   g20440(.A1(new_n17986_), .A2(new_n10721_), .A3(pi0763), .ZN(new_n22877_));
  NAND2_X1   g20441(.A1(new_n22877_), .A2(new_n22876_), .ZN(new_n22878_));
  OAI22_X1   g20442(.A1(new_n14065_), .A2(pi0763), .B1(new_n10721_), .B2(new_n14067_), .ZN(new_n22879_));
  AOI21_X1   g20443(.A1(pi0039), .A2(new_n22879_), .B(new_n22878_), .ZN(new_n22880_));
  NAND2_X1   g20444(.A1(new_n13397_), .A2(new_n10721_), .ZN(new_n22881_));
  NAND2_X1   g20445(.A1(new_n22881_), .A2(pi0038), .ZN(new_n22882_));
  NOR2_X1    g20446(.A1(new_n13342_), .A2(new_n16945_), .ZN(new_n22883_));
  OAI22_X1   g20447(.A1(new_n22880_), .A2(pi0038), .B1(new_n22882_), .B2(new_n22883_), .ZN(new_n22884_));
  AOI21_X1   g20448(.A1(new_n22884_), .A2(new_n2609_), .B(new_n22875_), .ZN(new_n22885_));
  NOR2_X1    g20449(.A1(new_n22885_), .A2(new_n12760_), .ZN(new_n22886_));
  NOR2_X1    g20450(.A1(new_n22870_), .A2(new_n12761_), .ZN(new_n22887_));
  NOR3_X1    g20451(.A1(new_n22886_), .A2(pi0785), .A3(new_n22887_), .ZN(new_n22888_));
  AOI22_X1   g20452(.A1(new_n22886_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n22873_), .ZN(new_n22889_));
  NOR2_X1    g20453(.A1(new_n22889_), .A2(pi1155), .ZN(new_n22890_));
  AOI22_X1   g20454(.A1(new_n22886_), .A2(pi0609), .B1(new_n13357_), .B2(new_n22873_), .ZN(new_n22891_));
  NOR2_X1    g20455(.A1(new_n22891_), .A2(new_n12770_), .ZN(new_n22892_));
  NOR3_X1    g20456(.A1(new_n22892_), .A2(new_n22890_), .A3(new_n12764_), .ZN(new_n22893_));
  NOR2_X1    g20457(.A1(new_n22893_), .A2(new_n22888_), .ZN(new_n22894_));
  NAND2_X1   g20458(.A1(new_n22894_), .A2(new_n12781_), .ZN(new_n22895_));
  NOR2_X1    g20459(.A1(new_n22870_), .A2(new_n12781_), .ZN(new_n22896_));
  INV_X1     g20460(.I(new_n22896_), .ZN(new_n22897_));
  AOI21_X1   g20461(.A1(new_n22895_), .A2(new_n22897_), .B(pi1154), .ZN(new_n22898_));
  NAND2_X1   g20462(.A1(new_n22894_), .A2(pi0618), .ZN(new_n22899_));
  NAND2_X1   g20463(.A1(new_n22873_), .A2(new_n12781_), .ZN(new_n22900_));
  AOI21_X1   g20464(.A1(new_n22899_), .A2(new_n22900_), .B(new_n12785_), .ZN(new_n22901_));
  OR2_X2     g20465(.A1(new_n22901_), .A2(new_n12779_), .Z(new_n22902_));
  OAI22_X1   g20466(.A1(new_n22902_), .A2(new_n22898_), .B1(pi0781), .B2(new_n22894_), .ZN(new_n22903_));
  NAND2_X1   g20467(.A1(new_n22873_), .A2(pi0619), .ZN(new_n22904_));
  OAI21_X1   g20468(.A1(new_n22903_), .A2(pi0619), .B(new_n22904_), .ZN(new_n22905_));
  NAND2_X1   g20469(.A1(new_n22905_), .A2(new_n12791_), .ZN(new_n22906_));
  NOR2_X1    g20470(.A1(new_n22903_), .A2(new_n12793_), .ZN(new_n22907_));
  AOI21_X1   g20471(.A1(new_n12793_), .A2(new_n22873_), .B(new_n22907_), .ZN(new_n22908_));
  NOR2_X1    g20472(.A1(new_n22908_), .A2(new_n12791_), .ZN(new_n22909_));
  NOR2_X1    g20473(.A1(new_n22909_), .A2(new_n12796_), .ZN(new_n22910_));
  AOI22_X1   g20474(.A1(new_n22910_), .A2(new_n22906_), .B1(new_n12796_), .B2(new_n22903_), .ZN(new_n22911_));
  NOR2_X1    g20475(.A1(new_n22870_), .A2(new_n17504_), .ZN(new_n22912_));
  AOI21_X1   g20476(.A1(new_n22911_), .A2(new_n17504_), .B(new_n22912_), .ZN(new_n22913_));
  OAI21_X1   g20477(.A1(new_n22913_), .A2(new_n12943_), .B(new_n22874_), .ZN(new_n22914_));
  AOI21_X1   g20478(.A1(new_n22914_), .A2(new_n12985_), .B(new_n22872_), .ZN(new_n22915_));
  NAND2_X1   g20479(.A1(new_n22915_), .A2(new_n12975_), .ZN(new_n22916_));
  AOI21_X1   g20480(.A1(new_n22916_), .A2(new_n22871_), .B(pi1160), .ZN(new_n22917_));
  NAND2_X1   g20481(.A1(new_n22873_), .A2(new_n12741_), .ZN(new_n22918_));
  NOR2_X1    g20482(.A1(new_n22870_), .A2(pi0628), .ZN(new_n22919_));
  NAND2_X1   g20483(.A1(new_n22870_), .A2(new_n12869_), .ZN(new_n22920_));
  INV_X1     g20484(.I(new_n22875_), .ZN(new_n22921_));
  NAND3_X1   g20485(.A1(new_n13395_), .A2(new_n10721_), .A3(new_n22761_), .ZN(new_n22922_));
  NOR2_X1    g20486(.A1(new_n18033_), .A2(new_n10721_), .ZN(new_n22923_));
  AOI21_X1   g20487(.A1(new_n10721_), .A2(new_n14118_), .B(new_n22923_), .ZN(new_n22924_));
  AOI21_X1   g20488(.A1(new_n13399_), .A2(new_n22881_), .B(new_n22761_), .ZN(new_n22925_));
  OAI21_X1   g20489(.A1(new_n22924_), .A2(pi0038), .B(new_n22925_), .ZN(new_n22926_));
  NAND3_X1   g20490(.A1(new_n22926_), .A2(new_n2609_), .A3(new_n22922_), .ZN(new_n22927_));
  NAND2_X1   g20491(.A1(new_n22927_), .A2(new_n22921_), .ZN(new_n22928_));
  NAND2_X1   g20492(.A1(new_n22873_), .A2(pi0625), .ZN(new_n22929_));
  NAND2_X1   g20493(.A1(new_n22928_), .A2(new_n13521_), .ZN(new_n22930_));
  AOI21_X1   g20494(.A1(new_n22930_), .A2(new_n22929_), .B(pi1153), .ZN(new_n22931_));
  NAND2_X1   g20495(.A1(new_n22873_), .A2(new_n13521_), .ZN(new_n22932_));
  NAND2_X1   g20496(.A1(new_n22928_), .A2(pi0625), .ZN(new_n22933_));
  AOI21_X1   g20497(.A1(new_n22933_), .A2(new_n22932_), .B(new_n12841_), .ZN(new_n22934_));
  OR2_X2     g20498(.A1(new_n22934_), .A2(new_n12758_), .Z(new_n22935_));
  OAI22_X1   g20499(.A1(new_n22935_), .A2(new_n22931_), .B1(pi0778), .B2(new_n22928_), .ZN(new_n22936_));
  NAND2_X1   g20500(.A1(new_n22936_), .A2(new_n12870_), .ZN(new_n22937_));
  NAND2_X1   g20501(.A1(new_n22937_), .A2(new_n22920_), .ZN(new_n22938_));
  NAND2_X1   g20502(.A1(new_n22873_), .A2(new_n12887_), .ZN(new_n22939_));
  OAI21_X1   g20503(.A1(new_n22938_), .A2(new_n12887_), .B(new_n22939_), .ZN(new_n22940_));
  NAND2_X1   g20504(.A1(new_n22870_), .A2(new_n12910_), .ZN(new_n22941_));
  OAI21_X1   g20505(.A1(new_n22940_), .A2(new_n12910_), .B(new_n22941_), .ZN(new_n22942_));
  NAND2_X1   g20506(.A1(new_n22873_), .A2(new_n12817_), .ZN(new_n22943_));
  OAI21_X1   g20507(.A1(new_n22942_), .A2(new_n12817_), .B(new_n22943_), .ZN(new_n22944_));
  AOI21_X1   g20508(.A1(new_n22944_), .A2(pi0628), .B(new_n22919_), .ZN(new_n22945_));
  NOR2_X1    g20509(.A1(new_n22945_), .A2(new_n12742_), .ZN(new_n22946_));
  NOR2_X1    g20510(.A1(new_n22870_), .A2(new_n12920_), .ZN(new_n22947_));
  AOI21_X1   g20511(.A1(new_n22944_), .A2(new_n12920_), .B(new_n22947_), .ZN(new_n22948_));
  NOR2_X1    g20512(.A1(new_n22948_), .A2(pi1156), .ZN(new_n22949_));
  OAI21_X1   g20513(.A1(new_n22946_), .A2(new_n22949_), .B(pi0792), .ZN(new_n22950_));
  NAND2_X1   g20514(.A1(new_n22944_), .A2(new_n12937_), .ZN(new_n22951_));
  NAND2_X1   g20515(.A1(new_n22950_), .A2(new_n22951_), .ZN(new_n22952_));
  NAND2_X1   g20516(.A1(new_n22952_), .A2(pi0647), .ZN(new_n22953_));
  AOI21_X1   g20517(.A1(new_n22953_), .A2(new_n22918_), .B(new_n12965_), .ZN(new_n22954_));
  NAND2_X1   g20518(.A1(new_n22873_), .A2(pi0647), .ZN(new_n22955_));
  NAND2_X1   g20519(.A1(new_n22952_), .A2(new_n12741_), .ZN(new_n22956_));
  AOI21_X1   g20520(.A1(new_n22956_), .A2(new_n22955_), .B(pi1157), .ZN(new_n22957_));
  OAI21_X1   g20521(.A1(new_n22954_), .A2(new_n22957_), .B(pi0787), .ZN(new_n22958_));
  NAND2_X1   g20522(.A1(new_n22952_), .A2(new_n12972_), .ZN(new_n22959_));
  NAND2_X1   g20523(.A1(new_n22958_), .A2(new_n22959_), .ZN(new_n22960_));
  OAI21_X1   g20524(.A1(new_n22960_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n22961_));
  AOI21_X1   g20525(.A1(new_n22870_), .A2(new_n12975_), .B(pi0715), .ZN(new_n22962_));
  NAND2_X1   g20526(.A1(new_n22915_), .A2(pi0644), .ZN(new_n22963_));
  AOI21_X1   g20527(.A1(new_n22963_), .A2(new_n22962_), .B(new_n12739_), .ZN(new_n22964_));
  OAI21_X1   g20528(.A1(new_n22960_), .A2(pi0644), .B(pi0715), .ZN(new_n22965_));
  AOI22_X1   g20529(.A1(new_n22917_), .A2(new_n22961_), .B1(new_n22964_), .B2(new_n22965_), .ZN(new_n22966_));
  NOR2_X1    g20530(.A1(new_n22966_), .A2(new_n13000_), .ZN(new_n22967_));
  OR2_X2     g20531(.A1(new_n22964_), .A2(new_n12975_), .Z(new_n22968_));
  OR2_X2     g20532(.A1(new_n22917_), .A2(pi0644), .Z(new_n22969_));
  AOI21_X1   g20533(.A1(new_n22968_), .A2(new_n22969_), .B(new_n13000_), .ZN(new_n22970_));
  NAND2_X1   g20534(.A1(new_n22953_), .A2(new_n22918_), .ZN(new_n22971_));
  NAND2_X1   g20535(.A1(new_n22956_), .A2(new_n22955_), .ZN(new_n22972_));
  AOI22_X1   g20536(.A1(new_n12980_), .A2(new_n22971_), .B1(new_n22972_), .B2(new_n12982_), .ZN(new_n22973_));
  NAND2_X1   g20537(.A1(new_n22914_), .A2(new_n15608_), .ZN(new_n22974_));
  AOI21_X1   g20538(.A1(new_n22974_), .A2(new_n22973_), .B(new_n12972_), .ZN(new_n22975_));
  OAI22_X1   g20539(.A1(new_n18087_), .A2(new_n22945_), .B1(new_n22948_), .B2(new_n18088_), .ZN(new_n22976_));
  NOR2_X1    g20540(.A1(new_n22913_), .A2(new_n15821_), .ZN(new_n22977_));
  OAI21_X1   g20541(.A1(new_n22977_), .A2(new_n22976_), .B(pi0792), .ZN(new_n22978_));
  NOR2_X1    g20542(.A1(new_n22911_), .A2(pi0626), .ZN(new_n22979_));
  AOI21_X1   g20543(.A1(pi0626), .A2(new_n22870_), .B(new_n22979_), .ZN(new_n22980_));
  NAND2_X1   g20544(.A1(new_n22870_), .A2(new_n12747_), .ZN(new_n22981_));
  OAI21_X1   g20545(.A1(new_n22911_), .A2(new_n12747_), .B(new_n22981_), .ZN(new_n22982_));
  AOI22_X1   g20546(.A1(new_n22982_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n22942_), .ZN(new_n22983_));
  OAI21_X1   g20547(.A1(new_n12816_), .A2(new_n22980_), .B(new_n22983_), .ZN(new_n22984_));
  AOI21_X1   g20548(.A1(new_n22984_), .A2(pi0788), .B(new_n15340_), .ZN(new_n22985_));
  OR2_X2     g20549(.A1(new_n22936_), .A2(pi0609), .Z(new_n22986_));
  OAI21_X1   g20550(.A1(new_n13562_), .A2(new_n22736_), .B(pi0190), .ZN(new_n22987_));
  OAI21_X1   g20551(.A1(new_n18102_), .A2(pi0763), .B(new_n13566_), .ZN(new_n22988_));
  NAND2_X1   g20552(.A1(new_n22988_), .A2(new_n2627_), .ZN(new_n22989_));
  AOI21_X1   g20553(.A1(new_n22989_), .A2(new_n10721_), .B(new_n3265_), .ZN(new_n22990_));
  OAI21_X1   g20554(.A1(new_n5337_), .A2(new_n22987_), .B(new_n22990_), .ZN(new_n22991_));
  NOR2_X1    g20555(.A1(new_n14172_), .A2(new_n10721_), .ZN(new_n22992_));
  NOR2_X1    g20556(.A1(new_n14174_), .A2(pi0190), .ZN(new_n22993_));
  OAI21_X1   g20557(.A1(new_n22992_), .A2(new_n22993_), .B(pi0763), .ZN(new_n22994_));
  NAND2_X1   g20558(.A1(new_n18110_), .A2(new_n10721_), .ZN(new_n22995_));
  OAI21_X1   g20559(.A1(new_n10721_), .A2(new_n15835_), .B(new_n22995_), .ZN(new_n22996_));
  NAND2_X1   g20560(.A1(new_n22996_), .A2(new_n16945_), .ZN(new_n22997_));
  NAND3_X1   g20561(.A1(new_n22997_), .A2(new_n2627_), .A3(new_n22994_), .ZN(new_n22998_));
  NOR2_X1    g20562(.A1(new_n14182_), .A2(pi0190), .ZN(new_n22999_));
  NOR2_X1    g20563(.A1(new_n14184_), .A2(new_n10721_), .ZN(new_n23000_));
  OAI21_X1   g20564(.A1(new_n22999_), .A2(new_n23000_), .B(new_n16945_), .ZN(new_n23001_));
  NOR2_X1    g20565(.A1(new_n14187_), .A2(new_n10721_), .ZN(new_n23002_));
  NOR2_X1    g20566(.A1(new_n14189_), .A2(pi0190), .ZN(new_n23003_));
  OAI21_X1   g20567(.A1(new_n23002_), .A2(new_n23003_), .B(pi0763), .ZN(new_n23004_));
  NAND3_X1   g20568(.A1(new_n23004_), .A2(new_n23001_), .A3(pi0039), .ZN(new_n23005_));
  NAND3_X1   g20569(.A1(new_n22998_), .A2(new_n23005_), .A3(new_n3265_), .ZN(new_n23006_));
  NAND3_X1   g20570(.A1(new_n23006_), .A2(pi0699), .A3(new_n22991_), .ZN(new_n23007_));
  NAND2_X1   g20571(.A1(new_n23007_), .A2(new_n2609_), .ZN(new_n23008_));
  NOR2_X1    g20572(.A1(new_n22884_), .A2(pi0699), .ZN(new_n23009_));
  OAI21_X1   g20573(.A1(new_n23008_), .A2(new_n23009_), .B(new_n22921_), .ZN(new_n23010_));
  OR2_X2     g20574(.A1(new_n22885_), .A2(new_n13521_), .Z(new_n23011_));
  NAND2_X1   g20575(.A1(new_n23010_), .A2(new_n13521_), .ZN(new_n23012_));
  AOI21_X1   g20576(.A1(new_n23012_), .A2(new_n23011_), .B(pi1153), .ZN(new_n23013_));
  NOR3_X1    g20577(.A1(new_n23013_), .A2(pi0608), .A3(new_n22934_), .ZN(new_n23014_));
  NOR2_X1    g20578(.A1(new_n22885_), .A2(pi0625), .ZN(new_n23015_));
  AOI21_X1   g20579(.A1(new_n23010_), .A2(pi0625), .B(new_n23015_), .ZN(new_n23016_));
  NOR2_X1    g20580(.A1(new_n23016_), .A2(new_n12841_), .ZN(new_n23017_));
  NOR3_X1    g20581(.A1(new_n23017_), .A2(new_n13560_), .A3(new_n22931_), .ZN(new_n23018_));
  NOR3_X1    g20582(.A1(new_n23018_), .A2(new_n23014_), .A3(new_n12758_), .ZN(new_n23019_));
  AOI21_X1   g20583(.A1(new_n12758_), .A2(new_n23010_), .B(new_n23019_), .ZN(new_n23020_));
  OAI21_X1   g20584(.A1(new_n23020_), .A2(new_n12766_), .B(new_n22986_), .ZN(new_n23021_));
  AOI21_X1   g20585(.A1(new_n23021_), .A2(pi1155), .B(new_n22890_), .ZN(new_n23022_));
  NOR2_X1    g20586(.A1(new_n23020_), .A2(pi0609), .ZN(new_n23023_));
  NOR2_X1    g20587(.A1(new_n22936_), .A2(new_n12766_), .ZN(new_n23024_));
  OAI21_X1   g20588(.A1(new_n23023_), .A2(new_n23024_), .B(new_n12770_), .ZN(new_n23025_));
  NOR2_X1    g20589(.A1(new_n22892_), .A2(pi0660), .ZN(new_n23026_));
  AOI22_X1   g20590(.A1(new_n23022_), .A2(pi0660), .B1(new_n23025_), .B2(new_n23026_), .ZN(new_n23027_));
  AND2_X2    g20591(.A1(new_n23027_), .A2(pi0785), .Z(new_n23028_));
  NOR2_X1    g20592(.A1(new_n23020_), .A2(pi0785), .ZN(new_n23029_));
  NOR2_X1    g20593(.A1(new_n23028_), .A2(new_n23029_), .ZN(new_n23030_));
  NOR2_X1    g20594(.A1(new_n23030_), .A2(pi0781), .ZN(new_n23031_));
  NOR2_X1    g20595(.A1(new_n22938_), .A2(pi0618), .ZN(new_n23032_));
  INV_X1     g20596(.I(new_n23032_), .ZN(new_n23033_));
  OAI21_X1   g20597(.A1(new_n23028_), .A2(new_n23029_), .B(pi0618), .ZN(new_n23034_));
  AOI21_X1   g20598(.A1(new_n23034_), .A2(new_n23033_), .B(new_n12785_), .ZN(new_n23035_));
  NOR3_X1    g20599(.A1(new_n23035_), .A2(new_n12880_), .A3(new_n22898_), .ZN(new_n23036_));
  OAI21_X1   g20600(.A1(new_n23028_), .A2(new_n23029_), .B(new_n12781_), .ZN(new_n23037_));
  NAND3_X1   g20601(.A1(new_n22937_), .A2(pi0618), .A3(new_n22920_), .ZN(new_n23038_));
  AOI21_X1   g20602(.A1(new_n23037_), .A2(new_n23038_), .B(pi1154), .ZN(new_n23039_));
  NOR3_X1    g20603(.A1(new_n23039_), .A2(pi0627), .A3(new_n22901_), .ZN(new_n23040_));
  NOR3_X1    g20604(.A1(new_n23036_), .A2(new_n23040_), .A3(new_n12779_), .ZN(new_n23041_));
  OAI21_X1   g20605(.A1(new_n23041_), .A2(new_n23031_), .B(new_n12796_), .ZN(new_n23042_));
  NAND2_X1   g20606(.A1(new_n23042_), .A2(new_n12819_), .ZN(new_n23043_));
  NAND2_X1   g20607(.A1(new_n22940_), .A2(pi0619), .ZN(new_n23044_));
  OAI21_X1   g20608(.A1(new_n23041_), .A2(new_n23031_), .B(new_n12793_), .ZN(new_n23045_));
  AOI21_X1   g20609(.A1(new_n23045_), .A2(new_n23044_), .B(pi1159), .ZN(new_n23046_));
  NOR3_X1    g20610(.A1(new_n23046_), .A2(pi0648), .A3(new_n22909_), .ZN(new_n23047_));
  INV_X1     g20611(.I(new_n22906_), .ZN(new_n23048_));
  OAI21_X1   g20612(.A1(new_n23041_), .A2(new_n23031_), .B(pi0619), .ZN(new_n23049_));
  NAND2_X1   g20613(.A1(new_n22940_), .A2(new_n12793_), .ZN(new_n23050_));
  AOI21_X1   g20614(.A1(new_n23049_), .A2(new_n23050_), .B(new_n12791_), .ZN(new_n23051_));
  NOR3_X1    g20615(.A1(new_n23051_), .A2(new_n12895_), .A3(new_n23048_), .ZN(new_n23052_));
  NOR3_X1    g20616(.A1(new_n23047_), .A2(new_n23052_), .A3(new_n12796_), .ZN(new_n23053_));
  OAI21_X1   g20617(.A1(new_n23053_), .A2(new_n23043_), .B(new_n22985_), .ZN(new_n23054_));
  AOI21_X1   g20618(.A1(new_n23054_), .A2(new_n22978_), .B(new_n15341_), .ZN(new_n23055_));
  NOR3_X1    g20619(.A1(new_n22970_), .A2(new_n22975_), .A3(new_n23055_), .ZN(new_n23056_));
  OAI21_X1   g20620(.A1(new_n23056_), .A2(new_n22967_), .B(new_n6643_), .ZN(new_n23057_));
  AOI21_X1   g20621(.A1(po1038), .A2(new_n10721_), .B(pi0832), .ZN(new_n23058_));
  AOI21_X1   g20622(.A1(new_n23057_), .A2(new_n23058_), .B(new_n22869_), .ZN(po0347));
  NOR2_X1    g20623(.A1(new_n3042_), .A2(pi0191), .ZN(new_n23060_));
  NOR2_X1    g20624(.A1(new_n13340_), .A2(new_n16996_), .ZN(new_n23061_));
  NOR2_X1    g20625(.A1(new_n23061_), .A2(new_n23060_), .ZN(new_n23062_));
  NOR3_X1    g20626(.A1(new_n23062_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n23063_));
  INV_X1     g20627(.I(new_n23061_), .ZN(new_n23064_));
  NOR2_X1    g20628(.A1(new_n23064_), .A2(new_n13354_), .ZN(new_n23065_));
  NOR3_X1    g20629(.A1(new_n23065_), .A2(new_n12762_), .A3(new_n23062_), .ZN(new_n23066_));
  NOR2_X1    g20630(.A1(new_n23066_), .A2(new_n12770_), .ZN(new_n23067_));
  NOR3_X1    g20631(.A1(new_n23065_), .A2(pi1155), .A3(new_n23060_), .ZN(new_n23068_));
  NOR3_X1    g20632(.A1(new_n23067_), .A2(new_n12764_), .A3(new_n23068_), .ZN(new_n23069_));
  NOR2_X1    g20633(.A1(new_n23069_), .A2(new_n23063_), .ZN(new_n23070_));
  NOR2_X1    g20634(.A1(new_n23070_), .A2(pi0781), .ZN(new_n23071_));
  INV_X1     g20635(.I(new_n23070_), .ZN(new_n23072_));
  AOI21_X1   g20636(.A1(new_n23072_), .A2(new_n12783_), .B(pi1154), .ZN(new_n23073_));
  AOI21_X1   g20637(.A1(new_n23072_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n23074_));
  NOR3_X1    g20638(.A1(new_n23073_), .A2(new_n23074_), .A3(new_n12779_), .ZN(new_n23075_));
  NOR2_X1    g20639(.A1(new_n23075_), .A2(new_n23071_), .ZN(new_n23076_));
  NOR2_X1    g20640(.A1(new_n23076_), .A2(new_n17229_), .ZN(new_n23077_));
  NOR2_X1    g20641(.A1(new_n23077_), .A2(pi1159), .ZN(new_n23078_));
  OAI21_X1   g20642(.A1(new_n23076_), .A2(new_n17232_), .B(pi1159), .ZN(new_n23079_));
  NAND2_X1   g20643(.A1(new_n23079_), .A2(pi0789), .ZN(new_n23080_));
  OAI22_X1   g20644(.A1(new_n23080_), .A2(new_n23078_), .B1(pi0789), .B2(new_n23076_), .ZN(new_n23081_));
  INV_X1     g20645(.I(new_n23060_), .ZN(new_n23082_));
  NAND2_X1   g20646(.A1(new_n12818_), .A2(new_n23082_), .ZN(new_n23083_));
  OAI21_X1   g20647(.A1(new_n23081_), .A2(new_n12818_), .B(new_n23083_), .ZN(new_n23084_));
  AOI21_X1   g20648(.A1(new_n12826_), .A2(pi0729), .B(new_n23060_), .ZN(new_n23085_));
  INV_X1     g20649(.I(pi0729), .ZN(new_n23086_));
  NOR2_X1    g20650(.A1(new_n12834_), .A2(new_n23086_), .ZN(new_n23087_));
  INV_X1     g20651(.I(new_n23087_), .ZN(new_n23088_));
  NOR2_X1    g20652(.A1(new_n23060_), .A2(pi1153), .ZN(new_n23089_));
  NAND2_X1   g20653(.A1(new_n23088_), .A2(new_n23089_), .ZN(new_n23090_));
  NOR2_X1    g20654(.A1(new_n23087_), .A2(new_n23085_), .ZN(new_n23091_));
  NOR2_X1    g20655(.A1(new_n23091_), .A2(new_n12841_), .ZN(new_n23092_));
  INV_X1     g20656(.I(new_n23092_), .ZN(new_n23093_));
  NAND3_X1   g20657(.A1(new_n23093_), .A2(pi0778), .A3(new_n23090_), .ZN(new_n23094_));
  OAI21_X1   g20658(.A1(pi0778), .A2(new_n23085_), .B(new_n23094_), .ZN(new_n23095_));
  NAND2_X1   g20659(.A1(new_n23095_), .A2(new_n17187_), .ZN(new_n23096_));
  NOR2_X1    g20660(.A1(new_n23096_), .A2(new_n12889_), .ZN(new_n23097_));
  INV_X1     g20661(.I(new_n23097_), .ZN(new_n23098_));
  NOR2_X1    g20662(.A1(new_n23098_), .A2(new_n12912_), .ZN(new_n23099_));
  INV_X1     g20663(.I(new_n23099_), .ZN(new_n23100_));
  NOR2_X1    g20664(.A1(new_n23100_), .A2(new_n17884_), .ZN(new_n23101_));
  INV_X1     g20665(.I(new_n23101_), .ZN(new_n23102_));
  OAI22_X1   g20666(.A1(new_n23084_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n23102_), .ZN(new_n23103_));
  NAND2_X1   g20667(.A1(new_n23103_), .A2(new_n12919_), .ZN(new_n23104_));
  OAI22_X1   g20668(.A1(new_n23084_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n23102_), .ZN(new_n23105_));
  NAND2_X1   g20669(.A1(new_n23105_), .A2(pi0629), .ZN(new_n23106_));
  AOI21_X1   g20670(.A1(new_n23104_), .A2(new_n23106_), .B(new_n12937_), .ZN(new_n23107_));
  INV_X1     g20671(.I(new_n23068_), .ZN(new_n23108_));
  NOR2_X1    g20672(.A1(new_n23085_), .A2(new_n12754_), .ZN(new_n23109_));
  NOR3_X1    g20673(.A1(new_n23109_), .A2(new_n23060_), .A3(new_n23061_), .ZN(new_n23110_));
  NAND2_X1   g20674(.A1(new_n23110_), .A2(new_n12758_), .ZN(new_n23111_));
  NAND2_X1   g20675(.A1(new_n23109_), .A2(pi0625), .ZN(new_n23112_));
  NAND3_X1   g20676(.A1(new_n23112_), .A2(pi1153), .A3(new_n23062_), .ZN(new_n23113_));
  NAND3_X1   g20677(.A1(new_n23090_), .A2(pi0608), .A3(new_n23113_), .ZN(new_n23114_));
  INV_X1     g20678(.I(new_n23112_), .ZN(new_n23115_));
  OAI21_X1   g20679(.A1(new_n23115_), .A2(new_n23110_), .B(new_n23089_), .ZN(new_n23116_));
  NAND3_X1   g20680(.A1(new_n23093_), .A2(new_n13560_), .A3(new_n23116_), .ZN(new_n23117_));
  NAND3_X1   g20681(.A1(new_n23117_), .A2(pi0778), .A3(new_n23114_), .ZN(new_n23118_));
  AOI21_X1   g20682(.A1(new_n23118_), .A2(new_n23111_), .B(new_n12766_), .ZN(new_n23119_));
  NOR2_X1    g20683(.A1(new_n23095_), .A2(pi0609), .ZN(new_n23120_));
  OAI21_X1   g20684(.A1(new_n23120_), .A2(new_n23119_), .B(pi1155), .ZN(new_n23121_));
  NAND3_X1   g20685(.A1(new_n23121_), .A2(pi0660), .A3(new_n23108_), .ZN(new_n23122_));
  NAND2_X1   g20686(.A1(new_n23118_), .A2(new_n23111_), .ZN(new_n23123_));
  NOR2_X1    g20687(.A1(new_n23095_), .A2(new_n12766_), .ZN(new_n23124_));
  AOI21_X1   g20688(.A1(new_n23123_), .A2(new_n12766_), .B(new_n23124_), .ZN(new_n23125_));
  NOR2_X1    g20689(.A1(new_n23067_), .A2(pi0660), .ZN(new_n23126_));
  OAI21_X1   g20690(.A1(new_n23125_), .A2(pi1155), .B(new_n23126_), .ZN(new_n23127_));
  NAND3_X1   g20691(.A1(new_n23127_), .A2(new_n23122_), .A3(pi0785), .ZN(new_n23128_));
  NAND2_X1   g20692(.A1(new_n23123_), .A2(new_n12764_), .ZN(new_n23129_));
  NAND2_X1   g20693(.A1(new_n23128_), .A2(new_n23129_), .ZN(new_n23130_));
  NAND2_X1   g20694(.A1(new_n23130_), .A2(new_n12781_), .ZN(new_n23131_));
  NAND2_X1   g20695(.A1(new_n23096_), .A2(pi0618), .ZN(new_n23132_));
  AOI21_X1   g20696(.A1(new_n23131_), .A2(new_n23132_), .B(pi1154), .ZN(new_n23133_));
  NOR3_X1    g20697(.A1(new_n23133_), .A2(pi0627), .A3(new_n23074_), .ZN(new_n23134_));
  NAND2_X1   g20698(.A1(new_n23096_), .A2(new_n12781_), .ZN(new_n23135_));
  NAND2_X1   g20699(.A1(new_n23130_), .A2(pi0618), .ZN(new_n23136_));
  AOI21_X1   g20700(.A1(new_n23136_), .A2(new_n23135_), .B(new_n12785_), .ZN(new_n23137_));
  NOR3_X1    g20701(.A1(new_n23137_), .A2(new_n12880_), .A3(new_n23073_), .ZN(new_n23138_));
  OR3_X2     g20702(.A1(new_n23134_), .A2(new_n23138_), .A3(new_n12779_), .Z(new_n23139_));
  NAND2_X1   g20703(.A1(new_n23130_), .A2(new_n12779_), .ZN(new_n23140_));
  NAND2_X1   g20704(.A1(new_n23139_), .A2(new_n23140_), .ZN(new_n23141_));
  AOI21_X1   g20705(.A1(new_n23141_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n23142_));
  NAND2_X1   g20706(.A1(new_n23098_), .A2(new_n12793_), .ZN(new_n23143_));
  NAND2_X1   g20707(.A1(new_n23141_), .A2(pi0619), .ZN(new_n23144_));
  AOI21_X1   g20708(.A1(new_n23144_), .A2(new_n23143_), .B(new_n12791_), .ZN(new_n23145_));
  NOR3_X1    g20709(.A1(new_n23145_), .A2(new_n12895_), .A3(new_n23078_), .ZN(new_n23146_));
  AOI21_X1   g20710(.A1(new_n23139_), .A2(new_n23140_), .B(pi0619), .ZN(new_n23147_));
  NOR2_X1    g20711(.A1(new_n23097_), .A2(new_n12793_), .ZN(new_n23148_));
  OAI21_X1   g20712(.A1(new_n23147_), .A2(new_n23148_), .B(new_n12791_), .ZN(new_n23149_));
  NAND3_X1   g20713(.A1(new_n23149_), .A2(new_n12895_), .A3(new_n23079_), .ZN(new_n23150_));
  NAND2_X1   g20714(.A1(new_n23150_), .A2(pi0789), .ZN(new_n23151_));
  OAI21_X1   g20715(.A1(new_n23151_), .A2(new_n23146_), .B(new_n23142_), .ZN(new_n23152_));
  NAND2_X1   g20716(.A1(new_n23060_), .A2(pi0626), .ZN(new_n23153_));
  NAND2_X1   g20717(.A1(new_n23081_), .A2(new_n12747_), .ZN(new_n23154_));
  AOI21_X1   g20718(.A1(new_n23154_), .A2(new_n23153_), .B(new_n12816_), .ZN(new_n23155_));
  NOR2_X1    g20719(.A1(new_n23082_), .A2(pi0626), .ZN(new_n23156_));
  AOI21_X1   g20720(.A1(new_n23081_), .A2(pi0626), .B(new_n23156_), .ZN(new_n23157_));
  OAI22_X1   g20721(.A1(new_n23157_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n23100_), .ZN(new_n23158_));
  OAI21_X1   g20722(.A1(new_n23158_), .A2(new_n23155_), .B(pi0788), .ZN(new_n23159_));
  AOI21_X1   g20723(.A1(new_n23152_), .A2(new_n23159_), .B(new_n15340_), .ZN(new_n23160_));
  OR2_X2     g20724(.A1(new_n23160_), .A2(new_n23107_), .Z(new_n23161_));
  NAND2_X1   g20725(.A1(new_n23084_), .A2(new_n13384_), .ZN(new_n23162_));
  NAND2_X1   g20726(.A1(new_n12943_), .A2(new_n23082_), .ZN(new_n23163_));
  AOI21_X1   g20727(.A1(new_n23162_), .A2(new_n23163_), .B(new_n17212_), .ZN(new_n23164_));
  NOR2_X1    g20728(.A1(new_n23102_), .A2(new_n12953_), .ZN(new_n23165_));
  NOR2_X1    g20729(.A1(new_n23165_), .A2(pi0647), .ZN(new_n23166_));
  NOR2_X1    g20730(.A1(new_n23060_), .A2(new_n12741_), .ZN(new_n23167_));
  OAI21_X1   g20731(.A1(new_n23166_), .A2(new_n23167_), .B(new_n12965_), .ZN(new_n23168_));
  NOR2_X1    g20732(.A1(new_n23082_), .A2(pi0647), .ZN(new_n23169_));
  AOI21_X1   g20733(.A1(new_n23165_), .A2(pi0647), .B(new_n23169_), .ZN(new_n23170_));
  INV_X1     g20734(.I(new_n23170_), .ZN(new_n23171_));
  OAI22_X1   g20735(.A1(new_n23168_), .A2(new_n12981_), .B1(new_n23171_), .B2(new_n15576_), .ZN(new_n23172_));
  NOR2_X1    g20736(.A1(new_n23172_), .A2(new_n23164_), .ZN(new_n23173_));
  OAI22_X1   g20737(.A1(new_n23161_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n23173_), .ZN(new_n23174_));
  OAI21_X1   g20738(.A1(new_n12965_), .A2(new_n23171_), .B(new_n23168_), .ZN(new_n23175_));
  NOR2_X1    g20739(.A1(new_n23175_), .A2(new_n12972_), .ZN(new_n23176_));
  AOI21_X1   g20740(.A1(new_n12972_), .A2(new_n23165_), .B(new_n23176_), .ZN(new_n23177_));
  AND2_X2    g20741(.A1(new_n23177_), .A2(pi0644), .Z(new_n23178_));
  AOI21_X1   g20742(.A1(new_n23174_), .A2(new_n12975_), .B(new_n23178_), .ZN(new_n23179_));
  NAND2_X1   g20743(.A1(new_n23082_), .A2(pi0644), .ZN(new_n23180_));
  NOR2_X1    g20744(.A1(new_n17611_), .A2(new_n23060_), .ZN(new_n23181_));
  AOI21_X1   g20745(.A1(new_n23084_), .A2(new_n17611_), .B(new_n23181_), .ZN(new_n23182_));
  OAI21_X1   g20746(.A1(new_n23182_), .A2(pi0644), .B(new_n23180_), .ZN(new_n23183_));
  NAND2_X1   g20747(.A1(new_n23183_), .A2(pi0715), .ZN(new_n23184_));
  OAI21_X1   g20748(.A1(new_n23179_), .A2(pi0715), .B(new_n23184_), .ZN(new_n23185_));
  NAND2_X1   g20749(.A1(new_n23174_), .A2(pi0644), .ZN(new_n23186_));
  NAND2_X1   g20750(.A1(new_n23177_), .A2(new_n12975_), .ZN(new_n23187_));
  AOI21_X1   g20751(.A1(new_n23186_), .A2(new_n23187_), .B(new_n12740_), .ZN(new_n23188_));
  OAI21_X1   g20752(.A1(new_n23082_), .A2(pi0644), .B(new_n12740_), .ZN(new_n23189_));
  AND2_X2    g20753(.A1(new_n23182_), .A2(pi0644), .Z(new_n23190_));
  OAI21_X1   g20754(.A1(new_n23190_), .A2(new_n23189_), .B(pi1160), .ZN(new_n23191_));
  OAI22_X1   g20755(.A1(new_n23185_), .A2(pi1160), .B1(new_n23188_), .B2(new_n23191_), .ZN(new_n23192_));
  OAI21_X1   g20756(.A1(new_n23174_), .A2(pi0790), .B(pi0832), .ZN(new_n23193_));
  AOI21_X1   g20757(.A1(new_n23192_), .A2(pi0790), .B(new_n23193_), .ZN(new_n23194_));
  NOR2_X1    g20758(.A1(new_n13193_), .A2(pi0191), .ZN(new_n23195_));
  AOI21_X1   g20759(.A1(new_n23195_), .A2(pi0644), .B(new_n12740_), .ZN(new_n23196_));
  NOR2_X1    g20760(.A1(new_n23195_), .A2(new_n12985_), .ZN(new_n23197_));
  INV_X1     g20761(.I(new_n23195_), .ZN(new_n23198_));
  NAND2_X1   g20762(.A1(new_n23198_), .A2(new_n12943_), .ZN(new_n23199_));
  NOR2_X1    g20763(.A1(new_n2609_), .A2(new_n12704_), .ZN(new_n23200_));
  OAI22_X1   g20764(.A1(new_n16992_), .A2(pi0191), .B1(new_n16996_), .B2(new_n13208_), .ZN(new_n23201_));
  NAND3_X1   g20765(.A1(new_n17986_), .A2(new_n12704_), .A3(pi0746), .ZN(new_n23202_));
  NAND2_X1   g20766(.A1(new_n23202_), .A2(new_n23201_), .ZN(new_n23203_));
  OAI22_X1   g20767(.A1(new_n14065_), .A2(pi0746), .B1(new_n12704_), .B2(new_n14067_), .ZN(new_n23204_));
  AOI21_X1   g20768(.A1(pi0039), .A2(new_n23204_), .B(new_n23203_), .ZN(new_n23205_));
  NAND2_X1   g20769(.A1(new_n13397_), .A2(new_n12704_), .ZN(new_n23206_));
  NAND2_X1   g20770(.A1(new_n23206_), .A2(pi0038), .ZN(new_n23207_));
  NOR2_X1    g20771(.A1(new_n13342_), .A2(new_n16996_), .ZN(new_n23208_));
  OAI22_X1   g20772(.A1(new_n23205_), .A2(pi0038), .B1(new_n23207_), .B2(new_n23208_), .ZN(new_n23209_));
  AOI21_X1   g20773(.A1(new_n23209_), .A2(new_n2609_), .B(new_n23200_), .ZN(new_n23210_));
  NOR2_X1    g20774(.A1(new_n23210_), .A2(new_n12760_), .ZN(new_n23211_));
  NOR2_X1    g20775(.A1(new_n23195_), .A2(new_n12761_), .ZN(new_n23212_));
  NOR3_X1    g20776(.A1(new_n23211_), .A2(pi0785), .A3(new_n23212_), .ZN(new_n23213_));
  AOI22_X1   g20777(.A1(new_n23211_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n23198_), .ZN(new_n23214_));
  NOR2_X1    g20778(.A1(new_n23214_), .A2(pi1155), .ZN(new_n23215_));
  AOI22_X1   g20779(.A1(new_n23211_), .A2(pi0609), .B1(new_n13357_), .B2(new_n23198_), .ZN(new_n23216_));
  NOR2_X1    g20780(.A1(new_n23216_), .A2(new_n12770_), .ZN(new_n23217_));
  NOR3_X1    g20781(.A1(new_n23217_), .A2(new_n23215_), .A3(new_n12764_), .ZN(new_n23218_));
  NOR2_X1    g20782(.A1(new_n23218_), .A2(new_n23213_), .ZN(new_n23219_));
  NAND2_X1   g20783(.A1(new_n23219_), .A2(new_n12781_), .ZN(new_n23220_));
  NOR2_X1    g20784(.A1(new_n23195_), .A2(new_n12781_), .ZN(new_n23221_));
  INV_X1     g20785(.I(new_n23221_), .ZN(new_n23222_));
  AOI21_X1   g20786(.A1(new_n23220_), .A2(new_n23222_), .B(pi1154), .ZN(new_n23223_));
  NAND2_X1   g20787(.A1(new_n23219_), .A2(pi0618), .ZN(new_n23224_));
  NAND2_X1   g20788(.A1(new_n23198_), .A2(new_n12781_), .ZN(new_n23225_));
  AOI21_X1   g20789(.A1(new_n23224_), .A2(new_n23225_), .B(new_n12785_), .ZN(new_n23226_));
  OR2_X2     g20790(.A1(new_n23226_), .A2(new_n12779_), .Z(new_n23227_));
  OAI22_X1   g20791(.A1(new_n23227_), .A2(new_n23223_), .B1(pi0781), .B2(new_n23219_), .ZN(new_n23228_));
  NAND2_X1   g20792(.A1(new_n23198_), .A2(pi0619), .ZN(new_n23229_));
  OAI21_X1   g20793(.A1(new_n23228_), .A2(pi0619), .B(new_n23229_), .ZN(new_n23230_));
  NAND2_X1   g20794(.A1(new_n23230_), .A2(new_n12791_), .ZN(new_n23231_));
  NOR2_X1    g20795(.A1(new_n23228_), .A2(new_n12793_), .ZN(new_n23232_));
  AOI21_X1   g20796(.A1(new_n12793_), .A2(new_n23198_), .B(new_n23232_), .ZN(new_n23233_));
  NOR2_X1    g20797(.A1(new_n23233_), .A2(new_n12791_), .ZN(new_n23234_));
  NOR2_X1    g20798(.A1(new_n23234_), .A2(new_n12796_), .ZN(new_n23235_));
  AOI22_X1   g20799(.A1(new_n23235_), .A2(new_n23231_), .B1(new_n12796_), .B2(new_n23228_), .ZN(new_n23236_));
  NOR2_X1    g20800(.A1(new_n23195_), .A2(new_n17504_), .ZN(new_n23237_));
  AOI21_X1   g20801(.A1(new_n23236_), .A2(new_n17504_), .B(new_n23237_), .ZN(new_n23238_));
  OAI21_X1   g20802(.A1(new_n23238_), .A2(new_n12943_), .B(new_n23199_), .ZN(new_n23239_));
  AOI21_X1   g20803(.A1(new_n23239_), .A2(new_n12985_), .B(new_n23197_), .ZN(new_n23240_));
  NAND2_X1   g20804(.A1(new_n23240_), .A2(new_n12975_), .ZN(new_n23241_));
  AOI21_X1   g20805(.A1(new_n23241_), .A2(new_n23196_), .B(pi1160), .ZN(new_n23242_));
  NAND2_X1   g20806(.A1(new_n23198_), .A2(new_n12741_), .ZN(new_n23243_));
  NOR2_X1    g20807(.A1(new_n23195_), .A2(pi0628), .ZN(new_n23244_));
  NAND2_X1   g20808(.A1(new_n23195_), .A2(new_n12869_), .ZN(new_n23245_));
  INV_X1     g20809(.I(new_n23200_), .ZN(new_n23246_));
  NAND3_X1   g20810(.A1(new_n13395_), .A2(new_n12704_), .A3(new_n23086_), .ZN(new_n23247_));
  NOR2_X1    g20811(.A1(new_n18033_), .A2(new_n12704_), .ZN(new_n23248_));
  AOI21_X1   g20812(.A1(new_n12704_), .A2(new_n14118_), .B(new_n23248_), .ZN(new_n23249_));
  AOI21_X1   g20813(.A1(new_n13399_), .A2(new_n23206_), .B(new_n23086_), .ZN(new_n23250_));
  OAI21_X1   g20814(.A1(new_n23249_), .A2(pi0038), .B(new_n23250_), .ZN(new_n23251_));
  NAND3_X1   g20815(.A1(new_n23251_), .A2(new_n2609_), .A3(new_n23247_), .ZN(new_n23252_));
  NAND2_X1   g20816(.A1(new_n23252_), .A2(new_n23246_), .ZN(new_n23253_));
  NAND2_X1   g20817(.A1(new_n23198_), .A2(pi0625), .ZN(new_n23254_));
  NAND2_X1   g20818(.A1(new_n23253_), .A2(new_n13521_), .ZN(new_n23255_));
  AOI21_X1   g20819(.A1(new_n23255_), .A2(new_n23254_), .B(pi1153), .ZN(new_n23256_));
  NAND2_X1   g20820(.A1(new_n23198_), .A2(new_n13521_), .ZN(new_n23257_));
  NAND2_X1   g20821(.A1(new_n23253_), .A2(pi0625), .ZN(new_n23258_));
  AOI21_X1   g20822(.A1(new_n23258_), .A2(new_n23257_), .B(new_n12841_), .ZN(new_n23259_));
  OR2_X2     g20823(.A1(new_n23259_), .A2(new_n12758_), .Z(new_n23260_));
  OAI22_X1   g20824(.A1(new_n23260_), .A2(new_n23256_), .B1(pi0778), .B2(new_n23253_), .ZN(new_n23261_));
  NAND2_X1   g20825(.A1(new_n23261_), .A2(new_n12870_), .ZN(new_n23262_));
  NAND2_X1   g20826(.A1(new_n23262_), .A2(new_n23245_), .ZN(new_n23263_));
  NAND2_X1   g20827(.A1(new_n23198_), .A2(new_n12887_), .ZN(new_n23264_));
  OAI21_X1   g20828(.A1(new_n23263_), .A2(new_n12887_), .B(new_n23264_), .ZN(new_n23265_));
  NAND2_X1   g20829(.A1(new_n23195_), .A2(new_n12910_), .ZN(new_n23266_));
  OAI21_X1   g20830(.A1(new_n23265_), .A2(new_n12910_), .B(new_n23266_), .ZN(new_n23267_));
  NAND2_X1   g20831(.A1(new_n23198_), .A2(new_n12817_), .ZN(new_n23268_));
  OAI21_X1   g20832(.A1(new_n23267_), .A2(new_n12817_), .B(new_n23268_), .ZN(new_n23269_));
  AOI21_X1   g20833(.A1(new_n23269_), .A2(pi0628), .B(new_n23244_), .ZN(new_n23270_));
  NOR2_X1    g20834(.A1(new_n23270_), .A2(new_n12742_), .ZN(new_n23271_));
  NOR2_X1    g20835(.A1(new_n23195_), .A2(new_n12920_), .ZN(new_n23272_));
  AOI21_X1   g20836(.A1(new_n23269_), .A2(new_n12920_), .B(new_n23272_), .ZN(new_n23273_));
  NOR2_X1    g20837(.A1(new_n23273_), .A2(pi1156), .ZN(new_n23274_));
  OAI21_X1   g20838(.A1(new_n23271_), .A2(new_n23274_), .B(pi0792), .ZN(new_n23275_));
  NAND2_X1   g20839(.A1(new_n23269_), .A2(new_n12937_), .ZN(new_n23276_));
  NAND2_X1   g20840(.A1(new_n23275_), .A2(new_n23276_), .ZN(new_n23277_));
  NAND2_X1   g20841(.A1(new_n23277_), .A2(pi0647), .ZN(new_n23278_));
  AOI21_X1   g20842(.A1(new_n23278_), .A2(new_n23243_), .B(new_n12965_), .ZN(new_n23279_));
  NAND2_X1   g20843(.A1(new_n23198_), .A2(pi0647), .ZN(new_n23280_));
  NAND2_X1   g20844(.A1(new_n23277_), .A2(new_n12741_), .ZN(new_n23281_));
  AOI21_X1   g20845(.A1(new_n23281_), .A2(new_n23280_), .B(pi1157), .ZN(new_n23282_));
  OAI21_X1   g20846(.A1(new_n23279_), .A2(new_n23282_), .B(pi0787), .ZN(new_n23283_));
  NAND2_X1   g20847(.A1(new_n23277_), .A2(new_n12972_), .ZN(new_n23284_));
  NAND2_X1   g20848(.A1(new_n23283_), .A2(new_n23284_), .ZN(new_n23285_));
  OAI21_X1   g20849(.A1(new_n23285_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n23286_));
  AOI21_X1   g20850(.A1(new_n23195_), .A2(new_n12975_), .B(pi0715), .ZN(new_n23287_));
  NAND2_X1   g20851(.A1(new_n23240_), .A2(pi0644), .ZN(new_n23288_));
  AOI21_X1   g20852(.A1(new_n23288_), .A2(new_n23287_), .B(new_n12739_), .ZN(new_n23289_));
  OAI21_X1   g20853(.A1(new_n23285_), .A2(pi0644), .B(pi0715), .ZN(new_n23290_));
  AOI22_X1   g20854(.A1(new_n23242_), .A2(new_n23286_), .B1(new_n23289_), .B2(new_n23290_), .ZN(new_n23291_));
  NOR2_X1    g20855(.A1(new_n23291_), .A2(new_n13000_), .ZN(new_n23292_));
  OR2_X2     g20856(.A1(new_n23289_), .A2(new_n12975_), .Z(new_n23293_));
  OR2_X2     g20857(.A1(new_n23242_), .A2(pi0644), .Z(new_n23294_));
  AOI21_X1   g20858(.A1(new_n23293_), .A2(new_n23294_), .B(new_n13000_), .ZN(new_n23295_));
  NAND2_X1   g20859(.A1(new_n23278_), .A2(new_n23243_), .ZN(new_n23296_));
  NAND2_X1   g20860(.A1(new_n23281_), .A2(new_n23280_), .ZN(new_n23297_));
  AOI22_X1   g20861(.A1(new_n12980_), .A2(new_n23296_), .B1(new_n23297_), .B2(new_n12982_), .ZN(new_n23298_));
  NAND2_X1   g20862(.A1(new_n23239_), .A2(new_n15608_), .ZN(new_n23299_));
  AOI21_X1   g20863(.A1(new_n23299_), .A2(new_n23298_), .B(new_n12972_), .ZN(new_n23300_));
  OAI22_X1   g20864(.A1(new_n18087_), .A2(new_n23270_), .B1(new_n23273_), .B2(new_n18088_), .ZN(new_n23301_));
  NOR2_X1    g20865(.A1(new_n23238_), .A2(new_n15821_), .ZN(new_n23302_));
  OAI21_X1   g20866(.A1(new_n23302_), .A2(new_n23301_), .B(pi0792), .ZN(new_n23303_));
  NOR2_X1    g20867(.A1(new_n23236_), .A2(pi0626), .ZN(new_n23304_));
  AOI21_X1   g20868(.A1(pi0626), .A2(new_n23195_), .B(new_n23304_), .ZN(new_n23305_));
  NAND2_X1   g20869(.A1(new_n23195_), .A2(new_n12747_), .ZN(new_n23306_));
  OAI21_X1   g20870(.A1(new_n23236_), .A2(new_n12747_), .B(new_n23306_), .ZN(new_n23307_));
  AOI22_X1   g20871(.A1(new_n23307_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n23267_), .ZN(new_n23308_));
  OAI21_X1   g20872(.A1(new_n12816_), .A2(new_n23305_), .B(new_n23308_), .ZN(new_n23309_));
  AOI21_X1   g20873(.A1(new_n23309_), .A2(pi0788), .B(new_n15340_), .ZN(new_n23310_));
  OR2_X2     g20874(.A1(new_n23261_), .A2(pi0609), .Z(new_n23311_));
  OAI21_X1   g20875(.A1(new_n13562_), .A2(new_n23061_), .B(pi0191), .ZN(new_n23312_));
  OAI21_X1   g20876(.A1(new_n18102_), .A2(pi0746), .B(new_n13566_), .ZN(new_n23313_));
  NAND2_X1   g20877(.A1(new_n23313_), .A2(new_n2627_), .ZN(new_n23314_));
  AOI21_X1   g20878(.A1(new_n23314_), .A2(new_n12704_), .B(new_n3265_), .ZN(new_n23315_));
  OAI21_X1   g20879(.A1(new_n5337_), .A2(new_n23312_), .B(new_n23315_), .ZN(new_n23316_));
  NOR2_X1    g20880(.A1(new_n14172_), .A2(new_n12704_), .ZN(new_n23317_));
  NOR2_X1    g20881(.A1(new_n14174_), .A2(pi0191), .ZN(new_n23318_));
  OAI21_X1   g20882(.A1(new_n23317_), .A2(new_n23318_), .B(pi0746), .ZN(new_n23319_));
  NAND2_X1   g20883(.A1(new_n18110_), .A2(new_n12704_), .ZN(new_n23320_));
  OAI21_X1   g20884(.A1(new_n12704_), .A2(new_n15835_), .B(new_n23320_), .ZN(new_n23321_));
  NAND2_X1   g20885(.A1(new_n23321_), .A2(new_n16996_), .ZN(new_n23322_));
  NAND3_X1   g20886(.A1(new_n23322_), .A2(new_n2627_), .A3(new_n23319_), .ZN(new_n23323_));
  NOR2_X1    g20887(.A1(new_n14182_), .A2(pi0191), .ZN(new_n23324_));
  NOR2_X1    g20888(.A1(new_n14184_), .A2(new_n12704_), .ZN(new_n23325_));
  OAI21_X1   g20889(.A1(new_n23324_), .A2(new_n23325_), .B(new_n16996_), .ZN(new_n23326_));
  NOR2_X1    g20890(.A1(new_n14187_), .A2(new_n12704_), .ZN(new_n23327_));
  NOR2_X1    g20891(.A1(new_n14189_), .A2(pi0191), .ZN(new_n23328_));
  OAI21_X1   g20892(.A1(new_n23327_), .A2(new_n23328_), .B(pi0746), .ZN(new_n23329_));
  NAND3_X1   g20893(.A1(new_n23329_), .A2(new_n23326_), .A3(pi0039), .ZN(new_n23330_));
  NAND3_X1   g20894(.A1(new_n23323_), .A2(new_n23330_), .A3(new_n3265_), .ZN(new_n23331_));
  NAND3_X1   g20895(.A1(new_n23331_), .A2(pi0729), .A3(new_n23316_), .ZN(new_n23332_));
  NAND2_X1   g20896(.A1(new_n23332_), .A2(new_n2609_), .ZN(new_n23333_));
  NOR2_X1    g20897(.A1(new_n23209_), .A2(pi0729), .ZN(new_n23334_));
  OAI21_X1   g20898(.A1(new_n23333_), .A2(new_n23334_), .B(new_n23246_), .ZN(new_n23335_));
  OR2_X2     g20899(.A1(new_n23210_), .A2(new_n13521_), .Z(new_n23336_));
  NAND2_X1   g20900(.A1(new_n23335_), .A2(new_n13521_), .ZN(new_n23337_));
  AOI21_X1   g20901(.A1(new_n23337_), .A2(new_n23336_), .B(pi1153), .ZN(new_n23338_));
  NOR3_X1    g20902(.A1(new_n23338_), .A2(pi0608), .A3(new_n23259_), .ZN(new_n23339_));
  NOR2_X1    g20903(.A1(new_n23210_), .A2(pi0625), .ZN(new_n23340_));
  AOI21_X1   g20904(.A1(new_n23335_), .A2(pi0625), .B(new_n23340_), .ZN(new_n23341_));
  NOR2_X1    g20905(.A1(new_n23341_), .A2(new_n12841_), .ZN(new_n23342_));
  NOR3_X1    g20906(.A1(new_n23342_), .A2(new_n13560_), .A3(new_n23256_), .ZN(new_n23343_));
  NOR3_X1    g20907(.A1(new_n23343_), .A2(new_n23339_), .A3(new_n12758_), .ZN(new_n23344_));
  AOI21_X1   g20908(.A1(new_n12758_), .A2(new_n23335_), .B(new_n23344_), .ZN(new_n23345_));
  OAI21_X1   g20909(.A1(new_n23345_), .A2(new_n12766_), .B(new_n23311_), .ZN(new_n23346_));
  AOI21_X1   g20910(.A1(new_n23346_), .A2(pi1155), .B(new_n23215_), .ZN(new_n23347_));
  NOR2_X1    g20911(.A1(new_n23345_), .A2(pi0609), .ZN(new_n23348_));
  NOR2_X1    g20912(.A1(new_n23261_), .A2(new_n12766_), .ZN(new_n23349_));
  OAI21_X1   g20913(.A1(new_n23348_), .A2(new_n23349_), .B(new_n12770_), .ZN(new_n23350_));
  NOR2_X1    g20914(.A1(new_n23217_), .A2(pi0660), .ZN(new_n23351_));
  AOI22_X1   g20915(.A1(new_n23347_), .A2(pi0660), .B1(new_n23350_), .B2(new_n23351_), .ZN(new_n23352_));
  AND2_X2    g20916(.A1(new_n23352_), .A2(pi0785), .Z(new_n23353_));
  NOR2_X1    g20917(.A1(new_n23345_), .A2(pi0785), .ZN(new_n23354_));
  NOR2_X1    g20918(.A1(new_n23353_), .A2(new_n23354_), .ZN(new_n23355_));
  NOR2_X1    g20919(.A1(new_n23355_), .A2(pi0781), .ZN(new_n23356_));
  NOR2_X1    g20920(.A1(new_n23263_), .A2(pi0618), .ZN(new_n23357_));
  INV_X1     g20921(.I(new_n23357_), .ZN(new_n23358_));
  OAI21_X1   g20922(.A1(new_n23353_), .A2(new_n23354_), .B(pi0618), .ZN(new_n23359_));
  AOI21_X1   g20923(.A1(new_n23359_), .A2(new_n23358_), .B(new_n12785_), .ZN(new_n23360_));
  NOR3_X1    g20924(.A1(new_n23360_), .A2(new_n12880_), .A3(new_n23223_), .ZN(new_n23361_));
  OAI21_X1   g20925(.A1(new_n23353_), .A2(new_n23354_), .B(new_n12781_), .ZN(new_n23362_));
  NAND3_X1   g20926(.A1(new_n23262_), .A2(pi0618), .A3(new_n23245_), .ZN(new_n23363_));
  AOI21_X1   g20927(.A1(new_n23362_), .A2(new_n23363_), .B(pi1154), .ZN(new_n23364_));
  NOR3_X1    g20928(.A1(new_n23364_), .A2(pi0627), .A3(new_n23226_), .ZN(new_n23365_));
  NOR3_X1    g20929(.A1(new_n23361_), .A2(new_n23365_), .A3(new_n12779_), .ZN(new_n23366_));
  OAI21_X1   g20930(.A1(new_n23366_), .A2(new_n23356_), .B(new_n12796_), .ZN(new_n23367_));
  NAND2_X1   g20931(.A1(new_n23367_), .A2(new_n12819_), .ZN(new_n23368_));
  NAND2_X1   g20932(.A1(new_n23265_), .A2(pi0619), .ZN(new_n23369_));
  OAI21_X1   g20933(.A1(new_n23366_), .A2(new_n23356_), .B(new_n12793_), .ZN(new_n23370_));
  AOI21_X1   g20934(.A1(new_n23370_), .A2(new_n23369_), .B(pi1159), .ZN(new_n23371_));
  NOR3_X1    g20935(.A1(new_n23371_), .A2(pi0648), .A3(new_n23234_), .ZN(new_n23372_));
  INV_X1     g20936(.I(new_n23231_), .ZN(new_n23373_));
  OAI21_X1   g20937(.A1(new_n23366_), .A2(new_n23356_), .B(pi0619), .ZN(new_n23374_));
  NAND2_X1   g20938(.A1(new_n23265_), .A2(new_n12793_), .ZN(new_n23375_));
  AOI21_X1   g20939(.A1(new_n23374_), .A2(new_n23375_), .B(new_n12791_), .ZN(new_n23376_));
  NOR3_X1    g20940(.A1(new_n23376_), .A2(new_n12895_), .A3(new_n23373_), .ZN(new_n23377_));
  NOR3_X1    g20941(.A1(new_n23372_), .A2(new_n23377_), .A3(new_n12796_), .ZN(new_n23378_));
  OAI21_X1   g20942(.A1(new_n23378_), .A2(new_n23368_), .B(new_n23310_), .ZN(new_n23379_));
  AOI21_X1   g20943(.A1(new_n23379_), .A2(new_n23303_), .B(new_n15341_), .ZN(new_n23380_));
  NOR3_X1    g20944(.A1(new_n23295_), .A2(new_n23300_), .A3(new_n23380_), .ZN(new_n23381_));
  OAI21_X1   g20945(.A1(new_n23381_), .A2(new_n23292_), .B(new_n6643_), .ZN(new_n23382_));
  AOI21_X1   g20946(.A1(po1038), .A2(new_n12704_), .B(pi0832), .ZN(new_n23383_));
  AOI21_X1   g20947(.A1(new_n23382_), .A2(new_n23383_), .B(new_n23194_), .ZN(po0348));
  NOR2_X1    g20948(.A1(new_n3042_), .A2(pi0192), .ZN(new_n23385_));
  NOR2_X1    g20949(.A1(new_n13340_), .A2(new_n17096_), .ZN(new_n23386_));
  NOR2_X1    g20950(.A1(new_n23386_), .A2(new_n23385_), .ZN(new_n23387_));
  NOR3_X1    g20951(.A1(new_n23387_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n23388_));
  INV_X1     g20952(.I(new_n23386_), .ZN(new_n23389_));
  NOR2_X1    g20953(.A1(new_n23389_), .A2(new_n13354_), .ZN(new_n23390_));
  NOR3_X1    g20954(.A1(new_n23390_), .A2(new_n12762_), .A3(new_n23387_), .ZN(new_n23391_));
  NOR2_X1    g20955(.A1(new_n23391_), .A2(new_n12770_), .ZN(new_n23392_));
  NOR3_X1    g20956(.A1(new_n23390_), .A2(pi1155), .A3(new_n23385_), .ZN(new_n23393_));
  NOR3_X1    g20957(.A1(new_n23392_), .A2(new_n12764_), .A3(new_n23393_), .ZN(new_n23394_));
  NOR2_X1    g20958(.A1(new_n23394_), .A2(new_n23388_), .ZN(new_n23395_));
  NOR2_X1    g20959(.A1(new_n23395_), .A2(pi0781), .ZN(new_n23396_));
  INV_X1     g20960(.I(new_n23395_), .ZN(new_n23397_));
  AOI21_X1   g20961(.A1(new_n23397_), .A2(new_n12783_), .B(pi1154), .ZN(new_n23398_));
  AOI21_X1   g20962(.A1(new_n23397_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n23399_));
  NOR3_X1    g20963(.A1(new_n23398_), .A2(new_n23399_), .A3(new_n12779_), .ZN(new_n23400_));
  NOR2_X1    g20964(.A1(new_n23400_), .A2(new_n23396_), .ZN(new_n23401_));
  NOR2_X1    g20965(.A1(new_n23401_), .A2(new_n17229_), .ZN(new_n23402_));
  NOR2_X1    g20966(.A1(new_n23402_), .A2(pi1159), .ZN(new_n23403_));
  OAI21_X1   g20967(.A1(new_n23401_), .A2(new_n17232_), .B(pi1159), .ZN(new_n23404_));
  NAND2_X1   g20968(.A1(new_n23404_), .A2(pi0789), .ZN(new_n23405_));
  OAI22_X1   g20969(.A1(new_n23405_), .A2(new_n23403_), .B1(pi0789), .B2(new_n23401_), .ZN(new_n23406_));
  INV_X1     g20970(.I(new_n23385_), .ZN(new_n23407_));
  NAND2_X1   g20971(.A1(new_n12818_), .A2(new_n23407_), .ZN(new_n23408_));
  OAI21_X1   g20972(.A1(new_n23406_), .A2(new_n12818_), .B(new_n23408_), .ZN(new_n23409_));
  AOI21_X1   g20973(.A1(new_n12826_), .A2(pi0691), .B(new_n23385_), .ZN(new_n23410_));
  INV_X1     g20974(.I(pi0691), .ZN(new_n23411_));
  NOR2_X1    g20975(.A1(new_n12834_), .A2(new_n23411_), .ZN(new_n23412_));
  INV_X1     g20976(.I(new_n23412_), .ZN(new_n23413_));
  NOR2_X1    g20977(.A1(new_n23385_), .A2(pi1153), .ZN(new_n23414_));
  NAND2_X1   g20978(.A1(new_n23413_), .A2(new_n23414_), .ZN(new_n23415_));
  NOR2_X1    g20979(.A1(new_n23412_), .A2(new_n23410_), .ZN(new_n23416_));
  NOR2_X1    g20980(.A1(new_n23416_), .A2(new_n12841_), .ZN(new_n23417_));
  INV_X1     g20981(.I(new_n23417_), .ZN(new_n23418_));
  NAND3_X1   g20982(.A1(new_n23418_), .A2(pi0778), .A3(new_n23415_), .ZN(new_n23419_));
  OAI21_X1   g20983(.A1(pi0778), .A2(new_n23410_), .B(new_n23419_), .ZN(new_n23420_));
  NAND2_X1   g20984(.A1(new_n23420_), .A2(new_n17187_), .ZN(new_n23421_));
  NOR2_X1    g20985(.A1(new_n23421_), .A2(new_n12889_), .ZN(new_n23422_));
  INV_X1     g20986(.I(new_n23422_), .ZN(new_n23423_));
  NOR2_X1    g20987(.A1(new_n23423_), .A2(new_n12912_), .ZN(new_n23424_));
  INV_X1     g20988(.I(new_n23424_), .ZN(new_n23425_));
  NOR2_X1    g20989(.A1(new_n23425_), .A2(new_n17884_), .ZN(new_n23426_));
  INV_X1     g20990(.I(new_n23426_), .ZN(new_n23427_));
  OAI22_X1   g20991(.A1(new_n23409_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n23427_), .ZN(new_n23428_));
  NAND2_X1   g20992(.A1(new_n23428_), .A2(new_n12919_), .ZN(new_n23429_));
  OAI22_X1   g20993(.A1(new_n23409_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n23427_), .ZN(new_n23430_));
  NAND2_X1   g20994(.A1(new_n23430_), .A2(pi0629), .ZN(new_n23431_));
  AOI21_X1   g20995(.A1(new_n23429_), .A2(new_n23431_), .B(new_n12937_), .ZN(new_n23432_));
  INV_X1     g20996(.I(new_n23393_), .ZN(new_n23433_));
  NOR2_X1    g20997(.A1(new_n23410_), .A2(new_n12754_), .ZN(new_n23434_));
  NOR3_X1    g20998(.A1(new_n23434_), .A2(new_n23385_), .A3(new_n23386_), .ZN(new_n23435_));
  NAND2_X1   g20999(.A1(new_n23435_), .A2(new_n12758_), .ZN(new_n23436_));
  NAND2_X1   g21000(.A1(new_n23434_), .A2(pi0625), .ZN(new_n23437_));
  NAND3_X1   g21001(.A1(new_n23437_), .A2(pi1153), .A3(new_n23387_), .ZN(new_n23438_));
  NAND3_X1   g21002(.A1(new_n23415_), .A2(pi0608), .A3(new_n23438_), .ZN(new_n23439_));
  INV_X1     g21003(.I(new_n23437_), .ZN(new_n23440_));
  OAI21_X1   g21004(.A1(new_n23440_), .A2(new_n23435_), .B(new_n23414_), .ZN(new_n23441_));
  NAND3_X1   g21005(.A1(new_n23418_), .A2(new_n13560_), .A3(new_n23441_), .ZN(new_n23442_));
  NAND3_X1   g21006(.A1(new_n23442_), .A2(pi0778), .A3(new_n23439_), .ZN(new_n23443_));
  AOI21_X1   g21007(.A1(new_n23443_), .A2(new_n23436_), .B(new_n12766_), .ZN(new_n23444_));
  NOR2_X1    g21008(.A1(new_n23420_), .A2(pi0609), .ZN(new_n23445_));
  OAI21_X1   g21009(.A1(new_n23445_), .A2(new_n23444_), .B(pi1155), .ZN(new_n23446_));
  NAND3_X1   g21010(.A1(new_n23446_), .A2(pi0660), .A3(new_n23433_), .ZN(new_n23447_));
  NAND2_X1   g21011(.A1(new_n23443_), .A2(new_n23436_), .ZN(new_n23448_));
  NOR2_X1    g21012(.A1(new_n23420_), .A2(new_n12766_), .ZN(new_n23449_));
  AOI21_X1   g21013(.A1(new_n23448_), .A2(new_n12766_), .B(new_n23449_), .ZN(new_n23450_));
  NOR2_X1    g21014(.A1(new_n23392_), .A2(pi0660), .ZN(new_n23451_));
  OAI21_X1   g21015(.A1(new_n23450_), .A2(pi1155), .B(new_n23451_), .ZN(new_n23452_));
  NAND3_X1   g21016(.A1(new_n23452_), .A2(new_n23447_), .A3(pi0785), .ZN(new_n23453_));
  NAND2_X1   g21017(.A1(new_n23448_), .A2(new_n12764_), .ZN(new_n23454_));
  NAND2_X1   g21018(.A1(new_n23453_), .A2(new_n23454_), .ZN(new_n23455_));
  NAND2_X1   g21019(.A1(new_n23455_), .A2(new_n12781_), .ZN(new_n23456_));
  NAND2_X1   g21020(.A1(new_n23421_), .A2(pi0618), .ZN(new_n23457_));
  AOI21_X1   g21021(.A1(new_n23456_), .A2(new_n23457_), .B(pi1154), .ZN(new_n23458_));
  NOR3_X1    g21022(.A1(new_n23458_), .A2(pi0627), .A3(new_n23399_), .ZN(new_n23459_));
  NAND2_X1   g21023(.A1(new_n23421_), .A2(new_n12781_), .ZN(new_n23460_));
  NAND2_X1   g21024(.A1(new_n23455_), .A2(pi0618), .ZN(new_n23461_));
  AOI21_X1   g21025(.A1(new_n23461_), .A2(new_n23460_), .B(new_n12785_), .ZN(new_n23462_));
  NOR3_X1    g21026(.A1(new_n23462_), .A2(new_n12880_), .A3(new_n23398_), .ZN(new_n23463_));
  OR3_X2     g21027(.A1(new_n23459_), .A2(new_n23463_), .A3(new_n12779_), .Z(new_n23464_));
  NAND2_X1   g21028(.A1(new_n23455_), .A2(new_n12779_), .ZN(new_n23465_));
  NAND2_X1   g21029(.A1(new_n23464_), .A2(new_n23465_), .ZN(new_n23466_));
  AOI21_X1   g21030(.A1(new_n23466_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n23467_));
  NAND2_X1   g21031(.A1(new_n23423_), .A2(new_n12793_), .ZN(new_n23468_));
  NAND2_X1   g21032(.A1(new_n23466_), .A2(pi0619), .ZN(new_n23469_));
  AOI21_X1   g21033(.A1(new_n23469_), .A2(new_n23468_), .B(new_n12791_), .ZN(new_n23470_));
  NOR3_X1    g21034(.A1(new_n23470_), .A2(new_n12895_), .A3(new_n23403_), .ZN(new_n23471_));
  AOI21_X1   g21035(.A1(new_n23464_), .A2(new_n23465_), .B(pi0619), .ZN(new_n23472_));
  NOR2_X1    g21036(.A1(new_n23422_), .A2(new_n12793_), .ZN(new_n23473_));
  OAI21_X1   g21037(.A1(new_n23472_), .A2(new_n23473_), .B(new_n12791_), .ZN(new_n23474_));
  NAND3_X1   g21038(.A1(new_n23474_), .A2(new_n12895_), .A3(new_n23404_), .ZN(new_n23475_));
  NAND2_X1   g21039(.A1(new_n23475_), .A2(pi0789), .ZN(new_n23476_));
  OAI21_X1   g21040(.A1(new_n23476_), .A2(new_n23471_), .B(new_n23467_), .ZN(new_n23477_));
  NAND2_X1   g21041(.A1(new_n23385_), .A2(pi0626), .ZN(new_n23478_));
  NAND2_X1   g21042(.A1(new_n23406_), .A2(new_n12747_), .ZN(new_n23479_));
  AOI21_X1   g21043(.A1(new_n23479_), .A2(new_n23478_), .B(new_n12816_), .ZN(new_n23480_));
  NOR2_X1    g21044(.A1(new_n23407_), .A2(pi0626), .ZN(new_n23481_));
  AOI21_X1   g21045(.A1(new_n23406_), .A2(pi0626), .B(new_n23481_), .ZN(new_n23482_));
  OAI22_X1   g21046(.A1(new_n23482_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n23425_), .ZN(new_n23483_));
  OAI21_X1   g21047(.A1(new_n23483_), .A2(new_n23480_), .B(pi0788), .ZN(new_n23484_));
  AOI21_X1   g21048(.A1(new_n23477_), .A2(new_n23484_), .B(new_n15340_), .ZN(new_n23485_));
  OR2_X2     g21049(.A1(new_n23485_), .A2(new_n23432_), .Z(new_n23486_));
  NAND2_X1   g21050(.A1(new_n23409_), .A2(new_n13384_), .ZN(new_n23487_));
  NAND2_X1   g21051(.A1(new_n12943_), .A2(new_n23407_), .ZN(new_n23488_));
  AOI21_X1   g21052(.A1(new_n23487_), .A2(new_n23488_), .B(new_n17212_), .ZN(new_n23489_));
  NOR2_X1    g21053(.A1(new_n23427_), .A2(new_n12953_), .ZN(new_n23490_));
  NOR2_X1    g21054(.A1(new_n23490_), .A2(pi0647), .ZN(new_n23491_));
  NOR2_X1    g21055(.A1(new_n23385_), .A2(new_n12741_), .ZN(new_n23492_));
  OAI21_X1   g21056(.A1(new_n23491_), .A2(new_n23492_), .B(new_n12965_), .ZN(new_n23493_));
  NOR2_X1    g21057(.A1(new_n23407_), .A2(pi0647), .ZN(new_n23494_));
  AOI21_X1   g21058(.A1(new_n23490_), .A2(pi0647), .B(new_n23494_), .ZN(new_n23495_));
  INV_X1     g21059(.I(new_n23495_), .ZN(new_n23496_));
  OAI22_X1   g21060(.A1(new_n23493_), .A2(new_n12981_), .B1(new_n23496_), .B2(new_n15576_), .ZN(new_n23497_));
  NOR2_X1    g21061(.A1(new_n23497_), .A2(new_n23489_), .ZN(new_n23498_));
  OAI22_X1   g21062(.A1(new_n23486_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n23498_), .ZN(new_n23499_));
  OAI21_X1   g21063(.A1(new_n12965_), .A2(new_n23496_), .B(new_n23493_), .ZN(new_n23500_));
  NOR2_X1    g21064(.A1(new_n23500_), .A2(new_n12972_), .ZN(new_n23501_));
  AOI21_X1   g21065(.A1(new_n12972_), .A2(new_n23490_), .B(new_n23501_), .ZN(new_n23502_));
  AND2_X2    g21066(.A1(new_n23502_), .A2(pi0644), .Z(new_n23503_));
  AOI21_X1   g21067(.A1(new_n23499_), .A2(new_n12975_), .B(new_n23503_), .ZN(new_n23504_));
  NAND2_X1   g21068(.A1(new_n23407_), .A2(pi0644), .ZN(new_n23505_));
  NOR2_X1    g21069(.A1(new_n17611_), .A2(new_n23385_), .ZN(new_n23506_));
  AOI21_X1   g21070(.A1(new_n23409_), .A2(new_n17611_), .B(new_n23506_), .ZN(new_n23507_));
  OAI21_X1   g21071(.A1(new_n23507_), .A2(pi0644), .B(new_n23505_), .ZN(new_n23508_));
  NAND2_X1   g21072(.A1(new_n23508_), .A2(pi0715), .ZN(new_n23509_));
  OAI21_X1   g21073(.A1(new_n23504_), .A2(pi0715), .B(new_n23509_), .ZN(new_n23510_));
  NAND2_X1   g21074(.A1(new_n23499_), .A2(pi0644), .ZN(new_n23511_));
  NAND2_X1   g21075(.A1(new_n23502_), .A2(new_n12975_), .ZN(new_n23512_));
  AOI21_X1   g21076(.A1(new_n23511_), .A2(new_n23512_), .B(new_n12740_), .ZN(new_n23513_));
  OAI21_X1   g21077(.A1(new_n23407_), .A2(pi0644), .B(new_n12740_), .ZN(new_n23514_));
  AND2_X2    g21078(.A1(new_n23507_), .A2(pi0644), .Z(new_n23515_));
  OAI21_X1   g21079(.A1(new_n23515_), .A2(new_n23514_), .B(pi1160), .ZN(new_n23516_));
  OAI22_X1   g21080(.A1(new_n23510_), .A2(pi1160), .B1(new_n23513_), .B2(new_n23516_), .ZN(new_n23517_));
  OAI21_X1   g21081(.A1(new_n23499_), .A2(pi0790), .B(pi0832), .ZN(new_n23518_));
  AOI21_X1   g21082(.A1(new_n23517_), .A2(pi0790), .B(new_n23518_), .ZN(new_n23519_));
  NOR2_X1    g21083(.A1(new_n13193_), .A2(pi0192), .ZN(new_n23520_));
  AOI21_X1   g21084(.A1(new_n23520_), .A2(pi0644), .B(new_n12740_), .ZN(new_n23521_));
  NOR2_X1    g21085(.A1(new_n23520_), .A2(new_n12985_), .ZN(new_n23522_));
  INV_X1     g21086(.I(new_n23520_), .ZN(new_n23523_));
  NAND2_X1   g21087(.A1(new_n23523_), .A2(new_n12943_), .ZN(new_n23524_));
  NOR2_X1    g21088(.A1(new_n2609_), .A2(new_n12412_), .ZN(new_n23525_));
  OAI22_X1   g21089(.A1(new_n17092_), .A2(pi0192), .B1(new_n17096_), .B2(new_n13208_), .ZN(new_n23526_));
  NAND3_X1   g21090(.A1(new_n17986_), .A2(new_n12412_), .A3(pi0764), .ZN(new_n23527_));
  NAND2_X1   g21091(.A1(new_n23527_), .A2(new_n23526_), .ZN(new_n23528_));
  OAI22_X1   g21092(.A1(new_n14065_), .A2(pi0764), .B1(new_n12412_), .B2(new_n14067_), .ZN(new_n23529_));
  AOI21_X1   g21093(.A1(pi0039), .A2(new_n23529_), .B(new_n23528_), .ZN(new_n23530_));
  NAND2_X1   g21094(.A1(new_n13397_), .A2(new_n12412_), .ZN(new_n23531_));
  NAND2_X1   g21095(.A1(new_n23531_), .A2(pi0038), .ZN(new_n23532_));
  NOR2_X1    g21096(.A1(new_n13342_), .A2(new_n17096_), .ZN(new_n23533_));
  OAI22_X1   g21097(.A1(new_n23530_), .A2(pi0038), .B1(new_n23532_), .B2(new_n23533_), .ZN(new_n23534_));
  AOI21_X1   g21098(.A1(new_n23534_), .A2(new_n2609_), .B(new_n23525_), .ZN(new_n23535_));
  NOR2_X1    g21099(.A1(new_n23535_), .A2(new_n12760_), .ZN(new_n23536_));
  NOR2_X1    g21100(.A1(new_n23520_), .A2(new_n12761_), .ZN(new_n23537_));
  NOR3_X1    g21101(.A1(new_n23536_), .A2(pi0785), .A3(new_n23537_), .ZN(new_n23538_));
  AOI22_X1   g21102(.A1(new_n23536_), .A2(new_n12766_), .B1(new_n13354_), .B2(new_n23523_), .ZN(new_n23539_));
  NOR2_X1    g21103(.A1(new_n23539_), .A2(pi1155), .ZN(new_n23540_));
  AOI22_X1   g21104(.A1(new_n23536_), .A2(pi0609), .B1(new_n13357_), .B2(new_n23523_), .ZN(new_n23541_));
  NOR2_X1    g21105(.A1(new_n23541_), .A2(new_n12770_), .ZN(new_n23542_));
  NOR3_X1    g21106(.A1(new_n23542_), .A2(new_n23540_), .A3(new_n12764_), .ZN(new_n23543_));
  NOR2_X1    g21107(.A1(new_n23543_), .A2(new_n23538_), .ZN(new_n23544_));
  NAND2_X1   g21108(.A1(new_n23544_), .A2(new_n12781_), .ZN(new_n23545_));
  NOR2_X1    g21109(.A1(new_n23520_), .A2(new_n12781_), .ZN(new_n23546_));
  INV_X1     g21110(.I(new_n23546_), .ZN(new_n23547_));
  AOI21_X1   g21111(.A1(new_n23545_), .A2(new_n23547_), .B(pi1154), .ZN(new_n23548_));
  NAND2_X1   g21112(.A1(new_n23544_), .A2(pi0618), .ZN(new_n23549_));
  NAND2_X1   g21113(.A1(new_n23523_), .A2(new_n12781_), .ZN(new_n23550_));
  AOI21_X1   g21114(.A1(new_n23549_), .A2(new_n23550_), .B(new_n12785_), .ZN(new_n23551_));
  OR2_X2     g21115(.A1(new_n23551_), .A2(new_n12779_), .Z(new_n23552_));
  OAI22_X1   g21116(.A1(new_n23552_), .A2(new_n23548_), .B1(pi0781), .B2(new_n23544_), .ZN(new_n23553_));
  NAND2_X1   g21117(.A1(new_n23523_), .A2(pi0619), .ZN(new_n23554_));
  OAI21_X1   g21118(.A1(new_n23553_), .A2(pi0619), .B(new_n23554_), .ZN(new_n23555_));
  NAND2_X1   g21119(.A1(new_n23555_), .A2(new_n12791_), .ZN(new_n23556_));
  NOR2_X1    g21120(.A1(new_n23553_), .A2(new_n12793_), .ZN(new_n23557_));
  AOI21_X1   g21121(.A1(new_n12793_), .A2(new_n23523_), .B(new_n23557_), .ZN(new_n23558_));
  NOR2_X1    g21122(.A1(new_n23558_), .A2(new_n12791_), .ZN(new_n23559_));
  NOR2_X1    g21123(.A1(new_n23559_), .A2(new_n12796_), .ZN(new_n23560_));
  AOI22_X1   g21124(.A1(new_n23560_), .A2(new_n23556_), .B1(new_n12796_), .B2(new_n23553_), .ZN(new_n23561_));
  NOR2_X1    g21125(.A1(new_n23520_), .A2(new_n17504_), .ZN(new_n23562_));
  AOI21_X1   g21126(.A1(new_n23561_), .A2(new_n17504_), .B(new_n23562_), .ZN(new_n23563_));
  OAI21_X1   g21127(.A1(new_n23563_), .A2(new_n12943_), .B(new_n23524_), .ZN(new_n23564_));
  AOI21_X1   g21128(.A1(new_n23564_), .A2(new_n12985_), .B(new_n23522_), .ZN(new_n23565_));
  NAND2_X1   g21129(.A1(new_n23565_), .A2(new_n12975_), .ZN(new_n23566_));
  AOI21_X1   g21130(.A1(new_n23566_), .A2(new_n23521_), .B(pi1160), .ZN(new_n23567_));
  NAND2_X1   g21131(.A1(new_n23523_), .A2(new_n12741_), .ZN(new_n23568_));
  NOR2_X1    g21132(.A1(new_n23520_), .A2(pi0628), .ZN(new_n23569_));
  NAND2_X1   g21133(.A1(new_n23520_), .A2(new_n12869_), .ZN(new_n23570_));
  INV_X1     g21134(.I(new_n23525_), .ZN(new_n23571_));
  NAND3_X1   g21135(.A1(new_n13395_), .A2(new_n12412_), .A3(new_n23411_), .ZN(new_n23572_));
  NOR2_X1    g21136(.A1(new_n18033_), .A2(new_n12412_), .ZN(new_n23573_));
  AOI21_X1   g21137(.A1(new_n12412_), .A2(new_n14118_), .B(new_n23573_), .ZN(new_n23574_));
  AOI21_X1   g21138(.A1(new_n13399_), .A2(new_n23531_), .B(new_n23411_), .ZN(new_n23575_));
  OAI21_X1   g21139(.A1(new_n23574_), .A2(pi0038), .B(new_n23575_), .ZN(new_n23576_));
  NAND3_X1   g21140(.A1(new_n23576_), .A2(new_n2609_), .A3(new_n23572_), .ZN(new_n23577_));
  NAND2_X1   g21141(.A1(new_n23577_), .A2(new_n23571_), .ZN(new_n23578_));
  NAND2_X1   g21142(.A1(new_n23523_), .A2(pi0625), .ZN(new_n23579_));
  NAND2_X1   g21143(.A1(new_n23578_), .A2(new_n13521_), .ZN(new_n23580_));
  AOI21_X1   g21144(.A1(new_n23580_), .A2(new_n23579_), .B(pi1153), .ZN(new_n23581_));
  NAND2_X1   g21145(.A1(new_n23523_), .A2(new_n13521_), .ZN(new_n23582_));
  NAND2_X1   g21146(.A1(new_n23578_), .A2(pi0625), .ZN(new_n23583_));
  AOI21_X1   g21147(.A1(new_n23583_), .A2(new_n23582_), .B(new_n12841_), .ZN(new_n23584_));
  OR2_X2     g21148(.A1(new_n23584_), .A2(new_n12758_), .Z(new_n23585_));
  OAI22_X1   g21149(.A1(new_n23585_), .A2(new_n23581_), .B1(pi0778), .B2(new_n23578_), .ZN(new_n23586_));
  NAND2_X1   g21150(.A1(new_n23586_), .A2(new_n12870_), .ZN(new_n23587_));
  NAND2_X1   g21151(.A1(new_n23587_), .A2(new_n23570_), .ZN(new_n23588_));
  NAND2_X1   g21152(.A1(new_n23523_), .A2(new_n12887_), .ZN(new_n23589_));
  OAI21_X1   g21153(.A1(new_n23588_), .A2(new_n12887_), .B(new_n23589_), .ZN(new_n23590_));
  NAND2_X1   g21154(.A1(new_n23520_), .A2(new_n12910_), .ZN(new_n23591_));
  OAI21_X1   g21155(.A1(new_n23590_), .A2(new_n12910_), .B(new_n23591_), .ZN(new_n23592_));
  NAND2_X1   g21156(.A1(new_n23523_), .A2(new_n12817_), .ZN(new_n23593_));
  OAI21_X1   g21157(.A1(new_n23592_), .A2(new_n12817_), .B(new_n23593_), .ZN(new_n23594_));
  AOI21_X1   g21158(.A1(new_n23594_), .A2(pi0628), .B(new_n23569_), .ZN(new_n23595_));
  NOR2_X1    g21159(.A1(new_n23595_), .A2(new_n12742_), .ZN(new_n23596_));
  NOR2_X1    g21160(.A1(new_n23520_), .A2(new_n12920_), .ZN(new_n23597_));
  AOI21_X1   g21161(.A1(new_n23594_), .A2(new_n12920_), .B(new_n23597_), .ZN(new_n23598_));
  NOR2_X1    g21162(.A1(new_n23598_), .A2(pi1156), .ZN(new_n23599_));
  OAI21_X1   g21163(.A1(new_n23596_), .A2(new_n23599_), .B(pi0792), .ZN(new_n23600_));
  NAND2_X1   g21164(.A1(new_n23594_), .A2(new_n12937_), .ZN(new_n23601_));
  NAND2_X1   g21165(.A1(new_n23600_), .A2(new_n23601_), .ZN(new_n23602_));
  NAND2_X1   g21166(.A1(new_n23602_), .A2(pi0647), .ZN(new_n23603_));
  AOI21_X1   g21167(.A1(new_n23603_), .A2(new_n23568_), .B(new_n12965_), .ZN(new_n23604_));
  NAND2_X1   g21168(.A1(new_n23523_), .A2(pi0647), .ZN(new_n23605_));
  NAND2_X1   g21169(.A1(new_n23602_), .A2(new_n12741_), .ZN(new_n23606_));
  AOI21_X1   g21170(.A1(new_n23606_), .A2(new_n23605_), .B(pi1157), .ZN(new_n23607_));
  OAI21_X1   g21171(.A1(new_n23604_), .A2(new_n23607_), .B(pi0787), .ZN(new_n23608_));
  NAND2_X1   g21172(.A1(new_n23602_), .A2(new_n12972_), .ZN(new_n23609_));
  NAND2_X1   g21173(.A1(new_n23608_), .A2(new_n23609_), .ZN(new_n23610_));
  OAI21_X1   g21174(.A1(new_n23610_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n23611_));
  AOI21_X1   g21175(.A1(new_n23520_), .A2(new_n12975_), .B(pi0715), .ZN(new_n23612_));
  NAND2_X1   g21176(.A1(new_n23565_), .A2(pi0644), .ZN(new_n23613_));
  AOI21_X1   g21177(.A1(new_n23613_), .A2(new_n23612_), .B(new_n12739_), .ZN(new_n23614_));
  OAI21_X1   g21178(.A1(new_n23610_), .A2(pi0644), .B(pi0715), .ZN(new_n23615_));
  AOI22_X1   g21179(.A1(new_n23567_), .A2(new_n23611_), .B1(new_n23614_), .B2(new_n23615_), .ZN(new_n23616_));
  NOR2_X1    g21180(.A1(new_n23616_), .A2(new_n13000_), .ZN(new_n23617_));
  OR2_X2     g21181(.A1(new_n23614_), .A2(new_n12975_), .Z(new_n23618_));
  OR2_X2     g21182(.A1(new_n23567_), .A2(pi0644), .Z(new_n23619_));
  AOI21_X1   g21183(.A1(new_n23618_), .A2(new_n23619_), .B(new_n13000_), .ZN(new_n23620_));
  NAND2_X1   g21184(.A1(new_n23603_), .A2(new_n23568_), .ZN(new_n23621_));
  NAND2_X1   g21185(.A1(new_n23606_), .A2(new_n23605_), .ZN(new_n23622_));
  AOI22_X1   g21186(.A1(new_n12980_), .A2(new_n23621_), .B1(new_n23622_), .B2(new_n12982_), .ZN(new_n23623_));
  NAND2_X1   g21187(.A1(new_n23564_), .A2(new_n15608_), .ZN(new_n23624_));
  AOI21_X1   g21188(.A1(new_n23624_), .A2(new_n23623_), .B(new_n12972_), .ZN(new_n23625_));
  OAI22_X1   g21189(.A1(new_n18087_), .A2(new_n23595_), .B1(new_n23598_), .B2(new_n18088_), .ZN(new_n23626_));
  NOR2_X1    g21190(.A1(new_n23563_), .A2(new_n15821_), .ZN(new_n23627_));
  OAI21_X1   g21191(.A1(new_n23627_), .A2(new_n23626_), .B(pi0792), .ZN(new_n23628_));
  NOR2_X1    g21192(.A1(new_n23561_), .A2(pi0626), .ZN(new_n23629_));
  AOI21_X1   g21193(.A1(pi0626), .A2(new_n23520_), .B(new_n23629_), .ZN(new_n23630_));
  NAND2_X1   g21194(.A1(new_n23520_), .A2(new_n12747_), .ZN(new_n23631_));
  OAI21_X1   g21195(.A1(new_n23561_), .A2(new_n12747_), .B(new_n23631_), .ZN(new_n23632_));
  AOI22_X1   g21196(.A1(new_n23632_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n23592_), .ZN(new_n23633_));
  OAI21_X1   g21197(.A1(new_n12816_), .A2(new_n23630_), .B(new_n23633_), .ZN(new_n23634_));
  AOI21_X1   g21198(.A1(new_n23634_), .A2(pi0788), .B(new_n15340_), .ZN(new_n23635_));
  OR2_X2     g21199(.A1(new_n23586_), .A2(pi0609), .Z(new_n23636_));
  OAI21_X1   g21200(.A1(new_n13562_), .A2(new_n23386_), .B(pi0192), .ZN(new_n23637_));
  OAI21_X1   g21201(.A1(new_n18102_), .A2(pi0764), .B(new_n13566_), .ZN(new_n23638_));
  NAND2_X1   g21202(.A1(new_n23638_), .A2(new_n2627_), .ZN(new_n23639_));
  AOI21_X1   g21203(.A1(new_n23639_), .A2(new_n12412_), .B(new_n3265_), .ZN(new_n23640_));
  OAI21_X1   g21204(.A1(new_n5337_), .A2(new_n23637_), .B(new_n23640_), .ZN(new_n23641_));
  NOR2_X1    g21205(.A1(new_n14172_), .A2(new_n12412_), .ZN(new_n23642_));
  NOR2_X1    g21206(.A1(new_n14174_), .A2(pi0192), .ZN(new_n23643_));
  OAI21_X1   g21207(.A1(new_n23642_), .A2(new_n23643_), .B(pi0764), .ZN(new_n23644_));
  NAND2_X1   g21208(.A1(new_n18110_), .A2(new_n12412_), .ZN(new_n23645_));
  OAI21_X1   g21209(.A1(new_n12412_), .A2(new_n15835_), .B(new_n23645_), .ZN(new_n23646_));
  NAND2_X1   g21210(.A1(new_n23646_), .A2(new_n17096_), .ZN(new_n23647_));
  NAND3_X1   g21211(.A1(new_n23647_), .A2(new_n2627_), .A3(new_n23644_), .ZN(new_n23648_));
  NOR2_X1    g21212(.A1(new_n14182_), .A2(pi0192), .ZN(new_n23649_));
  NOR2_X1    g21213(.A1(new_n14184_), .A2(new_n12412_), .ZN(new_n23650_));
  OAI21_X1   g21214(.A1(new_n23649_), .A2(new_n23650_), .B(new_n17096_), .ZN(new_n23651_));
  NOR2_X1    g21215(.A1(new_n14187_), .A2(new_n12412_), .ZN(new_n23652_));
  NOR2_X1    g21216(.A1(new_n14189_), .A2(pi0192), .ZN(new_n23653_));
  OAI21_X1   g21217(.A1(new_n23652_), .A2(new_n23653_), .B(pi0764), .ZN(new_n23654_));
  NAND3_X1   g21218(.A1(new_n23654_), .A2(new_n23651_), .A3(pi0039), .ZN(new_n23655_));
  NAND3_X1   g21219(.A1(new_n23648_), .A2(new_n23655_), .A3(new_n3265_), .ZN(new_n23656_));
  NAND3_X1   g21220(.A1(new_n23656_), .A2(pi0691), .A3(new_n23641_), .ZN(new_n23657_));
  NAND2_X1   g21221(.A1(new_n23657_), .A2(new_n2609_), .ZN(new_n23658_));
  NOR2_X1    g21222(.A1(new_n23534_), .A2(pi0691), .ZN(new_n23659_));
  OAI21_X1   g21223(.A1(new_n23658_), .A2(new_n23659_), .B(new_n23571_), .ZN(new_n23660_));
  OR2_X2     g21224(.A1(new_n23535_), .A2(new_n13521_), .Z(new_n23661_));
  NAND2_X1   g21225(.A1(new_n23660_), .A2(new_n13521_), .ZN(new_n23662_));
  AOI21_X1   g21226(.A1(new_n23662_), .A2(new_n23661_), .B(pi1153), .ZN(new_n23663_));
  NOR3_X1    g21227(.A1(new_n23663_), .A2(pi0608), .A3(new_n23584_), .ZN(new_n23664_));
  NOR2_X1    g21228(.A1(new_n23535_), .A2(pi0625), .ZN(new_n23665_));
  AOI21_X1   g21229(.A1(new_n23660_), .A2(pi0625), .B(new_n23665_), .ZN(new_n23666_));
  NOR2_X1    g21230(.A1(new_n23666_), .A2(new_n12841_), .ZN(new_n23667_));
  NOR3_X1    g21231(.A1(new_n23667_), .A2(new_n13560_), .A3(new_n23581_), .ZN(new_n23668_));
  NOR3_X1    g21232(.A1(new_n23668_), .A2(new_n23664_), .A3(new_n12758_), .ZN(new_n23669_));
  AOI21_X1   g21233(.A1(new_n12758_), .A2(new_n23660_), .B(new_n23669_), .ZN(new_n23670_));
  OAI21_X1   g21234(.A1(new_n23670_), .A2(new_n12766_), .B(new_n23636_), .ZN(new_n23671_));
  AOI21_X1   g21235(.A1(new_n23671_), .A2(pi1155), .B(new_n23540_), .ZN(new_n23672_));
  NOR2_X1    g21236(.A1(new_n23670_), .A2(pi0609), .ZN(new_n23673_));
  NOR2_X1    g21237(.A1(new_n23586_), .A2(new_n12766_), .ZN(new_n23674_));
  OAI21_X1   g21238(.A1(new_n23673_), .A2(new_n23674_), .B(new_n12770_), .ZN(new_n23675_));
  NOR2_X1    g21239(.A1(new_n23542_), .A2(pi0660), .ZN(new_n23676_));
  AOI22_X1   g21240(.A1(new_n23672_), .A2(pi0660), .B1(new_n23675_), .B2(new_n23676_), .ZN(new_n23677_));
  AND2_X2    g21241(.A1(new_n23677_), .A2(pi0785), .Z(new_n23678_));
  NOR2_X1    g21242(.A1(new_n23670_), .A2(pi0785), .ZN(new_n23679_));
  NOR2_X1    g21243(.A1(new_n23678_), .A2(new_n23679_), .ZN(new_n23680_));
  NOR2_X1    g21244(.A1(new_n23680_), .A2(pi0781), .ZN(new_n23681_));
  NOR2_X1    g21245(.A1(new_n23588_), .A2(pi0618), .ZN(new_n23682_));
  INV_X1     g21246(.I(new_n23682_), .ZN(new_n23683_));
  OAI21_X1   g21247(.A1(new_n23678_), .A2(new_n23679_), .B(pi0618), .ZN(new_n23684_));
  AOI21_X1   g21248(.A1(new_n23684_), .A2(new_n23683_), .B(new_n12785_), .ZN(new_n23685_));
  NOR3_X1    g21249(.A1(new_n23685_), .A2(new_n12880_), .A3(new_n23548_), .ZN(new_n23686_));
  OAI21_X1   g21250(.A1(new_n23678_), .A2(new_n23679_), .B(new_n12781_), .ZN(new_n23687_));
  NAND3_X1   g21251(.A1(new_n23587_), .A2(pi0618), .A3(new_n23570_), .ZN(new_n23688_));
  AOI21_X1   g21252(.A1(new_n23687_), .A2(new_n23688_), .B(pi1154), .ZN(new_n23689_));
  NOR3_X1    g21253(.A1(new_n23689_), .A2(pi0627), .A3(new_n23551_), .ZN(new_n23690_));
  NOR3_X1    g21254(.A1(new_n23686_), .A2(new_n23690_), .A3(new_n12779_), .ZN(new_n23691_));
  OAI21_X1   g21255(.A1(new_n23691_), .A2(new_n23681_), .B(new_n12796_), .ZN(new_n23692_));
  NAND2_X1   g21256(.A1(new_n23692_), .A2(new_n12819_), .ZN(new_n23693_));
  NAND2_X1   g21257(.A1(new_n23590_), .A2(pi0619), .ZN(new_n23694_));
  OAI21_X1   g21258(.A1(new_n23691_), .A2(new_n23681_), .B(new_n12793_), .ZN(new_n23695_));
  AOI21_X1   g21259(.A1(new_n23695_), .A2(new_n23694_), .B(pi1159), .ZN(new_n23696_));
  NOR3_X1    g21260(.A1(new_n23696_), .A2(pi0648), .A3(new_n23559_), .ZN(new_n23697_));
  INV_X1     g21261(.I(new_n23556_), .ZN(new_n23698_));
  OAI21_X1   g21262(.A1(new_n23691_), .A2(new_n23681_), .B(pi0619), .ZN(new_n23699_));
  NAND2_X1   g21263(.A1(new_n23590_), .A2(new_n12793_), .ZN(new_n23700_));
  AOI21_X1   g21264(.A1(new_n23699_), .A2(new_n23700_), .B(new_n12791_), .ZN(new_n23701_));
  NOR3_X1    g21265(.A1(new_n23701_), .A2(new_n12895_), .A3(new_n23698_), .ZN(new_n23702_));
  NOR3_X1    g21266(.A1(new_n23697_), .A2(new_n23702_), .A3(new_n12796_), .ZN(new_n23703_));
  OAI21_X1   g21267(.A1(new_n23703_), .A2(new_n23693_), .B(new_n23635_), .ZN(new_n23704_));
  AOI21_X1   g21268(.A1(new_n23704_), .A2(new_n23628_), .B(new_n15341_), .ZN(new_n23705_));
  NOR3_X1    g21269(.A1(new_n23620_), .A2(new_n23625_), .A3(new_n23705_), .ZN(new_n23706_));
  OAI21_X1   g21270(.A1(new_n23706_), .A2(new_n23617_), .B(new_n6643_), .ZN(new_n23707_));
  AOI21_X1   g21271(.A1(po1038), .A2(new_n12412_), .B(pi0832), .ZN(new_n23708_));
  AOI21_X1   g21272(.A1(new_n23707_), .A2(new_n23708_), .B(new_n23519_), .ZN(po0349));
  NOR2_X1    g21273(.A1(new_n13340_), .A2(new_n17135_), .ZN(new_n23710_));
  NOR2_X1    g21274(.A1(new_n3042_), .A2(pi0193), .ZN(new_n23711_));
  NOR2_X1    g21275(.A1(new_n23710_), .A2(new_n23711_), .ZN(new_n23712_));
  NOR3_X1    g21276(.A1(new_n23712_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n23713_));
  INV_X1     g21277(.I(new_n23710_), .ZN(new_n23714_));
  NOR2_X1    g21278(.A1(new_n23714_), .A2(new_n13354_), .ZN(new_n23715_));
  NOR3_X1    g21279(.A1(new_n23715_), .A2(new_n12762_), .A3(new_n23712_), .ZN(new_n23716_));
  NOR2_X1    g21280(.A1(new_n23716_), .A2(new_n12770_), .ZN(new_n23717_));
  NOR3_X1    g21281(.A1(new_n23715_), .A2(pi1155), .A3(new_n23711_), .ZN(new_n23718_));
  NOR3_X1    g21282(.A1(new_n23717_), .A2(new_n12764_), .A3(new_n23718_), .ZN(new_n23719_));
  NOR2_X1    g21283(.A1(new_n23719_), .A2(new_n23713_), .ZN(new_n23720_));
  INV_X1     g21284(.I(new_n23720_), .ZN(new_n23721_));
  AOI21_X1   g21285(.A1(new_n23721_), .A2(new_n12783_), .B(pi1154), .ZN(new_n23722_));
  AOI21_X1   g21286(.A1(new_n23721_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n23723_));
  NOR3_X1    g21287(.A1(new_n23722_), .A2(new_n23723_), .A3(new_n12779_), .ZN(new_n23724_));
  AOI21_X1   g21288(.A1(new_n12779_), .A2(new_n23721_), .B(new_n23724_), .ZN(new_n23725_));
  OAI21_X1   g21289(.A1(new_n23725_), .A2(new_n17229_), .B(new_n12791_), .ZN(new_n23726_));
  OAI21_X1   g21290(.A1(new_n23725_), .A2(new_n17232_), .B(pi1159), .ZN(new_n23727_));
  NAND3_X1   g21291(.A1(new_n23726_), .A2(new_n23727_), .A3(pi0789), .ZN(new_n23728_));
  OAI21_X1   g21292(.A1(pi0789), .A2(new_n23725_), .B(new_n23728_), .ZN(new_n23729_));
  INV_X1     g21293(.I(new_n23711_), .ZN(new_n23730_));
  NAND2_X1   g21294(.A1(new_n12818_), .A2(new_n23730_), .ZN(new_n23731_));
  OAI21_X1   g21295(.A1(new_n23729_), .A2(new_n12818_), .B(new_n23731_), .ZN(new_n23732_));
  AOI21_X1   g21296(.A1(new_n12826_), .A2(pi0690), .B(new_n23711_), .ZN(new_n23733_));
  NOR2_X1    g21297(.A1(new_n12834_), .A2(new_n17137_), .ZN(new_n23734_));
  INV_X1     g21298(.I(new_n23734_), .ZN(new_n23735_));
  NOR2_X1    g21299(.A1(new_n23711_), .A2(pi1153), .ZN(new_n23736_));
  NAND2_X1   g21300(.A1(new_n23735_), .A2(new_n23736_), .ZN(new_n23737_));
  NOR2_X1    g21301(.A1(new_n23734_), .A2(new_n23733_), .ZN(new_n23738_));
  NOR2_X1    g21302(.A1(new_n23738_), .A2(new_n12841_), .ZN(new_n23739_));
  INV_X1     g21303(.I(new_n23739_), .ZN(new_n23740_));
  NAND3_X1   g21304(.A1(new_n23740_), .A2(pi0778), .A3(new_n23737_), .ZN(new_n23741_));
  OAI21_X1   g21305(.A1(pi0778), .A2(new_n23733_), .B(new_n23741_), .ZN(new_n23742_));
  NAND2_X1   g21306(.A1(new_n23742_), .A2(new_n17187_), .ZN(new_n23743_));
  NOR2_X1    g21307(.A1(new_n23743_), .A2(new_n12889_), .ZN(new_n23744_));
  NAND2_X1   g21308(.A1(new_n23744_), .A2(new_n18203_), .ZN(new_n23745_));
  NOR2_X1    g21309(.A1(new_n23745_), .A2(new_n17884_), .ZN(new_n23746_));
  INV_X1     g21310(.I(new_n23746_), .ZN(new_n23747_));
  OAI22_X1   g21311(.A1(new_n23732_), .A2(new_n15694_), .B1(new_n15696_), .B2(new_n23747_), .ZN(new_n23748_));
  AND2_X2    g21312(.A1(new_n23748_), .A2(new_n12919_), .Z(new_n23749_));
  OAI22_X1   g21313(.A1(new_n23732_), .A2(new_n15699_), .B1(new_n15701_), .B2(new_n23747_), .ZN(new_n23750_));
  AOI21_X1   g21314(.A1(pi0629), .A2(new_n23750_), .B(new_n23749_), .ZN(new_n23751_));
  INV_X1     g21315(.I(new_n23718_), .ZN(new_n23752_));
  NOR2_X1    g21316(.A1(new_n23733_), .A2(new_n12754_), .ZN(new_n23753_));
  NOR3_X1    g21317(.A1(new_n23753_), .A2(new_n23710_), .A3(new_n23711_), .ZN(new_n23754_));
  NAND2_X1   g21318(.A1(new_n23754_), .A2(new_n12758_), .ZN(new_n23755_));
  NAND2_X1   g21319(.A1(new_n23753_), .A2(pi0625), .ZN(new_n23756_));
  NAND3_X1   g21320(.A1(new_n23756_), .A2(pi1153), .A3(new_n23712_), .ZN(new_n23757_));
  NAND3_X1   g21321(.A1(new_n23737_), .A2(pi0608), .A3(new_n23757_), .ZN(new_n23758_));
  INV_X1     g21322(.I(new_n23756_), .ZN(new_n23759_));
  OAI21_X1   g21323(.A1(new_n23759_), .A2(new_n23754_), .B(new_n23736_), .ZN(new_n23760_));
  NAND3_X1   g21324(.A1(new_n23740_), .A2(new_n13560_), .A3(new_n23760_), .ZN(new_n23761_));
  NAND3_X1   g21325(.A1(new_n23761_), .A2(pi0778), .A3(new_n23758_), .ZN(new_n23762_));
  AOI21_X1   g21326(.A1(new_n23762_), .A2(new_n23755_), .B(new_n12766_), .ZN(new_n23763_));
  NOR2_X1    g21327(.A1(new_n23742_), .A2(pi0609), .ZN(new_n23764_));
  OAI21_X1   g21328(.A1(new_n23764_), .A2(new_n23763_), .B(pi1155), .ZN(new_n23765_));
  NAND3_X1   g21329(.A1(new_n23765_), .A2(pi0660), .A3(new_n23752_), .ZN(new_n23766_));
  NAND2_X1   g21330(.A1(new_n23762_), .A2(new_n23755_), .ZN(new_n23767_));
  NOR2_X1    g21331(.A1(new_n23742_), .A2(new_n12766_), .ZN(new_n23768_));
  AOI21_X1   g21332(.A1(new_n23767_), .A2(new_n12766_), .B(new_n23768_), .ZN(new_n23769_));
  NOR2_X1    g21333(.A1(new_n23717_), .A2(pi0660), .ZN(new_n23770_));
  OAI21_X1   g21334(.A1(new_n23769_), .A2(pi1155), .B(new_n23770_), .ZN(new_n23771_));
  NAND3_X1   g21335(.A1(new_n23771_), .A2(new_n23766_), .A3(pi0785), .ZN(new_n23772_));
  NAND2_X1   g21336(.A1(new_n23767_), .A2(new_n12764_), .ZN(new_n23773_));
  NAND2_X1   g21337(.A1(new_n23772_), .A2(new_n23773_), .ZN(new_n23774_));
  NAND2_X1   g21338(.A1(new_n23774_), .A2(new_n12781_), .ZN(new_n23775_));
  NAND2_X1   g21339(.A1(new_n23743_), .A2(pi0618), .ZN(new_n23776_));
  AOI21_X1   g21340(.A1(new_n23775_), .A2(new_n23776_), .B(pi1154), .ZN(new_n23777_));
  NOR3_X1    g21341(.A1(new_n23777_), .A2(pi0627), .A3(new_n23723_), .ZN(new_n23778_));
  NAND2_X1   g21342(.A1(new_n23743_), .A2(new_n12781_), .ZN(new_n23779_));
  NAND2_X1   g21343(.A1(new_n23774_), .A2(pi0618), .ZN(new_n23780_));
  AOI21_X1   g21344(.A1(new_n23780_), .A2(new_n23779_), .B(new_n12785_), .ZN(new_n23781_));
  NOR3_X1    g21345(.A1(new_n23781_), .A2(new_n12880_), .A3(new_n23722_), .ZN(new_n23782_));
  OR3_X2     g21346(.A1(new_n23778_), .A2(new_n23782_), .A3(new_n12779_), .Z(new_n23783_));
  NAND2_X1   g21347(.A1(new_n23774_), .A2(new_n12779_), .ZN(new_n23784_));
  NAND2_X1   g21348(.A1(new_n23783_), .A2(new_n23784_), .ZN(new_n23785_));
  AOI21_X1   g21349(.A1(new_n23785_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n23786_));
  NOR2_X1    g21350(.A1(new_n23744_), .A2(pi0619), .ZN(new_n23787_));
  AOI21_X1   g21351(.A1(new_n23783_), .A2(new_n23784_), .B(new_n12793_), .ZN(new_n23788_));
  OAI21_X1   g21352(.A1(new_n23788_), .A2(new_n23787_), .B(pi1159), .ZN(new_n23789_));
  NAND3_X1   g21353(.A1(new_n23789_), .A2(pi0648), .A3(new_n23726_), .ZN(new_n23790_));
  NAND2_X1   g21354(.A1(new_n23785_), .A2(new_n12793_), .ZN(new_n23791_));
  OAI21_X1   g21355(.A1(new_n12793_), .A2(new_n23744_), .B(new_n23791_), .ZN(new_n23792_));
  NAND2_X1   g21356(.A1(new_n23792_), .A2(new_n12791_), .ZN(new_n23793_));
  NAND3_X1   g21357(.A1(new_n23793_), .A2(new_n12895_), .A3(new_n23727_), .ZN(new_n23794_));
  NAND3_X1   g21358(.A1(new_n23794_), .A2(pi0789), .A3(new_n23790_), .ZN(new_n23795_));
  NOR2_X1    g21359(.A1(new_n23730_), .A2(new_n12747_), .ZN(new_n23796_));
  AND2_X2    g21360(.A1(new_n23729_), .A2(new_n12747_), .Z(new_n23797_));
  OAI21_X1   g21361(.A1(new_n23797_), .A2(new_n23796_), .B(new_n12815_), .ZN(new_n23798_));
  INV_X1     g21362(.I(new_n23745_), .ZN(new_n23799_));
  NAND2_X1   g21363(.A1(new_n23729_), .A2(pi0626), .ZN(new_n23800_));
  OAI21_X1   g21364(.A1(pi0626), .A2(new_n23730_), .B(new_n23800_), .ZN(new_n23801_));
  AOI22_X1   g21365(.A1(new_n23801_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n23799_), .ZN(new_n23802_));
  NAND2_X1   g21366(.A1(new_n23802_), .A2(new_n23798_), .ZN(new_n23803_));
  AOI22_X1   g21367(.A1(new_n23795_), .A2(new_n23786_), .B1(pi0788), .B2(new_n23803_), .ZN(new_n23804_));
  OAI22_X1   g21368(.A1(new_n23804_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n23751_), .ZN(new_n23805_));
  NAND2_X1   g21369(.A1(new_n23732_), .A2(new_n13384_), .ZN(new_n23806_));
  NAND2_X1   g21370(.A1(new_n12943_), .A2(new_n23730_), .ZN(new_n23807_));
  NAND2_X1   g21371(.A1(new_n23806_), .A2(new_n23807_), .ZN(new_n23808_));
  NOR2_X1    g21372(.A1(new_n23747_), .A2(new_n12953_), .ZN(new_n23809_));
  NOR2_X1    g21373(.A1(new_n23809_), .A2(pi0647), .ZN(new_n23810_));
  NOR2_X1    g21374(.A1(new_n23711_), .A2(new_n12741_), .ZN(new_n23811_));
  OAI21_X1   g21375(.A1(new_n23810_), .A2(new_n23811_), .B(new_n12965_), .ZN(new_n23812_));
  NAND2_X1   g21376(.A1(new_n23809_), .A2(pi0647), .ZN(new_n23813_));
  OAI21_X1   g21377(.A1(pi0647), .A2(new_n23730_), .B(new_n23813_), .ZN(new_n23814_));
  OAI22_X1   g21378(.A1(new_n23814_), .A2(new_n15576_), .B1(new_n23812_), .B2(new_n12981_), .ZN(new_n23815_));
  AOI21_X1   g21379(.A1(new_n23808_), .A2(new_n15608_), .B(new_n23815_), .ZN(new_n23816_));
  OAI22_X1   g21380(.A1(new_n23805_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n23816_), .ZN(new_n23817_));
  NAND2_X1   g21381(.A1(new_n23817_), .A2(new_n13000_), .ZN(new_n23818_));
  AND2_X2    g21382(.A1(new_n23817_), .A2(new_n12975_), .Z(new_n23819_));
  OAI21_X1   g21383(.A1(new_n23814_), .A2(new_n12965_), .B(new_n23812_), .ZN(new_n23820_));
  NAND2_X1   g21384(.A1(new_n23809_), .A2(new_n12972_), .ZN(new_n23821_));
  OAI21_X1   g21385(.A1(new_n23820_), .A2(new_n12972_), .B(new_n23821_), .ZN(new_n23822_));
  NOR2_X1    g21386(.A1(new_n23822_), .A2(new_n12975_), .ZN(new_n23823_));
  OAI21_X1   g21387(.A1(new_n23819_), .A2(new_n23823_), .B(new_n12740_), .ZN(new_n23824_));
  NAND2_X1   g21388(.A1(new_n23730_), .A2(pi0644), .ZN(new_n23825_));
  NOR2_X1    g21389(.A1(new_n17611_), .A2(new_n23711_), .ZN(new_n23826_));
  AOI21_X1   g21390(.A1(new_n23732_), .A2(new_n17611_), .B(new_n23826_), .ZN(new_n23827_));
  OAI21_X1   g21391(.A1(new_n23827_), .A2(pi0644), .B(new_n23825_), .ZN(new_n23828_));
  NAND2_X1   g21392(.A1(new_n23828_), .A2(pi0715), .ZN(new_n23829_));
  NAND3_X1   g21393(.A1(new_n23824_), .A2(new_n12739_), .A3(new_n23829_), .ZN(new_n23830_));
  NOR2_X1    g21394(.A1(new_n23822_), .A2(pi0644), .ZN(new_n23831_));
  AOI21_X1   g21395(.A1(new_n23817_), .A2(pi0644), .B(new_n23831_), .ZN(new_n23832_));
  NAND2_X1   g21396(.A1(new_n23730_), .A2(new_n12975_), .ZN(new_n23833_));
  OAI21_X1   g21397(.A1(new_n23827_), .A2(new_n12975_), .B(new_n23833_), .ZN(new_n23834_));
  AOI21_X1   g21398(.A1(new_n23834_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n23835_));
  OAI21_X1   g21399(.A1(new_n23832_), .A2(new_n12740_), .B(new_n23835_), .ZN(new_n23836_));
  NAND3_X1   g21400(.A1(new_n23830_), .A2(pi0790), .A3(new_n23836_), .ZN(new_n23837_));
  NAND2_X1   g21401(.A1(new_n23837_), .A2(new_n23818_), .ZN(new_n23838_));
  AOI21_X1   g21402(.A1(po1038), .A2(new_n7858_), .B(pi0832), .ZN(new_n23839_));
  NAND2_X1   g21403(.A1(new_n13192_), .A2(new_n7858_), .ZN(new_n23840_));
  INV_X1     g21404(.I(new_n23840_), .ZN(new_n23841_));
  AOI21_X1   g21405(.A1(new_n23841_), .A2(pi0644), .B(new_n12740_), .ZN(new_n23842_));
  NAND2_X1   g21406(.A1(new_n23840_), .A2(new_n12984_), .ZN(new_n23843_));
  NOR2_X1    g21407(.A1(new_n23841_), .A2(new_n13384_), .ZN(new_n23844_));
  NOR2_X1    g21408(.A1(new_n2609_), .A2(new_n7858_), .ZN(new_n23845_));
  NOR2_X1    g21409(.A1(new_n13342_), .A2(new_n17135_), .ZN(new_n23846_));
  NOR2_X1    g21410(.A1(new_n13344_), .A2(pi0193), .ZN(new_n23847_));
  NOR3_X1    g21411(.A1(new_n23846_), .A2(new_n3265_), .A3(new_n23847_), .ZN(new_n23848_));
  NAND2_X1   g21412(.A1(new_n13334_), .A2(new_n7858_), .ZN(new_n23849_));
  NAND2_X1   g21413(.A1(new_n13245_), .A2(pi0193), .ZN(new_n23850_));
  AOI21_X1   g21414(.A1(new_n23849_), .A2(new_n23850_), .B(new_n17135_), .ZN(new_n23851_));
  NOR3_X1    g21415(.A1(new_n15787_), .A2(pi0193), .A3(pi0739), .ZN(new_n23852_));
  NOR2_X1    g21416(.A1(new_n23851_), .A2(new_n23852_), .ZN(new_n23853_));
  AOI21_X1   g21417(.A1(new_n23853_), .A2(new_n3265_), .B(new_n23848_), .ZN(new_n23854_));
  NOR2_X1    g21418(.A1(new_n23854_), .A2(new_n2610_), .ZN(new_n23855_));
  NOR2_X1    g21419(.A1(new_n23855_), .A2(new_n23845_), .ZN(new_n23856_));
  NOR2_X1    g21420(.A1(new_n23856_), .A2(new_n12760_), .ZN(new_n23857_));
  INV_X1     g21421(.I(new_n23857_), .ZN(new_n23858_));
  OAI21_X1   g21422(.A1(new_n12761_), .A2(new_n23841_), .B(new_n23858_), .ZN(new_n23859_));
  OAI22_X1   g21423(.A1(new_n23858_), .A2(pi0609), .B1(new_n13353_), .B2(new_n23841_), .ZN(new_n23860_));
  NAND2_X1   g21424(.A1(new_n23860_), .A2(new_n12770_), .ZN(new_n23861_));
  INV_X1     g21425(.I(new_n23861_), .ZN(new_n23862_));
  AOI22_X1   g21426(.A1(new_n23857_), .A2(pi0609), .B1(new_n13357_), .B2(new_n23840_), .ZN(new_n23863_));
  OAI21_X1   g21427(.A1(new_n23863_), .A2(new_n12770_), .B(pi0785), .ZN(new_n23864_));
  OAI22_X1   g21428(.A1(new_n23862_), .A2(new_n23864_), .B1(pi0785), .B2(new_n23859_), .ZN(new_n23865_));
  NAND2_X1   g21429(.A1(new_n23865_), .A2(new_n12779_), .ZN(new_n23866_));
  NAND2_X1   g21430(.A1(new_n23840_), .A2(pi0618), .ZN(new_n23867_));
  OAI21_X1   g21431(.A1(new_n23865_), .A2(pi0618), .B(new_n23867_), .ZN(new_n23868_));
  NAND2_X1   g21432(.A1(new_n23868_), .A2(new_n12785_), .ZN(new_n23869_));
  NAND2_X1   g21433(.A1(new_n23840_), .A2(new_n12781_), .ZN(new_n23870_));
  OAI21_X1   g21434(.A1(new_n23865_), .A2(new_n12781_), .B(new_n23870_), .ZN(new_n23871_));
  NAND2_X1   g21435(.A1(new_n23871_), .A2(pi1154), .ZN(new_n23872_));
  NAND3_X1   g21436(.A1(new_n23869_), .A2(new_n23872_), .A3(pi0781), .ZN(new_n23873_));
  NAND2_X1   g21437(.A1(new_n23873_), .A2(new_n23866_), .ZN(new_n23874_));
  NAND2_X1   g21438(.A1(new_n23874_), .A2(new_n12796_), .ZN(new_n23875_));
  NAND2_X1   g21439(.A1(new_n23840_), .A2(pi0619), .ZN(new_n23876_));
  OAI21_X1   g21440(.A1(new_n23874_), .A2(pi0619), .B(new_n23876_), .ZN(new_n23877_));
  NAND2_X1   g21441(.A1(new_n23877_), .A2(new_n12791_), .ZN(new_n23878_));
  NAND2_X1   g21442(.A1(new_n23840_), .A2(new_n12793_), .ZN(new_n23879_));
  OAI21_X1   g21443(.A1(new_n23874_), .A2(new_n12793_), .B(new_n23879_), .ZN(new_n23880_));
  NAND2_X1   g21444(.A1(new_n23880_), .A2(pi1159), .ZN(new_n23881_));
  NAND3_X1   g21445(.A1(new_n23878_), .A2(new_n23881_), .A3(pi0789), .ZN(new_n23882_));
  NAND2_X1   g21446(.A1(new_n23882_), .A2(new_n23875_), .ZN(new_n23883_));
  NAND2_X1   g21447(.A1(new_n23840_), .A2(new_n12818_), .ZN(new_n23884_));
  OAI21_X1   g21448(.A1(new_n23883_), .A2(new_n12818_), .B(new_n23884_), .ZN(new_n23885_));
  AOI21_X1   g21449(.A1(new_n23885_), .A2(new_n13384_), .B(new_n23844_), .ZN(new_n23886_));
  OAI21_X1   g21450(.A1(new_n23886_), .A2(new_n12984_), .B(new_n23843_), .ZN(new_n23887_));
  OAI21_X1   g21451(.A1(new_n23887_), .A2(pi0644), .B(new_n23842_), .ZN(new_n23888_));
  AND2_X2    g21452(.A1(new_n23888_), .A2(new_n12739_), .Z(new_n23889_));
  OAI21_X1   g21453(.A1(new_n14125_), .A2(new_n23847_), .B(pi0690), .ZN(new_n23890_));
  OAI21_X1   g21454(.A1(new_n14122_), .A2(new_n7858_), .B(new_n3265_), .ZN(new_n23891_));
  NAND2_X1   g21455(.A1(new_n23891_), .A2(new_n2609_), .ZN(new_n23892_));
  NAND2_X1   g21456(.A1(new_n15744_), .A2(new_n7858_), .ZN(new_n23893_));
  AOI21_X1   g21457(.A1(new_n23893_), .A2(new_n23892_), .B(new_n23890_), .ZN(new_n23894_));
  NAND2_X1   g21458(.A1(new_n2609_), .A2(pi0690), .ZN(new_n23895_));
  AOI21_X1   g21459(.A1(new_n23841_), .A2(new_n23895_), .B(new_n23894_), .ZN(new_n23896_));
  NAND2_X1   g21460(.A1(new_n23896_), .A2(new_n13521_), .ZN(new_n23897_));
  NAND2_X1   g21461(.A1(new_n23840_), .A2(pi0625), .ZN(new_n23898_));
  AOI21_X1   g21462(.A1(new_n23897_), .A2(new_n23898_), .B(pi1153), .ZN(new_n23899_));
  NAND2_X1   g21463(.A1(new_n23840_), .A2(new_n13521_), .ZN(new_n23900_));
  NAND2_X1   g21464(.A1(new_n23896_), .A2(pi0625), .ZN(new_n23901_));
  AOI21_X1   g21465(.A1(new_n23901_), .A2(new_n23900_), .B(new_n12841_), .ZN(new_n23902_));
  NOR3_X1    g21466(.A1(new_n23899_), .A2(new_n23902_), .A3(new_n12758_), .ZN(new_n23903_));
  NOR2_X1    g21467(.A1(new_n23896_), .A2(pi0778), .ZN(new_n23904_));
  NOR2_X1    g21468(.A1(new_n23903_), .A2(new_n23904_), .ZN(new_n23905_));
  NOR2_X1    g21469(.A1(new_n23905_), .A2(new_n12869_), .ZN(new_n23906_));
  AOI21_X1   g21470(.A1(new_n12869_), .A2(new_n23841_), .B(new_n23906_), .ZN(new_n23907_));
  NAND2_X1   g21471(.A1(new_n23907_), .A2(new_n12888_), .ZN(new_n23908_));
  OAI21_X1   g21472(.A1(new_n12888_), .A2(new_n23841_), .B(new_n23908_), .ZN(new_n23909_));
  INV_X1     g21473(.I(new_n23909_), .ZN(new_n23910_));
  NOR2_X1    g21474(.A1(new_n23840_), .A2(new_n12911_), .ZN(new_n23911_));
  AOI21_X1   g21475(.A1(new_n23910_), .A2(new_n12911_), .B(new_n23911_), .ZN(new_n23912_));
  NAND2_X1   g21476(.A1(new_n23912_), .A2(new_n13392_), .ZN(new_n23913_));
  OAI21_X1   g21477(.A1(new_n13392_), .A2(new_n23841_), .B(new_n23913_), .ZN(new_n23914_));
  NAND2_X1   g21478(.A1(new_n23914_), .A2(new_n12920_), .ZN(new_n23915_));
  NAND2_X1   g21479(.A1(new_n23840_), .A2(pi0628), .ZN(new_n23916_));
  AOI21_X1   g21480(.A1(new_n23915_), .A2(new_n23916_), .B(pi1156), .ZN(new_n23917_));
  NAND2_X1   g21481(.A1(new_n23840_), .A2(new_n12920_), .ZN(new_n23918_));
  NAND2_X1   g21482(.A1(new_n23914_), .A2(pi0628), .ZN(new_n23919_));
  AOI21_X1   g21483(.A1(new_n23919_), .A2(new_n23918_), .B(new_n12742_), .ZN(new_n23920_));
  OR2_X2     g21484(.A1(new_n23920_), .A2(new_n12937_), .Z(new_n23921_));
  OAI22_X1   g21485(.A1(new_n23921_), .A2(new_n23917_), .B1(pi0792), .B2(new_n23914_), .ZN(new_n23922_));
  NAND2_X1   g21486(.A1(new_n23922_), .A2(new_n12741_), .ZN(new_n23923_));
  OAI21_X1   g21487(.A1(new_n12741_), .A2(new_n23840_), .B(new_n23923_), .ZN(new_n23924_));
  NOR2_X1    g21488(.A1(new_n23924_), .A2(pi1157), .ZN(new_n23925_));
  NAND2_X1   g21489(.A1(new_n23922_), .A2(pi0647), .ZN(new_n23926_));
  OAI21_X1   g21490(.A1(pi0647), .A2(new_n23840_), .B(new_n23926_), .ZN(new_n23927_));
  NOR2_X1    g21491(.A1(new_n23927_), .A2(new_n12965_), .ZN(new_n23928_));
  OAI21_X1   g21492(.A1(new_n23925_), .A2(new_n23928_), .B(pi0787), .ZN(new_n23929_));
  OAI21_X1   g21493(.A1(pi0787), .A2(new_n23922_), .B(new_n23929_), .ZN(new_n23930_));
  OAI21_X1   g21494(.A1(new_n23930_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n23931_));
  AOI21_X1   g21495(.A1(new_n23841_), .A2(new_n12975_), .B(pi0715), .ZN(new_n23932_));
  OAI21_X1   g21496(.A1(new_n23887_), .A2(new_n12975_), .B(new_n23932_), .ZN(new_n23933_));
  AND2_X2    g21497(.A1(new_n23933_), .A2(pi1160), .Z(new_n23934_));
  OAI21_X1   g21498(.A1(new_n23930_), .A2(pi0644), .B(pi0715), .ZN(new_n23935_));
  AOI22_X1   g21499(.A1(new_n23889_), .A2(new_n23931_), .B1(new_n23935_), .B2(new_n23934_), .ZN(new_n23936_));
  NOR2_X1    g21500(.A1(new_n23936_), .A2(new_n13000_), .ZN(new_n23937_));
  NAND2_X1   g21501(.A1(new_n23841_), .A2(pi0626), .ZN(new_n23938_));
  NAND2_X1   g21502(.A1(new_n23883_), .A2(new_n12747_), .ZN(new_n23939_));
  AOI21_X1   g21503(.A1(new_n23939_), .A2(new_n23938_), .B(new_n12816_), .ZN(new_n23940_));
  NOR2_X1    g21504(.A1(new_n23840_), .A2(pi0626), .ZN(new_n23941_));
  AOI21_X1   g21505(.A1(new_n23883_), .A2(pi0626), .B(new_n23941_), .ZN(new_n23942_));
  OAI22_X1   g21506(.A1(new_n23942_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n23912_), .ZN(new_n23943_));
  OAI21_X1   g21507(.A1(new_n23943_), .A2(new_n23940_), .B(pi0788), .ZN(new_n23944_));
  NAND2_X1   g21508(.A1(new_n23944_), .A2(new_n15824_), .ZN(new_n23945_));
  NAND2_X1   g21509(.A1(new_n23905_), .A2(new_n12766_), .ZN(new_n23946_));
  OAI21_X1   g21510(.A1(new_n13562_), .A2(new_n23710_), .B(pi0193), .ZN(new_n23947_));
  OAI21_X1   g21511(.A1(new_n18102_), .A2(pi0739), .B(new_n13566_), .ZN(new_n23948_));
  NAND2_X1   g21512(.A1(new_n23948_), .A2(new_n2627_), .ZN(new_n23949_));
  AOI21_X1   g21513(.A1(new_n23949_), .A2(new_n7858_), .B(new_n3265_), .ZN(new_n23950_));
  OAI21_X1   g21514(.A1(new_n5337_), .A2(new_n23947_), .B(new_n23950_), .ZN(new_n23951_));
  NAND2_X1   g21515(.A1(new_n15835_), .A2(pi0193), .ZN(new_n23952_));
  NAND2_X1   g21516(.A1(new_n14177_), .A2(new_n7858_), .ZN(new_n23953_));
  AOI21_X1   g21517(.A1(new_n23953_), .A2(new_n23952_), .B(pi0739), .ZN(new_n23954_));
  NAND2_X1   g21518(.A1(new_n14172_), .A2(pi0193), .ZN(new_n23955_));
  NAND2_X1   g21519(.A1(new_n14174_), .A2(new_n7858_), .ZN(new_n23956_));
  AOI21_X1   g21520(.A1(new_n23955_), .A2(new_n23956_), .B(new_n17135_), .ZN(new_n23957_));
  OAI21_X1   g21521(.A1(new_n23954_), .A2(new_n23957_), .B(new_n2627_), .ZN(new_n23958_));
  NOR2_X1    g21522(.A1(new_n14182_), .A2(pi0193), .ZN(new_n23959_));
  NOR2_X1    g21523(.A1(new_n14184_), .A2(new_n7858_), .ZN(new_n23960_));
  OAI21_X1   g21524(.A1(new_n23959_), .A2(new_n23960_), .B(new_n17135_), .ZN(new_n23961_));
  NOR2_X1    g21525(.A1(new_n14187_), .A2(new_n7858_), .ZN(new_n23962_));
  NOR2_X1    g21526(.A1(new_n14189_), .A2(pi0193), .ZN(new_n23963_));
  OAI21_X1   g21527(.A1(new_n23962_), .A2(new_n23963_), .B(pi0739), .ZN(new_n23964_));
  NAND3_X1   g21528(.A1(new_n23964_), .A2(new_n23961_), .A3(pi0039), .ZN(new_n23965_));
  NAND3_X1   g21529(.A1(new_n23965_), .A2(new_n3265_), .A3(new_n23958_), .ZN(new_n23966_));
  NAND3_X1   g21530(.A1(new_n23966_), .A2(pi0690), .A3(new_n23951_), .ZN(new_n23967_));
  NAND2_X1   g21531(.A1(new_n23854_), .A2(new_n17137_), .ZN(new_n23968_));
  NAND3_X1   g21532(.A1(new_n23967_), .A2(new_n2609_), .A3(new_n23968_), .ZN(new_n23969_));
  OAI21_X1   g21533(.A1(new_n7858_), .A2(new_n2609_), .B(new_n23969_), .ZN(new_n23970_));
  INV_X1     g21534(.I(new_n23902_), .ZN(new_n23971_));
  NOR2_X1    g21535(.A1(new_n23856_), .A2(new_n13521_), .ZN(new_n23972_));
  AOI21_X1   g21536(.A1(new_n23970_), .A2(new_n13521_), .B(new_n23972_), .ZN(new_n23973_));
  OAI21_X1   g21537(.A1(new_n23973_), .A2(pi1153), .B(new_n23971_), .ZN(new_n23974_));
  NOR2_X1    g21538(.A1(new_n23856_), .A2(pi0625), .ZN(new_n23975_));
  AOI21_X1   g21539(.A1(new_n23970_), .A2(pi0625), .B(new_n23975_), .ZN(new_n23976_));
  OAI21_X1   g21540(.A1(new_n23976_), .A2(new_n12841_), .B(pi0608), .ZN(new_n23977_));
  OAI22_X1   g21541(.A1(pi0608), .A2(new_n23974_), .B1(new_n23977_), .B2(new_n23899_), .ZN(new_n23978_));
  NOR2_X1    g21542(.A1(new_n23978_), .A2(new_n12758_), .ZN(new_n23979_));
  AOI21_X1   g21543(.A1(new_n12758_), .A2(new_n23970_), .B(new_n23979_), .ZN(new_n23980_));
  OAI21_X1   g21544(.A1(new_n23980_), .A2(new_n12766_), .B(new_n23946_), .ZN(new_n23981_));
  AOI21_X1   g21545(.A1(new_n23981_), .A2(pi1155), .B(new_n23862_), .ZN(new_n23982_));
  NOR2_X1    g21546(.A1(new_n23980_), .A2(pi0609), .ZN(new_n23983_));
  NOR3_X1    g21547(.A1(new_n23903_), .A2(new_n12766_), .A3(new_n23904_), .ZN(new_n23984_));
  OAI21_X1   g21548(.A1(new_n23983_), .A2(new_n23984_), .B(new_n12770_), .ZN(new_n23985_));
  NOR2_X1    g21549(.A1(new_n23863_), .A2(new_n12770_), .ZN(new_n23986_));
  NOR2_X1    g21550(.A1(new_n23986_), .A2(pi0660), .ZN(new_n23987_));
  AOI22_X1   g21551(.A1(new_n23982_), .A2(pi0660), .B1(new_n23985_), .B2(new_n23987_), .ZN(new_n23988_));
  NOR2_X1    g21552(.A1(new_n23980_), .A2(pi0785), .ZN(new_n23989_));
  AOI21_X1   g21553(.A1(new_n23988_), .A2(pi0785), .B(new_n23989_), .ZN(new_n23990_));
  NOR2_X1    g21554(.A1(new_n23990_), .A2(pi0781), .ZN(new_n23991_));
  AND2_X2    g21555(.A1(new_n23907_), .A2(new_n12781_), .Z(new_n23992_));
  NOR2_X1    g21556(.A1(new_n23990_), .A2(new_n12781_), .ZN(new_n23993_));
  OAI21_X1   g21557(.A1(new_n23993_), .A2(new_n23992_), .B(pi1154), .ZN(new_n23994_));
  NAND3_X1   g21558(.A1(new_n23994_), .A2(pi0627), .A3(new_n23869_), .ZN(new_n23995_));
  INV_X1     g21559(.I(new_n23872_), .ZN(new_n23996_));
  NAND2_X1   g21560(.A1(new_n23907_), .A2(pi0618), .ZN(new_n23997_));
  OAI21_X1   g21561(.A1(new_n23990_), .A2(pi0618), .B(new_n23997_), .ZN(new_n23998_));
  AOI21_X1   g21562(.A1(new_n23998_), .A2(new_n12785_), .B(new_n23996_), .ZN(new_n23999_));
  AOI21_X1   g21563(.A1(new_n23999_), .A2(new_n12880_), .B(new_n12779_), .ZN(new_n24000_));
  AOI21_X1   g21564(.A1(new_n24000_), .A2(new_n23995_), .B(new_n23991_), .ZN(new_n24001_));
  OAI21_X1   g21565(.A1(new_n24001_), .A2(pi0789), .B(new_n12819_), .ZN(new_n24002_));
  NOR2_X1    g21566(.A1(new_n23910_), .A2(new_n12793_), .ZN(new_n24003_));
  NOR2_X1    g21567(.A1(new_n24001_), .A2(pi0619), .ZN(new_n24004_));
  OAI21_X1   g21568(.A1(new_n24004_), .A2(new_n24003_), .B(new_n12791_), .ZN(new_n24005_));
  NAND3_X1   g21569(.A1(new_n24005_), .A2(new_n12895_), .A3(new_n23881_), .ZN(new_n24006_));
  NAND2_X1   g21570(.A1(new_n23909_), .A2(new_n12793_), .ZN(new_n24007_));
  OAI21_X1   g21571(.A1(new_n24001_), .A2(new_n12793_), .B(new_n24007_), .ZN(new_n24008_));
  AOI21_X1   g21572(.A1(new_n24008_), .A2(pi1159), .B(new_n12895_), .ZN(new_n24009_));
  AOI21_X1   g21573(.A1(new_n24009_), .A2(new_n23878_), .B(new_n12796_), .ZN(new_n24010_));
  AOI21_X1   g21574(.A1(new_n24010_), .A2(new_n24006_), .B(new_n24002_), .ZN(new_n24011_));
  NOR2_X1    g21575(.A1(new_n23920_), .A2(pi0629), .ZN(new_n24012_));
  NOR2_X1    g21576(.A1(new_n23917_), .A2(new_n12919_), .ZN(new_n24013_));
  NOR2_X1    g21577(.A1(new_n24012_), .A2(new_n24013_), .ZN(new_n24014_));
  AOI21_X1   g21578(.A1(new_n23885_), .A2(new_n19160_), .B(new_n24014_), .ZN(new_n24015_));
  OAI22_X1   g21579(.A1(new_n24011_), .A2(new_n23945_), .B1(new_n12937_), .B2(new_n24015_), .ZN(new_n24016_));
  NOR2_X1    g21580(.A1(new_n23934_), .A2(new_n12975_), .ZN(new_n24017_));
  NOR2_X1    g21581(.A1(new_n23889_), .A2(pi0644), .ZN(new_n24018_));
  NOR2_X1    g21582(.A1(new_n24017_), .A2(new_n24018_), .ZN(new_n24019_));
  OAI22_X1   g21583(.A1(new_n15576_), .A2(new_n23927_), .B1(new_n23924_), .B2(new_n15730_), .ZN(new_n24020_));
  NOR2_X1    g21584(.A1(new_n23886_), .A2(new_n17212_), .ZN(new_n24021_));
  NOR2_X1    g21585(.A1(new_n24020_), .A2(new_n24021_), .ZN(new_n24022_));
  OAI22_X1   g21586(.A1(new_n24019_), .A2(new_n13000_), .B1(new_n24022_), .B2(new_n12972_), .ZN(new_n24023_));
  AOI21_X1   g21587(.A1(new_n15693_), .A2(new_n24016_), .B(new_n24023_), .ZN(new_n24024_));
  OAI21_X1   g21588(.A1(new_n23937_), .A2(new_n24024_), .B(new_n6643_), .ZN(new_n24025_));
  AOI22_X1   g21589(.A1(new_n24025_), .A2(new_n23839_), .B1(pi0832), .B2(new_n23838_), .ZN(po0350));
  NOR2_X1    g21590(.A1(new_n3042_), .A2(pi0194), .ZN(new_n24027_));
  INV_X1     g21591(.I(new_n24027_), .ZN(new_n24028_));
  AOI21_X1   g21592(.A1(new_n12756_), .A2(pi0748), .B(new_n24027_), .ZN(new_n24029_));
  NOR3_X1    g21593(.A1(new_n24029_), .A2(pi0785), .A3(new_n12762_), .ZN(new_n24030_));
  NOR2_X1    g21594(.A1(new_n24029_), .A2(new_n12762_), .ZN(new_n24031_));
  AOI21_X1   g21595(.A1(new_n24031_), .A2(new_n12768_), .B(pi1155), .ZN(new_n24032_));
  INV_X1     g21596(.I(new_n24029_), .ZN(new_n24033_));
  AOI21_X1   g21597(.A1(new_n24033_), .A2(new_n12774_), .B(new_n12770_), .ZN(new_n24034_));
  NOR3_X1    g21598(.A1(new_n24032_), .A2(new_n24034_), .A3(new_n12764_), .ZN(new_n24035_));
  NOR2_X1    g21599(.A1(new_n24035_), .A2(new_n24030_), .ZN(new_n24036_));
  NOR2_X1    g21600(.A1(new_n24036_), .A2(pi0781), .ZN(new_n24037_));
  INV_X1     g21601(.I(new_n24036_), .ZN(new_n24038_));
  AOI21_X1   g21602(.A1(new_n24038_), .A2(new_n12783_), .B(pi1154), .ZN(new_n24039_));
  AOI21_X1   g21603(.A1(new_n24038_), .A2(new_n12787_), .B(new_n12785_), .ZN(new_n24040_));
  NOR3_X1    g21604(.A1(new_n24039_), .A2(new_n24040_), .A3(new_n12779_), .ZN(new_n24041_));
  NOR2_X1    g21605(.A1(new_n24041_), .A2(new_n24037_), .ZN(new_n24042_));
  NOR3_X1    g21606(.A1(new_n24041_), .A2(pi0619), .A3(new_n24037_), .ZN(new_n24043_));
  NOR2_X1    g21607(.A1(new_n24027_), .A2(new_n12793_), .ZN(new_n24044_));
  OAI21_X1   g21608(.A1(new_n24043_), .A2(new_n24044_), .B(new_n12791_), .ZN(new_n24045_));
  NAND2_X1   g21609(.A1(new_n24042_), .A2(pi0619), .ZN(new_n24046_));
  NAND2_X1   g21610(.A1(new_n24028_), .A2(new_n12793_), .ZN(new_n24047_));
  AOI21_X1   g21611(.A1(new_n24046_), .A2(new_n24047_), .B(new_n12791_), .ZN(new_n24048_));
  INV_X1     g21612(.I(new_n24048_), .ZN(new_n24049_));
  NAND3_X1   g21613(.A1(new_n24049_), .A2(pi0789), .A3(new_n24045_), .ZN(new_n24050_));
  OAI21_X1   g21614(.A1(pi0789), .A2(new_n24042_), .B(new_n24050_), .ZN(new_n24051_));
  NOR2_X1    g21615(.A1(new_n24051_), .A2(new_n12818_), .ZN(new_n24052_));
  AOI21_X1   g21616(.A1(new_n12818_), .A2(new_n24028_), .B(new_n24052_), .ZN(new_n24053_));
  AOI21_X1   g21617(.A1(new_n12826_), .A2(pi0730), .B(new_n24027_), .ZN(new_n24054_));
  NOR2_X1    g21618(.A1(new_n24054_), .A2(pi0778), .ZN(new_n24055_));
  INV_X1     g21619(.I(pi0730), .ZN(new_n24056_));
  NOR2_X1    g21620(.A1(new_n12834_), .A2(new_n24056_), .ZN(new_n24057_));
  INV_X1     g21621(.I(new_n24057_), .ZN(new_n24058_));
  NOR2_X1    g21622(.A1(new_n24027_), .A2(pi1153), .ZN(new_n24059_));
  NAND2_X1   g21623(.A1(new_n24058_), .A2(new_n24059_), .ZN(new_n24060_));
  INV_X1     g21624(.I(new_n24060_), .ZN(new_n24061_));
  NOR2_X1    g21625(.A1(new_n24057_), .A2(new_n24054_), .ZN(new_n24062_));
  NOR2_X1    g21626(.A1(new_n24062_), .A2(new_n12841_), .ZN(new_n24063_));
  NOR2_X1    g21627(.A1(new_n24061_), .A2(new_n24063_), .ZN(new_n24064_));
  AOI21_X1   g21628(.A1(new_n24064_), .A2(pi0778), .B(new_n24055_), .ZN(new_n24065_));
  NOR2_X1    g21629(.A1(new_n24065_), .A2(new_n12871_), .ZN(new_n24066_));
  INV_X1     g21630(.I(new_n24066_), .ZN(new_n24067_));
  NOR2_X1    g21631(.A1(new_n24067_), .A2(new_n12889_), .ZN(new_n24068_));
  NAND2_X1   g21632(.A1(new_n24068_), .A2(new_n18203_), .ZN(new_n24069_));
  NOR2_X1    g21633(.A1(new_n24069_), .A2(new_n17884_), .ZN(new_n24070_));
  AOI22_X1   g21634(.A1(new_n24053_), .A2(new_n12949_), .B1(new_n15695_), .B2(new_n24070_), .ZN(new_n24071_));
  NOR2_X1    g21635(.A1(new_n24071_), .A2(pi0629), .ZN(new_n24072_));
  AOI22_X1   g21636(.A1(new_n24053_), .A2(new_n12948_), .B1(new_n15700_), .B2(new_n24070_), .ZN(new_n24073_));
  NOR2_X1    g21637(.A1(new_n24073_), .A2(new_n12919_), .ZN(new_n24074_));
  NOR2_X1    g21638(.A1(new_n24072_), .A2(new_n24074_), .ZN(new_n24075_));
  NOR2_X1    g21639(.A1(new_n24054_), .A2(new_n12754_), .ZN(new_n24076_));
  NOR2_X1    g21640(.A1(new_n24076_), .A2(new_n24033_), .ZN(new_n24077_));
  NAND2_X1   g21641(.A1(new_n24077_), .A2(new_n12758_), .ZN(new_n24078_));
  NAND2_X1   g21642(.A1(new_n24076_), .A2(pi0625), .ZN(new_n24079_));
  NAND3_X1   g21643(.A1(new_n24079_), .A2(pi1153), .A3(new_n24029_), .ZN(new_n24080_));
  AND3_X2    g21644(.A1(new_n24060_), .A2(pi0608), .A3(new_n24080_), .Z(new_n24081_));
  NOR2_X1    g21645(.A1(new_n24063_), .A2(pi0608), .ZN(new_n24082_));
  INV_X1     g21646(.I(new_n24079_), .ZN(new_n24083_));
  OAI21_X1   g21647(.A1(new_n24083_), .A2(new_n24077_), .B(new_n24059_), .ZN(new_n24084_));
  NAND2_X1   g21648(.A1(new_n24082_), .A2(new_n24084_), .ZN(new_n24085_));
  NAND2_X1   g21649(.A1(new_n24085_), .A2(pi0778), .ZN(new_n24086_));
  OAI21_X1   g21650(.A1(new_n24086_), .A2(new_n24081_), .B(new_n24078_), .ZN(new_n24087_));
  INV_X1     g21651(.I(new_n24087_), .ZN(new_n24088_));
  NAND2_X1   g21652(.A1(new_n24065_), .A2(new_n12766_), .ZN(new_n24089_));
  OAI21_X1   g21653(.A1(new_n24088_), .A2(new_n12766_), .B(new_n24089_), .ZN(new_n24090_));
  AOI21_X1   g21654(.A1(new_n24090_), .A2(pi1155), .B(new_n24032_), .ZN(new_n24091_));
  NAND2_X1   g21655(.A1(new_n24087_), .A2(new_n12766_), .ZN(new_n24092_));
  NAND2_X1   g21656(.A1(new_n24065_), .A2(pi0609), .ZN(new_n24093_));
  AOI21_X1   g21657(.A1(new_n24092_), .A2(new_n24093_), .B(pi1155), .ZN(new_n24094_));
  NOR3_X1    g21658(.A1(new_n24094_), .A2(pi0660), .A3(new_n24034_), .ZN(new_n24095_));
  AOI21_X1   g21659(.A1(pi0660), .A2(new_n24091_), .B(new_n24095_), .ZN(new_n24096_));
  NAND2_X1   g21660(.A1(new_n24096_), .A2(pi0785), .ZN(new_n24097_));
  OAI21_X1   g21661(.A1(pi0785), .A2(new_n24088_), .B(new_n24097_), .ZN(new_n24098_));
  INV_X1     g21662(.I(new_n24098_), .ZN(new_n24099_));
  NAND2_X1   g21663(.A1(new_n24067_), .A2(pi0618), .ZN(new_n24100_));
  OAI21_X1   g21664(.A1(new_n24099_), .A2(pi0618), .B(new_n24100_), .ZN(new_n24101_));
  AOI21_X1   g21665(.A1(new_n24101_), .A2(new_n12785_), .B(new_n24040_), .ZN(new_n24102_));
  NOR2_X1    g21666(.A1(new_n24066_), .A2(pi0618), .ZN(new_n24103_));
  NOR2_X1    g21667(.A1(new_n24099_), .A2(new_n12781_), .ZN(new_n24104_));
  OAI21_X1   g21668(.A1(new_n24104_), .A2(new_n24103_), .B(pi1154), .ZN(new_n24105_));
  NOR2_X1    g21669(.A1(new_n24039_), .A2(new_n12880_), .ZN(new_n24106_));
  AOI22_X1   g21670(.A1(new_n24102_), .A2(new_n12880_), .B1(new_n24105_), .B2(new_n24106_), .ZN(new_n24107_));
  NAND2_X1   g21671(.A1(new_n24107_), .A2(pi0781), .ZN(new_n24108_));
  NAND2_X1   g21672(.A1(new_n24098_), .A2(new_n12779_), .ZN(new_n24109_));
  NAND2_X1   g21673(.A1(new_n24108_), .A2(new_n24109_), .ZN(new_n24110_));
  AOI21_X1   g21674(.A1(new_n24110_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n24111_));
  NOR2_X1    g21675(.A1(new_n24068_), .A2(pi0619), .ZN(new_n24112_));
  INV_X1     g21676(.I(new_n24110_), .ZN(new_n24113_));
  NOR2_X1    g21677(.A1(new_n24113_), .A2(new_n12793_), .ZN(new_n24114_));
  OAI21_X1   g21678(.A1(new_n24114_), .A2(new_n24112_), .B(pi1159), .ZN(new_n24115_));
  NAND3_X1   g21679(.A1(new_n24115_), .A2(pi0648), .A3(new_n24045_), .ZN(new_n24116_));
  NOR2_X1    g21680(.A1(new_n24113_), .A2(pi0619), .ZN(new_n24117_));
  NOR2_X1    g21681(.A1(new_n24068_), .A2(new_n12793_), .ZN(new_n24118_));
  OAI21_X1   g21682(.A1(new_n24117_), .A2(new_n24118_), .B(new_n12791_), .ZN(new_n24119_));
  NAND3_X1   g21683(.A1(new_n24119_), .A2(new_n12895_), .A3(new_n24049_), .ZN(new_n24120_));
  NAND3_X1   g21684(.A1(new_n24116_), .A2(new_n24120_), .A3(pi0789), .ZN(new_n24121_));
  NOR2_X1    g21685(.A1(new_n24028_), .A2(new_n12747_), .ZN(new_n24122_));
  INV_X1     g21686(.I(new_n24051_), .ZN(new_n24123_));
  NOR2_X1    g21687(.A1(new_n24123_), .A2(pi0626), .ZN(new_n24124_));
  OAI21_X1   g21688(.A1(new_n24124_), .A2(new_n24122_), .B(new_n12815_), .ZN(new_n24125_));
  INV_X1     g21689(.I(new_n24069_), .ZN(new_n24126_));
  NAND2_X1   g21690(.A1(new_n24027_), .A2(new_n12747_), .ZN(new_n24127_));
  OAI21_X1   g21691(.A1(new_n24123_), .A2(new_n12747_), .B(new_n24127_), .ZN(new_n24128_));
  AOI22_X1   g21692(.A1(new_n24128_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n24126_), .ZN(new_n24129_));
  NAND2_X1   g21693(.A1(new_n24129_), .A2(new_n24125_), .ZN(new_n24130_));
  AOI22_X1   g21694(.A1(new_n24121_), .A2(new_n24111_), .B1(pi0788), .B2(new_n24130_), .ZN(new_n24131_));
  OAI22_X1   g21695(.A1(new_n24131_), .A2(new_n15340_), .B1(new_n12937_), .B2(new_n24075_), .ZN(new_n24132_));
  INV_X1     g21696(.I(new_n24053_), .ZN(new_n24133_));
  NAND2_X1   g21697(.A1(new_n24133_), .A2(new_n13384_), .ZN(new_n24134_));
  NAND2_X1   g21698(.A1(new_n12943_), .A2(new_n24028_), .ZN(new_n24135_));
  NAND2_X1   g21699(.A1(new_n24134_), .A2(new_n24135_), .ZN(new_n24136_));
  NAND2_X1   g21700(.A1(new_n24070_), .A2(new_n12954_), .ZN(new_n24137_));
  NAND2_X1   g21701(.A1(new_n24137_), .A2(new_n12741_), .ZN(new_n24138_));
  NOR2_X1    g21702(.A1(new_n24027_), .A2(new_n12741_), .ZN(new_n24139_));
  INV_X1     g21703(.I(new_n24139_), .ZN(new_n24140_));
  AOI21_X1   g21704(.A1(new_n24138_), .A2(new_n24140_), .B(pi1157), .ZN(new_n24141_));
  INV_X1     g21705(.I(new_n24141_), .ZN(new_n24142_));
  NAND2_X1   g21706(.A1(new_n24027_), .A2(new_n12741_), .ZN(new_n24143_));
  OAI21_X1   g21707(.A1(new_n24137_), .A2(new_n12741_), .B(new_n24143_), .ZN(new_n24144_));
  OAI22_X1   g21708(.A1(new_n24142_), .A2(new_n12981_), .B1(new_n24144_), .B2(new_n15576_), .ZN(new_n24145_));
  AOI21_X1   g21709(.A1(new_n24136_), .A2(new_n15608_), .B(new_n24145_), .ZN(new_n24146_));
  OAI22_X1   g21710(.A1(new_n24132_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n24146_), .ZN(new_n24147_));
  NAND2_X1   g21711(.A1(new_n24147_), .A2(new_n13000_), .ZN(new_n24148_));
  AND2_X2    g21712(.A1(new_n24147_), .A2(new_n12975_), .Z(new_n24149_));
  OAI21_X1   g21713(.A1(new_n12965_), .A2(new_n24144_), .B(new_n24142_), .ZN(new_n24150_));
  NAND3_X1   g21714(.A1(new_n24070_), .A2(new_n12972_), .A3(new_n12954_), .ZN(new_n24151_));
  OAI21_X1   g21715(.A1(new_n24150_), .A2(new_n12972_), .B(new_n24151_), .ZN(new_n24152_));
  NOR2_X1    g21716(.A1(new_n24152_), .A2(new_n12975_), .ZN(new_n24153_));
  OAI21_X1   g21717(.A1(new_n24149_), .A2(new_n24153_), .B(new_n12740_), .ZN(new_n24154_));
  NOR2_X1    g21718(.A1(new_n24027_), .A2(new_n12975_), .ZN(new_n24155_));
  NOR2_X1    g21719(.A1(new_n17611_), .A2(new_n24027_), .ZN(new_n24156_));
  AOI21_X1   g21720(.A1(new_n24133_), .A2(new_n17611_), .B(new_n24156_), .ZN(new_n24157_));
  NOR2_X1    g21721(.A1(new_n24157_), .A2(pi0644), .ZN(new_n24158_));
  OAI21_X1   g21722(.A1(new_n24158_), .A2(new_n24155_), .B(pi0715), .ZN(new_n24159_));
  NAND3_X1   g21723(.A1(new_n24154_), .A2(new_n12739_), .A3(new_n24159_), .ZN(new_n24160_));
  NOR2_X1    g21724(.A1(new_n24152_), .A2(pi0644), .ZN(new_n24161_));
  AOI21_X1   g21725(.A1(new_n24147_), .A2(pi0644), .B(new_n24161_), .ZN(new_n24162_));
  NAND2_X1   g21726(.A1(new_n24028_), .A2(new_n12975_), .ZN(new_n24163_));
  OAI21_X1   g21727(.A1(new_n24157_), .A2(new_n12975_), .B(new_n24163_), .ZN(new_n24164_));
  AOI21_X1   g21728(.A1(new_n24164_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n24165_));
  OAI21_X1   g21729(.A1(new_n24162_), .A2(new_n12740_), .B(new_n24165_), .ZN(new_n24166_));
  NAND3_X1   g21730(.A1(new_n24160_), .A2(pi0790), .A3(new_n24166_), .ZN(new_n24167_));
  AOI21_X1   g21731(.A1(new_n24167_), .A2(new_n24148_), .B(new_n12738_), .ZN(new_n24168_));
  AOI21_X1   g21732(.A1(po1038), .A2(new_n12494_), .B(pi0832), .ZN(new_n24169_));
  NOR2_X1    g21733(.A1(new_n13193_), .A2(pi0194), .ZN(new_n24170_));
  AOI21_X1   g21734(.A1(new_n24170_), .A2(pi0644), .B(new_n12740_), .ZN(new_n24171_));
  NOR2_X1    g21735(.A1(new_n24170_), .A2(new_n13384_), .ZN(new_n24172_));
  INV_X1     g21736(.I(new_n24172_), .ZN(new_n24173_));
  INV_X1     g21737(.I(new_n24170_), .ZN(new_n24174_));
  NOR2_X1    g21738(.A1(new_n2609_), .A2(new_n12494_), .ZN(new_n24175_));
  INV_X1     g21739(.I(new_n24175_), .ZN(new_n24176_));
  OAI21_X1   g21740(.A1(new_n15012_), .A2(new_n15011_), .B(new_n12494_), .ZN(new_n24177_));
  NAND3_X1   g21741(.A1(new_n18324_), .A2(pi0194), .A3(new_n18326_), .ZN(new_n24178_));
  AOI21_X1   g21742(.A1(new_n24177_), .A2(new_n24178_), .B(new_n17036_), .ZN(new_n24179_));
  NOR3_X1    g21743(.A1(new_n13191_), .A2(pi0194), .A3(pi0748), .ZN(new_n24180_));
  OR3_X2     g21744(.A1(new_n24179_), .A2(new_n2610_), .A3(new_n24180_), .Z(new_n24181_));
  NAND2_X1   g21745(.A1(new_n24181_), .A2(new_n24176_), .ZN(new_n24182_));
  NAND2_X1   g21746(.A1(new_n24182_), .A2(new_n12761_), .ZN(new_n24183_));
  INV_X1     g21747(.I(new_n24183_), .ZN(new_n24184_));
  NOR2_X1    g21748(.A1(new_n24170_), .A2(new_n12761_), .ZN(new_n24185_));
  NOR3_X1    g21749(.A1(new_n24184_), .A2(pi0785), .A3(new_n24185_), .ZN(new_n24186_));
  OAI22_X1   g21750(.A1(new_n24183_), .A2(pi0609), .B1(new_n13353_), .B2(new_n24170_), .ZN(new_n24187_));
  NAND2_X1   g21751(.A1(new_n24187_), .A2(new_n12770_), .ZN(new_n24188_));
  AOI22_X1   g21752(.A1(new_n24184_), .A2(pi0609), .B1(new_n13357_), .B2(new_n24174_), .ZN(new_n24189_));
  NOR2_X1    g21753(.A1(new_n24189_), .A2(new_n12770_), .ZN(new_n24190_));
  NOR2_X1    g21754(.A1(new_n24190_), .A2(new_n12764_), .ZN(new_n24191_));
  AOI21_X1   g21755(.A1(new_n24191_), .A2(new_n24188_), .B(new_n24186_), .ZN(new_n24192_));
  NOR2_X1    g21756(.A1(new_n24170_), .A2(new_n12781_), .ZN(new_n24193_));
  AOI21_X1   g21757(.A1(new_n24192_), .A2(new_n12781_), .B(new_n24193_), .ZN(new_n24194_));
  NOR2_X1    g21758(.A1(new_n24194_), .A2(pi1154), .ZN(new_n24195_));
  NOR2_X1    g21759(.A1(new_n24170_), .A2(pi0618), .ZN(new_n24196_));
  AOI21_X1   g21760(.A1(new_n24192_), .A2(pi0618), .B(new_n24196_), .ZN(new_n24197_));
  OAI21_X1   g21761(.A1(new_n24197_), .A2(new_n12785_), .B(pi0781), .ZN(new_n24198_));
  OAI22_X1   g21762(.A1(new_n24198_), .A2(new_n24195_), .B1(pi0781), .B2(new_n24192_), .ZN(new_n24199_));
  NAND2_X1   g21763(.A1(new_n24199_), .A2(new_n12796_), .ZN(new_n24200_));
  NAND2_X1   g21764(.A1(new_n24174_), .A2(pi0619), .ZN(new_n24201_));
  OAI21_X1   g21765(.A1(new_n24199_), .A2(pi0619), .B(new_n24201_), .ZN(new_n24202_));
  NAND2_X1   g21766(.A1(new_n24202_), .A2(new_n12791_), .ZN(new_n24203_));
  NAND2_X1   g21767(.A1(new_n24174_), .A2(new_n12793_), .ZN(new_n24204_));
  OAI21_X1   g21768(.A1(new_n24199_), .A2(new_n12793_), .B(new_n24204_), .ZN(new_n24205_));
  AOI21_X1   g21769(.A1(new_n24205_), .A2(pi1159), .B(new_n12796_), .ZN(new_n24206_));
  NAND2_X1   g21770(.A1(new_n24206_), .A2(new_n24203_), .ZN(new_n24207_));
  AND3_X2    g21771(.A1(new_n24207_), .A2(new_n17504_), .A3(new_n24200_), .Z(new_n24208_));
  AOI21_X1   g21772(.A1(new_n12818_), .A2(new_n24174_), .B(new_n24208_), .ZN(new_n24209_));
  OAI21_X1   g21773(.A1(new_n24209_), .A2(new_n12943_), .B(new_n24173_), .ZN(new_n24210_));
  NAND2_X1   g21774(.A1(new_n24170_), .A2(new_n12984_), .ZN(new_n24211_));
  OAI21_X1   g21775(.A1(new_n24210_), .A2(new_n12984_), .B(new_n24211_), .ZN(new_n24212_));
  NAND2_X1   g21776(.A1(new_n24212_), .A2(new_n12975_), .ZN(new_n24213_));
  AOI21_X1   g21777(.A1(new_n24213_), .A2(new_n24171_), .B(pi1160), .ZN(new_n24214_));
  NOR2_X1    g21778(.A1(new_n24174_), .A2(new_n12870_), .ZN(new_n24215_));
  NAND2_X1   g21779(.A1(new_n18371_), .A2(pi0194), .ZN(new_n24216_));
  AOI22_X1   g21780(.A1(new_n14118_), .A2(new_n3265_), .B1(new_n12825_), .B2(new_n16468_), .ZN(new_n24217_));
  OAI21_X1   g21781(.A1(new_n24217_), .A2(pi0194), .B(pi0730), .ZN(new_n24218_));
  NAND3_X1   g21782(.A1(new_n13395_), .A2(new_n12494_), .A3(new_n24056_), .ZN(new_n24219_));
  NAND3_X1   g21783(.A1(new_n24218_), .A2(new_n24219_), .A3(new_n2609_), .ZN(new_n24220_));
  NAND2_X1   g21784(.A1(new_n24220_), .A2(new_n24216_), .ZN(new_n24221_));
  NAND2_X1   g21785(.A1(new_n24221_), .A2(new_n13521_), .ZN(new_n24222_));
  NAND2_X1   g21786(.A1(new_n24174_), .A2(pi0625), .ZN(new_n24223_));
  AOI21_X1   g21787(.A1(new_n24222_), .A2(new_n24223_), .B(pi1153), .ZN(new_n24224_));
  AOI21_X1   g21788(.A1(new_n24220_), .A2(new_n24216_), .B(new_n13521_), .ZN(new_n24225_));
  NOR2_X1    g21789(.A1(new_n24170_), .A2(pi0625), .ZN(new_n24226_));
  OAI21_X1   g21790(.A1(new_n24225_), .A2(new_n24226_), .B(pi1153), .ZN(new_n24227_));
  NAND2_X1   g21791(.A1(new_n24227_), .A2(pi0778), .ZN(new_n24228_));
  OAI22_X1   g21792(.A1(new_n24228_), .A2(new_n24224_), .B1(pi0778), .B2(new_n24221_), .ZN(new_n24229_));
  AOI21_X1   g21793(.A1(new_n24229_), .A2(new_n12870_), .B(new_n24215_), .ZN(new_n24230_));
  NOR2_X1    g21794(.A1(new_n24170_), .A2(new_n12888_), .ZN(new_n24231_));
  AOI21_X1   g21795(.A1(new_n24230_), .A2(new_n12888_), .B(new_n24231_), .ZN(new_n24232_));
  NOR2_X1    g21796(.A1(new_n24174_), .A2(new_n12911_), .ZN(new_n24233_));
  AOI21_X1   g21797(.A1(new_n24232_), .A2(new_n12911_), .B(new_n24233_), .ZN(new_n24234_));
  NAND2_X1   g21798(.A1(new_n24234_), .A2(new_n13392_), .ZN(new_n24235_));
  OAI21_X1   g21799(.A1(new_n13392_), .A2(new_n24170_), .B(new_n24235_), .ZN(new_n24236_));
  NAND2_X1   g21800(.A1(new_n24236_), .A2(new_n12920_), .ZN(new_n24237_));
  NAND2_X1   g21801(.A1(new_n24174_), .A2(pi0628), .ZN(new_n24238_));
  AOI21_X1   g21802(.A1(new_n24237_), .A2(new_n24238_), .B(pi1156), .ZN(new_n24239_));
  NAND2_X1   g21803(.A1(new_n24174_), .A2(new_n12920_), .ZN(new_n24240_));
  NAND2_X1   g21804(.A1(new_n24236_), .A2(pi0628), .ZN(new_n24241_));
  AOI21_X1   g21805(.A1(new_n24241_), .A2(new_n24240_), .B(new_n12742_), .ZN(new_n24242_));
  NOR3_X1    g21806(.A1(new_n24242_), .A2(new_n24239_), .A3(new_n12937_), .ZN(new_n24243_));
  NOR2_X1    g21807(.A1(new_n24236_), .A2(pi0792), .ZN(new_n24244_));
  NOR2_X1    g21808(.A1(new_n24243_), .A2(new_n24244_), .ZN(new_n24245_));
  NAND2_X1   g21809(.A1(new_n24245_), .A2(new_n12741_), .ZN(new_n24246_));
  NAND2_X1   g21810(.A1(new_n24174_), .A2(pi0647), .ZN(new_n24247_));
  AOI21_X1   g21811(.A1(new_n24246_), .A2(new_n24247_), .B(pi1157), .ZN(new_n24248_));
  NAND2_X1   g21812(.A1(new_n24245_), .A2(pi0647), .ZN(new_n24249_));
  OAI21_X1   g21813(.A1(pi0647), .A2(new_n24170_), .B(new_n24249_), .ZN(new_n24250_));
  NAND2_X1   g21814(.A1(new_n24250_), .A2(pi1157), .ZN(new_n24251_));
  NAND2_X1   g21815(.A1(new_n24251_), .A2(pi0787), .ZN(new_n24252_));
  OAI22_X1   g21816(.A1(new_n24252_), .A2(new_n24248_), .B1(pi0787), .B2(new_n24245_), .ZN(new_n24253_));
  AOI21_X1   g21817(.A1(new_n24253_), .A2(pi0644), .B(pi0715), .ZN(new_n24254_));
  NOR2_X1    g21818(.A1(new_n24239_), .A2(new_n12919_), .ZN(new_n24255_));
  AOI21_X1   g21819(.A1(new_n24209_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n24256_));
  AOI21_X1   g21820(.A1(new_n24174_), .A2(new_n12747_), .B(pi0641), .ZN(new_n24257_));
  NAND3_X1   g21821(.A1(new_n24207_), .A2(pi0626), .A3(new_n24200_), .ZN(new_n24258_));
  AOI21_X1   g21822(.A1(new_n24258_), .A2(new_n24257_), .B(new_n12745_), .ZN(new_n24259_));
  AOI21_X1   g21823(.A1(new_n24234_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n24260_));
  OAI21_X1   g21824(.A1(new_n15111_), .A2(pi0194), .B(pi0748), .ZN(new_n24261_));
  NOR3_X1    g21825(.A1(new_n15116_), .A2(new_n12494_), .A3(new_n15113_), .ZN(new_n24262_));
  OAI21_X1   g21826(.A1(new_n24262_), .A2(new_n24261_), .B(pi0730), .ZN(new_n24263_));
  AOI21_X1   g21827(.A1(new_n15121_), .A2(new_n18421_), .B(new_n12494_), .ZN(new_n24264_));
  AOI21_X1   g21828(.A1(new_n15129_), .A2(new_n15126_), .B(pi0194), .ZN(new_n24265_));
  NOR3_X1    g21829(.A1(new_n24265_), .A2(pi0748), .A3(new_n24264_), .ZN(new_n24266_));
  NOR2_X1    g21830(.A1(new_n24263_), .A2(new_n24266_), .ZN(new_n24267_));
  OAI21_X1   g21831(.A1(new_n24179_), .A2(new_n24180_), .B(new_n24056_), .ZN(new_n24268_));
  NAND2_X1   g21832(.A1(new_n24268_), .A2(new_n2609_), .ZN(new_n24269_));
  OAI21_X1   g21833(.A1(new_n24267_), .A2(new_n24269_), .B(new_n24176_), .ZN(new_n24270_));
  NAND2_X1   g21834(.A1(new_n24270_), .A2(pi0625), .ZN(new_n24271_));
  NAND2_X1   g21835(.A1(new_n24182_), .A2(new_n13521_), .ZN(new_n24272_));
  AOI21_X1   g21836(.A1(new_n24271_), .A2(new_n24272_), .B(new_n12841_), .ZN(new_n24273_));
  NOR3_X1    g21837(.A1(new_n24273_), .A2(new_n13560_), .A3(new_n24224_), .ZN(new_n24274_));
  AOI21_X1   g21838(.A1(new_n24181_), .A2(new_n24176_), .B(new_n13521_), .ZN(new_n24275_));
  AOI21_X1   g21839(.A1(new_n24270_), .A2(new_n13521_), .B(new_n24275_), .ZN(new_n24276_));
  OAI21_X1   g21840(.A1(new_n24276_), .A2(pi1153), .B(new_n24227_), .ZN(new_n24277_));
  OAI21_X1   g21841(.A1(new_n24277_), .A2(pi0608), .B(pi0778), .ZN(new_n24278_));
  NAND2_X1   g21842(.A1(new_n24270_), .A2(new_n12758_), .ZN(new_n24279_));
  OAI21_X1   g21843(.A1(new_n24278_), .A2(new_n24274_), .B(new_n24279_), .ZN(new_n24280_));
  NAND2_X1   g21844(.A1(new_n24280_), .A2(new_n12764_), .ZN(new_n24281_));
  INV_X1     g21845(.I(new_n24281_), .ZN(new_n24282_));
  AOI21_X1   g21846(.A1(new_n24187_), .A2(new_n12770_), .B(new_n13829_), .ZN(new_n24283_));
  AOI21_X1   g21847(.A1(new_n24229_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n24284_));
  OAI21_X1   g21848(.A1(new_n24280_), .A2(new_n12766_), .B(new_n24284_), .ZN(new_n24285_));
  NAND2_X1   g21849(.A1(new_n24285_), .A2(new_n24283_), .ZN(new_n24286_));
  NOR2_X1    g21850(.A1(new_n24190_), .A2(pi0660), .ZN(new_n24287_));
  AOI21_X1   g21851(.A1(new_n24229_), .A2(pi0609), .B(pi1155), .ZN(new_n24288_));
  OAI21_X1   g21852(.A1(new_n24280_), .A2(pi0609), .B(new_n24288_), .ZN(new_n24289_));
  AOI21_X1   g21853(.A1(new_n24289_), .A2(new_n24287_), .B(new_n12764_), .ZN(new_n24290_));
  AOI21_X1   g21854(.A1(new_n24290_), .A2(new_n24286_), .B(new_n24282_), .ZN(new_n24291_));
  OR2_X2     g21855(.A1(new_n24291_), .A2(pi0781), .Z(new_n24292_));
  OAI21_X1   g21856(.A1(new_n24194_), .A2(pi1154), .B(pi0627), .ZN(new_n24293_));
  NOR2_X1    g21857(.A1(new_n24230_), .A2(pi0618), .ZN(new_n24294_));
  NOR2_X1    g21858(.A1(new_n24294_), .A2(new_n12785_), .ZN(new_n24295_));
  NAND2_X1   g21859(.A1(new_n24291_), .A2(pi0618), .ZN(new_n24296_));
  AOI21_X1   g21860(.A1(new_n24296_), .A2(new_n24295_), .B(new_n24293_), .ZN(new_n24297_));
  OAI21_X1   g21861(.A1(new_n24197_), .A2(new_n12785_), .B(new_n12880_), .ZN(new_n24298_));
  OAI21_X1   g21862(.A1(new_n24230_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n24299_));
  AOI21_X1   g21863(.A1(new_n24291_), .A2(new_n12781_), .B(new_n24299_), .ZN(new_n24300_));
  OAI21_X1   g21864(.A1(new_n24300_), .A2(new_n24298_), .B(pi0781), .ZN(new_n24301_));
  OAI21_X1   g21865(.A1(new_n24301_), .A2(new_n24297_), .B(new_n24292_), .ZN(new_n24302_));
  AND2_X2    g21866(.A1(new_n24302_), .A2(new_n12796_), .Z(new_n24303_));
  AOI21_X1   g21867(.A1(new_n24202_), .A2(new_n12791_), .B(new_n12895_), .ZN(new_n24304_));
  AOI21_X1   g21868(.A1(new_n24232_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n24305_));
  OAI21_X1   g21869(.A1(new_n24302_), .A2(new_n12793_), .B(new_n24305_), .ZN(new_n24306_));
  NAND2_X1   g21870(.A1(new_n24306_), .A2(new_n24304_), .ZN(new_n24307_));
  AOI21_X1   g21871(.A1(new_n24205_), .A2(pi1159), .B(pi0648), .ZN(new_n24308_));
  AOI21_X1   g21872(.A1(new_n24232_), .A2(pi0619), .B(pi1159), .ZN(new_n24309_));
  OAI21_X1   g21873(.A1(new_n24302_), .A2(pi0619), .B(new_n24309_), .ZN(new_n24310_));
  AOI21_X1   g21874(.A1(new_n24310_), .A2(new_n24308_), .B(new_n12796_), .ZN(new_n24311_));
  AOI21_X1   g21875(.A1(new_n24311_), .A2(new_n24307_), .B(new_n24303_), .ZN(new_n24312_));
  OAI21_X1   g21876(.A1(new_n24312_), .A2(new_n12747_), .B(new_n24260_), .ZN(new_n24313_));
  NAND2_X1   g21877(.A1(new_n24313_), .A2(new_n24259_), .ZN(new_n24314_));
  AOI21_X1   g21878(.A1(new_n24174_), .A2(pi0626), .B(new_n12814_), .ZN(new_n24315_));
  NAND3_X1   g21879(.A1(new_n24207_), .A2(new_n12747_), .A3(new_n24200_), .ZN(new_n24316_));
  AOI21_X1   g21880(.A1(new_n24316_), .A2(new_n24315_), .B(pi1158), .ZN(new_n24317_));
  AOI21_X1   g21881(.A1(new_n24234_), .A2(pi0626), .B(pi0641), .ZN(new_n24318_));
  OAI21_X1   g21882(.A1(new_n24312_), .A2(pi0626), .B(new_n24318_), .ZN(new_n24319_));
  AOI21_X1   g21883(.A1(new_n24319_), .A2(new_n24317_), .B(new_n12808_), .ZN(new_n24320_));
  AND2_X2    g21884(.A1(new_n24312_), .A2(new_n12808_), .Z(new_n24321_));
  AOI21_X1   g21885(.A1(new_n24320_), .A2(new_n24314_), .B(new_n24321_), .ZN(new_n24322_));
  OAI21_X1   g21886(.A1(new_n24322_), .A2(new_n12920_), .B(new_n24256_), .ZN(new_n24323_));
  NAND2_X1   g21887(.A1(new_n24323_), .A2(new_n24255_), .ZN(new_n24324_));
  NOR2_X1    g21888(.A1(new_n24242_), .A2(pi0629), .ZN(new_n24325_));
  AOI21_X1   g21889(.A1(new_n24209_), .A2(pi0628), .B(pi1156), .ZN(new_n24326_));
  OAI21_X1   g21890(.A1(new_n24322_), .A2(pi0628), .B(new_n24326_), .ZN(new_n24327_));
  AOI21_X1   g21891(.A1(new_n24327_), .A2(new_n24325_), .B(new_n12937_), .ZN(new_n24328_));
  AND2_X2    g21892(.A1(new_n24322_), .A2(new_n12937_), .Z(new_n24329_));
  AOI21_X1   g21893(.A1(new_n24328_), .A2(new_n24324_), .B(new_n24329_), .ZN(new_n24330_));
  OR2_X2     g21894(.A1(new_n24330_), .A2(pi0787), .Z(new_n24331_));
  OR2_X2     g21895(.A1(new_n24248_), .A2(new_n12981_), .Z(new_n24332_));
  NOR2_X1    g21896(.A1(new_n24210_), .A2(pi0647), .ZN(new_n24333_));
  NOR2_X1    g21897(.A1(new_n24333_), .A2(new_n12965_), .ZN(new_n24334_));
  NAND2_X1   g21898(.A1(new_n24330_), .A2(pi0647), .ZN(new_n24335_));
  AOI21_X1   g21899(.A1(new_n24335_), .A2(new_n24334_), .B(new_n24332_), .ZN(new_n24336_));
  NAND2_X1   g21900(.A1(new_n24251_), .A2(new_n12981_), .ZN(new_n24337_));
  OAI21_X1   g21901(.A1(new_n24210_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n24338_));
  AOI21_X1   g21902(.A1(new_n24330_), .A2(new_n12741_), .B(new_n24338_), .ZN(new_n24339_));
  OAI21_X1   g21903(.A1(new_n24339_), .A2(new_n24337_), .B(pi0787), .ZN(new_n24340_));
  OAI21_X1   g21904(.A1(new_n24340_), .A2(new_n24336_), .B(new_n24331_), .ZN(new_n24341_));
  OAI21_X1   g21905(.A1(new_n24341_), .A2(pi0644), .B(new_n24254_), .ZN(new_n24342_));
  NAND2_X1   g21906(.A1(new_n24342_), .A2(new_n24214_), .ZN(new_n24343_));
  AOI21_X1   g21907(.A1(new_n24170_), .A2(new_n12975_), .B(pi0715), .ZN(new_n24344_));
  NAND2_X1   g21908(.A1(new_n24212_), .A2(pi0644), .ZN(new_n24345_));
  AOI21_X1   g21909(.A1(new_n24345_), .A2(new_n24344_), .B(new_n12739_), .ZN(new_n24346_));
  NOR2_X1    g21910(.A1(new_n24253_), .A2(pi0644), .ZN(new_n24347_));
  AOI21_X1   g21911(.A1(new_n24341_), .A2(pi0644), .B(new_n24347_), .ZN(new_n24348_));
  OAI21_X1   g21912(.A1(new_n24348_), .A2(new_n12740_), .B(new_n24346_), .ZN(new_n24349_));
  NAND3_X1   g21913(.A1(new_n24349_), .A2(new_n24343_), .A3(pi0790), .ZN(new_n24350_));
  AOI21_X1   g21914(.A1(new_n24341_), .A2(new_n13000_), .B(po1038), .ZN(new_n24351_));
  NAND2_X1   g21915(.A1(new_n24350_), .A2(new_n24351_), .ZN(new_n24352_));
  AOI21_X1   g21916(.A1(new_n24352_), .A2(new_n24169_), .B(new_n24168_), .ZN(po0351));
  OAI22_X1   g21917(.A1(new_n12697_), .A2(new_n3932_), .B1(new_n7814_), .B2(new_n12401_), .ZN(new_n24354_));
  OAI21_X1   g21918(.A1(new_n12631_), .A2(pi0192), .B(pi0232), .ZN(new_n24355_));
  AOI21_X1   g21919(.A1(new_n24354_), .A2(pi0299), .B(new_n24355_), .ZN(new_n24356_));
  NAND2_X1   g21920(.A1(new_n12643_), .A2(pi0192), .ZN(new_n24357_));
  AOI21_X1   g21921(.A1(new_n24356_), .A2(new_n24357_), .B(new_n12634_), .ZN(new_n24358_));
  NOR2_X1    g21922(.A1(new_n12648_), .A2(pi0192), .ZN(new_n24359_));
  NOR2_X1    g21923(.A1(new_n12658_), .A2(new_n12412_), .ZN(new_n24360_));
  AOI21_X1   g21924(.A1(new_n3932_), .A2(new_n7627_), .B(new_n12660_), .ZN(new_n24361_));
  NOR2_X1    g21925(.A1(new_n24361_), .A2(new_n8070_), .ZN(new_n24362_));
  OAI22_X1   g21926(.A1(new_n24360_), .A2(new_n24359_), .B1(new_n7637_), .B2(new_n24362_), .ZN(new_n24363_));
  AOI21_X1   g21927(.A1(new_n24363_), .A2(pi0232), .B(new_n12653_), .ZN(new_n24364_));
  OAI21_X1   g21928(.A1(new_n24364_), .A2(new_n2627_), .B(new_n3270_), .ZN(new_n24365_));
  OAI21_X1   g21929(.A1(new_n24358_), .A2(new_n24365_), .B(new_n3458_), .ZN(new_n24366_));
  AOI21_X1   g21930(.A1(new_n24366_), .A2(new_n12696_), .B(pi0092), .ZN(new_n24367_));
  OAI21_X1   g21931(.A1(new_n24367_), .A2(new_n12695_), .B(new_n2602_), .ZN(new_n24368_));
  AOI21_X1   g21932(.A1(new_n24368_), .A2(new_n12627_), .B(new_n2471_), .ZN(new_n24369_));
  NOR3_X1    g21933(.A1(new_n12625_), .A2(pi0138), .A3(pi0139), .ZN(new_n24370_));
  AOI21_X1   g21934(.A1(new_n24370_), .A2(new_n12690_), .B(new_n12689_), .ZN(new_n24371_));
  NAND2_X1   g21935(.A1(new_n8103_), .A2(new_n24371_), .ZN(new_n24372_));
  INV_X1     g21936(.I(new_n24371_), .ZN(new_n24373_));
  OAI21_X1   g21937(.A1(new_n12683_), .A2(new_n12415_), .B(new_n2627_), .ZN(new_n24374_));
  NAND2_X1   g21938(.A1(new_n6745_), .A2(new_n12411_), .ZN(new_n24375_));
  NOR2_X1    g21939(.A1(new_n9241_), .A2(pi0192), .ZN(new_n24376_));
  NOR2_X1    g21940(.A1(new_n12675_), .A2(new_n12412_), .ZN(new_n24377_));
  OAI21_X1   g21941(.A1(new_n24377_), .A2(new_n24376_), .B(new_n2628_), .ZN(new_n24378_));
  NAND4_X1   g21942(.A1(new_n24378_), .A2(pi0232), .A3(new_n12721_), .A4(new_n24375_), .ZN(new_n24379_));
  NAND3_X1   g21943(.A1(new_n24379_), .A2(pi0039), .A3(new_n12720_), .ZN(new_n24380_));
  NAND4_X1   g21944(.A1(new_n24380_), .A2(new_n8280_), .A3(new_n24373_), .A4(new_n24374_), .ZN(new_n24381_));
  OAI21_X1   g21945(.A1(new_n24369_), .A2(new_n24372_), .B(new_n24381_), .ZN(po0352));
  AOI21_X1   g21946(.A1(new_n4089_), .A2(new_n7627_), .B(new_n12660_), .ZN(new_n24383_));
  OAI21_X1   g21947(.A1(new_n24383_), .A2(new_n8070_), .B(new_n7620_), .ZN(new_n24384_));
  AOI21_X1   g21948(.A1(new_n24384_), .A2(new_n12654_), .B(new_n5666_), .ZN(new_n24385_));
  OAI21_X1   g21949(.A1(new_n24385_), .A2(new_n12653_), .B(pi0039), .ZN(new_n24386_));
  NAND3_X1   g21950(.A1(new_n24386_), .A2(new_n3265_), .A3(new_n12494_), .ZN(new_n24387_));
  NOR2_X1    g21951(.A1(new_n24385_), .A2(new_n12653_), .ZN(new_n24388_));
  NAND2_X1   g21952(.A1(new_n12658_), .A2(pi0232), .ZN(new_n24389_));
  AOI21_X1   g21953(.A1(new_n24388_), .A2(new_n24389_), .B(new_n2627_), .ZN(new_n24390_));
  NOR3_X1    g21954(.A1(new_n24390_), .A2(pi0038), .A3(new_n12494_), .ZN(new_n24391_));
  INV_X1     g21955(.I(new_n24391_), .ZN(new_n24392_));
  OAI22_X1   g21956(.A1(new_n12643_), .A2(new_n24392_), .B1(new_n12630_), .B2(new_n24387_), .ZN(new_n24393_));
  NAND2_X1   g21957(.A1(new_n7691_), .A2(new_n12491_), .ZN(new_n24394_));
  NAND2_X1   g21958(.A1(new_n7814_), .A2(new_n12492_), .ZN(new_n24395_));
  NAND3_X1   g21959(.A1(new_n24395_), .A2(pi0299), .A3(new_n24394_), .ZN(new_n24396_));
  AND3_X2    g21960(.A1(new_n24393_), .A2(pi0232), .A3(new_n24396_), .Z(new_n24397_));
  AOI21_X1   g21961(.A1(new_n24387_), .A2(new_n24392_), .B(new_n12635_), .ZN(new_n24398_));
  OAI21_X1   g21962(.A1(new_n24398_), .A2(new_n24397_), .B(new_n2702_), .ZN(new_n24399_));
  AOI21_X1   g21963(.A1(new_n24399_), .A2(new_n3458_), .B(new_n12629_), .ZN(new_n24400_));
  OAI21_X1   g21964(.A1(new_n24400_), .A2(pi0092), .B(new_n12669_), .ZN(new_n24401_));
  AOI21_X1   g21965(.A1(new_n24401_), .A2(new_n2602_), .B(new_n12628_), .ZN(new_n24402_));
  OAI21_X1   g21966(.A1(new_n24402_), .A2(new_n2471_), .B(new_n8103_), .ZN(new_n24403_));
  NOR2_X1    g21967(.A1(new_n24403_), .A2(new_n12690_), .ZN(new_n24404_));
  NOR2_X1    g21968(.A1(new_n8159_), .A2(pi0170), .ZN(new_n24405_));
  OAI21_X1   g21969(.A1(new_n24405_), .A2(new_n12673_), .B(new_n10332_), .ZN(new_n24406_));
  NOR2_X1    g21970(.A1(new_n12674_), .A2(new_n10849_), .ZN(new_n24407_));
  INV_X1     g21971(.I(new_n24407_), .ZN(new_n24408_));
  AOI21_X1   g21972(.A1(new_n24406_), .A2(new_n24408_), .B(new_n5666_), .ZN(new_n24409_));
  NOR2_X1    g21973(.A1(new_n24409_), .A2(new_n12719_), .ZN(new_n24410_));
  AOI21_X1   g21974(.A1(new_n24410_), .A2(pi0299), .B(new_n9242_), .ZN(new_n24411_));
  AND2_X2    g21975(.A1(new_n24411_), .A2(pi0039), .Z(new_n24412_));
  NOR3_X1    g21976(.A1(new_n12683_), .A2(pi0039), .A3(new_n12493_), .ZN(new_n24413_));
  NOR3_X1    g21977(.A1(new_n24412_), .A2(pi0194), .A3(new_n24413_), .ZN(new_n24414_));
  NOR2_X1    g21978(.A1(new_n24410_), .A2(new_n2627_), .ZN(new_n24415_));
  NOR3_X1    g21979(.A1(new_n12683_), .A2(pi0039), .A3(new_n12501_), .ZN(new_n24416_));
  NOR3_X1    g21980(.A1(new_n24415_), .A2(new_n12494_), .A3(new_n24416_), .ZN(new_n24417_));
  NOR3_X1    g21981(.A1(new_n24414_), .A2(new_n8281_), .A3(new_n24417_), .ZN(new_n24418_));
  AOI21_X1   g21982(.A1(new_n12690_), .A2(new_n24418_), .B(new_n24404_), .ZN(new_n24419_));
  NAND2_X1   g21983(.A1(new_n12690_), .A2(pi0195), .ZN(new_n24420_));
  NAND2_X1   g21984(.A1(new_n24418_), .A2(new_n24420_), .ZN(new_n24421_));
  OAI21_X1   g21985(.A1(new_n24403_), .A2(new_n24420_), .B(new_n24421_), .ZN(new_n24422_));
  NAND2_X1   g21986(.A1(new_n24422_), .A2(new_n24370_), .ZN(new_n24423_));
  OAI21_X1   g21987(.A1(new_n24419_), .A2(new_n24370_), .B(new_n24423_), .ZN(po0353));
  NOR2_X1    g21988(.A1(new_n16175_), .A2(new_n5636_), .ZN(new_n24425_));
  AOI21_X1   g21989(.A1(new_n16052_), .A2(new_n5636_), .B(new_n24425_), .ZN(new_n24426_));
  NAND2_X1   g21990(.A1(new_n16015_), .A2(new_n5636_), .ZN(new_n24427_));
  AOI21_X1   g21991(.A1(new_n24427_), .A2(new_n16025_), .B(new_n15782_), .ZN(new_n24428_));
  NOR2_X1    g21992(.A1(new_n16010_), .A2(pi0197), .ZN(new_n24429_));
  NOR2_X1    g21993(.A1(new_n16032_), .A2(new_n5636_), .ZN(new_n24430_));
  OAI21_X1   g21994(.A1(new_n24429_), .A2(new_n24430_), .B(pi0299), .ZN(new_n24431_));
  AOI21_X1   g21995(.A1(new_n24431_), .A2(new_n24428_), .B(new_n2627_), .ZN(new_n24432_));
  OAI21_X1   g21996(.A1(new_n24426_), .A2(pi0767), .B(new_n24432_), .ZN(new_n24433_));
  NOR2_X1    g21997(.A1(new_n5692_), .A2(pi0767), .ZN(new_n24434_));
  NOR2_X1    g21998(.A1(new_n13060_), .A2(new_n24434_), .ZN(new_n24435_));
  NOR2_X1    g21999(.A1(new_n16102_), .A2(new_n5636_), .ZN(new_n24436_));
  OAI21_X1   g22000(.A1(new_n24436_), .A2(new_n24435_), .B(new_n2627_), .ZN(new_n24437_));
  OR2_X2     g22001(.A1(new_n24437_), .A2(new_n16023_), .Z(new_n24438_));
  AOI21_X1   g22002(.A1(new_n24433_), .A2(new_n24438_), .B(pi0038), .ZN(new_n24439_));
  NOR2_X1    g22003(.A1(new_n15782_), .A2(new_n5692_), .ZN(new_n24440_));
  NOR3_X1    g22004(.A1(new_n16186_), .A2(pi0039), .A3(new_n24440_), .ZN(new_n24441_));
  OAI21_X1   g22005(.A1(new_n13344_), .A2(pi0197), .B(pi0038), .ZN(new_n24442_));
  OAI21_X1   g22006(.A1(new_n24441_), .A2(new_n24442_), .B(new_n15577_), .ZN(new_n24443_));
  NOR2_X1    g22007(.A1(new_n15782_), .A2(pi0197), .ZN(new_n24444_));
  AOI21_X1   g22008(.A1(new_n14065_), .A2(new_n24444_), .B(new_n2627_), .ZN(new_n24445_));
  NOR2_X1    g22009(.A1(new_n16646_), .A2(new_n5636_), .ZN(new_n24446_));
  NOR2_X1    g22010(.A1(new_n16114_), .A2(pi0197), .ZN(new_n24447_));
  OAI21_X1   g22011(.A1(new_n24447_), .A2(new_n24446_), .B(pi0299), .ZN(new_n24448_));
  NAND2_X1   g22012(.A1(new_n16086_), .A2(new_n24427_), .ZN(new_n24449_));
  NAND3_X1   g22013(.A1(new_n24448_), .A2(new_n15782_), .A3(new_n24449_), .ZN(new_n24450_));
  AOI21_X1   g22014(.A1(new_n24450_), .A2(new_n24445_), .B(pi0038), .ZN(new_n24451_));
  INV_X1     g22015(.I(new_n24434_), .ZN(new_n24452_));
  AOI21_X1   g22016(.A1(new_n13344_), .A2(new_n24452_), .B(new_n3265_), .ZN(new_n24453_));
  NAND2_X1   g22017(.A1(new_n16073_), .A2(pi0197), .ZN(new_n24454_));
  AOI22_X1   g22018(.A1(new_n24451_), .A2(new_n24437_), .B1(new_n24453_), .B2(new_n24454_), .ZN(new_n24455_));
  OAI22_X1   g22019(.A1(new_n24455_), .A2(new_n15577_), .B1(new_n24439_), .B2(new_n24443_), .ZN(new_n24456_));
  NAND2_X1   g22020(.A1(new_n8265_), .A2(pi0197), .ZN(new_n24457_));
  OAI21_X1   g22021(.A1(new_n24456_), .A2(new_n8265_), .B(new_n24457_), .ZN(new_n24458_));
  NAND2_X1   g22022(.A1(new_n15936_), .A2(new_n15577_), .ZN(new_n24459_));
  NAND3_X1   g22023(.A1(new_n24459_), .A2(new_n24452_), .A3(new_n3042_), .ZN(new_n24460_));
  NAND2_X1   g22024(.A1(new_n3043_), .A2(pi0197), .ZN(new_n24461_));
  AOI21_X1   g22025(.A1(new_n24460_), .A2(new_n24461_), .B(new_n12738_), .ZN(new_n24462_));
  AOI21_X1   g22026(.A1(new_n24458_), .A2(new_n12738_), .B(new_n24462_), .ZN(po0354));
  OAI21_X1   g22027(.A1(new_n16102_), .A2(new_n2573_), .B(new_n14460_), .ZN(new_n24464_));
  NOR2_X1    g22028(.A1(new_n13150_), .A2(new_n2672_), .ZN(new_n24465_));
  NOR2_X1    g22029(.A1(new_n13098_), .A2(new_n2672_), .ZN(new_n24466_));
  OAI21_X1   g22030(.A1(po1101), .A2(new_n24466_), .B(new_n24465_), .ZN(new_n24467_));
  OAI21_X1   g22031(.A1(new_n13149_), .A2(new_n5724_), .B(new_n13484_), .ZN(new_n24468_));
  NOR2_X1    g22032(.A1(new_n24468_), .A2(new_n2672_), .ZN(new_n24469_));
  NAND2_X1   g22033(.A1(new_n24469_), .A2(new_n6764_), .ZN(new_n24470_));
  AOI21_X1   g22034(.A1(new_n24470_), .A2(new_n24467_), .B(new_n2436_), .ZN(new_n24471_));
  OAI21_X1   g22035(.A1(new_n24466_), .A2(new_n3304_), .B(new_n2436_), .ZN(new_n24472_));
  OAI21_X1   g22036(.A1(new_n13226_), .A2(new_n2672_), .B(new_n6764_), .ZN(new_n24473_));
  NOR2_X1    g22037(.A1(new_n13098_), .A2(po1101), .ZN(new_n24474_));
  AOI21_X1   g22038(.A1(new_n13109_), .A2(po1101), .B(new_n24474_), .ZN(new_n24475_));
  OAI21_X1   g22039(.A1(new_n24475_), .A2(new_n2672_), .B(new_n5422_), .ZN(new_n24476_));
  AOI21_X1   g22040(.A1(new_n24473_), .A2(new_n24476_), .B(new_n3303_), .ZN(new_n24477_));
  OAI21_X1   g22041(.A1(new_n24477_), .A2(new_n24472_), .B(pi0299), .ZN(new_n24478_));
  NOR2_X1    g22042(.A1(new_n24478_), .A2(new_n24471_), .ZN(new_n24479_));
  NAND2_X1   g22043(.A1(new_n24469_), .A2(new_n5445_), .ZN(new_n24480_));
  AOI21_X1   g22044(.A1(new_n24480_), .A2(new_n24467_), .B(new_n2668_), .ZN(new_n24481_));
  OAI21_X1   g22045(.A1(new_n24466_), .A2(new_n2642_), .B(new_n2668_), .ZN(new_n24482_));
  OAI21_X1   g22046(.A1(new_n13226_), .A2(new_n2672_), .B(new_n5445_), .ZN(new_n24483_));
  OAI21_X1   g22047(.A1(new_n24475_), .A2(new_n2672_), .B(new_n5446_), .ZN(new_n24484_));
  AOI21_X1   g22048(.A1(new_n24483_), .A2(new_n24484_), .B(new_n2641_), .ZN(new_n24485_));
  OAI21_X1   g22049(.A1(new_n24485_), .A2(new_n24482_), .B(new_n2628_), .ZN(new_n24486_));
  NOR2_X1    g22050(.A1(new_n24486_), .A2(new_n24481_), .ZN(new_n24487_));
  NOR4_X1    g22051(.A1(new_n24479_), .A2(new_n2610_), .A3(new_n24487_), .A4(new_n8896_), .ZN(new_n24488_));
  AOI21_X1   g22052(.A1(new_n24464_), .A2(pi0198), .B(new_n24488_), .ZN(new_n24489_));
  NOR2_X1    g22053(.A1(new_n2609_), .A2(new_n2672_), .ZN(new_n24490_));
  NOR2_X1    g22054(.A1(new_n2627_), .A2(pi0198), .ZN(new_n24491_));
  NOR2_X1    g22055(.A1(new_n13136_), .A2(new_n2672_), .ZN(new_n24492_));
  INV_X1     g22056(.I(pi0634), .ZN(new_n24493_));
  NOR3_X1    g22057(.A1(new_n13568_), .A2(new_n24493_), .A3(new_n12825_), .ZN(new_n24494_));
  NOR3_X1    g22058(.A1(new_n24494_), .A2(pi0039), .A3(new_n24492_), .ZN(new_n24495_));
  OAI21_X1   g22059(.A1(new_n24495_), .A2(new_n24491_), .B(pi0038), .ZN(new_n24496_));
  INV_X1     g22060(.I(new_n24496_), .ZN(new_n24497_));
  NOR2_X1    g22061(.A1(new_n24493_), .A2(new_n12821_), .ZN(new_n24498_));
  INV_X1     g22062(.I(new_n24498_), .ZN(new_n24499_));
  OAI21_X1   g22063(.A1(new_n14557_), .A2(new_n2672_), .B(new_n24499_), .ZN(new_n24500_));
  AND2_X2    g22064(.A1(new_n13248_), .A2(pi0665), .Z(new_n24501_));
  NOR2_X1    g22065(.A1(new_n14655_), .A2(pi0198), .ZN(new_n24502_));
  AOI21_X1   g22066(.A1(pi0198), .A2(new_n24501_), .B(new_n24502_), .ZN(new_n24503_));
  OR2_X2     g22067(.A1(new_n24503_), .A2(new_n24499_), .Z(new_n24504_));
  AOI21_X1   g22068(.A1(new_n24504_), .A2(new_n24500_), .B(new_n2628_), .ZN(new_n24505_));
  NAND2_X1   g22069(.A1(new_n13054_), .A2(pi0198), .ZN(new_n24506_));
  INV_X1     g22070(.I(new_n24506_), .ZN(new_n24507_));
  NAND3_X1   g22071(.A1(new_n13053_), .A2(pi0198), .A3(new_n13049_), .ZN(new_n24508_));
  NAND3_X1   g22072(.A1(new_n13409_), .A2(new_n2672_), .A3(new_n13039_), .ZN(new_n24509_));
  NAND2_X1   g22073(.A1(new_n24509_), .A2(new_n24498_), .ZN(new_n24510_));
  NOR2_X1    g22074(.A1(new_n13053_), .A2(new_n12822_), .ZN(new_n24511_));
  AOI22_X1   g22075(.A1(new_n24507_), .A2(new_n24511_), .B1(new_n24508_), .B2(new_n24510_), .ZN(new_n24512_));
  NOR2_X1    g22076(.A1(new_n24512_), .A2(pi0299), .ZN(new_n24513_));
  OAI21_X1   g22077(.A1(new_n24505_), .A2(new_n24513_), .B(new_n2627_), .ZN(new_n24514_));
  NOR2_X1    g22078(.A1(new_n13274_), .A2(new_n2672_), .ZN(new_n24515_));
  NOR3_X1    g22079(.A1(new_n13149_), .A2(new_n13420_), .A3(new_n24493_), .ZN(new_n24516_));
  NOR2_X1    g22080(.A1(new_n24515_), .A2(new_n24516_), .ZN(new_n24517_));
  NOR2_X1    g22081(.A1(new_n24517_), .A2(new_n5409_), .ZN(new_n24518_));
  INV_X1     g22082(.I(new_n24517_), .ZN(new_n24519_));
  NOR2_X1    g22083(.A1(new_n13420_), .A2(new_n24493_), .ZN(new_n24520_));
  NOR2_X1    g22084(.A1(new_n24520_), .A2(new_n24466_), .ZN(new_n24521_));
  NOR2_X1    g22085(.A1(new_n24521_), .A2(new_n5398_), .ZN(new_n24522_));
  AOI21_X1   g22086(.A1(new_n24519_), .A2(new_n5398_), .B(new_n24522_), .ZN(new_n24523_));
  NOR2_X1    g22087(.A1(new_n24523_), .A2(new_n5410_), .ZN(new_n24524_));
  OAI21_X1   g22088(.A1(new_n24524_), .A2(new_n24518_), .B(new_n13584_), .ZN(new_n24525_));
  NOR3_X1    g22089(.A1(new_n24468_), .A2(new_n2672_), .A3(pi0680), .ZN(new_n24526_));
  AOI21_X1   g22090(.A1(new_n24519_), .A2(new_n5404_), .B(new_n24526_), .ZN(new_n24527_));
  NAND2_X1   g22091(.A1(new_n24525_), .A2(new_n24527_), .ZN(new_n24528_));
  NAND2_X1   g22092(.A1(new_n24528_), .A2(new_n6764_), .ZN(new_n24529_));
  NAND2_X1   g22093(.A1(new_n24521_), .A2(new_n5398_), .ZN(new_n24530_));
  OAI21_X1   g22094(.A1(new_n24519_), .A2(new_n5398_), .B(new_n24530_), .ZN(new_n24531_));
  INV_X1     g22095(.I(new_n24521_), .ZN(new_n24532_));
  NAND2_X1   g22096(.A1(new_n24532_), .A2(new_n5409_), .ZN(new_n24533_));
  OAI21_X1   g22097(.A1(new_n24531_), .A2(new_n5409_), .B(new_n24533_), .ZN(new_n24534_));
  AOI22_X1   g22098(.A1(new_n24534_), .A2(new_n13584_), .B1(new_n24465_), .B2(new_n24526_), .ZN(new_n24535_));
  OAI21_X1   g22099(.A1(new_n5403_), .A2(new_n24531_), .B(new_n24535_), .ZN(new_n24536_));
  NAND2_X1   g22100(.A1(new_n24536_), .A2(new_n5422_), .ZN(new_n24537_));
  AOI21_X1   g22101(.A1(new_n24537_), .A2(new_n24529_), .B(new_n2436_), .ZN(new_n24538_));
  INV_X1     g22102(.I(new_n24466_), .ZN(new_n24539_));
  OAI21_X1   g22103(.A1(new_n13420_), .A2(new_n24499_), .B(new_n24539_), .ZN(new_n24540_));
  OAI21_X1   g22104(.A1(new_n24540_), .A2(new_n3304_), .B(new_n2436_), .ZN(new_n24541_));
  NAND3_X1   g22105(.A1(new_n13109_), .A2(pi0198), .A3(new_n5410_), .ZN(new_n24542_));
  NAND2_X1   g22106(.A1(new_n24466_), .A2(new_n5409_), .ZN(new_n24543_));
  AOI21_X1   g22107(.A1(new_n24542_), .A2(new_n24543_), .B(pi0680), .ZN(new_n24544_));
  INV_X1     g22108(.I(new_n13428_), .ZN(new_n24545_));
  NOR2_X1    g22109(.A1(new_n13082_), .A2(new_n2672_), .ZN(new_n24546_));
  AOI21_X1   g22110(.A1(new_n24545_), .A2(pi0634), .B(new_n24546_), .ZN(new_n24547_));
  INV_X1     g22111(.I(new_n24547_), .ZN(new_n24548_));
  OAI21_X1   g22112(.A1(new_n24548_), .A2(new_n5398_), .B(new_n24530_), .ZN(new_n24549_));
  OR2_X2     g22113(.A1(new_n24549_), .A2(new_n5409_), .Z(new_n24550_));
  AOI21_X1   g22114(.A1(new_n24550_), .A2(new_n24533_), .B(new_n13585_), .ZN(new_n24551_));
  NOR2_X1    g22115(.A1(new_n24549_), .A2(new_n5403_), .ZN(new_n24552_));
  NOR3_X1    g22116(.A1(new_n24551_), .A2(new_n24544_), .A3(new_n24552_), .ZN(new_n24553_));
  NAND2_X1   g22117(.A1(new_n24553_), .A2(new_n5422_), .ZN(new_n24554_));
  NOR3_X1    g22118(.A1(new_n13485_), .A2(new_n2672_), .A3(pi0680), .ZN(new_n24555_));
  NAND2_X1   g22119(.A1(new_n24548_), .A2(new_n5410_), .ZN(new_n24556_));
  INV_X1     g22120(.I(new_n24522_), .ZN(new_n24557_));
  OAI21_X1   g22121(.A1(new_n24547_), .A2(new_n5437_), .B(new_n24557_), .ZN(new_n24558_));
  NAND2_X1   g22122(.A1(new_n24558_), .A2(new_n5409_), .ZN(new_n24559_));
  AOI21_X1   g22123(.A1(new_n24559_), .A2(new_n24556_), .B(new_n13585_), .ZN(new_n24560_));
  NOR2_X1    g22124(.A1(new_n24547_), .A2(new_n5403_), .ZN(new_n24561_));
  NOR3_X1    g22125(.A1(new_n24560_), .A2(new_n24555_), .A3(new_n24561_), .ZN(new_n24562_));
  NAND2_X1   g22126(.A1(new_n24562_), .A2(new_n6764_), .ZN(new_n24563_));
  AOI21_X1   g22127(.A1(new_n24554_), .A2(new_n24563_), .B(new_n3303_), .ZN(new_n24564_));
  OAI21_X1   g22128(.A1(new_n24564_), .A2(new_n24541_), .B(pi0299), .ZN(new_n24565_));
  NAND2_X1   g22129(.A1(new_n24553_), .A2(new_n5446_), .ZN(new_n24566_));
  NAND2_X1   g22130(.A1(new_n24562_), .A2(new_n5445_), .ZN(new_n24567_));
  AOI21_X1   g22131(.A1(new_n24566_), .A2(new_n24567_), .B(new_n2641_), .ZN(new_n24568_));
  OAI21_X1   g22132(.A1(new_n24540_), .A2(new_n2642_), .B(new_n2668_), .ZN(new_n24569_));
  NAND2_X1   g22133(.A1(new_n24528_), .A2(new_n5445_), .ZN(new_n24570_));
  NAND2_X1   g22134(.A1(new_n24536_), .A2(new_n5446_), .ZN(new_n24571_));
  NAND2_X1   g22135(.A1(new_n24571_), .A2(new_n24570_), .ZN(new_n24572_));
  AOI21_X1   g22136(.A1(new_n24572_), .A2(pi0223), .B(pi0299), .ZN(new_n24573_));
  OAI21_X1   g22137(.A1(new_n24568_), .A2(new_n24569_), .B(new_n24573_), .ZN(new_n24574_));
  OAI21_X1   g22138(.A1(new_n24538_), .A2(new_n24565_), .B(new_n24574_), .ZN(new_n24575_));
  NAND2_X1   g22139(.A1(new_n24575_), .A2(pi0039), .ZN(new_n24576_));
  AOI21_X1   g22140(.A1(new_n24576_), .A2(new_n24514_), .B(pi0038), .ZN(new_n24577_));
  NOR3_X1    g22141(.A1(new_n24577_), .A2(new_n2610_), .A3(new_n24497_), .ZN(new_n24578_));
  NOR2_X1    g22142(.A1(new_n24578_), .A2(new_n24490_), .ZN(new_n24579_));
  INV_X1     g22143(.I(new_n24579_), .ZN(new_n24580_));
  INV_X1     g22144(.I(new_n24489_), .ZN(new_n24581_));
  NAND2_X1   g22145(.A1(new_n24581_), .A2(pi0625), .ZN(new_n24582_));
  OAI21_X1   g22146(.A1(new_n24579_), .A2(pi0625), .B(new_n24582_), .ZN(new_n24583_));
  NAND2_X1   g22147(.A1(new_n24583_), .A2(new_n12841_), .ZN(new_n24584_));
  NAND2_X1   g22148(.A1(new_n24580_), .A2(pi0625), .ZN(new_n24585_));
  NAND2_X1   g22149(.A1(new_n24581_), .A2(new_n13521_), .ZN(new_n24586_));
  AOI21_X1   g22150(.A1(new_n24585_), .A2(new_n24586_), .B(new_n12841_), .ZN(new_n24587_));
  NOR2_X1    g22151(.A1(new_n24587_), .A2(new_n12758_), .ZN(new_n24588_));
  NAND2_X1   g22152(.A1(new_n24588_), .A2(new_n24584_), .ZN(new_n24589_));
  OAI21_X1   g22153(.A1(pi0778), .A2(new_n24580_), .B(new_n24589_), .ZN(new_n24590_));
  NOR2_X1    g22154(.A1(new_n24489_), .A2(new_n12870_), .ZN(new_n24591_));
  INV_X1     g22155(.I(new_n24591_), .ZN(new_n24592_));
  OAI21_X1   g22156(.A1(new_n24590_), .A2(new_n12869_), .B(new_n24592_), .ZN(new_n24593_));
  NOR2_X1    g22157(.A1(new_n24593_), .A2(new_n12887_), .ZN(new_n24594_));
  AOI21_X1   g22158(.A1(new_n12887_), .A2(new_n24489_), .B(new_n24594_), .ZN(new_n24595_));
  NAND2_X1   g22159(.A1(new_n24595_), .A2(new_n12923_), .ZN(new_n24596_));
  OAI21_X1   g22160(.A1(new_n12923_), .A2(new_n24489_), .B(new_n24596_), .ZN(new_n24597_));
  NOR2_X1    g22161(.A1(new_n24597_), .A2(pi0792), .ZN(new_n24598_));
  NAND2_X1   g22162(.A1(new_n24597_), .A2(new_n12920_), .ZN(new_n24599_));
  NAND2_X1   g22163(.A1(new_n24581_), .A2(pi0628), .ZN(new_n24600_));
  AOI21_X1   g22164(.A1(new_n24599_), .A2(new_n24600_), .B(pi1156), .ZN(new_n24601_));
  NOR2_X1    g22165(.A1(new_n24489_), .A2(pi0628), .ZN(new_n24602_));
  AOI21_X1   g22166(.A1(new_n24597_), .A2(pi0628), .B(new_n24602_), .ZN(new_n24603_));
  NOR2_X1    g22167(.A1(new_n24603_), .A2(new_n12742_), .ZN(new_n24604_));
  NOR3_X1    g22168(.A1(new_n24604_), .A2(new_n24601_), .A3(new_n12937_), .ZN(new_n24605_));
  NOR2_X1    g22169(.A1(new_n24605_), .A2(new_n24598_), .ZN(new_n24606_));
  NAND2_X1   g22170(.A1(new_n24606_), .A2(new_n12741_), .ZN(new_n24607_));
  OAI21_X1   g22171(.A1(new_n12741_), .A2(new_n24489_), .B(new_n24607_), .ZN(new_n24608_));
  NAND2_X1   g22172(.A1(new_n24608_), .A2(new_n12965_), .ZN(new_n24609_));
  NOR2_X1    g22173(.A1(new_n24609_), .A2(new_n12981_), .ZN(new_n24610_));
  INV_X1     g22174(.I(pi0633), .ZN(new_n24611_));
  NOR3_X1    g22175(.A1(new_n13568_), .A2(new_n24611_), .A3(new_n12755_), .ZN(new_n24612_));
  NOR3_X1    g22176(.A1(new_n24612_), .A2(pi0039), .A3(new_n24492_), .ZN(new_n24613_));
  OAI21_X1   g22177(.A1(new_n24613_), .A2(new_n24491_), .B(pi0038), .ZN(new_n24614_));
  NOR2_X1    g22178(.A1(new_n13803_), .A2(new_n2672_), .ZN(new_n24615_));
  AOI21_X1   g22179(.A1(new_n2672_), .A2(new_n13201_), .B(new_n24615_), .ZN(new_n24616_));
  INV_X1     g22180(.I(new_n24616_), .ZN(new_n24617_));
  NAND2_X1   g22181(.A1(pi0603), .A2(pi0633), .ZN(new_n24618_));
  NAND3_X1   g22182(.A1(new_n13055_), .A2(pi0198), .A3(new_n24618_), .ZN(new_n24619_));
  OAI21_X1   g22183(.A1(new_n24617_), .A2(new_n24618_), .B(new_n24619_), .ZN(new_n24620_));
  NOR2_X1    g22184(.A1(new_n24620_), .A2(new_n2628_), .ZN(new_n24621_));
  AND2_X2    g22185(.A1(new_n13199_), .A2(new_n13039_), .Z(new_n24622_));
  NOR2_X1    g22186(.A1(new_n13053_), .A2(new_n2672_), .ZN(new_n24623_));
  AOI22_X1   g22187(.A1(new_n24622_), .A2(new_n2672_), .B1(pi0621), .B2(new_n24623_), .ZN(new_n24624_));
  NAND2_X1   g22188(.A1(new_n24624_), .A2(pi0633), .ZN(new_n24625_));
  NAND2_X1   g22189(.A1(new_n24625_), .A2(new_n24508_), .ZN(new_n24626_));
  AOI21_X1   g22190(.A1(new_n24626_), .A2(new_n13251_), .B(pi0299), .ZN(new_n24627_));
  NOR2_X1    g22191(.A1(new_n24621_), .A2(new_n24627_), .ZN(new_n24628_));
  NOR3_X1    g22192(.A1(new_n13088_), .A2(new_n24611_), .A3(new_n12753_), .ZN(new_n24629_));
  NOR2_X1    g22193(.A1(new_n24629_), .A2(new_n24466_), .ZN(new_n24630_));
  NOR2_X1    g22194(.A1(new_n24630_), .A2(new_n5437_), .ZN(new_n24631_));
  NAND2_X1   g22195(.A1(new_n24629_), .A2(new_n13274_), .ZN(new_n24632_));
  INV_X1     g22196(.I(new_n24632_), .ZN(new_n24633_));
  NOR3_X1    g22197(.A1(new_n24631_), .A2(new_n24633_), .A3(new_n24465_), .ZN(new_n24634_));
  NOR2_X1    g22198(.A1(new_n24634_), .A2(new_n12751_), .ZN(new_n24635_));
  NOR3_X1    g22199(.A1(new_n24635_), .A2(new_n5403_), .A3(new_n24465_), .ZN(new_n24636_));
  NOR2_X1    g22200(.A1(new_n13088_), .A2(new_n24611_), .ZN(new_n24637_));
  AOI21_X1   g22201(.A1(new_n24637_), .A2(new_n12754_), .B(new_n24466_), .ZN(new_n24638_));
  NOR2_X1    g22202(.A1(new_n24539_), .A2(pi0603), .ZN(new_n24639_));
  INV_X1     g22203(.I(new_n24639_), .ZN(new_n24640_));
  NOR2_X1    g22204(.A1(new_n24635_), .A2(new_n13264_), .ZN(new_n24641_));
  AOI22_X1   g22205(.A1(new_n24641_), .A2(new_n24640_), .B1(new_n13264_), .B2(new_n24638_), .ZN(new_n24642_));
  NOR2_X1    g22206(.A1(new_n24642_), .A2(new_n5404_), .ZN(new_n24643_));
  NOR3_X1    g22207(.A1(new_n24643_), .A2(new_n5445_), .A3(new_n24636_), .ZN(new_n24644_));
  INV_X1     g22208(.I(new_n13276_), .ZN(new_n24645_));
  NOR2_X1    g22209(.A1(new_n24633_), .A2(new_n24515_), .ZN(new_n24646_));
  INV_X1     g22210(.I(new_n13215_), .ZN(new_n24647_));
  NOR2_X1    g22211(.A1(new_n24647_), .A2(new_n24611_), .ZN(new_n24648_));
  AOI21_X1   g22212(.A1(new_n24648_), .A2(new_n13213_), .B(new_n24469_), .ZN(new_n24649_));
  OAI22_X1   g22213(.A1(new_n24649_), .A2(new_n5404_), .B1(new_n24645_), .B2(new_n24646_), .ZN(new_n24650_));
  AND2_X2    g22214(.A1(new_n24650_), .A2(new_n5445_), .Z(new_n24651_));
  OAI21_X1   g22215(.A1(new_n24644_), .A2(new_n24651_), .B(pi0223), .ZN(new_n24652_));
  NOR2_X1    g22216(.A1(new_n24630_), .A2(new_n12751_), .ZN(new_n24653_));
  NAND2_X1   g22217(.A1(new_n24653_), .A2(new_n13096_), .ZN(new_n24654_));
  NAND2_X1   g22218(.A1(new_n24654_), .A2(new_n24640_), .ZN(new_n24655_));
  OAI21_X1   g22219(.A1(new_n24653_), .A2(new_n5406_), .B(new_n13095_), .ZN(new_n24656_));
  AOI21_X1   g22220(.A1(new_n13608_), .A2(pi0633), .B(new_n24546_), .ZN(new_n24657_));
  NOR2_X1    g22221(.A1(new_n24657_), .A2(new_n5398_), .ZN(new_n24658_));
  OAI21_X1   g22222(.A1(new_n24658_), .A2(new_n24631_), .B(pi0603), .ZN(new_n24659_));
  AOI21_X1   g22223(.A1(new_n24659_), .A2(new_n5406_), .B(new_n24656_), .ZN(new_n24660_));
  NOR2_X1    g22224(.A1(new_n24660_), .A2(new_n24655_), .ZN(new_n24661_));
  NAND3_X1   g22225(.A1(new_n13109_), .A2(pi0198), .A3(new_n12751_), .ZN(new_n24662_));
  AND3_X2    g22226(.A1(new_n24659_), .A2(new_n5404_), .A3(new_n24662_), .Z(new_n24663_));
  AOI21_X1   g22227(.A1(new_n24661_), .A2(new_n5403_), .B(new_n24663_), .ZN(new_n24664_));
  NOR2_X1    g22228(.A1(new_n24664_), .A2(new_n5445_), .ZN(new_n24665_));
  INV_X1     g22229(.I(new_n24657_), .ZN(new_n24666_));
  NAND2_X1   g22230(.A1(new_n24666_), .A2(pi0603), .ZN(new_n24667_));
  NAND2_X1   g22231(.A1(new_n13316_), .A2(new_n12751_), .ZN(new_n24668_));
  NAND2_X1   g22232(.A1(new_n24630_), .A2(new_n5437_), .ZN(new_n24669_));
  NAND3_X1   g22233(.A1(new_n24669_), .A2(pi0603), .A3(new_n13264_), .ZN(new_n24670_));
  NOR2_X1    g22234(.A1(new_n24666_), .A2(new_n5437_), .ZN(new_n24671_));
  OAI22_X1   g22235(.A1(new_n24671_), .A2(new_n24670_), .B1(new_n2672_), .B2(new_n24668_), .ZN(new_n24672_));
  NOR2_X1    g22236(.A1(new_n24667_), .A2(new_n13264_), .ZN(new_n24673_));
  NOR2_X1    g22237(.A1(new_n24672_), .A2(new_n24673_), .ZN(new_n24674_));
  NOR2_X1    g22238(.A1(new_n24546_), .A2(new_n5403_), .ZN(new_n24675_));
  AOI22_X1   g22239(.A1(new_n24674_), .A2(new_n5403_), .B1(new_n24667_), .B2(new_n24675_), .ZN(new_n24676_));
  NOR2_X1    g22240(.A1(new_n24676_), .A2(new_n5446_), .ZN(new_n24677_));
  OAI21_X1   g22241(.A1(new_n24677_), .A2(new_n24665_), .B(new_n2642_), .ZN(new_n24678_));
  AOI21_X1   g22242(.A1(new_n24638_), .A2(new_n2641_), .B(pi0223), .ZN(new_n24679_));
  NAND2_X1   g22243(.A1(new_n24678_), .A2(new_n24679_), .ZN(new_n24680_));
  AOI21_X1   g22244(.A1(new_n24680_), .A2(new_n24652_), .B(pi0299), .ZN(new_n24681_));
  OR3_X2     g22245(.A1(new_n24643_), .A2(new_n6764_), .A3(new_n24636_), .Z(new_n24682_));
  NAND2_X1   g22246(.A1(new_n24650_), .A2(new_n6764_), .ZN(new_n24683_));
  NAND2_X1   g22247(.A1(new_n24682_), .A2(new_n24683_), .ZN(new_n24684_));
  NOR2_X1    g22248(.A1(new_n24664_), .A2(new_n6764_), .ZN(new_n24685_));
  NOR2_X1    g22249(.A1(new_n24676_), .A2(new_n5422_), .ZN(new_n24686_));
  OAI21_X1   g22250(.A1(new_n24686_), .A2(new_n24685_), .B(new_n3304_), .ZN(new_n24687_));
  AOI21_X1   g22251(.A1(new_n24638_), .A2(new_n3303_), .B(pi0215), .ZN(new_n24688_));
  AOI22_X1   g22252(.A1(new_n24687_), .A2(new_n24688_), .B1(pi0215), .B2(new_n24684_), .ZN(new_n24689_));
  OAI21_X1   g22253(.A1(new_n24689_), .A2(new_n2628_), .B(pi0039), .ZN(new_n24690_));
  OAI22_X1   g22254(.A1(new_n24690_), .A2(new_n24681_), .B1(pi0039), .B2(new_n24628_), .ZN(new_n24691_));
  NAND2_X1   g22255(.A1(new_n24691_), .A2(new_n3265_), .ZN(new_n24692_));
  NAND3_X1   g22256(.A1(new_n24692_), .A2(new_n2609_), .A3(new_n24614_), .ZN(new_n24693_));
  OAI21_X1   g22257(.A1(new_n2672_), .A2(new_n2609_), .B(new_n24693_), .ZN(new_n24694_));
  NOR2_X1    g22258(.A1(new_n24694_), .A2(new_n12760_), .ZN(new_n24695_));
  AOI21_X1   g22259(.A1(new_n12760_), .A2(new_n24489_), .B(new_n24695_), .ZN(new_n24696_));
  NAND2_X1   g22260(.A1(new_n24489_), .A2(new_n13354_), .ZN(new_n24697_));
  OAI21_X1   g22261(.A1(new_n24694_), .A2(new_n13354_), .B(new_n24697_), .ZN(new_n24698_));
  NOR2_X1    g22262(.A1(new_n24698_), .A2(pi1155), .ZN(new_n24699_));
  NOR2_X1    g22263(.A1(new_n24694_), .A2(new_n13357_), .ZN(new_n24700_));
  AOI21_X1   g22264(.A1(new_n13357_), .A2(new_n24489_), .B(new_n24700_), .ZN(new_n24701_));
  NAND2_X1   g22265(.A1(new_n24701_), .A2(pi1155), .ZN(new_n24702_));
  NAND2_X1   g22266(.A1(new_n24702_), .A2(pi0785), .ZN(new_n24703_));
  OAI22_X1   g22267(.A1(new_n24703_), .A2(new_n24699_), .B1(pi0785), .B2(new_n24696_), .ZN(new_n24704_));
  NAND2_X1   g22268(.A1(new_n24704_), .A2(new_n12779_), .ZN(new_n24705_));
  NAND2_X1   g22269(.A1(new_n24581_), .A2(pi0618), .ZN(new_n24706_));
  OAI21_X1   g22270(.A1(new_n24704_), .A2(pi0618), .B(new_n24706_), .ZN(new_n24707_));
  NAND2_X1   g22271(.A1(new_n24707_), .A2(new_n12785_), .ZN(new_n24708_));
  NOR2_X1    g22272(.A1(new_n24704_), .A2(new_n12781_), .ZN(new_n24709_));
  NOR2_X1    g22273(.A1(new_n24489_), .A2(pi0618), .ZN(new_n24710_));
  NOR2_X1    g22274(.A1(new_n24709_), .A2(new_n24710_), .ZN(new_n24711_));
  NOR2_X1    g22275(.A1(new_n24711_), .A2(new_n12785_), .ZN(new_n24712_));
  NOR2_X1    g22276(.A1(new_n24712_), .A2(new_n12779_), .ZN(new_n24713_));
  NAND2_X1   g22277(.A1(new_n24713_), .A2(new_n24708_), .ZN(new_n24714_));
  NAND2_X1   g22278(.A1(new_n24714_), .A2(new_n24705_), .ZN(new_n24715_));
  NAND2_X1   g22279(.A1(new_n24715_), .A2(new_n12796_), .ZN(new_n24716_));
  NAND2_X1   g22280(.A1(new_n24581_), .A2(pi0619), .ZN(new_n24717_));
  OAI21_X1   g22281(.A1(new_n24715_), .A2(pi0619), .B(new_n24717_), .ZN(new_n24718_));
  NAND2_X1   g22282(.A1(new_n24718_), .A2(new_n12791_), .ZN(new_n24719_));
  NOR2_X1    g22283(.A1(new_n24715_), .A2(new_n12793_), .ZN(new_n24720_));
  NOR2_X1    g22284(.A1(new_n24489_), .A2(pi0619), .ZN(new_n24721_));
  NOR2_X1    g22285(.A1(new_n24720_), .A2(new_n24721_), .ZN(new_n24722_));
  NOR2_X1    g22286(.A1(new_n24722_), .A2(new_n12791_), .ZN(new_n24723_));
  NOR2_X1    g22287(.A1(new_n24723_), .A2(new_n12796_), .ZN(new_n24724_));
  NAND2_X1   g22288(.A1(new_n24724_), .A2(new_n24719_), .ZN(new_n24725_));
  NAND2_X1   g22289(.A1(new_n24725_), .A2(new_n24716_), .ZN(new_n24726_));
  NOR2_X1    g22290(.A1(new_n24489_), .A2(new_n17504_), .ZN(new_n24727_));
  INV_X1     g22291(.I(new_n24727_), .ZN(new_n24728_));
  OAI21_X1   g22292(.A1(new_n24726_), .A2(new_n12818_), .B(new_n24728_), .ZN(new_n24729_));
  NOR2_X1    g22293(.A1(new_n24581_), .A2(new_n13384_), .ZN(new_n24730_));
  INV_X1     g22294(.I(new_n24730_), .ZN(new_n24731_));
  OAI21_X1   g22295(.A1(new_n24729_), .A2(new_n12943_), .B(new_n24731_), .ZN(new_n24732_));
  NAND2_X1   g22296(.A1(new_n24489_), .A2(new_n12741_), .ZN(new_n24733_));
  OAI21_X1   g22297(.A1(new_n24606_), .A2(new_n12741_), .B(new_n24733_), .ZN(new_n24734_));
  OAI22_X1   g22298(.A1(new_n24732_), .A2(new_n17212_), .B1(new_n15576_), .B2(new_n24734_), .ZN(new_n24735_));
  NOR2_X1    g22299(.A1(new_n24735_), .A2(new_n24610_), .ZN(new_n24736_));
  NAND2_X1   g22300(.A1(new_n24601_), .A2(pi0629), .ZN(new_n24737_));
  NAND2_X1   g22301(.A1(new_n24729_), .A2(new_n19160_), .ZN(new_n24738_));
  NAND2_X1   g22302(.A1(new_n24738_), .A2(new_n24737_), .ZN(new_n24739_));
  NOR2_X1    g22303(.A1(new_n24603_), .A2(new_n18087_), .ZN(new_n24740_));
  NOR2_X1    g22304(.A1(new_n24739_), .A2(new_n24740_), .ZN(new_n24741_));
  NAND2_X1   g22305(.A1(new_n24741_), .A2(new_n15340_), .ZN(new_n24742_));
  NAND2_X1   g22306(.A1(new_n24742_), .A2(new_n15693_), .ZN(new_n24743_));
  NOR2_X1    g22307(.A1(new_n24741_), .A2(new_n12937_), .ZN(new_n24744_));
  INV_X1     g22308(.I(new_n24613_), .ZN(new_n24745_));
  NOR2_X1    g22309(.A1(new_n13572_), .A2(new_n24493_), .ZN(new_n24746_));
  AOI21_X1   g22310(.A1(new_n13136_), .A2(new_n24746_), .B(new_n24745_), .ZN(new_n24747_));
  OAI21_X1   g22311(.A1(new_n24747_), .A2(new_n24491_), .B(pi0038), .ZN(new_n24748_));
  INV_X1     g22312(.I(new_n24748_), .ZN(new_n24749_));
  NOR4_X1    g22313(.A1(new_n13088_), .A2(new_n24493_), .A3(pi0665), .A4(new_n13290_), .ZN(new_n24750_));
  NOR3_X1    g22314(.A1(new_n24750_), .A2(new_n24629_), .A3(new_n24466_), .ZN(new_n24751_));
  OR2_X2     g22315(.A1(new_n24751_), .A2(new_n5437_), .Z(new_n24752_));
  NOR3_X1    g22316(.A1(new_n13261_), .A2(pi0198), .A3(pi0665), .ZN(new_n24753_));
  NOR3_X1    g22317(.A1(new_n13290_), .A2(new_n2672_), .A3(pi0665), .ZN(new_n24754_));
  OAI21_X1   g22318(.A1(new_n24753_), .A2(new_n24754_), .B(pi0634), .ZN(new_n24755_));
  NAND2_X1   g22319(.A1(new_n24646_), .A2(new_n24755_), .ZN(new_n24756_));
  NAND2_X1   g22320(.A1(new_n24756_), .A2(new_n5437_), .ZN(new_n24757_));
  NAND2_X1   g22321(.A1(new_n24757_), .A2(new_n24752_), .ZN(new_n24758_));
  NAND2_X1   g22322(.A1(new_n24758_), .A2(pi0603), .ZN(new_n24759_));
  OR2_X2     g22323(.A1(new_n24531_), .A2(pi0603), .Z(new_n24760_));
  AOI21_X1   g22324(.A1(new_n24759_), .A2(new_n24760_), .B(new_n5403_), .ZN(new_n24761_));
  INV_X1     g22325(.I(new_n24642_), .ZN(new_n24762_));
  NOR2_X1    g22326(.A1(new_n24751_), .A2(new_n12751_), .ZN(new_n24763_));
  INV_X1     g22327(.I(new_n24763_), .ZN(new_n24764_));
  NAND2_X1   g22328(.A1(new_n24532_), .A2(new_n12751_), .ZN(new_n24765_));
  NAND2_X1   g22329(.A1(new_n24764_), .A2(new_n24765_), .ZN(new_n24766_));
  OAI21_X1   g22330(.A1(new_n24766_), .A2(new_n5408_), .B(new_n13584_), .ZN(new_n24767_));
  AND3_X2    g22331(.A1(new_n24759_), .A2(new_n5408_), .A3(new_n24765_), .Z(new_n24768_));
  OAI22_X1   g22332(.A1(new_n24768_), .A2(new_n24767_), .B1(pi0680), .B2(new_n24762_), .ZN(new_n24769_));
  NOR2_X1    g22333(.A1(new_n24769_), .A2(new_n24761_), .ZN(new_n24770_));
  NOR2_X1    g22334(.A1(new_n24770_), .A2(new_n6764_), .ZN(new_n24771_));
  INV_X1     g22335(.I(new_n24670_), .ZN(new_n24772_));
  AOI21_X1   g22336(.A1(new_n13264_), .A2(new_n24763_), .B(new_n24772_), .ZN(new_n24773_));
  NAND2_X1   g22337(.A1(new_n24773_), .A2(new_n5409_), .ZN(new_n24774_));
  NAND2_X1   g22338(.A1(new_n24774_), .A2(new_n24756_), .ZN(new_n24775_));
  NOR2_X1    g22339(.A1(new_n24773_), .A2(new_n5398_), .ZN(new_n24776_));
  NOR2_X1    g22340(.A1(new_n24523_), .A2(pi0603), .ZN(new_n24777_));
  NOR2_X1    g22341(.A1(new_n24776_), .A2(new_n24777_), .ZN(new_n24778_));
  NAND2_X1   g22342(.A1(new_n24778_), .A2(new_n24775_), .ZN(new_n24779_));
  NOR2_X1    g22343(.A1(new_n24517_), .A2(pi0603), .ZN(new_n24780_));
  AOI21_X1   g22344(.A1(new_n24756_), .A2(pi0603), .B(new_n24780_), .ZN(new_n24781_));
  OAI22_X1   g22345(.A1(new_n24649_), .A2(pi0680), .B1(new_n24781_), .B2(new_n5403_), .ZN(new_n24782_));
  AOI21_X1   g22346(.A1(new_n24779_), .A2(new_n13584_), .B(new_n24782_), .ZN(new_n24783_));
  NOR2_X1    g22347(.A1(new_n24783_), .A2(new_n5422_), .ZN(new_n24784_));
  OAI21_X1   g22348(.A1(new_n24771_), .A2(new_n24784_), .B(pi0215), .ZN(new_n24785_));
  OAI21_X1   g22349(.A1(new_n24493_), .A2(new_n14710_), .B(new_n24657_), .ZN(new_n24786_));
  NAND2_X1   g22350(.A1(new_n24786_), .A2(new_n5437_), .ZN(new_n24787_));
  AOI21_X1   g22351(.A1(new_n24787_), .A2(new_n24752_), .B(new_n12751_), .ZN(new_n24788_));
  NOR2_X1    g22352(.A1(new_n24549_), .A2(pi0603), .ZN(new_n24789_));
  OR3_X2     g22353(.A1(new_n24788_), .A2(new_n13119_), .A3(new_n24789_), .Z(new_n24790_));
  NAND2_X1   g22354(.A1(new_n24764_), .A2(pi0642), .ZN(new_n24791_));
  OAI21_X1   g22355(.A1(new_n24788_), .A2(pi0642), .B(new_n24791_), .ZN(new_n24792_));
  NAND3_X1   g22356(.A1(new_n24792_), .A2(new_n13095_), .A3(new_n24765_), .ZN(new_n24793_));
  OAI21_X1   g22357(.A1(new_n13095_), .A2(new_n24766_), .B(new_n24793_), .ZN(new_n24794_));
  AOI21_X1   g22358(.A1(new_n24794_), .A2(new_n13119_), .B(new_n12821_), .ZN(new_n24795_));
  NOR2_X1    g22359(.A1(new_n24661_), .A2(pi0680), .ZN(new_n24796_));
  AOI21_X1   g22360(.A1(new_n24795_), .A2(new_n24790_), .B(new_n24796_), .ZN(new_n24797_));
  AOI22_X1   g22361(.A1(new_n24548_), .A2(new_n12755_), .B1(new_n24666_), .B2(pi0603), .ZN(new_n24798_));
  AOI21_X1   g22362(.A1(new_n24774_), .A2(new_n24786_), .B(new_n24776_), .ZN(new_n24799_));
  NAND2_X1   g22363(.A1(new_n24558_), .A2(new_n12751_), .ZN(new_n24800_));
  AOI21_X1   g22364(.A1(new_n24799_), .A2(new_n24800_), .B(new_n13585_), .ZN(new_n24801_));
  NOR2_X1    g22365(.A1(new_n24674_), .A2(pi0680), .ZN(new_n24802_));
  NOR2_X1    g22366(.A1(new_n24801_), .A2(new_n24802_), .ZN(new_n24803_));
  OAI21_X1   g22367(.A1(new_n5403_), .A2(new_n24798_), .B(new_n24803_), .ZN(new_n24804_));
  NOR2_X1    g22368(.A1(new_n24804_), .A2(new_n5422_), .ZN(new_n24805_));
  AOI21_X1   g22369(.A1(new_n24797_), .A2(new_n5422_), .B(new_n24805_), .ZN(new_n24806_));
  INV_X1     g22370(.I(new_n24638_), .ZN(new_n24807_));
  AOI21_X1   g22371(.A1(new_n13421_), .A2(new_n24746_), .B(new_n24807_), .ZN(new_n24808_));
  AOI21_X1   g22372(.A1(new_n24808_), .A2(new_n3303_), .B(pi0215), .ZN(new_n24809_));
  OAI21_X1   g22373(.A1(new_n24806_), .A2(new_n3303_), .B(new_n24809_), .ZN(new_n24810_));
  AOI21_X1   g22374(.A1(new_n24810_), .A2(new_n24785_), .B(new_n2628_), .ZN(new_n24811_));
  NOR2_X1    g22375(.A1(new_n24804_), .A2(new_n5446_), .ZN(new_n24812_));
  AOI21_X1   g22376(.A1(new_n24797_), .A2(new_n5446_), .B(new_n24812_), .ZN(new_n24813_));
  AOI21_X1   g22377(.A1(new_n24808_), .A2(new_n2641_), .B(pi0223), .ZN(new_n24814_));
  OAI21_X1   g22378(.A1(new_n24813_), .A2(new_n2641_), .B(new_n24814_), .ZN(new_n24815_));
  NOR2_X1    g22379(.A1(new_n24770_), .A2(new_n5445_), .ZN(new_n24816_));
  NOR2_X1    g22380(.A1(new_n24783_), .A2(new_n5446_), .ZN(new_n24817_));
  OAI21_X1   g22381(.A1(new_n24816_), .A2(new_n24817_), .B(pi0223), .ZN(new_n24818_));
  AOI21_X1   g22382(.A1(new_n24815_), .A2(new_n24818_), .B(pi0299), .ZN(new_n24819_));
  OR3_X2     g22383(.A1(new_n24811_), .A2(new_n24819_), .A3(new_n2627_), .Z(new_n24820_));
  OAI21_X1   g22384(.A1(new_n24512_), .A2(pi0603), .B(pi0680), .ZN(new_n24821_));
  NOR2_X1    g22385(.A1(new_n13038_), .A2(new_n12752_), .ZN(new_n24822_));
  NOR2_X1    g22386(.A1(new_n24822_), .A2(pi0198), .ZN(new_n24823_));
  NAND2_X1   g22387(.A1(new_n24611_), .A2(pi0198), .ZN(new_n24824_));
  NAND3_X1   g22388(.A1(new_n24824_), .A2(pi0634), .A3(new_n12822_), .ZN(new_n24825_));
  OAI21_X1   g22389(.A1(new_n24823_), .A2(new_n24825_), .B(pi0603), .ZN(new_n24826_));
  AOI21_X1   g22390(.A1(new_n24624_), .A2(pi0633), .B(new_n24826_), .ZN(new_n24827_));
  NOR2_X1    g22391(.A1(new_n24508_), .A2(pi0634), .ZN(new_n24828_));
  NOR4_X1    g22392(.A1(new_n13198_), .A2(new_n24511_), .A3(new_n2672_), .A4(new_n24493_), .ZN(new_n24829_));
  OAI21_X1   g22393(.A1(new_n24829_), .A2(new_n24828_), .B(new_n24611_), .ZN(new_n24830_));
  AOI21_X1   g22394(.A1(new_n24827_), .A2(new_n24830_), .B(new_n24821_), .ZN(new_n24831_));
  AND3_X2    g22395(.A1(new_n24626_), .A2(new_n12821_), .A3(new_n13251_), .Z(new_n24832_));
  NOR3_X1    g22396(.A1(new_n24831_), .A2(new_n24832_), .A3(pi0299), .ZN(new_n24833_));
  INV_X1     g22397(.I(new_n24833_), .ZN(new_n24834_));
  AOI21_X1   g22398(.A1(new_n24620_), .A2(new_n24499_), .B(new_n2628_), .ZN(new_n24835_));
  AOI21_X1   g22399(.A1(pi0198), .A2(pi0665), .B(new_n24502_), .ZN(new_n24836_));
  NOR3_X1    g22400(.A1(new_n24836_), .A2(new_n24616_), .A3(new_n24611_), .ZN(new_n24837_));
  INV_X1     g22401(.I(new_n24837_), .ZN(new_n24838_));
  NOR2_X1    g22402(.A1(pi0198), .A2(pi0665), .ZN(new_n24839_));
  AOI21_X1   g22403(.A1(new_n14558_), .A2(new_n24839_), .B(pi0633), .ZN(new_n24840_));
  INV_X1     g22404(.I(new_n13201_), .ZN(new_n24841_));
  NOR3_X1    g22405(.A1(new_n24841_), .A2(new_n24501_), .A3(new_n2672_), .ZN(new_n24842_));
  INV_X1     g22406(.I(new_n24842_), .ZN(new_n24843_));
  AOI21_X1   g22407(.A1(new_n24843_), .A2(new_n24840_), .B(new_n12751_), .ZN(new_n24844_));
  AOI22_X1   g22408(.A1(new_n24838_), .A2(new_n24844_), .B1(new_n12751_), .B2(new_n24503_), .ZN(new_n24845_));
  OAI21_X1   g22409(.A1(new_n24845_), .A2(new_n24499_), .B(new_n24835_), .ZN(new_n24846_));
  AOI21_X1   g22410(.A1(new_n24846_), .A2(new_n24834_), .B(pi0039), .ZN(new_n24847_));
  INV_X1     g22411(.I(new_n24847_), .ZN(new_n24848_));
  AOI21_X1   g22412(.A1(new_n24820_), .A2(new_n24848_), .B(pi0038), .ZN(new_n24849_));
  NOR3_X1    g22413(.A1(new_n24849_), .A2(new_n2610_), .A3(new_n24749_), .ZN(new_n24850_));
  NOR2_X1    g22414(.A1(new_n24850_), .A2(new_n24490_), .ZN(new_n24851_));
  NOR2_X1    g22415(.A1(new_n24851_), .A2(pi0778), .ZN(new_n24852_));
  OAI21_X1   g22416(.A1(new_n24850_), .A2(new_n24490_), .B(new_n13521_), .ZN(new_n24853_));
  NAND2_X1   g22417(.A1(new_n24694_), .A2(pi0625), .ZN(new_n24854_));
  AOI21_X1   g22418(.A1(new_n24853_), .A2(new_n24854_), .B(pi1153), .ZN(new_n24855_));
  NOR3_X1    g22419(.A1(new_n24855_), .A2(pi0608), .A3(new_n24587_), .ZN(new_n24856_));
  NAND2_X1   g22420(.A1(new_n24694_), .A2(new_n13521_), .ZN(new_n24857_));
  OAI21_X1   g22421(.A1(new_n24851_), .A2(new_n13521_), .B(new_n24857_), .ZN(new_n24858_));
  NAND2_X1   g22422(.A1(new_n24584_), .A2(pi0608), .ZN(new_n24859_));
  AOI21_X1   g22423(.A1(new_n24858_), .A2(pi1153), .B(new_n24859_), .ZN(new_n24860_));
  NOR3_X1    g22424(.A1(new_n24856_), .A2(new_n24860_), .A3(new_n12758_), .ZN(new_n24861_));
  NOR2_X1    g22425(.A1(new_n24861_), .A2(new_n24852_), .ZN(new_n24862_));
  NOR2_X1    g22426(.A1(new_n24862_), .A2(pi0785), .ZN(new_n24863_));
  NOR2_X1    g22427(.A1(new_n24699_), .A2(new_n13829_), .ZN(new_n24864_));
  NAND2_X1   g22428(.A1(new_n24590_), .A2(new_n12766_), .ZN(new_n24865_));
  NAND2_X1   g22429(.A1(new_n24865_), .A2(pi1155), .ZN(new_n24866_));
  NOR3_X1    g22430(.A1(new_n24861_), .A2(new_n12766_), .A3(new_n24852_), .ZN(new_n24867_));
  OAI21_X1   g22431(.A1(new_n24866_), .A2(new_n24867_), .B(new_n24864_), .ZN(new_n24868_));
  AOI21_X1   g22432(.A1(new_n24590_), .A2(pi0609), .B(pi1155), .ZN(new_n24869_));
  NAND2_X1   g22433(.A1(new_n24862_), .A2(new_n12766_), .ZN(new_n24870_));
  NAND2_X1   g22434(.A1(new_n24870_), .A2(new_n24869_), .ZN(new_n24871_));
  NAND3_X1   g22435(.A1(new_n24871_), .A2(new_n13829_), .A3(new_n24702_), .ZN(new_n24872_));
  AND3_X2    g22436(.A1(new_n24872_), .A2(new_n24868_), .A3(pi0785), .Z(new_n24873_));
  NOR2_X1    g22437(.A1(new_n24873_), .A2(new_n24863_), .ZN(new_n24874_));
  NOR2_X1    g22438(.A1(new_n24874_), .A2(pi0781), .ZN(new_n24875_));
  NAND2_X1   g22439(.A1(new_n24708_), .A2(pi0627), .ZN(new_n24876_));
  OAI21_X1   g22440(.A1(new_n24593_), .A2(pi0618), .B(pi1154), .ZN(new_n24877_));
  AOI21_X1   g22441(.A1(new_n24874_), .A2(pi0618), .B(new_n24877_), .ZN(new_n24878_));
  NOR2_X1    g22442(.A1(new_n24878_), .A2(new_n24876_), .ZN(new_n24879_));
  OAI21_X1   g22443(.A1(new_n24593_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n24880_));
  NOR3_X1    g22444(.A1(new_n24873_), .A2(pi0618), .A3(new_n24863_), .ZN(new_n24881_));
  NOR2_X1    g22445(.A1(new_n24881_), .A2(new_n24880_), .ZN(new_n24882_));
  NOR3_X1    g22446(.A1(new_n24882_), .A2(pi0627), .A3(new_n24712_), .ZN(new_n24883_));
  NOR3_X1    g22447(.A1(new_n24883_), .A2(new_n24879_), .A3(new_n12779_), .ZN(new_n24884_));
  NOR2_X1    g22448(.A1(new_n24884_), .A2(new_n24875_), .ZN(new_n24885_));
  NOR2_X1    g22449(.A1(new_n24885_), .A2(pi0789), .ZN(new_n24886_));
  NOR2_X1    g22450(.A1(new_n24886_), .A2(new_n14303_), .ZN(new_n24887_));
  NAND2_X1   g22451(.A1(new_n24719_), .A2(pi0648), .ZN(new_n24888_));
  NOR2_X1    g22452(.A1(new_n24595_), .A2(pi0619), .ZN(new_n24889_));
  NOR2_X1    g22453(.A1(new_n24889_), .A2(new_n12791_), .ZN(new_n24890_));
  NAND2_X1   g22454(.A1(new_n24885_), .A2(pi0619), .ZN(new_n24891_));
  AOI21_X1   g22455(.A1(new_n24891_), .A2(new_n24890_), .B(new_n24888_), .ZN(new_n24892_));
  OAI21_X1   g22456(.A1(new_n24722_), .A2(new_n12791_), .B(new_n12895_), .ZN(new_n24893_));
  OAI21_X1   g22457(.A1(new_n24595_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n24894_));
  AOI21_X1   g22458(.A1(new_n24885_), .A2(new_n12793_), .B(new_n24894_), .ZN(new_n24895_));
  OAI21_X1   g22459(.A1(new_n24895_), .A2(new_n24893_), .B(pi0789), .ZN(new_n24896_));
  OAI21_X1   g22460(.A1(new_n24896_), .A2(new_n24892_), .B(new_n24887_), .ZN(new_n24897_));
  NAND2_X1   g22461(.A1(new_n24726_), .A2(pi0626), .ZN(new_n24898_));
  NAND2_X1   g22462(.A1(new_n24489_), .A2(new_n12747_), .ZN(new_n24899_));
  AOI21_X1   g22463(.A1(new_n24898_), .A2(new_n24899_), .B(new_n12813_), .ZN(new_n24900_));
  NOR2_X1    g22464(.A1(new_n24595_), .A2(new_n12910_), .ZN(new_n24901_));
  AOI21_X1   g22465(.A1(new_n12910_), .A2(new_n24489_), .B(new_n24901_), .ZN(new_n24902_));
  NOR2_X1    g22466(.A1(new_n24581_), .A2(new_n12747_), .ZN(new_n24903_));
  AOI21_X1   g22467(.A1(new_n24726_), .A2(new_n12747_), .B(new_n24903_), .ZN(new_n24904_));
  OAI22_X1   g22468(.A1(new_n24904_), .A2(new_n12816_), .B1(new_n12906_), .B2(new_n24902_), .ZN(new_n24905_));
  OAI21_X1   g22469(.A1(new_n24905_), .A2(new_n24900_), .B(pi0788), .ZN(new_n24906_));
  AOI21_X1   g22470(.A1(new_n24897_), .A2(new_n24906_), .B(new_n24744_), .ZN(new_n24907_));
  OAI22_X1   g22471(.A1(new_n24907_), .A2(new_n24743_), .B1(new_n12972_), .B2(new_n24736_), .ZN(new_n24908_));
  NAND2_X1   g22472(.A1(new_n24581_), .A2(pi0644), .ZN(new_n24909_));
  NOR2_X1    g22473(.A1(new_n24732_), .A2(new_n12984_), .ZN(new_n24910_));
  AOI21_X1   g22474(.A1(new_n12984_), .A2(new_n24581_), .B(new_n24910_), .ZN(new_n24911_));
  OAI21_X1   g22475(.A1(new_n24911_), .A2(pi0644), .B(new_n24909_), .ZN(new_n24912_));
  AOI21_X1   g22476(.A1(new_n24912_), .A2(pi0715), .B(pi1160), .ZN(new_n24913_));
  OR2_X2     g22477(.A1(new_n24734_), .A2(new_n12965_), .Z(new_n24914_));
  NAND3_X1   g22478(.A1(new_n24609_), .A2(pi0787), .A3(new_n24914_), .ZN(new_n24915_));
  OAI21_X1   g22479(.A1(pi0787), .A2(new_n24606_), .B(new_n24915_), .ZN(new_n24916_));
  NAND2_X1   g22480(.A1(new_n24916_), .A2(pi0644), .ZN(new_n24917_));
  NAND2_X1   g22481(.A1(new_n24917_), .A2(new_n12740_), .ZN(new_n24918_));
  NOR2_X1    g22482(.A1(new_n24908_), .A2(pi0644), .ZN(new_n24919_));
  OAI21_X1   g22483(.A1(new_n24919_), .A2(new_n24918_), .B(new_n24913_), .ZN(new_n24920_));
  NAND2_X1   g22484(.A1(new_n24581_), .A2(new_n12975_), .ZN(new_n24921_));
  OAI21_X1   g22485(.A1(new_n24911_), .A2(new_n12975_), .B(new_n24921_), .ZN(new_n24922_));
  AOI21_X1   g22486(.A1(new_n24922_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n24923_));
  AOI21_X1   g22487(.A1(new_n24916_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n24924_));
  OAI21_X1   g22488(.A1(new_n24908_), .A2(new_n12975_), .B(new_n24924_), .ZN(new_n24925_));
  AOI21_X1   g22489(.A1(new_n24925_), .A2(new_n24923_), .B(new_n13000_), .ZN(new_n24926_));
  AOI22_X1   g22490(.A1(new_n24926_), .A2(new_n24920_), .B1(new_n13000_), .B2(new_n24908_), .ZN(new_n24927_));
  NAND2_X1   g22491(.A1(po1038), .A2(pi0198), .ZN(new_n24928_));
  OAI21_X1   g22492(.A1(new_n24927_), .A2(po1038), .B(new_n24928_), .ZN(po0355));
  NOR2_X1    g22493(.A1(new_n2609_), .A2(pi0199), .ZN(new_n24930_));
  INV_X1     g22494(.I(new_n13398_), .ZN(new_n24931_));
  NAND2_X1   g22495(.A1(new_n13397_), .A2(pi0199), .ZN(new_n24932_));
  AOI21_X1   g22496(.A1(new_n24931_), .A2(new_n24932_), .B(new_n3265_), .ZN(new_n24933_));
  NAND2_X1   g22497(.A1(new_n13416_), .A2(new_n8525_), .ZN(new_n24934_));
  NAND2_X1   g22498(.A1(new_n13406_), .A2(pi0199), .ZN(new_n24935_));
  AOI21_X1   g22499(.A1(new_n24935_), .A2(new_n24934_), .B(pi0039), .ZN(new_n24936_));
  NAND2_X1   g22500(.A1(new_n15743_), .A2(pi0199), .ZN(new_n24937_));
  NAND3_X1   g22501(.A1(new_n13442_), .A2(new_n13452_), .A3(new_n8525_), .ZN(new_n24938_));
  AOI21_X1   g22502(.A1(new_n24937_), .A2(new_n24938_), .B(new_n2627_), .ZN(new_n24939_));
  NOR3_X1    g22503(.A1(new_n24939_), .A2(pi0038), .A3(new_n24936_), .ZN(new_n24940_));
  NOR3_X1    g22504(.A1(new_n24940_), .A2(new_n2610_), .A3(new_n24933_), .ZN(new_n24941_));
  OAI21_X1   g22505(.A1(new_n24941_), .A2(new_n24930_), .B(pi0637), .ZN(new_n24942_));
  INV_X1     g22506(.I(pi0637), .ZN(new_n24943_));
  NOR2_X1    g22507(.A1(new_n13193_), .A2(new_n8525_), .ZN(new_n24944_));
  INV_X1     g22508(.I(new_n24944_), .ZN(new_n24945_));
  NAND2_X1   g22509(.A1(new_n24945_), .A2(new_n24943_), .ZN(new_n24946_));
  NAND2_X1   g22510(.A1(new_n24942_), .A2(new_n24946_), .ZN(new_n24947_));
  INV_X1     g22511(.I(new_n24947_), .ZN(new_n24948_));
  OAI21_X1   g22512(.A1(new_n24944_), .A2(pi0625), .B(pi1153), .ZN(new_n24949_));
  AOI21_X1   g22513(.A1(new_n24947_), .A2(pi0625), .B(new_n24949_), .ZN(new_n24950_));
  OAI21_X1   g22514(.A1(new_n24944_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n24951_));
  AOI21_X1   g22515(.A1(new_n24942_), .A2(new_n24946_), .B(pi0625), .ZN(new_n24952_));
  OAI21_X1   g22516(.A1(new_n24952_), .A2(new_n24951_), .B(pi0778), .ZN(new_n24953_));
  OAI22_X1   g22517(.A1(new_n24953_), .A2(new_n24950_), .B1(pi0778), .B2(new_n24948_), .ZN(new_n24954_));
  NAND2_X1   g22518(.A1(new_n24944_), .A2(new_n12869_), .ZN(new_n24955_));
  OAI21_X1   g22519(.A1(new_n24954_), .A2(new_n12869_), .B(new_n24955_), .ZN(new_n24956_));
  INV_X1     g22520(.I(new_n24956_), .ZN(new_n24957_));
  NOR2_X1    g22521(.A1(new_n24944_), .A2(new_n12888_), .ZN(new_n24958_));
  AOI21_X1   g22522(.A1(new_n24957_), .A2(new_n12888_), .B(new_n24958_), .ZN(new_n24959_));
  NOR2_X1    g22523(.A1(new_n24945_), .A2(new_n12911_), .ZN(new_n24960_));
  AOI21_X1   g22524(.A1(new_n24959_), .A2(new_n12911_), .B(new_n24960_), .ZN(new_n24961_));
  INV_X1     g22525(.I(new_n24961_), .ZN(new_n24962_));
  NAND2_X1   g22526(.A1(new_n24945_), .A2(new_n12817_), .ZN(new_n24963_));
  OAI21_X1   g22527(.A1(new_n24962_), .A2(new_n12817_), .B(new_n24963_), .ZN(new_n24964_));
  NAND2_X1   g22528(.A1(new_n24944_), .A2(pi0628), .ZN(new_n24965_));
  OAI21_X1   g22529(.A1(new_n24964_), .A2(pi0628), .B(new_n24965_), .ZN(new_n24966_));
  AOI21_X1   g22530(.A1(new_n24966_), .A2(new_n12742_), .B(new_n12919_), .ZN(new_n24967_));
  NAND2_X1   g22531(.A1(new_n24945_), .A2(new_n12818_), .ZN(new_n24968_));
  NAND2_X1   g22532(.A1(new_n24944_), .A2(pi0609), .ZN(new_n24969_));
  INV_X1     g22533(.I(pi0617), .ZN(new_n24970_));
  INV_X1     g22534(.I(new_n24930_), .ZN(new_n24971_));
  NOR2_X1    g22535(.A1(new_n17986_), .A2(new_n8525_), .ZN(new_n24972_));
  NOR2_X1    g22536(.A1(new_n15784_), .A2(pi0199), .ZN(new_n24973_));
  OAI21_X1   g22537(.A1(new_n24972_), .A2(new_n24973_), .B(new_n3265_), .ZN(new_n24974_));
  OAI21_X1   g22538(.A1(new_n15006_), .A2(pi0199), .B(new_n15011_), .ZN(new_n24975_));
  NAND3_X1   g22539(.A1(new_n24974_), .A2(new_n2609_), .A3(new_n24975_), .ZN(new_n24976_));
  AOI21_X1   g22540(.A1(new_n24976_), .A2(new_n24971_), .B(new_n24970_), .ZN(new_n24977_));
  NOR2_X1    g22541(.A1(new_n24944_), .A2(pi0617), .ZN(new_n24978_));
  NOR2_X1    g22542(.A1(new_n24977_), .A2(new_n24978_), .ZN(new_n24979_));
  NAND2_X1   g22543(.A1(new_n24979_), .A2(new_n12761_), .ZN(new_n24980_));
  OAI21_X1   g22544(.A1(new_n12761_), .A2(new_n24945_), .B(new_n24980_), .ZN(new_n24981_));
  NAND2_X1   g22545(.A1(new_n24981_), .A2(new_n12766_), .ZN(new_n24982_));
  AOI21_X1   g22546(.A1(new_n24982_), .A2(new_n24969_), .B(pi1155), .ZN(new_n24983_));
  NAND2_X1   g22547(.A1(new_n24981_), .A2(pi0609), .ZN(new_n24984_));
  NAND2_X1   g22548(.A1(new_n24944_), .A2(new_n12766_), .ZN(new_n24985_));
  AOI21_X1   g22549(.A1(new_n24984_), .A2(new_n24985_), .B(new_n12770_), .ZN(new_n24986_));
  NOR3_X1    g22550(.A1(new_n24983_), .A2(new_n24986_), .A3(new_n12764_), .ZN(new_n24987_));
  NOR2_X1    g22551(.A1(new_n24981_), .A2(pi0785), .ZN(new_n24988_));
  NOR2_X1    g22552(.A1(new_n24987_), .A2(new_n24988_), .ZN(new_n24989_));
  NOR2_X1    g22553(.A1(new_n24945_), .A2(new_n12781_), .ZN(new_n24990_));
  AOI21_X1   g22554(.A1(new_n24989_), .A2(new_n12781_), .B(new_n24990_), .ZN(new_n24991_));
  NOR2_X1    g22555(.A1(new_n24991_), .A2(pi1154), .ZN(new_n24992_));
  NOR2_X1    g22556(.A1(new_n24945_), .A2(pi0618), .ZN(new_n24993_));
  AOI21_X1   g22557(.A1(new_n24989_), .A2(pi0618), .B(new_n24993_), .ZN(new_n24994_));
  OAI21_X1   g22558(.A1(new_n24994_), .A2(new_n12785_), .B(pi0781), .ZN(new_n24995_));
  OAI22_X1   g22559(.A1(new_n24995_), .A2(new_n24992_), .B1(pi0781), .B2(new_n24989_), .ZN(new_n24996_));
  NAND2_X1   g22560(.A1(new_n24944_), .A2(pi0619), .ZN(new_n24997_));
  OAI21_X1   g22561(.A1(new_n24996_), .A2(pi0619), .B(new_n24997_), .ZN(new_n24998_));
  NAND2_X1   g22562(.A1(new_n24998_), .A2(new_n12791_), .ZN(new_n24999_));
  NOR2_X1    g22563(.A1(new_n24945_), .A2(pi0619), .ZN(new_n25000_));
  INV_X1     g22564(.I(new_n25000_), .ZN(new_n25001_));
  OAI21_X1   g22565(.A1(new_n24996_), .A2(new_n12793_), .B(new_n25001_), .ZN(new_n25002_));
  AOI21_X1   g22566(.A1(new_n25002_), .A2(pi1159), .B(new_n12796_), .ZN(new_n25003_));
  AOI22_X1   g22567(.A1(new_n25003_), .A2(new_n24999_), .B1(new_n12796_), .B2(new_n24996_), .ZN(new_n25004_));
  OAI21_X1   g22568(.A1(new_n25004_), .A2(new_n12818_), .B(new_n24968_), .ZN(new_n25005_));
  AOI21_X1   g22569(.A1(new_n25005_), .A2(new_n12920_), .B(new_n12742_), .ZN(new_n25006_));
  AOI21_X1   g22570(.A1(new_n24944_), .A2(new_n12747_), .B(pi0641), .ZN(new_n25007_));
  NAND2_X1   g22571(.A1(new_n25004_), .A2(pi0626), .ZN(new_n25008_));
  AOI21_X1   g22572(.A1(new_n25008_), .A2(new_n25007_), .B(new_n12745_), .ZN(new_n25009_));
  AOI21_X1   g22573(.A1(new_n24962_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n25010_));
  OAI21_X1   g22574(.A1(new_n24977_), .A2(new_n24978_), .B(new_n24943_), .ZN(new_n25011_));
  AOI21_X1   g22575(.A1(new_n15111_), .A2(pi0199), .B(new_n24970_), .ZN(new_n25012_));
  NOR2_X1    g22576(.A1(new_n18438_), .A2(new_n2610_), .ZN(new_n25013_));
  OAI22_X1   g22577(.A1(new_n25013_), .A2(pi0199), .B1(new_n2610_), .B2(new_n25012_), .ZN(new_n25014_));
  NAND2_X1   g22578(.A1(new_n15124_), .A2(pi0038), .ZN(new_n25015_));
  OAI21_X1   g22579(.A1(new_n21986_), .A2(new_n15123_), .B(new_n2609_), .ZN(new_n25016_));
  NAND2_X1   g22580(.A1(new_n25016_), .A2(new_n8525_), .ZN(new_n25017_));
  NAND2_X1   g22581(.A1(new_n15128_), .A2(new_n15127_), .ZN(new_n25018_));
  NAND3_X1   g22582(.A1(new_n25018_), .A2(new_n3265_), .A3(pi0199), .ZN(new_n25019_));
  NAND4_X1   g22583(.A1(new_n25017_), .A2(new_n24970_), .A3(new_n25015_), .A4(new_n25019_), .ZN(new_n25020_));
  NAND3_X1   g22584(.A1(new_n25020_), .A2(pi0637), .A3(new_n25014_), .ZN(new_n25021_));
  NAND2_X1   g22585(.A1(new_n25011_), .A2(new_n25021_), .ZN(new_n25022_));
  NOR2_X1    g22586(.A1(new_n24952_), .A2(new_n24951_), .ZN(new_n25023_));
  OAI21_X1   g22587(.A1(new_n24979_), .A2(pi0625), .B(pi1153), .ZN(new_n25024_));
  AOI21_X1   g22588(.A1(new_n25022_), .A2(pi0625), .B(new_n25024_), .ZN(new_n25025_));
  NOR3_X1    g22589(.A1(new_n25025_), .A2(new_n13560_), .A3(new_n25023_), .ZN(new_n25026_));
  OAI21_X1   g22590(.A1(new_n24979_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n25027_));
  AOI21_X1   g22591(.A1(new_n25011_), .A2(new_n25021_), .B(pi0625), .ZN(new_n25028_));
  OAI21_X1   g22592(.A1(new_n25028_), .A2(new_n25027_), .B(new_n13560_), .ZN(new_n25029_));
  OAI21_X1   g22593(.A1(new_n25029_), .A2(new_n24950_), .B(pi0778), .ZN(new_n25030_));
  OAI22_X1   g22594(.A1(new_n25026_), .A2(new_n25030_), .B1(pi0778), .B2(new_n25022_), .ZN(new_n25031_));
  NAND2_X1   g22595(.A1(new_n25031_), .A2(new_n12764_), .ZN(new_n25032_));
  INV_X1     g22596(.I(new_n25032_), .ZN(new_n25033_));
  NOR2_X1    g22597(.A1(new_n24983_), .A2(new_n13829_), .ZN(new_n25034_));
  AOI21_X1   g22598(.A1(new_n24954_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n25035_));
  OAI21_X1   g22599(.A1(new_n25031_), .A2(new_n12766_), .B(new_n25035_), .ZN(new_n25036_));
  NAND2_X1   g22600(.A1(new_n25036_), .A2(new_n25034_), .ZN(new_n25037_));
  NOR2_X1    g22601(.A1(new_n24986_), .A2(pi0660), .ZN(new_n25038_));
  AOI21_X1   g22602(.A1(new_n24954_), .A2(pi0609), .B(pi1155), .ZN(new_n25039_));
  OAI21_X1   g22603(.A1(new_n25031_), .A2(pi0609), .B(new_n25039_), .ZN(new_n25040_));
  AOI21_X1   g22604(.A1(new_n25040_), .A2(new_n25038_), .B(new_n12764_), .ZN(new_n25041_));
  AOI21_X1   g22605(.A1(new_n25041_), .A2(new_n25037_), .B(new_n25033_), .ZN(new_n25042_));
  OR2_X2     g22606(.A1(new_n25042_), .A2(pi0781), .Z(new_n25043_));
  OAI21_X1   g22607(.A1(new_n24991_), .A2(pi1154), .B(pi0627), .ZN(new_n25044_));
  AOI21_X1   g22608(.A1(new_n24957_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n25045_));
  NAND2_X1   g22609(.A1(new_n25042_), .A2(pi0618), .ZN(new_n25046_));
  AOI21_X1   g22610(.A1(new_n25046_), .A2(new_n25045_), .B(new_n25044_), .ZN(new_n25047_));
  OAI21_X1   g22611(.A1(new_n24994_), .A2(new_n12785_), .B(new_n12880_), .ZN(new_n25048_));
  OAI21_X1   g22612(.A1(new_n24956_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n25049_));
  AOI21_X1   g22613(.A1(new_n25042_), .A2(new_n12781_), .B(new_n25049_), .ZN(new_n25050_));
  OAI21_X1   g22614(.A1(new_n25050_), .A2(new_n25048_), .B(pi0781), .ZN(new_n25051_));
  OAI21_X1   g22615(.A1(new_n25051_), .A2(new_n25047_), .B(new_n25043_), .ZN(new_n25052_));
  AND2_X2    g22616(.A1(new_n25052_), .A2(new_n12796_), .Z(new_n25053_));
  INV_X1     g22617(.I(new_n24959_), .ZN(new_n25054_));
  AOI21_X1   g22618(.A1(new_n25054_), .A2(new_n12793_), .B(new_n12791_), .ZN(new_n25055_));
  OAI21_X1   g22619(.A1(new_n25052_), .A2(new_n12793_), .B(new_n25055_), .ZN(new_n25056_));
  NAND3_X1   g22620(.A1(new_n25056_), .A2(pi0648), .A3(new_n24999_), .ZN(new_n25057_));
  AOI21_X1   g22621(.A1(new_n25002_), .A2(pi1159), .B(pi0648), .ZN(new_n25058_));
  AOI21_X1   g22622(.A1(new_n25054_), .A2(pi0619), .B(pi1159), .ZN(new_n25059_));
  OAI21_X1   g22623(.A1(new_n25052_), .A2(pi0619), .B(new_n25059_), .ZN(new_n25060_));
  AOI21_X1   g22624(.A1(new_n25060_), .A2(new_n25058_), .B(new_n12796_), .ZN(new_n25061_));
  AOI21_X1   g22625(.A1(new_n25061_), .A2(new_n25057_), .B(new_n25053_), .ZN(new_n25062_));
  OAI21_X1   g22626(.A1(new_n25062_), .A2(new_n12747_), .B(new_n25010_), .ZN(new_n25063_));
  NAND2_X1   g22627(.A1(new_n25063_), .A2(new_n25009_), .ZN(new_n25064_));
  AOI21_X1   g22628(.A1(new_n24944_), .A2(pi0626), .B(new_n12814_), .ZN(new_n25065_));
  NAND2_X1   g22629(.A1(new_n25004_), .A2(new_n12747_), .ZN(new_n25066_));
  AOI21_X1   g22630(.A1(new_n25066_), .A2(new_n25065_), .B(pi1158), .ZN(new_n25067_));
  AOI21_X1   g22631(.A1(new_n24962_), .A2(pi0626), .B(pi0641), .ZN(new_n25068_));
  OAI21_X1   g22632(.A1(new_n25062_), .A2(pi0626), .B(new_n25068_), .ZN(new_n25069_));
  AOI21_X1   g22633(.A1(new_n25069_), .A2(new_n25067_), .B(new_n12808_), .ZN(new_n25070_));
  AND2_X2    g22634(.A1(new_n25062_), .A2(new_n12808_), .Z(new_n25071_));
  AOI21_X1   g22635(.A1(new_n25070_), .A2(new_n25064_), .B(new_n25071_), .ZN(new_n25072_));
  OAI21_X1   g22636(.A1(new_n25072_), .A2(new_n12920_), .B(new_n25006_), .ZN(new_n25073_));
  NAND2_X1   g22637(.A1(new_n25073_), .A2(new_n24967_), .ZN(new_n25074_));
  NOR2_X1    g22638(.A1(new_n24964_), .A2(new_n12920_), .ZN(new_n25075_));
  AOI21_X1   g22639(.A1(new_n12920_), .A2(new_n24944_), .B(new_n25075_), .ZN(new_n25076_));
  NOR2_X1    g22640(.A1(new_n25076_), .A2(new_n12742_), .ZN(new_n25077_));
  NOR2_X1    g22641(.A1(new_n25077_), .A2(pi0629), .ZN(new_n25078_));
  AOI21_X1   g22642(.A1(new_n25005_), .A2(pi0628), .B(pi1156), .ZN(new_n25079_));
  OAI21_X1   g22643(.A1(new_n25072_), .A2(pi0628), .B(new_n25079_), .ZN(new_n25080_));
  AOI21_X1   g22644(.A1(new_n25080_), .A2(new_n25078_), .B(new_n12937_), .ZN(new_n25081_));
  AND2_X2    g22645(.A1(new_n25072_), .A2(new_n12937_), .Z(new_n25082_));
  AOI21_X1   g22646(.A1(new_n25081_), .A2(new_n25074_), .B(new_n25082_), .ZN(new_n25083_));
  OR2_X2     g22647(.A1(new_n25083_), .A2(pi0787), .Z(new_n25084_));
  NAND2_X1   g22648(.A1(new_n24966_), .A2(new_n12742_), .ZN(new_n25085_));
  NOR2_X1    g22649(.A1(new_n25077_), .A2(new_n12937_), .ZN(new_n25086_));
  AOI22_X1   g22650(.A1(new_n25086_), .A2(new_n25085_), .B1(new_n12937_), .B2(new_n24964_), .ZN(new_n25087_));
  NAND2_X1   g22651(.A1(new_n25087_), .A2(new_n12741_), .ZN(new_n25088_));
  NAND2_X1   g22652(.A1(new_n24944_), .A2(pi0647), .ZN(new_n25089_));
  AOI21_X1   g22653(.A1(new_n25088_), .A2(new_n25089_), .B(pi1157), .ZN(new_n25090_));
  OR2_X2     g22654(.A1(new_n25090_), .A2(new_n12981_), .Z(new_n25091_));
  NOR2_X1    g22655(.A1(new_n24944_), .A2(new_n13384_), .ZN(new_n25092_));
  AOI21_X1   g22656(.A1(new_n25005_), .A2(new_n13384_), .B(new_n25092_), .ZN(new_n25093_));
  NOR2_X1    g22657(.A1(new_n25093_), .A2(pi0647), .ZN(new_n25094_));
  NOR2_X1    g22658(.A1(new_n25094_), .A2(new_n12965_), .ZN(new_n25095_));
  NAND2_X1   g22659(.A1(new_n25083_), .A2(pi0647), .ZN(new_n25096_));
  AOI21_X1   g22660(.A1(new_n25096_), .A2(new_n25095_), .B(new_n25091_), .ZN(new_n25097_));
  NAND2_X1   g22661(.A1(new_n25087_), .A2(pi0647), .ZN(new_n25098_));
  OAI21_X1   g22662(.A1(pi0647), .A2(new_n24945_), .B(new_n25098_), .ZN(new_n25099_));
  NAND2_X1   g22663(.A1(new_n25099_), .A2(pi1157), .ZN(new_n25100_));
  NAND2_X1   g22664(.A1(new_n25100_), .A2(new_n12981_), .ZN(new_n25101_));
  OAI21_X1   g22665(.A1(new_n25093_), .A2(new_n12741_), .B(new_n12965_), .ZN(new_n25102_));
  AOI21_X1   g22666(.A1(new_n25083_), .A2(new_n12741_), .B(new_n25102_), .ZN(new_n25103_));
  OAI21_X1   g22667(.A1(new_n25103_), .A2(new_n25101_), .B(pi0787), .ZN(new_n25104_));
  OAI21_X1   g22668(.A1(new_n25104_), .A2(new_n25097_), .B(new_n25084_), .ZN(new_n25105_));
  AND2_X2    g22669(.A1(new_n25105_), .A2(new_n13000_), .Z(new_n25106_));
  AOI21_X1   g22670(.A1(new_n24945_), .A2(pi0644), .B(new_n12740_), .ZN(new_n25107_));
  NOR2_X1    g22671(.A1(new_n24945_), .A2(new_n12985_), .ZN(new_n25108_));
  AOI21_X1   g22672(.A1(new_n25093_), .A2(new_n12985_), .B(new_n25108_), .ZN(new_n25109_));
  NAND2_X1   g22673(.A1(new_n25109_), .A2(new_n12975_), .ZN(new_n25110_));
  AOI21_X1   g22674(.A1(new_n25110_), .A2(new_n25107_), .B(pi1160), .ZN(new_n25111_));
  NAND2_X1   g22675(.A1(new_n25100_), .A2(pi0787), .ZN(new_n25112_));
  OAI22_X1   g22676(.A1(new_n25112_), .A2(new_n25090_), .B1(pi0787), .B2(new_n25087_), .ZN(new_n25113_));
  AOI21_X1   g22677(.A1(new_n25113_), .A2(pi0644), .B(pi0715), .ZN(new_n25114_));
  OAI21_X1   g22678(.A1(new_n25105_), .A2(pi0644), .B(new_n25114_), .ZN(new_n25115_));
  NAND2_X1   g22679(.A1(new_n25115_), .A2(new_n25111_), .ZN(new_n25116_));
  AOI21_X1   g22680(.A1(new_n24945_), .A2(new_n12975_), .B(pi0715), .ZN(new_n25117_));
  NAND2_X1   g22681(.A1(new_n25109_), .A2(pi0644), .ZN(new_n25118_));
  AOI21_X1   g22682(.A1(new_n25118_), .A2(new_n25117_), .B(new_n12739_), .ZN(new_n25119_));
  AOI21_X1   g22683(.A1(new_n25113_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n25120_));
  OAI21_X1   g22684(.A1(new_n25105_), .A2(new_n12975_), .B(new_n25120_), .ZN(new_n25121_));
  AOI21_X1   g22685(.A1(new_n25121_), .A2(new_n25119_), .B(new_n13000_), .ZN(new_n25122_));
  AOI21_X1   g22686(.A1(new_n25122_), .A2(new_n25116_), .B(new_n25106_), .ZN(new_n25123_));
  NAND2_X1   g22687(.A1(po1038), .A2(pi0199), .ZN(new_n25124_));
  OAI21_X1   g22688(.A1(new_n25123_), .A2(po1038), .B(new_n25124_), .ZN(po0356));
  NAND2_X1   g22689(.A1(po1038), .A2(pi0200), .ZN(new_n25126_));
  NOR2_X1    g22690(.A1(new_n13193_), .A2(new_n8531_), .ZN(new_n25127_));
  NOR2_X1    g22691(.A1(new_n25127_), .A2(new_n13384_), .ZN(new_n25128_));
  INV_X1     g22692(.I(new_n25127_), .ZN(new_n25129_));
  NAND2_X1   g22693(.A1(new_n25129_), .A2(new_n12818_), .ZN(new_n25130_));
  INV_X1     g22694(.I(pi0606), .ZN(new_n25131_));
  NOR2_X1    g22695(.A1(new_n2609_), .A2(pi0200), .ZN(new_n25132_));
  INV_X1     g22696(.I(new_n25132_), .ZN(new_n25133_));
  NOR2_X1    g22697(.A1(new_n17986_), .A2(new_n8531_), .ZN(new_n25134_));
  NOR2_X1    g22698(.A1(new_n15784_), .A2(pi0200), .ZN(new_n25135_));
  OAI21_X1   g22699(.A1(new_n25134_), .A2(new_n25135_), .B(new_n3265_), .ZN(new_n25136_));
  OAI21_X1   g22700(.A1(new_n15006_), .A2(pi0200), .B(new_n15011_), .ZN(new_n25137_));
  NAND3_X1   g22701(.A1(new_n25136_), .A2(new_n2609_), .A3(new_n25137_), .ZN(new_n25138_));
  AOI21_X1   g22702(.A1(new_n25138_), .A2(new_n25133_), .B(new_n25131_), .ZN(new_n25139_));
  NOR2_X1    g22703(.A1(new_n25127_), .A2(pi0606), .ZN(new_n25140_));
  NOR3_X1    g22704(.A1(new_n25139_), .A2(new_n12760_), .A3(new_n25140_), .ZN(new_n25141_));
  AOI21_X1   g22705(.A1(new_n12760_), .A2(new_n25127_), .B(new_n25141_), .ZN(new_n25142_));
  NOR2_X1    g22706(.A1(new_n25129_), .A2(new_n12766_), .ZN(new_n25143_));
  NOR2_X1    g22707(.A1(new_n25142_), .A2(pi0609), .ZN(new_n25144_));
  OAI21_X1   g22708(.A1(new_n25144_), .A2(new_n25143_), .B(new_n12770_), .ZN(new_n25145_));
  INV_X1     g22709(.I(new_n25142_), .ZN(new_n25146_));
  NAND2_X1   g22710(.A1(new_n25146_), .A2(pi0609), .ZN(new_n25147_));
  NAND2_X1   g22711(.A1(new_n25127_), .A2(new_n12766_), .ZN(new_n25148_));
  AOI21_X1   g22712(.A1(new_n25147_), .A2(new_n25148_), .B(new_n12770_), .ZN(new_n25149_));
  NOR2_X1    g22713(.A1(new_n25149_), .A2(new_n12764_), .ZN(new_n25150_));
  AOI22_X1   g22714(.A1(new_n25150_), .A2(new_n25145_), .B1(new_n12764_), .B2(new_n25142_), .ZN(new_n25151_));
  NOR2_X1    g22715(.A1(new_n25151_), .A2(new_n15803_), .ZN(new_n25152_));
  NOR3_X1    g22716(.A1(new_n25127_), .A2(new_n12779_), .A3(new_n15238_), .ZN(new_n25153_));
  NOR2_X1    g22717(.A1(new_n25152_), .A2(new_n25153_), .ZN(new_n25154_));
  NOR2_X1    g22718(.A1(new_n25154_), .A2(pi0789), .ZN(new_n25155_));
  NAND2_X1   g22719(.A1(new_n25154_), .A2(new_n12793_), .ZN(new_n25156_));
  NAND2_X1   g22720(.A1(new_n25127_), .A2(pi0619), .ZN(new_n25157_));
  AOI21_X1   g22721(.A1(new_n25156_), .A2(new_n25157_), .B(pi1159), .ZN(new_n25158_));
  NAND2_X1   g22722(.A1(new_n25154_), .A2(pi0619), .ZN(new_n25159_));
  NAND2_X1   g22723(.A1(new_n25127_), .A2(new_n12793_), .ZN(new_n25160_));
  AOI21_X1   g22724(.A1(new_n25159_), .A2(new_n25160_), .B(new_n12791_), .ZN(new_n25161_));
  NOR3_X1    g22725(.A1(new_n25158_), .A2(new_n25161_), .A3(new_n12796_), .ZN(new_n25162_));
  NOR2_X1    g22726(.A1(new_n25162_), .A2(new_n25155_), .ZN(new_n25163_));
  OAI21_X1   g22727(.A1(new_n25163_), .A2(new_n12818_), .B(new_n25130_), .ZN(new_n25164_));
  AOI21_X1   g22728(.A1(new_n25164_), .A2(new_n13384_), .B(new_n25128_), .ZN(new_n25165_));
  NAND2_X1   g22729(.A1(new_n25127_), .A2(pi0625), .ZN(new_n25166_));
  INV_X1     g22730(.I(pi0643), .ZN(new_n25167_));
  NAND2_X1   g22731(.A1(new_n13397_), .A2(pi0200), .ZN(new_n25168_));
  AOI21_X1   g22732(.A1(new_n24931_), .A2(new_n25168_), .B(new_n3265_), .ZN(new_n25169_));
  INV_X1     g22733(.I(new_n25169_), .ZN(new_n25170_));
  NAND2_X1   g22734(.A1(new_n13405_), .A2(pi0200), .ZN(new_n25171_));
  OR2_X2     g22735(.A1(new_n13416_), .A2(pi0200), .Z(new_n25172_));
  AOI21_X1   g22736(.A1(new_n25172_), .A2(new_n25171_), .B(pi0039), .ZN(new_n25173_));
  NOR2_X1    g22737(.A1(new_n13451_), .A2(new_n13445_), .ZN(new_n25174_));
  NOR2_X1    g22738(.A1(new_n25174_), .A2(pi0200), .ZN(new_n25175_));
  AOI21_X1   g22739(.A1(new_n15741_), .A2(new_n13506_), .B(new_n8531_), .ZN(new_n25176_));
  OAI21_X1   g22740(.A1(new_n25176_), .A2(new_n25175_), .B(pi0299), .ZN(new_n25177_));
  AND2_X2    g22741(.A1(new_n13441_), .A2(new_n8531_), .Z(new_n25178_));
  AOI21_X1   g22742(.A1(new_n15739_), .A2(new_n13476_), .B(new_n8531_), .ZN(new_n25179_));
  OAI21_X1   g22743(.A1(new_n25179_), .A2(new_n25178_), .B(new_n2628_), .ZN(new_n25180_));
  AOI21_X1   g22744(.A1(new_n25177_), .A2(new_n25180_), .B(new_n2627_), .ZN(new_n25181_));
  OAI21_X1   g22745(.A1(new_n25181_), .A2(new_n25173_), .B(new_n3265_), .ZN(new_n25182_));
  NAND3_X1   g22746(.A1(new_n25182_), .A2(new_n2609_), .A3(new_n25170_), .ZN(new_n25183_));
  AOI21_X1   g22747(.A1(new_n25183_), .A2(new_n25133_), .B(new_n25167_), .ZN(new_n25184_));
  AOI21_X1   g22748(.A1(new_n25167_), .A2(new_n25129_), .B(new_n25184_), .ZN(new_n25185_));
  NAND2_X1   g22749(.A1(new_n25185_), .A2(new_n13521_), .ZN(new_n25186_));
  AOI21_X1   g22750(.A1(new_n25186_), .A2(new_n25166_), .B(pi1153), .ZN(new_n25187_));
  NAND2_X1   g22751(.A1(new_n25185_), .A2(pi0625), .ZN(new_n25188_));
  NAND2_X1   g22752(.A1(new_n25127_), .A2(new_n13521_), .ZN(new_n25189_));
  AOI21_X1   g22753(.A1(new_n25188_), .A2(new_n25189_), .B(new_n12841_), .ZN(new_n25190_));
  NOR3_X1    g22754(.A1(new_n25187_), .A2(new_n25190_), .A3(new_n12758_), .ZN(new_n25191_));
  NOR2_X1    g22755(.A1(new_n25185_), .A2(pi0778), .ZN(new_n25192_));
  NOR2_X1    g22756(.A1(new_n25191_), .A2(new_n25192_), .ZN(new_n25193_));
  INV_X1     g22757(.I(new_n25193_), .ZN(new_n25194_));
  NAND2_X1   g22758(.A1(new_n25127_), .A2(new_n12869_), .ZN(new_n25195_));
  OAI21_X1   g22759(.A1(new_n25194_), .A2(new_n12869_), .B(new_n25195_), .ZN(new_n25196_));
  NOR2_X1    g22760(.A1(new_n25196_), .A2(new_n12887_), .ZN(new_n25197_));
  AOI21_X1   g22761(.A1(new_n12887_), .A2(new_n25129_), .B(new_n25197_), .ZN(new_n25198_));
  NOR2_X1    g22762(.A1(new_n25129_), .A2(new_n12911_), .ZN(new_n25199_));
  AOI21_X1   g22763(.A1(new_n25198_), .A2(new_n12911_), .B(new_n25199_), .ZN(new_n25200_));
  NOR2_X1    g22764(.A1(new_n25127_), .A2(new_n13392_), .ZN(new_n25201_));
  AOI21_X1   g22765(.A1(new_n25200_), .A2(new_n13392_), .B(new_n25201_), .ZN(new_n25202_));
  NOR2_X1    g22766(.A1(new_n25202_), .A2(pi0792), .ZN(new_n25203_));
  NAND2_X1   g22767(.A1(new_n25202_), .A2(new_n12920_), .ZN(new_n25204_));
  NAND2_X1   g22768(.A1(new_n25127_), .A2(pi0628), .ZN(new_n25205_));
  AOI21_X1   g22769(.A1(new_n25204_), .A2(new_n25205_), .B(pi1156), .ZN(new_n25206_));
  NAND2_X1   g22770(.A1(new_n25202_), .A2(pi0628), .ZN(new_n25207_));
  NAND2_X1   g22771(.A1(new_n25127_), .A2(new_n12920_), .ZN(new_n25208_));
  AOI21_X1   g22772(.A1(new_n25207_), .A2(new_n25208_), .B(new_n12742_), .ZN(new_n25209_));
  NOR3_X1    g22773(.A1(new_n25206_), .A2(new_n25209_), .A3(new_n12937_), .ZN(new_n25210_));
  NOR2_X1    g22774(.A1(new_n25210_), .A2(new_n25203_), .ZN(new_n25211_));
  INV_X1     g22775(.I(new_n25211_), .ZN(new_n25212_));
  NOR2_X1    g22776(.A1(new_n25212_), .A2(pi0647), .ZN(new_n25213_));
  NOR2_X1    g22777(.A1(new_n25129_), .A2(new_n12741_), .ZN(new_n25214_));
  OAI21_X1   g22778(.A1(new_n25213_), .A2(new_n25214_), .B(new_n12965_), .ZN(new_n25215_));
  NAND2_X1   g22779(.A1(new_n25129_), .A2(new_n12741_), .ZN(new_n25216_));
  NAND2_X1   g22780(.A1(new_n25212_), .A2(pi0647), .ZN(new_n25217_));
  NAND2_X1   g22781(.A1(new_n25217_), .A2(new_n25216_), .ZN(new_n25218_));
  OAI22_X1   g22782(.A1(new_n25215_), .A2(new_n12981_), .B1(new_n25218_), .B2(new_n15576_), .ZN(new_n25219_));
  AOI21_X1   g22783(.A1(new_n15608_), .A2(new_n25165_), .B(new_n25219_), .ZN(new_n25220_));
  NOR2_X1    g22784(.A1(new_n25209_), .A2(pi0629), .ZN(new_n25221_));
  NOR2_X1    g22785(.A1(new_n25206_), .A2(new_n12919_), .ZN(new_n25222_));
  OAI22_X1   g22786(.A1(new_n25221_), .A2(new_n25222_), .B1(new_n25164_), .B2(new_n15821_), .ZN(new_n25223_));
  NOR2_X1    g22787(.A1(new_n25163_), .A2(pi0626), .ZN(new_n25224_));
  AOI21_X1   g22788(.A1(pi0626), .A2(new_n25129_), .B(new_n25224_), .ZN(new_n25225_));
  NAND2_X1   g22789(.A1(new_n25129_), .A2(new_n12747_), .ZN(new_n25226_));
  OAI21_X1   g22790(.A1(new_n25163_), .A2(new_n12747_), .B(new_n25226_), .ZN(new_n25227_));
  AOI22_X1   g22791(.A1(new_n25227_), .A2(new_n12812_), .B1(new_n14386_), .B2(new_n25200_), .ZN(new_n25228_));
  OAI21_X1   g22792(.A1(new_n12816_), .A2(new_n25225_), .B(new_n25228_), .ZN(new_n25229_));
  AOI21_X1   g22793(.A1(new_n25229_), .A2(pi0788), .B(new_n15340_), .ZN(new_n25230_));
  NOR2_X1    g22794(.A1(new_n25139_), .A2(new_n25140_), .ZN(new_n25231_));
  NOR2_X1    g22795(.A1(new_n25231_), .A2(pi0643), .ZN(new_n25232_));
  AOI21_X1   g22796(.A1(new_n15115_), .A2(new_n18424_), .B(pi0200), .ZN(new_n25233_));
  NOR2_X1    g22797(.A1(new_n2610_), .A2(pi0606), .ZN(new_n25234_));
  AND3_X2    g22798(.A1(new_n18755_), .A2(pi0200), .A3(new_n18754_), .Z(new_n25235_));
  NOR2_X1    g22799(.A1(new_n15114_), .A2(pi0200), .ZN(new_n25236_));
  OAI21_X1   g22800(.A1(new_n25235_), .A2(new_n25236_), .B(new_n3265_), .ZN(new_n25237_));
  NOR2_X1    g22801(.A1(new_n15109_), .A2(new_n8531_), .ZN(new_n25238_));
  INV_X1     g22802(.I(new_n25238_), .ZN(new_n25239_));
  AOI21_X1   g22803(.A1(new_n25237_), .A2(new_n25239_), .B(new_n2610_), .ZN(new_n25240_));
  NOR4_X1    g22804(.A1(new_n25240_), .A2(new_n25132_), .A3(new_n25233_), .A4(new_n25234_), .ZN(new_n25241_));
  NOR2_X1    g22805(.A1(new_n25018_), .A2(new_n8531_), .ZN(new_n25242_));
  NOR2_X1    g22806(.A1(new_n15119_), .A2(new_n15120_), .ZN(new_n25243_));
  NOR2_X1    g22807(.A1(new_n25243_), .A2(pi0200), .ZN(new_n25244_));
  NOR2_X1    g22808(.A1(new_n25242_), .A2(new_n25244_), .ZN(new_n25245_));
  NOR2_X1    g22809(.A1(new_n13399_), .A2(new_n13571_), .ZN(new_n25246_));
  OAI22_X1   g22810(.A1(new_n25245_), .A2(pi0038), .B1(new_n25170_), .B2(new_n25246_), .ZN(new_n25247_));
  AND2_X2    g22811(.A1(new_n25247_), .A2(new_n25234_), .Z(new_n25248_));
  NOR3_X1    g22812(.A1(new_n25248_), .A2(new_n25241_), .A3(new_n25167_), .ZN(new_n25249_));
  NOR2_X1    g22813(.A1(new_n25249_), .A2(new_n25232_), .ZN(new_n25250_));
  NAND2_X1   g22814(.A1(new_n25250_), .A2(new_n12758_), .ZN(new_n25251_));
  INV_X1     g22815(.I(new_n25251_), .ZN(new_n25252_));
  NAND2_X1   g22816(.A1(new_n25250_), .A2(new_n13521_), .ZN(new_n25253_));
  NAND2_X1   g22817(.A1(new_n25231_), .A2(pi0625), .ZN(new_n25254_));
  AOI21_X1   g22818(.A1(new_n25253_), .A2(new_n25254_), .B(pi1153), .ZN(new_n25255_));
  NOR3_X1    g22819(.A1(new_n25255_), .A2(pi0608), .A3(new_n25190_), .ZN(new_n25256_));
  NAND2_X1   g22820(.A1(new_n25250_), .A2(pi0625), .ZN(new_n25257_));
  NAND2_X1   g22821(.A1(new_n25231_), .A2(new_n13521_), .ZN(new_n25258_));
  AOI21_X1   g22822(.A1(new_n25257_), .A2(new_n25258_), .B(new_n12841_), .ZN(new_n25259_));
  NOR3_X1    g22823(.A1(new_n25259_), .A2(new_n13560_), .A3(new_n25187_), .ZN(new_n25260_));
  NOR3_X1    g22824(.A1(new_n25256_), .A2(new_n25260_), .A3(new_n12758_), .ZN(new_n25261_));
  NOR2_X1    g22825(.A1(new_n25261_), .A2(new_n25252_), .ZN(new_n25262_));
  NOR2_X1    g22826(.A1(new_n25262_), .A2(pi0785), .ZN(new_n25263_));
  NOR2_X1    g22827(.A1(new_n25194_), .A2(pi0609), .ZN(new_n25264_));
  NOR2_X1    g22828(.A1(new_n25262_), .A2(new_n12766_), .ZN(new_n25265_));
  OAI21_X1   g22829(.A1(new_n25265_), .A2(new_n25264_), .B(pi1155), .ZN(new_n25266_));
  NAND3_X1   g22830(.A1(new_n25266_), .A2(pi0660), .A3(new_n25145_), .ZN(new_n25267_));
  OAI21_X1   g22831(.A1(new_n25261_), .A2(new_n25252_), .B(new_n12766_), .ZN(new_n25268_));
  NAND2_X1   g22832(.A1(new_n25193_), .A2(pi0609), .ZN(new_n25269_));
  AOI21_X1   g22833(.A1(new_n25268_), .A2(new_n25269_), .B(pi1155), .ZN(new_n25270_));
  NOR3_X1    g22834(.A1(new_n25270_), .A2(pi0660), .A3(new_n25149_), .ZN(new_n25271_));
  NOR2_X1    g22835(.A1(new_n25271_), .A2(new_n12764_), .ZN(new_n25272_));
  AOI21_X1   g22836(.A1(new_n25272_), .A2(new_n25267_), .B(new_n25263_), .ZN(new_n25273_));
  OAI21_X1   g22837(.A1(new_n25127_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n25274_));
  NOR2_X1    g22838(.A1(new_n25151_), .A2(pi0618), .ZN(new_n25275_));
  OAI21_X1   g22839(.A1(new_n25275_), .A2(new_n25274_), .B(pi0627), .ZN(new_n25276_));
  NOR2_X1    g22840(.A1(new_n25196_), .A2(pi0618), .ZN(new_n25277_));
  NOR2_X1    g22841(.A1(new_n25277_), .A2(new_n12785_), .ZN(new_n25278_));
  NAND2_X1   g22842(.A1(new_n25273_), .A2(pi0618), .ZN(new_n25279_));
  AOI21_X1   g22843(.A1(new_n25279_), .A2(new_n25278_), .B(new_n25276_), .ZN(new_n25280_));
  OAI21_X1   g22844(.A1(new_n25127_), .A2(pi0618), .B(pi1154), .ZN(new_n25281_));
  NOR2_X1    g22845(.A1(new_n25151_), .A2(new_n12781_), .ZN(new_n25282_));
  OAI21_X1   g22846(.A1(new_n25282_), .A2(new_n25281_), .B(new_n12880_), .ZN(new_n25283_));
  OAI21_X1   g22847(.A1(new_n25196_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n25284_));
  AOI21_X1   g22848(.A1(new_n25273_), .A2(new_n12781_), .B(new_n25284_), .ZN(new_n25285_));
  OAI21_X1   g22849(.A1(new_n25285_), .A2(new_n25283_), .B(pi0781), .ZN(new_n25286_));
  OAI22_X1   g22850(.A1(new_n25286_), .A2(new_n25280_), .B1(pi0781), .B2(new_n25273_), .ZN(new_n25287_));
  AOI21_X1   g22851(.A1(new_n25287_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n25288_));
  NAND2_X1   g22852(.A1(new_n25287_), .A2(new_n12793_), .ZN(new_n25289_));
  NAND2_X1   g22853(.A1(new_n25198_), .A2(pi0619), .ZN(new_n25290_));
  AOI21_X1   g22854(.A1(new_n25289_), .A2(new_n25290_), .B(pi1159), .ZN(new_n25291_));
  NOR3_X1    g22855(.A1(new_n25291_), .A2(pi0648), .A3(new_n25161_), .ZN(new_n25292_));
  AND2_X2    g22856(.A1(new_n25198_), .A2(new_n12793_), .Z(new_n25293_));
  AOI21_X1   g22857(.A1(new_n25287_), .A2(pi0619), .B(new_n25293_), .ZN(new_n25294_));
  OAI21_X1   g22858(.A1(new_n25294_), .A2(new_n12791_), .B(pi0648), .ZN(new_n25295_));
  OAI21_X1   g22859(.A1(new_n25295_), .A2(new_n25158_), .B(pi0789), .ZN(new_n25296_));
  OAI21_X1   g22860(.A1(new_n25296_), .A2(new_n25292_), .B(new_n25288_), .ZN(new_n25297_));
  AOI22_X1   g22861(.A1(new_n25297_), .A2(new_n25230_), .B1(pi0792), .B2(new_n25223_), .ZN(new_n25298_));
  OAI22_X1   g22862(.A1(new_n25298_), .A2(new_n15341_), .B1(new_n12972_), .B2(new_n25220_), .ZN(new_n25299_));
  AOI21_X1   g22863(.A1(new_n25129_), .A2(new_n12975_), .B(pi0715), .ZN(new_n25300_));
  NAND2_X1   g22864(.A1(new_n25129_), .A2(new_n12984_), .ZN(new_n25301_));
  OAI21_X1   g22865(.A1(new_n25165_), .A2(new_n12984_), .B(new_n25301_), .ZN(new_n25302_));
  NAND2_X1   g22866(.A1(new_n25302_), .A2(pi0644), .ZN(new_n25303_));
  AOI21_X1   g22867(.A1(new_n25303_), .A2(new_n25300_), .B(new_n12739_), .ZN(new_n25304_));
  NAND3_X1   g22868(.A1(new_n25217_), .A2(pi1157), .A3(new_n25216_), .ZN(new_n25305_));
  NAND3_X1   g22869(.A1(new_n25215_), .A2(new_n25305_), .A3(pi0787), .ZN(new_n25306_));
  OAI21_X1   g22870(.A1(pi0787), .A2(new_n25211_), .B(new_n25306_), .ZN(new_n25307_));
  AOI21_X1   g22871(.A1(new_n25307_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n25308_));
  OAI21_X1   g22872(.A1(new_n25299_), .A2(new_n12975_), .B(new_n25308_), .ZN(new_n25309_));
  NAND2_X1   g22873(.A1(new_n25309_), .A2(new_n25304_), .ZN(new_n25310_));
  AOI21_X1   g22874(.A1(new_n25129_), .A2(pi0644), .B(new_n12740_), .ZN(new_n25311_));
  NAND2_X1   g22875(.A1(new_n25302_), .A2(new_n12975_), .ZN(new_n25312_));
  AOI21_X1   g22876(.A1(new_n25312_), .A2(new_n25311_), .B(pi1160), .ZN(new_n25313_));
  AOI21_X1   g22877(.A1(new_n25307_), .A2(pi0644), .B(pi0715), .ZN(new_n25314_));
  OAI21_X1   g22878(.A1(new_n25299_), .A2(pi0644), .B(new_n25314_), .ZN(new_n25315_));
  AOI21_X1   g22879(.A1(new_n25315_), .A2(new_n25313_), .B(new_n13000_), .ZN(new_n25316_));
  AOI22_X1   g22880(.A1(new_n25316_), .A2(new_n25310_), .B1(new_n13000_), .B2(new_n25299_), .ZN(new_n25317_));
  OAI21_X1   g22881(.A1(new_n25317_), .A2(po1038), .B(new_n25126_), .ZN(po0357));
  INV_X1     g22882(.I(new_n12618_), .ZN(new_n25319_));
  NAND2_X1   g22883(.A1(pi0096), .A2(pi0210), .ZN(new_n25320_));
  OAI21_X1   g22884(.A1(new_n5694_), .A2(new_n25320_), .B(new_n25319_), .ZN(new_n25321_));
  NOR2_X1    g22885(.A1(new_n2742_), .A2(new_n2672_), .ZN(new_n25322_));
  INV_X1     g22886(.I(new_n25322_), .ZN(new_n25323_));
  OAI21_X1   g22887(.A1(new_n5702_), .A2(new_n25323_), .B(new_n12618_), .ZN(new_n25324_));
  NAND2_X1   g22888(.A1(new_n25321_), .A2(new_n25324_), .ZN(new_n25325_));
  INV_X1     g22889(.I(pi0233), .ZN(new_n25326_));
  INV_X1     g22890(.I(pi0237), .ZN(new_n25327_));
  NOR2_X1    g22891(.A1(new_n25326_), .A2(new_n25327_), .ZN(new_n25328_));
  INV_X1     g22892(.I(new_n25328_), .ZN(new_n25329_));
  NOR2_X1    g22893(.A1(new_n25325_), .A2(new_n25329_), .ZN(new_n25330_));
  NAND2_X1   g22894(.A1(new_n25330_), .A2(pi0201), .ZN(new_n25331_));
  NOR2_X1    g22895(.A1(new_n10534_), .A2(pi0332), .ZN(new_n25332_));
  INV_X1     g22896(.I(new_n25332_), .ZN(new_n25333_));
  NOR2_X1    g22897(.A1(new_n2835_), .A2(pi0032), .ZN(new_n25334_));
  AOI21_X1   g22898(.A1(new_n25334_), .A2(new_n2742_), .B(pi0332), .ZN(new_n25335_));
  NOR3_X1    g22899(.A1(new_n2725_), .A2(pi0070), .A3(pi0841), .ZN(new_n25336_));
  NOR2_X1    g22900(.A1(new_n25336_), .A2(new_n25334_), .ZN(new_n25337_));
  OAI21_X1   g22901(.A1(pi0210), .A2(new_n25337_), .B(new_n25335_), .ZN(new_n25338_));
  OAI21_X1   g22902(.A1(new_n25338_), .A2(pi0468), .B(new_n25333_), .ZN(new_n25339_));
  NOR2_X1    g22903(.A1(new_n25339_), .A2(new_n5410_), .ZN(new_n25340_));
  NOR3_X1    g22904(.A1(new_n2742_), .A2(new_n2709_), .A3(new_n2630_), .ZN(new_n25341_));
  INV_X1     g22905(.I(new_n25341_), .ZN(new_n25342_));
  NAND2_X1   g22906(.A1(new_n25338_), .A2(new_n25342_), .ZN(new_n25343_));
  NOR2_X1    g22907(.A1(new_n25343_), .A2(new_n5409_), .ZN(new_n25344_));
  OAI21_X1   g22908(.A1(new_n25340_), .A2(new_n25344_), .B(pi0947), .ZN(new_n25345_));
  NOR2_X1    g22909(.A1(new_n5410_), .A2(pi0332), .ZN(new_n25346_));
  NOR2_X1    g22910(.A1(new_n25346_), .A2(pi0947), .ZN(new_n25347_));
  NOR2_X1    g22911(.A1(new_n25343_), .A2(new_n5398_), .ZN(new_n25348_));
  OAI21_X1   g22912(.A1(new_n25348_), .A2(new_n5409_), .B(new_n25347_), .ZN(new_n25349_));
  NAND2_X1   g22913(.A1(new_n25349_), .A2(new_n25345_), .ZN(new_n25350_));
  NAND2_X1   g22914(.A1(new_n25350_), .A2(new_n5476_), .ZN(new_n25351_));
  OAI21_X1   g22915(.A1(new_n2815_), .A2(pi0095), .B(new_n2835_), .ZN(new_n25352_));
  NAND3_X1   g22916(.A1(new_n25352_), .A2(new_n2725_), .A3(new_n2742_), .ZN(new_n25353_));
  NAND2_X1   g22917(.A1(new_n25353_), .A2(pi0210), .ZN(new_n25354_));
  INV_X1     g22918(.I(new_n25337_), .ZN(new_n25355_));
  AOI21_X1   g22919(.A1(new_n2835_), .A2(new_n3179_), .B(new_n2725_), .ZN(new_n25356_));
  NOR3_X1    g22920(.A1(new_n3079_), .A2(pi0095), .A3(new_n25356_), .ZN(new_n25357_));
  AOI21_X1   g22921(.A1(new_n2814_), .A2(new_n25357_), .B(new_n25355_), .ZN(new_n25358_));
  NAND2_X1   g22922(.A1(new_n25358_), .A2(new_n2709_), .ZN(new_n25359_));
  AOI21_X1   g22923(.A1(new_n25354_), .A2(new_n25359_), .B(pi0332), .ZN(new_n25360_));
  AOI21_X1   g22924(.A1(new_n25360_), .A2(new_n10534_), .B(new_n25332_), .ZN(new_n25361_));
  NAND2_X1   g22925(.A1(new_n25361_), .A2(new_n5409_), .ZN(new_n25362_));
  NOR2_X1    g22926(.A1(new_n25360_), .A2(new_n25341_), .ZN(new_n25363_));
  INV_X1     g22927(.I(new_n25363_), .ZN(new_n25364_));
  OAI21_X1   g22928(.A1(new_n5409_), .A2(new_n25364_), .B(new_n25362_), .ZN(new_n25365_));
  NOR2_X1    g22929(.A1(new_n25364_), .A2(new_n5398_), .ZN(new_n25366_));
  INV_X1     g22930(.I(new_n25366_), .ZN(new_n25367_));
  NAND2_X1   g22931(.A1(new_n25367_), .A2(new_n5410_), .ZN(new_n25368_));
  AOI22_X1   g22932(.A1(new_n25368_), .A2(new_n25347_), .B1(pi0947), .B2(new_n25365_), .ZN(new_n25369_));
  NOR2_X1    g22933(.A1(new_n25369_), .A2(new_n2612_), .ZN(new_n25370_));
  AOI21_X1   g22934(.A1(new_n2612_), .A2(new_n25350_), .B(new_n25370_), .ZN(new_n25371_));
  OR2_X2     g22935(.A1(new_n25371_), .A2(new_n5476_), .Z(new_n25372_));
  AOI21_X1   g22936(.A1(new_n25372_), .A2(new_n25351_), .B(new_n2469_), .ZN(new_n25373_));
  NOR2_X1    g22937(.A1(new_n2661_), .A2(pi0074), .ZN(new_n25374_));
  OAI21_X1   g22938(.A1(pi0198), .A2(new_n25337_), .B(new_n25335_), .ZN(new_n25375_));
  NAND2_X1   g22939(.A1(new_n5727_), .A2(new_n25375_), .ZN(new_n25376_));
  NAND2_X1   g22940(.A1(new_n25376_), .A2(new_n25346_), .ZN(new_n25377_));
  AND3_X2    g22941(.A1(new_n25377_), .A2(new_n2628_), .A3(new_n5701_), .Z(new_n25378_));
  OAI21_X1   g22942(.A1(new_n2630_), .A2(new_n25323_), .B(new_n25375_), .ZN(new_n25379_));
  NAND2_X1   g22943(.A1(new_n25379_), .A2(new_n5410_), .ZN(new_n25380_));
  AOI21_X1   g22944(.A1(new_n25378_), .A2(new_n25380_), .B(new_n25374_), .ZN(new_n25381_));
  NAND2_X1   g22945(.A1(new_n25350_), .A2(pi0299), .ZN(new_n25382_));
  AOI21_X1   g22946(.A1(new_n25381_), .A2(new_n25382_), .B(pi0055), .ZN(new_n25383_));
  NAND2_X1   g22947(.A1(new_n25369_), .A2(pi0299), .ZN(new_n25384_));
  NOR2_X1    g22948(.A1(new_n25346_), .A2(pi0587), .ZN(new_n25385_));
  NOR2_X1    g22949(.A1(new_n25323_), .A2(new_n2630_), .ZN(new_n25386_));
  NAND2_X1   g22950(.A1(new_n25353_), .A2(pi0198), .ZN(new_n25387_));
  NAND2_X1   g22951(.A1(new_n25358_), .A2(new_n2672_), .ZN(new_n25388_));
  AOI21_X1   g22952(.A1(new_n25387_), .A2(new_n25388_), .B(pi0332), .ZN(new_n25389_));
  NOR2_X1    g22953(.A1(new_n25389_), .A2(new_n25386_), .ZN(new_n25390_));
  INV_X1     g22954(.I(new_n25390_), .ZN(new_n25391_));
  OAI21_X1   g22955(.A1(new_n25391_), .A2(new_n5398_), .B(new_n5410_), .ZN(new_n25392_));
  NAND2_X1   g22956(.A1(new_n25392_), .A2(new_n25385_), .ZN(new_n25393_));
  AOI21_X1   g22957(.A1(pi0332), .A2(pi0468), .B(new_n5410_), .ZN(new_n25394_));
  OAI21_X1   g22958(.A1(new_n25389_), .A2(pi0468), .B(new_n25394_), .ZN(new_n25395_));
  NAND2_X1   g22959(.A1(new_n25391_), .A2(new_n5410_), .ZN(new_n25396_));
  NAND3_X1   g22960(.A1(new_n25396_), .A2(pi0587), .A3(new_n25395_), .ZN(new_n25397_));
  NAND3_X1   g22961(.A1(new_n25393_), .A2(new_n25397_), .A3(new_n2628_), .ZN(new_n25398_));
  AOI21_X1   g22962(.A1(new_n25384_), .A2(new_n25398_), .B(new_n12095_), .ZN(new_n25399_));
  INV_X1     g22963(.I(new_n6227_), .ZN(new_n25400_));
  NOR2_X1    g22964(.A1(new_n2800_), .A2(new_n2761_), .ZN(new_n25401_));
  NAND3_X1   g22965(.A1(new_n25401_), .A2(new_n2462_), .A3(new_n2524_), .ZN(new_n25402_));
  NAND2_X1   g22966(.A1(new_n25402_), .A2(new_n2835_), .ZN(new_n25403_));
  NAND3_X1   g22967(.A1(new_n25403_), .A2(new_n2725_), .A3(new_n2742_), .ZN(new_n25404_));
  NAND2_X1   g22968(.A1(new_n25404_), .A2(pi0210), .ZN(new_n25405_));
  AOI21_X1   g22969(.A1(new_n25401_), .A2(new_n25357_), .B(new_n25355_), .ZN(new_n25406_));
  NAND2_X1   g22970(.A1(new_n25406_), .A2(new_n2709_), .ZN(new_n25407_));
  AOI21_X1   g22971(.A1(new_n25405_), .A2(new_n25407_), .B(pi0332), .ZN(new_n25408_));
  NOR2_X1    g22972(.A1(new_n25408_), .A2(new_n25341_), .ZN(new_n25409_));
  INV_X1     g22973(.I(new_n25409_), .ZN(new_n25410_));
  NOR2_X1    g22974(.A1(new_n25410_), .A2(new_n5398_), .ZN(new_n25411_));
  OAI21_X1   g22975(.A1(new_n25411_), .A2(new_n5409_), .B(new_n25347_), .ZN(new_n25412_));
  AOI21_X1   g22976(.A1(new_n25408_), .A2(new_n10534_), .B(new_n25332_), .ZN(new_n25413_));
  AND2_X2    g22977(.A1(new_n25413_), .A2(new_n5409_), .Z(new_n25414_));
  NOR2_X1    g22978(.A1(new_n25410_), .A2(new_n5409_), .ZN(new_n25415_));
  OAI21_X1   g22979(.A1(new_n25414_), .A2(new_n25415_), .B(pi0947), .ZN(new_n25416_));
  NAND3_X1   g22980(.A1(new_n25416_), .A2(new_n25412_), .A3(pi0299), .ZN(new_n25417_));
  NAND2_X1   g22981(.A1(new_n25404_), .A2(pi0198), .ZN(new_n25418_));
  NAND2_X1   g22982(.A1(new_n25406_), .A2(new_n2672_), .ZN(new_n25419_));
  AOI21_X1   g22983(.A1(new_n25418_), .A2(new_n25419_), .B(pi0332), .ZN(new_n25420_));
  NOR2_X1    g22984(.A1(new_n25420_), .A2(new_n25386_), .ZN(new_n25421_));
  INV_X1     g22985(.I(new_n25421_), .ZN(new_n25422_));
  OAI21_X1   g22986(.A1(new_n25422_), .A2(new_n5398_), .B(new_n5410_), .ZN(new_n25423_));
  NAND2_X1   g22987(.A1(new_n25423_), .A2(new_n25385_), .ZN(new_n25424_));
  OAI21_X1   g22988(.A1(new_n25420_), .A2(pi0468), .B(new_n25394_), .ZN(new_n25425_));
  NAND2_X1   g22989(.A1(new_n25422_), .A2(new_n5410_), .ZN(new_n25426_));
  NAND3_X1   g22990(.A1(new_n25426_), .A2(pi0587), .A3(new_n25425_), .ZN(new_n25427_));
  NAND3_X1   g22991(.A1(new_n25424_), .A2(new_n25427_), .A3(new_n2628_), .ZN(new_n25428_));
  AOI21_X1   g22992(.A1(new_n25417_), .A2(new_n25428_), .B(new_n25400_), .ZN(new_n25429_));
  OAI21_X1   g22993(.A1(new_n25429_), .A2(new_n25399_), .B(new_n2625_), .ZN(new_n25430_));
  OAI21_X1   g22994(.A1(new_n25371_), .A2(new_n2602_), .B(new_n2470_), .ZN(new_n25431_));
  AOI21_X1   g22995(.A1(new_n25430_), .A2(new_n25383_), .B(new_n25431_), .ZN(new_n25432_));
  OAI21_X1   g22996(.A1(new_n25350_), .A2(new_n2470_), .B(new_n2469_), .ZN(new_n25433_));
  OAI21_X1   g22997(.A1(new_n25432_), .A2(new_n25433_), .B(new_n2582_), .ZN(new_n25434_));
  OAI22_X1   g22998(.A1(new_n25434_), .A2(new_n25373_), .B1(new_n2582_), .B2(new_n25350_), .ZN(new_n25435_));
  NAND3_X1   g22999(.A1(new_n2531_), .A2(new_n2611_), .A3(new_n5699_), .ZN(new_n25436_));
  OAI21_X1   g23000(.A1(new_n25436_), .A2(new_n5476_), .B(new_n2630_), .ZN(new_n25437_));
  NOR2_X1    g23001(.A1(new_n25437_), .A2(new_n2469_), .ZN(new_n25438_));
  NOR3_X1    g23002(.A1(new_n5704_), .A2(new_n2530_), .A3(new_n2661_), .ZN(new_n25439_));
  OAI22_X1   g23003(.A1(new_n25439_), .A2(pi0332), .B1(pi0054), .B2(new_n2661_), .ZN(new_n25440_));
  NOR2_X1    g23004(.A1(new_n2628_), .A2(pi0947), .ZN(new_n25441_));
  NOR2_X1    g23005(.A1(pi0299), .A2(pi0587), .ZN(new_n25442_));
  NOR3_X1    g23006(.A1(new_n25441_), .A2(pi0468), .A3(new_n25442_), .ZN(new_n25443_));
  AOI21_X1   g23007(.A1(new_n5410_), .A2(pi0468), .B(new_n25443_), .ZN(new_n25444_));
  NOR3_X1    g23008(.A1(new_n2800_), .A2(new_n9142_), .A3(new_n25444_), .ZN(new_n25445_));
  OAI21_X1   g23009(.A1(new_n25445_), .A2(pi0332), .B(new_n6227_), .ZN(new_n25446_));
  NAND3_X1   g23010(.A1(new_n25446_), .A2(new_n2625_), .A3(new_n25440_), .ZN(new_n25447_));
  NAND2_X1   g23011(.A1(new_n2630_), .A2(pi0074), .ZN(new_n25448_));
  AOI21_X1   g23012(.A1(new_n25447_), .A2(new_n25448_), .B(pi0055), .ZN(new_n25449_));
  NAND3_X1   g23013(.A1(new_n25436_), .A2(pi0055), .A3(new_n2630_), .ZN(new_n25450_));
  NAND2_X1   g23014(.A1(new_n25450_), .A2(new_n2470_), .ZN(new_n25451_));
  OAI22_X1   g23015(.A1(new_n25449_), .A2(new_n25451_), .B1(new_n2630_), .B2(new_n2470_), .ZN(new_n25452_));
  OAI21_X1   g23016(.A1(new_n25452_), .A2(pi0059), .B(new_n2582_), .ZN(new_n25453_));
  OAI22_X1   g23017(.A1(new_n25453_), .A2(new_n25438_), .B1(new_n2582_), .B2(new_n2630_), .ZN(new_n25454_));
  NOR2_X1    g23018(.A1(new_n25454_), .A2(new_n25328_), .ZN(new_n25455_));
  AOI21_X1   g23019(.A1(new_n25435_), .A2(new_n25328_), .B(new_n25455_), .ZN(new_n25456_));
  OAI21_X1   g23020(.A1(new_n25456_), .A2(pi0201), .B(new_n25331_), .ZN(po0358));
  NOR2_X1    g23021(.A1(new_n25327_), .A2(pi0233), .ZN(new_n25458_));
  INV_X1     g23022(.I(new_n25458_), .ZN(new_n25459_));
  NOR2_X1    g23023(.A1(new_n25325_), .A2(new_n25459_), .ZN(new_n25460_));
  NAND2_X1   g23024(.A1(new_n25460_), .A2(pi0202), .ZN(new_n25461_));
  NOR2_X1    g23025(.A1(new_n25454_), .A2(new_n25458_), .ZN(new_n25462_));
  AOI21_X1   g23026(.A1(new_n25435_), .A2(new_n25458_), .B(new_n25462_), .ZN(new_n25463_));
  OAI21_X1   g23027(.A1(new_n25463_), .A2(pi0202), .B(new_n25461_), .ZN(po0359));
  NOR2_X1    g23028(.A1(pi0233), .A2(pi0237), .ZN(new_n25465_));
  INV_X1     g23029(.I(new_n25465_), .ZN(new_n25466_));
  NOR2_X1    g23030(.A1(new_n25325_), .A2(new_n25466_), .ZN(new_n25467_));
  NAND2_X1   g23031(.A1(new_n25467_), .A2(pi0203), .ZN(new_n25468_));
  NOR2_X1    g23032(.A1(new_n25454_), .A2(new_n25465_), .ZN(new_n25469_));
  AOI21_X1   g23033(.A1(new_n25435_), .A2(new_n25465_), .B(new_n25469_), .ZN(new_n25470_));
  OAI21_X1   g23034(.A1(new_n25470_), .A2(pi0203), .B(new_n25468_), .ZN(po0360));
  NOR2_X1    g23035(.A1(new_n5475_), .A2(new_n25320_), .ZN(new_n25472_));
  OAI21_X1   g23036(.A1(new_n5488_), .A2(new_n25323_), .B(new_n12618_), .ZN(new_n25473_));
  OAI21_X1   g23037(.A1(new_n12618_), .A2(new_n25472_), .B(new_n25473_), .ZN(new_n25474_));
  NOR2_X1    g23038(.A1(new_n25474_), .A2(new_n25329_), .ZN(new_n25475_));
  NAND2_X1   g23039(.A1(new_n25475_), .A2(pi0204), .ZN(new_n25476_));
  NOR2_X1    g23040(.A1(new_n25339_), .A2(new_n5404_), .ZN(new_n25477_));
  NOR2_X1    g23041(.A1(new_n25343_), .A2(new_n5403_), .ZN(new_n25478_));
  OAI21_X1   g23042(.A1(new_n25477_), .A2(new_n25478_), .B(pi0907), .ZN(new_n25479_));
  AOI21_X1   g23043(.A1(new_n5403_), .A2(new_n2630_), .B(pi0907), .ZN(new_n25480_));
  OAI21_X1   g23044(.A1(new_n25348_), .A2(new_n5403_), .B(new_n25480_), .ZN(new_n25481_));
  NAND2_X1   g23045(.A1(new_n25479_), .A2(new_n25481_), .ZN(new_n25482_));
  INV_X1     g23046(.I(new_n25482_), .ZN(new_n25483_));
  NOR2_X1    g23047(.A1(new_n25483_), .A2(new_n5864_), .ZN(new_n25484_));
  NAND2_X1   g23048(.A1(new_n25361_), .A2(new_n5403_), .ZN(new_n25485_));
  NAND2_X1   g23049(.A1(new_n25363_), .A2(new_n5404_), .ZN(new_n25486_));
  NAND2_X1   g23050(.A1(new_n25485_), .A2(new_n25486_), .ZN(new_n25487_));
  AOI21_X1   g23051(.A1(new_n13119_), .A2(pi0332), .B(new_n12821_), .ZN(new_n25488_));
  NAND2_X1   g23052(.A1(new_n25367_), .A2(new_n25488_), .ZN(new_n25489_));
  AOI22_X1   g23053(.A1(new_n25489_), .A2(new_n25480_), .B1(pi0907), .B2(new_n25487_), .ZN(new_n25490_));
  INV_X1     g23054(.I(new_n25490_), .ZN(new_n25491_));
  NOR2_X1    g23055(.A1(new_n25483_), .A2(new_n2611_), .ZN(new_n25492_));
  AOI21_X1   g23056(.A1(new_n25491_), .A2(new_n2611_), .B(new_n25492_), .ZN(new_n25493_));
  NOR2_X1    g23057(.A1(new_n25493_), .A2(new_n5476_), .ZN(new_n25494_));
  OAI21_X1   g23058(.A1(new_n25494_), .A2(new_n25484_), .B(pi0059), .ZN(new_n25495_));
  NAND2_X1   g23059(.A1(new_n25483_), .A2(pi0299), .ZN(new_n25496_));
  NOR2_X1    g23060(.A1(new_n5403_), .A2(new_n25323_), .ZN(new_n25497_));
  OAI21_X1   g23061(.A1(new_n25497_), .A2(new_n2630_), .B(new_n2628_), .ZN(new_n25498_));
  INV_X1     g23062(.I(new_n25498_), .ZN(new_n25499_));
  NAND2_X1   g23063(.A1(new_n10534_), .A2(new_n5486_), .ZN(new_n25500_));
  OAI21_X1   g23064(.A1(new_n5404_), .A2(new_n10534_), .B(new_n25500_), .ZN(new_n25501_));
  OAI21_X1   g23065(.A1(new_n25501_), .A2(new_n25379_), .B(new_n25499_), .ZN(new_n25502_));
  AOI21_X1   g23066(.A1(new_n25496_), .A2(new_n25502_), .B(new_n25374_), .ZN(new_n25503_));
  OAI21_X1   g23067(.A1(new_n25411_), .A2(new_n5403_), .B(new_n25480_), .ZN(new_n25504_));
  NAND2_X1   g23068(.A1(new_n25413_), .A2(new_n5403_), .ZN(new_n25505_));
  NAND2_X1   g23069(.A1(new_n25409_), .A2(new_n5404_), .ZN(new_n25506_));
  NAND2_X1   g23070(.A1(new_n25505_), .A2(new_n25506_), .ZN(new_n25507_));
  NAND2_X1   g23071(.A1(new_n25507_), .A2(pi0907), .ZN(new_n25508_));
  AND3_X2    g23072(.A1(new_n25508_), .A2(pi0299), .A3(new_n25504_), .Z(new_n25509_));
  AOI21_X1   g23073(.A1(new_n25421_), .A2(new_n5489_), .B(new_n25498_), .ZN(new_n25510_));
  OAI21_X1   g23074(.A1(new_n25509_), .A2(new_n25510_), .B(new_n6227_), .ZN(new_n25511_));
  NOR2_X1    g23075(.A1(new_n25491_), .A2(new_n2628_), .ZN(new_n25512_));
  AOI21_X1   g23076(.A1(new_n25390_), .A2(new_n5489_), .B(new_n25498_), .ZN(new_n25513_));
  OAI21_X1   g23077(.A1(new_n25512_), .A2(new_n25513_), .B(new_n12094_), .ZN(new_n25514_));
  AOI21_X1   g23078(.A1(new_n25511_), .A2(new_n25514_), .B(pi0074), .ZN(new_n25515_));
  NOR3_X1    g23079(.A1(new_n25515_), .A2(pi0055), .A3(new_n25503_), .ZN(new_n25516_));
  OAI21_X1   g23080(.A1(new_n25493_), .A2(new_n2602_), .B(new_n2470_), .ZN(new_n25517_));
  AOI21_X1   g23081(.A1(new_n25483_), .A2(new_n2471_), .B(pi0059), .ZN(new_n25518_));
  OAI21_X1   g23082(.A1(new_n25516_), .A2(new_n25517_), .B(new_n25518_), .ZN(new_n25519_));
  NAND3_X1   g23083(.A1(new_n25519_), .A2(new_n2582_), .A3(new_n25495_), .ZN(new_n25520_));
  OAI21_X1   g23084(.A1(new_n2582_), .A2(new_n25482_), .B(new_n25520_), .ZN(new_n25521_));
  NAND3_X1   g23085(.A1(new_n2531_), .A2(new_n2611_), .A3(new_n5548_), .ZN(new_n25522_));
  OAI21_X1   g23086(.A1(new_n25522_), .A2(new_n5476_), .B(new_n2630_), .ZN(new_n25523_));
  NOR2_X1    g23087(.A1(new_n25523_), .A2(new_n2469_), .ZN(new_n25524_));
  NOR2_X1    g23088(.A1(new_n2470_), .A2(new_n2630_), .ZN(new_n25525_));
  NAND3_X1   g23089(.A1(new_n25522_), .A2(pi0055), .A3(new_n2630_), .ZN(new_n25526_));
  NAND2_X1   g23090(.A1(new_n25526_), .A2(new_n2470_), .ZN(new_n25527_));
  NOR2_X1    g23091(.A1(new_n25374_), .A2(new_n2630_), .ZN(new_n25528_));
  NOR2_X1    g23092(.A1(new_n25528_), .A2(pi0055), .ZN(new_n25529_));
  NOR2_X1    g23093(.A1(new_n25501_), .A2(pi0299), .ZN(new_n25530_));
  OAI21_X1   g23094(.A1(new_n5485_), .A2(new_n25530_), .B(new_n2531_), .ZN(new_n25531_));
  AOI21_X1   g23095(.A1(new_n25531_), .A2(new_n2630_), .B(new_n12095_), .ZN(new_n25532_));
  NOR2_X1    g23096(.A1(new_n2628_), .A2(new_n5473_), .ZN(new_n25533_));
  NOR2_X1    g23097(.A1(new_n5486_), .A2(pi0299), .ZN(new_n25534_));
  NOR3_X1    g23098(.A1(new_n25533_), .A2(new_n25534_), .A3(pi0468), .ZN(new_n25535_));
  AOI21_X1   g23099(.A1(new_n5403_), .A2(pi0468), .B(new_n25535_), .ZN(new_n25536_));
  NAND3_X1   g23100(.A1(new_n2801_), .A2(new_n8970_), .A3(new_n25536_), .ZN(new_n25537_));
  AOI21_X1   g23101(.A1(new_n25537_), .A2(new_n2630_), .B(new_n25400_), .ZN(new_n25538_));
  OAI21_X1   g23102(.A1(new_n25538_), .A2(new_n25532_), .B(new_n2625_), .ZN(new_n25539_));
  AOI21_X1   g23103(.A1(new_n25539_), .A2(new_n25529_), .B(new_n25527_), .ZN(new_n25540_));
  OR3_X2     g23104(.A1(new_n25540_), .A2(pi0059), .A3(new_n25525_), .Z(new_n25541_));
  NAND2_X1   g23105(.A1(new_n25541_), .A2(new_n2582_), .ZN(new_n25542_));
  OAI22_X1   g23106(.A1(new_n25542_), .A2(new_n25524_), .B1(new_n2582_), .B2(new_n2630_), .ZN(new_n25543_));
  NOR2_X1    g23107(.A1(new_n25543_), .A2(new_n25328_), .ZN(new_n25544_));
  AOI21_X1   g23108(.A1(new_n25521_), .A2(new_n25328_), .B(new_n25544_), .ZN(new_n25545_));
  OAI21_X1   g23109(.A1(new_n25545_), .A2(pi0204), .B(new_n25476_), .ZN(po0361));
  NOR2_X1    g23110(.A1(new_n25474_), .A2(new_n25459_), .ZN(new_n25547_));
  NAND2_X1   g23111(.A1(new_n25547_), .A2(pi0205), .ZN(new_n25548_));
  NOR2_X1    g23112(.A1(new_n25543_), .A2(new_n25458_), .ZN(new_n25549_));
  AOI21_X1   g23113(.A1(new_n25521_), .A2(new_n25458_), .B(new_n25549_), .ZN(new_n25550_));
  OAI21_X1   g23114(.A1(new_n25550_), .A2(pi0205), .B(new_n25548_), .ZN(po0362));
  NOR2_X1    g23115(.A1(new_n25326_), .A2(pi0237), .ZN(new_n25552_));
  INV_X1     g23116(.I(new_n25552_), .ZN(new_n25553_));
  NOR2_X1    g23117(.A1(new_n25474_), .A2(new_n25553_), .ZN(new_n25554_));
  NAND2_X1   g23118(.A1(new_n25554_), .A2(pi0206), .ZN(new_n25555_));
  NOR2_X1    g23119(.A1(new_n25543_), .A2(new_n25552_), .ZN(new_n25556_));
  AOI21_X1   g23120(.A1(new_n25521_), .A2(new_n25552_), .B(new_n25556_), .ZN(new_n25557_));
  OAI21_X1   g23121(.A1(new_n25557_), .A2(pi0206), .B(new_n25555_), .ZN(po0363));
  NOR2_X1    g23122(.A1(new_n18327_), .A2(new_n2610_), .ZN(new_n25559_));
  NAND2_X1   g23123(.A1(new_n25559_), .A2(new_n12761_), .ZN(new_n25560_));
  NOR2_X1    g23124(.A1(new_n25560_), .A2(new_n15232_), .ZN(new_n25561_));
  INV_X1     g23125(.I(new_n25561_), .ZN(new_n25562_));
  NOR3_X1    g23126(.A1(new_n25562_), .A2(new_n15239_), .A3(new_n15244_), .ZN(new_n25563_));
  NAND2_X1   g23127(.A1(new_n25563_), .A2(new_n17504_), .ZN(new_n25564_));
  NOR2_X1    g23128(.A1(new_n25564_), .A2(new_n12943_), .ZN(new_n25565_));
  NAND2_X1   g23129(.A1(new_n25565_), .A2(pi0207), .ZN(new_n25566_));
  NOR2_X1    g23130(.A1(new_n13193_), .A2(new_n13384_), .ZN(new_n25567_));
  NAND2_X1   g23131(.A1(new_n15013_), .A2(new_n2609_), .ZN(new_n25568_));
  NAND2_X1   g23132(.A1(new_n25568_), .A2(new_n12761_), .ZN(new_n25569_));
  OAI21_X1   g23133(.A1(new_n12761_), .A2(new_n13193_), .B(new_n25569_), .ZN(new_n25570_));
  NOR2_X1    g23134(.A1(new_n25570_), .A2(pi0785), .ZN(new_n25571_));
  NOR2_X1    g23135(.A1(new_n25569_), .A2(pi0609), .ZN(new_n25572_));
  NOR2_X1    g23136(.A1(new_n13193_), .A2(new_n13353_), .ZN(new_n25573_));
  OAI21_X1   g23137(.A1(new_n25572_), .A2(new_n25573_), .B(new_n12770_), .ZN(new_n25574_));
  OAI22_X1   g23138(.A1(new_n25569_), .A2(new_n12766_), .B1(new_n13193_), .B2(new_n12772_), .ZN(new_n25575_));
  AOI21_X1   g23139(.A1(new_n25575_), .A2(pi1155), .B(new_n12764_), .ZN(new_n25576_));
  AOI21_X1   g23140(.A1(new_n25576_), .A2(new_n25574_), .B(new_n25571_), .ZN(new_n25577_));
  NOR2_X1    g23141(.A1(new_n25577_), .A2(pi0781), .ZN(new_n25578_));
  NAND2_X1   g23142(.A1(new_n25577_), .A2(pi0618), .ZN(new_n25579_));
  NAND2_X1   g23143(.A1(new_n13192_), .A2(new_n12781_), .ZN(new_n25580_));
  AOI21_X1   g23144(.A1(new_n25579_), .A2(new_n25580_), .B(new_n12785_), .ZN(new_n25581_));
  NOR2_X1    g23145(.A1(new_n13193_), .A2(new_n12781_), .ZN(new_n25582_));
  AOI21_X1   g23146(.A1(new_n25577_), .A2(new_n12781_), .B(new_n25582_), .ZN(new_n25583_));
  OAI21_X1   g23147(.A1(new_n25583_), .A2(pi1154), .B(pi0781), .ZN(new_n25584_));
  NOR2_X1    g23148(.A1(new_n25584_), .A2(new_n25581_), .ZN(new_n25585_));
  NOR2_X1    g23149(.A1(new_n25585_), .A2(new_n25578_), .ZN(new_n25586_));
  INV_X1     g23150(.I(new_n25586_), .ZN(new_n25587_));
  NAND2_X1   g23151(.A1(new_n13192_), .A2(new_n12793_), .ZN(new_n25588_));
  OAI21_X1   g23152(.A1(new_n25587_), .A2(new_n12793_), .B(new_n25588_), .ZN(new_n25589_));
  NAND2_X1   g23153(.A1(new_n25589_), .A2(pi1159), .ZN(new_n25590_));
  NOR2_X1    g23154(.A1(new_n13193_), .A2(new_n12793_), .ZN(new_n25591_));
  AOI21_X1   g23155(.A1(new_n25586_), .A2(new_n12793_), .B(new_n25591_), .ZN(new_n25592_));
  NOR2_X1    g23156(.A1(new_n25592_), .A2(pi1159), .ZN(new_n25593_));
  NOR2_X1    g23157(.A1(new_n25593_), .A2(new_n12796_), .ZN(new_n25594_));
  AOI22_X1   g23158(.A1(new_n25594_), .A2(new_n25590_), .B1(new_n12796_), .B2(new_n25587_), .ZN(new_n25595_));
  INV_X1     g23159(.I(new_n25595_), .ZN(new_n25596_));
  NAND2_X1   g23160(.A1(new_n13192_), .A2(new_n12818_), .ZN(new_n25597_));
  OAI21_X1   g23161(.A1(new_n25596_), .A2(new_n12818_), .B(new_n25597_), .ZN(new_n25598_));
  AND2_X2    g23162(.A1(new_n25598_), .A2(new_n13384_), .Z(new_n25599_));
  NOR2_X1    g23163(.A1(new_n25599_), .A2(new_n25567_), .ZN(new_n25600_));
  OAI21_X1   g23164(.A1(new_n25600_), .A2(pi0207), .B(new_n25566_), .ZN(new_n25601_));
  NOR2_X1    g23165(.A1(new_n13193_), .A2(pi0207), .ZN(new_n25602_));
  INV_X1     g23166(.I(new_n25602_), .ZN(new_n25603_));
  NOR2_X1    g23167(.A1(new_n25603_), .A2(pi0623), .ZN(new_n25604_));
  AOI21_X1   g23168(.A1(new_n25601_), .A2(pi0623), .B(new_n25604_), .ZN(new_n25605_));
  INV_X1     g23169(.I(new_n25605_), .ZN(new_n25606_));
  INV_X1     g23170(.I(pi0710), .ZN(new_n25607_));
  NOR2_X1    g23171(.A1(new_n18371_), .A2(new_n14285_), .ZN(new_n25608_));
  INV_X1     g23172(.I(new_n25608_), .ZN(new_n25609_));
  NOR2_X1    g23173(.A1(new_n25609_), .A2(new_n14292_), .ZN(new_n25610_));
  NAND2_X1   g23174(.A1(new_n25610_), .A2(new_n12952_), .ZN(new_n25611_));
  INV_X1     g23175(.I(new_n25611_), .ZN(new_n25612_));
  NAND2_X1   g23176(.A1(new_n25612_), .A2(pi0207), .ZN(new_n25613_));
  NOR2_X1    g23177(.A1(new_n24217_), .A2(new_n2610_), .ZN(new_n25614_));
  NOR2_X1    g23178(.A1(new_n25614_), .A2(pi0625), .ZN(new_n25615_));
  OAI21_X1   g23179(.A1(new_n25615_), .A2(new_n14163_), .B(new_n12841_), .ZN(new_n25616_));
  NAND2_X1   g23180(.A1(new_n18367_), .A2(new_n2609_), .ZN(new_n25617_));
  NAND2_X1   g23181(.A1(new_n25617_), .A2(pi0625), .ZN(new_n25618_));
  AOI21_X1   g23182(.A1(new_n25618_), .A2(new_n19435_), .B(new_n12841_), .ZN(new_n25619_));
  NOR2_X1    g23183(.A1(new_n25619_), .A2(new_n12758_), .ZN(new_n25620_));
  AOI22_X1   g23184(.A1(new_n25620_), .A2(new_n25616_), .B1(new_n12758_), .B2(new_n25614_), .ZN(new_n25621_));
  NOR2_X1    g23185(.A1(new_n25621_), .A2(new_n12869_), .ZN(new_n25622_));
  AOI21_X1   g23186(.A1(new_n12869_), .A2(new_n13193_), .B(new_n25622_), .ZN(new_n25623_));
  NAND2_X1   g23187(.A1(new_n25623_), .A2(new_n12888_), .ZN(new_n25624_));
  OAI21_X1   g23188(.A1(new_n12888_), .A2(new_n13193_), .B(new_n25624_), .ZN(new_n25625_));
  NOR2_X1    g23189(.A1(new_n25625_), .A2(new_n12910_), .ZN(new_n25626_));
  AOI21_X1   g23190(.A1(new_n12910_), .A2(new_n13193_), .B(new_n25626_), .ZN(new_n25627_));
  INV_X1     g23191(.I(new_n25627_), .ZN(new_n25628_));
  NAND2_X1   g23192(.A1(new_n13192_), .A2(new_n12817_), .ZN(new_n25629_));
  OAI21_X1   g23193(.A1(new_n25628_), .A2(new_n12817_), .B(new_n25629_), .ZN(new_n25630_));
  NOR2_X1    g23194(.A1(new_n25630_), .A2(new_n12951_), .ZN(new_n25631_));
  AOI21_X1   g23195(.A1(new_n12951_), .A2(new_n13193_), .B(new_n25631_), .ZN(new_n25632_));
  NAND2_X1   g23196(.A1(new_n25632_), .A2(new_n8521_), .ZN(new_n25633_));
  AOI21_X1   g23197(.A1(new_n25633_), .A2(new_n25613_), .B(new_n25607_), .ZN(new_n25634_));
  NOR2_X1    g23198(.A1(new_n25603_), .A2(pi0710), .ZN(new_n25635_));
  NOR2_X1    g23199(.A1(new_n25634_), .A2(new_n25635_), .ZN(new_n25636_));
  NAND2_X1   g23200(.A1(new_n25636_), .A2(new_n12741_), .ZN(new_n25637_));
  NAND2_X1   g23201(.A1(new_n25603_), .A2(pi0647), .ZN(new_n25638_));
  AOI21_X1   g23202(.A1(new_n25637_), .A2(new_n25638_), .B(pi1157), .ZN(new_n25639_));
  INV_X1     g23203(.I(new_n25636_), .ZN(new_n25640_));
  NOR2_X1    g23204(.A1(new_n25640_), .A2(new_n12741_), .ZN(new_n25641_));
  NOR2_X1    g23205(.A1(new_n25602_), .A2(pi0647), .ZN(new_n25642_));
  OAI21_X1   g23206(.A1(new_n25641_), .A2(new_n25642_), .B(pi1157), .ZN(new_n25643_));
  NAND2_X1   g23207(.A1(new_n25643_), .A2(new_n12981_), .ZN(new_n25644_));
  OAI21_X1   g23208(.A1(new_n12981_), .A2(new_n25639_), .B(new_n25644_), .ZN(new_n25645_));
  OAI21_X1   g23209(.A1(new_n17212_), .A2(new_n25606_), .B(new_n25645_), .ZN(new_n25646_));
  AOI21_X1   g23210(.A1(new_n25606_), .A2(new_n25607_), .B(new_n15341_), .ZN(new_n25647_));
  INV_X1     g23211(.I(pi0623), .ZN(new_n25648_));
  NAND3_X1   g23212(.A1(new_n25610_), .A2(new_n12943_), .A3(new_n18389_), .ZN(new_n25649_));
  NOR2_X1    g23213(.A1(new_n25609_), .A2(new_n12869_), .ZN(new_n25650_));
  INV_X1     g23214(.I(new_n25650_), .ZN(new_n25651_));
  AOI21_X1   g23215(.A1(new_n25651_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n25652_));
  NOR2_X1    g23216(.A1(new_n18371_), .A2(pi0625), .ZN(new_n25653_));
  OAI21_X1   g23217(.A1(new_n25653_), .A2(pi1153), .B(pi0608), .ZN(new_n25654_));
  INV_X1     g23218(.I(new_n25654_), .ZN(new_n25655_));
  OAI21_X1   g23219(.A1(new_n25016_), .A2(new_n13521_), .B(pi1153), .ZN(new_n25656_));
  NAND2_X1   g23220(.A1(new_n25655_), .A2(new_n25656_), .ZN(new_n25657_));
  NOR2_X1    g23221(.A1(new_n18371_), .A2(new_n13521_), .ZN(new_n25658_));
  OAI21_X1   g23222(.A1(new_n25658_), .A2(new_n12841_), .B(new_n13560_), .ZN(new_n25659_));
  INV_X1     g23223(.I(new_n25659_), .ZN(new_n25660_));
  OAI21_X1   g23224(.A1(new_n25016_), .A2(pi0625), .B(new_n12841_), .ZN(new_n25661_));
  AOI21_X1   g23225(.A1(new_n25660_), .A2(new_n25661_), .B(new_n12758_), .ZN(new_n25662_));
  AOI22_X1   g23226(.A1(new_n25662_), .A2(new_n25657_), .B1(new_n12758_), .B2(new_n25016_), .ZN(new_n25663_));
  AOI21_X1   g23227(.A1(new_n25609_), .A2(new_n12766_), .B(new_n12770_), .ZN(new_n25664_));
  INV_X1     g23228(.I(new_n25663_), .ZN(new_n25665_));
  NAND2_X1   g23229(.A1(new_n25665_), .A2(pi0609), .ZN(new_n25666_));
  NAND3_X1   g23230(.A1(new_n25666_), .A2(pi0660), .A3(new_n25664_), .ZN(new_n25667_));
  AOI21_X1   g23231(.A1(new_n25609_), .A2(pi0609), .B(pi1155), .ZN(new_n25668_));
  NAND2_X1   g23232(.A1(new_n25665_), .A2(new_n12766_), .ZN(new_n25669_));
  NAND3_X1   g23233(.A1(new_n25669_), .A2(new_n13829_), .A3(new_n25668_), .ZN(new_n25670_));
  NAND3_X1   g23234(.A1(new_n25667_), .A2(new_n25670_), .A3(pi0785), .ZN(new_n25671_));
  OAI21_X1   g23235(.A1(pi0785), .A2(new_n25663_), .B(new_n25671_), .ZN(new_n25672_));
  NAND2_X1   g23236(.A1(new_n25672_), .A2(pi0618), .ZN(new_n25673_));
  NAND3_X1   g23237(.A1(new_n25673_), .A2(pi0627), .A3(new_n25652_), .ZN(new_n25674_));
  AOI21_X1   g23238(.A1(new_n25651_), .A2(pi0618), .B(pi1154), .ZN(new_n25675_));
  NAND2_X1   g23239(.A1(new_n25672_), .A2(new_n12781_), .ZN(new_n25676_));
  NAND3_X1   g23240(.A1(new_n25676_), .A2(new_n12880_), .A3(new_n25675_), .ZN(new_n25677_));
  NAND3_X1   g23241(.A1(new_n25677_), .A2(new_n25674_), .A3(pi0781), .ZN(new_n25678_));
  AOI21_X1   g23242(.A1(new_n25672_), .A2(new_n12779_), .B(new_n17591_), .ZN(new_n25679_));
  NAND2_X1   g23243(.A1(new_n25678_), .A2(new_n25679_), .ZN(new_n25680_));
  NOR2_X1    g23244(.A1(new_n25609_), .A2(new_n14290_), .ZN(new_n25681_));
  NAND3_X1   g23245(.A1(new_n25681_), .A2(pi0789), .A3(new_n17599_), .ZN(new_n25682_));
  NAND2_X1   g23246(.A1(new_n25680_), .A2(new_n25682_), .ZN(new_n25683_));
  OAI21_X1   g23247(.A1(new_n25683_), .A2(pi0788), .B(new_n15824_), .ZN(new_n25684_));
  NOR3_X1    g23248(.A1(new_n25609_), .A2(new_n12910_), .A3(new_n14290_), .ZN(new_n25685_));
  OAI21_X1   g23249(.A1(new_n25685_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n25686_));
  NOR2_X1    g23250(.A1(new_n25683_), .A2(pi0626), .ZN(new_n25687_));
  NOR3_X1    g23251(.A1(new_n25687_), .A2(pi1158), .A3(new_n25686_), .ZN(new_n25688_));
  NAND2_X1   g23252(.A1(new_n25685_), .A2(new_n12747_), .ZN(new_n25689_));
  INV_X1     g23253(.I(new_n25689_), .ZN(new_n25690_));
  AOI21_X1   g23254(.A1(new_n25683_), .A2(pi0626), .B(new_n25690_), .ZN(new_n25691_));
  OAI21_X1   g23255(.A1(new_n25691_), .A2(new_n13557_), .B(pi0788), .ZN(new_n25692_));
  NOR2_X1    g23256(.A1(new_n25692_), .A2(new_n25688_), .ZN(new_n25693_));
  OAI21_X1   g23257(.A1(new_n25693_), .A2(new_n25684_), .B(new_n25649_), .ZN(new_n25694_));
  INV_X1     g23258(.I(new_n25694_), .ZN(new_n25695_));
  OAI21_X1   g23259(.A1(new_n25695_), .A2(new_n8521_), .B(new_n25648_), .ZN(new_n25696_));
  NAND2_X1   g23260(.A1(new_n13192_), .A2(pi0628), .ZN(new_n25697_));
  NAND2_X1   g23261(.A1(new_n25630_), .A2(new_n12920_), .ZN(new_n25698_));
  AOI21_X1   g23262(.A1(new_n25698_), .A2(new_n25697_), .B(new_n18088_), .ZN(new_n25699_));
  AOI21_X1   g23263(.A1(new_n12949_), .A2(new_n13192_), .B(new_n25699_), .ZN(new_n25700_));
  NOR2_X1    g23264(.A1(new_n25630_), .A2(new_n12920_), .ZN(new_n25701_));
  AOI21_X1   g23265(.A1(new_n12920_), .A2(new_n13193_), .B(new_n25701_), .ZN(new_n25702_));
  AOI21_X1   g23266(.A1(pi0628), .A2(pi0629), .B(new_n12742_), .ZN(new_n25703_));
  NAND2_X1   g23267(.A1(new_n25702_), .A2(new_n25703_), .ZN(new_n25704_));
  NAND2_X1   g23268(.A1(new_n25700_), .A2(new_n25704_), .ZN(new_n25705_));
  NAND2_X1   g23269(.A1(new_n25621_), .A2(new_n12766_), .ZN(new_n25706_));
  NOR2_X1    g23270(.A1(new_n18418_), .A2(new_n2610_), .ZN(new_n25707_));
  INV_X1     g23271(.I(new_n25707_), .ZN(new_n25708_));
  NOR2_X1    g23272(.A1(new_n25707_), .A2(new_n13521_), .ZN(new_n25709_));
  OAI21_X1   g23273(.A1(new_n25709_), .A2(new_n14199_), .B(pi1153), .ZN(new_n25710_));
  NAND3_X1   g23274(.A1(new_n25616_), .A2(new_n25710_), .A3(pi0608), .ZN(new_n25711_));
  OAI21_X1   g23275(.A1(new_n25707_), .A2(pi0625), .B(new_n19427_), .ZN(new_n25712_));
  AOI21_X1   g23276(.A1(new_n25712_), .A2(new_n12841_), .B(new_n25619_), .ZN(new_n25713_));
  AOI21_X1   g23277(.A1(new_n25713_), .A2(new_n13560_), .B(new_n12758_), .ZN(new_n25714_));
  AOI22_X1   g23278(.A1(new_n25714_), .A2(new_n25711_), .B1(new_n12758_), .B2(new_n25708_), .ZN(new_n25715_));
  OAI21_X1   g23279(.A1(new_n25715_), .A2(new_n12766_), .B(new_n25706_), .ZN(new_n25716_));
  NAND2_X1   g23280(.A1(new_n13193_), .A2(new_n12770_), .ZN(new_n25717_));
  OAI21_X1   g23281(.A1(new_n25716_), .A2(new_n12770_), .B(new_n25717_), .ZN(new_n25718_));
  NAND2_X1   g23282(.A1(new_n25718_), .A2(pi0660), .ZN(new_n25719_));
  NAND2_X1   g23283(.A1(new_n13193_), .A2(pi1155), .ZN(new_n25720_));
  NAND2_X1   g23284(.A1(new_n25621_), .A2(pi0609), .ZN(new_n25721_));
  OAI21_X1   g23285(.A1(new_n25715_), .A2(pi0609), .B(new_n25721_), .ZN(new_n25722_));
  OAI21_X1   g23286(.A1(new_n25722_), .A2(pi1155), .B(new_n25720_), .ZN(new_n25723_));
  AOI21_X1   g23287(.A1(new_n25723_), .A2(new_n13829_), .B(new_n12764_), .ZN(new_n25724_));
  NOR2_X1    g23288(.A1(new_n25715_), .A2(pi0785), .ZN(new_n25725_));
  AOI21_X1   g23289(.A1(new_n25724_), .A2(new_n25719_), .B(new_n25725_), .ZN(new_n25726_));
  NOR2_X1    g23290(.A1(new_n25726_), .A2(pi0781), .ZN(new_n25727_));
  NAND2_X1   g23291(.A1(new_n25623_), .A2(new_n12781_), .ZN(new_n25728_));
  OAI21_X1   g23292(.A1(new_n25726_), .A2(new_n12781_), .B(new_n25728_), .ZN(new_n25729_));
  NAND2_X1   g23293(.A1(new_n13193_), .A2(new_n12785_), .ZN(new_n25730_));
  OAI21_X1   g23294(.A1(new_n25729_), .A2(new_n12785_), .B(new_n25730_), .ZN(new_n25731_));
  NAND2_X1   g23295(.A1(new_n25731_), .A2(pi0627), .ZN(new_n25732_));
  NAND2_X1   g23296(.A1(new_n13193_), .A2(pi1154), .ZN(new_n25733_));
  NAND2_X1   g23297(.A1(new_n25623_), .A2(pi0618), .ZN(new_n25734_));
  OAI21_X1   g23298(.A1(new_n25726_), .A2(pi0618), .B(new_n25734_), .ZN(new_n25735_));
  OAI21_X1   g23299(.A1(new_n25735_), .A2(pi1154), .B(new_n25733_), .ZN(new_n25736_));
  AOI21_X1   g23300(.A1(new_n25736_), .A2(new_n12880_), .B(new_n12779_), .ZN(new_n25737_));
  AOI21_X1   g23301(.A1(new_n25737_), .A2(new_n25732_), .B(new_n25727_), .ZN(new_n25738_));
  OR2_X2     g23302(.A1(new_n25738_), .A2(pi0789), .Z(new_n25739_));
  INV_X1     g23303(.I(new_n25625_), .ZN(new_n25740_));
  NOR2_X1    g23304(.A1(new_n25740_), .A2(pi0619), .ZN(new_n25741_));
  INV_X1     g23305(.I(new_n25741_), .ZN(new_n25742_));
  OAI21_X1   g23306(.A1(new_n25738_), .A2(new_n12793_), .B(new_n25742_), .ZN(new_n25743_));
  NAND2_X1   g23307(.A1(new_n13193_), .A2(new_n12791_), .ZN(new_n25744_));
  OAI21_X1   g23308(.A1(new_n25743_), .A2(new_n12791_), .B(new_n25744_), .ZN(new_n25745_));
  NAND2_X1   g23309(.A1(new_n25745_), .A2(pi0648), .ZN(new_n25746_));
  NAND2_X1   g23310(.A1(new_n13193_), .A2(pi1159), .ZN(new_n25747_));
  NOR2_X1    g23311(.A1(new_n25740_), .A2(new_n12793_), .ZN(new_n25748_));
  INV_X1     g23312(.I(new_n25748_), .ZN(new_n25749_));
  OAI21_X1   g23313(.A1(new_n25738_), .A2(pi0619), .B(new_n25749_), .ZN(new_n25750_));
  OAI21_X1   g23314(.A1(new_n25750_), .A2(pi1159), .B(new_n25747_), .ZN(new_n25751_));
  AOI21_X1   g23315(.A1(new_n25751_), .A2(new_n12895_), .B(new_n12796_), .ZN(new_n25752_));
  NAND2_X1   g23316(.A1(new_n25752_), .A2(new_n25746_), .ZN(new_n25753_));
  AND3_X2    g23317(.A1(new_n25753_), .A2(new_n12808_), .A3(new_n25739_), .Z(new_n25754_));
  NOR2_X1    g23318(.A1(new_n25754_), .A2(new_n15340_), .ZN(new_n25755_));
  AOI21_X1   g23319(.A1(new_n13192_), .A2(new_n12814_), .B(new_n12745_), .ZN(new_n25756_));
  INV_X1     g23320(.I(new_n25756_), .ZN(new_n25757_));
  AOI21_X1   g23321(.A1(new_n25628_), .A2(new_n12747_), .B(new_n12814_), .ZN(new_n25758_));
  NAND3_X1   g23322(.A1(new_n25753_), .A2(pi0626), .A3(new_n25739_), .ZN(new_n25759_));
  AOI21_X1   g23323(.A1(new_n25759_), .A2(new_n25758_), .B(new_n25757_), .ZN(new_n25760_));
  AOI21_X1   g23324(.A1(new_n13192_), .A2(pi0641), .B(pi1158), .ZN(new_n25761_));
  INV_X1     g23325(.I(new_n25761_), .ZN(new_n25762_));
  AOI21_X1   g23326(.A1(new_n25628_), .A2(pi0626), .B(pi0641), .ZN(new_n25763_));
  NAND3_X1   g23327(.A1(new_n25753_), .A2(new_n12747_), .A3(new_n25739_), .ZN(new_n25764_));
  AOI21_X1   g23328(.A1(new_n25764_), .A2(new_n25763_), .B(new_n25762_), .ZN(new_n25765_));
  OAI21_X1   g23329(.A1(new_n25760_), .A2(new_n25765_), .B(pi0788), .ZN(new_n25766_));
  AOI22_X1   g23330(.A1(new_n25766_), .A2(new_n25755_), .B1(pi0792), .B2(new_n25705_), .ZN(new_n25767_));
  NOR2_X1    g23331(.A1(new_n25767_), .A2(pi0207), .ZN(new_n25768_));
  NOR2_X1    g23332(.A1(new_n25610_), .A2(new_n12742_), .ZN(new_n25769_));
  INV_X1     g23333(.I(new_n25564_), .ZN(new_n25770_));
  NOR2_X1    g23334(.A1(new_n25770_), .A2(pi1156), .ZN(new_n25771_));
  NOR4_X1    g23335(.A1(new_n25771_), .A2(new_n12920_), .A3(pi0629), .A4(new_n25769_), .ZN(new_n25772_));
  NOR2_X1    g23336(.A1(new_n25610_), .A2(pi1156), .ZN(new_n25773_));
  NOR2_X1    g23337(.A1(new_n25770_), .A2(new_n12742_), .ZN(new_n25774_));
  NOR4_X1    g23338(.A1(new_n25774_), .A2(pi0628), .A3(new_n12919_), .A4(new_n25773_), .ZN(new_n25775_));
  OAI21_X1   g23339(.A1(new_n25772_), .A2(new_n25775_), .B(pi0792), .ZN(new_n25776_));
  NAND3_X1   g23340(.A1(new_n25563_), .A2(new_n12747_), .A3(pi0641), .ZN(new_n25777_));
  NAND2_X1   g23341(.A1(new_n25777_), .A2(new_n12745_), .ZN(new_n25778_));
  AOI21_X1   g23342(.A1(new_n25559_), .A2(new_n13521_), .B(new_n12841_), .ZN(new_n25779_));
  NAND2_X1   g23343(.A1(new_n25013_), .A2(pi0625), .ZN(new_n25780_));
  AOI21_X1   g23344(.A1(new_n25780_), .A2(new_n25779_), .B(new_n25654_), .ZN(new_n25781_));
  AOI21_X1   g23345(.A1(new_n25559_), .A2(pi0625), .B(pi1153), .ZN(new_n25782_));
  NAND2_X1   g23346(.A1(new_n25013_), .A2(new_n13521_), .ZN(new_n25783_));
  AOI21_X1   g23347(.A1(new_n25783_), .A2(new_n25782_), .B(new_n25659_), .ZN(new_n25784_));
  NOR3_X1    g23348(.A1(new_n25781_), .A2(new_n25784_), .A3(new_n12758_), .ZN(new_n25785_));
  NOR2_X1    g23349(.A1(new_n25013_), .A2(pi0778), .ZN(new_n25786_));
  NOR2_X1    g23350(.A1(new_n25785_), .A2(new_n25786_), .ZN(new_n25787_));
  NAND2_X1   g23351(.A1(new_n25787_), .A2(new_n12764_), .ZN(new_n25788_));
  NOR2_X1    g23352(.A1(new_n25560_), .A2(pi1155), .ZN(new_n25789_));
  AOI21_X1   g23353(.A1(new_n25789_), .A2(new_n12766_), .B(new_n13829_), .ZN(new_n25790_));
  OAI21_X1   g23354(.A1(new_n25787_), .A2(new_n12766_), .B(new_n25664_), .ZN(new_n25791_));
  NAND2_X1   g23355(.A1(new_n25791_), .A2(new_n25790_), .ZN(new_n25792_));
  NOR2_X1    g23356(.A1(new_n25560_), .A2(new_n12770_), .ZN(new_n25793_));
  AOI21_X1   g23357(.A1(new_n25793_), .A2(pi0609), .B(pi0660), .ZN(new_n25794_));
  OAI21_X1   g23358(.A1(new_n25787_), .A2(pi0609), .B(new_n25668_), .ZN(new_n25795_));
  AOI21_X1   g23359(.A1(new_n25795_), .A2(new_n25794_), .B(new_n12764_), .ZN(new_n25796_));
  NAND2_X1   g23360(.A1(new_n25796_), .A2(new_n25792_), .ZN(new_n25797_));
  NAND2_X1   g23361(.A1(new_n25797_), .A2(new_n25788_), .ZN(new_n25798_));
  NOR3_X1    g23362(.A1(new_n25562_), .A2(new_n12781_), .A3(new_n12785_), .ZN(new_n25799_));
  NOR3_X1    g23363(.A1(new_n25675_), .A2(pi0627), .A3(new_n25799_), .ZN(new_n25800_));
  AOI21_X1   g23364(.A1(new_n25561_), .A2(new_n15802_), .B(new_n12880_), .ZN(new_n25801_));
  OAI21_X1   g23365(.A1(new_n25798_), .A2(new_n12781_), .B(new_n25652_), .ZN(new_n25802_));
  AOI21_X1   g23366(.A1(new_n25802_), .A2(new_n25801_), .B(new_n25800_), .ZN(new_n25803_));
  AOI21_X1   g23367(.A1(new_n12781_), .A2(new_n12880_), .B(new_n12779_), .ZN(new_n25804_));
  OAI22_X1   g23368(.A1(new_n25803_), .A2(new_n12779_), .B1(new_n25798_), .B2(new_n25804_), .ZN(new_n25805_));
  NOR2_X1    g23369(.A1(new_n25681_), .A2(pi1159), .ZN(new_n25806_));
  NOR2_X1    g23370(.A1(new_n25562_), .A2(new_n15239_), .ZN(new_n25807_));
  NOR2_X1    g23371(.A1(new_n25807_), .A2(new_n12791_), .ZN(new_n25808_));
  NOR4_X1    g23372(.A1(new_n25808_), .A2(new_n25806_), .A3(new_n12793_), .A4(pi0648), .ZN(new_n25809_));
  NOR2_X1    g23373(.A1(new_n25681_), .A2(new_n12791_), .ZN(new_n25810_));
  NOR2_X1    g23374(.A1(new_n25807_), .A2(pi1159), .ZN(new_n25811_));
  NOR4_X1    g23375(.A1(new_n25811_), .A2(new_n25810_), .A3(pi0619), .A4(new_n12895_), .ZN(new_n25812_));
  NOR4_X1    g23376(.A1(new_n25809_), .A2(new_n25812_), .A3(new_n12796_), .A4(new_n17590_), .ZN(new_n25813_));
  NOR2_X1    g23377(.A1(new_n25805_), .A2(new_n25813_), .ZN(new_n25814_));
  NOR3_X1    g23378(.A1(new_n25809_), .A2(new_n25812_), .A3(new_n12796_), .ZN(new_n25815_));
  NOR2_X1    g23379(.A1(new_n25815_), .A2(new_n12796_), .ZN(new_n25816_));
  NOR2_X1    g23380(.A1(new_n25814_), .A2(new_n25816_), .ZN(new_n25817_));
  AOI21_X1   g23381(.A1(new_n25817_), .A2(new_n12747_), .B(new_n25686_), .ZN(new_n25818_));
  NOR2_X1    g23382(.A1(new_n25818_), .A2(new_n25778_), .ZN(new_n25819_));
  OAI21_X1   g23383(.A1(new_n25817_), .A2(new_n12747_), .B(new_n25689_), .ZN(new_n25820_));
  NAND3_X1   g23384(.A1(new_n25563_), .A2(pi0626), .A3(new_n12814_), .ZN(new_n25821_));
  NAND2_X1   g23385(.A1(new_n25821_), .A2(pi1158), .ZN(new_n25822_));
  AOI21_X1   g23386(.A1(new_n25820_), .A2(pi0641), .B(new_n25822_), .ZN(new_n25823_));
  OAI21_X1   g23387(.A1(new_n25823_), .A2(new_n25819_), .B(pi0788), .ZN(new_n25824_));
  AOI21_X1   g23388(.A1(new_n25817_), .A2(new_n12808_), .B(new_n15340_), .ZN(new_n25825_));
  NAND2_X1   g23389(.A1(new_n25824_), .A2(new_n25825_), .ZN(new_n25826_));
  NAND2_X1   g23390(.A1(new_n25826_), .A2(new_n25776_), .ZN(new_n25827_));
  AOI21_X1   g23391(.A1(new_n25827_), .A2(pi0207), .B(new_n25648_), .ZN(new_n25828_));
  AOI21_X1   g23392(.A1(new_n25702_), .A2(new_n12940_), .B(new_n25699_), .ZN(new_n25829_));
  NAND2_X1   g23393(.A1(new_n25598_), .A2(new_n19160_), .ZN(new_n25830_));
  AND2_X2    g23394(.A1(new_n25829_), .A2(new_n25830_), .Z(new_n25831_));
  NAND2_X1   g23395(.A1(new_n12815_), .A2(new_n12747_), .ZN(new_n25832_));
  OAI21_X1   g23396(.A1(new_n12747_), .A2(new_n12813_), .B(new_n25832_), .ZN(new_n25833_));
  OAI21_X1   g23397(.A1(new_n13193_), .A2(new_n12814_), .B(new_n12748_), .ZN(new_n25834_));
  NOR2_X1    g23398(.A1(new_n25628_), .A2(pi0641), .ZN(new_n25835_));
  OAI21_X1   g23399(.A1(new_n13193_), .A2(pi0641), .B(new_n12746_), .ZN(new_n25836_));
  NOR2_X1    g23400(.A1(new_n25628_), .A2(new_n12814_), .ZN(new_n25837_));
  OAI22_X1   g23401(.A1(new_n25834_), .A2(new_n25835_), .B1(new_n25837_), .B2(new_n25836_), .ZN(new_n25838_));
  AOI21_X1   g23402(.A1(new_n25596_), .A2(new_n25833_), .B(new_n25838_), .ZN(new_n25839_));
  OAI21_X1   g23403(.A1(new_n25839_), .A2(new_n12808_), .B(new_n15824_), .ZN(new_n25840_));
  NOR2_X1    g23404(.A1(new_n25593_), .A2(new_n12895_), .ZN(new_n25841_));
  NOR2_X1    g23405(.A1(new_n25614_), .A2(new_n13521_), .ZN(new_n25842_));
  OAI21_X1   g23406(.A1(new_n25842_), .A2(new_n14199_), .B(pi1153), .ZN(new_n25843_));
  NAND2_X1   g23407(.A1(new_n25568_), .A2(pi0625), .ZN(new_n25844_));
  NAND2_X1   g23408(.A1(new_n15111_), .A2(new_n2609_), .ZN(new_n25845_));
  NAND2_X1   g23409(.A1(new_n25845_), .A2(new_n13521_), .ZN(new_n25846_));
  NAND2_X1   g23410(.A1(new_n25846_), .A2(new_n25844_), .ZN(new_n25847_));
  NAND2_X1   g23411(.A1(new_n25847_), .A2(new_n12841_), .ZN(new_n25848_));
  NAND3_X1   g23412(.A1(new_n25843_), .A2(new_n25848_), .A3(new_n13560_), .ZN(new_n25849_));
  NAND2_X1   g23413(.A1(new_n25568_), .A2(new_n13521_), .ZN(new_n25850_));
  NAND2_X1   g23414(.A1(new_n25845_), .A2(pi0625), .ZN(new_n25851_));
  NAND2_X1   g23415(.A1(new_n25851_), .A2(new_n25850_), .ZN(new_n25852_));
  NAND2_X1   g23416(.A1(new_n25852_), .A2(pi1153), .ZN(new_n25853_));
  NAND3_X1   g23417(.A1(new_n25616_), .A2(new_n25853_), .A3(pi0608), .ZN(new_n25854_));
  NAND3_X1   g23418(.A1(new_n25849_), .A2(new_n25854_), .A3(pi0778), .ZN(new_n25855_));
  NAND2_X1   g23419(.A1(new_n25845_), .A2(new_n12758_), .ZN(new_n25856_));
  NAND2_X1   g23420(.A1(new_n25855_), .A2(new_n25856_), .ZN(new_n25857_));
  NAND2_X1   g23421(.A1(new_n25857_), .A2(new_n12764_), .ZN(new_n25858_));
  INV_X1     g23422(.I(new_n25574_), .ZN(new_n25859_));
  NAND2_X1   g23423(.A1(new_n25857_), .A2(pi0609), .ZN(new_n25860_));
  AOI21_X1   g23424(.A1(new_n25860_), .A2(new_n25706_), .B(new_n12770_), .ZN(new_n25861_));
  NOR3_X1    g23425(.A1(new_n25861_), .A2(new_n13829_), .A3(new_n25859_), .ZN(new_n25862_));
  NAND2_X1   g23426(.A1(new_n25857_), .A2(new_n12766_), .ZN(new_n25863_));
  NAND2_X1   g23427(.A1(new_n25863_), .A2(new_n25721_), .ZN(new_n25864_));
  NAND2_X1   g23428(.A1(new_n25575_), .A2(pi1155), .ZN(new_n25865_));
  NAND2_X1   g23429(.A1(new_n25865_), .A2(new_n13829_), .ZN(new_n25866_));
  AOI21_X1   g23430(.A1(new_n25864_), .A2(new_n12770_), .B(new_n25866_), .ZN(new_n25867_));
  OR3_X2     g23431(.A1(new_n25862_), .A2(new_n12764_), .A3(new_n25867_), .Z(new_n25868_));
  NAND2_X1   g23432(.A1(new_n25868_), .A2(new_n25858_), .ZN(new_n25869_));
  NAND2_X1   g23433(.A1(new_n25869_), .A2(new_n12781_), .ZN(new_n25870_));
  AOI21_X1   g23434(.A1(new_n25870_), .A2(new_n25734_), .B(pi1154), .ZN(new_n25871_));
  NOR3_X1    g23435(.A1(new_n25871_), .A2(pi0627), .A3(new_n25581_), .ZN(new_n25872_));
  NAND2_X1   g23436(.A1(new_n25869_), .A2(pi0618), .ZN(new_n25873_));
  NAND2_X1   g23437(.A1(new_n25873_), .A2(new_n25728_), .ZN(new_n25874_));
  OAI21_X1   g23438(.A1(new_n25583_), .A2(pi1154), .B(pi0627), .ZN(new_n25875_));
  AOI21_X1   g23439(.A1(new_n25874_), .A2(pi1154), .B(new_n25875_), .ZN(new_n25876_));
  OR3_X2     g23440(.A1(new_n25872_), .A2(new_n12779_), .A3(new_n25876_), .Z(new_n25877_));
  NAND2_X1   g23441(.A1(new_n25869_), .A2(new_n12779_), .ZN(new_n25878_));
  NAND2_X1   g23442(.A1(new_n25877_), .A2(new_n25878_), .ZN(new_n25879_));
  AOI21_X1   g23443(.A1(new_n25879_), .A2(pi0619), .B(new_n25741_), .ZN(new_n25880_));
  OAI21_X1   g23444(.A1(new_n25880_), .A2(new_n12791_), .B(new_n25841_), .ZN(new_n25881_));
  AOI21_X1   g23445(.A1(new_n25589_), .A2(pi1159), .B(pi0648), .ZN(new_n25882_));
  AOI21_X1   g23446(.A1(new_n25877_), .A2(new_n25878_), .B(pi0619), .ZN(new_n25883_));
  OAI21_X1   g23447(.A1(new_n25883_), .A2(new_n25748_), .B(new_n12791_), .ZN(new_n25884_));
  AOI21_X1   g23448(.A1(new_n25884_), .A2(new_n25882_), .B(new_n12796_), .ZN(new_n25885_));
  NAND2_X1   g23449(.A1(new_n25879_), .A2(new_n12796_), .ZN(new_n25886_));
  NAND2_X1   g23450(.A1(new_n25886_), .A2(new_n12819_), .ZN(new_n25887_));
  AOI21_X1   g23451(.A1(new_n25885_), .A2(new_n25881_), .B(new_n25887_), .ZN(new_n25888_));
  OAI22_X1   g23452(.A1(new_n25888_), .A2(new_n25840_), .B1(new_n12937_), .B2(new_n25831_), .ZN(new_n25889_));
  NAND2_X1   g23453(.A1(new_n25889_), .A2(new_n8521_), .ZN(new_n25890_));
  AOI21_X1   g23454(.A1(new_n25890_), .A2(new_n25828_), .B(new_n25607_), .ZN(new_n25891_));
  OAI21_X1   g23455(.A1(new_n25768_), .A2(new_n25696_), .B(new_n25891_), .ZN(new_n25892_));
  AOI22_X1   g23456(.A1(new_n25892_), .A2(new_n25647_), .B1(pi0787), .B2(new_n25646_), .ZN(new_n25893_));
  OAI21_X1   g23457(.A1(new_n25603_), .A2(new_n12975_), .B(pi0715), .ZN(new_n25894_));
  NOR2_X1    g23458(.A1(new_n25603_), .A2(new_n12985_), .ZN(new_n25895_));
  AOI21_X1   g23459(.A1(new_n25606_), .A2(new_n12985_), .B(new_n25895_), .ZN(new_n25896_));
  NOR2_X1    g23460(.A1(new_n25896_), .A2(pi0644), .ZN(new_n25897_));
  OAI21_X1   g23461(.A1(new_n25897_), .A2(new_n25894_), .B(new_n12739_), .ZN(new_n25898_));
  NOR2_X1    g23462(.A1(new_n25639_), .A2(new_n12972_), .ZN(new_n25899_));
  AOI22_X1   g23463(.A1(new_n25899_), .A2(new_n25643_), .B1(new_n12972_), .B2(new_n25640_), .ZN(new_n25900_));
  NOR2_X1    g23464(.A1(new_n25900_), .A2(new_n12975_), .ZN(new_n25901_));
  NOR2_X1    g23465(.A1(new_n25901_), .A2(pi0715), .ZN(new_n25902_));
  NAND2_X1   g23466(.A1(new_n25893_), .A2(new_n12975_), .ZN(new_n25903_));
  AOI21_X1   g23467(.A1(new_n25903_), .A2(new_n25902_), .B(new_n25898_), .ZN(new_n25904_));
  OAI21_X1   g23468(.A1(new_n25603_), .A2(pi0644), .B(new_n12740_), .ZN(new_n25905_));
  NOR2_X1    g23469(.A1(new_n25896_), .A2(new_n12975_), .ZN(new_n25906_));
  OAI21_X1   g23470(.A1(new_n25906_), .A2(new_n25905_), .B(pi1160), .ZN(new_n25907_));
  OAI21_X1   g23471(.A1(new_n25900_), .A2(pi0644), .B(pi0715), .ZN(new_n25908_));
  AOI21_X1   g23472(.A1(new_n25893_), .A2(pi0644), .B(new_n25908_), .ZN(new_n25909_));
  OAI21_X1   g23473(.A1(new_n25909_), .A2(new_n25907_), .B(pi0790), .ZN(new_n25910_));
  OAI22_X1   g23474(.A1(new_n25910_), .A2(new_n25904_), .B1(pi0790), .B2(new_n25893_), .ZN(new_n25911_));
  NAND2_X1   g23475(.A1(po1038), .A2(new_n8521_), .ZN(new_n25912_));
  OAI21_X1   g23476(.A1(new_n25911_), .A2(po1038), .B(new_n25912_), .ZN(po0364));
  NAND2_X1   g23477(.A1(new_n25565_), .A2(pi0208), .ZN(new_n25914_));
  OAI21_X1   g23478(.A1(new_n25600_), .A2(pi0208), .B(new_n25914_), .ZN(new_n25915_));
  NOR2_X1    g23479(.A1(new_n13193_), .A2(pi0208), .ZN(new_n25916_));
  INV_X1     g23480(.I(new_n25916_), .ZN(new_n25917_));
  NOR2_X1    g23481(.A1(new_n25917_), .A2(pi0607), .ZN(new_n25918_));
  AOI21_X1   g23482(.A1(new_n25915_), .A2(pi0607), .B(new_n25918_), .ZN(new_n25919_));
  INV_X1     g23483(.I(new_n25919_), .ZN(new_n25920_));
  INV_X1     g23484(.I(pi0638), .ZN(new_n25921_));
  NAND2_X1   g23485(.A1(new_n25612_), .A2(pi0208), .ZN(new_n25922_));
  NAND2_X1   g23486(.A1(new_n25632_), .A2(new_n8522_), .ZN(new_n25923_));
  AOI21_X1   g23487(.A1(new_n25923_), .A2(new_n25922_), .B(new_n25921_), .ZN(new_n25924_));
  NOR2_X1    g23488(.A1(new_n25917_), .A2(pi0638), .ZN(new_n25925_));
  NOR2_X1    g23489(.A1(new_n25924_), .A2(new_n25925_), .ZN(new_n25926_));
  NAND2_X1   g23490(.A1(new_n25926_), .A2(new_n12741_), .ZN(new_n25927_));
  NAND2_X1   g23491(.A1(new_n25917_), .A2(pi0647), .ZN(new_n25928_));
  AOI21_X1   g23492(.A1(new_n25927_), .A2(new_n25928_), .B(pi1157), .ZN(new_n25929_));
  INV_X1     g23493(.I(new_n25926_), .ZN(new_n25930_));
  NOR2_X1    g23494(.A1(new_n25930_), .A2(new_n12741_), .ZN(new_n25931_));
  NOR2_X1    g23495(.A1(new_n25916_), .A2(pi0647), .ZN(new_n25932_));
  OAI21_X1   g23496(.A1(new_n25931_), .A2(new_n25932_), .B(pi1157), .ZN(new_n25933_));
  NAND2_X1   g23497(.A1(new_n25933_), .A2(new_n12981_), .ZN(new_n25934_));
  OAI21_X1   g23498(.A1(new_n12981_), .A2(new_n25929_), .B(new_n25934_), .ZN(new_n25935_));
  OAI21_X1   g23499(.A1(new_n17212_), .A2(new_n25920_), .B(new_n25935_), .ZN(new_n25936_));
  AOI21_X1   g23500(.A1(new_n25920_), .A2(new_n25921_), .B(new_n15341_), .ZN(new_n25937_));
  INV_X1     g23501(.I(pi0607), .ZN(new_n25938_));
  OAI21_X1   g23502(.A1(new_n25695_), .A2(new_n8522_), .B(new_n25938_), .ZN(new_n25939_));
  NOR2_X1    g23503(.A1(new_n25767_), .A2(pi0208), .ZN(new_n25940_));
  AOI21_X1   g23504(.A1(new_n25827_), .A2(pi0208), .B(new_n25938_), .ZN(new_n25941_));
  NAND2_X1   g23505(.A1(new_n25889_), .A2(new_n8522_), .ZN(new_n25942_));
  AOI21_X1   g23506(.A1(new_n25942_), .A2(new_n25941_), .B(new_n25921_), .ZN(new_n25943_));
  OAI21_X1   g23507(.A1(new_n25940_), .A2(new_n25939_), .B(new_n25943_), .ZN(new_n25944_));
  AOI22_X1   g23508(.A1(new_n25944_), .A2(new_n25937_), .B1(pi0787), .B2(new_n25936_), .ZN(new_n25945_));
  OAI21_X1   g23509(.A1(new_n25917_), .A2(new_n12975_), .B(pi0715), .ZN(new_n25946_));
  NOR2_X1    g23510(.A1(new_n25917_), .A2(new_n12985_), .ZN(new_n25947_));
  AOI21_X1   g23511(.A1(new_n25920_), .A2(new_n12985_), .B(new_n25947_), .ZN(new_n25948_));
  NOR2_X1    g23512(.A1(new_n25948_), .A2(pi0644), .ZN(new_n25949_));
  OAI21_X1   g23513(.A1(new_n25949_), .A2(new_n25946_), .B(new_n12739_), .ZN(new_n25950_));
  NOR2_X1    g23514(.A1(new_n25929_), .A2(new_n12972_), .ZN(new_n25951_));
  AOI22_X1   g23515(.A1(new_n25951_), .A2(new_n25933_), .B1(new_n12972_), .B2(new_n25930_), .ZN(new_n25952_));
  NOR2_X1    g23516(.A1(new_n25952_), .A2(new_n12975_), .ZN(new_n25953_));
  NOR2_X1    g23517(.A1(new_n25953_), .A2(pi0715), .ZN(new_n25954_));
  NAND2_X1   g23518(.A1(new_n25945_), .A2(new_n12975_), .ZN(new_n25955_));
  AOI21_X1   g23519(.A1(new_n25955_), .A2(new_n25954_), .B(new_n25950_), .ZN(new_n25956_));
  OAI21_X1   g23520(.A1(new_n25917_), .A2(pi0644), .B(new_n12740_), .ZN(new_n25957_));
  NOR2_X1    g23521(.A1(new_n25948_), .A2(new_n12975_), .ZN(new_n25958_));
  OAI21_X1   g23522(.A1(new_n25958_), .A2(new_n25957_), .B(pi1160), .ZN(new_n25959_));
  OAI21_X1   g23523(.A1(new_n25952_), .A2(pi0644), .B(pi0715), .ZN(new_n25960_));
  AOI21_X1   g23524(.A1(new_n25945_), .A2(pi0644), .B(new_n25960_), .ZN(new_n25961_));
  OAI21_X1   g23525(.A1(new_n25961_), .A2(new_n25959_), .B(pi0790), .ZN(new_n25962_));
  OAI22_X1   g23526(.A1(new_n25962_), .A2(new_n25956_), .B1(pi0790), .B2(new_n25945_), .ZN(new_n25963_));
  NAND2_X1   g23527(.A1(po1038), .A2(new_n8522_), .ZN(new_n25964_));
  OAI21_X1   g23528(.A1(new_n25963_), .A2(po1038), .B(new_n25964_), .ZN(po0365));
  INV_X1     g23529(.I(pi0639), .ZN(new_n25966_));
  NAND2_X1   g23530(.A1(new_n12975_), .A2(pi1160), .ZN(new_n25967_));
  NAND2_X1   g23531(.A1(new_n12739_), .A2(pi0644), .ZN(new_n25968_));
  AOI21_X1   g23532(.A1(new_n25967_), .A2(new_n25968_), .B(new_n13000_), .ZN(new_n25969_));
  NOR4_X1    g23533(.A1(new_n25564_), .A2(po1038), .A3(new_n17612_), .A4(new_n25969_), .ZN(new_n25970_));
  NAND2_X1   g23534(.A1(new_n25970_), .A2(pi0622), .ZN(new_n25971_));
  NAND2_X1   g23535(.A1(new_n25971_), .A2(new_n25966_), .ZN(new_n25972_));
  INV_X1     g23536(.I(pi0622), .ZN(new_n25973_));
  NAND2_X1   g23537(.A1(new_n12984_), .A2(new_n14299_), .ZN(new_n25974_));
  OAI22_X1   g23538(.A1(new_n25695_), .A2(new_n15341_), .B1(new_n25611_), .B2(new_n25974_), .ZN(new_n25975_));
  NOR2_X1    g23539(.A1(new_n25975_), .A2(pi0790), .ZN(new_n25976_));
  NOR2_X1    g23540(.A1(new_n25976_), .A2(po1038), .ZN(new_n25977_));
  NOR2_X1    g23541(.A1(new_n25611_), .A2(new_n14300_), .ZN(new_n25978_));
  INV_X1     g23542(.I(new_n25978_), .ZN(new_n25979_));
  AOI21_X1   g23543(.A1(new_n25979_), .A2(pi0644), .B(pi0715), .ZN(new_n25980_));
  OAI21_X1   g23544(.A1(new_n25975_), .A2(pi0644), .B(new_n25980_), .ZN(new_n25981_));
  NOR2_X1    g23545(.A1(new_n25981_), .A2(pi1160), .ZN(new_n25982_));
  AOI21_X1   g23546(.A1(new_n25979_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n25983_));
  INV_X1     g23547(.I(new_n25983_), .ZN(new_n25984_));
  OAI21_X1   g23548(.A1(new_n25975_), .A2(new_n12975_), .B(pi1160), .ZN(new_n25985_));
  OAI21_X1   g23549(.A1(new_n25985_), .A2(new_n25984_), .B(pi0790), .ZN(new_n25986_));
  OAI21_X1   g23550(.A1(new_n25986_), .A2(new_n25982_), .B(new_n25977_), .ZN(new_n25987_));
  NAND2_X1   g23551(.A1(new_n25987_), .A2(new_n25973_), .ZN(new_n25988_));
  INV_X1     g23552(.I(new_n25827_), .ZN(new_n25989_));
  NOR2_X1    g23553(.A1(new_n25565_), .A2(pi0647), .ZN(new_n25990_));
  AOI21_X1   g23554(.A1(new_n25989_), .A2(pi0647), .B(new_n25990_), .ZN(new_n25991_));
  NAND2_X1   g23555(.A1(new_n25612_), .A2(new_n12741_), .ZN(new_n25992_));
  AOI21_X1   g23556(.A1(new_n25992_), .A2(new_n12965_), .B(new_n12981_), .ZN(new_n25993_));
  OAI21_X1   g23557(.A1(new_n25991_), .A2(new_n12965_), .B(new_n25993_), .ZN(new_n25994_));
  NOR2_X1    g23558(.A1(new_n25565_), .A2(new_n12741_), .ZN(new_n25995_));
  AOI21_X1   g23559(.A1(new_n25989_), .A2(new_n12741_), .B(new_n25995_), .ZN(new_n25996_));
  NAND2_X1   g23560(.A1(new_n25612_), .A2(pi0647), .ZN(new_n25997_));
  AOI21_X1   g23561(.A1(new_n25997_), .A2(pi1157), .B(pi0630), .ZN(new_n25998_));
  OAI21_X1   g23562(.A1(new_n25996_), .A2(pi1157), .B(new_n25998_), .ZN(new_n25999_));
  NAND3_X1   g23563(.A1(new_n25994_), .A2(new_n25999_), .A3(pi0787), .ZN(new_n26000_));
  OAI21_X1   g23564(.A1(pi0787), .A2(new_n25827_), .B(new_n26000_), .ZN(new_n26001_));
  AOI21_X1   g23565(.A1(new_n26001_), .A2(new_n13000_), .B(po1038), .ZN(new_n26002_));
  NOR2_X1    g23566(.A1(new_n25564_), .A2(new_n17612_), .ZN(new_n26003_));
  NAND3_X1   g23567(.A1(new_n26003_), .A2(pi0644), .A3(new_n12740_), .ZN(new_n26004_));
  NAND2_X1   g23568(.A1(new_n26004_), .A2(pi1160), .ZN(new_n26005_));
  NAND2_X1   g23569(.A1(new_n26001_), .A2(pi0644), .ZN(new_n26006_));
  AOI21_X1   g23570(.A1(new_n26006_), .A2(new_n25983_), .B(new_n26005_), .ZN(new_n26007_));
  NAND3_X1   g23571(.A1(new_n26003_), .A2(new_n12975_), .A3(pi0715), .ZN(new_n26008_));
  NAND2_X1   g23572(.A1(new_n26008_), .A2(new_n12739_), .ZN(new_n26009_));
  NAND2_X1   g23573(.A1(new_n26001_), .A2(new_n12975_), .ZN(new_n26010_));
  AOI21_X1   g23574(.A1(new_n26010_), .A2(new_n25980_), .B(new_n26009_), .ZN(new_n26011_));
  OAI21_X1   g23575(.A1(new_n26007_), .A2(new_n26011_), .B(pi0790), .ZN(new_n26012_));
  NAND2_X1   g23576(.A1(new_n26012_), .A2(new_n26002_), .ZN(new_n26013_));
  NAND3_X1   g23577(.A1(new_n26013_), .A2(pi0622), .A3(pi0639), .ZN(new_n26014_));
  NAND4_X1   g23578(.A1(new_n26014_), .A2(pi0209), .A3(new_n25972_), .A4(new_n25988_), .ZN(new_n26015_));
  NOR2_X1    g23579(.A1(new_n13193_), .A2(pi0647), .ZN(new_n26016_));
  AOI21_X1   g23580(.A1(new_n25632_), .A2(pi0647), .B(new_n26016_), .ZN(new_n26017_));
  NOR2_X1    g23581(.A1(new_n26017_), .A2(pi0630), .ZN(new_n26018_));
  NOR2_X1    g23582(.A1(new_n13192_), .A2(new_n12741_), .ZN(new_n26019_));
  INV_X1     g23583(.I(new_n26019_), .ZN(new_n26020_));
  OAI21_X1   g23584(.A1(new_n25632_), .A2(pi0647), .B(new_n26020_), .ZN(new_n26021_));
  INV_X1     g23585(.I(new_n26021_), .ZN(new_n26022_));
  AOI22_X1   g23586(.A1(new_n26018_), .A2(pi1157), .B1(new_n26022_), .B2(new_n12982_), .ZN(new_n26023_));
  OAI21_X1   g23587(.A1(new_n17212_), .A2(new_n25600_), .B(new_n26023_), .ZN(new_n26024_));
  AOI22_X1   g23588(.A1(new_n25889_), .A2(new_n15693_), .B1(pi0787), .B2(new_n26024_), .ZN(new_n26025_));
  OAI21_X1   g23589(.A1(new_n26025_), .A2(pi0790), .B(new_n6643_), .ZN(new_n26026_));
  NOR2_X1    g23590(.A1(new_n13192_), .A2(new_n12985_), .ZN(new_n26027_));
  AOI21_X1   g23591(.A1(new_n25600_), .A2(new_n12985_), .B(new_n26027_), .ZN(new_n26028_));
  NAND2_X1   g23592(.A1(new_n13193_), .A2(new_n12975_), .ZN(new_n26029_));
  OAI21_X1   g23593(.A1(new_n26028_), .A2(new_n12975_), .B(new_n26029_), .ZN(new_n26030_));
  AOI21_X1   g23594(.A1(new_n26030_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n26031_));
  NOR2_X1    g23595(.A1(new_n25632_), .A2(new_n14300_), .ZN(new_n26032_));
  AOI21_X1   g23596(.A1(new_n13193_), .A2(new_n14300_), .B(new_n26032_), .ZN(new_n26033_));
  AOI21_X1   g23597(.A1(new_n26033_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n26034_));
  OAI21_X1   g23598(.A1(new_n26025_), .A2(new_n12975_), .B(new_n26034_), .ZN(new_n26035_));
  NAND2_X1   g23599(.A1(new_n13193_), .A2(pi0644), .ZN(new_n26036_));
  OAI21_X1   g23600(.A1(new_n26028_), .A2(pi0644), .B(new_n26036_), .ZN(new_n26037_));
  AOI21_X1   g23601(.A1(new_n26037_), .A2(pi0715), .B(pi1160), .ZN(new_n26038_));
  AOI21_X1   g23602(.A1(new_n26033_), .A2(pi0644), .B(pi0715), .ZN(new_n26039_));
  OAI21_X1   g23603(.A1(new_n26025_), .A2(pi0644), .B(new_n26039_), .ZN(new_n26040_));
  AOI22_X1   g23604(.A1(new_n26031_), .A2(new_n26035_), .B1(new_n26040_), .B2(new_n26038_), .ZN(new_n26041_));
  NOR2_X1    g23605(.A1(new_n26041_), .A2(new_n13000_), .ZN(new_n26042_));
  OAI21_X1   g23606(.A1(new_n26042_), .A2(new_n26026_), .B(pi0639), .ZN(new_n26043_));
  NOR2_X1    g23607(.A1(new_n26037_), .A2(pi1160), .ZN(new_n26044_));
  NOR2_X1    g23608(.A1(new_n26030_), .A2(new_n12739_), .ZN(new_n26045_));
  OAI21_X1   g23609(.A1(new_n26044_), .A2(new_n26045_), .B(pi0790), .ZN(new_n26046_));
  NAND2_X1   g23610(.A1(new_n26028_), .A2(new_n13000_), .ZN(new_n26047_));
  NAND3_X1   g23611(.A1(new_n26046_), .A2(new_n6643_), .A3(new_n26047_), .ZN(new_n26048_));
  NAND2_X1   g23612(.A1(new_n26048_), .A2(new_n25966_), .ZN(new_n26049_));
  AOI21_X1   g23613(.A1(new_n26043_), .A2(new_n26049_), .B(new_n25973_), .ZN(new_n26050_));
  OAI22_X1   g23614(.A1(new_n26021_), .A2(new_n15730_), .B1(new_n13193_), .B2(new_n15606_), .ZN(new_n26051_));
  INV_X1     g23615(.I(new_n26051_), .ZN(new_n26052_));
  OAI21_X1   g23616(.A1(new_n26018_), .A2(new_n26016_), .B(pi1157), .ZN(new_n26053_));
  AOI21_X1   g23617(.A1(new_n26052_), .A2(new_n26053_), .B(new_n12972_), .ZN(new_n26054_));
  INV_X1     g23618(.I(new_n26054_), .ZN(new_n26055_));
  OAI21_X1   g23619(.A1(new_n25767_), .A2(new_n15341_), .B(new_n26055_), .ZN(new_n26056_));
  NAND2_X1   g23620(.A1(new_n26056_), .A2(new_n13000_), .ZN(new_n26057_));
  NAND2_X1   g23621(.A1(new_n26057_), .A2(new_n6643_), .ZN(new_n26058_));
  OAI21_X1   g23622(.A1(new_n13192_), .A2(pi0715), .B(pi1160), .ZN(new_n26059_));
  INV_X1     g23623(.I(new_n26034_), .ZN(new_n26060_));
  AOI21_X1   g23624(.A1(new_n26056_), .A2(pi0644), .B(new_n26060_), .ZN(new_n26061_));
  OAI21_X1   g23625(.A1(new_n13192_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n26062_));
  INV_X1     g23626(.I(new_n26039_), .ZN(new_n26063_));
  AOI21_X1   g23627(.A1(new_n26056_), .A2(new_n12975_), .B(new_n26063_), .ZN(new_n26064_));
  OAI22_X1   g23628(.A1(new_n26059_), .A2(new_n26061_), .B1(new_n26064_), .B2(new_n26062_), .ZN(new_n26065_));
  AOI21_X1   g23629(.A1(new_n26065_), .A2(pi0790), .B(new_n26058_), .ZN(new_n26066_));
  OAI21_X1   g23630(.A1(new_n13395_), .A2(new_n8265_), .B(new_n25966_), .ZN(new_n26067_));
  OAI21_X1   g23631(.A1(new_n26066_), .A2(new_n25966_), .B(new_n26067_), .ZN(new_n26068_));
  AOI21_X1   g23632(.A1(new_n26068_), .A2(new_n25973_), .B(new_n26050_), .ZN(new_n26069_));
  OAI21_X1   g23633(.A1(new_n26069_), .A2(pi0209), .B(new_n26015_), .ZN(po0366));
  NAND2_X1   g23634(.A1(new_n13397_), .A2(new_n2709_), .ZN(new_n26071_));
  AOI22_X1   g23635(.A1(new_n15936_), .A2(pi0634), .B1(pi0633), .B2(pi0947), .ZN(new_n26072_));
  NAND2_X1   g23636(.A1(new_n13344_), .A2(new_n26072_), .ZN(new_n26073_));
  AOI21_X1   g23637(.A1(new_n26071_), .A2(new_n26073_), .B(new_n3265_), .ZN(new_n26074_));
  INV_X1     g23638(.I(new_n26072_), .ZN(new_n26075_));
  NAND3_X1   g23639(.A1(new_n13038_), .A2(new_n13039_), .A3(new_n2709_), .ZN(new_n26076_));
  AOI21_X1   g23640(.A1(new_n26076_), .A2(new_n26075_), .B(new_n2628_), .ZN(new_n26077_));
  OAI21_X1   g23641(.A1(new_n2709_), .A2(new_n13054_), .B(new_n26077_), .ZN(new_n26078_));
  NOR2_X1    g23642(.A1(new_n15945_), .A2(pi0210), .ZN(new_n26079_));
  NOR2_X1    g23643(.A1(new_n13058_), .A2(new_n26075_), .ZN(new_n26080_));
  OAI21_X1   g23644(.A1(new_n26079_), .A2(new_n26080_), .B(new_n2628_), .ZN(new_n26081_));
  NAND3_X1   g23645(.A1(new_n26081_), .A2(new_n2627_), .A3(new_n26078_), .ZN(new_n26082_));
  NAND2_X1   g23646(.A1(new_n26082_), .A2(new_n3265_), .ZN(new_n26083_));
  NOR2_X1    g23647(.A1(new_n13098_), .A2(pi0210), .ZN(new_n26084_));
  AOI21_X1   g23648(.A1(new_n24611_), .A2(new_n13098_), .B(new_n26084_), .ZN(new_n26085_));
  INV_X1     g23649(.I(new_n26085_), .ZN(new_n26086_));
  NOR2_X1    g23650(.A1(new_n26086_), .A2(new_n5427_), .ZN(new_n26087_));
  INV_X1     g23651(.I(new_n26087_), .ZN(new_n26088_));
  NOR2_X1    g23652(.A1(new_n13082_), .A2(pi0210), .ZN(new_n26089_));
  INV_X1     g23653(.I(new_n26089_), .ZN(new_n26090_));
  OAI21_X1   g23654(.A1(pi0633), .A2(new_n13303_), .B(new_n26090_), .ZN(new_n26091_));
  OAI21_X1   g23655(.A1(new_n26091_), .A2(new_n5413_), .B(new_n26088_), .ZN(new_n26092_));
  NAND2_X1   g23656(.A1(new_n26092_), .A2(pi0947), .ZN(new_n26093_));
  AOI21_X1   g23657(.A1(new_n24493_), .A2(new_n13098_), .B(new_n26084_), .ZN(new_n26094_));
  AND2_X2    g23658(.A1(new_n26094_), .A2(new_n5413_), .Z(new_n26095_));
  AOI21_X1   g23659(.A1(new_n24493_), .A2(new_n13082_), .B(new_n26089_), .ZN(new_n26096_));
  AOI21_X1   g23660(.A1(new_n26096_), .A2(new_n5427_), .B(new_n26095_), .ZN(new_n26097_));
  NOR2_X1    g23661(.A1(new_n26097_), .A2(new_n5473_), .ZN(new_n26098_));
  NOR2_X1    g23662(.A1(new_n24475_), .A2(new_n2709_), .ZN(new_n26099_));
  OAI21_X1   g23663(.A1(new_n26099_), .A2(new_n5419_), .B(new_n5473_), .ZN(new_n26100_));
  AOI21_X1   g23664(.A1(new_n13308_), .A2(pi0210), .B(new_n5418_), .ZN(new_n26101_));
  NOR2_X1    g23665(.A1(new_n26100_), .A2(new_n26101_), .ZN(new_n26102_));
  OAI21_X1   g23666(.A1(new_n26102_), .A2(new_n26098_), .B(new_n5692_), .ZN(new_n26103_));
  NAND3_X1   g23667(.A1(new_n26103_), .A2(new_n3304_), .A3(new_n26093_), .ZN(new_n26104_));
  AOI21_X1   g23668(.A1(new_n13098_), .A2(new_n26072_), .B(new_n26084_), .ZN(new_n26105_));
  NOR2_X1    g23669(.A1(new_n26105_), .A2(new_n3304_), .ZN(new_n26106_));
  NOR2_X1    g23670(.A1(new_n26106_), .A2(pi0215), .ZN(new_n26107_));
  NOR2_X1    g23671(.A1(new_n13274_), .A2(pi0210), .ZN(new_n26108_));
  AOI21_X1   g23672(.A1(new_n24611_), .A2(new_n13274_), .B(new_n26108_), .ZN(new_n26109_));
  NAND2_X1   g23673(.A1(new_n26109_), .A2(new_n5427_), .ZN(new_n26110_));
  AOI21_X1   g23674(.A1(new_n26110_), .A2(new_n26088_), .B(new_n5692_), .ZN(new_n26111_));
  INV_X1     g23675(.I(new_n26108_), .ZN(new_n26112_));
  OAI21_X1   g23676(.A1(pi0634), .A2(new_n13149_), .B(new_n26112_), .ZN(new_n26113_));
  NOR2_X1    g23677(.A1(new_n26113_), .A2(new_n5413_), .ZN(new_n26114_));
  OAI21_X1   g23678(.A1(new_n26114_), .A2(new_n26095_), .B(pi0907), .ZN(new_n26115_));
  INV_X1     g23679(.I(new_n13150_), .ZN(new_n26116_));
  AOI21_X1   g23680(.A1(new_n26116_), .A2(po1101), .B(new_n24474_), .ZN(new_n26117_));
  NOR2_X1    g23681(.A1(new_n26117_), .A2(new_n2709_), .ZN(new_n26118_));
  NAND2_X1   g23682(.A1(new_n13098_), .A2(new_n5413_), .ZN(new_n26119_));
  NAND3_X1   g23683(.A1(new_n13149_), .A2(new_n26119_), .A3(pi0210), .ZN(new_n26120_));
  NOR2_X1    g23684(.A1(new_n26120_), .A2(new_n5418_), .ZN(new_n26121_));
  AOI21_X1   g23685(.A1(new_n26118_), .A2(new_n5418_), .B(new_n26121_), .ZN(new_n26122_));
  OAI21_X1   g23686(.A1(new_n26122_), .A2(pi0907), .B(new_n26115_), .ZN(new_n26123_));
  AOI21_X1   g23687(.A1(new_n26123_), .A2(new_n5692_), .B(new_n26111_), .ZN(new_n26124_));
  OAI21_X1   g23688(.A1(new_n26124_), .A2(new_n2436_), .B(pi0299), .ZN(new_n26125_));
  AOI21_X1   g23689(.A1(new_n26104_), .A2(new_n26107_), .B(new_n26125_), .ZN(new_n26126_));
  NOR3_X1    g23690(.A1(new_n13226_), .A2(new_n2709_), .A3(pi0907), .ZN(new_n26127_));
  OAI21_X1   g23691(.A1(new_n26098_), .A2(new_n26127_), .B(new_n5692_), .ZN(new_n26128_));
  NAND3_X1   g23692(.A1(new_n26128_), .A2(new_n5445_), .A3(new_n26093_), .ZN(new_n26129_));
  NOR2_X1    g23693(.A1(new_n26094_), .A2(new_n5449_), .ZN(new_n26130_));
  INV_X1     g23694(.I(new_n26130_), .ZN(new_n26131_));
  OAI21_X1   g23695(.A1(new_n26096_), .A2(new_n6745_), .B(new_n26131_), .ZN(new_n26132_));
  NAND2_X1   g23696(.A1(new_n26132_), .A2(pi0907), .ZN(new_n26133_));
  OAI21_X1   g23697(.A1(new_n24475_), .A2(new_n2709_), .B(new_n5473_), .ZN(new_n26134_));
  NAND3_X1   g23698(.A1(new_n26133_), .A2(new_n5692_), .A3(new_n26134_), .ZN(new_n26135_));
  AOI21_X1   g23699(.A1(new_n26086_), .A2(new_n5411_), .B(new_n5692_), .ZN(new_n26136_));
  AOI21_X1   g23700(.A1(new_n26085_), .A2(new_n5398_), .B(new_n5411_), .ZN(new_n26137_));
  OAI21_X1   g23701(.A1(new_n26091_), .A2(new_n5398_), .B(new_n26137_), .ZN(new_n26138_));
  AOI21_X1   g23702(.A1(new_n26138_), .A2(new_n26136_), .B(new_n5445_), .ZN(new_n26139_));
  NAND2_X1   g23703(.A1(new_n26135_), .A2(new_n26139_), .ZN(new_n26140_));
  NAND3_X1   g23704(.A1(new_n26129_), .A2(new_n26140_), .A3(new_n2642_), .ZN(new_n26141_));
  NAND2_X1   g23705(.A1(new_n26105_), .A2(new_n2641_), .ZN(new_n26142_));
  AOI21_X1   g23706(.A1(new_n26141_), .A2(new_n26142_), .B(pi0223), .ZN(new_n26143_));
  INV_X1     g23707(.I(new_n26136_), .ZN(new_n26144_));
  NAND2_X1   g23708(.A1(new_n26109_), .A2(new_n5437_), .ZN(new_n26145_));
  AOI21_X1   g23709(.A1(new_n26145_), .A2(new_n26137_), .B(new_n26144_), .ZN(new_n26146_));
  NAND2_X1   g23710(.A1(new_n26113_), .A2(new_n5449_), .ZN(new_n26147_));
  NAND2_X1   g23711(.A1(new_n26147_), .A2(new_n26131_), .ZN(new_n26148_));
  OAI21_X1   g23712(.A1(new_n26118_), .A2(pi0907), .B(new_n5692_), .ZN(new_n26149_));
  AOI21_X1   g23713(.A1(new_n26148_), .A2(pi0907), .B(new_n26149_), .ZN(new_n26150_));
  NOR3_X1    g23714(.A1(new_n26150_), .A2(new_n5445_), .A3(new_n26146_), .ZN(new_n26151_));
  AOI21_X1   g23715(.A1(new_n26115_), .A2(new_n26120_), .B(pi0947), .ZN(new_n26152_));
  NOR3_X1    g23716(.A1(new_n26152_), .A2(new_n5446_), .A3(new_n26111_), .ZN(new_n26153_));
  NOR3_X1    g23717(.A1(new_n26153_), .A2(new_n26151_), .A3(new_n2668_), .ZN(new_n26154_));
  NOR3_X1    g23718(.A1(new_n26143_), .A2(pi0299), .A3(new_n26154_), .ZN(new_n26155_));
  NOR3_X1    g23719(.A1(new_n26155_), .A2(new_n2627_), .A3(new_n26126_), .ZN(new_n26156_));
  OAI21_X1   g23720(.A1(new_n26156_), .A2(new_n26083_), .B(new_n8264_), .ZN(new_n26157_));
  OAI22_X1   g23721(.A1(new_n26157_), .A2(new_n26074_), .B1(new_n2709_), .B2(new_n8264_), .ZN(po0367));
  NOR2_X1    g23722(.A1(new_n16477_), .A2(new_n2610_), .ZN(new_n26159_));
  NAND2_X1   g23723(.A1(new_n26159_), .A2(pi0606), .ZN(new_n26160_));
  NOR2_X1    g23724(.A1(new_n16481_), .A2(new_n2610_), .ZN(new_n26161_));
  NAND2_X1   g23725(.A1(new_n26161_), .A2(new_n25131_), .ZN(new_n26162_));
  AOI21_X1   g23726(.A1(new_n26162_), .A2(new_n26160_), .B(new_n25167_), .ZN(new_n26163_));
  NAND2_X1   g23727(.A1(new_n16098_), .A2(new_n2609_), .ZN(new_n26164_));
  NOR3_X1    g23728(.A1(new_n26164_), .A2(new_n25131_), .A3(pi0643), .ZN(new_n26165_));
  NOR2_X1    g23729(.A1(new_n26163_), .A2(new_n26165_), .ZN(new_n26166_));
  NAND2_X1   g23730(.A1(new_n6643_), .A2(new_n8510_), .ZN(new_n26167_));
  NAND2_X1   g23731(.A1(new_n16470_), .A2(new_n2609_), .ZN(new_n26168_));
  NAND2_X1   g23732(.A1(new_n26168_), .A2(new_n25131_), .ZN(new_n26169_));
  NAND2_X1   g23733(.A1(new_n16473_), .A2(new_n2609_), .ZN(new_n26170_));
  NAND2_X1   g23734(.A1(new_n26170_), .A2(pi0606), .ZN(new_n26171_));
  AOI21_X1   g23735(.A1(new_n26171_), .A2(new_n26169_), .B(new_n25167_), .ZN(new_n26172_));
  NAND2_X1   g23736(.A1(new_n16119_), .A2(new_n2609_), .ZN(new_n26173_));
  NAND2_X1   g23737(.A1(new_n26173_), .A2(pi0606), .ZN(new_n26174_));
  NAND2_X1   g23738(.A1(new_n13192_), .A2(new_n25131_), .ZN(new_n26175_));
  AOI21_X1   g23739(.A1(new_n26174_), .A2(new_n26175_), .B(pi0643), .ZN(new_n26176_));
  NOR3_X1    g23740(.A1(new_n26176_), .A2(po1038), .A3(new_n26172_), .ZN(new_n26177_));
  OAI22_X1   g23741(.A1(new_n26177_), .A2(new_n8510_), .B1(new_n26166_), .B2(new_n26167_), .ZN(po0368));
  NAND2_X1   g23742(.A1(new_n26159_), .A2(pi0607), .ZN(new_n26179_));
  NAND2_X1   g23743(.A1(new_n26161_), .A2(new_n25938_), .ZN(new_n26180_));
  AOI21_X1   g23744(.A1(new_n26180_), .A2(new_n26179_), .B(new_n25921_), .ZN(new_n26181_));
  NOR3_X1    g23745(.A1(new_n26164_), .A2(new_n25938_), .A3(pi0638), .ZN(new_n26182_));
  NOR2_X1    g23746(.A1(new_n26181_), .A2(new_n26182_), .ZN(new_n26183_));
  NAND2_X1   g23747(.A1(new_n6643_), .A2(pi0212), .ZN(new_n26184_));
  NAND2_X1   g23748(.A1(new_n26168_), .A2(new_n25938_), .ZN(new_n26185_));
  NAND2_X1   g23749(.A1(new_n26170_), .A2(pi0607), .ZN(new_n26186_));
  AOI21_X1   g23750(.A1(new_n26186_), .A2(new_n26185_), .B(new_n25921_), .ZN(new_n26187_));
  NAND2_X1   g23751(.A1(new_n26173_), .A2(pi0607), .ZN(new_n26188_));
  NAND2_X1   g23752(.A1(new_n13192_), .A2(new_n25938_), .ZN(new_n26189_));
  AOI21_X1   g23753(.A1(new_n26188_), .A2(new_n26189_), .B(pi0638), .ZN(new_n26190_));
  NOR3_X1    g23754(.A1(new_n26190_), .A2(po1038), .A3(new_n26187_), .ZN(new_n26191_));
  OAI22_X1   g23755(.A1(new_n26191_), .A2(pi0212), .B1(new_n26183_), .B2(new_n26184_), .ZN(po0369));
  NAND2_X1   g23756(.A1(new_n26159_), .A2(pi0622), .ZN(new_n26193_));
  NAND2_X1   g23757(.A1(new_n26161_), .A2(new_n25973_), .ZN(new_n26194_));
  AOI21_X1   g23758(.A1(new_n26194_), .A2(new_n26193_), .B(new_n25966_), .ZN(new_n26195_));
  NOR3_X1    g23759(.A1(new_n26164_), .A2(new_n25973_), .A3(pi0639), .ZN(new_n26196_));
  NOR2_X1    g23760(.A1(new_n26195_), .A2(new_n26196_), .ZN(new_n26197_));
  INV_X1     g23761(.I(pi0213), .ZN(new_n26198_));
  NOR2_X1    g23762(.A1(po1038), .A2(new_n26198_), .ZN(new_n26199_));
  INV_X1     g23763(.I(new_n26199_), .ZN(new_n26200_));
  NAND2_X1   g23764(.A1(new_n26173_), .A2(new_n25966_), .ZN(new_n26201_));
  NAND2_X1   g23765(.A1(new_n26170_), .A2(pi0639), .ZN(new_n26202_));
  AOI21_X1   g23766(.A1(new_n26201_), .A2(new_n26202_), .B(new_n25973_), .ZN(new_n26203_));
  NAND2_X1   g23767(.A1(new_n26168_), .A2(pi0639), .ZN(new_n26204_));
  NAND2_X1   g23768(.A1(new_n13192_), .A2(new_n25966_), .ZN(new_n26205_));
  AOI21_X1   g23769(.A1(new_n26204_), .A2(new_n26205_), .B(pi0622), .ZN(new_n26206_));
  NOR3_X1    g23770(.A1(new_n26203_), .A2(po1038), .A3(new_n26206_), .ZN(new_n26207_));
  OAI22_X1   g23771(.A1(new_n26207_), .A2(pi0213), .B1(new_n26197_), .B2(new_n26200_), .ZN(po0370));
  NAND2_X1   g23772(.A1(new_n26159_), .A2(pi0623), .ZN(new_n26209_));
  NAND2_X1   g23773(.A1(new_n26161_), .A2(new_n25648_), .ZN(new_n26210_));
  AOI21_X1   g23774(.A1(new_n26210_), .A2(new_n26209_), .B(new_n25607_), .ZN(new_n26211_));
  NOR3_X1    g23775(.A1(new_n26164_), .A2(new_n25648_), .A3(pi0710), .ZN(new_n26212_));
  NOR2_X1    g23776(.A1(new_n26211_), .A2(new_n26212_), .ZN(new_n26213_));
  NAND2_X1   g23777(.A1(new_n6643_), .A2(pi0214), .ZN(new_n26214_));
  NAND2_X1   g23778(.A1(new_n26168_), .A2(new_n25648_), .ZN(new_n26215_));
  NAND2_X1   g23779(.A1(new_n26170_), .A2(pi0623), .ZN(new_n26216_));
  AOI21_X1   g23780(.A1(new_n26216_), .A2(new_n26215_), .B(new_n25607_), .ZN(new_n26217_));
  NAND2_X1   g23781(.A1(new_n26173_), .A2(pi0623), .ZN(new_n26218_));
  NAND2_X1   g23782(.A1(new_n13192_), .A2(new_n25648_), .ZN(new_n26219_));
  AOI21_X1   g23783(.A1(new_n26218_), .A2(new_n26219_), .B(pi0710), .ZN(new_n26220_));
  NOR3_X1    g23784(.A1(new_n26220_), .A2(po1038), .A3(new_n26217_), .ZN(new_n26221_));
  OAI22_X1   g23785(.A1(new_n26221_), .A2(pi0214), .B1(new_n26213_), .B2(new_n26214_), .ZN(po0371));
  NAND2_X1   g23786(.A1(new_n13397_), .A2(new_n2436_), .ZN(new_n26223_));
  NOR2_X1    g23787(.A1(new_n5399_), .A2(new_n5473_), .ZN(new_n26224_));
  NOR2_X1    g23788(.A1(new_n26224_), .A2(pi0947), .ZN(new_n26225_));
  AOI21_X1   g23789(.A1(new_n5406_), .A2(pi0947), .B(new_n26225_), .ZN(new_n26226_));
  INV_X1     g23790(.I(new_n26226_), .ZN(new_n26227_));
  NAND2_X1   g23791(.A1(new_n13344_), .A2(new_n26227_), .ZN(new_n26228_));
  AOI21_X1   g23792(.A1(new_n26223_), .A2(new_n26228_), .B(new_n3265_), .ZN(new_n26229_));
  NAND2_X1   g23793(.A1(new_n13058_), .A2(new_n2436_), .ZN(new_n26230_));
  NAND2_X1   g23794(.A1(new_n15945_), .A2(new_n26227_), .ZN(new_n26231_));
  AOI21_X1   g23795(.A1(new_n26231_), .A2(new_n26230_), .B(pi0299), .ZN(new_n26232_));
  NOR2_X1    g23796(.A1(new_n14557_), .A2(pi0215), .ZN(new_n26233_));
  NOR2_X1    g23797(.A1(new_n13055_), .A2(new_n26226_), .ZN(new_n26234_));
  OAI21_X1   g23798(.A1(new_n26233_), .A2(new_n26234_), .B(pi0299), .ZN(new_n26235_));
  NAND2_X1   g23799(.A1(new_n26235_), .A2(new_n2627_), .ZN(new_n26236_));
  OAI21_X1   g23800(.A1(new_n26236_), .A2(new_n26232_), .B(new_n3265_), .ZN(new_n26237_));
  NOR2_X1    g23801(.A1(new_n13144_), .A2(new_n5445_), .ZN(new_n26238_));
  INV_X1     g23802(.I(new_n26238_), .ZN(new_n26239_));
  AOI21_X1   g23803(.A1(new_n26239_), .A2(new_n26224_), .B(pi0947), .ZN(new_n26240_));
  NOR2_X1    g23804(.A1(new_n13120_), .A2(new_n5406_), .ZN(new_n26241_));
  NAND2_X1   g23805(.A1(new_n13122_), .A2(pi0642), .ZN(new_n26242_));
  NOR2_X1    g23806(.A1(new_n13151_), .A2(new_n26242_), .ZN(new_n26243_));
  NOR3_X1    g23807(.A1(new_n26243_), .A2(new_n5692_), .A3(new_n26241_), .ZN(new_n26244_));
  NAND2_X1   g23808(.A1(new_n13169_), .A2(pi0947), .ZN(new_n26245_));
  AND3_X2    g23809(.A1(new_n13466_), .A2(new_n5445_), .A3(new_n26245_), .Z(new_n26246_));
  OR3_X2     g23810(.A1(new_n26240_), .A2(new_n26246_), .A3(new_n26244_), .Z(new_n26247_));
  NOR2_X1    g23811(.A1(new_n13304_), .A2(new_n12821_), .ZN(new_n26248_));
  NOR2_X1    g23812(.A1(new_n26248_), .A2(new_n26242_), .ZN(new_n26249_));
  OAI21_X1   g23813(.A1(new_n26249_), .A2(new_n26241_), .B(pi0947), .ZN(new_n26250_));
  NOR2_X1    g23814(.A1(new_n13103_), .A2(new_n13105_), .ZN(new_n26251_));
  INV_X1     g23815(.I(new_n26251_), .ZN(new_n26252_));
  INV_X1     g23816(.I(new_n26224_), .ZN(new_n26253_));
  NOR2_X1    g23817(.A1(new_n26253_), .A2(pi0947), .ZN(new_n26254_));
  AOI21_X1   g23818(.A1(new_n26252_), .A2(new_n26254_), .B(new_n5445_), .ZN(new_n26255_));
  NAND2_X1   g23819(.A1(new_n26255_), .A2(new_n26250_), .ZN(new_n26256_));
  INV_X1     g23820(.I(new_n13225_), .ZN(new_n26257_));
  AOI21_X1   g23821(.A1(new_n13603_), .A2(new_n5403_), .B(new_n26257_), .ZN(new_n26258_));
  NOR3_X1    g23822(.A1(new_n26258_), .A2(new_n5406_), .A3(new_n13119_), .ZN(new_n26259_));
  NAND3_X1   g23823(.A1(new_n13603_), .A2(pi0642), .A3(new_n13119_), .ZN(new_n26260_));
  NAND2_X1   g23824(.A1(new_n26260_), .A2(pi0947), .ZN(new_n26261_));
  NOR2_X1    g23825(.A1(new_n13090_), .A2(new_n26253_), .ZN(new_n26262_));
  OAI22_X1   g23826(.A1(new_n26259_), .A2(new_n26261_), .B1(pi0947), .B2(new_n26262_), .ZN(new_n26263_));
  NAND2_X1   g23827(.A1(new_n26263_), .A2(new_n5445_), .ZN(new_n26264_));
  NAND3_X1   g23828(.A1(new_n26264_), .A2(new_n2642_), .A3(new_n26256_), .ZN(new_n26265_));
  AOI21_X1   g23829(.A1(new_n13185_), .A2(new_n26226_), .B(pi0223), .ZN(new_n26266_));
  AOI22_X1   g23830(.A1(new_n26265_), .A2(new_n26266_), .B1(pi0223), .B2(new_n26247_), .ZN(new_n26267_));
  AOI21_X1   g23831(.A1(new_n13639_), .A2(new_n26226_), .B(new_n2628_), .ZN(new_n26268_));
  OR2_X2     g23832(.A1(new_n26263_), .A2(new_n3303_), .Z(new_n26269_));
  AOI21_X1   g23833(.A1(new_n26269_), .A2(new_n26268_), .B(pi0215), .ZN(new_n26270_));
  OAI21_X1   g23834(.A1(new_n26267_), .A2(pi0299), .B(new_n26270_), .ZN(new_n26271_));
  NAND2_X1   g23835(.A1(new_n13098_), .A2(new_n26227_), .ZN(new_n26272_));
  AOI21_X1   g23836(.A1(new_n26272_), .A2(new_n2641_), .B(pi0223), .ZN(new_n26273_));
  INV_X1     g23837(.I(new_n13730_), .ZN(new_n26274_));
  OAI21_X1   g23838(.A1(new_n13104_), .A2(pi0642), .B(new_n5403_), .ZN(new_n26275_));
  AOI21_X1   g23839(.A1(new_n26274_), .A2(new_n5408_), .B(new_n26275_), .ZN(new_n26276_));
  AOI21_X1   g23840(.A1(new_n13304_), .A2(new_n5406_), .B(new_n5403_), .ZN(new_n26277_));
  NOR3_X1    g23841(.A1(new_n26276_), .A2(new_n5445_), .A3(new_n26277_), .ZN(new_n26278_));
  NOR3_X1    g23842(.A1(new_n13308_), .A2(pi0642), .A3(new_n5446_), .ZN(new_n26279_));
  OAI21_X1   g23843(.A1(new_n26279_), .A2(new_n26278_), .B(pi0947), .ZN(new_n26280_));
  NAND2_X1   g23844(.A1(new_n16315_), .A2(new_n26225_), .ZN(new_n26281_));
  NAND3_X1   g23845(.A1(new_n26281_), .A2(new_n2642_), .A3(new_n26280_), .ZN(new_n26282_));
  OAI21_X1   g23846(.A1(new_n13143_), .A2(new_n5404_), .B(new_n13271_), .ZN(new_n26283_));
  NAND3_X1   g23847(.A1(new_n26283_), .A2(new_n5406_), .A3(new_n5446_), .ZN(new_n26284_));
  NAND3_X1   g23848(.A1(new_n13149_), .A2(new_n13163_), .A3(new_n13116_), .ZN(new_n26285_));
  NAND2_X1   g23849(.A1(new_n13466_), .A2(new_n5403_), .ZN(new_n26286_));
  NAND4_X1   g23850(.A1(new_n26286_), .A2(new_n5406_), .A3(new_n5445_), .A4(new_n26285_), .ZN(new_n26287_));
  AOI21_X1   g23851(.A1(new_n26287_), .A2(new_n26284_), .B(new_n5692_), .ZN(new_n26288_));
  OAI21_X1   g23852(.A1(new_n16042_), .A2(new_n26288_), .B(pi0223), .ZN(new_n26289_));
  OAI21_X1   g23853(.A1(new_n26289_), .A2(new_n26254_), .B(new_n2628_), .ZN(new_n26290_));
  AOI21_X1   g23854(.A1(new_n26273_), .A2(new_n26282_), .B(new_n26290_), .ZN(new_n26291_));
  NAND2_X1   g23855(.A1(new_n16254_), .A2(new_n5692_), .ZN(new_n26292_));
  NAND4_X1   g23856(.A1(new_n26286_), .A2(new_n5406_), .A3(pi0947), .A4(new_n26285_), .ZN(new_n26293_));
  OAI21_X1   g23857(.A1(pi0947), .A2(new_n26224_), .B(new_n26293_), .ZN(new_n26294_));
  AOI21_X1   g23858(.A1(new_n26292_), .A2(new_n26294_), .B(new_n2628_), .ZN(new_n26295_));
  OAI21_X1   g23859(.A1(new_n26291_), .A2(new_n26295_), .B(pi0215), .ZN(new_n26296_));
  AOI21_X1   g23860(.A1(new_n26296_), .A2(new_n26271_), .B(new_n2627_), .ZN(new_n26297_));
  OAI21_X1   g23861(.A1(new_n26297_), .A2(new_n26237_), .B(new_n8264_), .ZN(new_n26298_));
  OAI22_X1   g23862(.A1(new_n26298_), .A2(new_n26229_), .B1(new_n2436_), .B2(new_n8264_), .ZN(po0372));
  NOR2_X1    g23863(.A1(new_n13344_), .A2(pi0216), .ZN(new_n26300_));
  NOR2_X1    g23864(.A1(new_n15994_), .A2(new_n5400_), .ZN(new_n26301_));
  NOR2_X1    g23865(.A1(new_n5405_), .A2(new_n5692_), .ZN(new_n26302_));
  NOR2_X1    g23866(.A1(new_n26301_), .A2(new_n26302_), .ZN(new_n26303_));
  INV_X1     g23867(.I(new_n26303_), .ZN(new_n26304_));
  NOR2_X1    g23868(.A1(new_n13397_), .A2(new_n26304_), .ZN(new_n26305_));
  OAI21_X1   g23869(.A1(new_n26305_), .A2(new_n26300_), .B(pi0038), .ZN(new_n26306_));
  NOR2_X1    g23870(.A1(new_n15945_), .A2(pi0216), .ZN(new_n26307_));
  NOR2_X1    g23871(.A1(new_n13058_), .A2(new_n26304_), .ZN(new_n26308_));
  OAI21_X1   g23872(.A1(new_n26307_), .A2(new_n26308_), .B(new_n2628_), .ZN(new_n26309_));
  NAND2_X1   g23873(.A1(new_n13055_), .A2(new_n2614_), .ZN(new_n26310_));
  OAI21_X1   g23874(.A1(new_n13055_), .A2(new_n26304_), .B(new_n26310_), .ZN(new_n26311_));
  AOI21_X1   g23875(.A1(new_n26311_), .A2(pi0299), .B(pi0039), .ZN(new_n26312_));
  AOI21_X1   g23876(.A1(new_n26312_), .A2(new_n26309_), .B(pi0038), .ZN(new_n26313_));
  NOR2_X1    g23877(.A1(new_n5400_), .A2(new_n5473_), .ZN(new_n26314_));
  NAND2_X1   g23878(.A1(new_n26239_), .A2(new_n26314_), .ZN(new_n26315_));
  NAND2_X1   g23879(.A1(new_n26315_), .A2(new_n5692_), .ZN(new_n26316_));
  OAI21_X1   g23880(.A1(new_n13151_), .A2(new_n13123_), .B(pi0947), .ZN(new_n26317_));
  NOR2_X1    g23881(.A1(new_n26317_), .A2(new_n13121_), .ZN(new_n26318_));
  NOR2_X1    g23882(.A1(new_n26246_), .A2(new_n26318_), .ZN(new_n26319_));
  AOI21_X1   g23883(.A1(new_n26319_), .A2(new_n26316_), .B(new_n2668_), .ZN(new_n26320_));
  OAI21_X1   g23884(.A1(new_n16045_), .A2(new_n26303_), .B(new_n2668_), .ZN(new_n26321_));
  OAI21_X1   g23885(.A1(new_n13124_), .A2(new_n13121_), .B(pi0947), .ZN(new_n26322_));
  NAND2_X1   g23886(.A1(new_n26252_), .A2(new_n26301_), .ZN(new_n26323_));
  NAND3_X1   g23887(.A1(new_n26323_), .A2(new_n5446_), .A3(new_n26322_), .ZN(new_n26324_));
  INV_X1     g23888(.I(new_n26258_), .ZN(new_n26325_));
  AOI22_X1   g23889(.A1(new_n26325_), .A2(new_n26302_), .B1(new_n13485_), .B2(new_n26301_), .ZN(new_n26326_));
  AOI21_X1   g23890(.A1(new_n26326_), .A2(new_n5445_), .B(new_n2641_), .ZN(new_n26327_));
  AOI21_X1   g23891(.A1(new_n26327_), .A2(new_n26324_), .B(new_n26321_), .ZN(new_n26328_));
  NOR3_X1    g23892(.A1(new_n26328_), .A2(pi0216), .A3(new_n26320_), .ZN(new_n26329_));
  INV_X1     g23893(.I(new_n26301_), .ZN(new_n26330_));
  NAND2_X1   g23894(.A1(new_n26330_), .A2(pi0223), .ZN(new_n26331_));
  NOR2_X1    g23895(.A1(new_n5405_), .A2(pi0616), .ZN(new_n26332_));
  NOR2_X1    g23896(.A1(new_n24468_), .A2(new_n26332_), .ZN(new_n26333_));
  NOR2_X1    g23897(.A1(new_n26333_), .A2(new_n5404_), .ZN(new_n26334_));
  AOI21_X1   g23898(.A1(new_n5404_), .A2(new_n13274_), .B(new_n26334_), .ZN(new_n26335_));
  NOR2_X1    g23899(.A1(new_n26335_), .A2(pi0614), .ZN(new_n26336_));
  NAND2_X1   g23900(.A1(new_n26336_), .A2(new_n5445_), .ZN(new_n26337_));
  OAI21_X1   g23901(.A1(new_n13142_), .A2(pi0616), .B(new_n13112_), .ZN(new_n26338_));
  OAI21_X1   g23902(.A1(new_n26338_), .A2(new_n5404_), .B(new_n13271_), .ZN(new_n26339_));
  NAND3_X1   g23903(.A1(new_n26339_), .A2(new_n5405_), .A3(new_n5446_), .ZN(new_n26340_));
  AOI21_X1   g23904(.A1(new_n26337_), .A2(new_n26340_), .B(new_n5692_), .ZN(new_n26341_));
  NOR2_X1    g23905(.A1(new_n16042_), .A2(new_n26341_), .ZN(new_n26342_));
  OAI21_X1   g23906(.A1(new_n26342_), .A2(new_n26331_), .B(pi0216), .ZN(new_n26343_));
  OAI21_X1   g23907(.A1(new_n13088_), .A2(new_n26304_), .B(new_n2641_), .ZN(new_n26344_));
  NAND2_X1   g23908(.A1(new_n26344_), .A2(new_n2668_), .ZN(new_n26345_));
  NOR3_X1    g23909(.A1(new_n14577_), .A2(pi0947), .A3(new_n26314_), .ZN(new_n26346_));
  NOR2_X1    g23910(.A1(new_n13115_), .A2(new_n5692_), .ZN(new_n26347_));
  OAI21_X1   g23911(.A1(new_n26346_), .A2(new_n26347_), .B(new_n5446_), .ZN(new_n26348_));
  AOI21_X1   g23912(.A1(new_n13226_), .A2(new_n5405_), .B(new_n5692_), .ZN(new_n26349_));
  NOR3_X1    g23913(.A1(new_n26349_), .A2(new_n5446_), .A3(new_n26301_), .ZN(new_n26350_));
  NAND2_X1   g23914(.A1(new_n13093_), .A2(new_n5692_), .ZN(new_n26351_));
  AOI21_X1   g23915(.A1(new_n26350_), .A2(new_n26351_), .B(new_n2641_), .ZN(new_n26352_));
  AOI21_X1   g23916(.A1(new_n26348_), .A2(new_n26352_), .B(new_n26345_), .ZN(new_n26353_));
  OAI21_X1   g23917(.A1(new_n26343_), .A2(new_n26353_), .B(new_n2628_), .ZN(new_n26354_));
  OAI21_X1   g23918(.A1(new_n26354_), .A2(new_n26329_), .B(pi0039), .ZN(new_n26355_));
  INV_X1     g23919(.I(new_n26326_), .ZN(new_n26356_));
  AOI22_X1   g23920(.A1(new_n26356_), .A2(new_n5056_), .B1(new_n13639_), .B2(new_n26304_), .ZN(new_n26357_));
  AOI21_X1   g23921(.A1(new_n16108_), .A2(new_n5692_), .B(new_n26349_), .ZN(new_n26358_));
  OAI21_X1   g23922(.A1(new_n5400_), .A2(new_n15994_), .B(new_n26358_), .ZN(new_n26359_));
  NAND2_X1   g23923(.A1(new_n26359_), .A2(pi0216), .ZN(new_n26360_));
  NAND2_X1   g23924(.A1(new_n26360_), .A2(new_n26357_), .ZN(new_n26361_));
  NAND2_X1   g23925(.A1(new_n13171_), .A2(new_n26301_), .ZN(new_n26362_));
  AOI21_X1   g23926(.A1(new_n26362_), .A2(new_n26245_), .B(new_n26318_), .ZN(new_n26363_));
  OAI21_X1   g23927(.A1(new_n26363_), .A2(pi0216), .B(pi0215), .ZN(new_n26364_));
  INV_X1     g23928(.I(new_n26292_), .ZN(new_n26365_));
  NOR2_X1    g23929(.A1(new_n26336_), .A2(new_n5692_), .ZN(new_n26366_));
  NOR4_X1    g23930(.A1(new_n26365_), .A2(new_n2614_), .A3(new_n26301_), .A4(new_n26366_), .ZN(new_n26367_));
  OAI21_X1   g23931(.A1(new_n26367_), .A2(new_n26364_), .B(pi0299), .ZN(new_n26368_));
  AOI21_X1   g23932(.A1(new_n26361_), .A2(new_n2436_), .B(new_n26368_), .ZN(new_n26369_));
  OAI21_X1   g23933(.A1(new_n26369_), .A2(new_n26355_), .B(new_n26313_), .ZN(new_n26370_));
  NAND3_X1   g23934(.A1(new_n26370_), .A2(new_n8264_), .A3(new_n26306_), .ZN(new_n26371_));
  OAI21_X1   g23935(.A1(new_n2614_), .A2(new_n8264_), .B(new_n26371_), .ZN(po0373));
  INV_X1     g23936(.I(pi0612), .ZN(new_n26373_));
  OAI21_X1   g23937(.A1(new_n25987_), .A2(pi0695), .B(pi0217), .ZN(new_n26374_));
  NAND2_X1   g23938(.A1(new_n26374_), .A2(new_n26373_), .ZN(new_n26375_));
  INV_X1     g23939(.I(pi0695), .ZN(new_n26376_));
  AOI21_X1   g23940(.A1(new_n13191_), .A2(new_n8264_), .B(new_n26376_), .ZN(new_n26377_));
  NOR2_X1    g23941(.A1(new_n26066_), .A2(pi0695), .ZN(new_n26378_));
  NOR3_X1    g23942(.A1(new_n26378_), .A2(pi0217), .A3(new_n26377_), .ZN(new_n26379_));
  NOR2_X1    g23943(.A1(new_n26048_), .A2(new_n26376_), .ZN(new_n26380_));
  NOR3_X1    g23944(.A1(new_n26042_), .A2(pi0695), .A3(new_n26026_), .ZN(new_n26381_));
  OAI21_X1   g23945(.A1(new_n26381_), .A2(new_n26380_), .B(new_n9751_), .ZN(new_n26382_));
  AOI21_X1   g23946(.A1(new_n26012_), .A2(new_n26002_), .B(pi0695), .ZN(new_n26383_));
  NOR2_X1    g23947(.A1(new_n25970_), .A2(new_n26376_), .ZN(new_n26384_));
  OAI21_X1   g23948(.A1(new_n26383_), .A2(new_n26384_), .B(pi0217), .ZN(new_n26385_));
  NAND3_X1   g23949(.A1(new_n26385_), .A2(pi0612), .A3(new_n26382_), .ZN(new_n26386_));
  OAI21_X1   g23950(.A1(new_n26375_), .A2(new_n26379_), .B(new_n26386_), .ZN(po0374));
  NOR2_X1    g23951(.A1(new_n25474_), .A2(new_n25466_), .ZN(new_n26388_));
  NAND2_X1   g23952(.A1(new_n26388_), .A2(pi0218), .ZN(new_n26389_));
  NOR2_X1    g23953(.A1(new_n25543_), .A2(new_n25465_), .ZN(new_n26390_));
  AOI21_X1   g23954(.A1(new_n25521_), .A2(new_n25465_), .B(new_n26390_), .ZN(new_n26391_));
  OAI21_X1   g23955(.A1(new_n26391_), .A2(pi0218), .B(new_n26389_), .ZN(po0375));
  NAND2_X1   g23956(.A1(new_n26159_), .A2(pi0617), .ZN(new_n26393_));
  NAND2_X1   g23957(.A1(new_n26161_), .A2(new_n24970_), .ZN(new_n26394_));
  AOI21_X1   g23958(.A1(new_n26394_), .A2(new_n26393_), .B(new_n24943_), .ZN(new_n26395_));
  NOR3_X1    g23959(.A1(new_n26164_), .A2(new_n24970_), .A3(pi0637), .ZN(new_n26396_));
  NOR2_X1    g23960(.A1(po1038), .A2(pi0219), .ZN(new_n26397_));
  OAI21_X1   g23961(.A1(new_n26395_), .A2(new_n26396_), .B(new_n26397_), .ZN(new_n26398_));
  NAND2_X1   g23962(.A1(new_n26168_), .A2(new_n24970_), .ZN(new_n26399_));
  NAND2_X1   g23963(.A1(new_n26170_), .A2(pi0617), .ZN(new_n26400_));
  AOI21_X1   g23964(.A1(new_n26400_), .A2(new_n26399_), .B(new_n24943_), .ZN(new_n26401_));
  NAND2_X1   g23965(.A1(new_n26173_), .A2(pi0617), .ZN(new_n26402_));
  NAND2_X1   g23966(.A1(new_n13192_), .A2(new_n24970_), .ZN(new_n26403_));
  AOI21_X1   g23967(.A1(new_n26402_), .A2(new_n26403_), .B(pi0637), .ZN(new_n26404_));
  NOR3_X1    g23968(.A1(new_n26404_), .A2(po1038), .A3(new_n26401_), .ZN(new_n26405_));
  OAI21_X1   g23969(.A1(new_n26405_), .A2(new_n8807_), .B(new_n26398_), .ZN(po0376));
  NOR2_X1    g23970(.A1(new_n25325_), .A2(new_n25553_), .ZN(new_n26407_));
  NAND2_X1   g23971(.A1(new_n26407_), .A2(pi0220), .ZN(new_n26408_));
  NOR2_X1    g23972(.A1(new_n25454_), .A2(new_n25552_), .ZN(new_n26409_));
  AOI21_X1   g23973(.A1(new_n25435_), .A2(new_n25552_), .B(new_n26409_), .ZN(new_n26410_));
  OAI21_X1   g23974(.A1(new_n26410_), .A2(pi0220), .B(new_n26408_), .ZN(po0377));
  NAND2_X1   g23975(.A1(new_n13397_), .A2(new_n2441_), .ZN(new_n26412_));
  INV_X1     g23976(.I(pi0661), .ZN(new_n26413_));
  NOR2_X1    g23977(.A1(new_n15994_), .A2(new_n26413_), .ZN(new_n26414_));
  NOR2_X1    g23978(.A1(new_n13111_), .A2(new_n5692_), .ZN(new_n26415_));
  NOR2_X1    g23979(.A1(new_n26414_), .A2(new_n26415_), .ZN(new_n26416_));
  NAND2_X1   g23980(.A1(new_n13344_), .A2(new_n26416_), .ZN(new_n26417_));
  AOI21_X1   g23981(.A1(new_n26412_), .A2(new_n26417_), .B(new_n3265_), .ZN(new_n26418_));
  NAND2_X1   g23982(.A1(new_n13058_), .A2(new_n2441_), .ZN(new_n26419_));
  NAND2_X1   g23983(.A1(new_n15945_), .A2(new_n26416_), .ZN(new_n26420_));
  AOI21_X1   g23984(.A1(new_n26420_), .A2(new_n26419_), .B(pi0299), .ZN(new_n26421_));
  NOR2_X1    g23985(.A1(new_n14557_), .A2(pi0221), .ZN(new_n26422_));
  INV_X1     g23986(.I(new_n26416_), .ZN(new_n26423_));
  NOR2_X1    g23987(.A1(new_n13055_), .A2(new_n26423_), .ZN(new_n26424_));
  OAI21_X1   g23988(.A1(new_n26422_), .A2(new_n26424_), .B(pi0299), .ZN(new_n26425_));
  NAND2_X1   g23989(.A1(new_n26425_), .A2(new_n2627_), .ZN(new_n26426_));
  OAI21_X1   g23990(.A1(new_n26426_), .A2(new_n26421_), .B(new_n3265_), .ZN(new_n26427_));
  NOR2_X1    g23991(.A1(new_n13088_), .A2(pi0216), .ZN(new_n26428_));
  AOI21_X1   g23992(.A1(new_n26428_), .A2(new_n26423_), .B(pi0221), .ZN(new_n26429_));
  AOI22_X1   g23993(.A1(new_n26325_), .A2(new_n26415_), .B1(new_n13485_), .B2(new_n26414_), .ZN(new_n26430_));
  OR2_X2     g23994(.A1(new_n26430_), .A2(new_n2614_), .Z(new_n26431_));
  AOI21_X1   g23995(.A1(new_n26431_), .A2(new_n26429_), .B(pi0215), .ZN(new_n26432_));
  NOR2_X1    g23996(.A1(new_n13308_), .A2(pi0642), .ZN(new_n26433_));
  OAI21_X1   g23997(.A1(new_n26259_), .A2(new_n26433_), .B(new_n13157_), .ZN(new_n26434_));
  NAND2_X1   g23998(.A1(new_n13082_), .A2(new_n5398_), .ZN(new_n26435_));
  OAI21_X1   g23999(.A1(new_n13303_), .A2(new_n13099_), .B(new_n13100_), .ZN(new_n26436_));
  AOI21_X1   g24000(.A1(new_n26436_), .A2(new_n5405_), .B(new_n13153_), .ZN(new_n26437_));
  OAI21_X1   g24001(.A1(new_n26437_), .A2(new_n5398_), .B(new_n26435_), .ZN(new_n26438_));
  NAND3_X1   g24002(.A1(new_n26438_), .A2(new_n13111_), .A3(new_n13119_), .ZN(new_n26439_));
  NAND3_X1   g24003(.A1(new_n26434_), .A2(new_n26439_), .A3(pi0947), .ZN(new_n26440_));
  NOR2_X1    g24004(.A1(new_n26413_), .A2(new_n5473_), .ZN(new_n26441_));
  OAI21_X1   g24005(.A1(new_n16108_), .A2(new_n26441_), .B(new_n5692_), .ZN(new_n26442_));
  NAND3_X1   g24006(.A1(new_n26442_), .A2(pi0221), .A3(new_n26440_), .ZN(new_n26443_));
  AND2_X2    g24007(.A1(new_n13152_), .A2(pi0947), .Z(new_n26444_));
  NOR2_X1    g24008(.A1(new_n26444_), .A2(new_n26414_), .ZN(new_n26445_));
  AOI21_X1   g24009(.A1(new_n13466_), .A2(new_n26245_), .B(new_n26445_), .ZN(new_n26446_));
  OAI21_X1   g24010(.A1(new_n26446_), .A2(pi0221), .B(pi0215), .ZN(new_n26447_));
  OAI21_X1   g24011(.A1(pi0614), .A2(new_n13142_), .B(new_n13169_), .ZN(new_n26448_));
  AOI21_X1   g24012(.A1(new_n26448_), .A2(new_n5403_), .B(pi0616), .ZN(new_n26449_));
  AOI21_X1   g24013(.A1(new_n26449_), .A2(new_n26285_), .B(new_n5692_), .ZN(new_n26450_));
  NOR4_X1    g24014(.A1(new_n26365_), .A2(new_n2441_), .A3(new_n26414_), .A4(new_n26450_), .ZN(new_n26451_));
  OAI21_X1   g24015(.A1(new_n26451_), .A2(new_n26447_), .B(pi0299), .ZN(new_n26452_));
  AOI21_X1   g24016(.A1(new_n26432_), .A2(new_n26443_), .B(new_n26452_), .ZN(new_n26453_));
  AOI21_X1   g24017(.A1(new_n26239_), .A2(new_n26414_), .B(new_n26444_), .ZN(new_n26454_));
  OAI21_X1   g24018(.A1(new_n26454_), .A2(new_n26246_), .B(pi0223), .ZN(new_n26455_));
  NAND2_X1   g24019(.A1(new_n26455_), .A2(new_n2441_), .ZN(new_n26456_));
  AOI21_X1   g24020(.A1(new_n13185_), .A2(new_n26423_), .B(pi0223), .ZN(new_n26457_));
  INV_X1     g24021(.I(new_n26457_), .ZN(new_n26458_));
  OAI22_X1   g24022(.A1(new_n26248_), .A2(new_n13146_), .B1(new_n13111_), .B2(new_n13120_), .ZN(new_n26459_));
  NAND2_X1   g24023(.A1(new_n26459_), .A2(pi0947), .ZN(new_n26460_));
  AOI21_X1   g24024(.A1(new_n26252_), .A2(new_n26414_), .B(new_n5445_), .ZN(new_n26461_));
  NAND2_X1   g24025(.A1(new_n26461_), .A2(new_n26460_), .ZN(new_n26462_));
  AOI21_X1   g24026(.A1(new_n26430_), .A2(new_n5445_), .B(new_n2641_), .ZN(new_n26463_));
  AOI21_X1   g24027(.A1(new_n26463_), .A2(new_n26462_), .B(new_n26458_), .ZN(new_n26464_));
  OAI21_X1   g24028(.A1(new_n26464_), .A2(new_n26456_), .B(new_n2628_), .ZN(new_n26465_));
  NAND2_X1   g24029(.A1(new_n14577_), .A2(new_n5692_), .ZN(new_n26466_));
  OAI21_X1   g24030(.A1(new_n13123_), .A2(new_n26248_), .B(new_n13115_), .ZN(new_n26467_));
  NOR2_X1    g24031(.A1(new_n26437_), .A2(new_n13118_), .ZN(new_n26468_));
  AOI21_X1   g24032(.A1(new_n26467_), .A2(new_n13118_), .B(new_n26468_), .ZN(new_n26469_));
  OAI21_X1   g24033(.A1(new_n26469_), .A2(pi0616), .B(pi0947), .ZN(new_n26470_));
  AOI21_X1   g24034(.A1(new_n26470_), .A2(new_n26466_), .B(new_n5445_), .ZN(new_n26471_));
  AOI21_X1   g24035(.A1(new_n26440_), .A2(new_n26351_), .B(new_n5446_), .ZN(new_n26472_));
  NOR4_X1    g24036(.A1(new_n26471_), .A2(new_n2641_), .A3(new_n26472_), .A4(new_n26414_), .ZN(new_n26473_));
  OAI21_X1   g24037(.A1(new_n26473_), .A2(new_n13185_), .B(new_n26457_), .ZN(new_n26474_));
  AOI21_X1   g24038(.A1(new_n15956_), .A2(new_n5692_), .B(new_n26450_), .ZN(new_n26475_));
  NOR2_X1    g24039(.A1(new_n26475_), .A2(new_n5446_), .ZN(new_n26476_));
  NAND2_X1   g24040(.A1(new_n15953_), .A2(new_n5692_), .ZN(new_n26477_));
  OR3_X2     g24041(.A1(new_n13160_), .A2(new_n5692_), .A3(new_n13156_), .Z(new_n26478_));
  AOI21_X1   g24042(.A1(new_n26477_), .A2(new_n26478_), .B(new_n5445_), .ZN(new_n26479_));
  NOR4_X1    g24043(.A1(new_n26479_), .A2(new_n2668_), .A3(new_n26414_), .A4(new_n26476_), .ZN(new_n26480_));
  NOR2_X1    g24044(.A1(new_n26480_), .A2(new_n2441_), .ZN(new_n26481_));
  AOI21_X1   g24045(.A1(new_n26474_), .A2(new_n26481_), .B(new_n26465_), .ZN(new_n26482_));
  NOR3_X1    g24046(.A1(new_n26453_), .A2(new_n2627_), .A3(new_n26482_), .ZN(new_n26483_));
  OAI21_X1   g24047(.A1(new_n26483_), .A2(new_n26427_), .B(new_n8264_), .ZN(new_n26484_));
  OAI22_X1   g24048(.A1(new_n26484_), .A2(new_n26418_), .B1(new_n2441_), .B2(new_n8264_), .ZN(po0378));
  NAND2_X1   g24049(.A1(po1038), .A2(pi0222), .ZN(new_n26486_));
  NAND2_X1   g24050(.A1(new_n13184_), .A2(new_n2668_), .ZN(new_n26487_));
  AOI21_X1   g24051(.A1(new_n26487_), .A2(new_n13182_), .B(pi0299), .ZN(new_n26488_));
  NOR3_X1    g24052(.A1(new_n13178_), .A2(new_n2627_), .A3(new_n26488_), .ZN(new_n26489_));
  NOR3_X1    g24053(.A1(new_n26489_), .A2(pi0038), .A3(new_n13061_), .ZN(new_n26490_));
  NOR3_X1    g24054(.A1(new_n26490_), .A2(new_n2610_), .A3(new_n13005_), .ZN(new_n26491_));
  NOR2_X1    g24055(.A1(new_n26491_), .A2(new_n2629_), .ZN(new_n26492_));
  NAND2_X1   g24056(.A1(new_n26492_), .A2(pi0644), .ZN(new_n26493_));
  NOR2_X1    g24057(.A1(new_n2609_), .A2(new_n2629_), .ZN(new_n26494_));
  AOI21_X1   g24058(.A1(new_n13397_), .A2(pi0222), .B(new_n3265_), .ZN(new_n26495_));
  NAND2_X1   g24059(.A1(new_n13341_), .A2(pi0616), .ZN(new_n26496_));
  AOI21_X1   g24060(.A1(new_n26495_), .A2(new_n26496_), .B(new_n2610_), .ZN(new_n26497_));
  NOR2_X1    g24061(.A1(new_n13214_), .A2(new_n13111_), .ZN(new_n26498_));
  INV_X1     g24062(.I(new_n26498_), .ZN(new_n26499_));
  AOI21_X1   g24063(.A1(new_n13088_), .A2(pi0222), .B(new_n3304_), .ZN(new_n26500_));
  NAND2_X1   g24064(.A1(new_n26499_), .A2(new_n26500_), .ZN(new_n26501_));
  NAND2_X1   g24065(.A1(new_n26501_), .A2(new_n2436_), .ZN(new_n26502_));
  NOR2_X1    g24066(.A1(new_n13214_), .A2(new_n5404_), .ZN(new_n26503_));
  AOI21_X1   g24067(.A1(new_n13228_), .A2(new_n5404_), .B(new_n26503_), .ZN(new_n26504_));
  OR2_X2     g24068(.A1(new_n26504_), .A2(new_n13111_), .Z(new_n26505_));
  NOR2_X1    g24069(.A1(new_n26505_), .A2(new_n6764_), .ZN(new_n26506_));
  NOR2_X1    g24070(.A1(new_n13316_), .A2(new_n12755_), .ZN(new_n26507_));
  NAND2_X1   g24071(.A1(new_n26507_), .A2(pi0616), .ZN(new_n26508_));
  INV_X1     g24072(.I(new_n26508_), .ZN(new_n26509_));
  NOR2_X1    g24073(.A1(new_n5401_), .A2(new_n13111_), .ZN(new_n26510_));
  AOI21_X1   g24074(.A1(new_n13721_), .A2(new_n26510_), .B(new_n13117_), .ZN(new_n26511_));
  OAI21_X1   g24075(.A1(new_n26508_), .A2(new_n13163_), .B(new_n26511_), .ZN(new_n26512_));
  OAI21_X1   g24076(.A1(new_n13116_), .A2(new_n26509_), .B(new_n26512_), .ZN(new_n26513_));
  NOR2_X1    g24077(.A1(new_n26513_), .A2(new_n5422_), .ZN(new_n26514_));
  OAI21_X1   g24078(.A1(new_n26514_), .A2(new_n26506_), .B(new_n2629_), .ZN(new_n26515_));
  NAND2_X1   g24079(.A1(new_n26438_), .A2(new_n13111_), .ZN(new_n26516_));
  NAND2_X1   g24080(.A1(new_n13317_), .A2(pi0616), .ZN(new_n26517_));
  NAND3_X1   g24081(.A1(new_n26516_), .A2(new_n5401_), .A3(new_n26517_), .ZN(new_n26518_));
  NOR2_X1    g24082(.A1(new_n12755_), .A2(new_n13111_), .ZN(new_n26519_));
  INV_X1     g24083(.I(new_n26519_), .ZN(new_n26520_));
  NAND2_X1   g24084(.A1(new_n13608_), .A2(new_n26520_), .ZN(new_n26521_));
  NAND3_X1   g24085(.A1(new_n26521_), .A2(new_n13163_), .A3(new_n13309_), .ZN(new_n26522_));
  AOI21_X1   g24086(.A1(new_n26518_), .A2(new_n26522_), .B(new_n13117_), .ZN(new_n26523_));
  NAND2_X1   g24087(.A1(new_n26516_), .A2(new_n26517_), .ZN(new_n26524_));
  NOR2_X1    g24088(.A1(new_n26524_), .A2(new_n13116_), .ZN(new_n26525_));
  NOR2_X1    g24089(.A1(new_n26523_), .A2(new_n26525_), .ZN(new_n26526_));
  NOR2_X1    g24090(.A1(new_n26526_), .A2(new_n5422_), .ZN(new_n26527_));
  NOR2_X1    g24091(.A1(new_n13265_), .A2(new_n13111_), .ZN(new_n26528_));
  AOI21_X1   g24092(.A1(new_n26437_), .A2(new_n13111_), .B(new_n26528_), .ZN(new_n26529_));
  INV_X1     g24093(.I(new_n26529_), .ZN(new_n26530_));
  OAI21_X1   g24094(.A1(new_n26530_), .A2(new_n13163_), .B(new_n13116_), .ZN(new_n26531_));
  NAND2_X1   g24095(.A1(new_n13304_), .A2(new_n13163_), .ZN(new_n26532_));
  NOR2_X1    g24096(.A1(new_n26532_), .A2(new_n26519_), .ZN(new_n26533_));
  OAI22_X1   g24097(.A1(new_n26531_), .A2(new_n26533_), .B1(new_n13116_), .B2(new_n26529_), .ZN(new_n26534_));
  AND2_X2    g24098(.A1(new_n26534_), .A2(new_n5422_), .Z(new_n26535_));
  OAI21_X1   g24099(.A1(new_n26527_), .A2(new_n26535_), .B(pi0222), .ZN(new_n26536_));
  AND3_X2    g24100(.A1(new_n26536_), .A2(new_n3304_), .A3(new_n26515_), .Z(new_n26537_));
  NOR2_X1    g24101(.A1(new_n13275_), .A2(new_n13111_), .ZN(new_n26538_));
  AOI21_X1   g24102(.A1(new_n13149_), .A2(new_n13163_), .B(new_n26538_), .ZN(new_n26539_));
  NOR2_X1    g24103(.A1(new_n13171_), .A2(new_n13163_), .ZN(new_n26540_));
  INV_X1     g24104(.I(new_n26540_), .ZN(new_n26541_));
  AOI21_X1   g24105(.A1(new_n26541_), .A2(new_n26539_), .B(new_n13117_), .ZN(new_n26542_));
  NOR2_X1    g24106(.A1(new_n13466_), .A2(new_n26538_), .ZN(new_n26543_));
  INV_X1     g24107(.I(new_n26543_), .ZN(new_n26544_));
  AOI21_X1   g24108(.A1(new_n13117_), .A2(new_n26544_), .B(new_n26542_), .ZN(new_n26545_));
  NOR2_X1    g24109(.A1(new_n26545_), .A2(new_n5422_), .ZN(new_n26546_));
  NAND3_X1   g24110(.A1(new_n13150_), .A2(new_n13163_), .A3(new_n26520_), .ZN(new_n26547_));
  NOR2_X1    g24111(.A1(new_n13159_), .A2(new_n26528_), .ZN(new_n26548_));
  NAND2_X1   g24112(.A1(new_n26548_), .A2(new_n5401_), .ZN(new_n26549_));
  NAND3_X1   g24113(.A1(new_n26549_), .A2(new_n13116_), .A3(new_n26547_), .ZN(new_n26550_));
  OAI21_X1   g24114(.A1(new_n13159_), .A2(new_n26528_), .B(new_n13117_), .ZN(new_n26551_));
  AND2_X2    g24115(.A1(new_n26550_), .A2(new_n26551_), .Z(new_n26552_));
  NOR2_X1    g24116(.A1(new_n26552_), .A2(new_n6764_), .ZN(new_n26553_));
  NOR2_X1    g24117(.A1(new_n26546_), .A2(new_n26553_), .ZN(new_n26554_));
  NOR2_X1    g24118(.A1(new_n13209_), .A2(new_n5403_), .ZN(new_n26555_));
  NOR2_X1    g24119(.A1(new_n26555_), .A2(new_n26499_), .ZN(new_n26556_));
  NAND2_X1   g24120(.A1(new_n26556_), .A2(new_n2629_), .ZN(new_n26557_));
  OAI22_X1   g24121(.A1(new_n26554_), .A2(new_n2629_), .B1(new_n13218_), .B2(new_n26557_), .ZN(new_n26558_));
  AOI21_X1   g24122(.A1(new_n26558_), .A2(pi0215), .B(new_n2628_), .ZN(new_n26559_));
  OAI21_X1   g24123(.A1(new_n26537_), .A2(new_n26502_), .B(new_n26559_), .ZN(new_n26560_));
  OR2_X2     g24124(.A1(new_n26552_), .A2(new_n5445_), .Z(new_n26561_));
  OAI21_X1   g24125(.A1(new_n5446_), .A2(new_n26545_), .B(new_n26561_), .ZN(new_n26562_));
  OAI21_X1   g24126(.A1(new_n26557_), .A2(new_n13235_), .B(pi0223), .ZN(new_n26563_));
  AOI21_X1   g24127(.A1(new_n26562_), .A2(pi0222), .B(new_n26563_), .ZN(new_n26564_));
  NAND2_X1   g24128(.A1(new_n26513_), .A2(new_n5445_), .ZN(new_n26565_));
  NAND2_X1   g24129(.A1(new_n26505_), .A2(new_n5446_), .ZN(new_n26566_));
  AOI21_X1   g24130(.A1(new_n26565_), .A2(new_n26566_), .B(new_n2631_), .ZN(new_n26567_));
  NOR2_X1    g24131(.A1(new_n26498_), .A2(pi0224), .ZN(new_n26568_));
  NOR3_X1    g24132(.A1(new_n26567_), .A2(pi0222), .A3(new_n26568_), .ZN(new_n26569_));
  OAI21_X1   g24133(.A1(new_n26523_), .A2(new_n26525_), .B(new_n5445_), .ZN(new_n26570_));
  NAND2_X1   g24134(.A1(new_n26534_), .A2(new_n5446_), .ZN(new_n26571_));
  AOI21_X1   g24135(.A1(new_n26570_), .A2(new_n26571_), .B(new_n2629_), .ZN(new_n26572_));
  NOR3_X1    g24136(.A1(new_n26572_), .A2(pi0223), .A3(new_n26569_), .ZN(new_n26573_));
  OAI21_X1   g24137(.A1(new_n26573_), .A2(new_n26564_), .B(new_n2628_), .ZN(new_n26574_));
  NAND3_X1   g24138(.A1(new_n26560_), .A2(pi0039), .A3(new_n26574_), .ZN(new_n26575_));
  NAND2_X1   g24139(.A1(new_n19651_), .A2(pi0616), .ZN(new_n26576_));
  NAND2_X1   g24140(.A1(new_n13798_), .A2(pi0222), .ZN(new_n26577_));
  AOI21_X1   g24141(.A1(new_n26576_), .A2(new_n26577_), .B(pi0039), .ZN(new_n26578_));
  NAND3_X1   g24142(.A1(new_n13255_), .A2(new_n13250_), .A3(pi0222), .ZN(new_n26579_));
  AOI21_X1   g24143(.A1(new_n26578_), .A2(new_n26579_), .B(pi0038), .ZN(new_n26580_));
  NAND2_X1   g24144(.A1(new_n26575_), .A2(new_n26580_), .ZN(new_n26581_));
  AOI21_X1   g24145(.A1(new_n26581_), .A2(new_n26497_), .B(new_n26494_), .ZN(new_n26582_));
  NAND2_X1   g24146(.A1(new_n26582_), .A2(new_n12761_), .ZN(new_n26583_));
  OAI21_X1   g24147(.A1(new_n12761_), .A2(new_n26492_), .B(new_n26583_), .ZN(new_n26584_));
  NAND2_X1   g24148(.A1(new_n26584_), .A2(new_n12764_), .ZN(new_n26585_));
  NAND2_X1   g24149(.A1(new_n26492_), .A2(pi0609), .ZN(new_n26586_));
  OAI21_X1   g24150(.A1(new_n26584_), .A2(pi0609), .B(new_n26586_), .ZN(new_n26587_));
  AND2_X2    g24151(.A1(new_n26587_), .A2(new_n12770_), .Z(new_n26588_));
  NAND2_X1   g24152(.A1(new_n26492_), .A2(new_n12766_), .ZN(new_n26589_));
  OAI21_X1   g24153(.A1(new_n26584_), .A2(new_n12766_), .B(new_n26589_), .ZN(new_n26590_));
  NAND2_X1   g24154(.A1(new_n26590_), .A2(pi1155), .ZN(new_n26591_));
  NAND2_X1   g24155(.A1(new_n26591_), .A2(pi0785), .ZN(new_n26592_));
  OAI21_X1   g24156(.A1(new_n26592_), .A2(new_n26588_), .B(new_n26585_), .ZN(new_n26593_));
  NAND2_X1   g24157(.A1(new_n26492_), .A2(pi0618), .ZN(new_n26594_));
  OAI21_X1   g24158(.A1(new_n26593_), .A2(pi0618), .B(new_n26594_), .ZN(new_n26595_));
  NAND2_X1   g24159(.A1(new_n26595_), .A2(new_n12785_), .ZN(new_n26596_));
  NAND2_X1   g24160(.A1(new_n26492_), .A2(new_n12781_), .ZN(new_n26597_));
  OAI21_X1   g24161(.A1(new_n26593_), .A2(new_n12781_), .B(new_n26597_), .ZN(new_n26598_));
  AOI21_X1   g24162(.A1(new_n26598_), .A2(pi1154), .B(new_n12779_), .ZN(new_n26599_));
  AOI22_X1   g24163(.A1(new_n26599_), .A2(new_n26596_), .B1(new_n12779_), .B2(new_n26593_), .ZN(new_n26600_));
  NAND2_X1   g24164(.A1(new_n26600_), .A2(new_n12793_), .ZN(new_n26601_));
  NAND2_X1   g24165(.A1(new_n26492_), .A2(pi0619), .ZN(new_n26602_));
  AOI21_X1   g24166(.A1(new_n26601_), .A2(new_n26602_), .B(pi1159), .ZN(new_n26603_));
  INV_X1     g24167(.I(new_n26492_), .ZN(new_n26604_));
  NAND2_X1   g24168(.A1(new_n26600_), .A2(pi0619), .ZN(new_n26605_));
  OAI21_X1   g24169(.A1(pi0619), .A2(new_n26604_), .B(new_n26605_), .ZN(new_n26606_));
  NAND2_X1   g24170(.A1(new_n26606_), .A2(pi1159), .ZN(new_n26607_));
  NAND2_X1   g24171(.A1(new_n26607_), .A2(pi0789), .ZN(new_n26608_));
  OAI22_X1   g24172(.A1(new_n26608_), .A2(new_n26603_), .B1(pi0789), .B2(new_n26600_), .ZN(new_n26609_));
  NAND2_X1   g24173(.A1(new_n26492_), .A2(new_n12818_), .ZN(new_n26610_));
  OAI21_X1   g24174(.A1(new_n26609_), .A2(new_n12818_), .B(new_n26610_), .ZN(new_n26611_));
  NAND2_X1   g24175(.A1(new_n26604_), .A2(new_n12943_), .ZN(new_n26612_));
  OAI21_X1   g24176(.A1(new_n26611_), .A2(new_n12943_), .B(new_n26612_), .ZN(new_n26613_));
  NOR2_X1    g24177(.A1(new_n26613_), .A2(new_n12984_), .ZN(new_n26614_));
  AOI21_X1   g24178(.A1(new_n12984_), .A2(new_n26492_), .B(new_n26614_), .ZN(new_n26615_));
  OAI21_X1   g24179(.A1(new_n26615_), .A2(pi0644), .B(new_n26493_), .ZN(new_n26616_));
  AOI21_X1   g24180(.A1(new_n26616_), .A2(pi0715), .B(pi1160), .ZN(new_n26617_));
  NAND2_X1   g24181(.A1(new_n26492_), .A2(pi0647), .ZN(new_n26618_));
  NOR2_X1    g24182(.A1(new_n26492_), .A2(new_n12952_), .ZN(new_n26619_));
  NOR2_X1    g24183(.A1(new_n26604_), .A2(new_n12923_), .ZN(new_n26620_));
  NAND2_X1   g24184(.A1(new_n26604_), .A2(new_n12887_), .ZN(new_n26621_));
  NOR2_X1    g24185(.A1(new_n26492_), .A2(new_n12870_), .ZN(new_n26622_));
  INV_X1     g24186(.I(new_n26494_), .ZN(new_n26623_));
  OAI21_X1   g24187(.A1(new_n24931_), .A2(new_n26413_), .B(new_n26495_), .ZN(new_n26624_));
  NAND2_X1   g24188(.A1(new_n26624_), .A2(new_n2609_), .ZN(new_n26625_));
  NAND2_X1   g24189(.A1(new_n13253_), .A2(pi0665), .ZN(new_n26626_));
  INV_X1     g24190(.I(new_n26626_), .ZN(new_n26627_));
  AOI21_X1   g24191(.A1(new_n26627_), .A2(pi0222), .B(pi0299), .ZN(new_n26628_));
  NOR2_X1    g24192(.A1(new_n26413_), .A2(new_n12821_), .ZN(new_n26629_));
  INV_X1     g24193(.I(new_n26629_), .ZN(new_n26630_));
  NOR2_X1    g24194(.A1(new_n13414_), .A2(new_n26630_), .ZN(new_n26631_));
  NOR2_X1    g24195(.A1(new_n14667_), .A2(new_n2629_), .ZN(new_n26632_));
  OAI21_X1   g24196(.A1(new_n26632_), .A2(new_n26631_), .B(new_n26628_), .ZN(new_n26633_));
  AOI21_X1   g24197(.A1(new_n24501_), .A2(pi0222), .B(new_n2628_), .ZN(new_n26634_));
  NOR2_X1    g24198(.A1(new_n13411_), .A2(new_n26630_), .ZN(new_n26635_));
  NOR2_X1    g24199(.A1(new_n14655_), .A2(new_n2629_), .ZN(new_n26636_));
  OAI21_X1   g24200(.A1(new_n26636_), .A2(new_n26635_), .B(new_n26634_), .ZN(new_n26637_));
  NAND3_X1   g24201(.A1(new_n26633_), .A2(new_n26637_), .A3(new_n2627_), .ZN(new_n26638_));
  NAND2_X1   g24202(.A1(new_n13446_), .A2(pi0661), .ZN(new_n26639_));
  AOI21_X1   g24203(.A1(new_n26639_), .A2(new_n26500_), .B(pi0215), .ZN(new_n26640_));
  NAND2_X1   g24204(.A1(new_n13436_), .A2(new_n13437_), .ZN(new_n26641_));
  INV_X1     g24205(.I(new_n26641_), .ZN(new_n26642_));
  NAND2_X1   g24206(.A1(new_n26642_), .A2(new_n26629_), .ZN(new_n26643_));
  NOR2_X1    g24207(.A1(new_n26643_), .A2(new_n6764_), .ZN(new_n26644_));
  NOR4_X1    g24208(.A1(new_n13090_), .A2(new_n26413_), .A3(new_n5422_), .A4(new_n12825_), .ZN(new_n26645_));
  OAI21_X1   g24209(.A1(new_n26644_), .A2(new_n26645_), .B(new_n2629_), .ZN(new_n26646_));
  NOR2_X1    g24210(.A1(new_n5399_), .A2(pi0661), .ZN(new_n26647_));
  INV_X1     g24211(.I(new_n26647_), .ZN(new_n26648_));
  OAI22_X1   g24212(.A1(new_n13496_), .A2(new_n26413_), .B1(new_n26252_), .B2(new_n26648_), .ZN(new_n26649_));
  NAND2_X1   g24213(.A1(new_n26252_), .A2(new_n5401_), .ZN(new_n26650_));
  AND3_X2    g24214(.A1(new_n26650_), .A2(new_n13116_), .A3(new_n26532_), .Z(new_n26651_));
  NOR2_X1    g24215(.A1(new_n26651_), .A2(new_n26649_), .ZN(new_n26652_));
  NOR2_X1    g24216(.A1(new_n26652_), .A2(new_n6764_), .ZN(new_n26653_));
  NOR2_X1    g24217(.A1(new_n13481_), .A2(new_n12821_), .ZN(new_n26654_));
  AOI21_X1   g24218(.A1(new_n12821_), .A2(new_n13485_), .B(new_n26654_), .ZN(new_n26655_));
  NOR2_X1    g24219(.A1(new_n26655_), .A2(new_n26413_), .ZN(new_n26656_));
  AOI21_X1   g24220(.A1(new_n26413_), .A2(new_n14452_), .B(new_n26656_), .ZN(new_n26657_));
  AND2_X2    g24221(.A1(new_n26657_), .A2(new_n6764_), .Z(new_n26658_));
  OAI21_X1   g24222(.A1(new_n26653_), .A2(new_n26658_), .B(pi0222), .ZN(new_n26659_));
  NAND3_X1   g24223(.A1(new_n26659_), .A2(new_n3304_), .A3(new_n26646_), .ZN(new_n26660_));
  INV_X1     g24224(.I(new_n13166_), .ZN(new_n26661_));
  AOI22_X1   g24225(.A1(new_n13468_), .A2(pi0661), .B1(new_n13466_), .B2(new_n26647_), .ZN(new_n26662_));
  NAND2_X1   g24226(.A1(new_n26662_), .A2(new_n26661_), .ZN(new_n26663_));
  NAND2_X1   g24227(.A1(new_n26663_), .A2(new_n6764_), .ZN(new_n26664_));
  OAI21_X1   g24228(.A1(new_n13455_), .A2(new_n13460_), .B(new_n13472_), .ZN(new_n26665_));
  NOR2_X1    g24229(.A1(new_n26665_), .A2(new_n26413_), .ZN(new_n26666_));
  AOI21_X1   g24230(.A1(new_n13179_), .A2(new_n26413_), .B(new_n26666_), .ZN(new_n26667_));
  NAND2_X1   g24231(.A1(new_n26667_), .A2(new_n5422_), .ZN(new_n26668_));
  AOI21_X1   g24232(.A1(new_n26664_), .A2(new_n26668_), .B(new_n2629_), .ZN(new_n26669_));
  NOR3_X1    g24233(.A1(new_n13444_), .A2(pi0222), .A3(new_n26413_), .ZN(new_n26670_));
  OAI21_X1   g24234(.A1(new_n26669_), .A2(new_n26670_), .B(pi0215), .ZN(new_n26671_));
  NAND2_X1   g24235(.A1(new_n26671_), .A2(pi0299), .ZN(new_n26672_));
  AOI21_X1   g24236(.A1(new_n26660_), .A2(new_n26640_), .B(new_n26672_), .ZN(new_n26673_));
  NAND2_X1   g24237(.A1(new_n26657_), .A2(new_n5445_), .ZN(new_n26674_));
  OAI21_X1   g24238(.A1(new_n26652_), .A2(new_n5445_), .B(new_n26674_), .ZN(new_n26675_));
  NAND2_X1   g24239(.A1(new_n26675_), .A2(pi0222), .ZN(new_n26676_));
  AOI21_X1   g24240(.A1(new_n26639_), .A2(new_n2631_), .B(pi0222), .ZN(new_n26677_));
  AOI21_X1   g24241(.A1(new_n13430_), .A2(pi0661), .B(new_n5446_), .ZN(new_n26678_));
  AOI21_X1   g24242(.A1(new_n26643_), .A2(new_n5446_), .B(new_n26678_), .ZN(new_n26679_));
  OAI21_X1   g24243(.A1(new_n26679_), .A2(new_n2631_), .B(new_n26677_), .ZN(new_n26680_));
  NAND3_X1   g24244(.A1(new_n26676_), .A2(new_n2668_), .A3(new_n26680_), .ZN(new_n26681_));
  NOR2_X1    g24245(.A1(new_n13425_), .A2(new_n26413_), .ZN(new_n26682_));
  AOI21_X1   g24246(.A1(new_n26682_), .A2(new_n2629_), .B(new_n2668_), .ZN(new_n26683_));
  AOI21_X1   g24247(.A1(new_n26662_), .A2(new_n26661_), .B(new_n5446_), .ZN(new_n26684_));
  AOI21_X1   g24248(.A1(new_n5446_), .A2(new_n26667_), .B(new_n26684_), .ZN(new_n26685_));
  OAI21_X1   g24249(.A1(new_n26685_), .A2(new_n2629_), .B(new_n26683_), .ZN(new_n26686_));
  AOI21_X1   g24250(.A1(new_n26681_), .A2(new_n26686_), .B(pi0299), .ZN(new_n26687_));
  OAI21_X1   g24251(.A1(new_n26673_), .A2(new_n26687_), .B(pi0039), .ZN(new_n26688_));
  AOI21_X1   g24252(.A1(new_n26688_), .A2(new_n26638_), .B(pi0038), .ZN(new_n26689_));
  OAI21_X1   g24253(.A1(new_n26689_), .A2(new_n26625_), .B(new_n26623_), .ZN(new_n26690_));
  NAND2_X1   g24254(.A1(new_n26690_), .A2(new_n13521_), .ZN(new_n26691_));
  NAND2_X1   g24255(.A1(new_n26492_), .A2(pi0625), .ZN(new_n26692_));
  AOI21_X1   g24256(.A1(new_n26691_), .A2(new_n26692_), .B(pi1153), .ZN(new_n26693_));
  NAND2_X1   g24257(.A1(new_n26690_), .A2(pi0625), .ZN(new_n26694_));
  OAI21_X1   g24258(.A1(pi0625), .A2(new_n26604_), .B(new_n26694_), .ZN(new_n26695_));
  NAND2_X1   g24259(.A1(new_n26695_), .A2(pi1153), .ZN(new_n26696_));
  NAND2_X1   g24260(.A1(new_n26696_), .A2(pi0778), .ZN(new_n26697_));
  OAI22_X1   g24261(.A1(new_n26697_), .A2(new_n26693_), .B1(pi0778), .B2(new_n26690_), .ZN(new_n26698_));
  AOI21_X1   g24262(.A1(new_n26698_), .A2(new_n12870_), .B(new_n26622_), .ZN(new_n26699_));
  INV_X1     g24263(.I(new_n26699_), .ZN(new_n26700_));
  NAND2_X1   g24264(.A1(new_n26700_), .A2(new_n12888_), .ZN(new_n26701_));
  NAND2_X1   g24265(.A1(new_n26701_), .A2(new_n26621_), .ZN(new_n26702_));
  INV_X1     g24266(.I(new_n26702_), .ZN(new_n26703_));
  AOI21_X1   g24267(.A1(new_n26703_), .A2(new_n12923_), .B(new_n26620_), .ZN(new_n26704_));
  AOI21_X1   g24268(.A1(new_n26704_), .A2(new_n12952_), .B(new_n26619_), .ZN(new_n26705_));
  NAND2_X1   g24269(.A1(new_n26705_), .A2(new_n12741_), .ZN(new_n26706_));
  AOI21_X1   g24270(.A1(new_n26706_), .A2(new_n26618_), .B(pi1157), .ZN(new_n26707_));
  NOR2_X1    g24271(.A1(new_n26604_), .A2(pi0647), .ZN(new_n26708_));
  AOI21_X1   g24272(.A1(new_n26705_), .A2(pi0647), .B(new_n26708_), .ZN(new_n26709_));
  NOR2_X1    g24273(.A1(new_n26709_), .A2(new_n12965_), .ZN(new_n26710_));
  NOR3_X1    g24274(.A1(new_n26710_), .A2(new_n26707_), .A3(new_n12972_), .ZN(new_n26711_));
  NOR2_X1    g24275(.A1(new_n26705_), .A2(pi0787), .ZN(new_n26712_));
  NOR2_X1    g24276(.A1(new_n26711_), .A2(new_n26712_), .ZN(new_n26713_));
  OAI21_X1   g24277(.A1(new_n26713_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n26714_));
  NOR2_X1    g24278(.A1(new_n26710_), .A2(pi0630), .ZN(new_n26715_));
  NOR2_X1    g24279(.A1(new_n26707_), .A2(new_n12981_), .ZN(new_n26716_));
  OAI22_X1   g24280(.A1(new_n26613_), .A2(new_n17212_), .B1(new_n26715_), .B2(new_n26716_), .ZN(new_n26717_));
  NAND2_X1   g24281(.A1(new_n26717_), .A2(pi0787), .ZN(new_n26718_));
  NAND2_X1   g24282(.A1(new_n26611_), .A2(new_n19160_), .ZN(new_n26719_));
  NAND2_X1   g24283(.A1(new_n26704_), .A2(pi0628), .ZN(new_n26720_));
  AOI21_X1   g24284(.A1(new_n26604_), .A2(new_n12920_), .B(new_n18087_), .ZN(new_n26721_));
  AOI21_X1   g24285(.A1(new_n26604_), .A2(pi0628), .B(new_n18088_), .ZN(new_n26722_));
  NAND2_X1   g24286(.A1(new_n26704_), .A2(new_n12920_), .ZN(new_n26723_));
  AOI22_X1   g24287(.A1(new_n26720_), .A2(new_n26721_), .B1(new_n26723_), .B2(new_n26722_), .ZN(new_n26724_));
  AOI21_X1   g24288(.A1(new_n26719_), .A2(new_n26724_), .B(new_n12937_), .ZN(new_n26725_));
  NOR2_X1    g24289(.A1(new_n26604_), .A2(new_n12911_), .ZN(new_n26726_));
  AOI21_X1   g24290(.A1(new_n26703_), .A2(new_n12911_), .B(new_n26726_), .ZN(new_n26727_));
  NAND2_X1   g24291(.A1(new_n26492_), .A2(pi0626), .ZN(new_n26728_));
  OAI21_X1   g24292(.A1(new_n26609_), .A2(pi0626), .B(new_n26728_), .ZN(new_n26729_));
  NAND2_X1   g24293(.A1(new_n26492_), .A2(new_n12747_), .ZN(new_n26730_));
  OAI21_X1   g24294(.A1(new_n26609_), .A2(new_n12747_), .B(new_n26730_), .ZN(new_n26731_));
  AOI22_X1   g24295(.A1(new_n12812_), .A2(new_n26731_), .B1(new_n26729_), .B2(new_n12815_), .ZN(new_n26732_));
  OAI21_X1   g24296(.A1(new_n12906_), .A2(new_n26727_), .B(new_n26732_), .ZN(new_n26733_));
  NOR2_X1    g24297(.A1(new_n26733_), .A2(new_n12819_), .ZN(new_n26734_));
  NOR2_X1    g24298(.A1(new_n26734_), .A2(new_n15340_), .ZN(new_n26735_));
  NAND2_X1   g24299(.A1(new_n26629_), .A2(pi0616), .ZN(new_n26736_));
  OAI22_X1   g24300(.A1(new_n26736_), .A2(pi0039), .B1(pi0222), .B2(pi0616), .ZN(new_n26737_));
  NOR2_X1    g24301(.A1(new_n13568_), .A2(new_n13672_), .ZN(new_n26738_));
  NAND2_X1   g24302(.A1(new_n26738_), .A2(new_n26737_), .ZN(new_n26739_));
  NAND2_X1   g24303(.A1(new_n13397_), .A2(pi0222), .ZN(new_n26740_));
  NAND2_X1   g24304(.A1(new_n13572_), .A2(new_n13111_), .ZN(new_n26741_));
  AOI21_X1   g24305(.A1(new_n26741_), .A2(new_n26629_), .B(new_n26519_), .ZN(new_n26742_));
  OAI21_X1   g24306(.A1(new_n13397_), .A2(new_n26742_), .B(new_n26740_), .ZN(new_n26743_));
  AOI21_X1   g24307(.A1(new_n26743_), .A2(new_n26739_), .B(new_n3265_), .ZN(new_n26744_));
  NAND2_X1   g24308(.A1(new_n24501_), .A2(new_n13659_), .ZN(new_n26745_));
  OAI21_X1   g24309(.A1(new_n14554_), .A2(pi0616), .B(new_n26745_), .ZN(new_n26746_));
  AND2_X2    g24310(.A1(new_n13804_), .A2(new_n26630_), .Z(new_n26747_));
  OAI21_X1   g24311(.A1(new_n26747_), .A2(new_n26746_), .B(pi0222), .ZN(new_n26748_));
  AOI21_X1   g24312(.A1(new_n14553_), .A2(pi0616), .B(pi0222), .ZN(new_n26749_));
  OAI21_X1   g24313(.A1(new_n14652_), .A2(new_n26413_), .B(new_n26749_), .ZN(new_n26750_));
  NAND3_X1   g24314(.A1(new_n26748_), .A2(pi0299), .A3(new_n26750_), .ZN(new_n26751_));
  OAI22_X1   g24315(.A1(new_n14666_), .A2(pi0616), .B1(new_n26626_), .B2(new_n13586_), .ZN(new_n26752_));
  INV_X1     g24316(.I(new_n13806_), .ZN(new_n26753_));
  NOR2_X1    g24317(.A1(new_n26753_), .A2(new_n26629_), .ZN(new_n26754_));
  OAI21_X1   g24318(.A1(new_n26754_), .A2(new_n26752_), .B(pi0222), .ZN(new_n26755_));
  AOI21_X1   g24319(.A1(new_n14546_), .A2(pi0616), .B(pi0222), .ZN(new_n26756_));
  OAI21_X1   g24320(.A1(new_n14663_), .A2(new_n26413_), .B(new_n26756_), .ZN(new_n26757_));
  NAND3_X1   g24321(.A1(new_n26755_), .A2(new_n2628_), .A3(new_n26757_), .ZN(new_n26758_));
  AOI21_X1   g24322(.A1(new_n26758_), .A2(new_n26751_), .B(pi0039), .ZN(new_n26759_));
  NAND2_X1   g24323(.A1(new_n26498_), .A2(new_n13274_), .ZN(new_n26760_));
  NOR2_X1    g24324(.A1(new_n24647_), .A2(new_n13111_), .ZN(new_n26761_));
  INV_X1     g24325(.I(new_n26761_), .ZN(new_n26762_));
  AOI22_X1   g24326(.A1(new_n26762_), .A2(new_n26413_), .B1(new_n5404_), .B2(new_n26760_), .ZN(new_n26763_));
  AOI21_X1   g24327(.A1(new_n13781_), .A2(new_n13779_), .B(pi0616), .ZN(new_n26764_));
  AOI21_X1   g24328(.A1(new_n26761_), .A2(new_n12821_), .B(new_n26413_), .ZN(new_n26765_));
  NOR2_X1    g24329(.A1(new_n13215_), .A2(new_n13578_), .ZN(new_n26766_));
  NAND2_X1   g24330(.A1(new_n26766_), .A2(pi0616), .ZN(new_n26767_));
  NAND2_X1   g24331(.A1(new_n26767_), .A2(pi0680), .ZN(new_n26768_));
  OAI21_X1   g24332(.A1(new_n26768_), .A2(new_n26764_), .B(new_n26765_), .ZN(new_n26769_));
  NAND2_X1   g24333(.A1(new_n26769_), .A2(new_n26763_), .ZN(new_n26770_));
  NAND2_X1   g24334(.A1(new_n26770_), .A2(new_n5445_), .ZN(new_n26771_));
  AOI21_X1   g24335(.A1(new_n13774_), .A2(new_n26629_), .B(new_n26556_), .ZN(new_n26772_));
  NAND2_X1   g24336(.A1(new_n26772_), .A2(new_n5446_), .ZN(new_n26773_));
  AOI21_X1   g24337(.A1(new_n26771_), .A2(new_n26773_), .B(pi0222), .ZN(new_n26774_));
  AOI21_X1   g24338(.A1(new_n26548_), .A2(new_n12821_), .B(new_n26413_), .ZN(new_n26775_));
  NOR2_X1    g24339(.A1(new_n13665_), .A2(new_n13111_), .ZN(new_n26776_));
  NOR2_X1    g24340(.A1(new_n26776_), .A2(new_n12821_), .ZN(new_n26777_));
  NAND2_X1   g24341(.A1(new_n13708_), .A2(new_n26777_), .ZN(new_n26778_));
  OAI21_X1   g24342(.A1(new_n26548_), .A2(new_n26648_), .B(new_n26550_), .ZN(new_n26779_));
  AOI21_X1   g24343(.A1(new_n26775_), .A2(new_n26778_), .B(new_n26779_), .ZN(new_n26780_));
  INV_X1     g24344(.I(new_n26542_), .ZN(new_n26781_));
  INV_X1     g24345(.I(new_n13716_), .ZN(new_n26782_));
  AOI21_X1   g24346(.A1(new_n13653_), .A2(new_n13457_), .B(new_n13672_), .ZN(new_n26783_));
  OAI21_X1   g24347(.A1(new_n26783_), .A2(new_n13111_), .B(pi0680), .ZN(new_n26784_));
  AOI21_X1   g24348(.A1(new_n26543_), .A2(new_n12821_), .B(new_n26413_), .ZN(new_n26785_));
  OAI21_X1   g24349(.A1(new_n26782_), .A2(new_n26784_), .B(new_n26785_), .ZN(new_n26786_));
  NAND2_X1   g24350(.A1(new_n26544_), .A2(new_n26647_), .ZN(new_n26787_));
  NAND3_X1   g24351(.A1(new_n26786_), .A2(new_n26781_), .A3(new_n26787_), .ZN(new_n26788_));
  NOR2_X1    g24352(.A1(new_n26788_), .A2(new_n5446_), .ZN(new_n26789_));
  AOI21_X1   g24353(.A1(new_n26780_), .A2(new_n5446_), .B(new_n26789_), .ZN(new_n26790_));
  OAI21_X1   g24354(.A1(new_n26790_), .A2(new_n2629_), .B(pi0223), .ZN(new_n26791_));
  OAI21_X1   g24355(.A1(new_n26791_), .A2(new_n26774_), .B(new_n2628_), .ZN(new_n26792_));
  NOR2_X1    g24356(.A1(new_n13303_), .A2(new_n12751_), .ZN(new_n26793_));
  AOI21_X1   g24357(.A1(new_n13478_), .A2(new_n5398_), .B(new_n13462_), .ZN(new_n26794_));
  NOR2_X1    g24358(.A1(new_n26794_), .A2(pi0603), .ZN(new_n26795_));
  OAI22_X1   g24359(.A1(new_n26795_), .A2(new_n26793_), .B1(new_n13290_), .B2(new_n13626_), .ZN(new_n26796_));
  NAND2_X1   g24360(.A1(new_n26796_), .A2(new_n5406_), .ZN(new_n26797_));
  OAI21_X1   g24361(.A1(new_n12755_), .A2(new_n13316_), .B(new_n26794_), .ZN(new_n26798_));
  OAI21_X1   g24362(.A1(new_n5406_), .A2(new_n26798_), .B(new_n26797_), .ZN(new_n26799_));
  NAND2_X1   g24363(.A1(new_n26799_), .A2(new_n13095_), .ZN(new_n26800_));
  INV_X1     g24364(.I(new_n26798_), .ZN(new_n26801_));
  NOR2_X1    g24365(.A1(new_n26794_), .A2(new_n13672_), .ZN(new_n26802_));
  OAI21_X1   g24366(.A1(new_n26802_), .A2(new_n13111_), .B(pi0680), .ZN(new_n26803_));
  AOI21_X1   g24367(.A1(new_n26332_), .A2(new_n26801_), .B(new_n26803_), .ZN(new_n26804_));
  AND2_X2    g24368(.A1(new_n26800_), .A2(new_n26804_), .Z(new_n26805_));
  NAND2_X1   g24369(.A1(new_n26524_), .A2(new_n12821_), .ZN(new_n26806_));
  NAND2_X1   g24370(.A1(new_n26806_), .A2(pi0661), .ZN(new_n26807_));
  OAI22_X1   g24371(.A1(new_n26805_), .A2(new_n26807_), .B1(new_n26524_), .B2(new_n26648_), .ZN(new_n26808_));
  NOR2_X1    g24372(.A1(new_n26808_), .A2(new_n26523_), .ZN(new_n26809_));
  NOR2_X1    g24373(.A1(new_n26809_), .A2(new_n5446_), .ZN(new_n26810_));
  NOR2_X1    g24374(.A1(new_n26531_), .A2(new_n26533_), .ZN(new_n26811_));
  NAND2_X1   g24375(.A1(new_n13733_), .A2(new_n26777_), .ZN(new_n26812_));
  NAND2_X1   g24376(.A1(new_n26812_), .A2(pi0661), .ZN(new_n26813_));
  NOR2_X1    g24377(.A1(new_n26530_), .A2(pi0680), .ZN(new_n26814_));
  OAI22_X1   g24378(.A1(new_n26813_), .A2(new_n26814_), .B1(new_n26529_), .B2(new_n26648_), .ZN(new_n26815_));
  NOR2_X1    g24379(.A1(new_n26815_), .A2(new_n26811_), .ZN(new_n26816_));
  NOR2_X1    g24380(.A1(new_n26816_), .A2(new_n5445_), .ZN(new_n26817_));
  NOR2_X1    g24381(.A1(new_n26810_), .A2(new_n26817_), .ZN(new_n26818_));
  NAND2_X1   g24382(.A1(new_n13317_), .A2(new_n13605_), .ZN(new_n26819_));
  INV_X1     g24383(.I(new_n26819_), .ZN(new_n26820_));
  NOR2_X1    g24384(.A1(new_n26820_), .A2(new_n13758_), .ZN(new_n26821_));
  AOI21_X1   g24385(.A1(new_n13768_), .A2(new_n13609_), .B(new_n5407_), .ZN(new_n26822_));
  OAI21_X1   g24386(.A1(new_n26821_), .A2(new_n26822_), .B(new_n13111_), .ZN(new_n26823_));
  NAND2_X1   g24387(.A1(new_n13617_), .A2(new_n13603_), .ZN(new_n26824_));
  AOI21_X1   g24388(.A1(new_n26824_), .A2(pi0616), .B(new_n12821_), .ZN(new_n26825_));
  NAND2_X1   g24389(.A1(new_n26823_), .A2(new_n26825_), .ZN(new_n26826_));
  AOI21_X1   g24390(.A1(new_n26509_), .A2(new_n12821_), .B(new_n26413_), .ZN(new_n26827_));
  NAND2_X1   g24391(.A1(new_n26826_), .A2(new_n26827_), .ZN(new_n26828_));
  NAND2_X1   g24392(.A1(new_n26508_), .A2(new_n26647_), .ZN(new_n26829_));
  NAND3_X1   g24393(.A1(new_n26828_), .A2(new_n26512_), .A3(new_n26829_), .ZN(new_n26830_));
  NAND2_X1   g24394(.A1(new_n26830_), .A2(new_n5445_), .ZN(new_n26831_));
  AOI21_X1   g24395(.A1(new_n26498_), .A2(new_n12821_), .B(new_n26413_), .ZN(new_n26832_));
  NOR2_X1    g24396(.A1(new_n13761_), .A2(new_n12821_), .ZN(new_n26833_));
  INV_X1     g24397(.I(new_n26833_), .ZN(new_n26834_));
  NOR2_X1    g24398(.A1(new_n13588_), .A2(new_n13111_), .ZN(new_n26835_));
  OAI21_X1   g24399(.A1(new_n26834_), .A2(new_n26835_), .B(new_n26832_), .ZN(new_n26836_));
  AOI21_X1   g24400(.A1(new_n26498_), .A2(new_n5401_), .B(new_n13117_), .ZN(new_n26837_));
  NAND2_X1   g24401(.A1(new_n13228_), .A2(new_n26510_), .ZN(new_n26838_));
  AOI22_X1   g24402(.A1(new_n26838_), .A2(new_n26837_), .B1(new_n26499_), .B2(new_n26647_), .ZN(new_n26839_));
  NAND2_X1   g24403(.A1(new_n26836_), .A2(new_n26839_), .ZN(new_n26840_));
  NAND2_X1   g24404(.A1(new_n26840_), .A2(new_n5446_), .ZN(new_n26841_));
  AOI21_X1   g24405(.A1(new_n26831_), .A2(new_n26841_), .B(new_n2631_), .ZN(new_n26842_));
  AOI21_X1   g24406(.A1(new_n13111_), .A2(new_n13759_), .B(new_n26835_), .ZN(new_n26843_));
  NAND2_X1   g24407(.A1(new_n26843_), .A2(new_n26629_), .ZN(new_n26844_));
  OAI21_X1   g24408(.A1(new_n26499_), .A2(new_n26629_), .B(new_n26844_), .ZN(new_n26845_));
  OAI21_X1   g24409(.A1(new_n26845_), .A2(pi0224), .B(new_n2629_), .ZN(new_n26846_));
  OAI22_X1   g24410(.A1(new_n26818_), .A2(new_n2629_), .B1(new_n26842_), .B2(new_n26846_), .ZN(new_n26847_));
  AOI21_X1   g24411(.A1(new_n26847_), .A2(new_n2668_), .B(new_n26792_), .ZN(new_n26848_));
  NAND2_X1   g24412(.A1(new_n26770_), .A2(new_n6764_), .ZN(new_n26849_));
  NAND2_X1   g24413(.A1(new_n26772_), .A2(new_n5422_), .ZN(new_n26850_));
  AOI21_X1   g24414(.A1(new_n26849_), .A2(new_n26850_), .B(pi0222), .ZN(new_n26851_));
  NOR2_X1    g24415(.A1(new_n26788_), .A2(new_n5422_), .ZN(new_n26852_));
  AOI21_X1   g24416(.A1(new_n26780_), .A2(new_n5422_), .B(new_n26852_), .ZN(new_n26853_));
  OAI21_X1   g24417(.A1(new_n26853_), .A2(new_n2629_), .B(pi0215), .ZN(new_n26854_));
  OAI21_X1   g24418(.A1(new_n26854_), .A2(new_n26851_), .B(pi0299), .ZN(new_n26855_));
  NAND2_X1   g24419(.A1(new_n26830_), .A2(new_n6764_), .ZN(new_n26856_));
  NAND2_X1   g24420(.A1(new_n26840_), .A2(new_n5422_), .ZN(new_n26857_));
  AOI21_X1   g24421(.A1(new_n26856_), .A2(new_n26857_), .B(pi0222), .ZN(new_n26858_));
  NAND2_X1   g24422(.A1(new_n26816_), .A2(new_n5422_), .ZN(new_n26859_));
  NAND2_X1   g24423(.A1(new_n26809_), .A2(new_n6764_), .ZN(new_n26860_));
  AOI21_X1   g24424(.A1(new_n26860_), .A2(new_n26859_), .B(new_n2629_), .ZN(new_n26861_));
  OAI21_X1   g24425(.A1(new_n26861_), .A2(new_n26858_), .B(new_n3304_), .ZN(new_n26862_));
  OAI21_X1   g24426(.A1(new_n26519_), .A2(new_n26629_), .B(new_n26843_), .ZN(new_n26863_));
  AOI21_X1   g24427(.A1(new_n26863_), .A2(new_n26500_), .B(pi0215), .ZN(new_n26864_));
  AOI21_X1   g24428(.A1(new_n26862_), .A2(new_n26864_), .B(new_n26855_), .ZN(new_n26865_));
  NOR3_X1    g24429(.A1(new_n26848_), .A2(new_n26865_), .A3(new_n2627_), .ZN(new_n26866_));
  NOR3_X1    g24430(.A1(new_n26866_), .A2(pi0038), .A3(new_n26759_), .ZN(new_n26867_));
  OR3_X2     g24431(.A1(new_n26867_), .A2(new_n2610_), .A3(new_n26744_), .Z(new_n26868_));
  NAND2_X1   g24432(.A1(new_n26868_), .A2(new_n26623_), .ZN(new_n26869_));
  NAND2_X1   g24433(.A1(new_n26869_), .A2(new_n12758_), .ZN(new_n26870_));
  NOR2_X1    g24434(.A1(new_n26582_), .A2(new_n13521_), .ZN(new_n26871_));
  AOI21_X1   g24435(.A1(new_n26869_), .A2(new_n13521_), .B(new_n26871_), .ZN(new_n26872_));
  OAI21_X1   g24436(.A1(new_n26872_), .A2(pi1153), .B(new_n26696_), .ZN(new_n26873_));
  NOR2_X1    g24437(.A1(new_n26582_), .A2(pi0625), .ZN(new_n26874_));
  AOI21_X1   g24438(.A1(new_n26869_), .A2(pi0625), .B(new_n26874_), .ZN(new_n26875_));
  OAI21_X1   g24439(.A1(new_n26875_), .A2(new_n12841_), .B(pi0608), .ZN(new_n26876_));
  OAI22_X1   g24440(.A1(pi0608), .A2(new_n26873_), .B1(new_n26876_), .B2(new_n26693_), .ZN(new_n26877_));
  OR2_X2     g24441(.A1(new_n26877_), .A2(new_n12758_), .Z(new_n26878_));
  AOI21_X1   g24442(.A1(new_n26878_), .A2(new_n26870_), .B(pi0785), .ZN(new_n26879_));
  INV_X1     g24443(.I(new_n26588_), .ZN(new_n26880_));
  NOR2_X1    g24444(.A1(new_n26698_), .A2(pi0609), .ZN(new_n26881_));
  AOI21_X1   g24445(.A1(new_n26878_), .A2(new_n26870_), .B(new_n12766_), .ZN(new_n26882_));
  OAI21_X1   g24446(.A1(new_n26882_), .A2(new_n26881_), .B(pi1155), .ZN(new_n26883_));
  NAND3_X1   g24447(.A1(new_n26883_), .A2(pi0660), .A3(new_n26880_), .ZN(new_n26884_));
  INV_X1     g24448(.I(new_n26591_), .ZN(new_n26885_));
  AOI21_X1   g24449(.A1(new_n26878_), .A2(new_n26870_), .B(pi0609), .ZN(new_n26886_));
  NOR2_X1    g24450(.A1(new_n26698_), .A2(new_n12766_), .ZN(new_n26887_));
  OR2_X2     g24451(.A1(new_n26886_), .A2(new_n26887_), .Z(new_n26888_));
  AOI21_X1   g24452(.A1(new_n26888_), .A2(new_n12770_), .B(new_n26885_), .ZN(new_n26889_));
  AOI21_X1   g24453(.A1(new_n26889_), .A2(new_n13829_), .B(new_n12764_), .ZN(new_n26890_));
  AOI21_X1   g24454(.A1(new_n26890_), .A2(new_n26884_), .B(new_n26879_), .ZN(new_n26891_));
  OR2_X2     g24455(.A1(new_n26891_), .A2(pi0781), .Z(new_n26892_));
  NAND2_X1   g24456(.A1(new_n26596_), .A2(pi0627), .ZN(new_n26893_));
  AOI21_X1   g24457(.A1(new_n26700_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n26894_));
  NAND2_X1   g24458(.A1(new_n26891_), .A2(pi0618), .ZN(new_n26895_));
  AOI21_X1   g24459(.A1(new_n26895_), .A2(new_n26894_), .B(new_n26893_), .ZN(new_n26896_));
  NAND2_X1   g24460(.A1(new_n26598_), .A2(pi1154), .ZN(new_n26897_));
  NAND2_X1   g24461(.A1(new_n26897_), .A2(new_n12880_), .ZN(new_n26898_));
  OAI21_X1   g24462(.A1(new_n26699_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n26899_));
  AOI21_X1   g24463(.A1(new_n26891_), .A2(new_n12781_), .B(new_n26899_), .ZN(new_n26900_));
  OAI21_X1   g24464(.A1(new_n26900_), .A2(new_n26898_), .B(pi0781), .ZN(new_n26901_));
  OAI21_X1   g24465(.A1(new_n26901_), .A2(new_n26896_), .B(new_n26892_), .ZN(new_n26902_));
  AOI22_X1   g24466(.A1(new_n26733_), .A2(pi0788), .B1(new_n12796_), .B2(new_n26902_), .ZN(new_n26903_));
  INV_X1     g24467(.I(new_n26607_), .ZN(new_n26904_));
  NAND2_X1   g24468(.A1(new_n26902_), .A2(new_n12793_), .ZN(new_n26905_));
  NAND2_X1   g24469(.A1(new_n26703_), .A2(pi0619), .ZN(new_n26906_));
  AOI21_X1   g24470(.A1(new_n26905_), .A2(new_n26906_), .B(pi1159), .ZN(new_n26907_));
  NOR3_X1    g24471(.A1(new_n26907_), .A2(pi0648), .A3(new_n26904_), .ZN(new_n26908_));
  NOR2_X1    g24472(.A1(new_n26702_), .A2(pi0619), .ZN(new_n26909_));
  AOI21_X1   g24473(.A1(new_n26902_), .A2(pi0619), .B(new_n26909_), .ZN(new_n26910_));
  OAI21_X1   g24474(.A1(new_n26910_), .A2(new_n12791_), .B(pi0648), .ZN(new_n26911_));
  OAI21_X1   g24475(.A1(new_n26911_), .A2(new_n26603_), .B(pi0789), .ZN(new_n26912_));
  OAI21_X1   g24476(.A1(new_n26912_), .A2(new_n26908_), .B(new_n26903_), .ZN(new_n26913_));
  AOI21_X1   g24477(.A1(new_n26913_), .A2(new_n26735_), .B(new_n26725_), .ZN(new_n26914_));
  OAI21_X1   g24478(.A1(new_n26914_), .A2(new_n15341_), .B(new_n26718_), .ZN(new_n26915_));
  NOR2_X1    g24479(.A1(new_n26915_), .A2(pi0644), .ZN(new_n26916_));
  OAI21_X1   g24480(.A1(new_n26916_), .A2(new_n26714_), .B(new_n26617_), .ZN(new_n26917_));
  NAND2_X1   g24481(.A1(new_n26492_), .A2(new_n12975_), .ZN(new_n26918_));
  OAI21_X1   g24482(.A1(new_n26615_), .A2(new_n12975_), .B(new_n26918_), .ZN(new_n26919_));
  AOI21_X1   g24483(.A1(new_n26919_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n26920_));
  NOR2_X1    g24484(.A1(new_n26713_), .A2(pi0644), .ZN(new_n26921_));
  NOR2_X1    g24485(.A1(new_n26921_), .A2(new_n12740_), .ZN(new_n26922_));
  OAI21_X1   g24486(.A1(new_n26915_), .A2(new_n12975_), .B(new_n26922_), .ZN(new_n26923_));
  AOI21_X1   g24487(.A1(new_n26923_), .A2(new_n26920_), .B(new_n13000_), .ZN(new_n26924_));
  AND2_X2    g24488(.A1(new_n26915_), .A2(new_n13000_), .Z(new_n26925_));
  AOI21_X1   g24489(.A1(new_n26924_), .A2(new_n26917_), .B(new_n26925_), .ZN(new_n26926_));
  OAI21_X1   g24490(.A1(new_n26926_), .A2(po1038), .B(new_n26486_), .ZN(po0379));
  NAND2_X1   g24491(.A1(po1038), .A2(pi0223), .ZN(new_n26928_));
  NOR2_X1    g24492(.A1(new_n16040_), .A2(pi0299), .ZN(new_n26929_));
  NOR3_X1    g24493(.A1(new_n13178_), .A2(new_n2627_), .A3(new_n26929_), .ZN(new_n26930_));
  NAND2_X1   g24494(.A1(new_n13336_), .A2(new_n11503_), .ZN(new_n26931_));
  OAI21_X1   g24495(.A1(new_n26931_), .A2(new_n26930_), .B(new_n14460_), .ZN(new_n26932_));
  NAND2_X1   g24496(.A1(new_n26932_), .A2(pi0223), .ZN(new_n26933_));
  NOR2_X1    g24497(.A1(new_n26933_), .A2(new_n12766_), .ZN(new_n26934_));
  INV_X1     g24498(.I(new_n26933_), .ZN(new_n26935_));
  NOR2_X1    g24499(.A1(new_n2609_), .A2(new_n2668_), .ZN(new_n26936_));
  AOI21_X1   g24500(.A1(pi0039), .A2(pi0223), .B(new_n3265_), .ZN(new_n26937_));
  INV_X1     g24501(.I(new_n26937_), .ZN(new_n26938_));
  AOI21_X1   g24502(.A1(new_n13568_), .A2(new_n2668_), .B(pi0039), .ZN(new_n26939_));
  NOR2_X1    g24503(.A1(new_n12755_), .A2(new_n5406_), .ZN(new_n26940_));
  NOR2_X1    g24504(.A1(new_n13568_), .A2(new_n26940_), .ZN(new_n26941_));
  INV_X1     g24505(.I(new_n26941_), .ZN(new_n26942_));
  AOI21_X1   g24506(.A1(new_n26942_), .A2(new_n26939_), .B(new_n26938_), .ZN(new_n26943_));
  INV_X1     g24507(.I(new_n26943_), .ZN(new_n26944_));
  NOR2_X1    g24508(.A1(new_n14666_), .A2(new_n5406_), .ZN(new_n26945_));
  AOI21_X1   g24509(.A1(new_n26945_), .A2(new_n2668_), .B(pi0299), .ZN(new_n26946_));
  OAI21_X1   g24510(.A1(new_n14666_), .A2(pi0642), .B(pi0223), .ZN(new_n26947_));
  OAI21_X1   g24511(.A1(new_n14547_), .A2(new_n26947_), .B(new_n26946_), .ZN(new_n26948_));
  NOR2_X1    g24512(.A1(new_n14554_), .A2(new_n5406_), .ZN(new_n26949_));
  AOI21_X1   g24513(.A1(new_n26949_), .A2(new_n2668_), .B(new_n2628_), .ZN(new_n26950_));
  NAND3_X1   g24514(.A1(new_n24841_), .A2(pi0603), .A3(new_n5406_), .ZN(new_n26951_));
  NAND3_X1   g24515(.A1(new_n14559_), .A2(new_n26951_), .A3(pi0223), .ZN(new_n26952_));
  AOI21_X1   g24516(.A1(new_n26950_), .A2(new_n26952_), .B(pi0039), .ZN(new_n26953_));
  AOI21_X1   g24517(.A1(new_n26948_), .A2(new_n26953_), .B(pi0038), .ZN(new_n26954_));
  INV_X1     g24518(.I(new_n5402_), .ZN(new_n26955_));
  NOR3_X1    g24519(.A1(new_n26116_), .A2(new_n26955_), .A3(new_n26942_), .ZN(new_n26956_));
  OAI21_X1   g24520(.A1(new_n5406_), .A2(new_n13265_), .B(new_n26548_), .ZN(new_n26957_));
  NOR2_X1    g24521(.A1(new_n13104_), .A2(new_n26940_), .ZN(new_n26958_));
  INV_X1     g24522(.I(new_n26958_), .ZN(new_n26959_));
  NAND2_X1   g24523(.A1(new_n26957_), .A2(new_n26959_), .ZN(new_n26960_));
  AOI22_X1   g24524(.A1(new_n26960_), .A2(new_n5403_), .B1(new_n5399_), .B2(new_n26956_), .ZN(new_n26961_));
  AND2_X2    g24525(.A1(new_n26961_), .A2(new_n5446_), .Z(new_n26962_));
  NOR2_X1    g24526(.A1(new_n13277_), .A2(new_n5406_), .ZN(new_n26963_));
  AOI21_X1   g24527(.A1(new_n13171_), .A2(new_n5406_), .B(new_n26963_), .ZN(new_n26964_));
  NOR2_X1    g24528(.A1(new_n13275_), .A2(new_n5406_), .ZN(new_n26965_));
  NOR3_X1    g24529(.A1(new_n13149_), .A2(new_n26955_), .A3(new_n26965_), .ZN(new_n26966_));
  INV_X1     g24530(.I(new_n26966_), .ZN(new_n26967_));
  OAI22_X1   g24531(.A1(new_n26964_), .A2(new_n5404_), .B1(pi0681), .B2(new_n26967_), .ZN(new_n26968_));
  NOR2_X1    g24532(.A1(new_n26968_), .A2(new_n5446_), .ZN(new_n26969_));
  OAI21_X1   g24533(.A1(new_n26962_), .A2(new_n26969_), .B(pi0223), .ZN(new_n26970_));
  NAND2_X1   g24534(.A1(new_n13210_), .A2(pi0642), .ZN(new_n26971_));
  AOI21_X1   g24535(.A1(new_n26971_), .A2(new_n2641_), .B(pi0223), .ZN(new_n26972_));
  NOR2_X1    g24536(.A1(new_n26955_), .A2(new_n5406_), .ZN(new_n26973_));
  NAND2_X1   g24537(.A1(new_n13721_), .A2(new_n26973_), .ZN(new_n26974_));
  NOR3_X1    g24538(.A1(new_n13316_), .A2(new_n5406_), .A3(new_n12755_), .ZN(new_n26975_));
  NAND2_X1   g24539(.A1(new_n26975_), .A2(new_n26955_), .ZN(new_n26976_));
  AND3_X2    g24540(.A1(new_n26976_), .A2(new_n5399_), .A3(new_n26974_), .Z(new_n26977_));
  NOR2_X1    g24541(.A1(new_n26975_), .A2(new_n5399_), .ZN(new_n26978_));
  NOR2_X1    g24542(.A1(new_n26977_), .A2(new_n26978_), .ZN(new_n26979_));
  NOR2_X1    g24543(.A1(new_n26979_), .A2(new_n5446_), .ZN(new_n26980_));
  INV_X1     g24544(.I(new_n26971_), .ZN(new_n26981_));
  INV_X1     g24545(.I(new_n26973_), .ZN(new_n26982_));
  OAI21_X1   g24546(.A1(new_n26971_), .A2(new_n5402_), .B(new_n5399_), .ZN(new_n26983_));
  INV_X1     g24547(.I(new_n26983_), .ZN(new_n26984_));
  OAI21_X1   g24548(.A1(new_n13642_), .A2(new_n26982_), .B(new_n26984_), .ZN(new_n26985_));
  OAI21_X1   g24549(.A1(new_n5399_), .A2(new_n26981_), .B(new_n26985_), .ZN(new_n26986_));
  AOI21_X1   g24550(.A1(new_n5446_), .A2(new_n26986_), .B(new_n26980_), .ZN(new_n26987_));
  OAI21_X1   g24551(.A1(new_n26987_), .A2(new_n2641_), .B(new_n26972_), .ZN(new_n26988_));
  NAND3_X1   g24552(.A1(new_n26988_), .A2(new_n2628_), .A3(new_n26970_), .ZN(new_n26989_));
  AOI21_X1   g24553(.A1(new_n13088_), .A2(pi0223), .B(new_n3304_), .ZN(new_n26990_));
  AOI21_X1   g24554(.A1(new_n26971_), .A2(new_n26990_), .B(pi0215), .ZN(new_n26991_));
  INV_X1     g24555(.I(new_n15979_), .ZN(new_n26992_));
  OAI21_X1   g24556(.A1(pi0947), .A2(new_n26992_), .B(new_n26979_), .ZN(new_n26993_));
  OR3_X2     g24557(.A1(new_n26986_), .A2(pi0947), .A3(new_n26992_), .Z(new_n26994_));
  AOI21_X1   g24558(.A1(new_n26993_), .A2(new_n26994_), .B(pi0223), .ZN(new_n26995_));
  OAI21_X1   g24559(.A1(new_n13083_), .A2(new_n26940_), .B(new_n5399_), .ZN(new_n26996_));
  NOR2_X1    g24560(.A1(new_n13090_), .A2(pi0642), .ZN(new_n26997_));
  AOI21_X1   g24561(.A1(new_n13317_), .A2(pi0642), .B(new_n26997_), .ZN(new_n26998_));
  NOR2_X1    g24562(.A1(new_n26998_), .A2(new_n5402_), .ZN(new_n26999_));
  OAI21_X1   g24563(.A1(new_n26999_), .A2(new_n26996_), .B(new_n6764_), .ZN(new_n27000_));
  NAND2_X1   g24564(.A1(new_n26998_), .A2(pi0681), .ZN(new_n27001_));
  INV_X1     g24565(.I(new_n27001_), .ZN(new_n27002_));
  OAI21_X1   g24566(.A1(new_n27000_), .A2(new_n27002_), .B(pi0223), .ZN(new_n27003_));
  NOR2_X1    g24567(.A1(new_n13730_), .A2(pi0642), .ZN(new_n27004_));
  NOR2_X1    g24568(.A1(new_n13284_), .A2(new_n5406_), .ZN(new_n27005_));
  OAI21_X1   g24569(.A1(new_n27004_), .A2(new_n27005_), .B(new_n13095_), .ZN(new_n27006_));
  NAND2_X1   g24570(.A1(new_n27006_), .A2(new_n26959_), .ZN(new_n27007_));
  NOR2_X1    g24571(.A1(new_n27007_), .A2(new_n5399_), .ZN(new_n27008_));
  NAND3_X1   g24572(.A1(new_n13292_), .A2(pi0603), .A3(pi0642), .ZN(new_n27009_));
  AOI21_X1   g24573(.A1(new_n27009_), .A2(new_n13304_), .B(new_n26955_), .ZN(new_n27010_));
  NOR2_X1    g24574(.A1(new_n27007_), .A2(new_n5402_), .ZN(new_n27011_));
  OAI21_X1   g24575(.A1(new_n27011_), .A2(new_n27010_), .B(new_n5399_), .ZN(new_n27012_));
  NAND2_X1   g24576(.A1(new_n27012_), .A2(new_n5422_), .ZN(new_n27013_));
  NOR2_X1    g24577(.A1(new_n27013_), .A2(new_n27008_), .ZN(new_n27014_));
  OAI21_X1   g24578(.A1(new_n27014_), .A2(new_n27003_), .B(new_n3304_), .ZN(new_n27015_));
  OAI21_X1   g24579(.A1(new_n27015_), .A2(new_n26995_), .B(new_n26991_), .ZN(new_n27016_));
  NOR2_X1    g24580(.A1(new_n26968_), .A2(new_n5422_), .ZN(new_n27017_));
  AOI21_X1   g24581(.A1(new_n26961_), .A2(new_n5422_), .B(new_n27017_), .ZN(new_n27018_));
  NOR2_X1    g24582(.A1(new_n13211_), .A2(new_n26982_), .ZN(new_n27019_));
  NOR2_X1    g24583(.A1(new_n27019_), .A2(new_n26983_), .ZN(new_n27020_));
  NOR2_X1    g24584(.A1(new_n26966_), .A2(pi0681), .ZN(new_n27021_));
  AOI21_X1   g24585(.A1(new_n13170_), .A2(new_n27021_), .B(new_n27020_), .ZN(new_n27022_));
  NOR2_X1    g24586(.A1(new_n24647_), .A2(new_n5406_), .ZN(new_n27023_));
  OAI21_X1   g24587(.A1(new_n5399_), .A2(new_n27023_), .B(new_n27022_), .ZN(new_n27024_));
  OR2_X2     g24588(.A1(new_n27024_), .A2(new_n15979_), .Z(new_n27025_));
  NOR2_X1    g24589(.A1(new_n27020_), .A2(new_n6764_), .ZN(new_n27026_));
  NAND2_X1   g24590(.A1(new_n27026_), .A2(new_n26981_), .ZN(new_n27027_));
  NAND3_X1   g24591(.A1(new_n27025_), .A2(new_n5692_), .A3(new_n27027_), .ZN(new_n27028_));
  AOI21_X1   g24592(.A1(new_n27024_), .A2(pi0947), .B(pi0223), .ZN(new_n27029_));
  NAND2_X1   g24593(.A1(new_n27028_), .A2(new_n27029_), .ZN(new_n27030_));
  OAI21_X1   g24594(.A1(new_n27018_), .A2(new_n2668_), .B(new_n27030_), .ZN(new_n27031_));
  NAND2_X1   g24595(.A1(new_n27031_), .A2(pi0215), .ZN(new_n27032_));
  NAND3_X1   g24596(.A1(new_n27032_), .A2(pi0299), .A3(new_n27016_), .ZN(new_n27033_));
  NAND3_X1   g24597(.A1(new_n27033_), .A2(pi0039), .A3(new_n26989_), .ZN(new_n27034_));
  AOI21_X1   g24598(.A1(new_n27034_), .A2(new_n26954_), .B(new_n2610_), .ZN(new_n27035_));
  AOI21_X1   g24599(.A1(new_n27035_), .A2(new_n26944_), .B(new_n26936_), .ZN(new_n27036_));
  NOR2_X1    g24600(.A1(new_n27036_), .A2(new_n12760_), .ZN(new_n27037_));
  AOI21_X1   g24601(.A1(new_n12760_), .A2(new_n26935_), .B(new_n27037_), .ZN(new_n27038_));
  NOR2_X1    g24602(.A1(new_n27038_), .A2(pi0609), .ZN(new_n27039_));
  OAI21_X1   g24603(.A1(new_n27039_), .A2(new_n26934_), .B(new_n12770_), .ZN(new_n27040_));
  NOR2_X1    g24604(.A1(new_n27038_), .A2(new_n12766_), .ZN(new_n27041_));
  NOR2_X1    g24605(.A1(new_n26933_), .A2(pi0609), .ZN(new_n27042_));
  OAI21_X1   g24606(.A1(new_n27041_), .A2(new_n27042_), .B(pi1155), .ZN(new_n27043_));
  NAND3_X1   g24607(.A1(new_n27040_), .A2(new_n27043_), .A3(pi0785), .ZN(new_n27044_));
  NAND2_X1   g24608(.A1(new_n27038_), .A2(new_n12764_), .ZN(new_n27045_));
  NAND2_X1   g24609(.A1(new_n27044_), .A2(new_n27045_), .ZN(new_n27046_));
  NAND2_X1   g24610(.A1(new_n27046_), .A2(new_n12779_), .ZN(new_n27047_));
  NAND2_X1   g24611(.A1(new_n26935_), .A2(pi0618), .ZN(new_n27048_));
  OAI21_X1   g24612(.A1(new_n27046_), .A2(pi0618), .B(new_n27048_), .ZN(new_n27049_));
  NAND2_X1   g24613(.A1(new_n27049_), .A2(new_n12785_), .ZN(new_n27050_));
  NOR2_X1    g24614(.A1(new_n27046_), .A2(new_n12781_), .ZN(new_n27051_));
  AOI21_X1   g24615(.A1(new_n12781_), .A2(new_n26935_), .B(new_n27051_), .ZN(new_n27052_));
  NOR2_X1    g24616(.A1(new_n27052_), .A2(new_n12785_), .ZN(new_n27053_));
  NOR2_X1    g24617(.A1(new_n27053_), .A2(new_n12779_), .ZN(new_n27054_));
  NAND2_X1   g24618(.A1(new_n27054_), .A2(new_n27050_), .ZN(new_n27055_));
  NAND2_X1   g24619(.A1(new_n27055_), .A2(new_n27047_), .ZN(new_n27056_));
  INV_X1     g24620(.I(new_n27056_), .ZN(new_n27057_));
  NOR2_X1    g24621(.A1(new_n27056_), .A2(pi0619), .ZN(new_n27058_));
  NOR2_X1    g24622(.A1(new_n26933_), .A2(new_n12793_), .ZN(new_n27059_));
  OAI21_X1   g24623(.A1(new_n27058_), .A2(new_n27059_), .B(new_n12791_), .ZN(new_n27060_));
  INV_X1     g24624(.I(new_n27060_), .ZN(new_n27061_));
  NOR2_X1    g24625(.A1(new_n27056_), .A2(new_n12793_), .ZN(new_n27062_));
  NOR2_X1    g24626(.A1(new_n26933_), .A2(pi0619), .ZN(new_n27063_));
  OAI21_X1   g24627(.A1(new_n27062_), .A2(new_n27063_), .B(pi1159), .ZN(new_n27064_));
  NAND2_X1   g24628(.A1(new_n27064_), .A2(pi0789), .ZN(new_n27065_));
  OAI22_X1   g24629(.A1(new_n27065_), .A2(new_n27061_), .B1(pi0789), .B2(new_n27057_), .ZN(new_n27066_));
  NAND2_X1   g24630(.A1(new_n26935_), .A2(new_n12818_), .ZN(new_n27067_));
  OAI21_X1   g24631(.A1(new_n27066_), .A2(new_n12818_), .B(new_n27067_), .ZN(new_n27068_));
  NAND2_X1   g24632(.A1(new_n26933_), .A2(new_n12943_), .ZN(new_n27069_));
  OAI21_X1   g24633(.A1(new_n27068_), .A2(new_n12943_), .B(new_n27069_), .ZN(new_n27070_));
  NOR2_X1    g24634(.A1(new_n26933_), .A2(new_n12923_), .ZN(new_n27071_));
  OAI21_X1   g24635(.A1(new_n13344_), .A2(new_n2668_), .B(pi0038), .ZN(new_n27072_));
  AOI21_X1   g24636(.A1(new_n13398_), .A2(pi0681), .B(new_n27072_), .ZN(new_n27073_));
  OAI21_X1   g24637(.A1(new_n26626_), .A2(new_n2668_), .B(new_n2628_), .ZN(new_n27074_));
  NOR2_X1    g24638(.A1(new_n12821_), .A2(new_n5399_), .ZN(new_n27075_));
  NAND2_X1   g24639(.A1(new_n14667_), .A2(new_n27075_), .ZN(new_n27076_));
  NAND2_X1   g24640(.A1(new_n13414_), .A2(pi0223), .ZN(new_n27077_));
  AOI21_X1   g24641(.A1(new_n27076_), .A2(new_n27077_), .B(new_n27074_), .ZN(new_n27078_));
  NAND2_X1   g24642(.A1(new_n24501_), .A2(pi0223), .ZN(new_n27079_));
  NAND2_X1   g24643(.A1(new_n27079_), .A2(pi0299), .ZN(new_n27080_));
  NAND2_X1   g24644(.A1(new_n14655_), .A2(new_n27075_), .ZN(new_n27081_));
  NAND2_X1   g24645(.A1(new_n13411_), .A2(pi0223), .ZN(new_n27082_));
  AOI21_X1   g24646(.A1(new_n27081_), .A2(new_n27082_), .B(new_n27080_), .ZN(new_n27083_));
  OR3_X2     g24647(.A1(new_n27083_), .A2(pi0039), .A3(new_n27078_), .Z(new_n27084_));
  NOR2_X1    g24648(.A1(new_n13091_), .A2(pi0681), .ZN(new_n27085_));
  NOR2_X1    g24649(.A1(new_n27085_), .A2(new_n5422_), .ZN(new_n27086_));
  NAND2_X1   g24650(.A1(new_n26655_), .A2(pi0681), .ZN(new_n27087_));
  AOI21_X1   g24651(.A1(new_n27087_), .A2(new_n27086_), .B(new_n2668_), .ZN(new_n27088_));
  NAND2_X1   g24652(.A1(new_n13125_), .A2(new_n13115_), .ZN(new_n27089_));
  INV_X1     g24653(.I(new_n13496_), .ZN(new_n27090_));
  NAND2_X1   g24654(.A1(new_n27090_), .A2(pi0681), .ZN(new_n27091_));
  NAND3_X1   g24655(.A1(new_n27091_), .A2(new_n5422_), .A3(new_n27089_), .ZN(new_n27092_));
  INV_X1     g24656(.I(new_n27075_), .ZN(new_n27093_));
  NOR2_X1    g24657(.A1(new_n26641_), .A2(new_n27093_), .ZN(new_n27094_));
  NAND2_X1   g24658(.A1(new_n27094_), .A2(new_n5422_), .ZN(new_n27095_));
  NAND3_X1   g24659(.A1(new_n13430_), .A2(pi0681), .A3(new_n6764_), .ZN(new_n27096_));
  NAND2_X1   g24660(.A1(new_n27095_), .A2(new_n27096_), .ZN(new_n27097_));
  AOI22_X1   g24661(.A1(new_n27092_), .A2(new_n27088_), .B1(new_n2668_), .B2(new_n27097_), .ZN(new_n27098_));
  NAND2_X1   g24662(.A1(new_n13446_), .A2(pi0681), .ZN(new_n27099_));
  AOI22_X1   g24663(.A1(new_n27098_), .A2(new_n3304_), .B1(new_n26990_), .B2(new_n27099_), .ZN(new_n27100_));
  NOR2_X1    g24664(.A1(new_n5399_), .A2(pi0223), .ZN(new_n27101_));
  AOI21_X1   g24665(.A1(new_n13443_), .A2(new_n27101_), .B(new_n2436_), .ZN(new_n27102_));
  NOR2_X1    g24666(.A1(new_n13171_), .A2(new_n26413_), .ZN(new_n27103_));
  INV_X1     g24667(.I(new_n27103_), .ZN(new_n27104_));
  NAND2_X1   g24668(.A1(new_n13165_), .A2(new_n13164_), .ZN(new_n27105_));
  NAND2_X1   g24669(.A1(new_n27105_), .A2(new_n26413_), .ZN(new_n27106_));
  AOI21_X1   g24670(.A1(new_n27106_), .A2(new_n27104_), .B(pi0681), .ZN(new_n27107_));
  AOI21_X1   g24671(.A1(pi0681), .A2(new_n13468_), .B(new_n27107_), .ZN(new_n27108_));
  NOR2_X1    g24672(.A1(new_n27108_), .A2(new_n5422_), .ZN(new_n27109_));
  AOI21_X1   g24673(.A1(new_n26665_), .A2(pi0681), .B(new_n13161_), .ZN(new_n27110_));
  NOR2_X1    g24674(.A1(new_n27110_), .A2(new_n6764_), .ZN(new_n27111_));
  OAI21_X1   g24675(.A1(new_n27109_), .A2(new_n27111_), .B(pi0223), .ZN(new_n27112_));
  AOI21_X1   g24676(.A1(new_n27112_), .A2(new_n27102_), .B(new_n2628_), .ZN(new_n27113_));
  OAI21_X1   g24677(.A1(new_n27100_), .A2(pi0215), .B(new_n27113_), .ZN(new_n27114_));
  AND2_X2    g24678(.A1(new_n27110_), .A2(new_n5446_), .Z(new_n27115_));
  AND2_X2    g24679(.A1(new_n27108_), .A2(new_n5445_), .Z(new_n27116_));
  OAI21_X1   g24680(.A1(new_n27116_), .A2(new_n27115_), .B(pi0223), .ZN(new_n27117_));
  NOR2_X1    g24681(.A1(new_n27094_), .A2(new_n5445_), .ZN(new_n27118_));
  AOI21_X1   g24682(.A1(new_n13430_), .A2(pi0681), .B(new_n5446_), .ZN(new_n27119_));
  OAI21_X1   g24683(.A1(new_n27118_), .A2(new_n27119_), .B(new_n2642_), .ZN(new_n27120_));
  NAND2_X1   g24684(.A1(new_n27099_), .A2(new_n2641_), .ZN(new_n27121_));
  NAND2_X1   g24685(.A1(new_n27120_), .A2(new_n27121_), .ZN(new_n27122_));
  AOI21_X1   g24686(.A1(new_n27122_), .A2(new_n2668_), .B(pi0299), .ZN(new_n27123_));
  AOI21_X1   g24687(.A1(new_n27117_), .A2(new_n27123_), .B(new_n2627_), .ZN(new_n27124_));
  NAND2_X1   g24688(.A1(new_n27114_), .A2(new_n27124_), .ZN(new_n27125_));
  AOI21_X1   g24689(.A1(new_n27125_), .A2(new_n27084_), .B(pi0038), .ZN(new_n27126_));
  NOR3_X1    g24690(.A1(new_n27126_), .A2(new_n2610_), .A3(new_n27073_), .ZN(new_n27127_));
  NOR2_X1    g24691(.A1(new_n27127_), .A2(new_n26936_), .ZN(new_n27128_));
  INV_X1     g24692(.I(new_n27128_), .ZN(new_n27129_));
  NOR2_X1    g24693(.A1(new_n27128_), .A2(pi0625), .ZN(new_n27130_));
  NOR2_X1    g24694(.A1(new_n26933_), .A2(new_n13521_), .ZN(new_n27131_));
  OAI21_X1   g24695(.A1(new_n27130_), .A2(new_n27131_), .B(new_n12841_), .ZN(new_n27132_));
  NOR2_X1    g24696(.A1(new_n27128_), .A2(new_n13521_), .ZN(new_n27133_));
  NOR2_X1    g24697(.A1(new_n26933_), .A2(pi0625), .ZN(new_n27134_));
  OAI21_X1   g24698(.A1(new_n27133_), .A2(new_n27134_), .B(pi1153), .ZN(new_n27135_));
  NAND3_X1   g24699(.A1(new_n27132_), .A2(new_n27135_), .A3(pi0778), .ZN(new_n27136_));
  OAI21_X1   g24700(.A1(pi0778), .A2(new_n27129_), .B(new_n27136_), .ZN(new_n27137_));
  INV_X1     g24701(.I(new_n27137_), .ZN(new_n27138_));
  NOR2_X1    g24702(.A1(new_n26933_), .A2(new_n12870_), .ZN(new_n27139_));
  AOI21_X1   g24703(.A1(new_n27138_), .A2(new_n12870_), .B(new_n27139_), .ZN(new_n27140_));
  AND2_X2    g24704(.A1(new_n27140_), .A2(new_n12888_), .Z(new_n27141_));
  NOR2_X1    g24705(.A1(new_n26935_), .A2(new_n12888_), .ZN(new_n27142_));
  NOR2_X1    g24706(.A1(new_n27141_), .A2(new_n27142_), .ZN(new_n27143_));
  AOI21_X1   g24707(.A1(new_n27143_), .A2(new_n12923_), .B(new_n27071_), .ZN(new_n27144_));
  INV_X1     g24708(.I(new_n27144_), .ZN(new_n27145_));
  NOR2_X1    g24709(.A1(new_n27145_), .A2(new_n12951_), .ZN(new_n27146_));
  AOI21_X1   g24710(.A1(new_n12951_), .A2(new_n26933_), .B(new_n27146_), .ZN(new_n27147_));
  NAND2_X1   g24711(.A1(new_n27147_), .A2(pi0647), .ZN(new_n27148_));
  NAND2_X1   g24712(.A1(new_n26935_), .A2(new_n12741_), .ZN(new_n27149_));
  AOI21_X1   g24713(.A1(new_n27148_), .A2(new_n27149_), .B(new_n12965_), .ZN(new_n27150_));
  NOR2_X1    g24714(.A1(new_n26933_), .A2(new_n12741_), .ZN(new_n27151_));
  INV_X1     g24715(.I(new_n27147_), .ZN(new_n27152_));
  NOR2_X1    g24716(.A1(new_n27152_), .A2(pi0647), .ZN(new_n27153_));
  OAI21_X1   g24717(.A1(new_n27153_), .A2(new_n27151_), .B(new_n12965_), .ZN(new_n27154_));
  NAND2_X1   g24718(.A1(new_n27154_), .A2(pi0630), .ZN(new_n27155_));
  OAI21_X1   g24719(.A1(pi0630), .A2(new_n27150_), .B(new_n27155_), .ZN(new_n27156_));
  OAI21_X1   g24720(.A1(new_n27070_), .A2(new_n17212_), .B(new_n27156_), .ZN(new_n27157_));
  NAND2_X1   g24721(.A1(new_n27157_), .A2(pi0787), .ZN(new_n27158_));
  NOR2_X1    g24722(.A1(new_n27145_), .A2(new_n12920_), .ZN(new_n27159_));
  INV_X1     g24723(.I(new_n27159_), .ZN(new_n27160_));
  AOI21_X1   g24724(.A1(new_n26933_), .A2(new_n12920_), .B(new_n18087_), .ZN(new_n27161_));
  AOI21_X1   g24725(.A1(new_n26933_), .A2(pi0628), .B(new_n18088_), .ZN(new_n27162_));
  NOR2_X1    g24726(.A1(new_n27145_), .A2(pi0628), .ZN(new_n27163_));
  INV_X1     g24727(.I(new_n27163_), .ZN(new_n27164_));
  AOI22_X1   g24728(.A1(new_n27160_), .A2(new_n27161_), .B1(new_n27164_), .B2(new_n27162_), .ZN(new_n27165_));
  INV_X1     g24729(.I(new_n27165_), .ZN(new_n27166_));
  AOI21_X1   g24730(.A1(new_n27068_), .A2(new_n19160_), .B(new_n27166_), .ZN(new_n27167_));
  NAND2_X1   g24731(.A1(new_n27167_), .A2(new_n15340_), .ZN(new_n27168_));
  NAND2_X1   g24732(.A1(new_n27168_), .A2(new_n15693_), .ZN(new_n27169_));
  NOR2_X1    g24733(.A1(new_n27167_), .A2(new_n12937_), .ZN(new_n27170_));
  NAND2_X1   g24734(.A1(new_n26933_), .A2(pi0626), .ZN(new_n27171_));
  NAND2_X1   g24735(.A1(new_n27066_), .A2(new_n12747_), .ZN(new_n27172_));
  AOI21_X1   g24736(.A1(new_n27172_), .A2(new_n27171_), .B(new_n12816_), .ZN(new_n27173_));
  INV_X1     g24737(.I(new_n27143_), .ZN(new_n27174_));
  NOR2_X1    g24738(.A1(new_n26935_), .A2(new_n12911_), .ZN(new_n27175_));
  AOI21_X1   g24739(.A1(new_n27174_), .A2(new_n12911_), .B(new_n27175_), .ZN(new_n27176_));
  NOR2_X1    g24740(.A1(new_n26935_), .A2(pi0626), .ZN(new_n27177_));
  AOI21_X1   g24741(.A1(new_n27066_), .A2(pi0626), .B(new_n27177_), .ZN(new_n27178_));
  OAI22_X1   g24742(.A1(new_n27178_), .A2(new_n12813_), .B1(new_n12906_), .B2(new_n27176_), .ZN(new_n27179_));
  OAI21_X1   g24743(.A1(new_n27179_), .A2(new_n27173_), .B(pi0788), .ZN(new_n27180_));
  INV_X1     g24744(.I(new_n27043_), .ZN(new_n27181_));
  NAND2_X1   g24745(.A1(new_n26942_), .A2(new_n27093_), .ZN(new_n27182_));
  NOR2_X1    g24746(.A1(new_n13569_), .A2(pi0642), .ZN(new_n27183_));
  AOI21_X1   g24747(.A1(pi0642), .A2(new_n13587_), .B(new_n27183_), .ZN(new_n27184_));
  NOR2_X1    g24748(.A1(new_n13568_), .A2(new_n27184_), .ZN(new_n27185_));
  INV_X1     g24749(.I(new_n27185_), .ZN(new_n27186_));
  NAND2_X1   g24750(.A1(new_n27186_), .A2(new_n27075_), .ZN(new_n27187_));
  AOI21_X1   g24751(.A1(new_n27182_), .A2(new_n27187_), .B(new_n2668_), .ZN(new_n27188_));
  INV_X1     g24752(.I(new_n27183_), .ZN(new_n27189_));
  NOR2_X1    g24753(.A1(new_n26738_), .A2(new_n27093_), .ZN(new_n27190_));
  AOI22_X1   g24754(.A1(new_n27190_), .A2(new_n27189_), .B1(new_n26940_), .B2(new_n27093_), .ZN(new_n27191_));
  INV_X1     g24755(.I(new_n27191_), .ZN(new_n27192_));
  OAI21_X1   g24756(.A1(new_n27192_), .A2(new_n27188_), .B(new_n26939_), .ZN(new_n27193_));
  NAND2_X1   g24757(.A1(new_n27193_), .A2(new_n26937_), .ZN(new_n27194_));
  NOR2_X1    g24758(.A1(new_n26626_), .A2(new_n13586_), .ZN(new_n27195_));
  NOR2_X1    g24759(.A1(new_n26753_), .A2(new_n27075_), .ZN(new_n27196_));
  OR3_X2     g24760(.A1(new_n27196_), .A2(new_n27195_), .A3(new_n26947_), .Z(new_n27197_));
  NAND3_X1   g24761(.A1(new_n13806_), .A2(pi0680), .A3(new_n27101_), .ZN(new_n27198_));
  NAND3_X1   g24762(.A1(new_n27197_), .A2(new_n26946_), .A3(new_n27198_), .ZN(new_n27199_));
  NAND2_X1   g24763(.A1(new_n13804_), .A2(new_n27093_), .ZN(new_n27200_));
  NAND4_X1   g24764(.A1(new_n27200_), .A2(pi0223), .A3(new_n26745_), .A4(new_n26951_), .ZN(new_n27201_));
  NAND3_X1   g24765(.A1(new_n13804_), .A2(pi0680), .A3(new_n27101_), .ZN(new_n27202_));
  NAND3_X1   g24766(.A1(new_n26950_), .A2(new_n27201_), .A3(new_n27202_), .ZN(new_n27203_));
  NAND3_X1   g24767(.A1(new_n27199_), .A2(new_n2627_), .A3(new_n27203_), .ZN(new_n27204_));
  INV_X1     g24768(.I(new_n26960_), .ZN(new_n27205_));
  OAI21_X1   g24769(.A1(new_n27205_), .A2(new_n5402_), .B(new_n5399_), .ZN(new_n27206_));
  OAI21_X1   g24770(.A1(new_n27205_), .A2(pi0680), .B(pi0681), .ZN(new_n27207_));
  NOR2_X1    g24771(.A1(new_n27186_), .A2(new_n13678_), .ZN(new_n27208_));
  OAI21_X1   g24772(.A1(new_n27208_), .A2(new_n13095_), .B(pi0680), .ZN(new_n27209_));
  OAI22_X1   g24773(.A1(new_n13706_), .A2(pi0614), .B1(new_n5406_), .B2(new_n13665_), .ZN(new_n27210_));
  AOI21_X1   g24774(.A1(new_n27210_), .A2(new_n13111_), .B(new_n27209_), .ZN(new_n27211_));
  OAI22_X1   g24775(.A1(new_n26956_), .A2(new_n27206_), .B1(new_n27207_), .B2(new_n27211_), .ZN(new_n27212_));
  NAND2_X1   g24776(.A1(new_n27212_), .A2(new_n5446_), .ZN(new_n27213_));
  NOR3_X1    g24777(.A1(new_n13215_), .A2(new_n13095_), .A3(new_n13654_), .ZN(new_n27214_));
  NOR2_X1    g24778(.A1(new_n26783_), .A2(new_n5406_), .ZN(new_n27215_));
  NOR4_X1    g24779(.A1(new_n27214_), .A2(new_n13714_), .A3(new_n27215_), .A4(new_n12821_), .ZN(new_n27216_));
  NOR2_X1    g24780(.A1(new_n26964_), .A2(pi0680), .ZN(new_n27217_));
  NOR3_X1    g24781(.A1(new_n27217_), .A2(new_n27216_), .A3(new_n5399_), .ZN(new_n27218_));
  OR2_X2     g24782(.A1(new_n26964_), .A2(new_n5402_), .Z(new_n27219_));
  AOI21_X1   g24783(.A1(new_n27021_), .A2(new_n27219_), .B(new_n27218_), .ZN(new_n27220_));
  OR2_X2     g24784(.A1(new_n27220_), .A2(new_n5446_), .Z(new_n27221_));
  AOI21_X1   g24785(.A1(new_n27213_), .A2(new_n27221_), .B(new_n2668_), .ZN(new_n27222_));
  INV_X1     g24786(.I(new_n26977_), .ZN(new_n27223_));
  INV_X1     g24787(.I(new_n13769_), .ZN(new_n27224_));
  AOI21_X1   g24788(.A1(new_n26824_), .A2(pi0642), .B(new_n12821_), .ZN(new_n27225_));
  NAND2_X1   g24789(.A1(new_n27224_), .A2(new_n27225_), .ZN(new_n27226_));
  NOR2_X1    g24790(.A1(new_n13095_), .A2(pi0642), .ZN(new_n27227_));
  INV_X1     g24791(.I(new_n27227_), .ZN(new_n27228_));
  NOR2_X1    g24792(.A1(new_n26820_), .A2(new_n27228_), .ZN(new_n27229_));
  OAI22_X1   g24793(.A1(new_n27229_), .A2(new_n27226_), .B1(new_n26978_), .B2(new_n27075_), .ZN(new_n27230_));
  NAND2_X1   g24794(.A1(new_n27230_), .A2(new_n27223_), .ZN(new_n27231_));
  NAND2_X1   g24795(.A1(new_n27231_), .A2(new_n5445_), .ZN(new_n27232_));
  NOR2_X1    g24796(.A1(new_n26981_), .A2(pi0680), .ZN(new_n27233_));
  NOR2_X1    g24797(.A1(new_n13665_), .A2(new_n5406_), .ZN(new_n27234_));
  OAI21_X1   g24798(.A1(new_n27234_), .A2(new_n13569_), .B(new_n13105_), .ZN(new_n27235_));
  NAND2_X1   g24799(.A1(new_n27235_), .A2(pi0680), .ZN(new_n27236_));
  INV_X1     g24800(.I(new_n13588_), .ZN(new_n27237_));
  AOI21_X1   g24801(.A1(new_n27237_), .A2(pi0642), .B(new_n13096_), .ZN(new_n27238_));
  NOR2_X1    g24802(.A1(new_n13629_), .A2(pi0642), .ZN(new_n27239_));
  INV_X1     g24803(.I(new_n27239_), .ZN(new_n27240_));
  AOI21_X1   g24804(.A1(new_n27240_), .A2(new_n27238_), .B(new_n27236_), .ZN(new_n27241_));
  OAI21_X1   g24805(.A1(new_n27241_), .A2(new_n27233_), .B(pi0681), .ZN(new_n27242_));
  NAND2_X1   g24806(.A1(new_n27242_), .A2(new_n26985_), .ZN(new_n27243_));
  NAND2_X1   g24807(.A1(new_n27243_), .A2(new_n5446_), .ZN(new_n27244_));
  NAND2_X1   g24808(.A1(new_n27232_), .A2(new_n27244_), .ZN(new_n27245_));
  OAI21_X1   g24809(.A1(new_n27191_), .A2(new_n13088_), .B(new_n2641_), .ZN(new_n27246_));
  NAND2_X1   g24810(.A1(new_n27246_), .A2(new_n2668_), .ZN(new_n27247_));
  AOI21_X1   g24811(.A1(new_n27245_), .A2(new_n2642_), .B(new_n27247_), .ZN(new_n27248_));
  OR3_X2     g24812(.A1(new_n27248_), .A2(pi0299), .A3(new_n27222_), .Z(new_n27249_));
  INV_X1     g24813(.I(new_n26990_), .ZN(new_n27250_));
  NOR3_X1    g24814(.A1(new_n27191_), .A2(pi0223), .A3(new_n13088_), .ZN(new_n27251_));
  NOR3_X1    g24815(.A1(new_n27251_), .A2(new_n27250_), .A3(new_n27188_), .ZN(new_n27252_));
  NAND3_X1   g24816(.A1(new_n27242_), .A2(new_n5422_), .A3(new_n26985_), .ZN(new_n27253_));
  NAND3_X1   g24817(.A1(new_n27230_), .A2(new_n6764_), .A3(new_n27223_), .ZN(new_n27254_));
  AOI21_X1   g24818(.A1(new_n27254_), .A2(new_n27253_), .B(pi0223), .ZN(new_n27255_));
  OAI21_X1   g24819(.A1(new_n26802_), .A2(new_n5406_), .B(pi0680), .ZN(new_n27256_));
  AOI21_X1   g24820(.A1(new_n26801_), .A2(new_n27227_), .B(new_n27256_), .ZN(new_n27257_));
  NAND2_X1   g24821(.A1(new_n26796_), .A2(new_n5408_), .ZN(new_n27258_));
  AOI22_X1   g24822(.A1(new_n27001_), .A2(new_n27093_), .B1(new_n27257_), .B2(new_n27258_), .ZN(new_n27259_));
  NOR2_X1    g24823(.A1(new_n27259_), .A2(new_n27000_), .ZN(new_n27260_));
  INV_X1     g24824(.I(new_n27008_), .ZN(new_n27261_));
  INV_X1     g24825(.I(new_n27209_), .ZN(new_n27262_));
  AOI21_X1   g24826(.A1(new_n26274_), .A2(new_n13570_), .B(pi0642), .ZN(new_n27263_));
  OAI21_X1   g24827(.A1(new_n27263_), .A2(new_n27234_), .B(new_n13095_), .ZN(new_n27264_));
  AOI22_X1   g24828(.A1(new_n27261_), .A2(new_n27093_), .B1(new_n27262_), .B2(new_n27264_), .ZN(new_n27265_));
  OAI21_X1   g24829(.A1(new_n27265_), .A2(new_n27013_), .B(pi0223), .ZN(new_n27266_));
  OAI21_X1   g24830(.A1(new_n27266_), .A2(new_n27260_), .B(new_n3304_), .ZN(new_n27267_));
  OAI21_X1   g24831(.A1(new_n27267_), .A2(new_n27255_), .B(new_n2436_), .ZN(new_n27268_));
  AOI21_X1   g24832(.A1(new_n27023_), .A2(new_n12821_), .B(new_n5399_), .ZN(new_n27269_));
  AOI21_X1   g24833(.A1(new_n26766_), .A2(pi0642), .B(new_n12821_), .ZN(new_n27270_));
  OAI21_X1   g24834(.A1(new_n13779_), .A2(new_n27228_), .B(new_n27270_), .ZN(new_n27271_));
  NOR2_X1    g24835(.A1(new_n13579_), .A2(new_n13780_), .ZN(new_n27272_));
  NOR2_X1    g24836(.A1(new_n27272_), .A2(new_n13264_), .ZN(new_n27273_));
  OAI21_X1   g24837(.A1(new_n27271_), .A2(new_n27273_), .B(new_n27269_), .ZN(new_n27274_));
  NAND3_X1   g24838(.A1(new_n27274_), .A2(new_n6764_), .A3(new_n27022_), .ZN(new_n27275_));
  NAND2_X1   g24839(.A1(new_n13780_), .A2(new_n5406_), .ZN(new_n27276_));
  AOI21_X1   g24840(.A1(new_n27276_), .A2(new_n27238_), .B(new_n27236_), .ZN(new_n27277_));
  OAI21_X1   g24841(.A1(new_n27277_), .A2(new_n27233_), .B(pi0681), .ZN(new_n27278_));
  NAND2_X1   g24842(.A1(new_n27278_), .A2(new_n27026_), .ZN(new_n27279_));
  NAND3_X1   g24843(.A1(new_n27275_), .A2(new_n2668_), .A3(new_n27279_), .ZN(new_n27280_));
  NAND2_X1   g24844(.A1(new_n27220_), .A2(new_n6764_), .ZN(new_n27281_));
  OAI21_X1   g24845(.A1(new_n27212_), .A2(new_n6764_), .B(new_n27281_), .ZN(new_n27282_));
  AOI21_X1   g24846(.A1(new_n27282_), .A2(pi0223), .B(new_n2436_), .ZN(new_n27283_));
  AOI21_X1   g24847(.A1(new_n27283_), .A2(new_n27280_), .B(new_n2628_), .ZN(new_n27284_));
  OAI21_X1   g24848(.A1(new_n27252_), .A2(new_n27268_), .B(new_n27284_), .ZN(new_n27285_));
  NAND3_X1   g24849(.A1(new_n27249_), .A2(new_n27285_), .A3(pi0039), .ZN(new_n27286_));
  NAND3_X1   g24850(.A1(new_n27286_), .A2(new_n3265_), .A3(new_n27204_), .ZN(new_n27287_));
  NAND3_X1   g24851(.A1(new_n27287_), .A2(new_n2609_), .A3(new_n27194_), .ZN(new_n27288_));
  OAI21_X1   g24852(.A1(new_n2668_), .A2(new_n2609_), .B(new_n27288_), .ZN(new_n27289_));
  NAND2_X1   g24853(.A1(new_n27289_), .A2(new_n12758_), .ZN(new_n27290_));
  INV_X1     g24854(.I(new_n27132_), .ZN(new_n27291_));
  NOR2_X1    g24855(.A1(new_n27036_), .A2(new_n13521_), .ZN(new_n27292_));
  AOI21_X1   g24856(.A1(new_n27289_), .A2(new_n13521_), .B(new_n27292_), .ZN(new_n27293_));
  OAI21_X1   g24857(.A1(new_n27293_), .A2(pi1153), .B(new_n27135_), .ZN(new_n27294_));
  NOR2_X1    g24858(.A1(new_n27036_), .A2(pi0625), .ZN(new_n27295_));
  AOI21_X1   g24859(.A1(new_n27289_), .A2(pi0625), .B(new_n27295_), .ZN(new_n27296_));
  OAI21_X1   g24860(.A1(new_n27296_), .A2(new_n12841_), .B(pi0608), .ZN(new_n27297_));
  OAI22_X1   g24861(.A1(pi0608), .A2(new_n27294_), .B1(new_n27297_), .B2(new_n27291_), .ZN(new_n27298_));
  OAI21_X1   g24862(.A1(new_n27298_), .A2(new_n12758_), .B(new_n27290_), .ZN(new_n27299_));
  NAND2_X1   g24863(.A1(new_n27299_), .A2(new_n12766_), .ZN(new_n27300_));
  NAND2_X1   g24864(.A1(new_n27138_), .A2(pi0609), .ZN(new_n27301_));
  AOI21_X1   g24865(.A1(new_n27300_), .A2(new_n27301_), .B(pi1155), .ZN(new_n27302_));
  NOR3_X1    g24866(.A1(new_n27302_), .A2(pi0660), .A3(new_n27181_), .ZN(new_n27303_));
  NAND2_X1   g24867(.A1(new_n27299_), .A2(pi0609), .ZN(new_n27304_));
  OAI21_X1   g24868(.A1(pi0609), .A2(new_n27137_), .B(new_n27304_), .ZN(new_n27305_));
  NAND2_X1   g24869(.A1(new_n27040_), .A2(pi0660), .ZN(new_n27306_));
  AOI21_X1   g24870(.A1(new_n27305_), .A2(pi1155), .B(new_n27306_), .ZN(new_n27307_));
  NOR3_X1    g24871(.A1(new_n27307_), .A2(new_n27303_), .A3(new_n12764_), .ZN(new_n27308_));
  NAND2_X1   g24872(.A1(new_n27299_), .A2(new_n12764_), .ZN(new_n27309_));
  INV_X1     g24873(.I(new_n27309_), .ZN(new_n27310_));
  NOR2_X1    g24874(.A1(new_n27308_), .A2(new_n27310_), .ZN(new_n27311_));
  NAND2_X1   g24875(.A1(new_n27050_), .A2(pi0627), .ZN(new_n27312_));
  AOI21_X1   g24876(.A1(new_n27140_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n27313_));
  NAND2_X1   g24877(.A1(new_n27311_), .A2(pi0618), .ZN(new_n27314_));
  AOI21_X1   g24878(.A1(new_n27314_), .A2(new_n27313_), .B(new_n27312_), .ZN(new_n27315_));
  NOR2_X1    g24879(.A1(new_n27053_), .A2(pi0627), .ZN(new_n27316_));
  INV_X1     g24880(.I(new_n27311_), .ZN(new_n27317_));
  AOI21_X1   g24881(.A1(new_n27140_), .A2(pi0618), .B(pi1154), .ZN(new_n27318_));
  OAI21_X1   g24882(.A1(new_n27317_), .A2(pi0618), .B(new_n27318_), .ZN(new_n27319_));
  NAND2_X1   g24883(.A1(new_n27319_), .A2(new_n27316_), .ZN(new_n27320_));
  NAND2_X1   g24884(.A1(new_n27320_), .A2(pi0781), .ZN(new_n27321_));
  OAI22_X1   g24885(.A1(new_n27321_), .A2(new_n27315_), .B1(pi0781), .B2(new_n27311_), .ZN(new_n27322_));
  AOI21_X1   g24886(.A1(new_n27322_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n27323_));
  INV_X1     g24887(.I(new_n27064_), .ZN(new_n27324_));
  NAND2_X1   g24888(.A1(new_n27322_), .A2(new_n12793_), .ZN(new_n27325_));
  NAND2_X1   g24889(.A1(new_n27143_), .A2(pi0619), .ZN(new_n27326_));
  AOI21_X1   g24890(.A1(new_n27325_), .A2(new_n27326_), .B(pi1159), .ZN(new_n27327_));
  NOR3_X1    g24891(.A1(new_n27327_), .A2(pi0648), .A3(new_n27324_), .ZN(new_n27328_));
  NOR2_X1    g24892(.A1(new_n27174_), .A2(pi0619), .ZN(new_n27329_));
  AOI21_X1   g24893(.A1(new_n27322_), .A2(pi0619), .B(new_n27329_), .ZN(new_n27330_));
  OAI21_X1   g24894(.A1(new_n27330_), .A2(new_n12791_), .B(pi0648), .ZN(new_n27331_));
  OAI21_X1   g24895(.A1(new_n27331_), .A2(new_n27061_), .B(pi0789), .ZN(new_n27332_));
  OAI21_X1   g24896(.A1(new_n27332_), .A2(new_n27328_), .B(new_n27323_), .ZN(new_n27333_));
  AOI21_X1   g24897(.A1(new_n27333_), .A2(new_n27180_), .B(new_n27170_), .ZN(new_n27334_));
  OAI21_X1   g24898(.A1(new_n27334_), .A2(new_n27169_), .B(new_n27158_), .ZN(new_n27335_));
  NAND2_X1   g24899(.A1(new_n26935_), .A2(pi0644), .ZN(new_n27336_));
  NOR2_X1    g24900(.A1(new_n27070_), .A2(new_n12984_), .ZN(new_n27337_));
  AOI21_X1   g24901(.A1(new_n12984_), .A2(new_n26935_), .B(new_n27337_), .ZN(new_n27338_));
  OAI21_X1   g24902(.A1(new_n27338_), .A2(pi0644), .B(new_n27336_), .ZN(new_n27339_));
  AOI21_X1   g24903(.A1(new_n27339_), .A2(pi0715), .B(pi1160), .ZN(new_n27340_));
  NOR2_X1    g24904(.A1(new_n27150_), .A2(new_n12972_), .ZN(new_n27341_));
  AOI22_X1   g24905(.A1(new_n27341_), .A2(new_n27154_), .B1(new_n12972_), .B2(new_n27152_), .ZN(new_n27342_));
  OAI21_X1   g24906(.A1(new_n27342_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n27343_));
  NOR2_X1    g24907(.A1(new_n27335_), .A2(pi0644), .ZN(new_n27344_));
  OAI21_X1   g24908(.A1(new_n27344_), .A2(new_n27343_), .B(new_n27340_), .ZN(new_n27345_));
  NAND2_X1   g24909(.A1(new_n26935_), .A2(new_n12975_), .ZN(new_n27346_));
  OAI21_X1   g24910(.A1(new_n27338_), .A2(new_n12975_), .B(new_n27346_), .ZN(new_n27347_));
  AOI21_X1   g24911(.A1(new_n27347_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n27348_));
  NOR2_X1    g24912(.A1(new_n27342_), .A2(pi0644), .ZN(new_n27349_));
  NOR2_X1    g24913(.A1(new_n27349_), .A2(new_n12740_), .ZN(new_n27350_));
  OAI21_X1   g24914(.A1(new_n27335_), .A2(new_n12975_), .B(new_n27350_), .ZN(new_n27351_));
  AOI21_X1   g24915(.A1(new_n27351_), .A2(new_n27348_), .B(new_n13000_), .ZN(new_n27352_));
  AOI22_X1   g24916(.A1(new_n27352_), .A2(new_n27345_), .B1(new_n13000_), .B2(new_n27335_), .ZN(new_n27353_));
  OAI21_X1   g24917(.A1(new_n27353_), .A2(po1038), .B(new_n26928_), .ZN(po0380));
  NAND2_X1   g24918(.A1(po1038), .A2(pi0224), .ZN(new_n27355_));
  NOR2_X1    g24919(.A1(new_n26491_), .A2(new_n2631_), .ZN(new_n27356_));
  INV_X1     g24920(.I(new_n27356_), .ZN(new_n27357_));
  AOI21_X1   g24921(.A1(new_n13397_), .A2(pi0224), .B(new_n3265_), .ZN(new_n27358_));
  INV_X1     g24922(.I(new_n27358_), .ZN(new_n27359_));
  AOI21_X1   g24923(.A1(pi0614), .A2(new_n13341_), .B(new_n27359_), .ZN(new_n27360_));
  NOR2_X1    g24924(.A1(new_n14666_), .A2(new_n5405_), .ZN(new_n27361_));
  AOI21_X1   g24925(.A1(new_n27361_), .A2(new_n2631_), .B(pi0299), .ZN(new_n27362_));
  OAI21_X1   g24926(.A1(new_n14666_), .A2(pi0614), .B(pi0224), .ZN(new_n27363_));
  OAI21_X1   g24927(.A1(new_n14547_), .A2(new_n27363_), .B(new_n27362_), .ZN(new_n27364_));
  NAND2_X1   g24928(.A1(new_n14553_), .A2(pi0614), .ZN(new_n27365_));
  INV_X1     g24929(.I(new_n27365_), .ZN(new_n27366_));
  NAND2_X1   g24930(.A1(new_n14558_), .A2(pi0224), .ZN(new_n27367_));
  AOI22_X1   g24931(.A1(new_n27366_), .A2(new_n27367_), .B1(pi0224), .B2(new_n13055_), .ZN(new_n27368_));
  NAND2_X1   g24932(.A1(new_n27368_), .A2(pi0299), .ZN(new_n27369_));
  NAND3_X1   g24933(.A1(new_n27364_), .A2(new_n27369_), .A3(new_n2627_), .ZN(new_n27370_));
  NOR2_X1    g24934(.A1(new_n12755_), .A2(new_n5405_), .ZN(new_n27371_));
  INV_X1     g24935(.I(new_n27371_), .ZN(new_n27372_));
  AOI21_X1   g24936(.A1(new_n13098_), .A2(new_n27372_), .B(new_n5410_), .ZN(new_n27373_));
  NOR3_X1    g24937(.A1(new_n13159_), .A2(pi0680), .A3(new_n27373_), .ZN(new_n27374_));
  NOR3_X1    g24938(.A1(new_n26116_), .A2(new_n12821_), .A3(new_n27371_), .ZN(new_n27375_));
  NOR2_X1    g24939(.A1(new_n27374_), .A2(new_n27375_), .ZN(new_n27376_));
  NOR2_X1    g24940(.A1(new_n13159_), .A2(new_n27373_), .ZN(new_n27377_));
  NAND2_X1   g24941(.A1(new_n27377_), .A2(new_n13119_), .ZN(new_n27378_));
  OAI21_X1   g24942(.A1(new_n27376_), .A2(new_n13119_), .B(new_n27378_), .ZN(new_n27379_));
  NOR2_X1    g24943(.A1(new_n27379_), .A2(new_n5445_), .ZN(new_n27380_));
  AOI21_X1   g24944(.A1(pi0614), .A2(new_n13277_), .B(new_n26333_), .ZN(new_n27381_));
  INV_X1     g24945(.I(new_n13275_), .ZN(new_n27382_));
  NAND2_X1   g24946(.A1(new_n27382_), .A2(pi0614), .ZN(new_n27383_));
  AOI21_X1   g24947(.A1(new_n13274_), .A2(new_n27383_), .B(new_n12821_), .ZN(new_n27384_));
  NOR2_X1    g24948(.A1(new_n27381_), .A2(pi0680), .ZN(new_n27385_));
  OAI21_X1   g24949(.A1(new_n27385_), .A2(new_n27384_), .B(new_n13118_), .ZN(new_n27386_));
  OAI21_X1   g24950(.A1(new_n13118_), .A2(new_n27381_), .B(new_n27386_), .ZN(new_n27387_));
  AOI21_X1   g24951(.A1(new_n27387_), .A2(new_n5445_), .B(new_n27380_), .ZN(new_n27388_));
  NOR2_X1    g24952(.A1(new_n13214_), .A2(new_n5405_), .ZN(new_n27389_));
  INV_X1     g24953(.I(new_n27389_), .ZN(new_n27390_));
  NOR2_X1    g24954(.A1(new_n26555_), .A2(new_n27390_), .ZN(new_n27391_));
  INV_X1     g24955(.I(new_n27391_), .ZN(new_n27392_));
  NOR2_X1    g24956(.A1(new_n27392_), .A2(pi0224), .ZN(new_n27393_));
  INV_X1     g24957(.I(new_n27393_), .ZN(new_n27394_));
  NOR2_X1    g24958(.A1(new_n27394_), .A2(new_n13235_), .ZN(new_n27395_));
  NOR2_X1    g24959(.A1(new_n27395_), .A2(new_n2668_), .ZN(new_n27396_));
  OAI21_X1   g24960(.A1(new_n27388_), .A2(new_n2631_), .B(new_n27396_), .ZN(new_n27397_));
  NAND3_X1   g24961(.A1(new_n13185_), .A2(pi0614), .A3(new_n12754_), .ZN(new_n27398_));
  NAND2_X1   g24962(.A1(new_n26437_), .A2(new_n13111_), .ZN(new_n27399_));
  INV_X1     g24963(.I(new_n27373_), .ZN(new_n27400_));
  NAND3_X1   g24964(.A1(new_n27399_), .A2(new_n12821_), .A3(new_n27400_), .ZN(new_n27401_));
  NOR2_X1    g24965(.A1(new_n27371_), .A2(new_n12821_), .ZN(new_n27402_));
  NAND2_X1   g24966(.A1(new_n13304_), .A2(new_n27402_), .ZN(new_n27403_));
  NAND2_X1   g24967(.A1(new_n27401_), .A2(new_n27403_), .ZN(new_n27404_));
  NAND2_X1   g24968(.A1(new_n27399_), .A2(new_n27400_), .ZN(new_n27405_));
  NOR2_X1    g24969(.A1(new_n27405_), .A2(new_n13118_), .ZN(new_n27406_));
  AOI21_X1   g24970(.A1(new_n27404_), .A2(new_n13118_), .B(new_n27406_), .ZN(new_n27407_));
  AND2_X2    g24971(.A1(new_n27407_), .A2(new_n5446_), .Z(new_n27408_));
  AOI21_X1   g24972(.A1(new_n13721_), .A2(pi0614), .B(new_n12821_), .ZN(new_n27409_));
  INV_X1     g24973(.I(new_n27409_), .ZN(new_n27410_));
  NAND2_X1   g24974(.A1(new_n5405_), .A2(pi0616), .ZN(new_n27411_));
  OAI22_X1   g24975(.A1(new_n13317_), .A2(new_n5405_), .B1(new_n13603_), .B2(new_n27411_), .ZN(new_n27412_));
  NAND2_X1   g24976(.A1(new_n26435_), .A2(new_n13095_), .ZN(new_n27413_));
  AOI21_X1   g24977(.A1(new_n5437_), .A2(new_n26436_), .B(new_n27413_), .ZN(new_n27414_));
  OR2_X2     g24978(.A1(new_n27412_), .A2(new_n27414_), .Z(new_n27415_));
  NOR2_X1    g24979(.A1(new_n27415_), .A2(pi0680), .ZN(new_n27416_));
  OAI22_X1   g24980(.A1(new_n27416_), .A2(new_n27402_), .B1(new_n13082_), .B2(new_n27410_), .ZN(new_n27417_));
  NAND2_X1   g24981(.A1(new_n27417_), .A2(new_n13118_), .ZN(new_n27418_));
  NAND2_X1   g24982(.A1(new_n27415_), .A2(new_n13119_), .ZN(new_n27419_));
  AOI21_X1   g24983(.A1(new_n27418_), .A2(new_n27419_), .B(new_n5446_), .ZN(new_n27420_));
  OAI21_X1   g24984(.A1(new_n27420_), .A2(new_n27408_), .B(pi0224), .ZN(new_n27421_));
  NOR2_X1    g24985(.A1(new_n26504_), .A2(new_n5405_), .ZN(new_n27422_));
  INV_X1     g24986(.I(new_n27422_), .ZN(new_n27423_));
  NOR2_X1    g24987(.A1(new_n27423_), .A2(new_n5445_), .ZN(new_n27424_));
  NOR2_X1    g24988(.A1(new_n13316_), .A2(new_n27372_), .ZN(new_n27425_));
  NOR2_X1    g24989(.A1(new_n27425_), .A2(pi0680), .ZN(new_n27426_));
  INV_X1     g24990(.I(new_n27426_), .ZN(new_n27427_));
  AOI21_X1   g24991(.A1(new_n27427_), .A2(new_n27410_), .B(new_n13119_), .ZN(new_n27428_));
  INV_X1     g24992(.I(new_n27428_), .ZN(new_n27429_));
  OAI21_X1   g24993(.A1(new_n13118_), .A2(new_n27425_), .B(new_n27429_), .ZN(new_n27430_));
  NOR2_X1    g24994(.A1(new_n27430_), .A2(new_n5446_), .ZN(new_n27431_));
  OAI21_X1   g24995(.A1(new_n27431_), .A2(new_n27424_), .B(new_n5081_), .ZN(new_n27432_));
  NAND4_X1   g24996(.A1(new_n27421_), .A2(new_n2668_), .A3(new_n27398_), .A4(new_n27432_), .ZN(new_n27433_));
  NAND2_X1   g24997(.A1(new_n27433_), .A2(new_n27397_), .ZN(new_n27434_));
  NAND2_X1   g24998(.A1(new_n27434_), .A2(new_n2628_), .ZN(new_n27435_));
  OAI21_X1   g24999(.A1(new_n13098_), .A2(new_n2631_), .B(new_n3303_), .ZN(new_n27436_));
  OAI21_X1   g25000(.A1(new_n27389_), .A2(new_n27436_), .B(new_n2436_), .ZN(new_n27437_));
  NAND2_X1   g25001(.A1(new_n27422_), .A2(new_n5422_), .ZN(new_n27438_));
  OR2_X2     g25002(.A1(new_n27430_), .A2(new_n5422_), .Z(new_n27439_));
  AOI21_X1   g25003(.A1(new_n27439_), .A2(new_n27438_), .B(pi0224), .ZN(new_n27440_));
  NAND2_X1   g25004(.A1(new_n27407_), .A2(new_n5422_), .ZN(new_n27441_));
  NAND2_X1   g25005(.A1(new_n27418_), .A2(new_n27419_), .ZN(new_n27442_));
  NAND2_X1   g25006(.A1(new_n27442_), .A2(new_n6764_), .ZN(new_n27443_));
  AOI21_X1   g25007(.A1(new_n27443_), .A2(new_n27441_), .B(new_n2631_), .ZN(new_n27444_));
  NOR3_X1    g25008(.A1(new_n27444_), .A2(new_n3303_), .A3(new_n27440_), .ZN(new_n27445_));
  NOR2_X1    g25009(.A1(new_n27379_), .A2(new_n6764_), .ZN(new_n27446_));
  AOI21_X1   g25010(.A1(new_n27387_), .A2(new_n6764_), .B(new_n27446_), .ZN(new_n27447_));
  OAI22_X1   g25011(.A1(new_n27447_), .A2(new_n2631_), .B1(new_n13218_), .B2(new_n27394_), .ZN(new_n27448_));
  AOI21_X1   g25012(.A1(new_n27448_), .A2(pi0215), .B(new_n2628_), .ZN(new_n27449_));
  OAI21_X1   g25013(.A1(new_n27445_), .A2(new_n27437_), .B(new_n27449_), .ZN(new_n27450_));
  NAND3_X1   g25014(.A1(new_n27435_), .A2(new_n27450_), .A3(pi0039), .ZN(new_n27451_));
  NAND3_X1   g25015(.A1(new_n27451_), .A2(new_n3265_), .A3(new_n27370_), .ZN(new_n27452_));
  NAND2_X1   g25016(.A1(new_n27452_), .A2(new_n2609_), .ZN(new_n27453_));
  OAI22_X1   g25017(.A1(new_n27453_), .A2(new_n27360_), .B1(new_n2631_), .B2(new_n2609_), .ZN(new_n27454_));
  NOR2_X1    g25018(.A1(new_n27454_), .A2(new_n12760_), .ZN(new_n27455_));
  AOI21_X1   g25019(.A1(new_n12760_), .A2(new_n27357_), .B(new_n27455_), .ZN(new_n27456_));
  INV_X1     g25020(.I(new_n27456_), .ZN(new_n27457_));
  NAND2_X1   g25021(.A1(new_n27456_), .A2(new_n12766_), .ZN(new_n27458_));
  NOR2_X1    g25022(.A1(new_n27357_), .A2(new_n12766_), .ZN(new_n27459_));
  INV_X1     g25023(.I(new_n27459_), .ZN(new_n27460_));
  AOI21_X1   g25024(.A1(new_n27458_), .A2(new_n27460_), .B(pi1155), .ZN(new_n27461_));
  INV_X1     g25025(.I(new_n27461_), .ZN(new_n27462_));
  NAND2_X1   g25026(.A1(new_n27456_), .A2(pi0609), .ZN(new_n27463_));
  NAND2_X1   g25027(.A1(new_n27356_), .A2(new_n12766_), .ZN(new_n27464_));
  AOI21_X1   g25028(.A1(new_n27463_), .A2(new_n27464_), .B(new_n12770_), .ZN(new_n27465_));
  NOR2_X1    g25029(.A1(new_n27465_), .A2(new_n12764_), .ZN(new_n27466_));
  AOI22_X1   g25030(.A1(new_n27466_), .A2(new_n27462_), .B1(new_n12764_), .B2(new_n27457_), .ZN(new_n27467_));
  NOR2_X1    g25031(.A1(new_n27467_), .A2(pi0781), .ZN(new_n27468_));
  NOR2_X1    g25032(.A1(new_n27357_), .A2(new_n12781_), .ZN(new_n27469_));
  AOI21_X1   g25033(.A1(new_n27467_), .A2(new_n12781_), .B(new_n27469_), .ZN(new_n27470_));
  NOR2_X1    g25034(.A1(new_n27470_), .A2(pi1154), .ZN(new_n27471_));
  NAND2_X1   g25035(.A1(new_n27467_), .A2(pi0618), .ZN(new_n27472_));
  NAND2_X1   g25036(.A1(new_n27356_), .A2(new_n12781_), .ZN(new_n27473_));
  AOI21_X1   g25037(.A1(new_n27472_), .A2(new_n27473_), .B(new_n12785_), .ZN(new_n27474_));
  NOR3_X1    g25038(.A1(new_n27471_), .A2(new_n27474_), .A3(new_n12779_), .ZN(new_n27475_));
  OAI21_X1   g25039(.A1(new_n27475_), .A2(new_n27468_), .B(new_n12796_), .ZN(new_n27476_));
  NOR3_X1    g25040(.A1(new_n27475_), .A2(pi0619), .A3(new_n27468_), .ZN(new_n27477_));
  NOR2_X1    g25041(.A1(new_n27357_), .A2(new_n12793_), .ZN(new_n27478_));
  OAI21_X1   g25042(.A1(new_n27477_), .A2(new_n27478_), .B(new_n12791_), .ZN(new_n27479_));
  NOR3_X1    g25043(.A1(new_n27475_), .A2(new_n12793_), .A3(new_n27468_), .ZN(new_n27480_));
  NOR2_X1    g25044(.A1(new_n27357_), .A2(pi0619), .ZN(new_n27481_));
  OAI21_X1   g25045(.A1(new_n27480_), .A2(new_n27481_), .B(pi1159), .ZN(new_n27482_));
  NAND3_X1   g25046(.A1(new_n27479_), .A2(new_n27482_), .A3(pi0789), .ZN(new_n27483_));
  NAND2_X1   g25047(.A1(new_n27483_), .A2(new_n27476_), .ZN(new_n27484_));
  NAND2_X1   g25048(.A1(new_n27356_), .A2(new_n12818_), .ZN(new_n27485_));
  OAI21_X1   g25049(.A1(new_n27484_), .A2(new_n12818_), .B(new_n27485_), .ZN(new_n27486_));
  NAND2_X1   g25050(.A1(new_n27357_), .A2(new_n12943_), .ZN(new_n27487_));
  OAI21_X1   g25051(.A1(new_n27486_), .A2(new_n12943_), .B(new_n27487_), .ZN(new_n27488_));
  NOR2_X1    g25052(.A1(new_n27356_), .A2(new_n12952_), .ZN(new_n27489_));
  NOR2_X1    g25053(.A1(new_n27357_), .A2(new_n12923_), .ZN(new_n27490_));
  NAND2_X1   g25054(.A1(new_n27357_), .A2(new_n12887_), .ZN(new_n27491_));
  NOR2_X1    g25055(.A1(new_n27356_), .A2(new_n12870_), .ZN(new_n27492_));
  NOR2_X1    g25056(.A1(new_n2609_), .A2(new_n2631_), .ZN(new_n27493_));
  AOI21_X1   g25057(.A1(pi0662), .A2(new_n13398_), .B(new_n27359_), .ZN(new_n27494_));
  NOR2_X1    g25058(.A1(new_n13425_), .A2(new_n5400_), .ZN(new_n27495_));
  AOI21_X1   g25059(.A1(new_n27495_), .A2(new_n2631_), .B(new_n2668_), .ZN(new_n27496_));
  NAND2_X1   g25060(.A1(new_n13175_), .A2(new_n5400_), .ZN(new_n27497_));
  OAI21_X1   g25061(.A1(new_n5400_), .A2(new_n13468_), .B(new_n27497_), .ZN(new_n27498_));
  NOR2_X1    g25062(.A1(new_n27498_), .A2(new_n5446_), .ZN(new_n27499_));
  NOR2_X1    g25063(.A1(new_n26665_), .A2(new_n5400_), .ZN(new_n27500_));
  AOI21_X1   g25064(.A1(new_n13179_), .A2(new_n5400_), .B(new_n27500_), .ZN(new_n27501_));
  AND2_X2    g25065(.A1(new_n27501_), .A2(new_n5446_), .Z(new_n27502_));
  OAI21_X1   g25066(.A1(new_n27502_), .A2(new_n27499_), .B(pi0224), .ZN(new_n27503_));
  AOI21_X1   g25067(.A1(new_n27503_), .A2(new_n27496_), .B(pi0299), .ZN(new_n27504_));
  NOR2_X1    g25068(.A1(new_n27090_), .A2(new_n5400_), .ZN(new_n27505_));
  AOI21_X1   g25069(.A1(new_n5400_), .A2(new_n13126_), .B(new_n27505_), .ZN(new_n27506_));
  AOI21_X1   g25070(.A1(new_n26655_), .A2(new_n5401_), .B(new_n13093_), .ZN(new_n27507_));
  NOR2_X1    g25071(.A1(new_n27507_), .A2(new_n5446_), .ZN(new_n27508_));
  AOI21_X1   g25072(.A1(new_n27506_), .A2(new_n5446_), .B(new_n27508_), .ZN(new_n27509_));
  NAND3_X1   g25073(.A1(new_n13185_), .A2(pi0662), .A3(new_n12824_), .ZN(new_n27510_));
  NAND2_X1   g25074(.A1(new_n27510_), .A2(new_n2668_), .ZN(new_n27511_));
  NOR2_X1    g25075(.A1(new_n5400_), .A2(new_n12821_), .ZN(new_n27512_));
  NAND2_X1   g25076(.A1(new_n26642_), .A2(new_n27512_), .ZN(new_n27513_));
  AOI21_X1   g25077(.A1(new_n27513_), .A2(new_n5446_), .B(new_n5082_), .ZN(new_n27514_));
  NAND2_X1   g25078(.A1(new_n13430_), .A2(pi0662), .ZN(new_n27515_));
  NAND2_X1   g25079(.A1(new_n27515_), .A2(new_n5445_), .ZN(new_n27516_));
  AOI21_X1   g25080(.A1(new_n27514_), .A2(new_n27516_), .B(new_n27511_), .ZN(new_n27517_));
  OAI21_X1   g25081(.A1(new_n27509_), .A2(new_n2631_), .B(new_n27517_), .ZN(new_n27518_));
  AOI21_X1   g25082(.A1(new_n27518_), .A2(new_n27504_), .B(new_n2627_), .ZN(new_n27519_));
  NAND3_X1   g25083(.A1(new_n13443_), .A2(new_n2631_), .A3(pi0662), .ZN(new_n27520_));
  NAND2_X1   g25084(.A1(new_n27501_), .A2(new_n5422_), .ZN(new_n27521_));
  OAI21_X1   g25085(.A1(new_n5422_), .A2(new_n27498_), .B(new_n27521_), .ZN(new_n27522_));
  AOI21_X1   g25086(.A1(new_n27522_), .A2(pi0224), .B(new_n2436_), .ZN(new_n27523_));
  AOI21_X1   g25087(.A1(new_n27523_), .A2(new_n27520_), .B(new_n2628_), .ZN(new_n27524_));
  AOI21_X1   g25088(.A1(new_n13421_), .A2(new_n27512_), .B(new_n27436_), .ZN(new_n27525_));
  NOR2_X1    g25089(.A1(new_n27513_), .A2(new_n6764_), .ZN(new_n27526_));
  NOR2_X1    g25090(.A1(new_n27515_), .A2(new_n5422_), .ZN(new_n27527_));
  OAI21_X1   g25091(.A1(new_n27526_), .A2(new_n27527_), .B(new_n2631_), .ZN(new_n27528_));
  NAND2_X1   g25092(.A1(new_n27506_), .A2(new_n5422_), .ZN(new_n27529_));
  OAI21_X1   g25093(.A1(new_n5422_), .A2(new_n27507_), .B(new_n27529_), .ZN(new_n27530_));
  AOI21_X1   g25094(.A1(new_n27530_), .A2(pi0224), .B(new_n3303_), .ZN(new_n27531_));
  AOI21_X1   g25095(.A1(new_n27531_), .A2(new_n27528_), .B(new_n27525_), .ZN(new_n27532_));
  OAI21_X1   g25096(.A1(new_n27532_), .A2(pi0215), .B(new_n27524_), .ZN(new_n27533_));
  NAND2_X1   g25097(.A1(new_n27533_), .A2(new_n27519_), .ZN(new_n27534_));
  AOI21_X1   g25098(.A1(new_n26627_), .A2(pi0224), .B(pi0299), .ZN(new_n27535_));
  INV_X1     g25099(.I(new_n27512_), .ZN(new_n27536_));
  NOR2_X1    g25100(.A1(new_n13414_), .A2(new_n27536_), .ZN(new_n27537_));
  NOR2_X1    g25101(.A1(new_n14667_), .A2(new_n2631_), .ZN(new_n27538_));
  OAI21_X1   g25102(.A1(new_n27538_), .A2(new_n27537_), .B(new_n27535_), .ZN(new_n27539_));
  NAND2_X1   g25103(.A1(new_n14655_), .A2(new_n2631_), .ZN(new_n27540_));
  OAI21_X1   g25104(.A1(new_n2631_), .A2(new_n24501_), .B(new_n27540_), .ZN(new_n27541_));
  NAND2_X1   g25105(.A1(new_n14655_), .A2(new_n27536_), .ZN(new_n27542_));
  NAND3_X1   g25106(.A1(new_n27541_), .A2(pi0299), .A3(new_n27542_), .ZN(new_n27543_));
  NAND3_X1   g25107(.A1(new_n27543_), .A2(new_n2627_), .A3(new_n27539_), .ZN(new_n27544_));
  AOI21_X1   g25108(.A1(new_n27534_), .A2(new_n27544_), .B(pi0038), .ZN(new_n27545_));
  NOR3_X1    g25109(.A1(new_n27545_), .A2(new_n2610_), .A3(new_n27494_), .ZN(new_n27546_));
  NOR2_X1    g25110(.A1(new_n27546_), .A2(new_n27493_), .ZN(new_n27547_));
  NAND2_X1   g25111(.A1(new_n27547_), .A2(new_n12758_), .ZN(new_n27548_));
  NOR2_X1    g25112(.A1(new_n27547_), .A2(pi0625), .ZN(new_n27549_));
  NOR2_X1    g25113(.A1(new_n27357_), .A2(new_n13521_), .ZN(new_n27550_));
  OAI21_X1   g25114(.A1(new_n27549_), .A2(new_n27550_), .B(new_n12841_), .ZN(new_n27551_));
  NOR2_X1    g25115(.A1(new_n27547_), .A2(new_n13521_), .ZN(new_n27552_));
  NOR2_X1    g25116(.A1(new_n27357_), .A2(pi0625), .ZN(new_n27553_));
  OAI21_X1   g25117(.A1(new_n27552_), .A2(new_n27553_), .B(pi1153), .ZN(new_n27554_));
  NAND3_X1   g25118(.A1(new_n27551_), .A2(new_n27554_), .A3(pi0778), .ZN(new_n27555_));
  NAND2_X1   g25119(.A1(new_n27555_), .A2(new_n27548_), .ZN(new_n27556_));
  AOI21_X1   g25120(.A1(new_n27556_), .A2(new_n12870_), .B(new_n27492_), .ZN(new_n27557_));
  INV_X1     g25121(.I(new_n27557_), .ZN(new_n27558_));
  NAND2_X1   g25122(.A1(new_n27558_), .A2(new_n12888_), .ZN(new_n27559_));
  NAND2_X1   g25123(.A1(new_n27559_), .A2(new_n27491_), .ZN(new_n27560_));
  INV_X1     g25124(.I(new_n27560_), .ZN(new_n27561_));
  AOI21_X1   g25125(.A1(new_n27561_), .A2(new_n12923_), .B(new_n27490_), .ZN(new_n27562_));
  AOI21_X1   g25126(.A1(new_n27562_), .A2(new_n12952_), .B(new_n27489_), .ZN(new_n27563_));
  NOR2_X1    g25127(.A1(new_n27357_), .A2(pi0647), .ZN(new_n27564_));
  AOI21_X1   g25128(.A1(new_n27563_), .A2(pi0647), .B(new_n27564_), .ZN(new_n27565_));
  NOR2_X1    g25129(.A1(new_n27565_), .A2(new_n12965_), .ZN(new_n27566_));
  NOR2_X1    g25130(.A1(new_n27566_), .A2(pi0630), .ZN(new_n27567_));
  NAND2_X1   g25131(.A1(new_n27356_), .A2(pi0647), .ZN(new_n27568_));
  NAND2_X1   g25132(.A1(new_n27563_), .A2(new_n12741_), .ZN(new_n27569_));
  AOI21_X1   g25133(.A1(new_n27569_), .A2(new_n27568_), .B(pi1157), .ZN(new_n27570_));
  NOR2_X1    g25134(.A1(new_n27570_), .A2(new_n12981_), .ZN(new_n27571_));
  OAI22_X1   g25135(.A1(new_n27488_), .A2(new_n17212_), .B1(new_n27567_), .B2(new_n27571_), .ZN(new_n27572_));
  NAND2_X1   g25136(.A1(new_n27572_), .A2(pi0787), .ZN(new_n27573_));
  NAND2_X1   g25137(.A1(new_n27486_), .A2(new_n19160_), .ZN(new_n27574_));
  NAND2_X1   g25138(.A1(new_n27562_), .A2(pi0628), .ZN(new_n27575_));
  AOI21_X1   g25139(.A1(new_n27357_), .A2(new_n12920_), .B(new_n18087_), .ZN(new_n27576_));
  AOI21_X1   g25140(.A1(new_n27357_), .A2(pi0628), .B(new_n18088_), .ZN(new_n27577_));
  NAND2_X1   g25141(.A1(new_n27562_), .A2(new_n12920_), .ZN(new_n27578_));
  AOI22_X1   g25142(.A1(new_n27575_), .A2(new_n27576_), .B1(new_n27578_), .B2(new_n27577_), .ZN(new_n27579_));
  NAND2_X1   g25143(.A1(new_n27574_), .A2(new_n27579_), .ZN(new_n27580_));
  NOR2_X1    g25144(.A1(new_n27356_), .A2(pi0626), .ZN(new_n27581_));
  AOI21_X1   g25145(.A1(new_n27483_), .A2(new_n27476_), .B(new_n12747_), .ZN(new_n27582_));
  OAI21_X1   g25146(.A1(new_n27582_), .A2(new_n27581_), .B(new_n12812_), .ZN(new_n27583_));
  NOR2_X1    g25147(.A1(new_n27356_), .A2(new_n12911_), .ZN(new_n27584_));
  NOR2_X1    g25148(.A1(new_n27561_), .A2(new_n12910_), .ZN(new_n27585_));
  OAI21_X1   g25149(.A1(new_n27585_), .A2(new_n27584_), .B(new_n14386_), .ZN(new_n27586_));
  AOI21_X1   g25150(.A1(new_n27356_), .A2(pi0626), .B(new_n12816_), .ZN(new_n27587_));
  OAI21_X1   g25151(.A1(new_n27484_), .A2(pi0626), .B(new_n27587_), .ZN(new_n27588_));
  NAND3_X1   g25152(.A1(new_n27583_), .A2(new_n27588_), .A3(new_n27586_), .ZN(new_n27589_));
  AOI21_X1   g25153(.A1(new_n27589_), .A2(pi0788), .B(new_n15340_), .ZN(new_n27590_));
  NAND3_X1   g25154(.A1(new_n13344_), .A2(pi0662), .A3(new_n13571_), .ZN(new_n27591_));
  NAND2_X1   g25155(.A1(new_n27360_), .A2(new_n27591_), .ZN(new_n27592_));
  NOR2_X1    g25156(.A1(new_n13665_), .A2(new_n5405_), .ZN(new_n27593_));
  OAI21_X1   g25157(.A1(new_n13707_), .A2(new_n27593_), .B(new_n13111_), .ZN(new_n27594_));
  NAND2_X1   g25158(.A1(new_n26738_), .A2(pi0614), .ZN(new_n27595_));
  OAI21_X1   g25159(.A1(pi0614), .A2(new_n18102_), .B(new_n27595_), .ZN(new_n27596_));
  NAND2_X1   g25160(.A1(new_n27596_), .A2(new_n13679_), .ZN(new_n27597_));
  AOI21_X1   g25161(.A1(new_n27597_), .A2(pi0616), .B(new_n12821_), .ZN(new_n27598_));
  AOI21_X1   g25162(.A1(new_n27594_), .A2(new_n27598_), .B(new_n27374_), .ZN(new_n27599_));
  AOI22_X1   g25163(.A1(new_n27599_), .A2(pi0662), .B1(new_n13118_), .B2(new_n27376_), .ZN(new_n27600_));
  NOR2_X1    g25164(.A1(new_n13116_), .A2(pi0662), .ZN(new_n27601_));
  INV_X1     g25165(.I(new_n27601_), .ZN(new_n27602_));
  OAI21_X1   g25166(.A1(new_n27377_), .A2(new_n27602_), .B(new_n27600_), .ZN(new_n27603_));
  NAND2_X1   g25167(.A1(new_n27603_), .A2(pi0224), .ZN(new_n27604_));
  INV_X1     g25168(.I(new_n13759_), .ZN(new_n27605_));
  OAI21_X1   g25169(.A1(new_n27605_), .A2(pi0614), .B(new_n13588_), .ZN(new_n27606_));
  NAND3_X1   g25170(.A1(new_n27606_), .A2(pi0616), .A3(pi0680), .ZN(new_n27607_));
  NAND2_X1   g25171(.A1(new_n27607_), .A2(pi0662), .ZN(new_n27608_));
  NOR2_X1    g25172(.A1(new_n13774_), .A2(pi0616), .ZN(new_n27609_));
  NOR2_X1    g25173(.A1(new_n27609_), .A2(new_n12821_), .ZN(new_n27610_));
  NOR2_X1    g25174(.A1(new_n27610_), .A2(new_n27389_), .ZN(new_n27611_));
  OAI22_X1   g25175(.A1(new_n27611_), .A2(new_n27608_), .B1(pi0662), .B2(new_n27392_), .ZN(new_n27612_));
  NAND2_X1   g25176(.A1(new_n27612_), .A2(new_n2631_), .ZN(new_n27613_));
  AOI21_X1   g25177(.A1(new_n27604_), .A2(new_n27613_), .B(new_n5445_), .ZN(new_n27614_));
  NOR2_X1    g25178(.A1(new_n26783_), .A2(new_n5405_), .ZN(new_n27615_));
  NOR2_X1    g25179(.A1(new_n26782_), .A2(new_n27615_), .ZN(new_n27616_));
  NOR2_X1    g25180(.A1(new_n27616_), .A2(new_n12821_), .ZN(new_n27617_));
  OAI21_X1   g25181(.A1(new_n27617_), .A2(new_n27385_), .B(pi0662), .ZN(new_n27618_));
  NAND2_X1   g25182(.A1(new_n27618_), .A2(new_n27386_), .ZN(new_n27619_));
  NOR2_X1    g25183(.A1(new_n27381_), .A2(new_n27602_), .ZN(new_n27620_));
  OAI21_X1   g25184(.A1(new_n27619_), .A2(new_n27620_), .B(pi0224), .ZN(new_n27621_));
  NAND2_X1   g25185(.A1(new_n27391_), .A2(new_n13169_), .ZN(new_n27622_));
  NOR2_X1    g25186(.A1(new_n24647_), .A2(new_n5405_), .ZN(new_n27623_));
  AOI21_X1   g25187(.A1(new_n27623_), .A2(new_n12821_), .B(new_n5400_), .ZN(new_n27624_));
  AOI21_X1   g25188(.A1(new_n27276_), .A2(new_n13779_), .B(new_n13096_), .ZN(new_n27625_));
  NOR2_X1    g25189(.A1(new_n13779_), .A2(new_n13111_), .ZN(new_n27626_));
  NOR2_X1    g25190(.A1(new_n27626_), .A2(pi0614), .ZN(new_n27627_));
  NOR2_X1    g25191(.A1(new_n26766_), .A2(new_n5405_), .ZN(new_n27628_));
  NOR2_X1    g25192(.A1(new_n27627_), .A2(new_n27628_), .ZN(new_n27629_));
  OR3_X2     g25193(.A1(new_n27629_), .A2(new_n12821_), .A3(new_n27625_), .Z(new_n27630_));
  AOI22_X1   g25194(.A1(new_n27630_), .A2(new_n27624_), .B1(new_n5400_), .B2(new_n27622_), .ZN(new_n27631_));
  NAND2_X1   g25195(.A1(new_n27631_), .A2(new_n2631_), .ZN(new_n27632_));
  AOI21_X1   g25196(.A1(new_n27621_), .A2(new_n27632_), .B(new_n5446_), .ZN(new_n27633_));
  NOR3_X1    g25197(.A1(new_n27633_), .A2(new_n27614_), .A3(new_n2668_), .ZN(new_n27634_));
  INV_X1     g25198(.I(new_n27404_), .ZN(new_n27635_));
  INV_X1     g25199(.I(new_n27401_), .ZN(new_n27636_));
  OAI21_X1   g25200(.A1(new_n13732_), .A2(new_n27593_), .B(new_n13111_), .ZN(new_n27637_));
  AOI21_X1   g25201(.A1(new_n27598_), .A2(new_n27637_), .B(new_n27636_), .ZN(new_n27638_));
  AOI22_X1   g25202(.A1(new_n27638_), .A2(pi0662), .B1(new_n13118_), .B2(new_n27635_), .ZN(new_n27639_));
  NAND2_X1   g25203(.A1(new_n27405_), .A2(new_n27601_), .ZN(new_n27640_));
  NAND2_X1   g25204(.A1(new_n27639_), .A2(new_n27640_), .ZN(new_n27641_));
  NAND2_X1   g25205(.A1(new_n27641_), .A2(new_n5446_), .ZN(new_n27642_));
  OAI22_X1   g25206(.A1(new_n26798_), .A2(new_n27411_), .B1(new_n26802_), .B2(new_n5405_), .ZN(new_n27643_));
  NOR2_X1    g25207(.A1(new_n27643_), .A2(new_n12821_), .ZN(new_n27644_));
  AOI21_X1   g25208(.A1(new_n26800_), .A2(new_n27644_), .B(new_n27416_), .ZN(new_n27645_));
  NAND2_X1   g25209(.A1(new_n27645_), .A2(pi0662), .ZN(new_n27646_));
  NAND2_X1   g25210(.A1(new_n27415_), .A2(new_n27601_), .ZN(new_n27647_));
  NAND3_X1   g25211(.A1(new_n27646_), .A2(new_n27418_), .A3(new_n27647_), .ZN(new_n27648_));
  NAND2_X1   g25212(.A1(new_n27648_), .A2(new_n5445_), .ZN(new_n27649_));
  AOI21_X1   g25213(.A1(new_n27649_), .A2(new_n27642_), .B(new_n2631_), .ZN(new_n27650_));
  NOR2_X1    g25214(.A1(new_n26833_), .A2(new_n27389_), .ZN(new_n27651_));
  OAI22_X1   g25215(.A1(new_n27651_), .A2(new_n27608_), .B1(pi0662), .B2(new_n27423_), .ZN(new_n27652_));
  NAND2_X1   g25216(.A1(new_n27652_), .A2(new_n5446_), .ZN(new_n27653_));
  OAI21_X1   g25217(.A1(new_n27425_), .A2(new_n27602_), .B(new_n27429_), .ZN(new_n27654_));
  NOR2_X1    g25218(.A1(new_n13770_), .A2(new_n13769_), .ZN(new_n27655_));
  NOR2_X1    g25219(.A1(new_n27655_), .A2(pi0614), .ZN(new_n27656_));
  AOI21_X1   g25220(.A1(new_n13617_), .A2(new_n13603_), .B(new_n5405_), .ZN(new_n27657_));
  OAI21_X1   g25221(.A1(new_n27656_), .A2(new_n27657_), .B(pi0680), .ZN(new_n27658_));
  NAND2_X1   g25222(.A1(new_n27658_), .A2(new_n27427_), .ZN(new_n27659_));
  AOI21_X1   g25223(.A1(new_n27659_), .A2(pi0662), .B(new_n27654_), .ZN(new_n27660_));
  NAND2_X1   g25224(.A1(new_n27660_), .A2(new_n5445_), .ZN(new_n27661_));
  AOI21_X1   g25225(.A1(new_n27661_), .A2(new_n27653_), .B(new_n5082_), .ZN(new_n27662_));
  NAND2_X1   g25226(.A1(new_n27605_), .A2(new_n27512_), .ZN(new_n27663_));
  AOI21_X1   g25227(.A1(new_n27663_), .A2(new_n27390_), .B(pi0224), .ZN(new_n27664_));
  AND2_X2    g25228(.A1(new_n27664_), .A2(new_n2629_), .Z(new_n27665_));
  NOR4_X1    g25229(.A1(new_n27650_), .A2(pi0223), .A3(new_n27662_), .A4(new_n27665_), .ZN(new_n27666_));
  OAI21_X1   g25230(.A1(new_n27666_), .A2(new_n27634_), .B(new_n2628_), .ZN(new_n27667_));
  NOR2_X1    g25231(.A1(new_n27612_), .A2(new_n6764_), .ZN(new_n27668_));
  NOR2_X1    g25232(.A1(new_n27631_), .A2(new_n5422_), .ZN(new_n27669_));
  OAI21_X1   g25233(.A1(new_n27669_), .A2(new_n27668_), .B(new_n2631_), .ZN(new_n27670_));
  OR3_X2     g25234(.A1(new_n27619_), .A2(new_n5422_), .A3(new_n27620_), .Z(new_n27671_));
  OAI21_X1   g25235(.A1(new_n6764_), .A2(new_n27603_), .B(new_n27671_), .ZN(new_n27672_));
  AOI21_X1   g25236(.A1(new_n27672_), .A2(pi0224), .B(new_n2436_), .ZN(new_n27673_));
  AOI21_X1   g25237(.A1(new_n27673_), .A2(new_n27670_), .B(new_n2628_), .ZN(new_n27674_));
  NAND3_X1   g25238(.A1(new_n13136_), .A2(new_n27372_), .A3(new_n27536_), .ZN(new_n27675_));
  NAND2_X1   g25239(.A1(new_n27596_), .A2(new_n27512_), .ZN(new_n27676_));
  NAND3_X1   g25240(.A1(new_n27676_), .A2(pi0224), .A3(new_n27675_), .ZN(new_n27677_));
  NOR2_X1    g25241(.A1(new_n27664_), .A2(new_n27436_), .ZN(new_n27678_));
  AOI21_X1   g25242(.A1(new_n27678_), .A2(new_n27677_), .B(pi0215), .ZN(new_n27679_));
  NAND2_X1   g25243(.A1(new_n27660_), .A2(new_n2631_), .ZN(new_n27680_));
  NAND2_X1   g25244(.A1(new_n27648_), .A2(pi0224), .ZN(new_n27681_));
  AOI21_X1   g25245(.A1(new_n27681_), .A2(new_n27680_), .B(new_n5422_), .ZN(new_n27682_));
  AOI21_X1   g25246(.A1(new_n27639_), .A2(new_n27640_), .B(new_n2631_), .ZN(new_n27683_));
  AOI21_X1   g25247(.A1(new_n2631_), .A2(new_n27652_), .B(new_n27683_), .ZN(new_n27684_));
  OAI21_X1   g25248(.A1(new_n27684_), .A2(new_n6764_), .B(new_n3304_), .ZN(new_n27685_));
  OAI21_X1   g25249(.A1(new_n27682_), .A2(new_n27685_), .B(new_n27679_), .ZN(new_n27686_));
  AOI21_X1   g25250(.A1(new_n27674_), .A2(new_n27686_), .B(new_n2627_), .ZN(new_n27687_));
  NOR2_X1    g25251(.A1(new_n27368_), .A2(new_n27512_), .ZN(new_n27688_));
  NOR3_X1    g25252(.A1(new_n27366_), .A2(pi0224), .A3(new_n13804_), .ZN(new_n27689_));
  NAND2_X1   g25253(.A1(new_n14553_), .A2(new_n5405_), .ZN(new_n27690_));
  AOI21_X1   g25254(.A1(new_n27690_), .A2(new_n26745_), .B(new_n2631_), .ZN(new_n27691_));
  NOR3_X1    g25255(.A1(new_n27689_), .A2(new_n27536_), .A3(new_n27691_), .ZN(new_n27692_));
  OAI21_X1   g25256(.A1(new_n27688_), .A2(new_n27692_), .B(pi0299), .ZN(new_n27693_));
  AOI21_X1   g25257(.A1(new_n13806_), .A2(new_n27512_), .B(new_n27361_), .ZN(new_n27694_));
  NOR2_X1    g25258(.A1(new_n27694_), .A2(pi0224), .ZN(new_n27695_));
  NOR2_X1    g25259(.A1(new_n26753_), .A2(new_n27512_), .ZN(new_n27696_));
  NOR3_X1    g25260(.A1(new_n27696_), .A2(new_n27195_), .A3(new_n27363_), .ZN(new_n27697_));
  OAI21_X1   g25261(.A1(new_n27695_), .A2(new_n27697_), .B(new_n2628_), .ZN(new_n27698_));
  NAND2_X1   g25262(.A1(new_n27693_), .A2(new_n27698_), .ZN(new_n27699_));
  AOI22_X1   g25263(.A1(new_n27667_), .A2(new_n27687_), .B1(new_n2627_), .B2(new_n27699_), .ZN(new_n27700_));
  AOI21_X1   g25264(.A1(new_n27700_), .A2(new_n3265_), .B(new_n2610_), .ZN(new_n27701_));
  AOI21_X1   g25265(.A1(new_n27701_), .A2(new_n27592_), .B(new_n27493_), .ZN(new_n27702_));
  NOR2_X1    g25266(.A1(new_n27702_), .A2(pi0778), .ZN(new_n27703_));
  INV_X1     g25267(.I(new_n27554_), .ZN(new_n27704_));
  NAND2_X1   g25268(.A1(new_n27454_), .A2(pi0625), .ZN(new_n27705_));
  OAI21_X1   g25269(.A1(new_n27702_), .A2(pi0625), .B(new_n27705_), .ZN(new_n27706_));
  AOI21_X1   g25270(.A1(new_n27706_), .A2(new_n12841_), .B(new_n27704_), .ZN(new_n27707_));
  NOR2_X1    g25271(.A1(new_n27702_), .A2(new_n13521_), .ZN(new_n27708_));
  AND2_X2    g25272(.A1(new_n27454_), .A2(new_n13521_), .Z(new_n27709_));
  OAI21_X1   g25273(.A1(new_n27709_), .A2(new_n27708_), .B(pi1153), .ZN(new_n27710_));
  AND2_X2    g25274(.A1(new_n27551_), .A2(pi0608), .Z(new_n27711_));
  AOI22_X1   g25275(.A1(new_n27707_), .A2(new_n13560_), .B1(new_n27710_), .B2(new_n27711_), .ZN(new_n27712_));
  AOI21_X1   g25276(.A1(new_n27712_), .A2(pi0778), .B(new_n27703_), .ZN(new_n27713_));
  NOR2_X1    g25277(.A1(new_n27713_), .A2(pi0785), .ZN(new_n27714_));
  NOR2_X1    g25278(.A1(new_n27556_), .A2(pi0609), .ZN(new_n27715_));
  NOR2_X1    g25279(.A1(new_n27713_), .A2(new_n12766_), .ZN(new_n27716_));
  OAI21_X1   g25280(.A1(new_n27716_), .A2(new_n27715_), .B(pi1155), .ZN(new_n27717_));
  NAND3_X1   g25281(.A1(new_n27717_), .A2(pi0660), .A3(new_n27462_), .ZN(new_n27718_));
  NAND3_X1   g25282(.A1(new_n27555_), .A2(pi0609), .A3(new_n27548_), .ZN(new_n27719_));
  OAI21_X1   g25283(.A1(new_n27713_), .A2(pi0609), .B(new_n27719_), .ZN(new_n27720_));
  AOI21_X1   g25284(.A1(new_n27720_), .A2(new_n12770_), .B(new_n27465_), .ZN(new_n27721_));
  AOI21_X1   g25285(.A1(new_n27721_), .A2(new_n13829_), .B(new_n12764_), .ZN(new_n27722_));
  AOI21_X1   g25286(.A1(new_n27722_), .A2(new_n27718_), .B(new_n27714_), .ZN(new_n27723_));
  OAI21_X1   g25287(.A1(new_n27470_), .A2(pi1154), .B(pi0627), .ZN(new_n27724_));
  AOI21_X1   g25288(.A1(new_n27558_), .A2(new_n12781_), .B(new_n12785_), .ZN(new_n27725_));
  NAND2_X1   g25289(.A1(new_n27723_), .A2(pi0618), .ZN(new_n27726_));
  AOI21_X1   g25290(.A1(new_n27726_), .A2(new_n27725_), .B(new_n27724_), .ZN(new_n27727_));
  OR2_X2     g25291(.A1(new_n27474_), .A2(pi0627), .Z(new_n27728_));
  AOI21_X1   g25292(.A1(new_n27558_), .A2(pi0618), .B(pi1154), .ZN(new_n27729_));
  INV_X1     g25293(.I(new_n27729_), .ZN(new_n27730_));
  AOI21_X1   g25294(.A1(new_n27723_), .A2(new_n12781_), .B(new_n27730_), .ZN(new_n27731_));
  OAI21_X1   g25295(.A1(new_n27731_), .A2(new_n27728_), .B(pi0781), .ZN(new_n27732_));
  OAI22_X1   g25296(.A1(new_n27732_), .A2(new_n27727_), .B1(pi0781), .B2(new_n27723_), .ZN(new_n27733_));
  AOI21_X1   g25297(.A1(new_n27733_), .A2(new_n12796_), .B(new_n14303_), .ZN(new_n27734_));
  INV_X1     g25298(.I(new_n27482_), .ZN(new_n27735_));
  NAND2_X1   g25299(.A1(new_n27733_), .A2(new_n12793_), .ZN(new_n27736_));
  NAND2_X1   g25300(.A1(new_n27561_), .A2(pi0619), .ZN(new_n27737_));
  AOI21_X1   g25301(.A1(new_n27736_), .A2(new_n27737_), .B(pi1159), .ZN(new_n27738_));
  NOR3_X1    g25302(.A1(new_n27738_), .A2(pi0648), .A3(new_n27735_), .ZN(new_n27739_));
  INV_X1     g25303(.I(new_n27479_), .ZN(new_n27740_));
  NOR2_X1    g25304(.A1(new_n27560_), .A2(pi0619), .ZN(new_n27741_));
  AOI21_X1   g25305(.A1(new_n27733_), .A2(pi0619), .B(new_n27741_), .ZN(new_n27742_));
  OAI21_X1   g25306(.A1(new_n27742_), .A2(new_n12791_), .B(pi0648), .ZN(new_n27743_));
  OAI21_X1   g25307(.A1(new_n27743_), .A2(new_n27740_), .B(pi0789), .ZN(new_n27744_));
  OAI21_X1   g25308(.A1(new_n27744_), .A2(new_n27739_), .B(new_n27734_), .ZN(new_n27745_));
  AOI22_X1   g25309(.A1(new_n27745_), .A2(new_n27590_), .B1(pi0792), .B2(new_n27580_), .ZN(new_n27746_));
  OAI21_X1   g25310(.A1(new_n27746_), .A2(new_n15341_), .B(new_n27573_), .ZN(new_n27747_));
  NAND2_X1   g25311(.A1(new_n27356_), .A2(pi0644), .ZN(new_n27748_));
  NOR2_X1    g25312(.A1(new_n27488_), .A2(new_n12984_), .ZN(new_n27749_));
  AOI21_X1   g25313(.A1(new_n12984_), .A2(new_n27356_), .B(new_n27749_), .ZN(new_n27750_));
  OAI21_X1   g25314(.A1(new_n27750_), .A2(pi0644), .B(new_n27748_), .ZN(new_n27751_));
  AOI21_X1   g25315(.A1(new_n27751_), .A2(pi0715), .B(pi1160), .ZN(new_n27752_));
  NOR3_X1    g25316(.A1(new_n27566_), .A2(new_n27570_), .A3(new_n12972_), .ZN(new_n27753_));
  NOR2_X1    g25317(.A1(new_n27563_), .A2(pi0787), .ZN(new_n27754_));
  NOR2_X1    g25318(.A1(new_n27753_), .A2(new_n27754_), .ZN(new_n27755_));
  OAI21_X1   g25319(.A1(new_n27755_), .A2(new_n12975_), .B(new_n12740_), .ZN(new_n27756_));
  NOR2_X1    g25320(.A1(new_n27747_), .A2(pi0644), .ZN(new_n27757_));
  OAI21_X1   g25321(.A1(new_n27757_), .A2(new_n27756_), .B(new_n27752_), .ZN(new_n27758_));
  NAND2_X1   g25322(.A1(new_n27356_), .A2(new_n12975_), .ZN(new_n27759_));
  OAI21_X1   g25323(.A1(new_n27750_), .A2(new_n12975_), .B(new_n27759_), .ZN(new_n27760_));
  AOI21_X1   g25324(.A1(new_n27760_), .A2(new_n12740_), .B(new_n12739_), .ZN(new_n27761_));
  NOR2_X1    g25325(.A1(new_n27755_), .A2(pi0644), .ZN(new_n27762_));
  NOR2_X1    g25326(.A1(new_n27762_), .A2(new_n12740_), .ZN(new_n27763_));
  OAI21_X1   g25327(.A1(new_n27747_), .A2(new_n12975_), .B(new_n27763_), .ZN(new_n27764_));
  AOI21_X1   g25328(.A1(new_n27764_), .A2(new_n27761_), .B(new_n13000_), .ZN(new_n27765_));
  AOI22_X1   g25329(.A1(new_n27765_), .A2(new_n27758_), .B1(new_n13000_), .B2(new_n27747_), .ZN(new_n27766_));
  OAI21_X1   g25330(.A1(new_n27766_), .A2(po1038), .B(new_n27355_), .ZN(po0381));
  NOR2_X1    g25331(.A1(new_n6173_), .A2(new_n3016_), .ZN(new_n27768_));
  INV_X1     g25332(.I(new_n27768_), .ZN(new_n27769_));
  NOR2_X1    g25333(.A1(new_n27769_), .A2(new_n3319_), .ZN(new_n27770_));
  AOI21_X1   g25334(.A1(new_n27770_), .A2(pi0062), .B(new_n3425_), .ZN(new_n27771_));
  INV_X1     g25335(.I(new_n6171_), .ZN(new_n27772_));
  NAND2_X1   g25336(.A1(new_n27768_), .A2(new_n2566_), .ZN(new_n27773_));
  AOI21_X1   g25337(.A1(new_n27773_), .A2(pi0054), .B(pi0074), .ZN(new_n27774_));
  NAND3_X1   g25338(.A1(new_n27768_), .A2(pi0092), .A3(new_n2564_), .ZN(new_n27775_));
  NAND2_X1   g25339(.A1(new_n27775_), .A2(new_n5499_), .ZN(new_n27776_));
  AOI21_X1   g25340(.A1(new_n5309_), .A2(new_n5350_), .B(pi0137), .ZN(new_n27777_));
  OAI21_X1   g25341(.A1(new_n9095_), .A2(new_n3016_), .B(new_n3265_), .ZN(new_n27778_));
  AOI21_X1   g25342(.A1(new_n2524_), .A2(new_n9203_), .B(new_n3068_), .ZN(new_n27779_));
  OR2_X2     g25343(.A1(new_n27779_), .A2(new_n3083_), .Z(new_n27780_));
  NOR2_X1    g25344(.A1(new_n6659_), .A2(new_n2726_), .ZN(new_n27781_));
  NAND4_X1   g25345(.A1(new_n27781_), .A2(pi0070), .A3(new_n2814_), .A4(new_n3083_), .ZN(new_n27782_));
  AOI21_X1   g25346(.A1(new_n27780_), .A2(new_n27782_), .B(new_n3038_), .ZN(new_n27783_));
  INV_X1     g25347(.I(new_n27783_), .ZN(new_n27784_));
  INV_X1     g25348(.I(new_n9350_), .ZN(new_n27785_));
  NAND2_X1   g25349(.A1(new_n3037_), .A2(new_n3083_), .ZN(new_n27786_));
  AOI21_X1   g25350(.A1(new_n2805_), .A2(new_n27781_), .B(pi0032), .ZN(new_n27787_));
  OAI21_X1   g25351(.A1(new_n27787_), .A2(new_n27786_), .B(new_n3041_), .ZN(new_n27788_));
  NOR2_X1    g25352(.A1(new_n3069_), .A2(new_n3083_), .ZN(new_n27789_));
  OR2_X2     g25353(.A1(new_n27788_), .A2(new_n27789_), .Z(new_n27790_));
  AOI21_X1   g25354(.A1(new_n3035_), .A2(new_n27781_), .B(pi0032), .ZN(new_n27791_));
  NOR2_X1    g25355(.A1(new_n27789_), .A2(new_n3041_), .ZN(new_n27792_));
  OAI21_X1   g25356(.A1(new_n27786_), .A2(new_n27791_), .B(new_n27792_), .ZN(new_n27793_));
  AOI21_X1   g25357(.A1(new_n27793_), .A2(new_n27790_), .B(new_n27785_), .ZN(new_n27794_));
  NOR2_X1    g25358(.A1(new_n27779_), .A2(new_n3038_), .ZN(new_n27795_));
  OAI22_X1   g25359(.A1(new_n27783_), .A2(new_n27788_), .B1(new_n3041_), .B2(new_n27795_), .ZN(new_n27796_));
  AOI22_X1   g25360(.A1(new_n27796_), .A2(new_n9344_), .B1(new_n27794_), .B2(new_n27784_), .ZN(new_n27797_));
  NOR3_X1    g25361(.A1(new_n2993_), .A2(new_n3191_), .A3(new_n9203_), .ZN(new_n27798_));
  OAI21_X1   g25362(.A1(new_n27798_), .A2(new_n3128_), .B(new_n2820_), .ZN(new_n27799_));
  AOI21_X1   g25363(.A1(new_n27799_), .A2(new_n3013_), .B(pi0095), .ZN(new_n27800_));
  OAI21_X1   g25364(.A1(new_n27800_), .A2(new_n3000_), .B(pi0137), .ZN(new_n27801_));
  AND2_X2    g25365(.A1(new_n27801_), .A2(new_n27797_), .Z(new_n27802_));
  OAI21_X1   g25366(.A1(new_n3014_), .A2(new_n3000_), .B(pi0137), .ZN(new_n27803_));
  INV_X1     g25367(.I(new_n9344_), .ZN(new_n27804_));
  NAND2_X1   g25368(.A1(new_n3069_), .A2(pi1093), .ZN(new_n27805_));
  AOI21_X1   g25369(.A1(new_n27790_), .A2(new_n27805_), .B(new_n27804_), .ZN(new_n27806_));
  NOR3_X1    g25370(.A1(new_n27794_), .A2(pi0332), .A3(new_n27806_), .ZN(new_n27807_));
  AOI22_X1   g25371(.A1(new_n27802_), .A2(pi0332), .B1(new_n27803_), .B2(new_n27807_), .ZN(new_n27808_));
  NAND2_X1   g25372(.A1(new_n27808_), .A2(new_n5504_), .ZN(new_n27809_));
  OAI21_X1   g25373(.A1(new_n27779_), .A2(new_n3038_), .B(new_n3016_), .ZN(new_n27810_));
  NAND3_X1   g25374(.A1(new_n27801_), .A2(pi0332), .A3(new_n27810_), .ZN(new_n27811_));
  NAND3_X1   g25375(.A1(new_n27803_), .A2(new_n2630_), .A3(new_n3070_), .ZN(new_n27812_));
  AND2_X2    g25376(.A1(new_n27811_), .A2(new_n27812_), .Z(new_n27813_));
  NAND2_X1   g25377(.A1(new_n27813_), .A2(new_n5306_), .ZN(new_n27814_));
  AOI21_X1   g25378(.A1(new_n27809_), .A2(new_n27814_), .B(pi0198), .ZN(new_n27815_));
  NAND2_X1   g25379(.A1(new_n27799_), .A2(new_n2754_), .ZN(new_n27816_));
  AOI21_X1   g25380(.A1(new_n27816_), .A2(new_n2462_), .B(new_n3163_), .ZN(new_n27817_));
  NOR4_X1    g25381(.A1(new_n27779_), .A2(pi0095), .A3(pi0137), .A4(new_n2753_), .ZN(new_n27818_));
  NOR3_X1    g25382(.A1(new_n27817_), .A2(new_n2630_), .A3(new_n27818_), .ZN(new_n27819_));
  AOI21_X1   g25383(.A1(new_n2997_), .A2(new_n3001_), .B(new_n3016_), .ZN(new_n27820_));
  OR2_X2     g25384(.A1(new_n27820_), .A2(new_n3062_), .Z(new_n27821_));
  AOI21_X1   g25385(.A1(new_n27821_), .A2(new_n2630_), .B(new_n27819_), .ZN(new_n27822_));
  OAI21_X1   g25386(.A1(new_n27822_), .A2(new_n2672_), .B(new_n2628_), .ZN(new_n27823_));
  NAND2_X1   g25387(.A1(new_n27808_), .A2(new_n2707_), .ZN(new_n27824_));
  NAND2_X1   g25388(.A1(new_n27813_), .A2(new_n2691_), .ZN(new_n27825_));
  AOI21_X1   g25389(.A1(new_n27824_), .A2(new_n27825_), .B(pi0210), .ZN(new_n27826_));
  OAI21_X1   g25390(.A1(new_n27822_), .A2(new_n2709_), .B(pi0299), .ZN(new_n27827_));
  OAI22_X1   g25391(.A1(new_n27815_), .A2(new_n27823_), .B1(new_n27826_), .B2(new_n27827_), .ZN(new_n27828_));
  AOI21_X1   g25392(.A1(new_n27828_), .A2(new_n2627_), .B(new_n27778_), .ZN(new_n27829_));
  OAI21_X1   g25393(.A1(new_n5346_), .A2(new_n3016_), .B(pi0038), .ZN(new_n27830_));
  NAND2_X1   g25394(.A1(new_n27830_), .A2(new_n2702_), .ZN(new_n27831_));
  OAI22_X1   g25395(.A1(new_n27829_), .A2(new_n27831_), .B1(new_n5339_), .B2(new_n27777_), .ZN(new_n27832_));
  NAND2_X1   g25396(.A1(new_n27769_), .A2(pi0087), .ZN(new_n27833_));
  OAI21_X1   g25397(.A1(new_n27832_), .A2(pi0087), .B(new_n27833_), .ZN(new_n27834_));
  OAI21_X1   g25398(.A1(new_n12043_), .A2(new_n27777_), .B(pi0075), .ZN(new_n27835_));
  NAND2_X1   g25399(.A1(new_n27835_), .A2(new_n3444_), .ZN(new_n27836_));
  AOI21_X1   g25400(.A1(new_n27834_), .A2(new_n3465_), .B(new_n27836_), .ZN(new_n27837_));
  OAI21_X1   g25401(.A1(new_n27837_), .A2(new_n27776_), .B(new_n27774_), .ZN(new_n27838_));
  NOR2_X1    g25402(.A1(new_n27769_), .A2(new_n6226_), .ZN(new_n27839_));
  AOI21_X1   g25403(.A1(new_n27839_), .A2(pi0074), .B(pi0055), .ZN(new_n27840_));
  AOI21_X1   g25404(.A1(new_n27838_), .A2(new_n27840_), .B(new_n27772_), .ZN(new_n27841_));
  NOR3_X1    g25405(.A1(new_n27769_), .A2(new_n3284_), .A3(new_n2571_), .ZN(new_n27842_));
  OAI21_X1   g25406(.A1(new_n27841_), .A2(new_n27842_), .B(new_n3471_), .ZN(new_n27843_));
  NOR3_X1    g25407(.A1(new_n27769_), .A2(pi0062), .A3(new_n3319_), .ZN(new_n27844_));
  OAI21_X1   g25408(.A1(new_n27844_), .A2(new_n3291_), .B(new_n5295_), .ZN(new_n27845_));
  AOI21_X1   g25409(.A1(new_n27843_), .A2(new_n27771_), .B(new_n27845_), .ZN(po0382));
  NAND2_X1   g25410(.A1(pi0228), .A2(pi0231), .ZN(new_n27847_));
  INV_X1     g25411(.I(new_n27847_), .ZN(new_n27848_));
  OAI21_X1   g25412(.A1(new_n27848_), .A2(new_n2602_), .B(new_n3284_), .ZN(new_n27849_));
  AOI21_X1   g25413(.A1(new_n6228_), .A2(new_n27847_), .B(new_n2625_), .ZN(new_n27850_));
  NAND2_X1   g25414(.A1(new_n27848_), .A2(pi0054), .ZN(new_n27851_));
  NAND3_X1   g25415(.A1(new_n10870_), .A2(pi0092), .A3(new_n27847_), .ZN(new_n27852_));
  OAI21_X1   g25416(.A1(new_n10872_), .A2(new_n27848_), .B(pi0075), .ZN(new_n27853_));
  NOR2_X1    g25417(.A1(new_n6234_), .A2(new_n3458_), .ZN(new_n27854_));
  AOI21_X1   g25418(.A1(new_n27854_), .A2(new_n27847_), .B(pi0075), .ZN(new_n27855_));
  OAI21_X1   g25419(.A1(new_n3212_), .A2(new_n2773_), .B(new_n2835_), .ZN(new_n27856_));
  AOI21_X1   g25420(.A1(new_n27856_), .A2(new_n2744_), .B(new_n2834_), .ZN(new_n27857_));
  OAI21_X1   g25421(.A1(new_n27857_), .A2(new_n3191_), .B(new_n2823_), .ZN(new_n27858_));
  AOI21_X1   g25422(.A1(new_n27858_), .A2(new_n2820_), .B(new_n5358_), .ZN(new_n27859_));
  OAI21_X1   g25423(.A1(new_n27859_), .A2(pi0095), .B(new_n3063_), .ZN(new_n27860_));
  NOR2_X1    g25424(.A1(new_n27860_), .A2(pi0039), .ZN(new_n27861_));
  NOR2_X1    g25425(.A1(new_n27861_), .A2(new_n3447_), .ZN(new_n27862_));
  NOR2_X1    g25426(.A1(new_n27862_), .A2(pi0038), .ZN(new_n27863_));
  NAND2_X1   g25427(.A1(new_n27863_), .A2(new_n2458_), .ZN(new_n27864_));
  AOI21_X1   g25428(.A1(new_n27864_), .A2(new_n27847_), .B(pi0100), .ZN(new_n27865_));
  AOI21_X1   g25429(.A1(new_n3322_), .A2(new_n2572_), .B(new_n27848_), .ZN(new_n27866_));
  OAI21_X1   g25430(.A1(new_n27866_), .A2(new_n2702_), .B(new_n3458_), .ZN(new_n27867_));
  OAI21_X1   g25431(.A1(new_n27865_), .A2(new_n27867_), .B(new_n27855_), .ZN(new_n27868_));
  NAND3_X1   g25432(.A1(new_n27868_), .A2(new_n3444_), .A3(new_n27853_), .ZN(new_n27869_));
  NAND3_X1   g25433(.A1(new_n27869_), .A2(new_n5499_), .A3(new_n27852_), .ZN(new_n27870_));
  AOI21_X1   g25434(.A1(new_n27870_), .A2(new_n27851_), .B(pi0074), .ZN(new_n27871_));
  NOR3_X1    g25435(.A1(new_n27871_), .A2(pi0055), .A3(new_n27850_), .ZN(new_n27872_));
  OAI21_X1   g25436(.A1(new_n3487_), .A2(new_n2577_), .B(new_n27847_), .ZN(new_n27873_));
  AOI21_X1   g25437(.A1(new_n27873_), .A2(pi0056), .B(pi0062), .ZN(new_n27874_));
  OAI21_X1   g25438(.A1(new_n27872_), .A2(new_n27849_), .B(new_n27874_), .ZN(new_n27875_));
  NAND3_X1   g25439(.A1(new_n6235_), .A2(pi0062), .A3(new_n27847_), .ZN(new_n27876_));
  NAND3_X1   g25440(.A1(new_n27875_), .A2(new_n3291_), .A3(new_n27876_), .ZN(new_n27877_));
  OAI21_X1   g25441(.A1(new_n3291_), .A2(new_n27847_), .B(new_n27877_), .ZN(po0383));
  NOR2_X1    g25442(.A1(new_n9233_), .A2(new_n8281_), .ZN(new_n27879_));
  NOR3_X1    g25443(.A1(new_n2758_), .A2(pi0824), .A3(new_n3082_), .ZN(new_n27880_));
  AOI21_X1   g25444(.A1(new_n8313_), .A2(new_n2755_), .B(pi0091), .ZN(new_n27881_));
  OAI21_X1   g25445(.A1(new_n8931_), .A2(new_n8913_), .B(new_n27881_), .ZN(new_n27882_));
  AOI21_X1   g25446(.A1(new_n8925_), .A2(new_n27880_), .B(new_n27882_), .ZN(new_n27883_));
  NOR2_X1    g25447(.A1(new_n5561_), .A2(new_n2749_), .ZN(new_n27884_));
  INV_X1     g25448(.I(new_n27884_), .ZN(new_n27885_));
  OAI21_X1   g25449(.A1(new_n27883_), .A2(new_n27885_), .B(new_n2821_), .ZN(new_n27886_));
  AOI21_X1   g25450(.A1(new_n27886_), .A2(new_n5558_), .B(new_n5429_), .ZN(new_n27887_));
  OAI21_X1   g25451(.A1(new_n27885_), .A2(new_n27881_), .B(new_n2821_), .ZN(new_n27888_));
  NOR2_X1    g25452(.A1(new_n27885_), .A2(new_n8931_), .ZN(new_n27889_));
  NOR2_X1    g25453(.A1(new_n27888_), .A2(new_n27889_), .ZN(new_n27890_));
  NOR2_X1    g25454(.A1(new_n27890_), .A2(new_n5559_), .ZN(new_n27891_));
  INV_X1     g25455(.I(new_n27888_), .ZN(new_n27892_));
  AOI22_X1   g25456(.A1(new_n27889_), .A2(new_n6259_), .B1(pi0829), .B2(new_n3041_), .ZN(new_n27893_));
  AOI21_X1   g25457(.A1(new_n27893_), .A2(new_n27892_), .B(new_n5559_), .ZN(new_n27894_));
  INV_X1     g25458(.I(new_n5539_), .ZN(new_n27895_));
  NAND4_X1   g25459(.A1(new_n5558_), .A2(new_n2748_), .A3(new_n6258_), .A4(new_n10327_), .ZN(new_n27896_));
  AOI21_X1   g25460(.A1(new_n27896_), .A2(new_n27895_), .B(new_n3041_), .ZN(new_n27897_));
  OAI22_X1   g25461(.A1(new_n27894_), .A2(new_n27897_), .B1(new_n10302_), .B2(new_n27891_), .ZN(new_n27898_));
  AOI21_X1   g25462(.A1(pi0829), .A2(new_n27887_), .B(new_n27898_), .ZN(new_n27899_));
  OAI21_X1   g25463(.A1(new_n27899_), .A2(pi0039), .B(new_n27879_), .ZN(po0384));
  OAI21_X1   g25464(.A1(new_n3080_), .A2(new_n7287_), .B(new_n2769_), .ZN(new_n27901_));
  NOR4_X1    g25465(.A1(new_n27901_), .A2(pi0032), .A3(pi0039), .A4(pi0095), .ZN(new_n27902_));
  NOR3_X1    g25466(.A1(new_n5527_), .A2(new_n3022_), .A3(new_n9211_), .ZN(new_n27903_));
  NOR2_X1    g25467(.A1(new_n9207_), .A2(new_n9208_), .ZN(new_n27904_));
  NOR2_X1    g25468(.A1(new_n27904_), .A2(new_n2627_), .ZN(new_n27905_));
  AOI22_X1   g25469(.A1(new_n27902_), .A2(new_n9252_), .B1(new_n27903_), .B2(new_n27905_), .ZN(new_n27906_));
  OAI22_X1   g25470(.A1(new_n27906_), .A2(new_n8281_), .B1(pi0039), .B2(new_n2458_), .ZN(po0385));
  NOR2_X1    g25471(.A1(new_n13019_), .A2(pi0047), .ZN(new_n27908_));
  NAND2_X1   g25472(.A1(new_n13016_), .A2(new_n5353_), .ZN(new_n27909_));
  OAI21_X1   g25473(.A1(new_n27908_), .A2(new_n27909_), .B(new_n2818_), .ZN(new_n27910_));
  NAND3_X1   g25474(.A1(new_n27910_), .A2(new_n2525_), .A3(new_n13044_), .ZN(new_n27911_));
  AOI21_X1   g25475(.A1(new_n27911_), .A2(pi0252), .B(new_n5331_), .ZN(new_n27912_));
  AOI21_X1   g25476(.A1(new_n27912_), .A2(new_n13013_), .B(pi1093), .ZN(new_n27913_));
  NAND2_X1   g25477(.A1(new_n13023_), .A2(new_n5331_), .ZN(new_n27914_));
  AOI21_X1   g25478(.A1(new_n27914_), .A2(new_n27913_), .B(pi0039), .ZN(new_n27915_));
  AOI21_X1   g25479(.A1(new_n6259_), .A2(new_n13023_), .B(new_n13035_), .ZN(new_n27916_));
  NOR3_X1    g25480(.A1(new_n27916_), .A2(new_n5351_), .A3(new_n5533_), .ZN(new_n27917_));
  NOR2_X1    g25481(.A1(new_n27917_), .A2(new_n3041_), .ZN(new_n27918_));
  NOR2_X1    g25482(.A1(new_n13046_), .A2(new_n5428_), .ZN(new_n27919_));
  NOR2_X1    g25483(.A1(new_n3044_), .A2(new_n3022_), .ZN(new_n27920_));
  AOI21_X1   g25484(.A1(new_n13050_), .A2(new_n27920_), .B(pi0824), .ZN(new_n27921_));
  NOR3_X1    g25485(.A1(new_n27921_), .A2(new_n27919_), .A3(new_n5533_), .ZN(new_n27922_));
  NOR2_X1    g25486(.A1(new_n27922_), .A2(new_n13023_), .ZN(new_n27923_));
  NOR4_X1    g25487(.A1(new_n13050_), .A2(pi0824), .A3(new_n3044_), .A4(new_n3022_), .ZN(new_n27924_));
  OAI21_X1   g25488(.A1(new_n27924_), .A2(new_n27919_), .B(new_n8913_), .ZN(new_n27925_));
  AOI21_X1   g25489(.A1(new_n27925_), .A2(new_n5351_), .B(new_n5533_), .ZN(new_n27926_));
  OAI21_X1   g25490(.A1(new_n27926_), .A2(new_n27923_), .B(new_n27918_), .ZN(new_n27927_));
  NAND2_X1   g25491(.A1(new_n5434_), .A2(pi0120), .ZN(new_n27928_));
  OAI21_X1   g25492(.A1(new_n6745_), .A2(new_n27928_), .B(new_n13087_), .ZN(new_n27929_));
  NAND2_X1   g25493(.A1(new_n27929_), .A2(new_n5422_), .ZN(new_n27930_));
  OAI21_X1   g25494(.A1(new_n5413_), .A2(new_n27928_), .B(new_n13087_), .ZN(new_n27931_));
  NAND2_X1   g25495(.A1(new_n27931_), .A2(new_n6764_), .ZN(new_n27932_));
  AOI21_X1   g25496(.A1(new_n27930_), .A2(new_n27932_), .B(new_n2436_), .ZN(new_n27933_));
  OAI21_X1   g25497(.A1(new_n13221_), .A2(new_n3304_), .B(new_n2436_), .ZN(new_n27934_));
  NOR2_X1    g25498(.A1(new_n13085_), .A2(new_n5528_), .ZN(new_n27935_));
  NOR2_X1    g25499(.A1(new_n13295_), .A2(new_n5529_), .ZN(new_n27936_));
  OAI21_X1   g25500(.A1(new_n27935_), .A2(new_n27936_), .B(new_n3022_), .ZN(new_n27937_));
  AOI21_X1   g25501(.A1(new_n13137_), .A2(new_n6712_), .B(new_n13085_), .ZN(new_n27938_));
  NOR3_X1    g25502(.A1(new_n13295_), .A2(new_n5329_), .A3(new_n6713_), .ZN(new_n27939_));
  OAI21_X1   g25503(.A1(new_n27938_), .A2(new_n27939_), .B(pi1091), .ZN(new_n27940_));
  NAND3_X1   g25504(.A1(new_n27940_), .A2(new_n10903_), .A3(new_n27937_), .ZN(new_n27941_));
  AND2_X2    g25505(.A1(new_n27941_), .A2(new_n13084_), .Z(new_n27942_));
  NAND2_X1   g25506(.A1(new_n27942_), .A2(new_n5427_), .ZN(new_n27943_));
  OAI21_X1   g25507(.A1(new_n5427_), .A2(new_n13087_), .B(new_n27943_), .ZN(new_n27944_));
  OR2_X2     g25508(.A1(new_n27944_), .A2(new_n5422_), .Z(new_n27945_));
  NAND2_X1   g25509(.A1(new_n27942_), .A2(new_n5449_), .ZN(new_n27946_));
  OAI21_X1   g25510(.A1(new_n5449_), .A2(new_n13087_), .B(new_n27946_), .ZN(new_n27947_));
  OR2_X2     g25511(.A1(new_n27947_), .A2(new_n6764_), .Z(new_n27948_));
  AOI21_X1   g25512(.A1(new_n27945_), .A2(new_n27948_), .B(new_n3303_), .ZN(new_n27949_));
  OAI21_X1   g25513(.A1(new_n27949_), .A2(new_n27934_), .B(pi0299), .ZN(new_n27950_));
  OR2_X2     g25514(.A1(new_n27944_), .A2(new_n5446_), .Z(new_n27951_));
  OR2_X2     g25515(.A1(new_n27947_), .A2(new_n5445_), .Z(new_n27952_));
  AOI21_X1   g25516(.A1(new_n27951_), .A2(new_n27952_), .B(new_n2641_), .ZN(new_n27953_));
  OAI21_X1   g25517(.A1(new_n13221_), .A2(new_n2642_), .B(new_n2668_), .ZN(new_n27954_));
  NAND2_X1   g25518(.A1(new_n27929_), .A2(new_n5446_), .ZN(new_n27955_));
  NAND2_X1   g25519(.A1(new_n27931_), .A2(new_n5445_), .ZN(new_n27956_));
  NAND2_X1   g25520(.A1(new_n27955_), .A2(new_n27956_), .ZN(new_n27957_));
  AOI21_X1   g25521(.A1(new_n27957_), .A2(pi0223), .B(pi0299), .ZN(new_n27958_));
  OAI21_X1   g25522(.A1(new_n27953_), .A2(new_n27954_), .B(new_n27958_), .ZN(new_n27959_));
  OAI21_X1   g25523(.A1(new_n27933_), .A2(new_n27950_), .B(new_n27959_), .ZN(new_n27960_));
  AOI22_X1   g25524(.A1(new_n27960_), .A2(pi0039), .B1(new_n27915_), .B2(new_n27927_), .ZN(new_n27961_));
  OAI21_X1   g25525(.A1(new_n5345_), .A2(new_n3265_), .B(new_n8264_), .ZN(new_n27962_));
  AOI21_X1   g25526(.A1(new_n27961_), .A2(new_n3265_), .B(new_n27962_), .ZN(po0387));
  INV_X1     g25527(.I(new_n2863_), .ZN(new_n27964_));
  NAND3_X1   g25528(.A1(new_n2959_), .A2(new_n2500_), .A3(new_n2893_), .ZN(new_n27965_));
  AOI21_X1   g25529(.A1(new_n27965_), .A2(new_n9178_), .B(pi0102), .ZN(new_n27966_));
  OAI21_X1   g25530(.A1(new_n27966_), .A2(new_n2850_), .B(new_n2889_), .ZN(new_n27967_));
  AOI21_X1   g25531(.A1(new_n27967_), .A2(new_n2883_), .B(new_n5593_), .ZN(new_n27968_));
  OAI21_X1   g25532(.A1(new_n27968_), .A2(new_n2880_), .B(new_n5566_), .ZN(new_n27969_));
  AOI21_X1   g25533(.A1(new_n27969_), .A2(new_n2879_), .B(new_n5563_), .ZN(new_n27970_));
  OAI21_X1   g25534(.A1(new_n27970_), .A2(new_n2877_), .B(new_n10883_), .ZN(new_n27971_));
  AOI21_X1   g25535(.A1(new_n27971_), .A2(new_n2849_), .B(new_n27964_), .ZN(new_n27972_));
  OAI21_X1   g25536(.A1(new_n27972_), .A2(new_n2981_), .B(new_n5366_), .ZN(new_n27973_));
  AOI21_X1   g25537(.A1(new_n27973_), .A2(new_n2847_), .B(new_n12052_), .ZN(new_n27974_));
  OAI21_X1   g25538(.A1(new_n27974_), .A2(new_n2841_), .B(new_n2987_), .ZN(new_n27975_));
  OAI22_X1   g25539(.A1(new_n27975_), .A2(new_n2537_), .B1(new_n2548_), .B2(new_n12049_), .ZN(new_n27976_));
  OAI21_X1   g25540(.A1(new_n27976_), .A2(pi0070), .B(new_n3192_), .ZN(new_n27977_));
  AOI21_X1   g25541(.A1(new_n27977_), .A2(new_n2744_), .B(new_n2834_), .ZN(new_n27978_));
  OAI21_X1   g25542(.A1(new_n27978_), .A2(new_n3191_), .B(new_n2823_), .ZN(new_n27979_));
  INV_X1     g25543(.I(pi1082), .ZN(new_n27980_));
  AOI21_X1   g25544(.A1(new_n2819_), .A2(new_n27980_), .B(pi0032), .ZN(new_n27981_));
  AOI22_X1   g25545(.A1(new_n27979_), .A2(new_n27981_), .B1(pi0032), .B2(new_n3178_), .ZN(new_n27982_));
  OAI21_X1   g25546(.A1(new_n27982_), .A2(pi0095), .B(new_n3001_), .ZN(new_n27983_));
  OAI21_X1   g25547(.A1(new_n27983_), .A2(pi0039), .B(new_n9095_), .ZN(new_n27984_));
  NOR2_X1    g25548(.A1(new_n5452_), .A2(pi0299), .ZN(new_n27985_));
  AOI21_X1   g25549(.A1(new_n6809_), .A2(pi0299), .B(new_n27985_), .ZN(new_n27986_));
  NAND4_X1   g25550(.A1(new_n27986_), .A2(pi0835), .A3(new_n5391_), .A4(new_n5432_), .ZN(new_n27987_));
  NAND4_X1   g25551(.A1(new_n27987_), .A2(pi0039), .A3(new_n5393_), .A4(new_n8303_), .ZN(new_n27988_));
  NAND3_X1   g25552(.A1(new_n27984_), .A2(new_n3265_), .A3(new_n27988_), .ZN(new_n27989_));
  NAND2_X1   g25553(.A1(new_n27989_), .A2(new_n5348_), .ZN(new_n27990_));
  AOI21_X1   g25554(.A1(new_n27990_), .A2(new_n2702_), .B(pi0087), .ZN(new_n27991_));
  AOI21_X1   g25555(.A1(new_n27991_), .A2(new_n5339_), .B(new_n5302_), .ZN(new_n27992_));
  OAI21_X1   g25556(.A1(new_n27992_), .A2(new_n2606_), .B(new_n6180_), .ZN(new_n27993_));
  AOI21_X1   g25557(.A1(new_n27993_), .A2(new_n5499_), .B(new_n6175_), .ZN(new_n27994_));
  OAI21_X1   g25558(.A1(new_n27994_), .A2(new_n7264_), .B(new_n12102_), .ZN(new_n27995_));
  AOI21_X1   g25559(.A1(new_n27995_), .A2(new_n3284_), .B(new_n5298_), .ZN(new_n27996_));
  OAI21_X1   g25560(.A1(new_n27996_), .A2(pi0062), .B(new_n5465_), .ZN(new_n27997_));
  AOI21_X1   g25561(.A1(new_n27997_), .A2(new_n3291_), .B(new_n5296_), .ZN(po0389));
  INV_X1     g25562(.I(pi0230), .ZN(new_n27999_));
  NOR2_X1    g25563(.A1(new_n8511_), .A2(pi0211), .ZN(new_n28000_));
  INV_X1     g25564(.I(new_n28000_), .ZN(new_n28001_));
  OAI21_X1   g25565(.A1(new_n28001_), .A2(new_n12770_), .B(new_n8509_), .ZN(new_n28002_));
  NOR2_X1    g25566(.A1(new_n12785_), .A2(pi0211), .ZN(new_n28003_));
  INV_X1     g25567(.I(new_n28003_), .ZN(new_n28004_));
  NOR2_X1    g25568(.A1(new_n12841_), .A2(pi0211), .ZN(new_n28005_));
  NOR2_X1    g25569(.A1(new_n8811_), .A2(new_n28005_), .ZN(new_n28006_));
  AOI21_X1   g25570(.A1(new_n8511_), .A2(new_n28004_), .B(new_n28006_), .ZN(new_n28007_));
  NAND2_X1   g25571(.A1(new_n28007_), .A2(new_n28002_), .ZN(new_n28008_));
  AOI21_X1   g25572(.A1(new_n28008_), .A2(pi0219), .B(new_n6643_), .ZN(new_n28009_));
  NOR2_X1    g25573(.A1(new_n12770_), .A2(pi0211), .ZN(new_n28010_));
  NOR2_X1    g25574(.A1(new_n8510_), .A2(new_n12785_), .ZN(new_n28011_));
  NOR3_X1    g25575(.A1(new_n28011_), .A2(new_n28010_), .A3(new_n8511_), .ZN(new_n28012_));
  NOR2_X1    g25576(.A1(new_n12742_), .A2(pi0211), .ZN(new_n28013_));
  NOR2_X1    g25577(.A1(new_n8510_), .A2(new_n12770_), .ZN(new_n28014_));
  NOR3_X1    g25578(.A1(new_n28014_), .A2(new_n28013_), .A3(pi0214), .ZN(new_n28015_));
  NOR3_X1    g25579(.A1(new_n28012_), .A2(new_n28015_), .A3(new_n8509_), .ZN(new_n28016_));
  NOR2_X1    g25580(.A1(new_n8510_), .A2(new_n12742_), .ZN(new_n28017_));
  NOR2_X1    g25581(.A1(new_n12965_), .A2(pi0211), .ZN(new_n28018_));
  NOR2_X1    g25582(.A1(new_n28017_), .A2(new_n28018_), .ZN(new_n28019_));
  NOR2_X1    g25583(.A1(new_n8511_), .A2(pi0212), .ZN(new_n28020_));
  INV_X1     g25584(.I(new_n28020_), .ZN(new_n28021_));
  NOR2_X1    g25585(.A1(new_n28019_), .A2(new_n28021_), .ZN(new_n28022_));
  NOR2_X1    g25586(.A1(new_n28016_), .A2(new_n28022_), .ZN(new_n28023_));
  NAND2_X1   g25587(.A1(new_n28023_), .A2(new_n8807_), .ZN(new_n28024_));
  AOI21_X1   g25588(.A1(new_n28009_), .A2(new_n28024_), .B(pi0213), .ZN(new_n28025_));
  NOR2_X1    g25589(.A1(new_n8521_), .A2(pi0299), .ZN(new_n28026_));
  INV_X1     g25590(.I(new_n28026_), .ZN(new_n28027_));
  NOR2_X1    g25591(.A1(new_n3768_), .A2(pi0199), .ZN(new_n28028_));
  NOR2_X1    g25592(.A1(new_n28028_), .A2(new_n8531_), .ZN(new_n28029_));
  AOI21_X1   g25593(.A1(pi0199), .A2(pi1142), .B(pi0200), .ZN(new_n28030_));
  INV_X1     g25594(.I(new_n28030_), .ZN(new_n28031_));
  NOR2_X1    g25595(.A1(new_n3605_), .A2(pi0199), .ZN(new_n28032_));
  NOR2_X1    g25596(.A1(new_n28031_), .A2(new_n28032_), .ZN(new_n28033_));
  NOR3_X1    g25597(.A1(new_n28033_), .A2(new_n28027_), .A3(new_n28029_), .ZN(new_n28034_));
  NOR2_X1    g25598(.A1(new_n28032_), .A2(new_n8531_), .ZN(new_n28035_));
  INV_X1     g25599(.I(new_n28035_), .ZN(new_n28036_));
  OAI21_X1   g25600(.A1(pi0199), .A2(new_n2446_), .B(new_n28030_), .ZN(new_n28037_));
  NAND2_X1   g25601(.A1(new_n28036_), .A2(new_n28037_), .ZN(new_n28038_));
  AOI21_X1   g25602(.A1(new_n28038_), .A2(new_n2628_), .B(pi0207), .ZN(new_n28039_));
  OAI21_X1   g25603(.A1(new_n28039_), .A2(new_n28034_), .B(pi0208), .ZN(new_n28040_));
  NOR2_X1    g25604(.A1(new_n8521_), .A2(pi0208), .ZN(new_n28041_));
  NAND3_X1   g25605(.A1(new_n28036_), .A2(new_n28037_), .A3(new_n28041_), .ZN(new_n28042_));
  AOI21_X1   g25606(.A1(new_n28040_), .A2(new_n28042_), .B(pi0299), .ZN(new_n28043_));
  INV_X1     g25607(.I(new_n8808_), .ZN(new_n28044_));
  INV_X1     g25608(.I(new_n10289_), .ZN(new_n28045_));
  NOR2_X1    g25609(.A1(new_n2628_), .A2(new_n12841_), .ZN(new_n28046_));
  NAND2_X1   g25610(.A1(new_n28046_), .A2(pi0214), .ZN(new_n28047_));
  NOR2_X1    g25611(.A1(new_n2628_), .A2(new_n12785_), .ZN(new_n28048_));
  NAND2_X1   g25612(.A1(new_n28048_), .A2(new_n8511_), .ZN(new_n28049_));
  NAND2_X1   g25613(.A1(new_n28047_), .A2(new_n28049_), .ZN(new_n28050_));
  NOR2_X1    g25614(.A1(new_n2628_), .A2(new_n12770_), .ZN(new_n28051_));
  AOI22_X1   g25615(.A1(new_n28050_), .A2(pi0212), .B1(new_n28020_), .B2(new_n28051_), .ZN(new_n28052_));
  OAI22_X1   g25616(.A1(new_n28044_), .A2(new_n28052_), .B1(new_n28023_), .B2(new_n28045_), .ZN(new_n28053_));
  OAI21_X1   g25617(.A1(new_n28043_), .A2(new_n28053_), .B(new_n6643_), .ZN(new_n28054_));
  NAND2_X1   g25618(.A1(new_n28054_), .A2(new_n28025_), .ZN(new_n28055_));
  NOR2_X1    g25619(.A1(pi0212), .A2(pi0214), .ZN(new_n28056_));
  NOR2_X1    g25620(.A1(new_n28056_), .A2(pi0211), .ZN(new_n28057_));
  NOR2_X1    g25621(.A1(new_n28057_), .A2(new_n8807_), .ZN(new_n28058_));
  NOR2_X1    g25622(.A1(new_n6643_), .A2(new_n28058_), .ZN(new_n28059_));
  INV_X1     g25623(.I(new_n28059_), .ZN(new_n28060_));
  NOR2_X1    g25624(.A1(new_n8510_), .A2(pi1143), .ZN(new_n28061_));
  NOR2_X1    g25625(.A1(pi0211), .A2(pi1144), .ZN(new_n28062_));
  NOR2_X1    g25626(.A1(new_n28061_), .A2(new_n28062_), .ZN(new_n28063_));
  INV_X1     g25627(.I(new_n28063_), .ZN(new_n28064_));
  NOR2_X1    g25628(.A1(new_n8809_), .A2(new_n28056_), .ZN(new_n28065_));
  INV_X1     g25629(.I(new_n28065_), .ZN(new_n28066_));
  NOR2_X1    g25630(.A1(new_n3605_), .A2(pi0211), .ZN(new_n28067_));
  INV_X1     g25631(.I(new_n28067_), .ZN(new_n28068_));
  OAI22_X1   g25632(.A1(new_n28066_), .A2(new_n28064_), .B1(new_n8811_), .B2(new_n28068_), .ZN(new_n28069_));
  NAND2_X1   g25633(.A1(new_n28069_), .A2(new_n8807_), .ZN(new_n28070_));
  NOR2_X1    g25634(.A1(new_n8515_), .A2(new_n3768_), .ZN(new_n28071_));
  INV_X1     g25635(.I(new_n28071_), .ZN(new_n28072_));
  AOI21_X1   g25636(.A1(new_n28070_), .A2(new_n28072_), .B(new_n28060_), .ZN(new_n28073_));
  NOR2_X1    g25637(.A1(new_n28064_), .A2(new_n2628_), .ZN(new_n28074_));
  INV_X1     g25638(.I(new_n28074_), .ZN(new_n28075_));
  NOR2_X1    g25639(.A1(new_n28075_), .A2(new_n8511_), .ZN(new_n28076_));
  OAI21_X1   g25640(.A1(new_n28043_), .A2(new_n28076_), .B(new_n8509_), .ZN(new_n28077_));
  NOR2_X1    g25641(.A1(new_n8510_), .A2(pi1142), .ZN(new_n28078_));
  NOR2_X1    g25642(.A1(pi0211), .A2(pi1143), .ZN(new_n28079_));
  NOR3_X1    g25643(.A1(new_n28078_), .A2(new_n2628_), .A3(new_n28079_), .ZN(new_n28080_));
  NOR3_X1    g25644(.A1(new_n28043_), .A2(new_n8511_), .A3(new_n28080_), .ZN(new_n28081_));
  NOR2_X1    g25645(.A1(new_n28081_), .A2(new_n8509_), .ZN(new_n28082_));
  INV_X1     g25646(.I(new_n28043_), .ZN(new_n28083_));
  NAND3_X1   g25647(.A1(new_n28083_), .A2(new_n8511_), .A3(new_n28075_), .ZN(new_n28084_));
  AOI21_X1   g25648(.A1(new_n28082_), .A2(new_n28084_), .B(pi0219), .ZN(new_n28085_));
  AOI21_X1   g25649(.A1(new_n28085_), .A2(new_n28077_), .B(po1038), .ZN(new_n28086_));
  NOR2_X1    g25650(.A1(new_n2628_), .A2(new_n3768_), .ZN(new_n28087_));
  NAND2_X1   g25651(.A1(new_n28057_), .A2(new_n28087_), .ZN(new_n28088_));
  NAND3_X1   g25652(.A1(new_n28083_), .A2(pi0219), .A3(new_n28088_), .ZN(new_n28089_));
  AOI21_X1   g25653(.A1(new_n28086_), .A2(new_n28089_), .B(new_n28073_), .ZN(new_n28090_));
  NAND2_X1   g25654(.A1(new_n28090_), .A2(pi0213), .ZN(new_n28091_));
  NAND3_X1   g25655(.A1(new_n28091_), .A2(pi0209), .A3(new_n28055_), .ZN(new_n28092_));
  INV_X1     g25656(.I(new_n28073_), .ZN(new_n28093_));
  NOR2_X1    g25657(.A1(new_n28056_), .A2(pi0219), .ZN(new_n28094_));
  NOR2_X1    g25658(.A1(new_n28057_), .A2(new_n28094_), .ZN(new_n28095_));
  NOR2_X1    g25659(.A1(pi0207), .A2(pi0299), .ZN(new_n28096_));
  NOR2_X1    g25660(.A1(new_n28096_), .A2(pi0208), .ZN(new_n28097_));
  INV_X1     g25661(.I(new_n28097_), .ZN(new_n28098_));
  NOR2_X1    g25662(.A1(new_n12770_), .A2(pi0200), .ZN(new_n28099_));
  NOR2_X1    g25663(.A1(new_n9172_), .A2(new_n28099_), .ZN(new_n28100_));
  NOR2_X1    g25664(.A1(new_n28100_), .A2(new_n12742_), .ZN(new_n28101_));
  NOR2_X1    g25665(.A1(new_n8531_), .A2(pi0299), .ZN(new_n28102_));
  NOR2_X1    g25666(.A1(new_n28102_), .A2(new_n12770_), .ZN(new_n28103_));
  NOR2_X1    g25667(.A1(new_n8780_), .A2(pi1155), .ZN(new_n28104_));
  NOR2_X1    g25668(.A1(new_n28104_), .A2(new_n28103_), .ZN(new_n28105_));
  INV_X1     g25669(.I(new_n28105_), .ZN(new_n28106_));
  AOI21_X1   g25670(.A1(new_n28106_), .A2(new_n12742_), .B(new_n28101_), .ZN(new_n28107_));
  AOI21_X1   g25671(.A1(new_n28107_), .A2(pi0207), .B(new_n28098_), .ZN(new_n28108_));
  NOR2_X1    g25672(.A1(new_n28108_), .A2(new_n12965_), .ZN(new_n28109_));
  INV_X1     g25673(.I(new_n28099_), .ZN(new_n28110_));
  NOR3_X1    g25674(.A1(new_n28110_), .A2(new_n8525_), .A3(pi0299), .ZN(new_n28111_));
  NOR2_X1    g25675(.A1(new_n8531_), .A2(pi0199), .ZN(new_n28112_));
  NOR2_X1    g25676(.A1(new_n28112_), .A2(pi0299), .ZN(new_n28113_));
  INV_X1     g25677(.I(new_n28113_), .ZN(new_n28114_));
  AOI21_X1   g25678(.A1(pi1156), .A2(new_n28114_), .B(new_n28111_), .ZN(new_n28115_));
  INV_X1     g25679(.I(new_n28115_), .ZN(new_n28116_));
  AOI21_X1   g25680(.A1(new_n28116_), .A2(pi0207), .B(pi0299), .ZN(new_n28117_));
  NOR2_X1    g25681(.A1(new_n28117_), .A2(pi0208), .ZN(new_n28118_));
  NOR2_X1    g25682(.A1(new_n28118_), .A2(pi1157), .ZN(new_n28119_));
  NOR2_X1    g25683(.A1(new_n2628_), .A2(pi1142), .ZN(new_n28120_));
  NOR3_X1    g25684(.A1(new_n28119_), .A2(new_n28109_), .A3(new_n28120_), .ZN(new_n28121_));
  INV_X1     g25685(.I(new_n28120_), .ZN(new_n28122_));
  NOR2_X1    g25686(.A1(new_n8525_), .A2(pi0200), .ZN(new_n28123_));
  NOR2_X1    g25687(.A1(new_n28112_), .A2(new_n28123_), .ZN(new_n28124_));
  NOR2_X1    g25688(.A1(new_n28124_), .A2(pi0299), .ZN(new_n28125_));
  INV_X1     g25689(.I(new_n28125_), .ZN(new_n28126_));
  NOR2_X1    g25690(.A1(new_n8525_), .A2(pi1153), .ZN(new_n28127_));
  NOR2_X1    g25691(.A1(new_n28126_), .A2(new_n28127_), .ZN(new_n28128_));
  NOR2_X1    g25692(.A1(new_n9171_), .A2(new_n12770_), .ZN(new_n28129_));
  NOR2_X1    g25693(.A1(new_n28128_), .A2(new_n28129_), .ZN(new_n28130_));
  INV_X1     g25694(.I(new_n28130_), .ZN(new_n28131_));
  INV_X1     g25695(.I(new_n28102_), .ZN(new_n28132_));
  NOR2_X1    g25696(.A1(new_n28132_), .A2(new_n12841_), .ZN(new_n28133_));
  AOI21_X1   g25697(.A1(new_n12841_), .A2(new_n8780_), .B(new_n28133_), .ZN(new_n28134_));
  INV_X1     g25698(.I(new_n28134_), .ZN(new_n28135_));
  INV_X1     g25699(.I(new_n8761_), .ZN(new_n28136_));
  NOR2_X1    g25700(.A1(new_n8525_), .A2(pi1155), .ZN(new_n28137_));
  INV_X1     g25701(.I(new_n28137_), .ZN(new_n28138_));
  NOR2_X1    g25702(.A1(new_n28138_), .A2(new_n28136_), .ZN(new_n28139_));
  AOI21_X1   g25703(.A1(new_n28139_), .A2(pi1153), .B(pi1154), .ZN(new_n28140_));
  OAI21_X1   g25704(.A1(new_n28135_), .A2(new_n12770_), .B(new_n28140_), .ZN(new_n28141_));
  OAI21_X1   g25705(.A1(new_n28131_), .A2(new_n12785_), .B(new_n28141_), .ZN(new_n28142_));
  NAND2_X1   g25706(.A1(new_n28142_), .A2(new_n2628_), .ZN(new_n28143_));
  AOI21_X1   g25707(.A1(new_n28143_), .A2(new_n28122_), .B(new_n8521_), .ZN(new_n28144_));
  NOR2_X1    g25708(.A1(new_n12770_), .A2(pi0199), .ZN(new_n28145_));
  INV_X1     g25709(.I(new_n28145_), .ZN(new_n28146_));
  NOR2_X1    g25710(.A1(new_n28132_), .A2(new_n28146_), .ZN(new_n28147_));
  NOR2_X1    g25711(.A1(new_n28147_), .A2(new_n28087_), .ZN(new_n28148_));
  NAND2_X1   g25712(.A1(new_n12785_), .A2(new_n12742_), .ZN(new_n28149_));
  OAI21_X1   g25713(.A1(new_n28148_), .A2(new_n28149_), .B(new_n8521_), .ZN(new_n28150_));
  NOR2_X1    g25714(.A1(new_n28123_), .A2(pi0299), .ZN(new_n28151_));
  NOR2_X1    g25715(.A1(new_n28151_), .A2(pi1155), .ZN(new_n28152_));
  INV_X1     g25716(.I(new_n28124_), .ZN(new_n28153_));
  NOR2_X1    g25717(.A1(new_n28153_), .A2(pi0299), .ZN(new_n28154_));
  NOR2_X1    g25718(.A1(new_n28154_), .A2(new_n12770_), .ZN(new_n28155_));
  NOR2_X1    g25719(.A1(new_n28155_), .A2(new_n28152_), .ZN(new_n28156_));
  NOR2_X1    g25720(.A1(new_n28156_), .A2(new_n12785_), .ZN(new_n28157_));
  NOR2_X1    g25721(.A1(new_n28104_), .A2(new_n28129_), .ZN(new_n28158_));
  NOR2_X1    g25722(.A1(new_n28158_), .A2(new_n12742_), .ZN(new_n28159_));
  NOR2_X1    g25723(.A1(new_n28157_), .A2(new_n28159_), .ZN(new_n28160_));
  INV_X1     g25724(.I(new_n28160_), .ZN(new_n28161_));
  AOI21_X1   g25725(.A1(new_n28161_), .A2(new_n28122_), .B(new_n28150_), .ZN(new_n28162_));
  NOR3_X1    g25726(.A1(new_n28144_), .A2(new_n28162_), .A3(new_n8522_), .ZN(new_n28163_));
  NOR4_X1    g25727(.A1(new_n28163_), .A2(new_n28121_), .A3(new_n8515_), .A4(new_n28095_), .ZN(new_n28164_));
  INV_X1     g25728(.I(new_n28095_), .ZN(new_n28165_));
  NOR2_X1    g25729(.A1(new_n28136_), .A2(new_n28127_), .ZN(new_n28166_));
  INV_X1     g25730(.I(new_n28166_), .ZN(new_n28167_));
  NOR2_X1    g25731(.A1(pi0199), .A2(pi1155), .ZN(new_n28168_));
  NOR3_X1    g25732(.A1(new_n28167_), .A2(pi1154), .A3(new_n28168_), .ZN(new_n28169_));
  NOR2_X1    g25733(.A1(new_n8691_), .A2(pi1153), .ZN(new_n28170_));
  NOR2_X1    g25734(.A1(new_n28110_), .A2(new_n9183_), .ZN(new_n28171_));
  AOI21_X1   g25735(.A1(new_n28153_), .A2(pi1154), .B(new_n28171_), .ZN(new_n28172_));
  NOR2_X1    g25736(.A1(new_n28172_), .A2(new_n28170_), .ZN(new_n28173_));
  NOR2_X1    g25737(.A1(new_n8525_), .A2(new_n8531_), .ZN(new_n28174_));
  NOR2_X1    g25738(.A1(new_n28174_), .A2(pi0299), .ZN(new_n28175_));
  NOR2_X1    g25739(.A1(new_n28175_), .A2(new_n12841_), .ZN(new_n28176_));
  NOR2_X1    g25740(.A1(new_n28176_), .A2(new_n12785_), .ZN(new_n28177_));
  AOI21_X1   g25741(.A1(new_n28173_), .A2(new_n28177_), .B(new_n28169_), .ZN(new_n28178_));
  INV_X1     g25742(.I(new_n28178_), .ZN(new_n28179_));
  NOR2_X1    g25743(.A1(new_n28179_), .A2(new_n8521_), .ZN(new_n28180_));
  NOR2_X1    g25744(.A1(new_n8531_), .A2(pi1155), .ZN(new_n28181_));
  NOR2_X1    g25745(.A1(new_n9183_), .A2(new_n28181_), .ZN(new_n28182_));
  NAND2_X1   g25746(.A1(new_n28182_), .A2(pi1156), .ZN(new_n28183_));
  INV_X1     g25747(.I(new_n28183_), .ZN(new_n28184_));
  NOR2_X1    g25748(.A1(new_n28147_), .A2(pi1154), .ZN(new_n28185_));
  NOR2_X1    g25749(.A1(new_n28145_), .A2(new_n8531_), .ZN(new_n28186_));
  NOR2_X1    g25750(.A1(new_n8781_), .A2(new_n28186_), .ZN(new_n28187_));
  INV_X1     g25751(.I(new_n28187_), .ZN(new_n28188_));
  NOR2_X1    g25752(.A1(new_n28185_), .A2(new_n28188_), .ZN(new_n28189_));
  NOR2_X1    g25753(.A1(new_n28189_), .A2(new_n28184_), .ZN(new_n28190_));
  INV_X1     g25754(.I(new_n28190_), .ZN(new_n28191_));
  NOR2_X1    g25755(.A1(new_n28191_), .A2(pi0207), .ZN(new_n28192_));
  OAI21_X1   g25756(.A1(new_n28180_), .A2(new_n28192_), .B(pi0208), .ZN(new_n28193_));
  NOR2_X1    g25757(.A1(new_n28111_), .A2(pi1156), .ZN(new_n28194_));
  INV_X1     g25758(.I(new_n28194_), .ZN(new_n28195_));
  NOR2_X1    g25759(.A1(pi0200), .A2(pi1155), .ZN(new_n28196_));
  NOR2_X1    g25760(.A1(new_n28126_), .A2(new_n28196_), .ZN(new_n28197_));
  NAND2_X1   g25761(.A1(new_n28197_), .A2(new_n28195_), .ZN(new_n28198_));
  NOR2_X1    g25762(.A1(new_n28198_), .A2(new_n8521_), .ZN(new_n28199_));
  NOR2_X1    g25763(.A1(new_n28199_), .A2(pi0208), .ZN(new_n28200_));
  NAND2_X1   g25764(.A1(new_n28175_), .A2(pi1156), .ZN(new_n28201_));
  NOR2_X1    g25765(.A1(new_n28136_), .A2(pi1156), .ZN(new_n28202_));
  INV_X1     g25766(.I(new_n28202_), .ZN(new_n28203_));
  AOI21_X1   g25767(.A1(new_n28201_), .A2(new_n28203_), .B(new_n28137_), .ZN(new_n28204_));
  INV_X1     g25768(.I(new_n28204_), .ZN(new_n28205_));
  NOR2_X1    g25769(.A1(new_n28205_), .A2(new_n8521_), .ZN(new_n28206_));
  OAI21_X1   g25770(.A1(new_n28206_), .A2(pi0208), .B(pi1157), .ZN(new_n28207_));
  OAI21_X1   g25771(.A1(new_n28200_), .A2(pi1157), .B(new_n28207_), .ZN(new_n28208_));
  AOI21_X1   g25772(.A1(new_n28193_), .A2(new_n28208_), .B(new_n28165_), .ZN(new_n28209_));
  NOR3_X1    g25773(.A1(new_n28164_), .A2(po1038), .A3(new_n28209_), .ZN(new_n28210_));
  NOR2_X1    g25774(.A1(new_n8509_), .A2(pi0214), .ZN(new_n28211_));
  NOR2_X1    g25775(.A1(new_n28020_), .A2(new_n28211_), .ZN(new_n28212_));
  INV_X1     g25776(.I(new_n28180_), .ZN(new_n28213_));
  NOR2_X1    g25777(.A1(new_n2628_), .A2(new_n2446_), .ZN(new_n28214_));
  INV_X1     g25778(.I(new_n28186_), .ZN(new_n28215_));
  NAND2_X1   g25779(.A1(new_n28215_), .A2(new_n2628_), .ZN(new_n28216_));
  NAND2_X1   g25780(.A1(new_n28216_), .A2(pi1154), .ZN(new_n28217_));
  OAI21_X1   g25781(.A1(new_n28217_), .A2(new_n28214_), .B(pi1156), .ZN(new_n28218_));
  NOR2_X1    g25782(.A1(new_n2628_), .A2(pi1144), .ZN(new_n28219_));
  NOR2_X1    g25783(.A1(new_n28158_), .A2(new_n28219_), .ZN(new_n28220_));
  NOR2_X1    g25784(.A1(new_n28220_), .A2(pi1154), .ZN(new_n28221_));
  NOR2_X1    g25785(.A1(new_n28218_), .A2(new_n28221_), .ZN(new_n28222_));
  INV_X1     g25786(.I(new_n28214_), .ZN(new_n28223_));
  NAND2_X1   g25787(.A1(new_n28185_), .A2(new_n28223_), .ZN(new_n28224_));
  INV_X1     g25788(.I(new_n28155_), .ZN(new_n28225_));
  NOR2_X1    g25789(.A1(new_n28139_), .A2(new_n12785_), .ZN(new_n28226_));
  INV_X1     g25790(.I(new_n28226_), .ZN(new_n28227_));
  AOI21_X1   g25791(.A1(new_n12770_), .A2(new_n28214_), .B(new_n28227_), .ZN(new_n28228_));
  OAI21_X1   g25792(.A1(new_n28225_), .A2(new_n28219_), .B(new_n28228_), .ZN(new_n28229_));
  AND3_X2    g25793(.A1(new_n28229_), .A2(new_n12742_), .A3(new_n28224_), .Z(new_n28230_));
  NOR2_X1    g25794(.A1(new_n28230_), .A2(new_n28222_), .ZN(new_n28231_));
  AOI21_X1   g25795(.A1(new_n28231_), .A2(new_n8521_), .B(new_n8522_), .ZN(new_n28232_));
  OAI21_X1   g25796(.A1(new_n28213_), .A2(new_n28214_), .B(new_n28232_), .ZN(new_n28233_));
  NOR2_X1    g25797(.A1(new_n28219_), .A2(pi1157), .ZN(new_n28234_));
  NOR2_X1    g25798(.A1(new_n12965_), .A2(pi0208), .ZN(new_n28235_));
  NOR2_X1    g25799(.A1(new_n28201_), .A2(new_n28137_), .ZN(new_n28236_));
  OAI21_X1   g25800(.A1(new_n28106_), .A2(new_n28236_), .B(new_n28026_), .ZN(new_n28237_));
  NAND2_X1   g25801(.A1(new_n28237_), .A2(new_n28223_), .ZN(new_n28238_));
  AOI22_X1   g25802(.A1(new_n28118_), .A2(new_n28234_), .B1(new_n28235_), .B2(new_n28238_), .ZN(new_n28239_));
  AOI21_X1   g25803(.A1(new_n28233_), .A2(new_n28239_), .B(pi0211), .ZN(new_n28240_));
  NOR2_X1    g25804(.A1(new_n2628_), .A2(new_n3605_), .ZN(new_n28241_));
  INV_X1     g25805(.I(new_n28241_), .ZN(new_n28242_));
  NOR2_X1    g25806(.A1(new_n2628_), .A2(pi1143), .ZN(new_n28243_));
  OAI21_X1   g25807(.A1(new_n28158_), .A2(new_n28243_), .B(new_n12785_), .ZN(new_n28244_));
  INV_X1     g25808(.I(new_n28217_), .ZN(new_n28245_));
  AOI21_X1   g25809(.A1(new_n28245_), .A2(new_n28242_), .B(new_n12742_), .ZN(new_n28246_));
  AOI21_X1   g25810(.A1(new_n12770_), .A2(new_n28241_), .B(new_n28227_), .ZN(new_n28247_));
  OAI21_X1   g25811(.A1(new_n28225_), .A2(new_n28243_), .B(new_n28247_), .ZN(new_n28248_));
  AOI21_X1   g25812(.A1(new_n28185_), .A2(new_n28242_), .B(pi1156), .ZN(new_n28249_));
  AOI22_X1   g25813(.A1(new_n28248_), .A2(new_n28249_), .B1(new_n28244_), .B2(new_n28246_), .ZN(new_n28250_));
  NAND2_X1   g25814(.A1(new_n28250_), .A2(new_n8521_), .ZN(new_n28251_));
  NAND2_X1   g25815(.A1(new_n28251_), .A2(pi0208), .ZN(new_n28252_));
  AOI21_X1   g25816(.A1(new_n28180_), .A2(new_n28242_), .B(new_n28252_), .ZN(new_n28253_));
  INV_X1     g25817(.I(new_n28118_), .ZN(new_n28254_));
  NOR3_X1    g25818(.A1(new_n28254_), .A2(pi1157), .A3(new_n28243_), .ZN(new_n28255_));
  INV_X1     g25819(.I(new_n28235_), .ZN(new_n28256_));
  AOI21_X1   g25820(.A1(new_n28237_), .A2(new_n28242_), .B(new_n28256_), .ZN(new_n28257_));
  NOR3_X1    g25821(.A1(new_n28253_), .A2(new_n28255_), .A3(new_n28257_), .ZN(new_n28258_));
  NOR2_X1    g25822(.A1(new_n28258_), .A2(new_n8510_), .ZN(new_n28259_));
  NOR3_X1    g25823(.A1(new_n28259_), .A2(new_n28212_), .A3(new_n28240_), .ZN(new_n28260_));
  NOR2_X1    g25824(.A1(new_n8811_), .A2(pi0211), .ZN(new_n28261_));
  INV_X1     g25825(.I(new_n28261_), .ZN(new_n28262_));
  NOR4_X1    g25826(.A1(new_n28253_), .A2(new_n28255_), .A3(new_n28257_), .A4(new_n28262_), .ZN(new_n28263_));
  OAI21_X1   g25827(.A1(new_n28260_), .A2(new_n28263_), .B(new_n8807_), .ZN(new_n28264_));
  AOI21_X1   g25828(.A1(new_n28264_), .A2(new_n28210_), .B(new_n26198_), .ZN(new_n28265_));
  AOI21_X1   g25829(.A1(new_n28265_), .A2(new_n28093_), .B(pi0209), .ZN(new_n28266_));
  NOR2_X1    g25830(.A1(pi0211), .A2(pi0214), .ZN(new_n28267_));
  INV_X1     g25831(.I(new_n28267_), .ZN(new_n28268_));
  NOR2_X1    g25832(.A1(new_n2628_), .A2(new_n12742_), .ZN(new_n28269_));
  NOR2_X1    g25833(.A1(new_n28189_), .A2(new_n28159_), .ZN(new_n28270_));
  NAND2_X1   g25834(.A1(new_n28270_), .A2(new_n8521_), .ZN(new_n28271_));
  OAI21_X1   g25835(.A1(new_n8521_), .A2(new_n28269_), .B(new_n28271_), .ZN(new_n28272_));
  OAI21_X1   g25836(.A1(new_n8521_), .A2(new_n28178_), .B(new_n28272_), .ZN(new_n28273_));
  OAI21_X1   g25837(.A1(new_n28206_), .A2(new_n28269_), .B(new_n28235_), .ZN(new_n28274_));
  OAI21_X1   g25838(.A1(new_n28254_), .A2(new_n28194_), .B(new_n28274_), .ZN(new_n28275_));
  AOI21_X1   g25839(.A1(new_n28273_), .A2(pi0208), .B(new_n28275_), .ZN(new_n28276_));
  NOR2_X1    g25840(.A1(new_n28276_), .A2(new_n28268_), .ZN(new_n28277_));
  NOR3_X1    g25841(.A1(new_n28191_), .A2(pi0207), .A3(new_n28051_), .ZN(new_n28278_));
  INV_X1     g25842(.I(new_n28142_), .ZN(new_n28279_));
  NOR2_X1    g25843(.A1(new_n28279_), .A2(new_n8521_), .ZN(new_n28280_));
  OR3_X2     g25844(.A1(new_n28280_), .A2(new_n8522_), .A3(new_n28278_), .Z(new_n28281_));
  INV_X1     g25845(.I(new_n28051_), .ZN(new_n28282_));
  AOI21_X1   g25846(.A1(new_n28282_), .A2(new_n8521_), .B(pi0208), .ZN(new_n28283_));
  INV_X1     g25847(.I(new_n28152_), .ZN(new_n28284_));
  NOR2_X1    g25848(.A1(new_n28102_), .A2(pi1156), .ZN(new_n28285_));
  INV_X1     g25849(.I(new_n28103_), .ZN(new_n28286_));
  NAND2_X1   g25850(.A1(new_n28286_), .A2(new_n9183_), .ZN(new_n28287_));
  AOI22_X1   g25851(.A1(new_n28284_), .A2(new_n28285_), .B1(new_n28287_), .B2(pi1156), .ZN(new_n28288_));
  NAND2_X1   g25852(.A1(new_n28288_), .A2(pi0207), .ZN(new_n28289_));
  NAND3_X1   g25853(.A1(new_n28289_), .A2(pi1157), .A3(new_n28283_), .ZN(new_n28290_));
  NOR2_X1    g25854(.A1(new_n8691_), .A2(pi1155), .ZN(new_n28291_));
  NAND2_X1   g25855(.A1(new_n28195_), .A2(new_n28153_), .ZN(new_n28292_));
  AOI21_X1   g25856(.A1(new_n28292_), .A2(new_n2628_), .B(new_n28291_), .ZN(new_n28293_));
  NAND2_X1   g25857(.A1(new_n28293_), .A2(new_n28283_), .ZN(new_n28294_));
  NAND3_X1   g25858(.A1(new_n28281_), .A2(new_n28290_), .A3(new_n28294_), .ZN(new_n28295_));
  NOR2_X1    g25859(.A1(new_n8510_), .A2(pi0214), .ZN(new_n28296_));
  NOR2_X1    g25860(.A1(new_n28000_), .A2(new_n28296_), .ZN(new_n28297_));
  INV_X1     g25861(.I(new_n28297_), .ZN(new_n28298_));
  AOI21_X1   g25862(.A1(new_n28295_), .A2(new_n28298_), .B(new_n28277_), .ZN(new_n28299_));
  NOR2_X1    g25863(.A1(new_n28157_), .A2(new_n28191_), .ZN(new_n28300_));
  NOR2_X1    g25864(.A1(new_n28300_), .A2(pi0207), .ZN(new_n28301_));
  INV_X1     g25865(.I(new_n28301_), .ZN(new_n28302_));
  NAND2_X1   g25866(.A1(new_n28130_), .A2(new_n2628_), .ZN(new_n28303_));
  AOI21_X1   g25867(.A1(new_n28303_), .A2(pi1154), .B(new_n28169_), .ZN(new_n28304_));
  NOR2_X1    g25868(.A1(new_n28304_), .A2(new_n8521_), .ZN(new_n28305_));
  INV_X1     g25869(.I(new_n28305_), .ZN(new_n28306_));
  AOI21_X1   g25870(.A1(new_n28306_), .A2(new_n28302_), .B(new_n8522_), .ZN(new_n28307_));
  OAI21_X1   g25871(.A1(new_n28199_), .A2(new_n28048_), .B(new_n8522_), .ZN(new_n28308_));
  INV_X1     g25872(.I(new_n28308_), .ZN(new_n28309_));
  NOR2_X1    g25873(.A1(new_n2628_), .A2(pi1154), .ZN(new_n28310_));
  NOR2_X1    g25874(.A1(new_n28310_), .A2(new_n12965_), .ZN(new_n28311_));
  AOI22_X1   g25875(.A1(new_n28309_), .A2(new_n12965_), .B1(new_n28108_), .B2(new_n28311_), .ZN(new_n28312_));
  INV_X1     g25876(.I(new_n28312_), .ZN(new_n28313_));
  OAI21_X1   g25877(.A1(new_n28307_), .A2(new_n28313_), .B(new_n8512_), .ZN(new_n28314_));
  AOI21_X1   g25878(.A1(new_n28299_), .A2(new_n28314_), .B(new_n8509_), .ZN(new_n28315_));
  NAND2_X1   g25879(.A1(new_n28193_), .A2(new_n28208_), .ZN(new_n28316_));
  AOI21_X1   g25880(.A1(new_n28316_), .A2(new_n8511_), .B(pi0212), .ZN(new_n28317_));
  INV_X1     g25881(.I(new_n28200_), .ZN(new_n28318_));
  AOI21_X1   g25882(.A1(new_n28193_), .A2(new_n28318_), .B(pi1157), .ZN(new_n28319_));
  INV_X1     g25883(.I(new_n28109_), .ZN(new_n28320_));
  INV_X1     g25884(.I(new_n28151_), .ZN(new_n28321_));
  AOI21_X1   g25885(.A1(pi1153), .A2(new_n28321_), .B(new_n28173_), .ZN(new_n28322_));
  INV_X1     g25886(.I(new_n28322_), .ZN(new_n28323_));
  NOR2_X1    g25887(.A1(new_n28323_), .A2(new_n28027_), .ZN(new_n28324_));
  NOR2_X1    g25888(.A1(new_n28113_), .A2(new_n12770_), .ZN(new_n28325_));
  INV_X1     g25889(.I(new_n28325_), .ZN(new_n28326_));
  NAND2_X1   g25890(.A1(new_n12770_), .A2(pi0299), .ZN(new_n28327_));
  NAND2_X1   g25891(.A1(new_n28326_), .A2(new_n28327_), .ZN(new_n28328_));
  NOR2_X1    g25892(.A1(new_n28161_), .A2(new_n28328_), .ZN(new_n28329_));
  INV_X1     g25893(.I(new_n28329_), .ZN(new_n28330_));
  NOR2_X1    g25894(.A1(new_n28330_), .A2(pi0207), .ZN(new_n28331_));
  NOR3_X1    g25895(.A1(new_n28331_), .A2(new_n8522_), .A3(new_n28324_), .ZN(new_n28332_));
  OAI21_X1   g25896(.A1(new_n28332_), .A2(new_n28320_), .B(new_n8510_), .ZN(new_n28333_));
  NOR2_X1    g25897(.A1(new_n28333_), .A2(new_n28319_), .ZN(new_n28334_));
  OAI21_X1   g25898(.A1(new_n28276_), .A2(new_n8510_), .B(pi0214), .ZN(new_n28335_));
  OAI21_X1   g25899(.A1(new_n28334_), .A2(new_n28335_), .B(new_n28317_), .ZN(new_n28336_));
  NAND2_X1   g25900(.A1(new_n28336_), .A2(new_n8807_), .ZN(new_n28337_));
  NOR2_X1    g25901(.A1(new_n2628_), .A2(pi1153), .ZN(new_n28338_));
  OR3_X2     g25902(.A1(new_n28119_), .A2(new_n28109_), .A3(new_n28338_), .Z(new_n28339_));
  NOR3_X1    g25903(.A1(new_n28329_), .A2(pi0207), .A3(new_n28338_), .ZN(new_n28340_));
  NOR2_X1    g25904(.A1(new_n28322_), .A2(new_n8521_), .ZN(new_n28341_));
  OAI21_X1   g25905(.A1(new_n28340_), .A2(new_n28341_), .B(pi0208), .ZN(new_n28342_));
  NAND3_X1   g25906(.A1(new_n28342_), .A2(new_n28339_), .A3(new_n28000_), .ZN(new_n28343_));
  OR3_X2     g25907(.A1(new_n28307_), .A2(new_n28268_), .A3(new_n28313_), .Z(new_n28344_));
  NAND3_X1   g25908(.A1(new_n28343_), .A2(new_n28344_), .A3(pi0212), .ZN(new_n28345_));
  OAI21_X1   g25909(.A1(new_n28295_), .A2(new_n28001_), .B(new_n28317_), .ZN(new_n28346_));
  AOI22_X1   g25910(.A1(new_n28345_), .A2(new_n28346_), .B1(pi0211), .B2(new_n28316_), .ZN(new_n28347_));
  OAI22_X1   g25911(.A1(new_n28337_), .A2(new_n28315_), .B1(new_n8807_), .B2(new_n28347_), .ZN(new_n28348_));
  OAI21_X1   g25912(.A1(new_n28348_), .A2(po1038), .B(new_n28025_), .ZN(new_n28349_));
  AOI21_X1   g25913(.A1(new_n28349_), .A2(new_n28266_), .B(new_n27999_), .ZN(new_n28350_));
  AOI22_X1   g25914(.A1(new_n28350_), .A2(new_n28092_), .B1(new_n27999_), .B2(pi0233), .ZN(po0390));
  NOR2_X1    g25915(.A1(new_n28003_), .A2(new_n8807_), .ZN(new_n28352_));
  INV_X1     g25916(.I(new_n28013_), .ZN(new_n28353_));
  INV_X1     g25917(.I(new_n28014_), .ZN(new_n28354_));
  AOI21_X1   g25918(.A1(new_n28354_), .A2(new_n28353_), .B(new_n8511_), .ZN(new_n28355_));
  INV_X1     g25919(.I(new_n28355_), .ZN(new_n28356_));
  NOR2_X1    g25920(.A1(new_n28356_), .A2(pi0212), .ZN(new_n28357_));
  NOR3_X1    g25921(.A1(new_n28357_), .A2(pi0219), .A3(new_n28016_), .ZN(new_n28358_));
  OR4_X2     g25922(.A1(new_n26198_), .A2(new_n28358_), .A3(new_n28060_), .A4(new_n28352_), .Z(new_n28359_));
  INV_X1     g25923(.I(pi0209), .ZN(new_n28360_));
  INV_X1     g25924(.I(new_n28094_), .ZN(new_n28361_));
  NOR2_X1    g25925(.A1(new_n8510_), .A2(pi1153), .ZN(new_n28362_));
  AOI21_X1   g25926(.A1(new_n8510_), .A2(new_n12785_), .B(new_n28362_), .ZN(new_n28363_));
  INV_X1     g25927(.I(new_n28363_), .ZN(new_n28364_));
  AOI21_X1   g25928(.A1(new_n28364_), .A2(new_n8811_), .B(new_n28361_), .ZN(new_n28365_));
  INV_X1     g25929(.I(new_n28365_), .ZN(new_n28366_));
  NOR2_X1    g25930(.A1(new_n28366_), .A2(new_n28006_), .ZN(new_n28367_));
  AOI21_X1   g25931(.A1(new_n28367_), .A2(po1038), .B(pi1152), .ZN(new_n28368_));
  INV_X1     g25932(.I(new_n28368_), .ZN(new_n28369_));
  NOR2_X1    g25933(.A1(new_n8522_), .A2(pi0207), .ZN(new_n28370_));
  NOR2_X1    g25934(.A1(new_n28041_), .A2(new_n28370_), .ZN(new_n28371_));
  INV_X1     g25935(.I(new_n28371_), .ZN(new_n28372_));
  INV_X1     g25936(.I(new_n9217_), .ZN(new_n28373_));
  NOR2_X1    g25937(.A1(new_n28373_), .A2(new_n12841_), .ZN(new_n28374_));
  NOR2_X1    g25938(.A1(new_n28374_), .A2(pi1154), .ZN(new_n28375_));
  AOI21_X1   g25939(.A1(pi0200), .A2(new_n12841_), .B(new_n9183_), .ZN(new_n28376_));
  INV_X1     g25940(.I(new_n28376_), .ZN(new_n28377_));
  AOI21_X1   g25941(.A1(pi1154), .A2(new_n28377_), .B(new_n28375_), .ZN(new_n28378_));
  NAND2_X1   g25942(.A1(new_n28378_), .A2(new_n28372_), .ZN(new_n28379_));
  NOR2_X1    g25943(.A1(new_n28027_), .A2(new_n8522_), .ZN(new_n28380_));
  NOR2_X1    g25944(.A1(new_n8780_), .A2(new_n12841_), .ZN(new_n28381_));
  NAND2_X1   g25945(.A1(new_n28380_), .A2(new_n28381_), .ZN(new_n28382_));
  NAND2_X1   g25946(.A1(new_n28379_), .A2(new_n28382_), .ZN(new_n28383_));
  INV_X1     g25947(.I(new_n28383_), .ZN(new_n28384_));
  NOR2_X1    g25948(.A1(new_n8514_), .A2(new_n28361_), .ZN(new_n28385_));
  INV_X1     g25949(.I(new_n28385_), .ZN(new_n28386_));
  AOI21_X1   g25950(.A1(new_n28384_), .A2(new_n28386_), .B(po1038), .ZN(new_n28387_));
  NOR2_X1    g25951(.A1(new_n8780_), .A2(pi1153), .ZN(new_n28388_));
  INV_X1     g25952(.I(new_n28388_), .ZN(new_n28389_));
  NOR2_X1    g25953(.A1(new_n9171_), .A2(new_n12841_), .ZN(new_n28390_));
  INV_X1     g25954(.I(new_n28390_), .ZN(new_n28391_));
  AOI21_X1   g25955(.A1(new_n28389_), .A2(new_n28391_), .B(new_n12785_), .ZN(new_n28392_));
  NOR2_X1    g25956(.A1(new_n28392_), .A2(new_n28374_), .ZN(new_n28393_));
  NAND2_X1   g25957(.A1(new_n28393_), .A2(new_n8521_), .ZN(new_n28394_));
  INV_X1     g25958(.I(new_n28310_), .ZN(new_n28395_));
  OAI21_X1   g25959(.A1(new_n8641_), .A2(new_n12841_), .B(new_n2628_), .ZN(new_n28396_));
  NAND2_X1   g25960(.A1(new_n28396_), .A2(new_n28395_), .ZN(new_n28397_));
  AOI21_X1   g25961(.A1(new_n28397_), .A2(pi0207), .B(new_n8522_), .ZN(new_n28398_));
  INV_X1     g25962(.I(new_n28048_), .ZN(new_n28399_));
  NOR3_X1    g25963(.A1(new_n28392_), .A2(new_n8521_), .A3(new_n28374_), .ZN(new_n28400_));
  AOI21_X1   g25964(.A1(new_n8521_), .A2(new_n28399_), .B(new_n28400_), .ZN(new_n28401_));
  AOI22_X1   g25965(.A1(new_n28401_), .A2(new_n8522_), .B1(new_n28394_), .B2(new_n28398_), .ZN(new_n28402_));
  NOR2_X1    g25966(.A1(new_n28402_), .A2(pi0211), .ZN(new_n28403_));
  NOR2_X1    g25967(.A1(new_n28381_), .A2(new_n8521_), .ZN(new_n28404_));
  NOR2_X1    g25968(.A1(new_n8761_), .A2(pi1153), .ZN(new_n28405_));
  NOR3_X1    g25969(.A1(new_n28405_), .A2(new_n12785_), .A3(new_n9171_), .ZN(new_n28406_));
  NOR3_X1    g25970(.A1(new_n28113_), .A2(new_n12841_), .A3(pi1154), .ZN(new_n28407_));
  NOR3_X1    g25971(.A1(new_n28407_), .A2(pi0207), .A3(new_n28406_), .ZN(new_n28408_));
  OAI21_X1   g25972(.A1(new_n28408_), .A2(new_n28404_), .B(pi0208), .ZN(new_n28409_));
  INV_X1     g25973(.I(new_n28409_), .ZN(new_n28410_));
  INV_X1     g25974(.I(new_n28046_), .ZN(new_n28411_));
  NOR2_X1    g25975(.A1(new_n28411_), .A2(pi0207), .ZN(new_n28412_));
  NOR2_X1    g25976(.A1(new_n28407_), .A2(new_n28406_), .ZN(new_n28413_));
  NOR2_X1    g25977(.A1(new_n28413_), .A2(new_n8521_), .ZN(new_n28414_));
  NOR3_X1    g25978(.A1(new_n28414_), .A2(pi0208), .A3(new_n28412_), .ZN(new_n28415_));
  NOR3_X1    g25979(.A1(new_n28415_), .A2(new_n28410_), .A3(new_n8510_), .ZN(new_n28416_));
  NOR3_X1    g25980(.A1(new_n28403_), .A2(new_n28212_), .A3(new_n28416_), .ZN(new_n28417_));
  NOR2_X1    g25981(.A1(new_n28415_), .A2(new_n28410_), .ZN(new_n28418_));
  NOR2_X1    g25982(.A1(new_n28418_), .A2(new_n28262_), .ZN(new_n28419_));
  OAI21_X1   g25983(.A1(new_n28417_), .A2(new_n28419_), .B(new_n8807_), .ZN(new_n28420_));
  AOI21_X1   g25984(.A1(new_n28420_), .A2(new_n28387_), .B(new_n28369_), .ZN(new_n28421_));
  INV_X1     g25985(.I(pi1152), .ZN(new_n28422_));
  NAND2_X1   g25986(.A1(new_n28267_), .A2(new_n12785_), .ZN(new_n28423_));
  NAND2_X1   g25987(.A1(new_n28298_), .A2(new_n12841_), .ZN(new_n28424_));
  NAND3_X1   g25988(.A1(new_n28424_), .A2(pi0212), .A3(new_n28423_), .ZN(new_n28425_));
  AOI21_X1   g25989(.A1(new_n28363_), .A2(new_n28020_), .B(pi0219), .ZN(new_n28426_));
  NAND2_X1   g25990(.A1(new_n28425_), .A2(new_n28426_), .ZN(new_n28427_));
  AOI21_X1   g25991(.A1(new_n28427_), .A2(new_n28059_), .B(new_n28422_), .ZN(new_n28428_));
  INV_X1     g25992(.I(new_n28428_), .ZN(new_n28429_));
  INV_X1     g25993(.I(new_n28056_), .ZN(new_n28430_));
  INV_X1     g25994(.I(new_n28375_), .ZN(new_n28431_));
  NAND2_X1   g25995(.A1(new_n8525_), .A2(pi1153), .ZN(new_n28432_));
  NAND3_X1   g25996(.A1(new_n28102_), .A2(new_n28432_), .A3(pi1154), .ZN(new_n28433_));
  AOI21_X1   g25997(.A1(new_n28431_), .A2(new_n28433_), .B(new_n28321_), .ZN(new_n28434_));
  INV_X1     g25998(.I(new_n28434_), .ZN(new_n28435_));
  NAND2_X1   g25999(.A1(new_n28435_), .A2(new_n8521_), .ZN(new_n28436_));
  NOR2_X1    g26000(.A1(pi0200), .A2(pi1153), .ZN(new_n28437_));
  NOR2_X1    g26001(.A1(new_n28437_), .A2(pi0199), .ZN(new_n28438_));
  NOR2_X1    g26002(.A1(new_n28438_), .A2(pi0299), .ZN(new_n28439_));
  INV_X1     g26003(.I(new_n28439_), .ZN(new_n28440_));
  NOR2_X1    g26004(.A1(new_n28440_), .A2(new_n28123_), .ZN(new_n28441_));
  NOR2_X1    g26005(.A1(new_n28441_), .A2(new_n8521_), .ZN(new_n28442_));
  INV_X1     g26006(.I(new_n28442_), .ZN(new_n28443_));
  AOI21_X1   g26007(.A1(new_n28436_), .A2(new_n28443_), .B(new_n8522_), .ZN(new_n28444_));
  INV_X1     g26008(.I(new_n28444_), .ZN(new_n28445_));
  NAND2_X1   g26009(.A1(new_n28435_), .A2(new_n28097_), .ZN(new_n28446_));
  NAND2_X1   g26010(.A1(new_n28445_), .A2(new_n28446_), .ZN(new_n28447_));
  INV_X1     g26011(.I(new_n28175_), .ZN(new_n28448_));
  NOR2_X1    g26012(.A1(new_n8641_), .A2(pi1153), .ZN(new_n28449_));
  NOR2_X1    g26013(.A1(new_n28448_), .A2(new_n28449_), .ZN(new_n28450_));
  NOR2_X1    g26014(.A1(pi0199), .A2(pi1153), .ZN(new_n28451_));
  NOR2_X1    g26015(.A1(new_n28126_), .A2(new_n28451_), .ZN(new_n28452_));
  OAI21_X1   g26016(.A1(pi1153), .A2(new_n10288_), .B(new_n28177_), .ZN(new_n28453_));
  INV_X1     g26017(.I(new_n28453_), .ZN(new_n28454_));
  NOR2_X1    g26018(.A1(new_n28454_), .A2(new_n28452_), .ZN(new_n28455_));
  INV_X1     g26019(.I(new_n28455_), .ZN(new_n28456_));
  AOI22_X1   g26020(.A1(new_n28456_), .A2(new_n28372_), .B1(new_n8523_), .B2(new_n28450_), .ZN(new_n28457_));
  NOR2_X1    g26021(.A1(new_n28457_), .A2(new_n8510_), .ZN(new_n28458_));
  AOI21_X1   g26022(.A1(new_n28447_), .A2(new_n8510_), .B(new_n28458_), .ZN(new_n28459_));
  INV_X1     g26023(.I(new_n28457_), .ZN(new_n28460_));
  NOR2_X1    g26024(.A1(new_n28460_), .A2(new_n28430_), .ZN(new_n28461_));
  AOI21_X1   g26025(.A1(new_n28459_), .A2(new_n28430_), .B(new_n28461_), .ZN(new_n28462_));
  OAI21_X1   g26026(.A1(new_n28462_), .A2(new_n8807_), .B(new_n6643_), .ZN(new_n28463_));
  INV_X1     g26027(.I(new_n28463_), .ZN(new_n28464_));
  NOR2_X1    g26028(.A1(new_n28132_), .A2(new_n8525_), .ZN(new_n28465_));
  NOR2_X1    g26029(.A1(new_n28465_), .A2(new_n8521_), .ZN(new_n28466_));
  INV_X1     g26030(.I(new_n28466_), .ZN(new_n28467_));
  NOR2_X1    g26031(.A1(new_n28154_), .A2(new_n28405_), .ZN(new_n28468_));
  NOR2_X1    g26032(.A1(new_n28468_), .A2(new_n28406_), .ZN(new_n28469_));
  OAI22_X1   g26033(.A1(new_n28469_), .A2(pi0207), .B1(new_n28388_), .B2(new_n28467_), .ZN(new_n28470_));
  NOR2_X1    g26034(.A1(new_n28470_), .A2(new_n8522_), .ZN(new_n28471_));
  NOR2_X1    g26035(.A1(new_n28046_), .A2(pi0207), .ZN(new_n28472_));
  INV_X1     g26036(.I(new_n28472_), .ZN(new_n28473_));
  NAND2_X1   g26037(.A1(new_n28469_), .A2(pi0207), .ZN(new_n28474_));
  AOI21_X1   g26038(.A1(new_n28474_), .A2(new_n28473_), .B(pi0208), .ZN(new_n28475_));
  NOR2_X1    g26039(.A1(new_n28471_), .A2(new_n28475_), .ZN(new_n28476_));
  NOR2_X1    g26040(.A1(new_n8780_), .A2(new_n12785_), .ZN(new_n28477_));
  NOR2_X1    g26041(.A1(new_n28454_), .A2(new_n28477_), .ZN(new_n28478_));
  INV_X1     g26042(.I(new_n28478_), .ZN(new_n28479_));
  OAI21_X1   g26043(.A1(new_n28479_), .A2(new_n28452_), .B(new_n8521_), .ZN(new_n28480_));
  OAI21_X1   g26044(.A1(new_n28310_), .A2(new_n28443_), .B(new_n28480_), .ZN(new_n28481_));
  NOR2_X1    g26045(.A1(new_n28481_), .A2(new_n8522_), .ZN(new_n28482_));
  AOI21_X1   g26046(.A1(new_n28456_), .A2(pi0207), .B(pi0208), .ZN(new_n28483_));
  INV_X1     g26047(.I(new_n28483_), .ZN(new_n28484_));
  NOR2_X1    g26048(.A1(new_n28484_), .A2(new_n28048_), .ZN(new_n28485_));
  NOR2_X1    g26049(.A1(new_n28482_), .A2(new_n28485_), .ZN(new_n28486_));
  INV_X1     g26050(.I(new_n28486_), .ZN(new_n28487_));
  NAND2_X1   g26051(.A1(new_n28487_), .A2(new_n8510_), .ZN(new_n28488_));
  OAI21_X1   g26052(.A1(new_n8510_), .A2(new_n28476_), .B(new_n28488_), .ZN(new_n28489_));
  NOR2_X1    g26053(.A1(new_n28457_), .A2(pi0214), .ZN(new_n28490_));
  INV_X1     g26054(.I(new_n28490_), .ZN(new_n28491_));
  OAI21_X1   g26055(.A1(new_n28489_), .A2(new_n8511_), .B(new_n28491_), .ZN(new_n28492_));
  NAND2_X1   g26056(.A1(new_n28492_), .A2(new_n8509_), .ZN(new_n28493_));
  NOR2_X1    g26057(.A1(new_n28447_), .A2(new_n8510_), .ZN(new_n28494_));
  NOR2_X1    g26058(.A1(new_n28476_), .A2(pi0211), .ZN(new_n28495_));
  OAI21_X1   g26059(.A1(new_n28494_), .A2(new_n28495_), .B(pi0214), .ZN(new_n28496_));
  NAND2_X1   g26060(.A1(new_n28489_), .A2(new_n8511_), .ZN(new_n28497_));
  NAND3_X1   g26061(.A1(new_n28497_), .A2(pi0212), .A3(new_n28496_), .ZN(new_n28498_));
  NAND3_X1   g26062(.A1(new_n28493_), .A2(new_n28498_), .A3(new_n8807_), .ZN(new_n28499_));
  AOI21_X1   g26063(.A1(new_n28499_), .A2(new_n28464_), .B(new_n28429_), .ZN(new_n28500_));
  NOR2_X1    g26064(.A1(new_n28500_), .A2(new_n28421_), .ZN(new_n28501_));
  NOR2_X1    g26065(.A1(new_n28501_), .A2(pi0213), .ZN(new_n28502_));
  INV_X1     g26066(.I(new_n28057_), .ZN(new_n28503_));
  NOR2_X1    g26067(.A1(new_n28486_), .A2(new_n28503_), .ZN(new_n28504_));
  NOR2_X1    g26068(.A1(new_n28460_), .A2(new_n28057_), .ZN(new_n28505_));
  NOR3_X1    g26069(.A1(new_n28504_), .A2(new_n8807_), .A3(new_n28505_), .ZN(new_n28506_));
  NOR2_X1    g26070(.A1(new_n8641_), .A2(pi1154), .ZN(new_n28507_));
  NAND2_X1   g26071(.A1(new_n28507_), .A2(new_n28096_), .ZN(new_n28508_));
  INV_X1     g26072(.I(new_n28283_), .ZN(new_n28509_));
  OAI21_X1   g26073(.A1(new_n28509_), .A2(new_n28434_), .B(new_n28445_), .ZN(new_n28510_));
  NAND3_X1   g26074(.A1(new_n28510_), .A2(new_n28327_), .A3(new_n28508_), .ZN(new_n28511_));
  NAND2_X1   g26075(.A1(new_n28511_), .A2(new_n8510_), .ZN(new_n28512_));
  NAND2_X1   g26076(.A1(new_n28487_), .A2(pi0211), .ZN(new_n28513_));
  AOI21_X1   g26077(.A1(new_n28513_), .A2(new_n28512_), .B(new_n8811_), .ZN(new_n28514_));
  OAI21_X1   g26078(.A1(new_n28484_), .A2(new_n28269_), .B(new_n8510_), .ZN(new_n28515_));
  INV_X1     g26079(.I(new_n28269_), .ZN(new_n28516_));
  NAND2_X1   g26080(.A1(new_n28455_), .A2(new_n28516_), .ZN(new_n28517_));
  NOR2_X1    g26081(.A1(new_n2628_), .A2(pi1156), .ZN(new_n28518_));
  OAI21_X1   g26082(.A1(new_n28443_), .A2(new_n28518_), .B(pi0208), .ZN(new_n28519_));
  AOI21_X1   g26083(.A1(new_n28517_), .A2(new_n8521_), .B(new_n28519_), .ZN(new_n28520_));
  OAI22_X1   g26084(.A1(new_n28511_), .A2(new_n8510_), .B1(new_n28515_), .B2(new_n28520_), .ZN(new_n28521_));
  NOR2_X1    g26085(.A1(new_n28521_), .A2(new_n28066_), .ZN(new_n28522_));
  NOR4_X1    g26086(.A1(new_n28514_), .A2(new_n28522_), .A3(pi0219), .A4(new_n28461_), .ZN(new_n28523_));
  OAI21_X1   g26087(.A1(new_n28523_), .A2(new_n28506_), .B(pi1152), .ZN(new_n28524_));
  NOR2_X1    g26088(.A1(new_n28056_), .A2(new_n8807_), .ZN(new_n28525_));
  NOR2_X1    g26089(.A1(new_n28384_), .A2(new_n8510_), .ZN(new_n28526_));
  OAI21_X1   g26090(.A1(new_n28526_), .A2(new_n28403_), .B(new_n28525_), .ZN(new_n28527_));
  NAND2_X1   g26091(.A1(new_n28383_), .A2(new_n28056_), .ZN(new_n28528_));
  NAND2_X1   g26092(.A1(new_n28527_), .A2(new_n28528_), .ZN(new_n28529_));
  NOR2_X1    g26093(.A1(new_n28383_), .A2(pi0211), .ZN(new_n28530_));
  AOI21_X1   g26094(.A1(new_n28530_), .A2(new_n28516_), .B(new_n28066_), .ZN(new_n28531_));
  INV_X1     g26095(.I(new_n28291_), .ZN(new_n28532_));
  INV_X1     g26096(.I(new_n28374_), .ZN(new_n28533_));
  NAND2_X1   g26097(.A1(new_n28533_), .A2(new_n28282_), .ZN(new_n28534_));
  AOI22_X1   g26098(.A1(new_n28534_), .A2(new_n12785_), .B1(new_n28532_), .B2(new_n28392_), .ZN(new_n28535_));
  NAND2_X1   g26099(.A1(new_n28535_), .A2(pi0207), .ZN(new_n28536_));
  NAND2_X1   g26100(.A1(new_n28536_), .A2(new_n28283_), .ZN(new_n28537_));
  AOI21_X1   g26101(.A1(new_n28396_), .A2(new_n28327_), .B(new_n8521_), .ZN(new_n28538_));
  NOR2_X1    g26102(.A1(new_n28538_), .A2(new_n8522_), .ZN(new_n28539_));
  NAND2_X1   g26103(.A1(new_n28535_), .A2(new_n8521_), .ZN(new_n28540_));
  NAND2_X1   g26104(.A1(new_n28540_), .A2(new_n28539_), .ZN(new_n28541_));
  NAND2_X1   g26105(.A1(new_n28537_), .A2(new_n28541_), .ZN(new_n28542_));
  OAI21_X1   g26106(.A1(new_n8510_), .A2(new_n28542_), .B(new_n28531_), .ZN(new_n28543_));
  AOI21_X1   g26107(.A1(new_n28402_), .A2(pi0211), .B(new_n8811_), .ZN(new_n28544_));
  OAI21_X1   g26108(.A1(new_n28542_), .A2(pi0211), .B(new_n28544_), .ZN(new_n28545_));
  AOI21_X1   g26109(.A1(new_n28543_), .A2(new_n28545_), .B(pi0219), .ZN(new_n28546_));
  OAI21_X1   g26110(.A1(new_n28546_), .A2(new_n28529_), .B(new_n28422_), .ZN(new_n28547_));
  NAND2_X1   g26111(.A1(new_n28524_), .A2(new_n28547_), .ZN(new_n28548_));
  AOI21_X1   g26112(.A1(new_n28548_), .A2(new_n6643_), .B(new_n26198_), .ZN(new_n28549_));
  OAI21_X1   g26113(.A1(new_n28502_), .A2(new_n28549_), .B(new_n28360_), .ZN(new_n28550_));
  NOR2_X1    g26114(.A1(new_n28171_), .A2(pi1154), .ZN(new_n28551_));
  NOR2_X1    g26115(.A1(new_n8641_), .A2(pi1155), .ZN(new_n28552_));
  NOR3_X1    g26116(.A1(new_n28551_), .A2(new_n28448_), .A3(new_n28552_), .ZN(new_n28553_));
  AOI22_X1   g26117(.A1(new_n28191_), .A2(new_n28372_), .B1(new_n8523_), .B2(new_n28553_), .ZN(new_n28554_));
  INV_X1     g26118(.I(new_n28554_), .ZN(new_n28555_));
  AOI21_X1   g26119(.A1(new_n28555_), .A2(new_n28503_), .B(new_n8807_), .ZN(new_n28556_));
  INV_X1     g26120(.I(new_n28331_), .ZN(new_n28557_));
  NAND2_X1   g26121(.A1(new_n28329_), .A2(pi0207), .ZN(new_n28558_));
  NOR2_X1    g26122(.A1(new_n28552_), .A2(new_n28174_), .ZN(new_n28559_));
  OAI22_X1   g26123(.A1(new_n28559_), .A2(pi0299), .B1(pi1154), .B2(new_n28171_), .ZN(new_n28560_));
  AOI21_X1   g26124(.A1(new_n28560_), .A2(new_n28026_), .B(new_n8522_), .ZN(new_n28561_));
  AOI22_X1   g26125(.A1(new_n28557_), .A2(new_n28561_), .B1(new_n28097_), .B2(new_n28558_), .ZN(new_n28562_));
  OAI21_X1   g26126(.A1(new_n28562_), .A2(new_n28503_), .B(new_n28556_), .ZN(new_n28563_));
  NOR2_X1    g26127(.A1(new_n28562_), .A2(new_n28338_), .ZN(new_n28564_));
  NOR2_X1    g26128(.A1(new_n28300_), .A2(new_n8521_), .ZN(new_n28565_));
  INV_X1     g26129(.I(new_n28565_), .ZN(new_n28566_));
  NOR2_X1    g26130(.A1(new_n28399_), .A2(pi0207), .ZN(new_n28567_));
  INV_X1     g26131(.I(new_n28567_), .ZN(new_n28568_));
  AOI21_X1   g26132(.A1(new_n28566_), .A2(new_n28568_), .B(pi0208), .ZN(new_n28569_));
  OR2_X2     g26133(.A1(new_n28560_), .A2(new_n8521_), .Z(new_n28570_));
  AOI21_X1   g26134(.A1(new_n28302_), .A2(new_n28570_), .B(new_n8522_), .ZN(new_n28571_));
  NOR2_X1    g26135(.A1(new_n28569_), .A2(new_n28571_), .ZN(new_n28572_));
  NAND2_X1   g26136(.A1(new_n28572_), .A2(new_n8510_), .ZN(new_n28573_));
  OAI21_X1   g26137(.A1(new_n28564_), .A2(new_n8510_), .B(new_n28573_), .ZN(new_n28574_));
  NOR2_X1    g26138(.A1(new_n28554_), .A2(pi0214), .ZN(new_n28575_));
  INV_X1     g26139(.I(new_n28575_), .ZN(new_n28576_));
  OAI21_X1   g26140(.A1(new_n28574_), .A2(new_n8511_), .B(new_n28576_), .ZN(new_n28577_));
  AOI21_X1   g26141(.A1(new_n28577_), .A2(new_n8509_), .B(pi0219), .ZN(new_n28578_));
  NOR2_X1    g26142(.A1(new_n28574_), .A2(pi0214), .ZN(new_n28579_));
  INV_X1     g26143(.I(new_n28338_), .ZN(new_n28580_));
  NOR2_X1    g26144(.A1(new_n28580_), .A2(pi0211), .ZN(new_n28581_));
  NOR3_X1    g26145(.A1(new_n28562_), .A2(new_n8511_), .A3(new_n28581_), .ZN(new_n28582_));
  OAI21_X1   g26146(.A1(new_n28579_), .A2(new_n28582_), .B(pi0212), .ZN(new_n28583_));
  AOI21_X1   g26147(.A1(new_n28578_), .A2(new_n28583_), .B(po1038), .ZN(new_n28584_));
  AOI21_X1   g26148(.A1(new_n28584_), .A2(new_n28563_), .B(new_n28429_), .ZN(new_n28585_));
  OAI21_X1   g26149(.A1(new_n28555_), .A2(new_n8807_), .B(new_n6643_), .ZN(new_n28586_));
  NAND2_X1   g26150(.A1(new_n28555_), .A2(pi0211), .ZN(new_n28587_));
  NAND2_X1   g26151(.A1(new_n28564_), .A2(new_n8510_), .ZN(new_n28588_));
  AOI21_X1   g26152(.A1(new_n28588_), .A2(new_n28587_), .B(new_n8511_), .ZN(new_n28589_));
  OAI21_X1   g26153(.A1(new_n28579_), .A2(new_n28589_), .B(pi0212), .ZN(new_n28590_));
  AOI21_X1   g26154(.A1(new_n28578_), .A2(new_n28590_), .B(new_n28586_), .ZN(new_n28591_));
  OAI21_X1   g26155(.A1(new_n28591_), .A2(new_n28369_), .B(new_n26198_), .ZN(new_n28592_));
  INV_X1     g26156(.I(new_n28572_), .ZN(new_n28593_));
  NOR2_X1    g26157(.A1(new_n28593_), .A2(new_n8510_), .ZN(new_n28594_));
  OAI21_X1   g26158(.A1(new_n28191_), .A2(new_n28051_), .B(new_n28283_), .ZN(new_n28595_));
  OR2_X2     g26159(.A1(new_n28553_), .A2(new_n28051_), .Z(new_n28596_));
  OAI21_X1   g26160(.A1(new_n28596_), .A2(new_n8521_), .B(pi0208), .ZN(new_n28597_));
  OAI21_X1   g26161(.A1(new_n28278_), .A2(new_n28597_), .B(new_n28595_), .ZN(new_n28598_));
  NOR2_X1    g26162(.A1(new_n28598_), .A2(pi0211), .ZN(new_n28599_));
  OAI21_X1   g26163(.A1(new_n28594_), .A2(new_n28599_), .B(pi0214), .ZN(new_n28600_));
  NAND2_X1   g26164(.A1(new_n28553_), .A2(pi0207), .ZN(new_n28601_));
  AOI21_X1   g26165(.A1(new_n28272_), .A2(new_n28601_), .B(new_n8522_), .ZN(new_n28602_));
  NOR2_X1    g26166(.A1(new_n28270_), .A2(new_n8521_), .ZN(new_n28603_));
  INV_X1     g26167(.I(new_n28603_), .ZN(new_n28604_));
  NAND2_X1   g26168(.A1(new_n28604_), .A2(new_n28516_), .ZN(new_n28605_));
  AOI21_X1   g26169(.A1(new_n28605_), .A2(new_n8522_), .B(pi0211), .ZN(new_n28606_));
  INV_X1     g26170(.I(new_n28606_), .ZN(new_n28607_));
  OAI22_X1   g26171(.A1(new_n28607_), .A2(new_n28602_), .B1(new_n8510_), .B2(new_n28598_), .ZN(new_n28608_));
  AOI21_X1   g26172(.A1(new_n28608_), .A2(new_n8511_), .B(new_n8509_), .ZN(new_n28609_));
  NAND2_X1   g26173(.A1(new_n28600_), .A2(new_n28609_), .ZN(new_n28610_));
  OAI21_X1   g26174(.A1(new_n28608_), .A2(new_n8511_), .B(new_n28576_), .ZN(new_n28611_));
  AOI21_X1   g26175(.A1(new_n28611_), .A2(new_n8509_), .B(pi0219), .ZN(new_n28612_));
  NAND2_X1   g26176(.A1(new_n28610_), .A2(new_n28612_), .ZN(new_n28613_));
  NAND2_X1   g26177(.A1(new_n28593_), .A2(new_n28057_), .ZN(new_n28614_));
  AOI21_X1   g26178(.A1(new_n28614_), .A2(new_n28556_), .B(new_n26200_), .ZN(new_n28615_));
  AOI21_X1   g26179(.A1(new_n28613_), .A2(new_n28615_), .B(new_n28360_), .ZN(new_n28616_));
  OAI21_X1   g26180(.A1(new_n28592_), .A2(new_n28585_), .B(new_n28616_), .ZN(new_n28617_));
  AOI21_X1   g26181(.A1(new_n28550_), .A2(new_n28617_), .B(new_n27999_), .ZN(new_n28618_));
  AOI22_X1   g26182(.A1(new_n28618_), .A2(new_n28359_), .B1(new_n27999_), .B2(new_n3097_), .ZN(po0391));
  NOR2_X1    g26183(.A1(pi0207), .A2(pi0208), .ZN(new_n28620_));
  INV_X1     g26184(.I(new_n28620_), .ZN(new_n28621_));
  AOI21_X1   g26185(.A1(new_n28204_), .A2(new_n28621_), .B(new_n8523_), .ZN(new_n28622_));
  INV_X1     g26186(.I(new_n28147_), .ZN(new_n28623_));
  NOR2_X1    g26187(.A1(new_n28623_), .A2(pi1156), .ZN(new_n28624_));
  NOR3_X1    g26188(.A1(new_n28624_), .A2(new_n8524_), .A3(new_n28184_), .ZN(new_n28625_));
  OR3_X2     g26189(.A1(new_n28625_), .A2(new_n12965_), .A3(new_n28622_), .Z(new_n28626_));
  INV_X1     g26190(.I(new_n28198_), .ZN(new_n28627_));
  AOI21_X1   g26191(.A1(new_n28627_), .A2(new_n28621_), .B(new_n8523_), .ZN(new_n28628_));
  NOR3_X1    g26192(.A1(new_n28628_), .A2(pi1157), .A3(new_n28625_), .ZN(new_n28629_));
  INV_X1     g26193(.I(new_n28629_), .ZN(new_n28630_));
  NAND2_X1   g26194(.A1(new_n28630_), .A2(new_n28626_), .ZN(new_n28631_));
  AOI21_X1   g26195(.A1(new_n28631_), .A2(new_n28066_), .B(new_n8807_), .ZN(new_n28632_));
  OAI21_X1   g26196(.A1(new_n28631_), .A2(new_n8510_), .B(new_n28065_), .ZN(new_n28633_));
  NOR2_X1    g26197(.A1(new_n28254_), .A2(new_n28194_), .ZN(new_n28634_));
  OAI21_X1   g26198(.A1(new_n28624_), .A2(new_n28159_), .B(pi0207), .ZN(new_n28635_));
  NOR2_X1    g26199(.A1(new_n28115_), .A2(pi0207), .ZN(new_n28636_));
  INV_X1     g26200(.I(new_n28636_), .ZN(new_n28637_));
  AOI21_X1   g26201(.A1(new_n28637_), .A2(new_n28635_), .B(new_n8522_), .ZN(new_n28638_));
  OAI21_X1   g26202(.A1(new_n28634_), .A2(new_n28638_), .B(new_n12965_), .ZN(new_n28639_));
  INV_X1     g26203(.I(new_n28639_), .ZN(new_n28640_));
  AOI21_X1   g26204(.A1(new_n28107_), .A2(new_n8521_), .B(new_n8522_), .ZN(new_n28641_));
  INV_X1     g26205(.I(new_n28641_), .ZN(new_n28642_));
  NOR3_X1    g26206(.A1(new_n28328_), .A2(new_n8521_), .A3(new_n28159_), .ZN(new_n28643_));
  NOR2_X1    g26207(.A1(new_n28642_), .A2(new_n28643_), .ZN(new_n28644_));
  NOR2_X1    g26208(.A1(new_n28644_), .A2(new_n28108_), .ZN(new_n28645_));
  NOR2_X1    g26209(.A1(new_n28645_), .A2(new_n12965_), .ZN(new_n28646_));
  NOR2_X1    g26210(.A1(new_n2628_), .A2(pi1157), .ZN(new_n28647_));
  NOR3_X1    g26211(.A1(new_n28640_), .A2(new_n28646_), .A3(new_n28647_), .ZN(new_n28648_));
  NOR2_X1    g26212(.A1(new_n28648_), .A2(new_n28338_), .ZN(new_n28649_));
  NOR2_X1    g26213(.A1(new_n28649_), .A2(pi0211), .ZN(new_n28650_));
  OAI21_X1   g26214(.A1(new_n28650_), .A2(new_n28633_), .B(new_n28632_), .ZN(new_n28651_));
  OAI21_X1   g26215(.A1(new_n28648_), .A2(new_n28338_), .B(pi0211), .ZN(new_n28652_));
  INV_X1     g26216(.I(new_n28645_), .ZN(new_n28653_));
  NOR2_X1    g26217(.A1(new_n28110_), .A2(new_n8525_), .ZN(new_n28654_));
  NOR3_X1    g26218(.A1(new_n28654_), .A2(new_n28114_), .A3(new_n12742_), .ZN(new_n28655_));
  OAI22_X1   g26219(.A1(new_n28655_), .A2(new_n12785_), .B1(new_n28126_), .B2(new_n28196_), .ZN(new_n28656_));
  NAND2_X1   g26220(.A1(new_n28194_), .A2(new_n2628_), .ZN(new_n28657_));
  NAND3_X1   g26221(.A1(new_n28656_), .A2(new_n8521_), .A3(new_n28657_), .ZN(new_n28658_));
  INV_X1     g26222(.I(new_n28185_), .ZN(new_n28659_));
  NAND2_X1   g26223(.A1(new_n28659_), .A2(new_n28328_), .ZN(new_n28660_));
  AOI21_X1   g26224(.A1(new_n28660_), .A2(new_n28183_), .B(new_n8521_), .ZN(new_n28661_));
  INV_X1     g26225(.I(new_n28661_), .ZN(new_n28662_));
  AOI21_X1   g26226(.A1(new_n28662_), .A2(new_n28658_), .B(new_n8522_), .ZN(new_n28663_));
  OR2_X2     g26227(.A1(new_n28663_), .A2(new_n28309_), .Z(new_n28664_));
  AOI22_X1   g26228(.A1(new_n28664_), .A2(new_n12965_), .B1(new_n28311_), .B2(new_n28653_), .ZN(new_n28665_));
  NAND2_X1   g26229(.A1(new_n28665_), .A2(new_n8510_), .ZN(new_n28666_));
  AOI21_X1   g26230(.A1(new_n28652_), .A2(new_n28666_), .B(new_n8811_), .ZN(new_n28667_));
  NAND3_X1   g26231(.A1(new_n28630_), .A2(new_n28056_), .A3(new_n28626_), .ZN(new_n28668_));
  INV_X1     g26232(.I(new_n28212_), .ZN(new_n28669_));
  NOR2_X1    g26233(.A1(new_n8522_), .A2(new_n12965_), .ZN(new_n28670_));
  AOI21_X1   g26234(.A1(new_n28326_), .A2(new_n28183_), .B(new_n8521_), .ZN(new_n28671_));
  NOR2_X1    g26235(.A1(new_n28288_), .A2(pi0207), .ZN(new_n28672_));
  OAI21_X1   g26236(.A1(new_n28672_), .A2(new_n28671_), .B(new_n28670_), .ZN(new_n28673_));
  NAND2_X1   g26237(.A1(new_n28293_), .A2(new_n8521_), .ZN(new_n28674_));
  INV_X1     g26238(.I(new_n28674_), .ZN(new_n28675_));
  OAI21_X1   g26239(.A1(new_n28675_), .A2(new_n28671_), .B(pi0208), .ZN(new_n28676_));
  NAND2_X1   g26240(.A1(new_n28676_), .A2(new_n28294_), .ZN(new_n28677_));
  NAND2_X1   g26241(.A1(new_n28677_), .A2(new_n12965_), .ZN(new_n28678_));
  NAND3_X1   g26242(.A1(new_n28678_), .A2(new_n28290_), .A3(new_n28673_), .ZN(new_n28679_));
  NOR2_X1    g26243(.A1(new_n28679_), .A2(pi0211), .ZN(new_n28680_));
  AND2_X2    g26244(.A1(new_n28665_), .A2(pi0211), .Z(new_n28681_));
  OAI21_X1   g26245(.A1(new_n28681_), .A2(new_n28680_), .B(new_n28669_), .ZN(new_n28682_));
  NAND2_X1   g26246(.A1(new_n28682_), .A2(new_n28668_), .ZN(new_n28683_));
  OAI21_X1   g26247(.A1(new_n28683_), .A2(new_n28667_), .B(new_n8807_), .ZN(new_n28684_));
  NAND3_X1   g26248(.A1(new_n28684_), .A2(pi0209), .A3(new_n28651_), .ZN(new_n28685_));
  AOI21_X1   g26249(.A1(new_n28178_), .A2(new_n8524_), .B(new_n28620_), .ZN(new_n28686_));
  OAI21_X1   g26250(.A1(new_n8524_), .A2(new_n28378_), .B(new_n28686_), .ZN(new_n28687_));
  AOI21_X1   g26251(.A1(new_n28687_), .A2(pi0211), .B(new_n28066_), .ZN(new_n28688_));
  NOR2_X1    g26252(.A1(new_n28341_), .A2(new_n28412_), .ZN(new_n28689_));
  NOR2_X1    g26253(.A1(new_n28689_), .A2(pi0208), .ZN(new_n28690_));
  INV_X1     g26254(.I(new_n28414_), .ZN(new_n28691_));
  NAND2_X1   g26255(.A1(new_n28323_), .A2(new_n8521_), .ZN(new_n28692_));
  AOI21_X1   g26256(.A1(new_n28692_), .A2(new_n28691_), .B(new_n8522_), .ZN(new_n28693_));
  OR2_X2     g26257(.A1(new_n28690_), .A2(new_n28693_), .Z(new_n28694_));
  OAI21_X1   g26258(.A1(new_n28694_), .A2(pi0211), .B(new_n28688_), .ZN(new_n28695_));
  INV_X1     g26259(.I(new_n28687_), .ZN(new_n28696_));
  AOI21_X1   g26260(.A1(new_n28696_), .A2(new_n28066_), .B(new_n8807_), .ZN(new_n28697_));
  NAND2_X1   g26261(.A1(new_n28695_), .A2(new_n28697_), .ZN(new_n28698_));
  AOI21_X1   g26262(.A1(new_n28306_), .A2(new_n28568_), .B(pi0208), .ZN(new_n28699_));
  NAND2_X1   g26263(.A1(new_n28304_), .A2(new_n8521_), .ZN(new_n28700_));
  INV_X1     g26264(.I(new_n28700_), .ZN(new_n28701_));
  NOR3_X1    g26265(.A1(new_n28701_), .A2(new_n8522_), .A3(new_n28400_), .ZN(new_n28702_));
  OR3_X2     g26266(.A1(new_n28699_), .A2(new_n28702_), .A3(new_n8510_), .Z(new_n28703_));
  NOR2_X1    g26267(.A1(new_n28142_), .A2(new_n28509_), .ZN(new_n28704_));
  INV_X1     g26268(.I(new_n28704_), .ZN(new_n28705_));
  NOR2_X1    g26269(.A1(new_n28279_), .A2(pi0207), .ZN(new_n28706_));
  INV_X1     g26270(.I(new_n28706_), .ZN(new_n28707_));
  NAND3_X1   g26271(.A1(new_n28707_), .A2(pi0208), .A3(new_n28536_), .ZN(new_n28708_));
  NAND3_X1   g26272(.A1(new_n28708_), .A2(new_n8510_), .A3(new_n28705_), .ZN(new_n28709_));
  AOI21_X1   g26273(.A1(new_n28703_), .A2(new_n28709_), .B(new_n28066_), .ZN(new_n28710_));
  NOR2_X1    g26274(.A1(new_n28694_), .A2(new_n8510_), .ZN(new_n28711_));
  NOR3_X1    g26275(.A1(new_n28699_), .A2(new_n28702_), .A3(pi0211), .ZN(new_n28712_));
  NOR2_X1    g26276(.A1(new_n28711_), .A2(new_n28712_), .ZN(new_n28713_));
  OAI22_X1   g26277(.A1(new_n28713_), .A2(new_n8811_), .B1(new_n28430_), .B2(new_n28696_), .ZN(new_n28714_));
  OAI21_X1   g26278(.A1(new_n28714_), .A2(new_n28710_), .B(new_n8807_), .ZN(new_n28715_));
  NAND3_X1   g26279(.A1(new_n28715_), .A2(new_n28360_), .A3(new_n28698_), .ZN(new_n28716_));
  NAND2_X1   g26280(.A1(new_n28685_), .A2(new_n28716_), .ZN(new_n28717_));
  NOR2_X1    g26281(.A1(new_n28011_), .A2(new_n28010_), .ZN(new_n28718_));
  AOI21_X1   g26282(.A1(new_n28363_), .A2(new_n8809_), .B(pi0219), .ZN(new_n28719_));
  OAI21_X1   g26283(.A1(new_n28718_), .A2(new_n28212_), .B(new_n28719_), .ZN(new_n28720_));
  OAI21_X1   g26284(.A1(new_n8807_), .A2(new_n28669_), .B(new_n28720_), .ZN(new_n28721_));
  OAI21_X1   g26285(.A1(new_n12841_), .A2(pi0211), .B(pi0219), .ZN(new_n28722_));
  NAND2_X1   g26286(.A1(po1038), .A2(new_n28722_), .ZN(new_n28723_));
  OAI21_X1   g26287(.A1(new_n28721_), .A2(new_n28723_), .B(new_n26198_), .ZN(new_n28724_));
  AOI21_X1   g26288(.A1(new_n28717_), .A2(new_n6643_), .B(new_n28724_), .ZN(new_n28725_));
  INV_X1     g26289(.I(new_n28010_), .ZN(new_n28726_));
  OAI21_X1   g26290(.A1(new_n28212_), .A2(new_n28726_), .B(pi0219), .ZN(new_n28727_));
  OAI21_X1   g26291(.A1(pi0214), .A2(new_n28019_), .B(new_n28356_), .ZN(new_n28728_));
  AOI21_X1   g26292(.A1(new_n28728_), .A2(pi0212), .B(pi0219), .ZN(new_n28729_));
  OAI21_X1   g26293(.A1(new_n28019_), .A2(new_n28021_), .B(new_n28729_), .ZN(new_n28730_));
  NAND3_X1   g26294(.A1(new_n28730_), .A2(po1038), .A3(new_n28727_), .ZN(new_n28731_));
  INV_X1     g26295(.I(new_n28697_), .ZN(new_n28732_));
  AOI21_X1   g26296(.A1(new_n28709_), .A2(new_n28688_), .B(new_n28732_), .ZN(new_n28733_));
  NAND2_X1   g26297(.A1(new_n28687_), .A2(new_n12965_), .ZN(new_n28734_));
  NAND2_X1   g26298(.A1(new_n28322_), .A2(new_n28096_), .ZN(new_n28735_));
  INV_X1     g26299(.I(new_n28112_), .ZN(new_n28736_));
  OAI21_X1   g26300(.A1(new_n28736_), .A2(new_n12841_), .B(new_n2628_), .ZN(new_n28737_));
  AOI21_X1   g26301(.A1(new_n12785_), .A2(new_n28737_), .B(new_n28392_), .ZN(new_n28738_));
  NAND2_X1   g26302(.A1(new_n28738_), .A2(pi0207), .ZN(new_n28739_));
  NAND3_X1   g26303(.A1(new_n28735_), .A2(pi0208), .A3(new_n28739_), .ZN(new_n28740_));
  NOR2_X1    g26304(.A1(new_n28324_), .A2(new_n28098_), .ZN(new_n28741_));
  INV_X1     g26305(.I(new_n28741_), .ZN(new_n28742_));
  NAND3_X1   g26306(.A1(new_n28742_), .A2(pi1157), .A3(new_n28740_), .ZN(new_n28743_));
  AOI21_X1   g26307(.A1(new_n28743_), .A2(new_n28734_), .B(pi0211), .ZN(new_n28744_));
  NOR3_X1    g26308(.A1(new_n28696_), .A2(new_n8510_), .A3(new_n28269_), .ZN(new_n28745_));
  OAI21_X1   g26309(.A1(new_n28744_), .A2(new_n28745_), .B(new_n28669_), .ZN(new_n28746_));
  NAND3_X1   g26310(.A1(new_n28708_), .A2(pi0211), .A3(new_n28705_), .ZN(new_n28747_));
  NAND3_X1   g26311(.A1(new_n28687_), .A2(new_n8510_), .A3(new_n28516_), .ZN(new_n28748_));
  NAND2_X1   g26312(.A1(new_n28747_), .A2(new_n28748_), .ZN(new_n28749_));
  AOI22_X1   g26313(.A1(new_n28749_), .A2(new_n8809_), .B1(new_n28056_), .B2(new_n28687_), .ZN(new_n28750_));
  AOI21_X1   g26314(.A1(new_n28750_), .A2(new_n28746_), .B(pi0219), .ZN(new_n28751_));
  NOR3_X1    g26315(.A1(new_n28751_), .A2(pi0209), .A3(new_n28733_), .ZN(new_n28752_));
  NOR2_X1    g26316(.A1(new_n28679_), .A2(new_n8510_), .ZN(new_n28753_));
  INV_X1     g26317(.I(new_n28635_), .ZN(new_n28754_));
  AOI21_X1   g26318(.A1(new_n28138_), .A2(new_n28202_), .B(new_n28101_), .ZN(new_n28755_));
  NOR2_X1    g26319(.A1(new_n28755_), .A2(pi0207), .ZN(new_n28756_));
  OAI21_X1   g26320(.A1(new_n28754_), .A2(new_n28756_), .B(new_n28670_), .ZN(new_n28757_));
  NAND3_X1   g26321(.A1(new_n28639_), .A2(new_n28274_), .A3(new_n28757_), .ZN(new_n28758_));
  NOR2_X1    g26322(.A1(new_n28758_), .A2(pi0211), .ZN(new_n28759_));
  OAI21_X1   g26323(.A1(new_n28753_), .A2(new_n28759_), .B(new_n8809_), .ZN(new_n28760_));
  OAI21_X1   g26324(.A1(new_n28646_), .A2(new_n28629_), .B(new_n8510_), .ZN(new_n28761_));
  NAND2_X1   g26325(.A1(new_n28758_), .A2(pi0211), .ZN(new_n28762_));
  NAND3_X1   g26326(.A1(new_n28762_), .A2(new_n28669_), .A3(new_n28761_), .ZN(new_n28763_));
  NAND3_X1   g26327(.A1(new_n28760_), .A2(new_n28668_), .A3(new_n28763_), .ZN(new_n28764_));
  OAI21_X1   g26328(.A1(new_n28680_), .A2(new_n28633_), .B(new_n28632_), .ZN(new_n28765_));
  NAND2_X1   g26329(.A1(new_n28765_), .A2(pi0209), .ZN(new_n28766_));
  AOI21_X1   g26330(.A1(new_n28764_), .A2(new_n8807_), .B(new_n28766_), .ZN(new_n28767_));
  OAI21_X1   g26331(.A1(new_n28767_), .A2(new_n28752_), .B(new_n6643_), .ZN(new_n28768_));
  NAND3_X1   g26332(.A1(new_n28768_), .A2(pi0213), .A3(new_n28731_), .ZN(new_n28769_));
  NAND2_X1   g26333(.A1(new_n28769_), .A2(pi0230), .ZN(new_n28770_));
  OAI22_X1   g26334(.A1(new_n28770_), .A2(new_n28725_), .B1(pi0230), .B2(new_n3479_), .ZN(po0392));
  INV_X1     g26335(.I(new_n5302_), .ZN(new_n28772_));
  NAND2_X1   g26336(.A1(new_n27863_), .A2(new_n2702_), .ZN(new_n28773_));
  NAND3_X1   g26337(.A1(new_n28773_), .A2(new_n3458_), .A3(new_n5339_), .ZN(new_n28774_));
  AOI21_X1   g26338(.A1(new_n28774_), .A2(new_n28772_), .B(pi0075), .ZN(new_n28775_));
  OAI21_X1   g26339(.A1(new_n28775_), .A2(new_n6178_), .B(new_n3444_), .ZN(new_n28776_));
  NAND2_X1   g26340(.A1(new_n28776_), .A2(new_n10652_), .ZN(new_n28777_));
  AOI21_X1   g26341(.A1(new_n28777_), .A2(new_n2625_), .B(new_n5300_), .ZN(new_n28778_));
  AOI21_X1   g26342(.A1(new_n28778_), .A2(new_n2602_), .B(pi0056), .ZN(new_n28779_));
  OAI21_X1   g26343(.A1(new_n28779_), .A2(new_n5298_), .B(new_n3471_), .ZN(new_n28780_));
  AND3_X2    g26344(.A1(new_n28780_), .A2(new_n3291_), .A3(new_n5465_), .Z(po0393));
  NOR2_X1    g26345(.A1(new_n28068_), .A2(new_n8807_), .ZN(new_n28782_));
  NOR2_X1    g26346(.A1(new_n8510_), .A2(pi1144), .ZN(new_n28783_));
  AOI21_X1   g26347(.A1(new_n8510_), .A2(new_n3512_), .B(new_n28783_), .ZN(new_n28784_));
  AOI22_X1   g26348(.A1(new_n28669_), .A2(new_n28784_), .B1(new_n8809_), .B2(new_n28063_), .ZN(new_n28785_));
  NOR2_X1    g26349(.A1(new_n28785_), .A2(pi0219), .ZN(new_n28786_));
  OAI21_X1   g26350(.A1(new_n28786_), .A2(new_n28782_), .B(new_n28059_), .ZN(new_n28787_));
  INV_X1     g26351(.I(new_n28787_), .ZN(new_n28788_));
  NOR2_X1    g26352(.A1(new_n8525_), .A2(pi1143), .ZN(new_n28789_));
  NOR2_X1    g26353(.A1(pi0199), .A2(pi1144), .ZN(new_n28790_));
  OAI21_X1   g26354(.A1(new_n28789_), .A2(new_n28790_), .B(new_n8531_), .ZN(new_n28791_));
  NAND3_X1   g26355(.A1(new_n28036_), .A2(new_n28380_), .A3(new_n28791_), .ZN(new_n28792_));
  OAI21_X1   g26356(.A1(new_n2446_), .A2(pi0199), .B(pi0200), .ZN(new_n28793_));
  NOR2_X1    g26357(.A1(new_n3512_), .A2(pi0199), .ZN(new_n28794_));
  INV_X1     g26358(.I(new_n28794_), .ZN(new_n28795_));
  NAND2_X1   g26359(.A1(new_n28795_), .A2(new_n8531_), .ZN(new_n28796_));
  NOR2_X1    g26360(.A1(new_n8525_), .A2(new_n3605_), .ZN(new_n28797_));
  NOR2_X1    g26361(.A1(new_n28796_), .A2(new_n28797_), .ZN(new_n28798_));
  INV_X1     g26362(.I(new_n28798_), .ZN(new_n28799_));
  NAND3_X1   g26363(.A1(new_n28799_), .A2(new_n28372_), .A3(new_n28793_), .ZN(new_n28800_));
  AOI21_X1   g26364(.A1(new_n28800_), .A2(new_n28792_), .B(pi0299), .ZN(new_n28801_));
  INV_X1     g26365(.I(new_n28801_), .ZN(new_n28802_));
  INV_X1     g26366(.I(new_n28785_), .ZN(new_n28803_));
  NOR2_X1    g26367(.A1(new_n28056_), .A2(new_n2628_), .ZN(new_n28804_));
  AOI22_X1   g26368(.A1(new_n28803_), .A2(new_n10289_), .B1(new_n28782_), .B2(new_n28804_), .ZN(new_n28805_));
  AOI21_X1   g26369(.A1(new_n28802_), .A2(new_n28805_), .B(po1038), .ZN(new_n28806_));
  OR3_X2     g26370(.A1(new_n28806_), .A2(new_n26198_), .A3(new_n28788_), .Z(new_n28807_));
  NOR2_X1    g26371(.A1(new_n8510_), .A2(new_n12965_), .ZN(new_n28808_));
  NOR2_X1    g26372(.A1(new_n12745_), .A2(pi0211), .ZN(new_n28809_));
  OAI21_X1   g26373(.A1(new_n28808_), .A2(new_n28809_), .B(new_n28020_), .ZN(new_n28810_));
  NAND2_X1   g26374(.A1(new_n28729_), .A2(new_n28810_), .ZN(new_n28811_));
  AOI21_X1   g26375(.A1(new_n28013_), .A2(new_n28020_), .B(new_n8807_), .ZN(new_n28812_));
  NAND2_X1   g26376(.A1(pi0214), .A2(pi1154), .ZN(new_n28813_));
  OAI21_X1   g26377(.A1(pi0214), .A2(new_n12770_), .B(new_n28813_), .ZN(new_n28814_));
  NAND4_X1   g26378(.A1(po1038), .A2(new_n28814_), .A3(new_n8510_), .A4(pi0212), .ZN(new_n28815_));
  OAI21_X1   g26379(.A1(new_n6643_), .A2(new_n28812_), .B(new_n28815_), .ZN(new_n28816_));
  AOI21_X1   g26380(.A1(new_n28811_), .A2(new_n28816_), .B(pi0213), .ZN(new_n28817_));
  NOR2_X1    g26381(.A1(new_n8509_), .A2(new_n2628_), .ZN(new_n28818_));
  AOI22_X1   g26382(.A1(new_n28814_), .A2(new_n28818_), .B1(new_n28020_), .B2(new_n28269_), .ZN(new_n28819_));
  NOR2_X1    g26383(.A1(new_n28819_), .A2(new_n28044_), .ZN(new_n28820_));
  AOI21_X1   g26384(.A1(new_n28729_), .A2(new_n28810_), .B(new_n28045_), .ZN(new_n28821_));
  NOR3_X1    g26385(.A1(new_n28821_), .A2(new_n28801_), .A3(new_n28820_), .ZN(new_n28822_));
  OAI21_X1   g26386(.A1(new_n28822_), .A2(po1038), .B(new_n28817_), .ZN(new_n28823_));
  NAND3_X1   g26387(.A1(new_n28807_), .A2(pi0209), .A3(new_n28823_), .ZN(new_n28824_));
  INV_X1     g26388(.I(new_n28041_), .ZN(new_n28825_));
  INV_X1     g26389(.I(new_n10288_), .ZN(new_n28826_));
  NOR2_X1    g26390(.A1(new_n28826_), .A2(new_n12745_), .ZN(new_n28827_));
  INV_X1     g26391(.I(new_n28827_), .ZN(new_n28828_));
  AOI22_X1   g26392(.A1(new_n28828_), .A2(new_n12742_), .B1(new_n8525_), .B2(new_n12745_), .ZN(new_n28829_));
  INV_X1     g26393(.I(new_n28829_), .ZN(new_n28830_));
  NOR3_X1    g26394(.A1(new_n28830_), .A2(new_n28136_), .A3(new_n28825_), .ZN(new_n28831_));
  NAND2_X1   g26395(.A1(new_n28191_), .A2(pi0207), .ZN(new_n28832_));
  NAND2_X1   g26396(.A1(new_n28627_), .A2(new_n8521_), .ZN(new_n28833_));
  AOI21_X1   g26397(.A1(new_n28832_), .A2(new_n28833_), .B(new_n8522_), .ZN(new_n28834_));
  OAI21_X1   g26398(.A1(new_n28834_), .A2(new_n28831_), .B(new_n12965_), .ZN(new_n28835_));
  NAND2_X1   g26399(.A1(new_n28204_), .A2(new_n8521_), .ZN(new_n28836_));
  AOI21_X1   g26400(.A1(new_n28832_), .A2(new_n28836_), .B(new_n8522_), .ZN(new_n28837_));
  NAND2_X1   g26401(.A1(new_n8531_), .A2(pi1156), .ZN(new_n28838_));
  AOI22_X1   g26402(.A1(new_n28838_), .A2(pi0199), .B1(new_n12745_), .B2(new_n8640_), .ZN(new_n28839_));
  INV_X1     g26403(.I(new_n28839_), .ZN(new_n28840_));
  NOR2_X1    g26404(.A1(new_n28840_), .A2(new_n28027_), .ZN(new_n28841_));
  INV_X1     g26405(.I(new_n28841_), .ZN(new_n28842_));
  NOR2_X1    g26406(.A1(new_n28842_), .A2(pi0208), .ZN(new_n28843_));
  OAI21_X1   g26407(.A1(new_n28837_), .A2(new_n28843_), .B(pi1157), .ZN(new_n28844_));
  NAND2_X1   g26408(.A1(new_n28835_), .A2(new_n28844_), .ZN(new_n28845_));
  INV_X1     g26409(.I(new_n28845_), .ZN(new_n28846_));
  NAND2_X1   g26410(.A1(new_n28846_), .A2(new_n28503_), .ZN(new_n28847_));
  INV_X1     g26411(.I(new_n28243_), .ZN(new_n28848_));
  OAI21_X1   g26412(.A1(new_n28250_), .A2(new_n8521_), .B(pi0208), .ZN(new_n28849_));
  NAND2_X1   g26413(.A1(new_n8640_), .A2(pi1157), .ZN(new_n28850_));
  NOR2_X1    g26414(.A1(new_n28116_), .A2(pi0299), .ZN(new_n28851_));
  AOI21_X1   g26415(.A1(new_n28851_), .A2(new_n28850_), .B(pi0207), .ZN(new_n28852_));
  AOI21_X1   g26416(.A1(new_n28848_), .A2(new_n28852_), .B(new_n28849_), .ZN(new_n28853_));
  INV_X1     g26417(.I(new_n28465_), .ZN(new_n28854_));
  AOI21_X1   g26418(.A1(new_n28126_), .A2(new_n12745_), .B(new_n12742_), .ZN(new_n28855_));
  NAND2_X1   g26419(.A1(new_n8531_), .A2(new_n12745_), .ZN(new_n28856_));
  AOI22_X1   g26420(.A1(new_n28855_), .A2(new_n28854_), .B1(new_n8525_), .B2(new_n28856_), .ZN(new_n28857_));
  NOR2_X1    g26421(.A1(new_n28857_), .A2(new_n28027_), .ZN(new_n28858_));
  NOR2_X1    g26422(.A1(new_n8521_), .A2(pi0200), .ZN(new_n28859_));
  INV_X1     g26423(.I(new_n28859_), .ZN(new_n28860_));
  NOR2_X1    g26424(.A1(new_n28830_), .A2(new_n28860_), .ZN(new_n28861_));
  OAI21_X1   g26425(.A1(new_n28861_), .A2(pi1157), .B(new_n28858_), .ZN(new_n28862_));
  NOR2_X1    g26426(.A1(new_n28862_), .A2(pi0208), .ZN(new_n28863_));
  NOR2_X1    g26427(.A1(new_n28863_), .A2(pi0208), .ZN(new_n28864_));
  AOI21_X1   g26428(.A1(new_n28864_), .A2(new_n28242_), .B(new_n28853_), .ZN(new_n28865_));
  OAI21_X1   g26429(.A1(new_n28865_), .A2(new_n28503_), .B(new_n28847_), .ZN(new_n28866_));
  AOI21_X1   g26430(.A1(new_n28866_), .A2(pi0219), .B(po1038), .ZN(new_n28867_));
  NOR2_X1    g26431(.A1(new_n28231_), .A2(new_n8521_), .ZN(new_n28868_));
  NOR2_X1    g26432(.A1(new_n28868_), .A2(new_n8522_), .ZN(new_n28869_));
  INV_X1     g26433(.I(new_n28219_), .ZN(new_n28870_));
  NAND2_X1   g26434(.A1(new_n28852_), .A2(new_n28870_), .ZN(new_n28871_));
  AOI22_X1   g26435(.A1(new_n28869_), .A2(new_n28871_), .B1(new_n28223_), .B2(new_n28864_), .ZN(new_n28872_));
  NOR2_X1    g26436(.A1(new_n28872_), .A2(pi0211), .ZN(new_n28873_));
  NOR2_X1    g26437(.A1(new_n28865_), .A2(new_n8510_), .ZN(new_n28874_));
  OAI21_X1   g26438(.A1(new_n28873_), .A2(new_n28874_), .B(pi0214), .ZN(new_n28875_));
  NOR2_X1    g26439(.A1(new_n2628_), .A2(pi1145), .ZN(new_n28876_));
  INV_X1     g26440(.I(new_n28876_), .ZN(new_n28877_));
  AOI21_X1   g26441(.A1(new_n28852_), .A2(new_n28877_), .B(new_n8522_), .ZN(new_n28878_));
  NOR2_X1    g26442(.A1(new_n2628_), .A2(new_n3512_), .ZN(new_n28879_));
  INV_X1     g26443(.I(new_n28879_), .ZN(new_n28880_));
  NAND2_X1   g26444(.A1(new_n28245_), .A2(new_n28880_), .ZN(new_n28881_));
  OAI21_X1   g26445(.A1(new_n28158_), .A2(new_n28876_), .B(new_n12785_), .ZN(new_n28882_));
  NAND3_X1   g26446(.A1(new_n28881_), .A2(pi1156), .A3(new_n28882_), .ZN(new_n28883_));
  AOI21_X1   g26447(.A1(new_n28185_), .A2(new_n28880_), .B(pi1156), .ZN(new_n28884_));
  OAI21_X1   g26448(.A1(new_n28156_), .A2(new_n28876_), .B(pi1154), .ZN(new_n28885_));
  NAND2_X1   g26449(.A1(new_n28885_), .A2(new_n28884_), .ZN(new_n28886_));
  NAND2_X1   g26450(.A1(new_n28886_), .A2(new_n28883_), .ZN(new_n28887_));
  NAND2_X1   g26451(.A1(new_n28887_), .A2(pi0207), .ZN(new_n28888_));
  NAND2_X1   g26452(.A1(new_n28888_), .A2(new_n28878_), .ZN(new_n28889_));
  NOR2_X1    g26453(.A1(new_n28126_), .A2(new_n28285_), .ZN(new_n28890_));
  INV_X1     g26454(.I(new_n28890_), .ZN(new_n28891_));
  NOR2_X1    g26455(.A1(new_n28827_), .A2(new_n12965_), .ZN(new_n28892_));
  AOI21_X1   g26456(.A1(new_n28891_), .A2(new_n28892_), .B(new_n8521_), .ZN(new_n28893_));
  INV_X1     g26457(.I(new_n28123_), .ZN(new_n28894_));
  NOR2_X1    g26458(.A1(new_n28894_), .A2(new_n12742_), .ZN(new_n28895_));
  AOI21_X1   g26459(.A1(new_n28895_), .A2(new_n2628_), .B(pi1157), .ZN(new_n28896_));
  NAND2_X1   g26460(.A1(new_n28828_), .A2(new_n28896_), .ZN(new_n28897_));
  AOI21_X1   g26461(.A1(new_n28893_), .A2(new_n28897_), .B(pi0208), .ZN(new_n28898_));
  AOI21_X1   g26462(.A1(new_n28898_), .A2(new_n28880_), .B(pi0211), .ZN(new_n28899_));
  AOI22_X1   g26463(.A1(new_n28872_), .A2(pi0211), .B1(new_n28889_), .B2(new_n28899_), .ZN(new_n28900_));
  NAND2_X1   g26464(.A1(new_n28900_), .A2(new_n8511_), .ZN(new_n28901_));
  NAND3_X1   g26465(.A1(new_n28901_), .A2(new_n28875_), .A3(pi0212), .ZN(new_n28902_));
  AOI21_X1   g26466(.A1(new_n28846_), .A2(new_n8511_), .B(pi0212), .ZN(new_n28903_));
  NAND2_X1   g26467(.A1(new_n28900_), .A2(pi0214), .ZN(new_n28904_));
  NAND2_X1   g26468(.A1(new_n28904_), .A2(new_n28903_), .ZN(new_n28905_));
  NAND3_X1   g26469(.A1(new_n28902_), .A2(new_n28905_), .A3(new_n8807_), .ZN(new_n28906_));
  AOI21_X1   g26470(.A1(new_n28906_), .A2(new_n28867_), .B(new_n26198_), .ZN(new_n28907_));
  AOI21_X1   g26471(.A1(new_n28907_), .A2(new_n28787_), .B(pi0209), .ZN(new_n28908_));
  NOR2_X1    g26472(.A1(new_n28831_), .A2(pi1157), .ZN(new_n28909_));
  NAND2_X1   g26473(.A1(new_n28909_), .A2(new_n28658_), .ZN(new_n28910_));
  OR2_X2     g26474(.A1(new_n28107_), .A2(new_n28310_), .Z(new_n28911_));
  OAI21_X1   g26475(.A1(new_n28911_), .A2(pi0207), .B(pi1157), .ZN(new_n28912_));
  NAND2_X1   g26476(.A1(new_n28566_), .A2(pi0208), .ZN(new_n28913_));
  AOI21_X1   g26477(.A1(new_n28910_), .A2(new_n28912_), .B(new_n28913_), .ZN(new_n28914_));
  NOR3_X1    g26478(.A1(new_n28909_), .A2(new_n28027_), .A3(new_n28857_), .ZN(new_n28915_));
  NOR3_X1    g26479(.A1(new_n28915_), .A2(pi0208), .A3(new_n28048_), .ZN(new_n28916_));
  NOR3_X1    g26480(.A1(new_n28914_), .A2(new_n8511_), .A3(new_n28916_), .ZN(new_n28917_));
  OAI21_X1   g26481(.A1(new_n28858_), .A2(new_n28051_), .B(new_n28235_), .ZN(new_n28918_));
  AOI21_X1   g26482(.A1(new_n28190_), .A2(new_n28282_), .B(new_n8521_), .ZN(new_n28919_));
  OAI21_X1   g26483(.A1(new_n28919_), .A2(new_n28672_), .B(new_n28670_), .ZN(new_n28920_));
  NOR3_X1    g26484(.A1(new_n28675_), .A2(new_n8522_), .A3(new_n28919_), .ZN(new_n28921_));
  AOI21_X1   g26485(.A1(new_n8522_), .A2(new_n28282_), .B(new_n28921_), .ZN(new_n28922_));
  OAI21_X1   g26486(.A1(new_n28922_), .A2(new_n28831_), .B(new_n12965_), .ZN(new_n28923_));
  AND3_X2    g26487(.A1(new_n28923_), .A2(new_n28918_), .A3(new_n28920_), .Z(new_n28924_));
  OAI21_X1   g26488(.A1(new_n28924_), .A2(pi0214), .B(pi0212), .ZN(new_n28925_));
  OAI21_X1   g26489(.A1(new_n28603_), .A2(new_n28756_), .B(new_n28670_), .ZN(new_n28926_));
  NAND2_X1   g26490(.A1(new_n28842_), .A2(new_n28516_), .ZN(new_n28927_));
  NOR2_X1    g26491(.A1(new_n28861_), .A2(pi0208), .ZN(new_n28928_));
  AOI21_X1   g26492(.A1(new_n28928_), .A2(new_n28516_), .B(pi1157), .ZN(new_n28929_));
  NAND3_X1   g26493(.A1(new_n28604_), .A2(new_n28637_), .A3(pi0208), .ZN(new_n28930_));
  AOI22_X1   g26494(.A1(new_n28929_), .A2(new_n28930_), .B1(new_n28235_), .B2(new_n28927_), .ZN(new_n28931_));
  NAND2_X1   g26495(.A1(new_n28931_), .A2(new_n28926_), .ZN(new_n28932_));
  OAI22_X1   g26496(.A1(new_n28925_), .A2(new_n28917_), .B1(new_n28021_), .B2(new_n28932_), .ZN(new_n28933_));
  NAND2_X1   g26497(.A1(new_n28933_), .A2(new_n8510_), .ZN(new_n28934_));
  AOI21_X1   g26498(.A1(new_n28934_), .A2(new_n28847_), .B(new_n8807_), .ZN(new_n28935_));
  AOI21_X1   g26499(.A1(new_n28840_), .A2(new_n2628_), .B(new_n28098_), .ZN(new_n28936_));
  AOI21_X1   g26500(.A1(new_n28558_), .A2(new_n28641_), .B(new_n28936_), .ZN(new_n28937_));
  OAI21_X1   g26501(.A1(new_n28937_), .A2(new_n12965_), .B(new_n28835_), .ZN(new_n28938_));
  AOI22_X1   g26502(.A1(new_n28938_), .A2(new_n28267_), .B1(new_n28298_), .B2(new_n28932_), .ZN(new_n28939_));
  OR2_X2     g26503(.A1(new_n28924_), .A2(new_n8513_), .Z(new_n28940_));
  AOI21_X1   g26504(.A1(new_n28940_), .A2(new_n28939_), .B(new_n8509_), .ZN(new_n28941_));
  INV_X1     g26505(.I(new_n28903_), .ZN(new_n28942_));
  AOI21_X1   g26506(.A1(new_n8640_), .A2(pi0207), .B(pi0299), .ZN(new_n28943_));
  INV_X1     g26507(.I(new_n28943_), .ZN(new_n28944_));
  NAND2_X1   g26508(.A1(new_n28944_), .A2(pi1158), .ZN(new_n28945_));
  NAND2_X1   g26509(.A1(new_n28895_), .A2(new_n28026_), .ZN(new_n28946_));
  NAND3_X1   g26510(.A1(new_n28946_), .A2(new_n8522_), .A3(new_n28945_), .ZN(new_n28947_));
  AOI21_X1   g26511(.A1(new_n12745_), .A2(pi0299), .B(pi0207), .ZN(new_n28948_));
  INV_X1     g26512(.I(new_n28948_), .ZN(new_n28949_));
  NOR2_X1    g26513(.A1(new_n28851_), .A2(new_n28949_), .ZN(new_n28950_));
  NOR2_X1    g26514(.A1(new_n28950_), .A2(new_n8522_), .ZN(new_n28951_));
  NOR2_X1    g26515(.A1(new_n28190_), .A2(pi1158), .ZN(new_n28952_));
  AOI21_X1   g26516(.A1(new_n28330_), .A2(pi1158), .B(new_n28952_), .ZN(new_n28953_));
  OAI21_X1   g26517(.A1(new_n28953_), .A2(new_n8521_), .B(new_n28951_), .ZN(new_n28954_));
  NAND3_X1   g26518(.A1(new_n28954_), .A2(new_n12965_), .A3(new_n28947_), .ZN(new_n28955_));
  INV_X1     g26519(.I(new_n28893_), .ZN(new_n28956_));
  NAND2_X1   g26520(.A1(new_n28956_), .A2(new_n28945_), .ZN(new_n28957_));
  AOI21_X1   g26521(.A1(new_n28957_), .A2(new_n28235_), .B(pi0211), .ZN(new_n28958_));
  OAI22_X1   g26522(.A1(new_n28953_), .A2(new_n8521_), .B1(new_n28107_), .B2(new_n28949_), .ZN(new_n28959_));
  NAND2_X1   g26523(.A1(new_n28959_), .A2(new_n28670_), .ZN(new_n28960_));
  NAND3_X1   g26524(.A1(new_n28960_), .A2(new_n28955_), .A3(new_n28958_), .ZN(new_n28961_));
  OR2_X2     g26525(.A1(new_n28938_), .A2(new_n8510_), .Z(new_n28962_));
  AOI21_X1   g26526(.A1(new_n28961_), .A2(new_n28962_), .B(new_n8511_), .ZN(new_n28963_));
  OAI21_X1   g26527(.A1(new_n28963_), .A2(new_n28942_), .B(new_n8807_), .ZN(new_n28964_));
  OAI21_X1   g26528(.A1(new_n28964_), .A2(new_n28941_), .B(new_n6643_), .ZN(new_n28965_));
  OAI21_X1   g26529(.A1(new_n28935_), .A2(new_n28965_), .B(new_n28817_), .ZN(new_n28966_));
  AOI21_X1   g26530(.A1(new_n28908_), .A2(new_n28966_), .B(new_n27999_), .ZN(new_n28967_));
  AOI22_X1   g26531(.A1(new_n28967_), .A2(new_n28824_), .B1(new_n27999_), .B2(pi0237), .ZN(po0394));
  NOR2_X1    g26532(.A1(pi0211), .A2(pi1153), .ZN(new_n28969_));
  NAND2_X1   g26533(.A1(new_n28969_), .A2(pi0219), .ZN(new_n28970_));
  AND3_X2    g26534(.A1(new_n28059_), .A2(new_n28720_), .A3(new_n28970_), .Z(new_n28971_));
  INV_X1     g26535(.I(new_n28686_), .ZN(new_n28972_));
  NOR3_X1    g26536(.A1(new_n28126_), .A2(new_n12841_), .A3(pi1154), .ZN(new_n28973_));
  NOR3_X1    g26537(.A1(new_n28454_), .A2(new_n8524_), .A3(new_n28973_), .ZN(new_n28974_));
  NOR2_X1    g26538(.A1(new_n28972_), .A2(new_n28974_), .ZN(new_n28975_));
  NOR2_X1    g26539(.A1(new_n28975_), .A2(new_n8510_), .ZN(new_n28976_));
  INV_X1     g26540(.I(new_n28976_), .ZN(new_n28977_));
  NOR2_X1    g26541(.A1(new_n28154_), .A2(new_n12841_), .ZN(new_n28978_));
  OAI21_X1   g26542(.A1(new_n28454_), .A2(new_n28978_), .B(pi0207), .ZN(new_n28979_));
  AOI21_X1   g26543(.A1(new_n28692_), .A2(new_n28979_), .B(new_n8522_), .ZN(new_n28980_));
  NOR2_X1    g26544(.A1(new_n28690_), .A2(new_n28980_), .ZN(new_n28981_));
  NAND2_X1   g26545(.A1(new_n28981_), .A2(new_n8510_), .ZN(new_n28982_));
  NAND2_X1   g26546(.A1(new_n28982_), .A2(new_n28977_), .ZN(new_n28983_));
  NAND2_X1   g26547(.A1(new_n28983_), .A2(new_n28525_), .ZN(new_n28984_));
  INV_X1     g26548(.I(new_n28973_), .ZN(new_n28985_));
  NOR2_X1    g26549(.A1(new_n28479_), .A2(new_n8521_), .ZN(new_n28986_));
  AOI21_X1   g26550(.A1(new_n28985_), .A2(new_n28986_), .B(new_n28701_), .ZN(new_n28987_));
  AOI21_X1   g26551(.A1(new_n28987_), .A2(pi0208), .B(new_n28699_), .ZN(new_n28988_));
  NAND2_X1   g26552(.A1(new_n28988_), .A2(pi0211), .ZN(new_n28989_));
  OAI21_X1   g26553(.A1(new_n28124_), .A2(new_n12841_), .B(new_n2628_), .ZN(new_n28990_));
  NAND2_X1   g26554(.A1(new_n28990_), .A2(new_n12785_), .ZN(new_n28991_));
  AOI21_X1   g26555(.A1(new_n28986_), .A2(new_n28991_), .B(new_n8522_), .ZN(new_n28992_));
  NAND2_X1   g26556(.A1(new_n28538_), .A2(new_n28448_), .ZN(new_n28993_));
  NAND2_X1   g26557(.A1(new_n28992_), .A2(new_n28993_), .ZN(new_n28994_));
  NAND2_X1   g26558(.A1(new_n28994_), .A2(new_n28705_), .ZN(new_n28995_));
  NAND2_X1   g26559(.A1(new_n28995_), .A2(new_n28707_), .ZN(new_n28996_));
  NAND2_X1   g26560(.A1(new_n28996_), .A2(new_n8510_), .ZN(new_n28997_));
  AOI21_X1   g26561(.A1(new_n28997_), .A2(new_n28989_), .B(new_n28021_), .ZN(new_n28998_));
  NOR2_X1    g26562(.A1(new_n28988_), .A2(new_n28297_), .ZN(new_n28999_));
  NOR2_X1    g26563(.A1(new_n28981_), .A2(new_n8513_), .ZN(new_n29000_));
  NOR2_X1    g26564(.A1(new_n28996_), .A2(new_n28268_), .ZN(new_n29001_));
  NOR4_X1    g26565(.A1(new_n29001_), .A2(new_n8509_), .A3(new_n28999_), .A4(new_n29000_), .ZN(new_n29002_));
  OAI21_X1   g26566(.A1(new_n29002_), .A2(new_n28998_), .B(new_n8807_), .ZN(new_n29003_));
  NOR2_X1    g26567(.A1(new_n28975_), .A2(new_n28430_), .ZN(new_n29004_));
  INV_X1     g26568(.I(new_n29004_), .ZN(new_n29005_));
  NAND4_X1   g26569(.A1(new_n29003_), .A2(new_n6643_), .A3(new_n28984_), .A4(new_n29005_), .ZN(new_n29006_));
  NOR2_X1    g26570(.A1(po1038), .A2(pi1151), .ZN(new_n29007_));
  INV_X1     g26571(.I(new_n28525_), .ZN(new_n29008_));
  AOI21_X1   g26572(.A1(new_n28371_), .A2(new_n28860_), .B(new_n9183_), .ZN(new_n29009_));
  INV_X1     g26573(.I(new_n29009_), .ZN(new_n29010_));
  AOI21_X1   g26574(.A1(new_n8524_), .A2(new_n28437_), .B(new_n29010_), .ZN(new_n29011_));
  INV_X1     g26575(.I(new_n29011_), .ZN(new_n29012_));
  NOR2_X1    g26576(.A1(new_n28411_), .A2(pi0211), .ZN(new_n29013_));
  INV_X1     g26577(.I(new_n29013_), .ZN(new_n29014_));
  OAI22_X1   g26578(.A1(new_n29012_), .A2(new_n28094_), .B1(new_n29008_), .B2(new_n29014_), .ZN(new_n29015_));
  AOI21_X1   g26579(.A1(new_n8521_), .A2(new_n28438_), .B(new_n28944_), .ZN(new_n29016_));
  OAI22_X1   g26580(.A1(new_n29016_), .A2(new_n8522_), .B1(new_n28098_), .B2(new_n28439_), .ZN(new_n29017_));
  INV_X1     g26581(.I(new_n29017_), .ZN(new_n29018_));
  NOR3_X1    g26582(.A1(new_n29018_), .A2(pi0211), .A3(new_n28310_), .ZN(new_n29019_));
  NOR2_X1    g26583(.A1(new_n8641_), .A2(pi0207), .ZN(new_n29020_));
  NOR2_X1    g26584(.A1(new_n29020_), .A2(pi0299), .ZN(new_n29021_));
  AOI21_X1   g26585(.A1(pi0200), .A2(pi0207), .B(pi0199), .ZN(new_n29022_));
  OAI21_X1   g26586(.A1(new_n29022_), .A2(pi0299), .B(pi0208), .ZN(new_n29023_));
  INV_X1     g26587(.I(new_n29023_), .ZN(new_n29024_));
  OAI21_X1   g26588(.A1(new_n29021_), .A2(pi1153), .B(new_n29024_), .ZN(new_n29025_));
  NAND3_X1   g26589(.A1(new_n28373_), .A2(new_n28391_), .A3(pi0207), .ZN(new_n29026_));
  NAND3_X1   g26590(.A1(new_n29026_), .A2(new_n8522_), .A3(new_n28473_), .ZN(new_n29027_));
  AOI21_X1   g26591(.A1(new_n29027_), .A2(new_n29025_), .B(new_n8510_), .ZN(new_n29028_));
  OAI21_X1   g26592(.A1(new_n29019_), .A2(new_n29028_), .B(new_n8809_), .ZN(new_n29029_));
  NAND2_X1   g26593(.A1(new_n28718_), .A2(pi0299), .ZN(new_n29030_));
  NOR2_X1    g26594(.A1(new_n29018_), .A2(new_n28066_), .ZN(new_n29031_));
  NAND2_X1   g26595(.A1(new_n29031_), .A2(new_n29030_), .ZN(new_n29032_));
  AOI21_X1   g26596(.A1(new_n29029_), .A2(new_n29032_), .B(pi0219), .ZN(new_n29033_));
  OAI21_X1   g26597(.A1(new_n29033_), .A2(new_n29015_), .B(new_n29007_), .ZN(new_n29034_));
  INV_X1     g26598(.I(pi1151), .ZN(new_n29035_));
  NOR2_X1    g26599(.A1(po1038), .A2(new_n29035_), .ZN(new_n29036_));
  INV_X1     g26600(.I(new_n29036_), .ZN(new_n29037_));
  NOR2_X1    g26601(.A1(new_n28826_), .A2(new_n28371_), .ZN(new_n29038_));
  NOR2_X1    g26602(.A1(new_n29038_), .A2(pi0214), .ZN(new_n29039_));
  INV_X1     g26603(.I(new_n29039_), .ZN(new_n29040_));
  NOR2_X1    g26604(.A1(new_n29040_), .A2(pi0212), .ZN(new_n29041_));
  NOR2_X1    g26605(.A1(new_n28371_), .A2(new_n8641_), .ZN(new_n29042_));
  NOR2_X1    g26606(.A1(new_n29042_), .A2(pi0299), .ZN(new_n29043_));
  NOR2_X1    g26607(.A1(new_n8510_), .A2(new_n2628_), .ZN(new_n29044_));
  NOR2_X1    g26608(.A1(new_n29043_), .A2(new_n29044_), .ZN(new_n29045_));
  INV_X1     g26609(.I(new_n29045_), .ZN(new_n29046_));
  NOR2_X1    g26610(.A1(new_n29041_), .A2(new_n29046_), .ZN(new_n29047_));
  INV_X1     g26611(.I(new_n29047_), .ZN(new_n29048_));
  NOR2_X1    g26612(.A1(new_n29048_), .A2(new_n12841_), .ZN(new_n29049_));
  INV_X1     g26613(.I(new_n29049_), .ZN(new_n29050_));
  NOR3_X1    g26614(.A1(new_n28448_), .A2(new_n8522_), .A3(new_n29020_), .ZN(new_n29051_));
  NOR2_X1    g26615(.A1(new_n28124_), .A2(new_n28027_), .ZN(new_n29052_));
  NOR2_X1    g26616(.A1(new_n29051_), .A2(new_n29052_), .ZN(new_n29053_));
  INV_X1     g26617(.I(new_n29053_), .ZN(new_n29054_));
  NOR2_X1    g26618(.A1(new_n29054_), .A2(new_n8807_), .ZN(new_n29055_));
  AOI21_X1   g26619(.A1(new_n29050_), .A2(new_n29055_), .B(new_n29037_), .ZN(new_n29056_));
  OR2_X2     g26620(.A1(new_n29019_), .A2(new_n29054_), .Z(new_n29057_));
  NOR3_X1    g26621(.A1(new_n29043_), .A2(new_n8510_), .A3(new_n12841_), .ZN(new_n29058_));
  OAI21_X1   g26622(.A1(new_n29057_), .A2(new_n29058_), .B(new_n8809_), .ZN(new_n29059_));
  INV_X1     g26623(.I(new_n29038_), .ZN(new_n29060_));
  NOR2_X1    g26624(.A1(new_n29060_), .A2(new_n12841_), .ZN(new_n29061_));
  NOR2_X1    g26625(.A1(new_n29054_), .A2(pi0214), .ZN(new_n29062_));
  INV_X1     g26626(.I(new_n29062_), .ZN(new_n29063_));
  NOR2_X1    g26627(.A1(new_n29063_), .A2(new_n29061_), .ZN(new_n29064_));
  NOR2_X1    g26628(.A1(new_n29064_), .A2(pi0212), .ZN(new_n29065_));
  NAND2_X1   g26629(.A1(new_n29065_), .A2(new_n8511_), .ZN(new_n29066_));
  AOI21_X1   g26630(.A1(new_n28467_), .A2(new_n28441_), .B(new_n8522_), .ZN(new_n29067_));
  AOI21_X1   g26631(.A1(new_n28441_), .A2(pi0207), .B(new_n28098_), .ZN(new_n29068_));
  NOR2_X1    g26632(.A1(new_n29067_), .A2(new_n29068_), .ZN(new_n29069_));
  INV_X1     g26633(.I(new_n29069_), .ZN(new_n29070_));
  NAND3_X1   g26634(.A1(new_n29070_), .A2(new_n28065_), .A3(new_n29030_), .ZN(new_n29071_));
  NAND4_X1   g26635(.A1(new_n29066_), .A2(new_n8807_), .A3(new_n29059_), .A4(new_n29071_), .ZN(new_n29072_));
  NAND2_X1   g26636(.A1(new_n29072_), .A2(new_n29056_), .ZN(new_n29073_));
  NAND3_X1   g26637(.A1(new_n29073_), .A2(pi1152), .A3(new_n29034_), .ZN(new_n29074_));
  NAND2_X1   g26638(.A1(new_n28153_), .A2(new_n28380_), .ZN(new_n29075_));
  NAND2_X1   g26639(.A1(new_n28621_), .A2(new_n8761_), .ZN(new_n29076_));
  OAI21_X1   g26640(.A1(new_n8523_), .A2(new_n29076_), .B(new_n29075_), .ZN(new_n29077_));
  INV_X1     g26641(.I(new_n29077_), .ZN(new_n29078_));
  NOR2_X1    g26642(.A1(new_n29078_), .A2(new_n28449_), .ZN(new_n29079_));
  NOR2_X1    g26643(.A1(new_n29079_), .A2(new_n28430_), .ZN(new_n29080_));
  INV_X1     g26644(.I(new_n29080_), .ZN(new_n29081_));
  AOI21_X1   g26645(.A1(new_n28124_), .A2(new_n28026_), .B(new_n8522_), .ZN(new_n29082_));
  INV_X1     g26646(.I(new_n29082_), .ZN(new_n29083_));
  AOI21_X1   g26647(.A1(new_n8521_), .A2(new_n28102_), .B(new_n29083_), .ZN(new_n29084_));
  AOI21_X1   g26648(.A1(new_n28860_), .A2(new_n2628_), .B(pi0208), .ZN(new_n29085_));
  NOR2_X1    g26649(.A1(new_n29084_), .A2(new_n29085_), .ZN(new_n29086_));
  NOR2_X1    g26650(.A1(new_n29086_), .A2(pi0211), .ZN(new_n29087_));
  NOR2_X1    g26651(.A1(new_n29078_), .A2(new_n8510_), .ZN(new_n29088_));
  NOR2_X1    g26652(.A1(new_n29087_), .A2(new_n29088_), .ZN(new_n29089_));
  NOR2_X1    g26653(.A1(new_n29089_), .A2(new_n28388_), .ZN(new_n29090_));
  NAND2_X1   g26654(.A1(new_n29090_), .A2(new_n29081_), .ZN(new_n29091_));
  INV_X1     g26655(.I(new_n29091_), .ZN(new_n29092_));
  OAI21_X1   g26656(.A1(new_n29092_), .A2(new_n8807_), .B(new_n29036_), .ZN(new_n29093_));
  NOR3_X1    g26657(.A1(new_n29079_), .A2(new_n28048_), .A3(new_n28297_), .ZN(new_n29094_));
  NOR2_X1    g26658(.A1(new_n29086_), .A2(new_n28388_), .ZN(new_n29095_));
  NOR2_X1    g26659(.A1(new_n29095_), .A2(new_n8513_), .ZN(new_n29096_));
  NOR2_X1    g26660(.A1(new_n28136_), .A2(new_n28451_), .ZN(new_n29097_));
  AOI21_X1   g26661(.A1(new_n12841_), .A2(new_n28151_), .B(new_n28133_), .ZN(new_n29098_));
  NAND2_X1   g26662(.A1(new_n29098_), .A2(pi1155), .ZN(new_n29099_));
  INV_X1     g26663(.I(new_n29099_), .ZN(new_n29100_));
  OAI22_X1   g26664(.A1(new_n29100_), .A2(new_n29097_), .B1(new_n28283_), .B2(new_n29082_), .ZN(new_n29101_));
  NAND2_X1   g26665(.A1(new_n29101_), .A2(new_n29075_), .ZN(new_n29102_));
  NOR2_X1    g26666(.A1(new_n29102_), .A2(new_n28268_), .ZN(new_n29103_));
  NOR4_X1    g26667(.A1(new_n29103_), .A2(new_n8509_), .A3(new_n29094_), .A4(new_n29096_), .ZN(new_n29104_));
  OAI21_X1   g26668(.A1(new_n29102_), .A2(pi0299), .B(new_n29030_), .ZN(new_n29105_));
  INV_X1     g26669(.I(new_n29079_), .ZN(new_n29106_));
  AOI21_X1   g26670(.A1(new_n29106_), .A2(new_n8511_), .B(pi0212), .ZN(new_n29107_));
  INV_X1     g26671(.I(new_n29107_), .ZN(new_n29108_));
  AOI21_X1   g26672(.A1(new_n29105_), .A2(pi0214), .B(new_n29108_), .ZN(new_n29109_));
  NOR3_X1    g26673(.A1(new_n29109_), .A2(pi0219), .A3(new_n29104_), .ZN(new_n29110_));
  INV_X1     g26674(.I(new_n29007_), .ZN(new_n29111_));
  AOI21_X1   g26675(.A1(new_n29050_), .A2(new_n28361_), .B(new_n29111_), .ZN(new_n29112_));
  NOR2_X1    g26676(.A1(new_n28718_), .A2(new_n2628_), .ZN(new_n29113_));
  NOR3_X1    g26677(.A1(new_n29061_), .A2(new_n28066_), .A3(new_n29113_), .ZN(new_n29114_));
  INV_X1     g26678(.I(new_n29061_), .ZN(new_n29115_));
  AOI21_X1   g26679(.A1(new_n29115_), .A2(new_n28399_), .B(pi0211), .ZN(new_n29116_));
  NOR3_X1    g26680(.A1(new_n29116_), .A2(new_n8811_), .A3(new_n29058_), .ZN(new_n29117_));
  OAI21_X1   g26681(.A1(new_n29117_), .A2(new_n29114_), .B(new_n8807_), .ZN(new_n29118_));
  AOI21_X1   g26682(.A1(new_n29112_), .A2(new_n29118_), .B(pi1152), .ZN(new_n29119_));
  OAI21_X1   g26683(.A1(new_n29110_), .A2(new_n29093_), .B(new_n29119_), .ZN(new_n29120_));
  AOI21_X1   g26684(.A1(new_n29074_), .A2(new_n29120_), .B(pi0209), .ZN(new_n29121_));
  AOI21_X1   g26685(.A1(new_n29006_), .A2(pi0209), .B(new_n29121_), .ZN(new_n29122_));
  OAI21_X1   g26686(.A1(new_n29122_), .A2(new_n28971_), .B(pi0213), .ZN(new_n29123_));
  NOR2_X1    g26687(.A1(new_n28060_), .A2(new_n8515_), .ZN(new_n29124_));
  NOR2_X1    g26688(.A1(new_n28386_), .A2(new_n6643_), .ZN(new_n29125_));
  INV_X1     g26689(.I(new_n29125_), .ZN(new_n29126_));
  NOR2_X1    g26690(.A1(new_n8813_), .A2(new_n28005_), .ZN(new_n29127_));
  NOR2_X1    g26691(.A1(new_n29126_), .A2(new_n29127_), .ZN(new_n29128_));
  NOR3_X1    g26692(.A1(new_n29128_), .A2(new_n29124_), .A3(new_n29035_), .ZN(new_n29129_));
  AOI21_X1   g26693(.A1(new_n28992_), .A2(new_n28735_), .B(new_n28741_), .ZN(new_n29130_));
  AOI21_X1   g26694(.A1(new_n29130_), .A2(new_n8510_), .B(new_n28976_), .ZN(new_n29131_));
  OAI21_X1   g26695(.A1(new_n29131_), .A2(new_n28056_), .B(new_n29005_), .ZN(new_n29132_));
  NAND2_X1   g26696(.A1(new_n29132_), .A2(pi0219), .ZN(new_n29133_));
  NAND2_X1   g26697(.A1(new_n29133_), .A2(new_n6643_), .ZN(new_n29134_));
  NAND2_X1   g26698(.A1(new_n29130_), .A2(pi0211), .ZN(new_n29135_));
  AND2_X2    g26699(.A1(new_n29135_), .A2(new_n28982_), .Z(new_n29136_));
  NAND2_X1   g26700(.A1(new_n29136_), .A2(new_n8511_), .ZN(new_n29137_));
  OR2_X2     g26701(.A1(new_n29130_), .A2(new_n8511_), .Z(new_n29138_));
  AOI21_X1   g26702(.A1(new_n29137_), .A2(new_n29138_), .B(new_n8509_), .ZN(new_n29139_));
  INV_X1     g26703(.I(new_n28975_), .ZN(new_n29140_));
  NOR2_X1    g26704(.A1(new_n29140_), .A2(pi0214), .ZN(new_n29141_));
  AOI21_X1   g26705(.A1(new_n29136_), .A2(pi0214), .B(new_n29141_), .ZN(new_n29142_));
  OAI21_X1   g26706(.A1(new_n29142_), .A2(pi0212), .B(new_n8807_), .ZN(new_n29143_));
  NOR2_X1    g26707(.A1(new_n29143_), .A2(new_n29139_), .ZN(new_n29144_));
  OAI21_X1   g26708(.A1(new_n29144_), .A2(new_n29134_), .B(new_n29129_), .ZN(new_n29145_));
  NOR2_X1    g26709(.A1(new_n29128_), .A2(pi1151), .ZN(new_n29146_));
  OAI21_X1   g26710(.A1(new_n28975_), .A2(new_n8807_), .B(new_n6643_), .ZN(new_n29147_));
  NAND2_X1   g26711(.A1(new_n29131_), .A2(pi0214), .ZN(new_n29148_));
  AOI21_X1   g26712(.A1(new_n29137_), .A2(new_n29148_), .B(new_n8509_), .ZN(new_n29149_));
  NOR2_X1    g26713(.A1(new_n29143_), .A2(new_n29149_), .ZN(new_n29150_));
  OAI21_X1   g26714(.A1(new_n29150_), .A2(new_n29147_), .B(new_n29146_), .ZN(new_n29151_));
  NAND3_X1   g26715(.A1(new_n29145_), .A2(new_n29151_), .A3(pi1152), .ZN(new_n29152_));
  NOR2_X1    g26716(.A1(new_n28212_), .A2(pi0211), .ZN(new_n29153_));
  INV_X1     g26717(.I(new_n29153_), .ZN(new_n29154_));
  NOR2_X1    g26718(.A1(new_n29154_), .A2(new_n12841_), .ZN(new_n29155_));
  NOR2_X1    g26719(.A1(new_n6643_), .A2(pi0219), .ZN(new_n29156_));
  AOI21_X1   g26720(.A1(new_n29156_), .A2(new_n29155_), .B(pi1151), .ZN(new_n29157_));
  NOR2_X1    g26721(.A1(new_n28212_), .A2(pi0219), .ZN(new_n29158_));
  INV_X1     g26722(.I(new_n29158_), .ZN(new_n29159_));
  NOR2_X1    g26723(.A1(new_n28983_), .A2(new_n29159_), .ZN(new_n29160_));
  NOR2_X1    g26724(.A1(new_n29140_), .A2(new_n29158_), .ZN(new_n29161_));
  OAI21_X1   g26725(.A1(new_n29160_), .A2(new_n29161_), .B(new_n6643_), .ZN(new_n29162_));
  AOI21_X1   g26726(.A1(new_n29162_), .A2(new_n29157_), .B(pi1152), .ZN(new_n29163_));
  NOR2_X1    g26727(.A1(new_n29155_), .A2(new_n8520_), .ZN(new_n29164_));
  OAI21_X1   g26728(.A1(new_n29164_), .A2(new_n28060_), .B(pi1151), .ZN(new_n29165_));
  INV_X1     g26729(.I(new_n29165_), .ZN(new_n29166_));
  NAND2_X1   g26730(.A1(new_n29140_), .A2(new_n8510_), .ZN(new_n29167_));
  AOI21_X1   g26731(.A1(new_n29135_), .A2(new_n29167_), .B(new_n8511_), .ZN(new_n29168_));
  AOI21_X1   g26732(.A1(new_n28982_), .A2(new_n28977_), .B(pi0214), .ZN(new_n29169_));
  OAI21_X1   g26733(.A1(new_n29168_), .A2(new_n29169_), .B(pi0212), .ZN(new_n29170_));
  NOR2_X1    g26734(.A1(new_n29141_), .A2(pi0212), .ZN(new_n29171_));
  OAI21_X1   g26735(.A1(new_n28983_), .A2(new_n8511_), .B(new_n29171_), .ZN(new_n29172_));
  AOI21_X1   g26736(.A1(new_n29170_), .A2(new_n29172_), .B(pi0219), .ZN(new_n29173_));
  OAI21_X1   g26737(.A1(new_n29173_), .A2(new_n29134_), .B(new_n29166_), .ZN(new_n29174_));
  NAND2_X1   g26738(.A1(new_n29174_), .A2(new_n29163_), .ZN(new_n29175_));
  NAND3_X1   g26739(.A1(new_n29152_), .A2(pi0209), .A3(new_n29175_), .ZN(new_n29176_));
  NOR2_X1    g26740(.A1(new_n29061_), .A2(new_n29044_), .ZN(new_n29177_));
  NOR2_X1    g26741(.A1(new_n29177_), .A2(new_n8509_), .ZN(new_n29178_));
  AOI21_X1   g26742(.A1(new_n29178_), .A2(new_n29040_), .B(pi0219), .ZN(new_n29179_));
  INV_X1     g26743(.I(new_n29179_), .ZN(new_n29180_));
  NOR2_X1    g26744(.A1(new_n29014_), .A2(new_n28021_), .ZN(new_n29181_));
  NOR2_X1    g26745(.A1(new_n29050_), .A2(new_n29040_), .ZN(new_n29182_));
  NOR4_X1    g26746(.A1(new_n29182_), .A2(new_n29038_), .A3(new_n29180_), .A4(new_n29181_), .ZN(new_n29183_));
  AOI21_X1   g26747(.A1(new_n29060_), .A2(pi0219), .B(po1038), .ZN(new_n29184_));
  NAND2_X1   g26748(.A1(new_n29049_), .A2(new_n29184_), .ZN(new_n29185_));
  OAI21_X1   g26749(.A1(new_n29183_), .A2(new_n29185_), .B(new_n29157_), .ZN(new_n29186_));
  NOR2_X1    g26750(.A1(new_n2628_), .A2(pi0211), .ZN(new_n29187_));
  INV_X1     g26751(.I(new_n29187_), .ZN(new_n29188_));
  NAND2_X1   g26752(.A1(new_n29115_), .A2(new_n29188_), .ZN(new_n29189_));
  AOI21_X1   g26753(.A1(new_n29189_), .A2(new_n28430_), .B(new_n29079_), .ZN(new_n29190_));
  NAND2_X1   g26754(.A1(new_n29190_), .A2(pi0219), .ZN(new_n29191_));
  NAND2_X1   g26755(.A1(new_n29106_), .A2(new_n29177_), .ZN(new_n29192_));
  NAND2_X1   g26756(.A1(new_n29192_), .A2(pi0214), .ZN(new_n29193_));
  NAND2_X1   g26757(.A1(new_n29193_), .A2(pi0212), .ZN(new_n29194_));
  AOI21_X1   g26758(.A1(new_n29090_), .A2(new_n8511_), .B(new_n29194_), .ZN(new_n29195_));
  NOR2_X1    g26759(.A1(new_n29092_), .A2(pi0212), .ZN(new_n29196_));
  OAI21_X1   g26760(.A1(new_n29196_), .A2(new_n29195_), .B(new_n8807_), .ZN(new_n29197_));
  NAND3_X1   g26761(.A1(new_n29197_), .A2(new_n6643_), .A3(new_n29191_), .ZN(new_n29198_));
  AOI21_X1   g26762(.A1(new_n29198_), .A2(new_n29166_), .B(pi1152), .ZN(new_n29199_));
  INV_X1     g26763(.I(new_n29146_), .ZN(new_n29200_));
  OAI21_X1   g26764(.A1(new_n8811_), .A2(new_n29188_), .B(new_n8807_), .ZN(new_n29201_));
  AOI21_X1   g26765(.A1(new_n29011_), .A2(new_n28212_), .B(new_n29201_), .ZN(new_n29202_));
  NAND3_X1   g26766(.A1(new_n29027_), .A2(new_n8510_), .A3(new_n29025_), .ZN(new_n29203_));
  NAND2_X1   g26767(.A1(new_n29031_), .A2(new_n29203_), .ZN(new_n29204_));
  AOI21_X1   g26768(.A1(new_n29012_), .A2(pi0219), .B(po1038), .ZN(new_n29205_));
  INV_X1     g26769(.I(new_n29205_), .ZN(new_n29206_));
  AOI21_X1   g26770(.A1(new_n29204_), .A2(new_n29202_), .B(new_n29206_), .ZN(new_n29207_));
  OAI21_X1   g26771(.A1(new_n29207_), .A2(new_n29200_), .B(pi1152), .ZN(new_n29208_));
  NOR2_X1    g26772(.A1(new_n29054_), .A2(new_n29061_), .ZN(new_n29209_));
  OAI21_X1   g26773(.A1(new_n29069_), .A2(pi0211), .B(new_n29209_), .ZN(new_n29210_));
  NOR2_X1    g26774(.A1(new_n29210_), .A2(new_n8511_), .ZN(new_n29211_));
  OAI21_X1   g26775(.A1(new_n29211_), .A2(new_n29064_), .B(new_n8509_), .ZN(new_n29212_));
  NAND2_X1   g26776(.A1(new_n29212_), .A2(new_n29210_), .ZN(new_n29213_));
  AOI21_X1   g26777(.A1(new_n29213_), .A2(pi0219), .B(po1038), .ZN(new_n29214_));
  INV_X1     g26778(.I(new_n29065_), .ZN(new_n29215_));
  INV_X1     g26779(.I(new_n29043_), .ZN(new_n29216_));
  AOI22_X1   g26780(.A1(new_n29070_), .A2(pi0211), .B1(pi1153), .B2(new_n29216_), .ZN(new_n29217_));
  NOR2_X1    g26781(.A1(new_n29054_), .A2(new_n8511_), .ZN(new_n29218_));
  AOI21_X1   g26782(.A1(new_n29217_), .A2(new_n29218_), .B(new_n29215_), .ZN(new_n29219_));
  NOR2_X1    g26783(.A1(new_n29070_), .A2(new_n8511_), .ZN(new_n29220_));
  NOR2_X1    g26784(.A1(new_n29220_), .A2(new_n8509_), .ZN(new_n29221_));
  NAND2_X1   g26785(.A1(new_n29217_), .A2(new_n29062_), .ZN(new_n29222_));
  NAND2_X1   g26786(.A1(new_n29222_), .A2(new_n29221_), .ZN(new_n29223_));
  NAND2_X1   g26787(.A1(new_n29223_), .A2(new_n8807_), .ZN(new_n29224_));
  OAI21_X1   g26788(.A1(new_n29219_), .A2(new_n29224_), .B(new_n29214_), .ZN(new_n29225_));
  AOI21_X1   g26789(.A1(new_n29225_), .A2(new_n29129_), .B(new_n29208_), .ZN(new_n29226_));
  AOI21_X1   g26790(.A1(new_n29199_), .A2(new_n29186_), .B(new_n29226_), .ZN(new_n29227_));
  AOI21_X1   g26791(.A1(new_n29227_), .A2(new_n28360_), .B(pi0213), .ZN(new_n29228_));
  AOI21_X1   g26792(.A1(new_n29176_), .A2(new_n29228_), .B(new_n27999_), .ZN(new_n29229_));
  AOI22_X1   g26793(.A1(new_n29229_), .A2(new_n29123_), .B1(new_n27999_), .B2(new_n3625_), .ZN(po0395));
  NOR2_X1    g26794(.A1(new_n6643_), .A2(new_n28352_), .ZN(new_n29231_));
  INV_X1     g26795(.I(new_n29231_), .ZN(new_n29232_));
  OAI21_X1   g26796(.A1(new_n28355_), .A2(pi0219), .B(new_n28020_), .ZN(new_n29233_));
  OAI21_X1   g26797(.A1(new_n29232_), .A2(new_n29233_), .B(new_n26198_), .ZN(new_n29234_));
  NOR2_X1    g26798(.A1(new_n28190_), .A2(new_n28825_), .ZN(new_n29235_));
  INV_X1     g26799(.I(new_n29235_), .ZN(new_n29236_));
  NOR2_X1    g26800(.A1(new_n29236_), .A2(pi0214), .ZN(new_n29237_));
  NOR3_X1    g26801(.A1(new_n29237_), .A2(pi0212), .A3(pi0219), .ZN(new_n29238_));
  INV_X1     g26802(.I(new_n29238_), .ZN(new_n29239_));
  NOR2_X1    g26803(.A1(new_n28051_), .A2(new_n8510_), .ZN(new_n29240_));
  AOI21_X1   g26804(.A1(new_n28595_), .A2(new_n29240_), .B(new_n8511_), .ZN(new_n29241_));
  NOR2_X1    g26805(.A1(new_n28607_), .A2(new_n28269_), .ZN(new_n29242_));
  INV_X1     g26806(.I(new_n29242_), .ZN(new_n29243_));
  AOI21_X1   g26807(.A1(new_n29243_), .A2(new_n29241_), .B(new_n29239_), .ZN(new_n29244_));
  AOI21_X1   g26808(.A1(new_n29236_), .A2(pi0212), .B(po1038), .ZN(new_n29245_));
  NOR3_X1    g26809(.A1(new_n29237_), .A2(pi0212), .A3(new_n8807_), .ZN(new_n29246_));
  OAI21_X1   g26810(.A1(new_n29235_), .A2(new_n8510_), .B(pi0214), .ZN(new_n29247_));
  NOR2_X1    g26811(.A1(new_n28569_), .A2(new_n28048_), .ZN(new_n29248_));
  OAI21_X1   g26812(.A1(new_n29248_), .A2(new_n29247_), .B(new_n29246_), .ZN(new_n29249_));
  NAND2_X1   g26813(.A1(new_n29249_), .A2(new_n29245_), .ZN(new_n29250_));
  OAI21_X1   g26814(.A1(new_n29250_), .A2(new_n29244_), .B(new_n28360_), .ZN(new_n29251_));
  NOR3_X1    g26815(.A1(new_n28909_), .A2(pi0208), .A3(new_n28842_), .ZN(new_n29252_));
  INV_X1     g26816(.I(new_n29252_), .ZN(new_n29253_));
  NOR2_X1    g26817(.A1(new_n29253_), .A2(pi0214), .ZN(new_n29254_));
  NOR3_X1    g26818(.A1(new_n29254_), .A2(pi0212), .A3(pi0219), .ZN(new_n29255_));
  NAND3_X1   g26819(.A1(new_n29253_), .A2(new_n8510_), .A3(new_n28516_), .ZN(new_n29256_));
  NAND2_X1   g26820(.A1(new_n29256_), .A2(pi0214), .ZN(new_n29257_));
  NOR3_X1    g26821(.A1(new_n28863_), .A2(new_n8510_), .A3(new_n28051_), .ZN(new_n29258_));
  OAI21_X1   g26822(.A1(new_n29258_), .A2(new_n29257_), .B(new_n29255_), .ZN(new_n29259_));
  AOI21_X1   g26823(.A1(new_n29253_), .A2(pi0212), .B(po1038), .ZN(new_n29260_));
  NOR3_X1    g26824(.A1(new_n29254_), .A2(pi0212), .A3(new_n8807_), .ZN(new_n29261_));
  NOR3_X1    g26825(.A1(new_n28863_), .A2(pi0211), .A3(new_n28048_), .ZN(new_n29262_));
  OAI21_X1   g26826(.A1(new_n29252_), .A2(new_n8510_), .B(pi0214), .ZN(new_n29263_));
  OAI21_X1   g26827(.A1(new_n29262_), .A2(new_n29263_), .B(new_n29261_), .ZN(new_n29264_));
  NAND3_X1   g26828(.A1(new_n29259_), .A2(new_n29264_), .A3(new_n29260_), .ZN(new_n29265_));
  NAND2_X1   g26829(.A1(new_n29265_), .A2(pi0209), .ZN(new_n29266_));
  AOI21_X1   g26830(.A1(new_n29266_), .A2(new_n29251_), .B(new_n29234_), .ZN(new_n29267_));
  NOR2_X1    g26831(.A1(new_n6643_), .A2(new_n28812_), .ZN(new_n29268_));
  NAND2_X1   g26832(.A1(new_n28810_), .A2(new_n8807_), .ZN(new_n29269_));
  AOI21_X1   g26833(.A1(new_n29268_), .A2(new_n29269_), .B(new_n26198_), .ZN(new_n29270_));
  NOR2_X1    g26834(.A1(new_n29252_), .A2(new_n8510_), .ZN(new_n29271_));
  OAI21_X1   g26835(.A1(new_n29257_), .A2(new_n29271_), .B(new_n29261_), .ZN(new_n29272_));
  NAND3_X1   g26836(.A1(new_n29272_), .A2(pi0209), .A3(new_n29260_), .ZN(new_n29273_));
  INV_X1     g26837(.I(new_n29255_), .ZN(new_n29274_));
  AOI21_X1   g26838(.A1(pi0208), .A2(pi0299), .B(new_n12965_), .ZN(new_n29275_));
  INV_X1     g26839(.I(new_n29275_), .ZN(new_n29276_));
  NOR2_X1    g26840(.A1(new_n28936_), .A2(new_n29276_), .ZN(new_n29277_));
  OAI21_X1   g26841(.A1(new_n28909_), .A2(new_n29277_), .B(pi0211), .ZN(new_n29278_));
  OAI21_X1   g26842(.A1(new_n2628_), .A2(new_n12745_), .B(pi0208), .ZN(new_n29279_));
  NAND3_X1   g26843(.A1(new_n28947_), .A2(new_n28256_), .A3(new_n29279_), .ZN(new_n29280_));
  AOI21_X1   g26844(.A1(new_n28958_), .A2(new_n29280_), .B(new_n8511_), .ZN(new_n29281_));
  AOI21_X1   g26845(.A1(new_n29278_), .A2(new_n29281_), .B(new_n29274_), .ZN(new_n29282_));
  OAI21_X1   g26846(.A1(new_n29273_), .A2(new_n29282_), .B(new_n29270_), .ZN(new_n29283_));
  OAI21_X1   g26847(.A1(new_n29242_), .A2(new_n29247_), .B(new_n29246_), .ZN(new_n29284_));
  NAND3_X1   g26848(.A1(new_n29284_), .A2(new_n28360_), .A3(new_n29245_), .ZN(new_n29285_));
  NAND2_X1   g26849(.A1(new_n28558_), .A2(new_n28097_), .ZN(new_n29286_));
  OAI21_X1   g26850(.A1(new_n29235_), .A2(pi1157), .B(pi0211), .ZN(new_n29287_));
  AOI21_X1   g26851(.A1(new_n29286_), .A2(new_n29275_), .B(new_n29287_), .ZN(new_n29288_));
  NAND3_X1   g26852(.A1(new_n28825_), .A2(pi0299), .A3(pi1158), .ZN(new_n29289_));
  OR2_X2     g26853(.A1(new_n28953_), .A2(new_n28825_), .Z(new_n29290_));
  AOI21_X1   g26854(.A1(new_n29290_), .A2(new_n29289_), .B(pi0211), .ZN(new_n29291_));
  OAI21_X1   g26855(.A1(new_n29291_), .A2(new_n29288_), .B(pi0214), .ZN(new_n29292_));
  AOI21_X1   g26856(.A1(new_n29292_), .A2(new_n29238_), .B(new_n29285_), .ZN(new_n29293_));
  OAI21_X1   g26857(.A1(new_n29283_), .A2(new_n29293_), .B(pi0230), .ZN(new_n29294_));
  OAI22_X1   g26858(.A1(new_n29294_), .A2(new_n29267_), .B1(pi0230), .B2(new_n3476_), .ZN(po0396));
  INV_X1     g26859(.I(pi1148), .ZN(new_n29296_));
  INV_X1     g26860(.I(pi1149), .ZN(new_n29297_));
  INV_X1     g26861(.I(new_n8810_), .ZN(new_n29298_));
  NOR2_X1    g26862(.A1(new_n29298_), .A2(new_n28361_), .ZN(new_n29299_));
  NOR2_X1    g26863(.A1(new_n28794_), .A2(new_n8531_), .ZN(new_n29300_));
  INV_X1     g26864(.I(new_n29300_), .ZN(new_n29301_));
  AOI21_X1   g26865(.A1(pi0199), .A2(pi1145), .B(pi0200), .ZN(new_n29302_));
  NOR2_X1    g26866(.A1(new_n3343_), .A2(pi0199), .ZN(new_n29303_));
  INV_X1     g26867(.I(new_n29303_), .ZN(new_n29304_));
  NAND2_X1   g26868(.A1(new_n29304_), .A2(new_n29302_), .ZN(new_n29305_));
  NAND3_X1   g26869(.A1(new_n29301_), .A2(new_n29305_), .A3(new_n28026_), .ZN(new_n29306_));
  NAND2_X1   g26870(.A1(new_n29306_), .A2(new_n28371_), .ZN(new_n29307_));
  INV_X1     g26871(.I(new_n29302_), .ZN(new_n29308_));
  AOI21_X1   g26872(.A1(new_n29304_), .A2(pi0200), .B(pi0299), .ZN(new_n29309_));
  NAND2_X1   g26873(.A1(new_n29309_), .A2(new_n29308_), .ZN(new_n29310_));
  NAND2_X1   g26874(.A1(new_n29310_), .A2(new_n8524_), .ZN(new_n29311_));
  NAND2_X1   g26875(.A1(new_n29307_), .A2(new_n29311_), .ZN(new_n29312_));
  INV_X1     g26876(.I(new_n29312_), .ZN(new_n29313_));
  AOI21_X1   g26877(.A1(new_n29313_), .A2(new_n6643_), .B(new_n29299_), .ZN(new_n29314_));
  INV_X1     g26878(.I(new_n29299_), .ZN(new_n29315_));
  NOR2_X1    g26879(.A1(new_n2628_), .A2(new_n3343_), .ZN(new_n29316_));
  INV_X1     g26880(.I(new_n29316_), .ZN(new_n29317_));
  INV_X1     g26881(.I(new_n29309_), .ZN(new_n29318_));
  AOI21_X1   g26882(.A1(new_n3512_), .A2(new_n28123_), .B(new_n29318_), .ZN(new_n29319_));
  NAND2_X1   g26883(.A1(new_n29319_), .A2(new_n8521_), .ZN(new_n29320_));
  NAND3_X1   g26884(.A1(new_n29320_), .A2(new_n29306_), .A3(new_n29317_), .ZN(new_n29321_));
  NAND2_X1   g26885(.A1(new_n29321_), .A2(pi0208), .ZN(new_n29322_));
  NOR2_X1    g26886(.A1(new_n29320_), .A2(new_n29308_), .ZN(new_n29323_));
  OAI22_X1   g26887(.A1(new_n29322_), .A2(new_n29323_), .B1(new_n28825_), .B2(new_n29310_), .ZN(new_n29324_));
  NOR3_X1    g26888(.A1(new_n29324_), .A2(new_n25319_), .A3(new_n29315_), .ZN(new_n29325_));
  NOR3_X1    g26889(.A1(new_n29325_), .A2(pi1147), .A3(new_n29314_), .ZN(new_n29326_));
  NOR2_X1    g26890(.A1(new_n8520_), .A2(new_n29153_), .ZN(new_n29327_));
  NOR2_X1    g26891(.A1(new_n28060_), .A2(new_n29327_), .ZN(new_n29328_));
  INV_X1     g26892(.I(new_n29328_), .ZN(new_n29329_));
  OR2_X2     g26893(.A1(new_n29319_), .A2(new_n8523_), .Z(new_n29330_));
  NAND2_X1   g26894(.A1(new_n29330_), .A2(new_n29307_), .ZN(new_n29331_));
  OAI21_X1   g26895(.A1(new_n29331_), .A2(new_n28057_), .B(pi0219), .ZN(new_n29332_));
  NAND2_X1   g26896(.A1(new_n29319_), .A2(new_n28041_), .ZN(new_n29333_));
  NAND2_X1   g26897(.A1(new_n29322_), .A2(new_n29333_), .ZN(new_n29334_));
  NOR2_X1    g26898(.A1(new_n29334_), .A2(pi0299), .ZN(new_n29335_));
  NOR2_X1    g26899(.A1(new_n29335_), .A2(pi0211), .ZN(new_n29336_));
  NAND2_X1   g26900(.A1(new_n29336_), .A2(new_n28430_), .ZN(new_n29337_));
  INV_X1     g26901(.I(new_n29337_), .ZN(new_n29338_));
  OAI21_X1   g26902(.A1(new_n29338_), .A2(new_n29332_), .B(new_n6643_), .ZN(new_n29339_));
  NAND2_X1   g26903(.A1(new_n29336_), .A2(pi0214), .ZN(new_n29340_));
  AOI21_X1   g26904(.A1(new_n29340_), .A2(new_n29331_), .B(pi0212), .ZN(new_n29341_));
  INV_X1     g26905(.I(new_n29331_), .ZN(new_n29342_));
  NOR3_X1    g26906(.A1(new_n29336_), .A2(pi0214), .A3(new_n29342_), .ZN(new_n29343_));
  NOR2_X1    g26907(.A1(new_n29335_), .A2(new_n8510_), .ZN(new_n29344_));
  NAND2_X1   g26908(.A1(new_n29331_), .A2(pi0214), .ZN(new_n29345_));
  NOR2_X1    g26909(.A1(new_n29344_), .A2(new_n29345_), .ZN(new_n29346_));
  NOR3_X1    g26910(.A1(new_n29343_), .A2(new_n29346_), .A3(new_n8509_), .ZN(new_n29347_));
  NOR3_X1    g26911(.A1(new_n29347_), .A2(new_n29341_), .A3(pi0219), .ZN(new_n29348_));
  OAI21_X1   g26912(.A1(new_n29348_), .A2(new_n29339_), .B(new_n29329_), .ZN(new_n29349_));
  AOI21_X1   g26913(.A1(new_n29349_), .A2(pi1147), .B(new_n29326_), .ZN(new_n29350_));
  OAI21_X1   g26914(.A1(new_n29350_), .A2(new_n29297_), .B(new_n29296_), .ZN(new_n29351_));
  NOR2_X1    g26915(.A1(new_n29324_), .A2(pi0299), .ZN(new_n29352_));
  INV_X1     g26916(.I(new_n29352_), .ZN(new_n29353_));
  AOI21_X1   g26917(.A1(new_n29353_), .A2(pi0214), .B(new_n29344_), .ZN(new_n29354_));
  OAI22_X1   g26918(.A1(new_n29354_), .A2(new_n8509_), .B1(new_n8513_), .B2(new_n29335_), .ZN(new_n29355_));
  NOR3_X1    g26919(.A1(new_n29355_), .A2(pi0219), .A3(new_n29342_), .ZN(new_n29356_));
  NOR3_X1    g26920(.A1(new_n29356_), .A2(new_n29339_), .A3(new_n29348_), .ZN(new_n29357_));
  OAI21_X1   g26921(.A1(new_n29357_), .A2(new_n29124_), .B(pi1147), .ZN(new_n29358_));
  NOR2_X1    g26922(.A1(po1038), .A2(pi1147), .ZN(new_n29359_));
  NAND2_X1   g26923(.A1(new_n29313_), .A2(new_n29359_), .ZN(new_n29360_));
  AOI21_X1   g26924(.A1(new_n29358_), .A2(new_n29360_), .B(pi1149), .ZN(new_n29361_));
  OAI21_X1   g26925(.A1(new_n29361_), .A2(new_n29351_), .B(pi0213), .ZN(new_n29362_));
  INV_X1     g26926(.I(pi1147), .ZN(new_n29363_));
  AOI21_X1   g26927(.A1(new_n29298_), .A2(new_n28430_), .B(pi0219), .ZN(new_n29364_));
  NOR2_X1    g26928(.A1(new_n28060_), .A2(new_n29364_), .ZN(new_n29365_));
  NOR2_X1    g26929(.A1(new_n29365_), .A2(new_n29363_), .ZN(new_n29366_));
  OAI21_X1   g26930(.A1(new_n29356_), .A2(new_n29339_), .B(new_n29366_), .ZN(new_n29367_));
  NAND2_X1   g26931(.A1(new_n29313_), .A2(pi0219), .ZN(new_n29368_));
  NOR2_X1    g26932(.A1(new_n29313_), .A2(pi0214), .ZN(new_n29369_));
  INV_X1     g26933(.I(new_n29369_), .ZN(new_n29370_));
  OAI21_X1   g26934(.A1(new_n29353_), .A2(new_n8511_), .B(new_n29370_), .ZN(new_n29371_));
  NAND2_X1   g26935(.A1(new_n29371_), .A2(new_n8509_), .ZN(new_n29372_));
  NOR2_X1    g26936(.A1(new_n29336_), .A2(new_n29345_), .ZN(new_n29373_));
  OAI21_X1   g26937(.A1(new_n29373_), .A2(new_n29352_), .B(pi0212), .ZN(new_n29374_));
  NAND3_X1   g26938(.A1(new_n29372_), .A2(new_n29374_), .A3(new_n8807_), .ZN(new_n29375_));
  AOI21_X1   g26939(.A1(new_n29375_), .A2(new_n29368_), .B(po1038), .ZN(new_n29376_));
  OAI21_X1   g26940(.A1(new_n28430_), .A2(new_n29312_), .B(new_n29356_), .ZN(new_n29377_));
  NAND2_X1   g26941(.A1(new_n29377_), .A2(new_n29376_), .ZN(new_n29378_));
  INV_X1     g26942(.I(new_n29156_), .ZN(new_n29379_));
  AOI21_X1   g26943(.A1(new_n28669_), .A2(pi0211), .B(new_n28261_), .ZN(new_n29380_));
  NOR2_X1    g26944(.A1(new_n29379_), .A2(new_n29380_), .ZN(new_n29381_));
  INV_X1     g26945(.I(new_n29381_), .ZN(new_n29382_));
  NAND3_X1   g26946(.A1(new_n29378_), .A2(new_n29363_), .A3(new_n29382_), .ZN(new_n29383_));
  AND3_X2    g26947(.A1(new_n29383_), .A2(new_n29297_), .A3(new_n29367_), .Z(new_n29384_));
  NOR2_X1    g26948(.A1(new_n8510_), .A2(new_n8807_), .ZN(new_n29385_));
  NOR2_X1    g26949(.A1(new_n6643_), .A2(new_n29385_), .ZN(new_n29386_));
  INV_X1     g26950(.I(new_n29386_), .ZN(new_n29387_));
  NOR2_X1    g26951(.A1(new_n29387_), .A2(new_n28056_), .ZN(new_n29388_));
  NOR3_X1    g26952(.A1(new_n29342_), .A2(pi0219), .A3(new_n28804_), .ZN(new_n29389_));
  OAI21_X1   g26953(.A1(new_n29339_), .A2(new_n29389_), .B(pi1147), .ZN(new_n29390_));
  OAI21_X1   g26954(.A1(new_n29390_), .A2(new_n29388_), .B(pi1149), .ZN(new_n29391_));
  NOR3_X1    g26955(.A1(new_n29376_), .A2(pi1147), .A3(new_n29125_), .ZN(new_n29392_));
  OAI21_X1   g26956(.A1(new_n29392_), .A2(new_n29391_), .B(pi1148), .ZN(new_n29393_));
  NOR2_X1    g26957(.A1(new_n29384_), .A2(new_n29393_), .ZN(new_n29394_));
  NAND2_X1   g26958(.A1(new_n29370_), .A2(new_n8509_), .ZN(new_n29395_));
  NOR2_X1    g26959(.A1(new_n29317_), .A2(new_n8510_), .ZN(new_n29396_));
  NOR2_X1    g26960(.A1(new_n29313_), .A2(new_n29396_), .ZN(new_n29397_));
  OAI21_X1   g26961(.A1(new_n29395_), .A2(new_n29397_), .B(new_n8807_), .ZN(new_n29398_));
  NOR2_X1    g26962(.A1(new_n29370_), .A2(new_n29396_), .ZN(new_n29399_));
  NOR2_X1    g26963(.A1(new_n29399_), .A2(new_n8509_), .ZN(new_n29400_));
  NAND2_X1   g26964(.A1(new_n29324_), .A2(new_n2628_), .ZN(new_n29401_));
  NOR2_X1    g26965(.A1(new_n8510_), .A2(pi1145), .ZN(new_n29402_));
  AOI21_X1   g26966(.A1(new_n8510_), .A2(new_n3343_), .B(new_n29402_), .ZN(new_n29403_));
  INV_X1     g26967(.I(new_n29403_), .ZN(new_n29404_));
  NOR2_X1    g26968(.A1(new_n29404_), .A2(new_n2628_), .ZN(new_n29405_));
  NOR2_X1    g26969(.A1(new_n29405_), .A2(new_n8511_), .ZN(new_n29406_));
  NAND2_X1   g26970(.A1(new_n29401_), .A2(new_n29406_), .ZN(new_n29407_));
  AOI21_X1   g26971(.A1(new_n29407_), .A2(new_n29400_), .B(new_n29398_), .ZN(new_n29408_));
  NOR2_X1    g26972(.A1(new_n29312_), .A2(new_n28430_), .ZN(new_n29409_));
  NOR2_X1    g26973(.A1(new_n29409_), .A2(new_n8807_), .ZN(new_n29410_));
  OAI21_X1   g26974(.A1(new_n29313_), .A2(new_n8510_), .B(new_n28430_), .ZN(new_n29411_));
  AND3_X2    g26975(.A1(new_n29401_), .A2(new_n8510_), .A3(new_n28880_), .Z(new_n29412_));
  OAI21_X1   g26976(.A1(new_n29412_), .A2(new_n29411_), .B(new_n29410_), .ZN(new_n29413_));
  NAND2_X1   g26977(.A1(new_n29413_), .A2(new_n6643_), .ZN(new_n29414_));
  NOR2_X1    g26978(.A1(new_n3512_), .A2(pi0211), .ZN(new_n29415_));
  OAI21_X1   g26979(.A1(new_n8807_), .A2(new_n29415_), .B(po1038), .ZN(new_n29416_));
  NOR2_X1    g26980(.A1(new_n8510_), .A2(new_n3343_), .ZN(new_n29417_));
  AOI22_X1   g26981(.A1(new_n28669_), .A2(new_n29417_), .B1(new_n8809_), .B2(new_n29403_), .ZN(new_n29418_));
  AOI21_X1   g26982(.A1(new_n29008_), .A2(new_n29418_), .B(new_n29416_), .ZN(new_n29419_));
  NOR2_X1    g26983(.A1(new_n29419_), .A2(pi1147), .ZN(new_n29420_));
  OAI21_X1   g26984(.A1(new_n29414_), .A2(new_n29408_), .B(new_n29420_), .ZN(new_n29421_));
  NOR2_X1    g26985(.A1(new_n29396_), .A2(new_n29187_), .ZN(new_n29422_));
  NAND4_X1   g26986(.A1(new_n29322_), .A2(new_n8511_), .A3(new_n29333_), .A4(new_n29422_), .ZN(new_n29423_));
  NAND2_X1   g26987(.A1(new_n29423_), .A2(pi0212), .ZN(new_n29424_));
  INV_X1     g26988(.I(new_n29406_), .ZN(new_n29425_));
  OAI22_X1   g26989(.A1(new_n29335_), .A2(new_n8513_), .B1(new_n29334_), .B2(new_n29425_), .ZN(new_n29426_));
  NAND2_X1   g26990(.A1(new_n29344_), .A2(new_n28877_), .ZN(new_n29427_));
  AOI21_X1   g26991(.A1(new_n29427_), .A2(new_n29426_), .B(new_n29424_), .ZN(new_n29428_));
  NOR3_X1    g26992(.A1(new_n29428_), .A2(new_n29341_), .A3(new_n29398_), .ZN(new_n29429_));
  NOR2_X1    g26993(.A1(new_n29337_), .A2(new_n28876_), .ZN(new_n29430_));
  OAI21_X1   g26994(.A1(new_n29430_), .A2(new_n29332_), .B(new_n6643_), .ZN(new_n29431_));
  NOR2_X1    g26995(.A1(new_n29315_), .A2(new_n6643_), .ZN(new_n29432_));
  NOR3_X1    g26996(.A1(new_n29419_), .A2(new_n29363_), .A3(new_n29432_), .ZN(new_n29433_));
  OAI21_X1   g26997(.A1(new_n29429_), .A2(new_n29431_), .B(new_n29433_), .ZN(new_n29434_));
  NAND2_X1   g26998(.A1(new_n29434_), .A2(new_n29421_), .ZN(new_n29435_));
  OAI22_X1   g26999(.A1(new_n29394_), .A2(new_n29362_), .B1(pi0213), .B2(new_n29435_), .ZN(new_n29436_));
  INV_X1     g27000(.I(new_n29089_), .ZN(new_n29437_));
  NAND2_X1   g27001(.A1(new_n29078_), .A2(new_n8511_), .ZN(new_n29438_));
  NAND2_X1   g27002(.A1(new_n29438_), .A2(new_n8509_), .ZN(new_n29439_));
  NOR2_X1    g27003(.A1(new_n29437_), .A2(new_n8511_), .ZN(new_n29440_));
  NOR2_X1    g27004(.A1(new_n29440_), .A2(new_n29439_), .ZN(new_n29441_));
  NOR2_X1    g27005(.A1(new_n29441_), .A2(pi0219), .ZN(new_n29442_));
  INV_X1     g27006(.I(new_n29442_), .ZN(new_n29443_));
  INV_X1     g27007(.I(new_n29086_), .ZN(new_n29444_));
  AOI21_X1   g27008(.A1(new_n29077_), .A2(new_n8510_), .B(new_n8511_), .ZN(new_n29445_));
  INV_X1     g27009(.I(new_n29445_), .ZN(new_n29446_));
  AOI21_X1   g27010(.A1(new_n29444_), .A2(pi0211), .B(new_n29446_), .ZN(new_n29447_));
  NOR2_X1    g27011(.A1(new_n29447_), .A2(new_n8509_), .ZN(new_n29448_));
  AOI21_X1   g27012(.A1(new_n29437_), .A2(new_n29448_), .B(new_n29443_), .ZN(new_n29449_));
  INV_X1     g27013(.I(new_n29449_), .ZN(new_n29450_));
  NOR2_X1    g27014(.A1(new_n29447_), .A2(new_n8811_), .ZN(new_n29451_));
  NOR2_X1    g27015(.A1(new_n29450_), .A2(new_n29451_), .ZN(new_n29452_));
  INV_X1     g27016(.I(new_n29441_), .ZN(new_n29453_));
  AOI21_X1   g27017(.A1(new_n29437_), .A2(pi0212), .B(new_n8807_), .ZN(new_n29454_));
  AOI21_X1   g27018(.A1(new_n29453_), .A2(new_n29454_), .B(po1038), .ZN(new_n29455_));
  INV_X1     g27019(.I(new_n29455_), .ZN(new_n29456_));
  NOR2_X1    g27020(.A1(new_n29452_), .A2(new_n29456_), .ZN(new_n29457_));
  NOR2_X1    g27021(.A1(new_n29457_), .A2(new_n29328_), .ZN(new_n29458_));
  NOR2_X1    g27022(.A1(new_n12618_), .A2(pi0219), .ZN(new_n29459_));
  INV_X1     g27023(.I(new_n29459_), .ZN(new_n29460_));
  NOR2_X1    g27024(.A1(new_n29460_), .A2(new_n29154_), .ZN(new_n29461_));
  NAND2_X1   g27025(.A1(new_n12618_), .A2(new_n29042_), .ZN(new_n29462_));
  INV_X1     g27026(.I(new_n29462_), .ZN(new_n29463_));
  NOR2_X1    g27027(.A1(new_n29461_), .A2(new_n29463_), .ZN(new_n29464_));
  INV_X1     g27028(.I(new_n29464_), .ZN(new_n29465_));
  NAND2_X1   g27029(.A1(new_n29465_), .A2(new_n29363_), .ZN(new_n29466_));
  OAI21_X1   g27030(.A1(new_n29458_), .A2(new_n29363_), .B(new_n29466_), .ZN(new_n29467_));
  OAI21_X1   g27031(.A1(new_n8531_), .A2(new_n8521_), .B(new_n28151_), .ZN(new_n29468_));
  AOI21_X1   g27032(.A1(new_n29468_), .A2(pi0208), .B(pi0199), .ZN(new_n29469_));
  NOR2_X1    g27033(.A1(new_n29053_), .A2(new_n29469_), .ZN(new_n29470_));
  NOR2_X1    g27034(.A1(new_n29470_), .A2(pi0299), .ZN(new_n29471_));
  INV_X1     g27035(.I(new_n29044_), .ZN(new_n29472_));
  AOI21_X1   g27036(.A1(new_n29062_), .A2(new_n29188_), .B(new_n8509_), .ZN(new_n29473_));
  INV_X1     g27037(.I(new_n29473_), .ZN(new_n29474_));
  AOI21_X1   g27038(.A1(new_n29472_), .A2(new_n29218_), .B(new_n29474_), .ZN(new_n29475_));
  AOI21_X1   g27039(.A1(pi0214), .A2(new_n29187_), .B(new_n29054_), .ZN(new_n29476_));
  INV_X1     g27040(.I(new_n29476_), .ZN(new_n29477_));
  AOI21_X1   g27041(.A1(new_n29477_), .A2(new_n8509_), .B(pi0219), .ZN(new_n29478_));
  INV_X1     g27042(.I(new_n29478_), .ZN(new_n29479_));
  NOR2_X1    g27043(.A1(new_n29475_), .A2(new_n29479_), .ZN(new_n29480_));
  NOR2_X1    g27044(.A1(new_n29053_), .A2(po1038), .ZN(new_n29481_));
  INV_X1     g27045(.I(new_n29481_), .ZN(new_n29482_));
  NOR2_X1    g27046(.A1(po1038), .A2(new_n28058_), .ZN(new_n29483_));
  INV_X1     g27047(.I(new_n29483_), .ZN(new_n29484_));
  AOI21_X1   g27048(.A1(pi0219), .A2(new_n29188_), .B(new_n29484_), .ZN(new_n29485_));
  INV_X1     g27049(.I(new_n29485_), .ZN(new_n29486_));
  AOI21_X1   g27050(.A1(new_n29482_), .A2(new_n29486_), .B(new_n29480_), .ZN(new_n29487_));
  INV_X1     g27051(.I(new_n29487_), .ZN(new_n29488_));
  NOR2_X1    g27052(.A1(new_n29488_), .A2(new_n29471_), .ZN(new_n29489_));
  INV_X1     g27053(.I(new_n29489_), .ZN(new_n29490_));
  INV_X1     g27054(.I(new_n29471_), .ZN(new_n29491_));
  AOI21_X1   g27055(.A1(new_n29044_), .A2(new_n8511_), .B(new_n8509_), .ZN(new_n29492_));
  NOR2_X1    g27056(.A1(new_n8513_), .A2(new_n2628_), .ZN(new_n29493_));
  NOR3_X1    g27057(.A1(new_n29054_), .A2(pi0212), .A3(new_n29493_), .ZN(new_n29494_));
  AOI21_X1   g27058(.A1(new_n29476_), .A2(new_n29492_), .B(new_n29494_), .ZN(new_n29495_));
  AOI21_X1   g27059(.A1(new_n29495_), .A2(new_n29491_), .B(pi0219), .ZN(new_n29496_));
  AOI21_X1   g27060(.A1(new_n8510_), .A2(new_n29496_), .B(new_n29490_), .ZN(new_n29497_));
  NOR2_X1    g27061(.A1(new_n29497_), .A2(new_n29124_), .ZN(new_n29498_));
  NOR3_X1    g27062(.A1(new_n29498_), .A2(new_n29363_), .A3(pi1149), .ZN(new_n29499_));
  AOI21_X1   g27063(.A1(new_n29467_), .A2(pi1149), .B(new_n29499_), .ZN(new_n29500_));
  AOI22_X1   g27064(.A1(new_n28372_), .A2(new_n28114_), .B1(new_n8523_), .B2(new_n8781_), .ZN(new_n29501_));
  INV_X1     g27065(.I(new_n29501_), .ZN(new_n29502_));
  NAND2_X1   g27066(.A1(new_n29502_), .A2(new_n29021_), .ZN(new_n29503_));
  INV_X1     g27067(.I(new_n29503_), .ZN(new_n29504_));
  NOR2_X1    g27068(.A1(new_n29504_), .A2(new_n29493_), .ZN(new_n29505_));
  OAI21_X1   g27069(.A1(new_n29505_), .A2(pi0212), .B(new_n8807_), .ZN(new_n29506_));
  NOR2_X1    g27070(.A1(new_n29504_), .A2(new_n29044_), .ZN(new_n29507_));
  NOR2_X1    g27071(.A1(new_n29502_), .A2(pi0299), .ZN(new_n29508_));
  NOR2_X1    g27072(.A1(new_n29508_), .A2(new_n8511_), .ZN(new_n29509_));
  INV_X1     g27073(.I(new_n29509_), .ZN(new_n29510_));
  AOI21_X1   g27074(.A1(new_n29510_), .A2(new_n29507_), .B(new_n8509_), .ZN(new_n29511_));
  INV_X1     g27075(.I(new_n29511_), .ZN(new_n29512_));
  OAI21_X1   g27076(.A1(new_n29503_), .A2(pi0214), .B(new_n8509_), .ZN(new_n29513_));
  NOR2_X1    g27077(.A1(new_n29508_), .A2(pi0211), .ZN(new_n29514_));
  NOR2_X1    g27078(.A1(new_n29514_), .A2(new_n29504_), .ZN(new_n29515_));
  INV_X1     g27079(.I(new_n29515_), .ZN(new_n29516_));
  AOI21_X1   g27080(.A1(new_n29516_), .A2(pi0214), .B(new_n8509_), .ZN(new_n29517_));
  OAI21_X1   g27081(.A1(pi0214), .A2(new_n29508_), .B(new_n29517_), .ZN(new_n29518_));
  OAI21_X1   g27082(.A1(new_n29509_), .A2(new_n29513_), .B(new_n29518_), .ZN(new_n29519_));
  NOR2_X1    g27083(.A1(new_n29519_), .A2(new_n29512_), .ZN(new_n29520_));
  NOR2_X1    g27084(.A1(new_n29520_), .A2(new_n29506_), .ZN(new_n29521_));
  NAND2_X1   g27085(.A1(new_n29503_), .A2(pi0219), .ZN(new_n29522_));
  NAND2_X1   g27086(.A1(new_n29522_), .A2(new_n6643_), .ZN(new_n29523_));
  NOR2_X1    g27087(.A1(new_n29521_), .A2(new_n29523_), .ZN(new_n29524_));
  NOR2_X1    g27088(.A1(new_n29524_), .A2(new_n29381_), .ZN(new_n29525_));
  NOR2_X1    g27089(.A1(new_n29525_), .A2(pi1147), .ZN(new_n29526_));
  INV_X1     g27090(.I(new_n28804_), .ZN(new_n29527_));
  NOR2_X1    g27091(.A1(new_n29484_), .A2(new_n29527_), .ZN(new_n29528_));
  INV_X1     g27092(.I(new_n29528_), .ZN(new_n29529_));
  AOI21_X1   g27093(.A1(new_n29529_), .A2(new_n28060_), .B(new_n29364_), .ZN(new_n29530_));
  NOR2_X1    g27094(.A1(new_n29530_), .A2(new_n29481_), .ZN(new_n29531_));
  NOR2_X1    g27095(.A1(new_n29531_), .A2(new_n29363_), .ZN(new_n29532_));
  OAI21_X1   g27096(.A1(new_n29526_), .A2(new_n29532_), .B(new_n29297_), .ZN(new_n29533_));
  NOR2_X1    g27097(.A1(new_n29010_), .A2(po1038), .ZN(new_n29534_));
  NOR2_X1    g27098(.A1(new_n29184_), .A2(new_n29534_), .ZN(new_n29535_));
  NOR2_X1    g27099(.A1(new_n28825_), .A2(new_n9183_), .ZN(new_n29536_));
  NOR2_X1    g27100(.A1(new_n29024_), .A2(pi0299), .ZN(new_n29537_));
  INV_X1     g27101(.I(new_n29537_), .ZN(new_n29538_));
  NOR2_X1    g27102(.A1(new_n29538_), .A2(new_n29536_), .ZN(new_n29539_));
  INV_X1     g27103(.I(new_n29539_), .ZN(new_n29540_));
  NOR2_X1    g27104(.A1(new_n29009_), .A2(pi0214), .ZN(new_n29541_));
  NOR2_X1    g27105(.A1(new_n29541_), .A2(pi0212), .ZN(new_n29542_));
  OAI21_X1   g27106(.A1(new_n29540_), .A2(new_n8511_), .B(new_n29542_), .ZN(new_n29543_));
  NAND2_X1   g27107(.A1(new_n29543_), .A2(new_n8807_), .ZN(new_n29544_));
  NOR2_X1    g27108(.A1(new_n29539_), .A2(pi0211), .ZN(new_n29545_));
  NOR2_X1    g27109(.A1(new_n29010_), .A2(new_n8510_), .ZN(new_n29546_));
  NOR3_X1    g27110(.A1(new_n29545_), .A2(new_n8511_), .A3(new_n29546_), .ZN(new_n29547_));
  NOR2_X1    g27111(.A1(new_n29547_), .A2(new_n8509_), .ZN(new_n29548_));
  AOI21_X1   g27112(.A1(new_n29548_), .A2(new_n29540_), .B(new_n29544_), .ZN(new_n29549_));
  NOR2_X1    g27113(.A1(new_n29549_), .A2(new_n29535_), .ZN(new_n29550_));
  NOR2_X1    g27114(.A1(new_n29550_), .A2(new_n29125_), .ZN(new_n29551_));
  NOR2_X1    g27115(.A1(new_n28448_), .A2(new_n28620_), .ZN(new_n29552_));
  INV_X1     g27116(.I(new_n29552_), .ZN(new_n29553_));
  NOR2_X1    g27117(.A1(new_n29388_), .A2(new_n29528_), .ZN(new_n29554_));
  OAI21_X1   g27118(.A1(po1038), .A2(new_n29553_), .B(new_n29554_), .ZN(new_n29555_));
  NAND2_X1   g27119(.A1(new_n29555_), .A2(pi1147), .ZN(new_n29556_));
  OAI21_X1   g27120(.A1(new_n29551_), .A2(pi1147), .B(new_n29556_), .ZN(new_n29557_));
  AOI21_X1   g27121(.A1(new_n29557_), .A2(pi1149), .B(new_n29296_), .ZN(new_n29558_));
  AOI22_X1   g27122(.A1(new_n29500_), .A2(new_n29296_), .B1(new_n29533_), .B2(new_n29558_), .ZN(new_n29559_));
  INV_X1     g27123(.I(new_n29433_), .ZN(new_n29560_));
  INV_X1     g27124(.I(new_n29405_), .ZN(new_n29561_));
  AOI21_X1   g27125(.A1(new_n29053_), .A2(new_n29561_), .B(new_n8811_), .ZN(new_n29562_));
  AOI21_X1   g27126(.A1(new_n29054_), .A2(new_n28056_), .B(pi0219), .ZN(new_n29563_));
  INV_X1     g27127(.I(new_n29563_), .ZN(new_n29564_));
  AOI21_X1   g27128(.A1(new_n29053_), .A2(new_n29422_), .B(new_n28212_), .ZN(new_n29565_));
  OR3_X2     g27129(.A1(new_n29564_), .A2(new_n29562_), .A3(new_n29565_), .Z(new_n29566_));
  NOR2_X1    g27130(.A1(new_n28880_), .A2(pi0211), .ZN(new_n29567_));
  OAI21_X1   g27131(.A1(new_n8807_), .A2(new_n29567_), .B(new_n29483_), .ZN(new_n29568_));
  NAND2_X1   g27132(.A1(new_n29482_), .A2(new_n29568_), .ZN(new_n29569_));
  AOI21_X1   g27133(.A1(new_n29566_), .A2(new_n29569_), .B(new_n29560_), .ZN(new_n29570_));
  INV_X1     g27134(.I(new_n29420_), .ZN(new_n29571_));
  NOR2_X1    g27135(.A1(new_n29418_), .A2(new_n2628_), .ZN(new_n29572_));
  NAND2_X1   g27136(.A1(new_n29572_), .A2(new_n26397_), .ZN(new_n29573_));
  OAI21_X1   g27137(.A1(new_n8807_), .A2(new_n29568_), .B(new_n29573_), .ZN(new_n29574_));
  NOR2_X1    g27138(.A1(new_n29503_), .A2(po1038), .ZN(new_n29575_));
  NOR3_X1    g27139(.A1(new_n29571_), .A2(new_n29574_), .A3(new_n29575_), .ZN(new_n29576_));
  NOR3_X1    g27140(.A1(new_n29570_), .A2(new_n29296_), .A3(new_n29576_), .ZN(new_n29577_));
  NOR2_X1    g27141(.A1(new_n29571_), .A2(new_n29574_), .ZN(new_n29578_));
  AOI21_X1   g27142(.A1(new_n3343_), .A2(new_n29044_), .B(new_n28212_), .ZN(new_n29579_));
  OAI21_X1   g27143(.A1(new_n29562_), .A2(new_n29579_), .B(new_n8807_), .ZN(new_n29580_));
  NOR3_X1    g27144(.A1(new_n29527_), .A2(new_n3512_), .A3(new_n28044_), .ZN(new_n29581_));
  AOI21_X1   g27145(.A1(new_n29470_), .A2(new_n28361_), .B(new_n29581_), .ZN(new_n29582_));
  OAI21_X1   g27146(.A1(new_n29580_), .A2(new_n29471_), .B(new_n29582_), .ZN(new_n29583_));
  AOI21_X1   g27147(.A1(new_n29583_), .A2(new_n6643_), .B(new_n29560_), .ZN(new_n29584_));
  NOR3_X1    g27148(.A1(new_n29584_), .A2(pi1148), .A3(new_n29578_), .ZN(new_n29585_));
  NOR3_X1    g27149(.A1(new_n29577_), .A2(pi1149), .A3(new_n29585_), .ZN(new_n29586_));
  NOR2_X1    g27150(.A1(new_n28825_), .A2(pi0200), .ZN(new_n29587_));
  OAI21_X1   g27151(.A1(new_n29084_), .A2(new_n29587_), .B(new_n2628_), .ZN(new_n29588_));
  NAND2_X1   g27152(.A1(new_n29588_), .A2(new_n29406_), .ZN(new_n29589_));
  NAND2_X1   g27153(.A1(new_n29589_), .A2(pi0212), .ZN(new_n29590_));
  AOI21_X1   g27154(.A1(new_n29588_), .A2(new_n29317_), .B(new_n8510_), .ZN(new_n29591_));
  NOR2_X1    g27155(.A1(new_n29591_), .A2(new_n29087_), .ZN(new_n29592_));
  AOI21_X1   g27156(.A1(new_n29592_), .A2(new_n8511_), .B(new_n29590_), .ZN(new_n29593_));
  NOR3_X1    g27157(.A1(new_n29591_), .A2(new_n8511_), .A3(new_n29087_), .ZN(new_n29594_));
  NOR2_X1    g27158(.A1(new_n29594_), .A2(new_n29439_), .ZN(new_n29595_));
  NOR3_X1    g27159(.A1(new_n29593_), .A2(new_n29595_), .A3(pi0219), .ZN(new_n29596_));
  INV_X1     g27160(.I(new_n29568_), .ZN(new_n29597_));
  NOR2_X1    g27161(.A1(new_n29077_), .A2(new_n8807_), .ZN(new_n29598_));
  NOR2_X1    g27162(.A1(new_n29598_), .A2(po1038), .ZN(new_n29599_));
  NOR2_X1    g27163(.A1(new_n29599_), .A2(new_n29597_), .ZN(new_n29600_));
  OAI21_X1   g27164(.A1(new_n29596_), .A2(new_n29600_), .B(new_n29433_), .ZN(new_n29601_));
  AOI21_X1   g27165(.A1(new_n29578_), .A2(new_n29462_), .B(pi1148), .ZN(new_n29602_));
  AOI21_X1   g27166(.A1(new_n29553_), .A2(pi0219), .B(po1038), .ZN(new_n29603_));
  INV_X1     g27167(.I(new_n29603_), .ZN(new_n29604_));
  NOR2_X1    g27168(.A1(new_n8511_), .A2(new_n2628_), .ZN(new_n29605_));
  INV_X1     g27169(.I(new_n29605_), .ZN(new_n29606_));
  AOI21_X1   g27170(.A1(new_n29553_), .A2(new_n29606_), .B(pi0212), .ZN(new_n29607_));
  INV_X1     g27171(.I(new_n29607_), .ZN(new_n29608_));
  NOR2_X1    g27172(.A1(new_n29552_), .A2(new_n8510_), .ZN(new_n29609_));
  NOR2_X1    g27173(.A1(new_n29608_), .A2(new_n29609_), .ZN(new_n29610_));
  INV_X1     g27174(.I(new_n29610_), .ZN(new_n29611_));
  AOI21_X1   g27175(.A1(new_n29553_), .A2(new_n2628_), .B(new_n8509_), .ZN(new_n29612_));
  INV_X1     g27176(.I(new_n28818_), .ZN(new_n29613_));
  NOR2_X1    g27177(.A1(new_n29613_), .A2(new_n28267_), .ZN(new_n29614_));
  INV_X1     g27178(.I(new_n29614_), .ZN(new_n29615_));
  AOI21_X1   g27179(.A1(new_n29612_), .A2(new_n29615_), .B(pi0219), .ZN(new_n29616_));
  AOI21_X1   g27180(.A1(new_n29611_), .A2(new_n29616_), .B(new_n29604_), .ZN(new_n29617_));
  INV_X1     g27181(.I(new_n29574_), .ZN(new_n29618_));
  NAND2_X1   g27182(.A1(new_n29618_), .A2(new_n29433_), .ZN(new_n29619_));
  OAI21_X1   g27183(.A1(new_n29617_), .A2(new_n29619_), .B(pi1148), .ZN(new_n29620_));
  AOI21_X1   g27184(.A1(new_n29009_), .A2(new_n28503_), .B(new_n8807_), .ZN(new_n29621_));
  OAI21_X1   g27185(.A1(new_n29539_), .A2(new_n28503_), .B(new_n29621_), .ZN(new_n29622_));
  NAND2_X1   g27186(.A1(new_n29622_), .A2(new_n6643_), .ZN(new_n29623_));
  OAI21_X1   g27187(.A1(new_n29623_), .A2(new_n9183_), .B(new_n29568_), .ZN(new_n29624_));
  NOR2_X1    g27188(.A1(new_n29539_), .A2(new_n8509_), .ZN(new_n29625_));
  NOR2_X1    g27189(.A1(new_n29404_), .A2(new_n8511_), .ZN(new_n29626_));
  INV_X1     g27190(.I(new_n29417_), .ZN(new_n29627_));
  OAI21_X1   g27191(.A1(pi0214), .A2(new_n29627_), .B(new_n29010_), .ZN(new_n29628_));
  OAI21_X1   g27192(.A1(new_n29626_), .A2(new_n29628_), .B(new_n29625_), .ZN(new_n29629_));
  OAI21_X1   g27193(.A1(new_n29009_), .A2(new_n29396_), .B(new_n29542_), .ZN(new_n29630_));
  NAND3_X1   g27194(.A1(new_n29629_), .A2(new_n29630_), .A3(new_n8807_), .ZN(new_n29631_));
  AOI21_X1   g27195(.A1(new_n29631_), .A2(new_n29624_), .B(new_n29571_), .ZN(new_n29632_));
  OAI21_X1   g27196(.A1(new_n29620_), .A2(new_n29632_), .B(pi1149), .ZN(new_n29633_));
  AOI21_X1   g27197(.A1(new_n29601_), .A2(new_n29602_), .B(new_n29633_), .ZN(new_n29634_));
  OAI21_X1   g27198(.A1(new_n29634_), .A2(new_n29586_), .B(new_n26198_), .ZN(new_n29635_));
  OAI21_X1   g27199(.A1(new_n29559_), .A2(new_n26198_), .B(new_n29635_), .ZN(new_n29636_));
  AOI21_X1   g27200(.A1(new_n29636_), .A2(pi0209), .B(new_n27999_), .ZN(new_n29637_));
  OAI21_X1   g27201(.A1(new_n29436_), .A2(pi0209), .B(new_n29637_), .ZN(new_n29638_));
  OAI21_X1   g27202(.A1(pi0230), .A2(new_n4587_), .B(new_n29638_), .ZN(po0397));
  NOR2_X1    g27203(.A1(new_n29035_), .A2(pi1150), .ZN(new_n29640_));
  AOI21_X1   g27204(.A1(new_n29465_), .A2(new_n29640_), .B(pi1149), .ZN(new_n29641_));
  INV_X1     g27205(.I(new_n29525_), .ZN(new_n29642_));
  NOR2_X1    g27206(.A1(new_n29642_), .A2(pi1151), .ZN(new_n29643_));
  INV_X1     g27207(.I(new_n29643_), .ZN(new_n29644_));
  NOR2_X1    g27208(.A1(new_n29125_), .A2(new_n29035_), .ZN(new_n29645_));
  INV_X1     g27209(.I(new_n29645_), .ZN(new_n29646_));
  NOR2_X1    g27210(.A1(new_n29550_), .A2(new_n29646_), .ZN(new_n29647_));
  INV_X1     g27211(.I(new_n29647_), .ZN(new_n29648_));
  NAND3_X1   g27212(.A1(new_n29644_), .A2(pi1150), .A3(new_n29648_), .ZN(new_n29649_));
  INV_X1     g27213(.I(pi1150), .ZN(new_n29650_));
  NOR2_X1    g27214(.A1(new_n29328_), .A2(new_n29035_), .ZN(new_n29651_));
  INV_X1     g27215(.I(new_n29651_), .ZN(new_n29652_));
  NOR2_X1    g27216(.A1(new_n29457_), .A2(new_n29652_), .ZN(new_n29653_));
  INV_X1     g27217(.I(new_n29653_), .ZN(new_n29654_));
  NOR2_X1    g27218(.A1(new_n29124_), .A2(pi1151), .ZN(new_n29655_));
  INV_X1     g27219(.I(new_n29655_), .ZN(new_n29656_));
  OR2_X2     g27220(.A1(new_n29497_), .A2(new_n29656_), .Z(new_n29657_));
  NAND3_X1   g27221(.A1(new_n29654_), .A2(new_n29657_), .A3(new_n29650_), .ZN(new_n29658_));
  AOI21_X1   g27222(.A1(new_n29531_), .A2(new_n29035_), .B(new_n29650_), .ZN(new_n29659_));
  NOR2_X1    g27223(.A1(new_n29553_), .A2(po1038), .ZN(new_n29660_));
  NOR2_X1    g27224(.A1(new_n29528_), .A2(new_n29660_), .ZN(new_n29661_));
  INV_X1     g27225(.I(new_n29661_), .ZN(new_n29662_));
  NOR2_X1    g27226(.A1(new_n29388_), .A2(new_n29035_), .ZN(new_n29663_));
  INV_X1     g27227(.I(new_n29663_), .ZN(new_n29664_));
  NOR2_X1    g27228(.A1(new_n29664_), .A2(new_n29662_), .ZN(new_n29665_));
  INV_X1     g27229(.I(new_n29665_), .ZN(new_n29666_));
  AOI21_X1   g27230(.A1(new_n29666_), .A2(new_n29659_), .B(new_n29297_), .ZN(new_n29667_));
  AOI22_X1   g27231(.A1(new_n29649_), .A2(new_n29641_), .B1(new_n29658_), .B2(new_n29667_), .ZN(new_n29668_));
  OR2_X2     g27232(.A1(new_n29668_), .A2(pi0213), .Z(new_n29669_));
  AOI21_X1   g27233(.A1(new_n29053_), .A2(new_n29188_), .B(new_n8811_), .ZN(new_n29670_));
  INV_X1     g27234(.I(new_n28969_), .ZN(new_n29671_));
  NOR2_X1    g27235(.A1(new_n29053_), .A2(pi0299), .ZN(new_n29672_));
  AOI21_X1   g27236(.A1(pi0299), .A2(new_n29671_), .B(new_n29672_), .ZN(new_n29673_));
  NOR2_X1    g27237(.A1(new_n29673_), .A2(new_n28066_), .ZN(new_n29674_));
  NOR3_X1    g27238(.A1(new_n29674_), .A2(new_n29564_), .A3(new_n29670_), .ZN(new_n29675_));
  NOR2_X1    g27239(.A1(new_n29055_), .A2(po1038), .ZN(new_n29676_));
  INV_X1     g27240(.I(new_n29676_), .ZN(new_n29677_));
  OAI21_X1   g27241(.A1(new_n29675_), .A2(new_n29677_), .B(new_n29146_), .ZN(new_n29678_));
  NOR2_X1    g27242(.A1(new_n29552_), .A2(pi0219), .ZN(new_n29679_));
  NAND3_X1   g27243(.A1(new_n29679_), .A2(new_n8510_), .A3(new_n29615_), .ZN(new_n29680_));
  NAND2_X1   g27244(.A1(new_n29662_), .A2(new_n29680_), .ZN(new_n29681_));
  NOR2_X1    g27245(.A1(new_n8513_), .A2(new_n29613_), .ZN(new_n29682_));
  NOR2_X1    g27246(.A1(new_n29682_), .A2(pi0219), .ZN(new_n29683_));
  NOR2_X1    g27247(.A1(new_n29486_), .A2(new_n29683_), .ZN(new_n29684_));
  NOR2_X1    g27248(.A1(new_n29617_), .A2(new_n29684_), .ZN(new_n29685_));
  INV_X1     g27249(.I(new_n29685_), .ZN(new_n29686_));
  NAND3_X1   g27250(.A1(new_n29679_), .A2(new_n12841_), .A3(new_n29615_), .ZN(new_n29687_));
  NAND2_X1   g27251(.A1(new_n29686_), .A2(new_n29687_), .ZN(new_n29688_));
  NAND3_X1   g27252(.A1(new_n29688_), .A2(new_n29129_), .A3(new_n29681_), .ZN(new_n29689_));
  NAND3_X1   g27253(.A1(new_n29689_), .A2(pi1152), .A3(new_n29678_), .ZN(new_n29690_));
  INV_X1     g27254(.I(new_n29157_), .ZN(new_n29691_));
  NOR2_X1    g27255(.A1(new_n29154_), .A2(new_n28045_), .ZN(new_n29692_));
  INV_X1     g27256(.I(new_n29692_), .ZN(new_n29693_));
  NOR2_X1    g27257(.A1(new_n29693_), .A2(new_n12841_), .ZN(new_n29694_));
  OAI21_X1   g27258(.A1(new_n29691_), .A2(new_n29694_), .B(new_n28422_), .ZN(new_n29695_));
  OAI21_X1   g27259(.A1(new_n29481_), .A2(pi1151), .B(new_n28422_), .ZN(new_n29696_));
  AOI22_X1   g27260(.A1(new_n29688_), .A2(new_n29166_), .B1(new_n29695_), .B2(new_n29696_), .ZN(new_n29697_));
  NOR2_X1    g27261(.A1(new_n29697_), .A2(new_n29650_), .ZN(new_n29698_));
  AOI21_X1   g27262(.A1(new_n29698_), .A2(new_n29690_), .B(new_n29297_), .ZN(new_n29699_));
  NOR3_X1    g27263(.A1(new_n29086_), .A2(pi0211), .A3(new_n28338_), .ZN(new_n29700_));
  NOR3_X1    g27264(.A1(new_n29451_), .A2(new_n29088_), .A3(new_n29700_), .ZN(new_n29701_));
  AOI21_X1   g27265(.A1(new_n8509_), .A2(new_n29438_), .B(new_n29448_), .ZN(new_n29702_));
  OAI21_X1   g27266(.A1(new_n29702_), .A2(new_n29701_), .B(new_n8807_), .ZN(new_n29703_));
  NAND2_X1   g27267(.A1(new_n29455_), .A2(new_n29703_), .ZN(new_n29704_));
  NOR2_X1    g27268(.A1(new_n29671_), .A2(new_n2628_), .ZN(new_n29705_));
  INV_X1     g27269(.I(new_n29470_), .ZN(new_n29706_));
  AOI21_X1   g27270(.A1(new_n29706_), .A2(new_n29693_), .B(po1038), .ZN(new_n29707_));
  INV_X1     g27271(.I(new_n29707_), .ZN(new_n29708_));
  OAI21_X1   g27272(.A1(new_n29708_), .A2(new_n29705_), .B(new_n29157_), .ZN(new_n29709_));
  NAND2_X1   g27273(.A1(new_n29709_), .A2(new_n28422_), .ZN(new_n29710_));
  AOI21_X1   g27274(.A1(new_n29704_), .A2(new_n29166_), .B(new_n29710_), .ZN(new_n29711_));
  NOR2_X1    g27275(.A1(new_n29470_), .A2(new_n28804_), .ZN(new_n29712_));
  AOI21_X1   g27276(.A1(new_n28126_), .A2(new_n29127_), .B(new_n29712_), .ZN(new_n29713_));
  NOR2_X1    g27277(.A1(new_n29713_), .A2(pi0219), .ZN(new_n29714_));
  OAI21_X1   g27278(.A1(new_n29470_), .A2(new_n8807_), .B(new_n6643_), .ZN(new_n29715_));
  OAI21_X1   g27279(.A1(new_n29714_), .A2(new_n29715_), .B(new_n29146_), .ZN(new_n29716_));
  NAND2_X1   g27280(.A1(new_n29716_), .A2(pi1152), .ZN(new_n29717_));
  INV_X1     g27281(.I(new_n29129_), .ZN(new_n29718_));
  INV_X1     g27282(.I(new_n29447_), .ZN(new_n29719_));
  NAND2_X1   g27283(.A1(new_n29719_), .A2(new_n29438_), .ZN(new_n29720_));
  NAND4_X1   g27284(.A1(new_n29720_), .A2(new_n29091_), .A3(new_n8807_), .A4(new_n29615_), .ZN(new_n29721_));
  AOI21_X1   g27285(.A1(new_n29455_), .A2(new_n29721_), .B(new_n29718_), .ZN(new_n29722_));
  OAI21_X1   g27286(.A1(new_n29722_), .A2(new_n29717_), .B(new_n29650_), .ZN(new_n29723_));
  OAI21_X1   g27287(.A1(new_n29723_), .A2(new_n29711_), .B(new_n29699_), .ZN(new_n29724_));
  AOI21_X1   g27288(.A1(new_n29048_), .A2(pi0219), .B(po1038), .ZN(new_n29725_));
  INV_X1     g27289(.I(new_n29725_), .ZN(new_n29726_));
  OR2_X2     g27290(.A1(new_n29183_), .A2(new_n29726_), .Z(new_n29727_));
  AOI21_X1   g27291(.A1(new_n29727_), .A2(new_n29166_), .B(new_n29695_), .ZN(new_n29728_));
  NOR2_X1    g27292(.A1(new_n29728_), .A2(pi1150), .ZN(new_n29729_));
  NOR2_X1    g27293(.A1(new_n28386_), .A2(new_n2628_), .ZN(new_n29730_));
  OAI21_X1   g27294(.A1(new_n8813_), .A2(new_n28005_), .B(new_n29730_), .ZN(new_n29731_));
  AOI21_X1   g27295(.A1(new_n29146_), .A2(new_n29731_), .B(new_n28422_), .ZN(new_n29732_));
  OAI21_X1   g27296(.A1(new_n29040_), .A2(pi0211), .B(pi0212), .ZN(new_n29733_));
  NOR2_X1    g27297(.A1(new_n29733_), .A2(new_n29043_), .ZN(new_n29734_));
  INV_X1     g27298(.I(new_n29734_), .ZN(new_n29735_));
  NOR2_X1    g27299(.A1(new_n29043_), .A2(pi0212), .ZN(new_n29736_));
  NAND2_X1   g27300(.A1(new_n29040_), .A2(new_n29736_), .ZN(new_n29737_));
  INV_X1     g27301(.I(new_n29737_), .ZN(new_n29738_));
  AOI21_X1   g27302(.A1(new_n29738_), .A2(new_n29188_), .B(pi0219), .ZN(new_n29739_));
  AOI21_X1   g27303(.A1(new_n29735_), .A2(new_n29739_), .B(new_n29726_), .ZN(new_n29740_));
  NAND2_X1   g27304(.A1(new_n29727_), .A2(new_n29129_), .ZN(new_n29741_));
  OAI21_X1   g27305(.A1(new_n29741_), .A2(new_n29740_), .B(new_n29732_), .ZN(new_n29742_));
  AOI21_X1   g27306(.A1(new_n29729_), .A2(new_n29742_), .B(pi1149), .ZN(new_n29743_));
  INV_X1     g27307(.I(new_n29523_), .ZN(new_n29744_));
  NOR2_X1    g27308(.A1(new_n29508_), .A2(new_n29705_), .ZN(new_n29745_));
  AOI21_X1   g27309(.A1(pi0214), .A2(new_n29745_), .B(new_n29513_), .ZN(new_n29746_));
  NAND2_X1   g27310(.A1(new_n29745_), .A2(new_n8511_), .ZN(new_n29747_));
  AOI21_X1   g27311(.A1(new_n29517_), .A2(new_n29747_), .B(new_n29746_), .ZN(new_n29748_));
  OAI21_X1   g27312(.A1(new_n29748_), .A2(pi0219), .B(new_n29744_), .ZN(new_n29749_));
  NOR2_X1    g27313(.A1(new_n29539_), .A2(new_n8510_), .ZN(new_n29750_));
  INV_X1     g27314(.I(new_n29750_), .ZN(new_n29751_));
  NOR2_X1    g27315(.A1(new_n28338_), .A2(pi0211), .ZN(new_n29752_));
  NOR2_X1    g27316(.A1(new_n28098_), .A2(new_n9171_), .ZN(new_n29753_));
  OAI21_X1   g27317(.A1(new_n29753_), .A2(new_n29024_), .B(new_n29752_), .ZN(new_n29754_));
  NAND2_X1   g27318(.A1(new_n29751_), .A2(new_n29754_), .ZN(new_n29755_));
  INV_X1     g27319(.I(new_n29755_), .ZN(new_n29756_));
  NAND2_X1   g27320(.A1(new_n29756_), .A2(new_n8511_), .ZN(new_n29757_));
  AOI21_X1   g27321(.A1(new_n29757_), .A2(new_n29625_), .B(pi0219), .ZN(new_n29758_));
  OAI21_X1   g27322(.A1(new_n29755_), .A2(new_n8511_), .B(new_n29542_), .ZN(new_n29759_));
  AOI21_X1   g27323(.A1(new_n29758_), .A2(new_n29759_), .B(new_n29623_), .ZN(new_n29760_));
  OAI21_X1   g27324(.A1(new_n29760_), .A2(new_n29718_), .B(pi1152), .ZN(new_n29761_));
  AOI21_X1   g27325(.A1(new_n29146_), .A2(new_n29749_), .B(new_n29761_), .ZN(new_n29762_));
  INV_X1     g27326(.I(new_n29754_), .ZN(new_n29763_));
  OAI21_X1   g27327(.A1(new_n29763_), .A2(new_n29546_), .B(new_n29542_), .ZN(new_n29764_));
  INV_X1     g27328(.I(new_n29541_), .ZN(new_n29765_));
  NOR2_X1    g27329(.A1(new_n29545_), .A2(new_n29765_), .ZN(new_n29766_));
  NOR2_X1    g27330(.A1(new_n29750_), .A2(new_n29009_), .ZN(new_n29767_));
  INV_X1     g27331(.I(new_n29767_), .ZN(new_n29768_));
  OAI21_X1   g27332(.A1(new_n29768_), .A2(new_n8511_), .B(pi0212), .ZN(new_n29769_));
  NOR2_X1    g27333(.A1(new_n29769_), .A2(new_n29766_), .ZN(new_n29770_));
  AOI21_X1   g27334(.A1(new_n29770_), .A2(new_n29755_), .B(pi0219), .ZN(new_n29771_));
  AOI21_X1   g27335(.A1(new_n29771_), .A2(new_n29764_), .B(new_n29623_), .ZN(new_n29772_));
  OAI21_X1   g27336(.A1(new_n29772_), .A2(new_n29165_), .B(new_n28422_), .ZN(new_n29773_));
  INV_X1     g27337(.I(new_n29508_), .ZN(new_n29774_));
  AOI21_X1   g27338(.A1(new_n29774_), .A2(new_n28580_), .B(pi0211), .ZN(new_n29775_));
  NAND2_X1   g27339(.A1(new_n29516_), .A2(new_n29158_), .ZN(new_n29776_));
  OAI22_X1   g27340(.A1(new_n29776_), .A2(new_n29775_), .B1(new_n29158_), .B2(new_n29503_), .ZN(new_n29777_));
  AOI21_X1   g27341(.A1(new_n29777_), .A2(new_n6643_), .B(new_n29691_), .ZN(new_n29778_));
  OAI21_X1   g27342(.A1(new_n29773_), .A2(new_n29778_), .B(pi1150), .ZN(new_n29779_));
  OAI21_X1   g27343(.A1(new_n29762_), .A2(new_n29779_), .B(new_n29743_), .ZN(new_n29780_));
  NAND3_X1   g27344(.A1(new_n29780_), .A2(pi0213), .A3(new_n29724_), .ZN(new_n29781_));
  AOI21_X1   g27345(.A1(new_n29669_), .A2(new_n29781_), .B(pi0209), .ZN(new_n29782_));
  AND2_X2    g27346(.A1(new_n29227_), .A2(pi0213), .Z(new_n29783_));
  INV_X1     g27347(.I(new_n29598_), .ZN(new_n29784_));
  NOR2_X1    g27348(.A1(new_n29095_), .A2(pi0299), .ZN(new_n29785_));
  INV_X1     g27349(.I(new_n29440_), .ZN(new_n29786_));
  AOI21_X1   g27350(.A1(new_n29086_), .A2(new_n8511_), .B(new_n8509_), .ZN(new_n29787_));
  AOI21_X1   g27351(.A1(new_n29786_), .A2(new_n29787_), .B(new_n29107_), .ZN(new_n29788_));
  OAI21_X1   g27352(.A1(new_n29788_), .A2(new_n29785_), .B(new_n8807_), .ZN(new_n29789_));
  NAND3_X1   g27353(.A1(new_n29789_), .A2(new_n28422_), .A3(new_n29784_), .ZN(new_n29790_));
  OAI21_X1   g27354(.A1(new_n29215_), .A2(new_n29220_), .B(new_n8807_), .ZN(new_n29791_));
  OAI21_X1   g27355(.A1(new_n29070_), .A2(pi0214), .B(pi0212), .ZN(new_n29792_));
  NOR2_X1    g27356(.A1(new_n29211_), .A2(new_n29792_), .ZN(new_n29793_));
  OAI21_X1   g27357(.A1(new_n29791_), .A2(new_n29793_), .B(pi1152), .ZN(new_n29794_));
  AOI21_X1   g27358(.A1(new_n29115_), .A2(pi0219), .B(po1038), .ZN(new_n29795_));
  INV_X1     g27359(.I(new_n29795_), .ZN(new_n29796_));
  AOI22_X1   g27360(.A1(new_n29790_), .A2(new_n29794_), .B1(new_n29482_), .B2(new_n29796_), .ZN(new_n29797_));
  NOR2_X1    g27361(.A1(new_n29797_), .A2(new_n29646_), .ZN(new_n29798_));
  INV_X1     g27362(.I(new_n29739_), .ZN(new_n29799_));
  NAND2_X1   g27363(.A1(new_n29046_), .A2(pi0214), .ZN(new_n29800_));
  AOI21_X1   g27364(.A1(new_n29734_), .A2(new_n29800_), .B(new_n29799_), .ZN(new_n29801_));
  NOR3_X1    g27365(.A1(new_n29180_), .A2(pi0299), .A3(new_n29061_), .ZN(new_n29802_));
  NOR2_X1    g27366(.A1(new_n29802_), .A2(new_n29801_), .ZN(new_n29803_));
  AOI21_X1   g27367(.A1(new_n29803_), .A2(new_n29795_), .B(pi1152), .ZN(new_n29804_));
  NOR3_X1    g27368(.A1(new_n29801_), .A2(new_n29802_), .A3(pi0219), .ZN(new_n29805_));
  OAI21_X1   g27369(.A1(new_n29805_), .A2(new_n29011_), .B(new_n6643_), .ZN(new_n29806_));
  AOI21_X1   g27370(.A1(new_n29806_), .A2(pi1152), .B(new_n29804_), .ZN(new_n29807_));
  NOR2_X1    g27371(.A1(new_n29381_), .A2(pi1151), .ZN(new_n29808_));
  INV_X1     g27372(.I(new_n29808_), .ZN(new_n29809_));
  OAI21_X1   g27373(.A1(new_n29807_), .A2(new_n29809_), .B(pi1150), .ZN(new_n29810_));
  NOR3_X1    g27374(.A1(new_n29012_), .A2(new_n28422_), .A3(new_n29111_), .ZN(new_n29811_));
  OAI21_X1   g27375(.A1(new_n6643_), .A2(new_n29299_), .B(pi1151), .ZN(new_n29812_));
  OAI21_X1   g27376(.A1(new_n29069_), .A2(new_n29315_), .B(new_n29209_), .ZN(new_n29813_));
  AOI21_X1   g27377(.A1(new_n29813_), .A2(pi1152), .B(po1038), .ZN(new_n29814_));
  AOI21_X1   g27378(.A1(new_n29106_), .A2(new_n29693_), .B(new_n29812_), .ZN(new_n29815_));
  AOI21_X1   g27379(.A1(new_n29007_), .A2(new_n29061_), .B(new_n29815_), .ZN(new_n29816_));
  OAI22_X1   g27380(.A1(new_n29816_), .A2(pi1152), .B1(new_n29812_), .B2(new_n29814_), .ZN(new_n29817_));
  NOR2_X1    g27381(.A1(new_n29817_), .A2(new_n29811_), .ZN(new_n29818_));
  OAI22_X1   g27382(.A1(new_n29798_), .A2(new_n29810_), .B1(pi1150), .B2(new_n29818_), .ZN(new_n29819_));
  NOR2_X1    g27383(.A1(new_n29795_), .A2(new_n29485_), .ZN(new_n29820_));
  INV_X1     g27384(.I(new_n29820_), .ZN(new_n29821_));
  NOR2_X1    g27385(.A1(new_n29017_), .A2(new_n8811_), .ZN(new_n29822_));
  NOR2_X1    g27386(.A1(new_n29177_), .A2(new_n29041_), .ZN(new_n29823_));
  NOR3_X1    g27387(.A1(new_n29823_), .A2(new_n8809_), .A3(new_n29011_), .ZN(new_n29824_));
  NOR2_X1    g27388(.A1(new_n29824_), .A2(new_n29822_), .ZN(new_n29825_));
  OAI22_X1   g27389(.A1(new_n29825_), .A2(pi0219), .B1(new_n29205_), .B2(new_n29821_), .ZN(new_n29826_));
  OAI21_X1   g27390(.A1(new_n29180_), .A2(new_n29061_), .B(new_n29821_), .ZN(new_n29827_));
  AOI22_X1   g27391(.A1(new_n29804_), .A2(new_n29827_), .B1(pi1152), .B2(new_n29826_), .ZN(new_n29828_));
  NOR3_X1    g27392(.A1(new_n29828_), .A2(pi1151), .A3(new_n29365_), .ZN(new_n29829_));
  NOR2_X1    g27393(.A1(new_n29785_), .A2(new_n29080_), .ZN(new_n29830_));
  NOR2_X1    g27394(.A1(new_n29830_), .A2(pi0219), .ZN(new_n29831_));
  NAND3_X1   g27395(.A1(new_n29191_), .A2(new_n28422_), .A3(new_n6643_), .ZN(new_n29832_));
  OAI21_X1   g27396(.A1(new_n29832_), .A2(new_n29831_), .B(new_n29663_), .ZN(new_n29833_));
  AOI21_X1   g27397(.A1(pi0212), .A2(new_n29070_), .B(new_n29791_), .ZN(new_n29834_));
  NOR2_X1    g27398(.A1(new_n29834_), .A2(new_n28422_), .ZN(new_n29835_));
  AOI21_X1   g27399(.A1(new_n29835_), .A2(new_n29214_), .B(new_n29833_), .ZN(new_n29836_));
  NOR3_X1    g27400(.A1(new_n29829_), .A2(new_n29650_), .A3(new_n29836_), .ZN(new_n29837_));
  OAI21_X1   g27401(.A1(new_n29180_), .A2(new_n29011_), .B(pi1152), .ZN(new_n29838_));
  AOI21_X1   g27402(.A1(new_n29206_), .A2(new_n29820_), .B(new_n29838_), .ZN(new_n29839_));
  OAI21_X1   g27403(.A1(new_n29827_), .A2(pi1152), .B(new_n29655_), .ZN(new_n29840_));
  NOR2_X1    g27404(.A1(new_n29839_), .A2(new_n29840_), .ZN(new_n29841_));
  NAND2_X1   g27405(.A1(new_n29190_), .A2(new_n8509_), .ZN(new_n29842_));
  OAI21_X1   g27406(.A1(new_n29189_), .A2(new_n29079_), .B(new_n8511_), .ZN(new_n29843_));
  NAND3_X1   g27407(.A1(new_n29193_), .A2(new_n29843_), .A3(pi0212), .ZN(new_n29844_));
  AOI21_X1   g27408(.A1(new_n29844_), .A2(new_n29842_), .B(pi0219), .ZN(new_n29845_));
  OAI21_X1   g27409(.A1(new_n29845_), .A2(new_n29832_), .B(new_n29651_), .ZN(new_n29846_));
  INV_X1     g27410(.I(new_n29214_), .ZN(new_n29847_));
  NAND2_X1   g27411(.A1(new_n29070_), .A2(new_n28297_), .ZN(new_n29848_));
  NAND3_X1   g27412(.A1(new_n29848_), .A2(pi0212), .A3(new_n29209_), .ZN(new_n29849_));
  AOI21_X1   g27413(.A1(new_n29212_), .A2(new_n29849_), .B(pi0219), .ZN(new_n29850_));
  NOR3_X1    g27414(.A1(new_n29847_), .A2(new_n28422_), .A3(new_n29850_), .ZN(new_n29851_));
  OAI21_X1   g27415(.A1(new_n29851_), .A2(new_n29846_), .B(new_n29650_), .ZN(new_n29852_));
  OAI21_X1   g27416(.A1(new_n29852_), .A2(new_n29841_), .B(pi1149), .ZN(new_n29853_));
  OAI22_X1   g27417(.A1(new_n29819_), .A2(pi1149), .B1(new_n29837_), .B2(new_n29853_), .ZN(new_n29854_));
  AOI21_X1   g27418(.A1(new_n29854_), .A2(new_n26198_), .B(new_n29783_), .ZN(new_n29855_));
  OAI21_X1   g27419(.A1(new_n29855_), .A2(new_n28360_), .B(pi0230), .ZN(new_n29856_));
  OAI22_X1   g27420(.A1(new_n29782_), .A2(new_n29856_), .B1(pi0230), .B2(new_n3948_), .ZN(po0398));
  NAND2_X1   g27421(.A1(new_n28793_), .A2(new_n2628_), .ZN(new_n29858_));
  AOI21_X1   g27422(.A1(pi0199), .A2(pi1144), .B(pi0200), .ZN(new_n29859_));
  AOI21_X1   g27423(.A1(new_n28795_), .A2(new_n29859_), .B(new_n29858_), .ZN(new_n29860_));
  NAND2_X1   g27424(.A1(new_n29860_), .A2(pi0207), .ZN(new_n29861_));
  NAND2_X1   g27425(.A1(new_n29304_), .A2(new_n29859_), .ZN(new_n29862_));
  NAND3_X1   g27426(.A1(new_n29301_), .A2(new_n29862_), .A3(new_n2628_), .ZN(new_n29863_));
  OAI21_X1   g27427(.A1(pi0207), .A2(new_n29863_), .B(new_n29861_), .ZN(new_n29864_));
  NAND2_X1   g27428(.A1(new_n29864_), .A2(pi0208), .ZN(new_n29865_));
  OAI22_X1   g27429(.A1(new_n28074_), .A2(new_n28212_), .B1(new_n8811_), .B2(new_n28080_), .ZN(new_n29866_));
  OAI21_X1   g27430(.A1(new_n28825_), .A2(new_n29863_), .B(new_n29866_), .ZN(new_n29867_));
  NOR2_X1    g27431(.A1(new_n29863_), .A2(new_n28371_), .ZN(new_n29868_));
  OAI22_X1   g27432(.A1(new_n29867_), .A2(pi0219), .B1(new_n28430_), .B2(new_n29868_), .ZN(new_n29869_));
  OAI21_X1   g27433(.A1(new_n29863_), .A2(new_n28371_), .B(pi0211), .ZN(new_n29870_));
  NOR2_X1    g27434(.A1(new_n29863_), .A2(new_n28825_), .ZN(new_n29871_));
  OR3_X2     g27435(.A1(new_n29871_), .A2(new_n28503_), .A3(new_n28087_), .Z(new_n29872_));
  AOI21_X1   g27436(.A1(new_n29872_), .A2(new_n29870_), .B(new_n8807_), .ZN(new_n29873_));
  OAI21_X1   g27437(.A1(new_n29873_), .A2(new_n29869_), .B(new_n29865_), .ZN(new_n29874_));
  NAND2_X1   g27438(.A1(new_n29874_), .A2(new_n6643_), .ZN(new_n29875_));
  NAND3_X1   g27439(.A1(new_n29875_), .A2(new_n26198_), .A3(new_n28093_), .ZN(new_n29876_));
  NOR2_X1    g27440(.A1(new_n29626_), .A2(pi0212), .ZN(new_n29877_));
  NOR2_X1    g27441(.A1(new_n28784_), .A2(new_n8511_), .ZN(new_n29878_));
  AOI21_X1   g27442(.A1(new_n8511_), .A2(new_n29404_), .B(new_n29878_), .ZN(new_n29879_));
  NOR2_X1    g27443(.A1(new_n29879_), .A2(new_n8509_), .ZN(new_n29880_));
  OAI21_X1   g27444(.A1(new_n29880_), .A2(new_n29877_), .B(new_n8807_), .ZN(new_n29881_));
  AOI21_X1   g27445(.A1(new_n8510_), .A2(pi1144), .B(new_n8807_), .ZN(new_n29882_));
  INV_X1     g27446(.I(new_n29882_), .ZN(new_n29883_));
  NAND2_X1   g27447(.A1(new_n29881_), .A2(new_n29883_), .ZN(new_n29884_));
  NOR2_X1    g27448(.A1(new_n29884_), .A2(new_n28060_), .ZN(new_n29885_));
  INV_X1     g27449(.I(new_n29865_), .ZN(new_n29886_));
  NOR2_X1    g27450(.A1(new_n29886_), .A2(new_n29868_), .ZN(new_n29887_));
  INV_X1     g27451(.I(new_n29887_), .ZN(new_n29888_));
  AOI21_X1   g27452(.A1(new_n29888_), .A2(new_n28503_), .B(new_n8807_), .ZN(new_n29889_));
  NOR2_X1    g27453(.A1(new_n29886_), .A2(new_n29871_), .ZN(new_n29890_));
  INV_X1     g27454(.I(new_n29890_), .ZN(new_n29891_));
  OAI21_X1   g27455(.A1(new_n29891_), .A2(new_n28214_), .B(new_n28057_), .ZN(new_n29892_));
  AOI21_X1   g27456(.A1(new_n29889_), .A2(new_n29892_), .B(po1038), .ZN(new_n29893_));
  NAND3_X1   g27457(.A1(new_n29890_), .A2(pi0211), .A3(new_n28223_), .ZN(new_n29894_));
  NOR2_X1    g27458(.A1(new_n29891_), .A2(new_n28879_), .ZN(new_n29895_));
  NAND2_X1   g27459(.A1(new_n29895_), .A2(new_n8510_), .ZN(new_n29896_));
  AOI21_X1   g27460(.A1(new_n29896_), .A2(new_n29894_), .B(new_n8511_), .ZN(new_n29897_));
  INV_X1     g27461(.I(new_n29895_), .ZN(new_n29898_));
  NOR2_X1    g27462(.A1(new_n29898_), .A2(new_n8510_), .ZN(new_n29899_));
  NOR2_X1    g27463(.A1(new_n29891_), .A2(new_n29316_), .ZN(new_n29900_));
  AOI21_X1   g27464(.A1(new_n8510_), .A2(new_n29900_), .B(new_n29899_), .ZN(new_n29901_));
  OAI21_X1   g27465(.A1(new_n29901_), .A2(pi0214), .B(pi0212), .ZN(new_n29902_));
  NAND2_X1   g27466(.A1(new_n29887_), .A2(new_n8511_), .ZN(new_n29903_));
  NAND2_X1   g27467(.A1(new_n29903_), .A2(new_n8509_), .ZN(new_n29904_));
  NOR2_X1    g27468(.A1(new_n29901_), .A2(new_n8511_), .ZN(new_n29905_));
  NOR2_X1    g27469(.A1(new_n29905_), .A2(new_n29904_), .ZN(new_n29906_));
  NOR2_X1    g27470(.A1(new_n29906_), .A2(pi0219), .ZN(new_n29907_));
  OAI21_X1   g27471(.A1(new_n29897_), .A2(new_n29902_), .B(new_n29907_), .ZN(new_n29908_));
  AOI21_X1   g27472(.A1(new_n29908_), .A2(new_n29893_), .B(new_n29885_), .ZN(new_n29909_));
  NAND2_X1   g27473(.A1(new_n29909_), .A2(pi0213), .ZN(new_n29910_));
  AOI21_X1   g27474(.A1(new_n29910_), .A2(new_n29876_), .B(new_n28360_), .ZN(new_n29911_));
  AOI21_X1   g27475(.A1(pi0219), .A2(new_n28056_), .B(new_n29884_), .ZN(new_n29912_));
  NAND2_X1   g27476(.A1(new_n29912_), .A2(pi0299), .ZN(new_n29913_));
  AOI21_X1   g27477(.A1(new_n29913_), .A2(new_n28083_), .B(po1038), .ZN(new_n29914_));
  NOR3_X1    g27478(.A1(new_n29914_), .A2(new_n26198_), .A3(new_n29885_), .ZN(new_n29915_));
  AOI21_X1   g27479(.A1(new_n28090_), .A2(new_n26198_), .B(new_n29915_), .ZN(new_n29916_));
  OAI21_X1   g27480(.A1(new_n29916_), .A2(pi0209), .B(pi0230), .ZN(new_n29917_));
  OAI22_X1   g27481(.A1(new_n29911_), .A2(new_n29917_), .B1(pi0230), .B2(new_n5143_), .ZN(po0399));
  OAI22_X1   g27482(.A1(new_n8641_), .A2(pi1155), .B1(new_n8531_), .B2(pi1156), .ZN(new_n29919_));
  AOI21_X1   g27483(.A1(new_n8531_), .A2(pi1157), .B(new_n8525_), .ZN(new_n29920_));
  OAI21_X1   g27484(.A1(new_n29919_), .A2(new_n29920_), .B(new_n12618_), .ZN(new_n29921_));
  NOR2_X1    g27485(.A1(new_n28017_), .A2(new_n28010_), .ZN(new_n29922_));
  INV_X1     g27486(.I(new_n29922_), .ZN(new_n29923_));
  AOI22_X1   g27487(.A1(new_n29923_), .A2(new_n8807_), .B1(pi1157), .B2(new_n8808_), .ZN(new_n29924_));
  NAND2_X1   g27488(.A1(new_n25319_), .A2(new_n29924_), .ZN(new_n29925_));
  NAND2_X1   g27489(.A1(new_n29925_), .A2(new_n29921_), .ZN(new_n29926_));
  INV_X1     g27490(.I(pi0268), .ZN(new_n29927_));
  INV_X1     g27491(.I(pi0272), .ZN(new_n29928_));
  INV_X1     g27492(.I(pi0275), .ZN(new_n29929_));
  INV_X1     g27493(.I(pi0283), .ZN(new_n29930_));
  NOR3_X1    g27494(.A1(new_n29928_), .A2(new_n29929_), .A3(new_n29930_), .ZN(new_n29931_));
  INV_X1     g27495(.I(new_n29931_), .ZN(new_n29932_));
  NOR2_X1    g27496(.A1(new_n29932_), .A2(new_n29927_), .ZN(new_n29933_));
  INV_X1     g27497(.I(new_n29933_), .ZN(new_n29934_));
  INV_X1     g27498(.I(pi0243), .ZN(new_n29935_));
  NOR2_X1    g27499(.A1(new_n29935_), .A2(pi1091), .ZN(new_n29936_));
  NOR2_X1    g27500(.A1(new_n28894_), .A2(pi0299), .ZN(new_n29937_));
  NOR2_X1    g27501(.A1(new_n29937_), .A2(new_n3022_), .ZN(new_n29938_));
  NOR2_X1    g27502(.A1(new_n29938_), .A2(new_n29936_), .ZN(new_n29939_));
  NAND2_X1   g27503(.A1(new_n29939_), .A2(new_n12770_), .ZN(new_n29940_));
  NOR2_X1    g27504(.A1(new_n28132_), .A2(new_n3022_), .ZN(new_n29941_));
  INV_X1     g27505(.I(new_n29941_), .ZN(new_n29942_));
  NOR2_X1    g27506(.A1(new_n29936_), .A2(new_n12770_), .ZN(new_n29943_));
  AOI21_X1   g27507(.A1(new_n29942_), .A2(new_n29943_), .B(pi1156), .ZN(new_n29944_));
  NOR2_X1    g27508(.A1(pi0243), .A2(pi1091), .ZN(new_n29945_));
  NOR2_X1    g27509(.A1(new_n3022_), .A2(pi0299), .ZN(new_n29946_));
  AOI21_X1   g27510(.A1(new_n28559_), .A2(new_n29946_), .B(new_n29945_), .ZN(new_n29947_));
  NOR2_X1    g27511(.A1(new_n9172_), .A2(new_n3022_), .ZN(new_n29948_));
  INV_X1     g27512(.I(new_n29948_), .ZN(new_n29949_));
  AOI21_X1   g27513(.A1(new_n29949_), .A2(new_n29943_), .B(new_n12742_), .ZN(new_n29950_));
  AOI22_X1   g27514(.A1(new_n29940_), .A2(new_n29944_), .B1(new_n29947_), .B2(new_n29950_), .ZN(new_n29951_));
  NAND2_X1   g27515(.A1(new_n29951_), .A2(pi1157), .ZN(new_n29952_));
  INV_X1     g27516(.I(new_n29936_), .ZN(new_n29953_));
  OAI21_X1   g27517(.A1(new_n9217_), .A2(new_n3022_), .B(new_n12770_), .ZN(new_n29954_));
  OAI21_X1   g27518(.A1(new_n12770_), .A2(new_n29948_), .B(new_n29954_), .ZN(new_n29955_));
  NAND3_X1   g27519(.A1(new_n29946_), .A2(pi0200), .A3(new_n12742_), .ZN(new_n29956_));
  NAND4_X1   g27520(.A1(new_n29955_), .A2(new_n12965_), .A3(new_n29953_), .A4(new_n29956_), .ZN(new_n29957_));
  AOI21_X1   g27521(.A1(new_n29952_), .A2(new_n29957_), .B(pi0211), .ZN(new_n29958_));
  NAND2_X1   g27522(.A1(new_n28736_), .A2(new_n29946_), .ZN(new_n29959_));
  NAND3_X1   g27523(.A1(new_n29959_), .A2(new_n12770_), .A3(new_n29953_), .ZN(new_n29960_));
  NAND2_X1   g27524(.A1(new_n29950_), .A2(new_n29960_), .ZN(new_n29961_));
  AOI21_X1   g27525(.A1(pi1091), .A2(pi1155), .B(new_n29945_), .ZN(new_n29962_));
  NOR2_X1    g27526(.A1(new_n10288_), .A2(new_n3022_), .ZN(new_n29963_));
  OAI21_X1   g27527(.A1(new_n29963_), .A2(new_n29962_), .B(new_n12742_), .ZN(new_n29964_));
  NAND3_X1   g27528(.A1(new_n29961_), .A2(new_n12965_), .A3(new_n29964_), .ZN(new_n29965_));
  NOR2_X1    g27529(.A1(new_n29962_), .A2(new_n28136_), .ZN(new_n29966_));
  OAI21_X1   g27530(.A1(new_n29939_), .A2(new_n29966_), .B(new_n12742_), .ZN(new_n29967_));
  INV_X1     g27531(.I(new_n29947_), .ZN(new_n29968_));
  INV_X1     g27532(.I(new_n29963_), .ZN(new_n29969_));
  NOR2_X1    g27533(.A1(new_n29969_), .A2(new_n28465_), .ZN(new_n29970_));
  OAI21_X1   g27534(.A1(new_n29968_), .A2(new_n29970_), .B(pi1156), .ZN(new_n29971_));
  NAND2_X1   g27535(.A1(new_n29971_), .A2(new_n29967_), .ZN(new_n29972_));
  NAND2_X1   g27536(.A1(new_n29972_), .A2(pi1157), .ZN(new_n29973_));
  AOI21_X1   g27537(.A1(new_n29973_), .A2(new_n29965_), .B(new_n8510_), .ZN(new_n29974_));
  OAI21_X1   g27538(.A1(new_n29974_), .A2(new_n29958_), .B(new_n8807_), .ZN(new_n29975_));
  NAND2_X1   g27539(.A1(new_n29968_), .A2(pi1156), .ZN(new_n29976_));
  NAND3_X1   g27540(.A1(new_n29976_), .A2(new_n29967_), .A3(new_n28808_), .ZN(new_n29977_));
  NOR2_X1    g27541(.A1(new_n2628_), .A2(new_n3022_), .ZN(new_n29978_));
  INV_X1     g27542(.I(new_n29978_), .ZN(new_n29979_));
  NAND4_X1   g27543(.A1(new_n29955_), .A2(new_n29953_), .A3(new_n29956_), .A4(new_n29979_), .ZN(new_n29980_));
  NAND2_X1   g27544(.A1(new_n29980_), .A2(new_n12965_), .ZN(new_n29981_));
  NAND3_X1   g27545(.A1(new_n28284_), .A2(pi1091), .A3(new_n28286_), .ZN(new_n29982_));
  NAND3_X1   g27546(.A1(new_n29982_), .A2(new_n12742_), .A3(new_n29953_), .ZN(new_n29983_));
  NAND3_X1   g27547(.A1(new_n29971_), .A2(new_n29983_), .A3(new_n28018_), .ZN(new_n29984_));
  NAND4_X1   g27548(.A1(new_n29984_), .A2(new_n29977_), .A3(new_n29981_), .A4(pi0219), .ZN(new_n29985_));
  AOI21_X1   g27549(.A1(new_n29975_), .A2(new_n29985_), .B(po1038), .ZN(new_n29986_));
  AOI21_X1   g27550(.A1(new_n29924_), .A2(pi1091), .B(new_n29936_), .ZN(new_n29987_));
  AND2_X2    g27551(.A1(new_n29987_), .A2(po1038), .Z(new_n29988_));
  OAI21_X1   g27552(.A1(new_n29986_), .A2(new_n29988_), .B(new_n29934_), .ZN(new_n29989_));
  INV_X1     g27553(.I(pi0267), .ZN(new_n29990_));
  INV_X1     g27554(.I(pi0253), .ZN(new_n29991_));
  INV_X1     g27555(.I(pi0254), .ZN(new_n29992_));
  NOR2_X1    g27556(.A1(new_n29991_), .A2(new_n29992_), .ZN(new_n29993_));
  INV_X1     g27557(.I(new_n29993_), .ZN(new_n29994_));
  NOR2_X1    g27558(.A1(new_n29994_), .A2(new_n29990_), .ZN(new_n29995_));
  INV_X1     g27559(.I(new_n29995_), .ZN(new_n29996_));
  NOR2_X1    g27560(.A1(new_n29996_), .A2(pi0263), .ZN(new_n29997_));
  INV_X1     g27561(.I(new_n29997_), .ZN(new_n29998_));
  INV_X1     g27562(.I(pi0273), .ZN(new_n29999_));
  INV_X1     g27563(.I(pi0271), .ZN(new_n30000_));
  INV_X1     g27564(.I(pi0802), .ZN(new_n30001_));
  NOR2_X1    g27565(.A1(pi0083), .A2(pi0085), .ZN(new_n30002_));
  AOI21_X1   g27566(.A1(new_n30002_), .A2(new_n2500_), .B(new_n5590_), .ZN(new_n30003_));
  INV_X1     g27567(.I(new_n30003_), .ZN(new_n30004_));
  NOR2_X1    g27568(.A1(new_n30004_), .A2(new_n30001_), .ZN(new_n30005_));
  NAND2_X1   g27569(.A1(new_n30005_), .A2(pi0276), .ZN(new_n30006_));
  NOR2_X1    g27570(.A1(new_n30006_), .A2(pi1091), .ZN(new_n30007_));
  INV_X1     g27571(.I(new_n30007_), .ZN(new_n30008_));
  NOR2_X1    g27572(.A1(new_n30008_), .A2(new_n30000_), .ZN(new_n30009_));
  INV_X1     g27573(.I(new_n30009_), .ZN(new_n30010_));
  NOR2_X1    g27574(.A1(new_n30010_), .A2(new_n29999_), .ZN(new_n30011_));
  INV_X1     g27575(.I(new_n30011_), .ZN(new_n30012_));
  OAI22_X1   g27576(.A1(new_n30012_), .A2(pi0243), .B1(new_n3022_), .B2(new_n29923_), .ZN(new_n30013_));
  NOR2_X1    g27577(.A1(new_n30002_), .A2(new_n5590_), .ZN(new_n30014_));
  INV_X1     g27578(.I(new_n30014_), .ZN(new_n30015_));
  NOR3_X1    g27579(.A1(new_n30015_), .A2(new_n3293_), .A3(new_n30001_), .ZN(new_n30016_));
  INV_X1     g27580(.I(new_n30016_), .ZN(new_n30017_));
  NOR2_X1    g27581(.A1(new_n30017_), .A2(new_n30000_), .ZN(new_n30018_));
  OAI21_X1   g27582(.A1(new_n30018_), .A2(pi1091), .B(pi0273), .ZN(new_n30019_));
  NAND2_X1   g27583(.A1(new_n30019_), .A2(new_n3022_), .ZN(new_n30020_));
  NOR2_X1    g27584(.A1(new_n30011_), .A2(new_n30020_), .ZN(new_n30021_));
  INV_X1     g27585(.I(new_n30021_), .ZN(new_n30022_));
  NOR2_X1    g27586(.A1(new_n30022_), .A2(new_n29935_), .ZN(new_n30023_));
  NOR3_X1    g27587(.A1(new_n30023_), .A2(pi0219), .A3(new_n30013_), .ZN(new_n30024_));
  NOR2_X1    g27588(.A1(new_n30017_), .A2(pi1091), .ZN(new_n30025_));
  INV_X1     g27589(.I(new_n30025_), .ZN(new_n30026_));
  NAND3_X1   g27590(.A1(new_n30026_), .A2(new_n28018_), .A3(new_n29953_), .ZN(new_n30027_));
  NAND2_X1   g27591(.A1(new_n30020_), .A2(new_n29935_), .ZN(new_n30028_));
  NOR3_X1    g27592(.A1(new_n30026_), .A2(new_n30000_), .A3(new_n29999_), .ZN(new_n30029_));
  OAI21_X1   g27593(.A1(new_n29935_), .A2(new_n30029_), .B(new_n30028_), .ZN(new_n30030_));
  AOI21_X1   g27594(.A1(new_n30030_), .A2(new_n30027_), .B(new_n8807_), .ZN(new_n30031_));
  NOR3_X1    g27595(.A1(new_n30024_), .A2(new_n29998_), .A3(new_n30031_), .ZN(new_n30032_));
  NOR2_X1    g27596(.A1(new_n29987_), .A2(new_n29997_), .ZN(new_n30033_));
  OAI21_X1   g27597(.A1(new_n30032_), .A2(new_n30033_), .B(po1038), .ZN(new_n30034_));
  NAND2_X1   g27598(.A1(new_n29975_), .A2(new_n29985_), .ZN(new_n30035_));
  AOI21_X1   g27599(.A1(new_n30035_), .A2(new_n29998_), .B(po1038), .ZN(new_n30036_));
  INV_X1     g27600(.I(new_n30020_), .ZN(new_n30037_));
  NOR2_X1    g27601(.A1(new_n30037_), .A2(new_n8525_), .ZN(new_n30038_));
  OAI21_X1   g27602(.A1(new_n30012_), .A2(pi0199), .B(new_n30037_), .ZN(new_n30039_));
  NAND2_X1   g27603(.A1(new_n30039_), .A2(new_n30007_), .ZN(new_n30040_));
  NAND2_X1   g27604(.A1(new_n30040_), .A2(new_n2628_), .ZN(new_n30041_));
  NOR2_X1    g27605(.A1(new_n30041_), .A2(new_n30038_), .ZN(new_n30042_));
  NAND2_X1   g27606(.A1(new_n30042_), .A2(pi0243), .ZN(new_n30043_));
  NOR2_X1    g27607(.A1(new_n30021_), .A2(pi0199), .ZN(new_n30044_));
  NAND2_X1   g27608(.A1(new_n30008_), .A2(new_n8531_), .ZN(new_n30045_));
  NAND2_X1   g27609(.A1(new_n30039_), .A2(new_n30045_), .ZN(new_n30046_));
  NAND2_X1   g27610(.A1(new_n30046_), .A2(new_n2628_), .ZN(new_n30047_));
  NOR2_X1    g27611(.A1(new_n30047_), .A2(new_n30044_), .ZN(new_n30048_));
  NOR2_X1    g27612(.A1(new_n30029_), .A2(new_n2628_), .ZN(new_n30049_));
  NOR2_X1    g27613(.A1(new_n30048_), .A2(new_n30049_), .ZN(new_n30050_));
  NAND2_X1   g27614(.A1(new_n30050_), .A2(new_n29935_), .ZN(new_n30051_));
  AOI21_X1   g27615(.A1(new_n30051_), .A2(new_n30043_), .B(pi1155), .ZN(new_n30052_));
  INV_X1     g27616(.I(new_n30047_), .ZN(new_n30053_));
  NOR2_X1    g27617(.A1(new_n30053_), .A2(new_n30049_), .ZN(new_n30054_));
  INV_X1     g27618(.I(new_n30054_), .ZN(new_n30055_));
  NOR3_X1    g27619(.A1(new_n30055_), .A2(pi0243), .A3(new_n12770_), .ZN(new_n30056_));
  NOR2_X1    g27620(.A1(new_n30037_), .A2(pi0200), .ZN(new_n30057_));
  NOR2_X1    g27621(.A1(new_n30041_), .A2(new_n30057_), .ZN(new_n30058_));
  NOR2_X1    g27622(.A1(new_n30020_), .A2(new_n2628_), .ZN(new_n30059_));
  NOR2_X1    g27623(.A1(new_n30058_), .A2(new_n30059_), .ZN(new_n30060_));
  NOR2_X1    g27624(.A1(new_n30060_), .A2(new_n29935_), .ZN(new_n30061_));
  NOR4_X1    g27625(.A1(new_n30052_), .A2(pi1156), .A3(new_n30056_), .A4(new_n30061_), .ZN(new_n30062_));
  NOR2_X1    g27626(.A1(new_n30047_), .A2(new_n30038_), .ZN(new_n30063_));
  INV_X1     g27627(.I(new_n30058_), .ZN(new_n30064_));
  NOR2_X1    g27628(.A1(new_n30064_), .A2(new_n30044_), .ZN(new_n30065_));
  NOR2_X1    g27629(.A1(new_n30065_), .A2(new_n30049_), .ZN(new_n30066_));
  INV_X1     g27630(.I(new_n30066_), .ZN(new_n30067_));
  NOR2_X1    g27631(.A1(new_n30067_), .A2(new_n30063_), .ZN(new_n30068_));
  INV_X1     g27632(.I(new_n30068_), .ZN(new_n30069_));
  AOI21_X1   g27633(.A1(new_n30069_), .A2(new_n30061_), .B(new_n12770_), .ZN(new_n30070_));
  INV_X1     g27634(.I(new_n30042_), .ZN(new_n30071_));
  NOR2_X1    g27635(.A1(new_n30071_), .A2(new_n30057_), .ZN(new_n30072_));
  NOR2_X1    g27636(.A1(new_n30072_), .A2(new_n30059_), .ZN(new_n30073_));
  NAND3_X1   g27637(.A1(new_n30073_), .A2(new_n29935_), .A3(new_n30054_), .ZN(new_n30074_));
  NAND2_X1   g27638(.A1(new_n30070_), .A2(new_n30074_), .ZN(new_n30075_));
  NAND2_X1   g27639(.A1(new_n30068_), .A2(pi0243), .ZN(new_n30076_));
  OAI21_X1   g27640(.A1(pi0243), .A2(new_n30073_), .B(new_n30076_), .ZN(new_n30077_));
  NOR2_X1    g27641(.A1(new_n30048_), .A2(new_n30059_), .ZN(new_n30078_));
  NOR2_X1    g27642(.A1(new_n30078_), .A2(pi0243), .ZN(new_n30079_));
  INV_X1     g27643(.I(new_n30079_), .ZN(new_n30080_));
  NOR2_X1    g27644(.A1(new_n30011_), .A2(new_n2628_), .ZN(new_n30081_));
  NOR2_X1    g27645(.A1(new_n30072_), .A2(new_n30081_), .ZN(new_n30082_));
  AOI21_X1   g27646(.A1(new_n30082_), .A2(new_n30080_), .B(new_n29936_), .ZN(new_n30083_));
  OAI21_X1   g27647(.A1(new_n30077_), .A2(new_n30083_), .B(new_n12770_), .ZN(new_n30084_));
  AOI21_X1   g27648(.A1(new_n30084_), .A2(new_n30075_), .B(new_n12742_), .ZN(new_n30085_));
  NOR4_X1    g27649(.A1(new_n30085_), .A2(pi0211), .A3(new_n12965_), .A4(new_n30062_), .ZN(new_n30086_));
  INV_X1     g27650(.I(new_n30077_), .ZN(new_n30087_));
  NOR2_X1    g27651(.A1(new_n30022_), .A2(new_n2628_), .ZN(new_n30088_));
  NOR2_X1    g27652(.A1(new_n30053_), .A2(new_n30088_), .ZN(new_n30089_));
  INV_X1     g27653(.I(new_n30089_), .ZN(new_n30090_));
  NOR2_X1    g27654(.A1(new_n30090_), .A2(pi0243), .ZN(new_n30091_));
  AOI21_X1   g27655(.A1(new_n30067_), .A2(pi0243), .B(new_n30091_), .ZN(new_n30092_));
  NAND2_X1   g27656(.A1(new_n30080_), .A2(new_n12770_), .ZN(new_n30093_));
  OAI21_X1   g27657(.A1(new_n30092_), .A2(new_n12770_), .B(new_n30093_), .ZN(new_n30094_));
  AOI21_X1   g27658(.A1(new_n30087_), .A2(new_n30094_), .B(new_n12742_), .ZN(new_n30095_));
  NOR2_X1    g27659(.A1(new_n30058_), .A2(new_n30049_), .ZN(new_n30096_));
  NOR2_X1    g27660(.A1(new_n30096_), .A2(new_n29935_), .ZN(new_n30097_));
  NOR3_X1    g27661(.A1(new_n30091_), .A2(new_n12770_), .A3(new_n30097_), .ZN(new_n30098_));
  INV_X1     g27662(.I(new_n30096_), .ZN(new_n30099_));
  NOR3_X1    g27663(.A1(new_n30099_), .A2(new_n29935_), .A3(new_n30042_), .ZN(new_n30100_));
  NOR3_X1    g27664(.A1(new_n30098_), .A2(new_n30100_), .A3(new_n30079_), .ZN(new_n30101_));
  OAI21_X1   g27665(.A1(new_n30101_), .A2(pi1156), .B(new_n28808_), .ZN(new_n30102_));
  NOR2_X1    g27666(.A1(new_n30041_), .A2(new_n30044_), .ZN(new_n30103_));
  NOR2_X1    g27667(.A1(new_n30103_), .A2(new_n30049_), .ZN(new_n30104_));
  INV_X1     g27668(.I(new_n30104_), .ZN(new_n30105_));
  NOR2_X1    g27669(.A1(new_n30105_), .A2(new_n30058_), .ZN(new_n30106_));
  INV_X1     g27670(.I(new_n30106_), .ZN(new_n30107_));
  NOR2_X1    g27671(.A1(new_n30107_), .A2(new_n29935_), .ZN(new_n30108_));
  NOR2_X1    g27672(.A1(new_n30063_), .A2(new_n30059_), .ZN(new_n30109_));
  OAI21_X1   g27673(.A1(new_n30109_), .A2(pi0243), .B(pi1155), .ZN(new_n30110_));
  OAI21_X1   g27674(.A1(new_n30108_), .A2(new_n30110_), .B(new_n12742_), .ZN(new_n30111_));
  INV_X1     g27675(.I(new_n30041_), .ZN(new_n30112_));
  NOR2_X1    g27676(.A1(new_n30112_), .A2(new_n30049_), .ZN(new_n30113_));
  NOR3_X1    g27677(.A1(new_n30113_), .A2(pi0243), .A3(pi1091), .ZN(new_n30114_));
  INV_X1     g27678(.I(new_n30113_), .ZN(new_n30115_));
  NOR2_X1    g27679(.A1(new_n30115_), .A2(new_n29935_), .ZN(new_n30116_));
  NOR3_X1    g27680(.A1(new_n30116_), .A2(pi1155), .A3(new_n30114_), .ZN(new_n30117_));
  OAI21_X1   g27681(.A1(new_n30111_), .A2(new_n30117_), .B(new_n12965_), .ZN(new_n30118_));
  NOR2_X1    g27682(.A1(new_n30058_), .A2(new_n30081_), .ZN(new_n30119_));
  INV_X1     g27683(.I(new_n30119_), .ZN(new_n30120_));
  NOR3_X1    g27684(.A1(new_n30120_), .A2(pi1155), .A3(new_n30007_), .ZN(new_n30121_));
  NOR2_X1    g27685(.A1(new_n30042_), .A2(new_n30059_), .ZN(new_n30122_));
  OR3_X2     g27686(.A1(new_n30121_), .A2(pi0243), .A3(new_n30122_), .Z(new_n30123_));
  NAND2_X1   g27687(.A1(new_n30053_), .A2(new_n12770_), .ZN(new_n30124_));
  NAND3_X1   g27688(.A1(new_n30104_), .A2(new_n30124_), .A3(pi0243), .ZN(new_n30125_));
  AOI21_X1   g27689(.A1(new_n30123_), .A2(new_n30125_), .B(new_n12742_), .ZN(new_n30126_));
  OAI22_X1   g27690(.A1(new_n30095_), .A2(new_n30102_), .B1(new_n30118_), .B2(new_n30126_), .ZN(new_n30127_));
  OAI21_X1   g27691(.A1(new_n30086_), .A2(new_n30127_), .B(pi0219), .ZN(new_n30128_));
  INV_X1     g27692(.I(new_n30082_), .ZN(new_n30129_));
  NOR2_X1    g27693(.A1(new_n30053_), .A2(new_n30081_), .ZN(new_n30130_));
  NOR2_X1    g27694(.A1(new_n30072_), .A2(pi0243), .ZN(new_n30131_));
  NOR2_X1    g27695(.A1(new_n30065_), .A2(new_n30088_), .ZN(new_n30132_));
  INV_X1     g27696(.I(new_n30132_), .ZN(new_n30133_));
  NOR2_X1    g27697(.A1(new_n30133_), .A2(new_n12770_), .ZN(new_n30134_));
  NOR2_X1    g27698(.A1(new_n30070_), .A2(new_n30134_), .ZN(new_n30135_));
  AOI21_X1   g27699(.A1(new_n30130_), .A2(new_n30131_), .B(new_n30135_), .ZN(new_n30136_));
  NOR2_X1    g27700(.A1(new_n30072_), .A2(new_n30048_), .ZN(new_n30137_));
  INV_X1     g27701(.I(new_n30137_), .ZN(new_n30138_));
  OAI21_X1   g27702(.A1(new_n30138_), .A2(new_n30088_), .B(new_n29935_), .ZN(new_n30139_));
  INV_X1     g27703(.I(new_n30065_), .ZN(new_n30140_));
  NOR2_X1    g27704(.A1(new_n30063_), .A2(new_n30081_), .ZN(new_n30141_));
  NAND3_X1   g27705(.A1(new_n30140_), .A2(pi0243), .A3(new_n30141_), .ZN(new_n30142_));
  AOI21_X1   g27706(.A1(new_n30139_), .A2(new_n30142_), .B(pi1155), .ZN(new_n30143_));
  NOR2_X1    g27707(.A1(new_n30136_), .A2(new_n30143_), .ZN(new_n30144_));
  INV_X1     g27708(.I(new_n30144_), .ZN(new_n30145_));
  AOI21_X1   g27709(.A1(new_n29953_), .A2(new_n30129_), .B(new_n30145_), .ZN(new_n30146_));
  NOR2_X1    g27710(.A1(new_n30119_), .A2(new_n29935_), .ZN(new_n30147_));
  OAI21_X1   g27711(.A1(new_n30091_), .A2(new_n30147_), .B(pi1155), .ZN(new_n30148_));
  NOR2_X1    g27712(.A1(new_n30042_), .A2(new_n30081_), .ZN(new_n30149_));
  INV_X1     g27713(.I(new_n30149_), .ZN(new_n30150_));
  NOR2_X1    g27714(.A1(new_n30150_), .A2(new_n30058_), .ZN(new_n30151_));
  NAND2_X1   g27715(.A1(new_n30151_), .A2(pi0243), .ZN(new_n30152_));
  NOR2_X1    g27716(.A1(new_n30112_), .A2(new_n30081_), .ZN(new_n30153_));
  NOR2_X1    g27717(.A1(new_n30080_), .A2(new_n30153_), .ZN(new_n30154_));
  NOR2_X1    g27718(.A1(new_n30154_), .A2(pi1155), .ZN(new_n30155_));
  AOI21_X1   g27719(.A1(new_n30155_), .A2(new_n30152_), .B(pi1156), .ZN(new_n30156_));
  AOI21_X1   g27720(.A1(new_n30156_), .A2(new_n30148_), .B(new_n12965_), .ZN(new_n30157_));
  OAI21_X1   g27721(.A1(new_n30146_), .A2(new_n12742_), .B(new_n30157_), .ZN(new_n30158_));
  NOR2_X1    g27722(.A1(new_n30149_), .A2(pi0243), .ZN(new_n30159_));
  NOR2_X1    g27723(.A1(new_n30103_), .A2(new_n30088_), .ZN(new_n30160_));
  AOI21_X1   g27724(.A1(pi0243), .A2(new_n30160_), .B(new_n30159_), .ZN(new_n30161_));
  NOR3_X1    g27725(.A1(new_n30161_), .A2(new_n12742_), .A3(new_n30121_), .ZN(new_n30162_));
  INV_X1     g27726(.I(new_n30162_), .ZN(new_n30163_));
  NAND2_X1   g27727(.A1(new_n30038_), .A2(new_n29943_), .ZN(new_n30164_));
  NAND2_X1   g27728(.A1(new_n30153_), .A2(new_n29935_), .ZN(new_n30165_));
  OAI21_X1   g27729(.A1(new_n30114_), .A2(new_n30153_), .B(new_n30165_), .ZN(new_n30166_));
  AOI21_X1   g27730(.A1(new_n30166_), .A2(new_n12770_), .B(pi1156), .ZN(new_n30167_));
  NAND3_X1   g27731(.A1(new_n30167_), .A2(new_n30148_), .A3(new_n30164_), .ZN(new_n30168_));
  NAND3_X1   g27732(.A1(new_n30168_), .A2(new_n30163_), .A3(new_n12965_), .ZN(new_n30169_));
  NAND3_X1   g27733(.A1(new_n30158_), .A2(pi0211), .A3(new_n30169_), .ZN(new_n30170_));
  NOR2_X1    g27734(.A1(new_n30130_), .A2(pi0243), .ZN(new_n30171_));
  NOR2_X1    g27735(.A1(new_n30058_), .A2(new_n30088_), .ZN(new_n30172_));
  AOI21_X1   g27736(.A1(pi0243), .A2(new_n30172_), .B(new_n30171_), .ZN(new_n30173_));
  OAI21_X1   g27737(.A1(new_n30161_), .A2(new_n30173_), .B(pi1155), .ZN(new_n30174_));
  NAND2_X1   g27738(.A1(new_n30174_), .A2(new_n30167_), .ZN(new_n30175_));
  NOR3_X1    g27739(.A1(new_n30058_), .A2(pi1155), .A3(new_n30088_), .ZN(new_n30176_));
  OAI21_X1   g27740(.A1(new_n30053_), .A2(new_n30081_), .B(new_n30176_), .ZN(new_n30177_));
  AOI21_X1   g27741(.A1(new_n30162_), .A2(new_n30177_), .B(pi1157), .ZN(new_n30178_));
  AOI21_X1   g27742(.A1(new_n30178_), .A2(new_n30175_), .B(pi0211), .ZN(new_n30179_));
  INV_X1     g27743(.I(new_n30173_), .ZN(new_n30180_));
  AOI21_X1   g27744(.A1(new_n30156_), .A2(new_n30180_), .B(new_n12965_), .ZN(new_n30181_));
  OAI21_X1   g27745(.A1(new_n30144_), .A2(new_n12742_), .B(new_n30181_), .ZN(new_n30182_));
  AOI21_X1   g27746(.A1(new_n30182_), .A2(new_n30179_), .B(pi0219), .ZN(new_n30183_));
  NAND2_X1   g27747(.A1(new_n30170_), .A2(new_n30183_), .ZN(new_n30184_));
  NAND3_X1   g27748(.A1(new_n30184_), .A2(new_n29997_), .A3(new_n30128_), .ZN(new_n30185_));
  AOI21_X1   g27749(.A1(new_n30185_), .A2(new_n30036_), .B(new_n29934_), .ZN(new_n30186_));
  AOI21_X1   g27750(.A1(new_n30186_), .A2(new_n30034_), .B(pi0230), .ZN(new_n30187_));
  AOI22_X1   g27751(.A1(new_n30187_), .A2(new_n29989_), .B1(pi0230), .B2(new_n29926_), .ZN(po0400));
  OAI21_X1   g27752(.A1(new_n29396_), .A2(new_n29187_), .B(new_n8811_), .ZN(new_n30189_));
  NAND2_X1   g27753(.A1(new_n29405_), .A2(new_n8809_), .ZN(new_n30190_));
  AOI21_X1   g27754(.A1(new_n30190_), .A2(new_n30189_), .B(new_n28361_), .ZN(new_n30191_));
  OAI21_X1   g27755(.A1(new_n29571_), .A2(new_n29572_), .B(new_n30191_), .ZN(new_n30192_));
  NOR2_X1    g27756(.A1(new_n28801_), .A2(new_n29581_), .ZN(new_n30193_));
  AOI21_X1   g27757(.A1(new_n30192_), .A2(new_n30193_), .B(po1038), .ZN(new_n30194_));
  AOI21_X1   g27758(.A1(new_n29420_), .A2(new_n29573_), .B(new_n29433_), .ZN(new_n30195_));
  NOR3_X1    g27759(.A1(new_n30194_), .A2(new_n26198_), .A3(new_n30195_), .ZN(new_n30196_));
  NOR3_X1    g27760(.A1(new_n28806_), .A2(pi0213), .A3(new_n28788_), .ZN(new_n30197_));
  OAI21_X1   g27761(.A1(new_n30196_), .A2(new_n30197_), .B(new_n28360_), .ZN(new_n30198_));
  NOR2_X1    g27762(.A1(new_n28784_), .A2(new_n2628_), .ZN(new_n30199_));
  NOR2_X1    g27763(.A1(new_n29335_), .A2(new_n30199_), .ZN(new_n30200_));
  NAND2_X1   g27764(.A1(new_n29353_), .A2(new_n30200_), .ZN(new_n30201_));
  AOI21_X1   g27765(.A1(new_n30201_), .A2(pi0214), .B(new_n29395_), .ZN(new_n30202_));
  AOI21_X1   g27766(.A1(new_n28064_), .A2(new_n29605_), .B(new_n8509_), .ZN(new_n30203_));
  OAI21_X1   g27767(.A1(new_n30200_), .A2(pi0214), .B(new_n30203_), .ZN(new_n30204_));
  OAI21_X1   g27768(.A1(new_n30204_), .A2(new_n29352_), .B(new_n8807_), .ZN(new_n30205_));
  NOR2_X1    g27769(.A1(new_n30202_), .A2(new_n30205_), .ZN(new_n30206_));
  INV_X1     g27770(.I(new_n29410_), .ZN(new_n30207_));
  NAND2_X1   g27771(.A1(new_n29353_), .A2(new_n28848_), .ZN(new_n30208_));
  AOI21_X1   g27772(.A1(new_n30208_), .A2(new_n8510_), .B(new_n29411_), .ZN(new_n30209_));
  OAI21_X1   g27773(.A1(new_n30209_), .A2(new_n30207_), .B(new_n29359_), .ZN(new_n30210_));
  NOR2_X1    g27774(.A1(new_n30210_), .A2(new_n30206_), .ZN(new_n30211_));
  NOR2_X1    g27775(.A1(new_n28067_), .A2(new_n8807_), .ZN(new_n30212_));
  INV_X1     g27776(.I(new_n30212_), .ZN(new_n30213_));
  NOR2_X1    g27777(.A1(new_n30213_), .A2(new_n2628_), .ZN(new_n30214_));
  NAND2_X1   g27778(.A1(new_n30200_), .A2(pi0214), .ZN(new_n30215_));
  NAND2_X1   g27779(.A1(new_n29342_), .A2(new_n8511_), .ZN(new_n30216_));
  AOI21_X1   g27780(.A1(new_n30215_), .A2(new_n30216_), .B(pi0212), .ZN(new_n30217_));
  NOR2_X1    g27781(.A1(new_n30204_), .A2(new_n29335_), .ZN(new_n30218_));
  NOR3_X1    g27782(.A1(new_n30218_), .A2(new_n30217_), .A3(pi0219), .ZN(new_n30219_));
  NOR4_X1    g27783(.A1(new_n30219_), .A2(new_n29363_), .A3(new_n29339_), .A4(new_n30214_), .ZN(new_n30220_));
  NOR4_X1    g27784(.A1(new_n30220_), .A2(new_n30211_), .A3(pi0213), .A4(new_n28788_), .ZN(new_n30221_));
  AOI21_X1   g27785(.A1(new_n29434_), .A2(new_n29421_), .B(new_n26198_), .ZN(new_n30222_));
  OAI21_X1   g27786(.A1(new_n30221_), .A2(new_n30222_), .B(pi0209), .ZN(new_n30223_));
  NAND3_X1   g27787(.A1(new_n30223_), .A2(pi0230), .A3(new_n30198_), .ZN(new_n30224_));
  OAI21_X1   g27788(.A1(pi0230), .A2(new_n5042_), .B(new_n30224_), .ZN(po0401));
  INV_X1     g27789(.I(new_n29124_), .ZN(new_n30226_));
  NOR2_X1    g27790(.A1(new_n30226_), .A2(new_n3343_), .ZN(new_n30227_));
  NOR2_X1    g27791(.A1(new_n30227_), .A2(pi1147), .ZN(new_n30228_));
  OAI21_X1   g27792(.A1(new_n29126_), .A2(new_n29327_), .B(new_n30228_), .ZN(new_n30229_));
  INV_X1     g27793(.I(new_n30229_), .ZN(new_n30230_));
  NOR2_X1    g27794(.A1(new_n29900_), .A2(new_n28503_), .ZN(new_n30231_));
  INV_X1     g27795(.I(new_n30231_), .ZN(new_n30232_));
  AOI21_X1   g27796(.A1(new_n30232_), .A2(new_n29889_), .B(po1038), .ZN(new_n30233_));
  INV_X1     g27797(.I(new_n30233_), .ZN(new_n30234_));
  NOR2_X1    g27798(.A1(new_n29396_), .A2(new_n8511_), .ZN(new_n30235_));
  NAND2_X1   g27799(.A1(new_n29901_), .A2(new_n2628_), .ZN(new_n30236_));
  AOI21_X1   g27800(.A1(new_n30236_), .A2(new_n30235_), .B(new_n8509_), .ZN(new_n30237_));
  NOR2_X1    g27801(.A1(new_n29898_), .A2(pi0299), .ZN(new_n30238_));
  NOR2_X1    g27802(.A1(new_n30238_), .A2(pi0211), .ZN(new_n30239_));
  NOR2_X1    g27803(.A1(new_n30239_), .A2(new_n29888_), .ZN(new_n30240_));
  NAND2_X1   g27804(.A1(new_n30240_), .A2(new_n8511_), .ZN(new_n30241_));
  OAI21_X1   g27805(.A1(new_n30240_), .A2(new_n29904_), .B(new_n8807_), .ZN(new_n30242_));
  AOI21_X1   g27806(.A1(new_n30237_), .A2(new_n30241_), .B(new_n30242_), .ZN(new_n30243_));
  OAI21_X1   g27807(.A1(new_n30243_), .A2(new_n30234_), .B(new_n30230_), .ZN(new_n30244_));
  NOR3_X1    g27808(.A1(new_n30227_), .A2(new_n29363_), .A3(new_n29125_), .ZN(new_n30245_));
  OAI21_X1   g27809(.A1(new_n30238_), .A2(new_n29904_), .B(new_n8807_), .ZN(new_n30246_));
  NOR2_X1    g27810(.A1(new_n29900_), .A2(new_n8510_), .ZN(new_n30247_));
  NOR3_X1    g27811(.A1(new_n30239_), .A2(new_n8511_), .A3(new_n30247_), .ZN(new_n30248_));
  NOR3_X1    g27812(.A1(new_n29898_), .A2(pi0214), .A3(pi0299), .ZN(new_n30249_));
  NOR3_X1    g27813(.A1(new_n30248_), .A2(new_n8509_), .A3(new_n30249_), .ZN(new_n30250_));
  OAI21_X1   g27814(.A1(new_n30250_), .A2(new_n30246_), .B(new_n30233_), .ZN(new_n30251_));
  AOI21_X1   g27815(.A1(new_n30251_), .A2(new_n30245_), .B(new_n29296_), .ZN(new_n30252_));
  NAND2_X1   g27816(.A1(new_n30244_), .A2(new_n30252_), .ZN(new_n30253_));
  OAI21_X1   g27817(.A1(new_n29887_), .A2(pi0212), .B(new_n8807_), .ZN(new_n30254_));
  AOI21_X1   g27818(.A1(new_n30237_), .A2(new_n29903_), .B(new_n30254_), .ZN(new_n30255_));
  OAI21_X1   g27819(.A1(new_n30255_), .A2(new_n30234_), .B(new_n30228_), .ZN(new_n30256_));
  NOR2_X1    g27820(.A1(new_n30245_), .A2(new_n29366_), .ZN(new_n30257_));
  INV_X1     g27821(.I(new_n30257_), .ZN(new_n30258_));
  NOR2_X1    g27822(.A1(new_n29888_), .A2(new_n29044_), .ZN(new_n30259_));
  OAI21_X1   g27823(.A1(new_n29904_), .A2(new_n30259_), .B(new_n8807_), .ZN(new_n30260_));
  NOR2_X1    g27824(.A1(new_n29903_), .A2(new_n29044_), .ZN(new_n30261_));
  NOR3_X1    g27825(.A1(new_n30248_), .A2(new_n8509_), .A3(new_n30261_), .ZN(new_n30262_));
  OAI21_X1   g27826(.A1(new_n30262_), .A2(new_n30260_), .B(new_n30233_), .ZN(new_n30263_));
  NAND2_X1   g27827(.A1(new_n30263_), .A2(new_n30258_), .ZN(new_n30264_));
  NAND3_X1   g27828(.A1(new_n30256_), .A2(new_n29296_), .A3(new_n30264_), .ZN(new_n30265_));
  NAND3_X1   g27829(.A1(new_n30265_), .A2(new_n30253_), .A3(pi0213), .ZN(new_n30266_));
  NAND2_X1   g27830(.A1(new_n29909_), .A2(new_n26198_), .ZN(new_n30267_));
  AOI21_X1   g27831(.A1(new_n30266_), .A2(new_n30267_), .B(pi0209), .ZN(new_n30268_));
  INV_X1     g27832(.I(new_n29885_), .ZN(new_n30269_));
  NOR3_X1    g27833(.A1(new_n8525_), .A2(pi0200), .A3(pi1146), .ZN(new_n30270_));
  NOR3_X1    g27834(.A1(new_n8523_), .A2(new_n30270_), .A3(new_n28136_), .ZN(new_n30271_));
  NOR2_X1    g27835(.A1(new_n29318_), .A2(new_n30270_), .ZN(new_n30272_));
  INV_X1     g27836(.I(new_n30272_), .ZN(new_n30273_));
  NOR2_X1    g27837(.A1(new_n30273_), .A2(new_n8522_), .ZN(new_n30274_));
  OAI21_X1   g27838(.A1(new_n30274_), .A2(pi0207), .B(new_n30271_), .ZN(new_n30275_));
  NOR2_X1    g27839(.A1(new_n28126_), .A2(new_n3343_), .ZN(new_n30276_));
  AOI22_X1   g27840(.A1(new_n30276_), .A2(pi0207), .B1(pi1146), .B2(new_n28321_), .ZN(new_n30277_));
  NAND2_X1   g27841(.A1(new_n30277_), .A2(pi0208), .ZN(new_n30278_));
  OAI21_X1   g27842(.A1(pi0208), .A2(new_n29316_), .B(new_n30278_), .ZN(new_n30279_));
  NAND2_X1   g27843(.A1(new_n30279_), .A2(new_n30275_), .ZN(new_n30280_));
  INV_X1     g27844(.I(new_n30280_), .ZN(new_n30281_));
  NOR2_X1    g27845(.A1(new_n30281_), .A2(pi0299), .ZN(new_n30282_));
  AOI21_X1   g27846(.A1(new_n30282_), .A2(new_n28503_), .B(new_n8807_), .ZN(new_n30283_));
  INV_X1     g27847(.I(new_n30283_), .ZN(new_n30284_));
  AOI21_X1   g27848(.A1(new_n30281_), .A2(new_n2628_), .B(new_n28503_), .ZN(new_n30285_));
  AOI21_X1   g27849(.A1(new_n28870_), .A2(new_n30285_), .B(new_n30284_), .ZN(new_n30286_));
  NOR3_X1    g27850(.A1(new_n30286_), .A2(pi1147), .A3(po1038), .ZN(new_n30287_));
  INV_X1     g27851(.I(new_n30282_), .ZN(new_n30288_));
  NAND2_X1   g27852(.A1(new_n29879_), .A2(pi0299), .ZN(new_n30289_));
  AOI21_X1   g27853(.A1(new_n30288_), .A2(new_n30289_), .B(new_n8509_), .ZN(new_n30290_));
  AOI21_X1   g27854(.A1(pi0214), .A2(new_n29405_), .B(new_n30282_), .ZN(new_n30291_));
  OAI21_X1   g27855(.A1(new_n30291_), .A2(pi0212), .B(new_n8807_), .ZN(new_n30292_));
  OAI21_X1   g27856(.A1(new_n30290_), .A2(new_n30292_), .B(new_n30287_), .ZN(new_n30293_));
  NOR2_X1    g27857(.A1(po1038), .A2(new_n29363_), .ZN(new_n30294_));
  INV_X1     g27858(.I(new_n30294_), .ZN(new_n30295_));
  NOR2_X1    g27859(.A1(new_n28448_), .A2(new_n30270_), .ZN(new_n30296_));
  NOR2_X1    g27860(.A1(new_n30273_), .A2(new_n8524_), .ZN(new_n30297_));
  AOI21_X1   g27861(.A1(new_n28372_), .A2(new_n30296_), .B(new_n30297_), .ZN(new_n30298_));
  INV_X1     g27862(.I(new_n30298_), .ZN(new_n30299_));
  AOI21_X1   g27863(.A1(new_n30299_), .A2(new_n28503_), .B(new_n8807_), .ZN(new_n30300_));
  AOI21_X1   g27864(.A1(new_n28041_), .A2(new_n30296_), .B(new_n30274_), .ZN(new_n30301_));
  NAND2_X1   g27865(.A1(new_n28123_), .A2(pi1146), .ZN(new_n30302_));
  AOI21_X1   g27866(.A1(new_n30302_), .A2(new_n28736_), .B(pi0299), .ZN(new_n30303_));
  AOI21_X1   g27867(.A1(new_n30303_), .A2(new_n8521_), .B(new_n29316_), .ZN(new_n30304_));
  NAND2_X1   g27868(.A1(new_n30272_), .A2(pi0207), .ZN(new_n30305_));
  AOI21_X1   g27869(.A1(new_n30305_), .A2(new_n30304_), .B(new_n8522_), .ZN(new_n30306_));
  NAND2_X1   g27870(.A1(new_n30306_), .A2(new_n2628_), .ZN(new_n30307_));
  NAND2_X1   g27871(.A1(new_n30301_), .A2(new_n30307_), .ZN(new_n30308_));
  OAI21_X1   g27872(.A1(new_n30308_), .A2(new_n28214_), .B(new_n28057_), .ZN(new_n30309_));
  AOI21_X1   g27873(.A1(new_n30309_), .A2(new_n30300_), .B(new_n30295_), .ZN(new_n30310_));
  INV_X1     g27874(.I(new_n30308_), .ZN(new_n30311_));
  AOI21_X1   g27875(.A1(new_n30311_), .A2(new_n30289_), .B(new_n8509_), .ZN(new_n30312_));
  NOR2_X1    g27876(.A1(new_n30299_), .A2(pi0214), .ZN(new_n30313_));
  NOR2_X1    g27877(.A1(new_n30313_), .A2(pi0212), .ZN(new_n30314_));
  INV_X1     g27878(.I(new_n30314_), .ZN(new_n30315_));
  NAND2_X1   g27879(.A1(new_n30311_), .A2(pi0214), .ZN(new_n30316_));
  NOR2_X1    g27880(.A1(new_n30316_), .A2(new_n29405_), .ZN(new_n30317_));
  OAI21_X1   g27881(.A1(new_n30317_), .A2(new_n30315_), .B(new_n8807_), .ZN(new_n30318_));
  OAI21_X1   g27882(.A1(new_n30318_), .A2(new_n30312_), .B(new_n30310_), .ZN(new_n30319_));
  NAND4_X1   g27883(.A1(new_n30293_), .A2(pi1148), .A3(new_n30269_), .A4(new_n30319_), .ZN(new_n30320_));
  NAND2_X1   g27884(.A1(new_n29076_), .A2(new_n8524_), .ZN(new_n30321_));
  NAND2_X1   g27885(.A1(new_n30276_), .A2(new_n30321_), .ZN(new_n30322_));
  INV_X1     g27886(.I(new_n30322_), .ZN(new_n30323_));
  AOI21_X1   g27887(.A1(new_n30323_), .A2(new_n28056_), .B(new_n8807_), .ZN(new_n30324_));
  OAI21_X1   g27888(.A1(new_n30323_), .A2(new_n8510_), .B(new_n28430_), .ZN(new_n30325_));
  NOR2_X1    g27889(.A1(new_n30276_), .A2(pi0299), .ZN(new_n30326_));
  NOR2_X1    g27890(.A1(new_n30281_), .A2(new_n30326_), .ZN(new_n30327_));
  NOR2_X1    g27891(.A1(new_n30327_), .A2(pi0299), .ZN(new_n30328_));
  NOR2_X1    g27892(.A1(new_n30328_), .A2(new_n28219_), .ZN(new_n30329_));
  NOR2_X1    g27893(.A1(new_n30329_), .A2(pi0211), .ZN(new_n30330_));
  OAI21_X1   g27894(.A1(new_n30330_), .A2(new_n30325_), .B(new_n30324_), .ZN(new_n30331_));
  INV_X1     g27895(.I(new_n30326_), .ZN(new_n30332_));
  AOI21_X1   g27896(.A1(new_n30290_), .A2(new_n30332_), .B(pi0219), .ZN(new_n30333_));
  NOR2_X1    g27897(.A1(new_n30322_), .A2(pi0214), .ZN(new_n30334_));
  NOR2_X1    g27898(.A1(new_n30328_), .A2(new_n8511_), .ZN(new_n30335_));
  INV_X1     g27899(.I(new_n30335_), .ZN(new_n30336_));
  AOI21_X1   g27900(.A1(new_n29561_), .A2(new_n30288_), .B(new_n30336_), .ZN(new_n30337_));
  OAI21_X1   g27901(.A1(new_n30337_), .A2(new_n30334_), .B(new_n8509_), .ZN(new_n30338_));
  NAND2_X1   g27902(.A1(new_n30338_), .A2(new_n30333_), .ZN(new_n30339_));
  NAND3_X1   g27903(.A1(new_n30339_), .A2(new_n29359_), .A3(new_n30331_), .ZN(new_n30340_));
  AOI21_X1   g27904(.A1(new_n28372_), .A2(new_n30303_), .B(new_n30297_), .ZN(new_n30341_));
  NOR2_X1    g27905(.A1(new_n30341_), .A2(pi0214), .ZN(new_n30342_));
  AOI21_X1   g27906(.A1(new_n30342_), .A2(new_n8509_), .B(new_n8807_), .ZN(new_n30343_));
  AOI21_X1   g27907(.A1(new_n30341_), .A2(pi0211), .B(new_n28056_), .ZN(new_n30344_));
  NAND2_X1   g27908(.A1(new_n30303_), .A2(pi0207), .ZN(new_n30345_));
  AOI21_X1   g27909(.A1(new_n30345_), .A2(new_n29317_), .B(pi0208), .ZN(new_n30346_));
  NOR2_X1    g27910(.A1(new_n30306_), .A2(new_n30346_), .ZN(new_n30347_));
  INV_X1     g27911(.I(new_n30347_), .ZN(new_n30348_));
  NOR2_X1    g27912(.A1(new_n30348_), .A2(pi0299), .ZN(new_n30349_));
  AOI21_X1   g27913(.A1(new_n30311_), .A2(new_n28223_), .B(new_n30349_), .ZN(new_n30350_));
  OAI21_X1   g27914(.A1(new_n30350_), .A2(pi0211), .B(new_n30344_), .ZN(new_n30351_));
  AOI21_X1   g27915(.A1(new_n30351_), .A2(new_n30343_), .B(new_n30295_), .ZN(new_n30352_));
  NOR2_X1    g27916(.A1(new_n30349_), .A2(new_n8511_), .ZN(new_n30353_));
  NAND2_X1   g27917(.A1(new_n30311_), .A2(new_n29561_), .ZN(new_n30354_));
  AOI21_X1   g27918(.A1(new_n30354_), .A2(new_n30353_), .B(new_n30342_), .ZN(new_n30355_));
  INV_X1     g27919(.I(new_n30349_), .ZN(new_n30356_));
  AOI21_X1   g27920(.A1(new_n30312_), .A2(new_n30356_), .B(pi0219), .ZN(new_n30357_));
  OAI21_X1   g27921(.A1(pi0212), .A2(new_n30355_), .B(new_n30357_), .ZN(new_n30358_));
  NAND2_X1   g27922(.A1(new_n30358_), .A2(new_n30352_), .ZN(new_n30359_));
  NAND4_X1   g27923(.A1(new_n30340_), .A2(new_n29296_), .A3(new_n30269_), .A4(new_n30359_), .ZN(new_n30360_));
  NAND3_X1   g27924(.A1(new_n30360_), .A2(new_n26198_), .A3(new_n30320_), .ZN(new_n30361_));
  INV_X1     g27925(.I(new_n30327_), .ZN(new_n30362_));
  OAI21_X1   g27926(.A1(new_n30362_), .A2(new_n30325_), .B(new_n30324_), .ZN(new_n30363_));
  NAND2_X1   g27927(.A1(new_n30363_), .A2(new_n6643_), .ZN(new_n30364_));
  NOR2_X1    g27928(.A1(new_n30282_), .A2(new_n29682_), .ZN(new_n30365_));
  NOR2_X1    g27929(.A1(new_n30365_), .A2(new_n30277_), .ZN(new_n30366_));
  NOR2_X1    g27930(.A1(new_n30366_), .A2(pi0219), .ZN(new_n30367_));
  OAI21_X1   g27931(.A1(new_n30367_), .A2(new_n30364_), .B(new_n30228_), .ZN(new_n30368_));
  NAND2_X1   g27932(.A1(new_n30368_), .A2(new_n29296_), .ZN(new_n30369_));
  AOI21_X1   g27933(.A1(new_n3343_), .A2(new_n28297_), .B(new_n29615_), .ZN(new_n30370_));
  INV_X1     g27934(.I(new_n30370_), .ZN(new_n30371_));
  NOR2_X1    g27935(.A1(new_n30342_), .A2(pi0212), .ZN(new_n30372_));
  INV_X1     g27936(.I(new_n30341_), .ZN(new_n30373_));
  NOR2_X1    g27937(.A1(new_n30373_), .A2(new_n29044_), .ZN(new_n30374_));
  OAI21_X1   g27938(.A1(new_n8511_), .A2(new_n30374_), .B(new_n30372_), .ZN(new_n30375_));
  INV_X1     g27939(.I(new_n30353_), .ZN(new_n30376_));
  NOR2_X1    g27940(.A1(new_n30308_), .A2(pi0299), .ZN(new_n30377_));
  INV_X1     g27941(.I(new_n30377_), .ZN(new_n30378_));
  AOI21_X1   g27942(.A1(new_n30378_), .A2(new_n8510_), .B(new_n30299_), .ZN(new_n30379_));
  OAI21_X1   g27943(.A1(new_n30379_), .A2(new_n30376_), .B(pi0212), .ZN(new_n30380_));
  NOR2_X1    g27944(.A1(new_n30374_), .A2(pi0214), .ZN(new_n30381_));
  OAI21_X1   g27945(.A1(new_n30380_), .A2(new_n30381_), .B(new_n30375_), .ZN(new_n30382_));
  NAND3_X1   g27946(.A1(new_n30382_), .A2(new_n8807_), .A3(new_n30371_), .ZN(new_n30383_));
  NAND2_X1   g27947(.A1(new_n30344_), .A2(new_n30348_), .ZN(new_n30384_));
  AOI21_X1   g27948(.A1(new_n30343_), .A2(new_n30384_), .B(po1038), .ZN(new_n30385_));
  AOI21_X1   g27949(.A1(new_n30383_), .A2(new_n30385_), .B(new_n30257_), .ZN(new_n30386_));
  NOR2_X1    g27950(.A1(new_n30323_), .A2(new_n8510_), .ZN(new_n30387_));
  AOI21_X1   g27951(.A1(new_n30328_), .A2(new_n8510_), .B(new_n30387_), .ZN(new_n30388_));
  AOI21_X1   g27952(.A1(new_n30388_), .A2(pi0214), .B(new_n30282_), .ZN(new_n30389_));
  OAI21_X1   g27953(.A1(new_n30389_), .A2(pi0212), .B(new_n8807_), .ZN(new_n30390_));
  NOR3_X1    g27954(.A1(new_n30388_), .A2(pi0214), .A3(new_n30282_), .ZN(new_n30391_));
  NOR2_X1    g27955(.A1(new_n30391_), .A2(new_n8509_), .ZN(new_n30392_));
  INV_X1     g27956(.I(new_n30392_), .ZN(new_n30393_));
  AOI21_X1   g27957(.A1(new_n30235_), .A2(new_n30288_), .B(new_n30393_), .ZN(new_n30394_));
  NAND2_X1   g27958(.A1(new_n30280_), .A2(new_n28057_), .ZN(new_n30395_));
  AOI21_X1   g27959(.A1(new_n30283_), .A2(new_n30395_), .B(po1038), .ZN(new_n30396_));
  OAI21_X1   g27960(.A1(new_n30394_), .A2(new_n30390_), .B(new_n30396_), .ZN(new_n30397_));
  NAND2_X1   g27961(.A1(new_n30397_), .A2(new_n30230_), .ZN(new_n30398_));
  INV_X1     g27962(.I(new_n30300_), .ZN(new_n30399_));
  NOR2_X1    g27963(.A1(new_n30308_), .A2(new_n29316_), .ZN(new_n30400_));
  NOR2_X1    g27964(.A1(new_n30400_), .A2(new_n28503_), .ZN(new_n30401_));
  OAI21_X1   g27965(.A1(new_n30401_), .A2(new_n30399_), .B(new_n6643_), .ZN(new_n30402_));
  AOI21_X1   g27966(.A1(new_n30378_), .A2(new_n30314_), .B(pi0219), .ZN(new_n30403_));
  INV_X1     g27967(.I(new_n30403_), .ZN(new_n30404_));
  NOR2_X1    g27968(.A1(new_n30377_), .A2(new_n8509_), .ZN(new_n30405_));
  INV_X1     g27969(.I(new_n30405_), .ZN(new_n30406_));
  AOI21_X1   g27970(.A1(new_n8512_), .A2(new_n30400_), .B(new_n30406_), .ZN(new_n30407_));
  NOR2_X1    g27971(.A1(new_n30407_), .A2(new_n30404_), .ZN(new_n30408_));
  OAI21_X1   g27972(.A1(new_n30408_), .A2(new_n30402_), .B(new_n30245_), .ZN(new_n30409_));
  NAND3_X1   g27973(.A1(new_n30398_), .A2(pi1148), .A3(new_n30409_), .ZN(new_n30410_));
  OAI21_X1   g27974(.A1(new_n30369_), .A2(new_n30386_), .B(new_n30410_), .ZN(new_n30411_));
  NAND2_X1   g27975(.A1(new_n30411_), .A2(pi0213), .ZN(new_n30412_));
  NAND3_X1   g27976(.A1(new_n30412_), .A2(pi0209), .A3(new_n30361_), .ZN(new_n30413_));
  NAND2_X1   g27977(.A1(new_n30413_), .A2(pi0230), .ZN(new_n30414_));
  OAI22_X1   g27978(.A1(new_n30414_), .A2(new_n30268_), .B1(pi0230), .B2(new_n4881_), .ZN(po0402));
  NOR2_X1    g27979(.A1(new_n29525_), .A2(pi1150), .ZN(new_n30416_));
  NOR2_X1    g27980(.A1(new_n29551_), .A2(new_n29650_), .ZN(new_n30417_));
  OAI21_X1   g27981(.A1(new_n30416_), .A2(new_n30417_), .B(pi1149), .ZN(new_n30418_));
  INV_X1     g27982(.I(new_n30418_), .ZN(new_n30419_));
  NOR3_X1    g27983(.A1(new_n29464_), .A2(pi1149), .A3(new_n29650_), .ZN(new_n30420_));
  NOR3_X1    g27984(.A1(new_n30419_), .A2(pi1148), .A3(new_n30420_), .ZN(new_n30421_));
  NOR2_X1    g27985(.A1(new_n29458_), .A2(new_n29650_), .ZN(new_n30422_));
  NOR2_X1    g27986(.A1(new_n29498_), .A2(pi1150), .ZN(new_n30423_));
  NOR2_X1    g27987(.A1(new_n30422_), .A2(new_n30423_), .ZN(new_n30424_));
  NAND2_X1   g27988(.A1(new_n29555_), .A2(pi1150), .ZN(new_n30425_));
  OAI21_X1   g27989(.A1(pi1150), .A2(new_n29531_), .B(new_n30425_), .ZN(new_n30426_));
  AOI21_X1   g27990(.A1(new_n30426_), .A2(pi1149), .B(new_n29296_), .ZN(new_n30427_));
  OAI21_X1   g27991(.A1(new_n30424_), .A2(pi1149), .B(new_n30427_), .ZN(new_n30428_));
  INV_X1     g27992(.I(new_n30428_), .ZN(new_n30429_));
  NOR2_X1    g27993(.A1(new_n30429_), .A2(new_n30421_), .ZN(new_n30430_));
  NOR2_X1    g27994(.A1(new_n30430_), .A2(new_n26198_), .ZN(new_n30431_));
  AOI21_X1   g27995(.A1(new_n29483_), .A2(new_n29774_), .B(new_n29744_), .ZN(new_n30432_));
  INV_X1     g27996(.I(new_n30432_), .ZN(new_n30433_));
  OAI21_X1   g27997(.A1(new_n29505_), .A2(new_n29736_), .B(new_n8807_), .ZN(new_n30434_));
  NAND2_X1   g27998(.A1(new_n30433_), .A2(new_n30434_), .ZN(new_n30435_));
  NOR2_X1    g27999(.A1(new_n29504_), .A2(pi1146), .ZN(new_n30436_));
  OAI21_X1   g28000(.A1(new_n30435_), .A2(new_n30436_), .B(new_n30228_), .ZN(new_n30437_));
  OAI21_X1   g28001(.A1(pi1146), .A2(new_n29522_), .B(new_n30433_), .ZN(new_n30438_));
  OAI21_X1   g28002(.A1(new_n29627_), .A2(new_n29606_), .B(new_n29521_), .ZN(new_n30439_));
  NOR2_X1    g28003(.A1(new_n30439_), .A2(new_n29504_), .ZN(new_n30440_));
  OAI21_X1   g28004(.A1(new_n30440_), .A2(new_n30438_), .B(new_n30258_), .ZN(new_n30441_));
  NAND3_X1   g28005(.A1(new_n30441_), .A2(new_n29650_), .A3(new_n30437_), .ZN(new_n30442_));
  OAI21_X1   g28006(.A1(pi0214), .A2(new_n29768_), .B(new_n29548_), .ZN(new_n30443_));
  NAND2_X1   g28007(.A1(new_n30443_), .A2(new_n8807_), .ZN(new_n30444_));
  AOI21_X1   g28008(.A1(new_n29765_), .A2(new_n29768_), .B(new_n30444_), .ZN(new_n30445_));
  NOR2_X1    g28009(.A1(new_n29623_), .A2(new_n9183_), .ZN(new_n30446_));
  AOI21_X1   g28010(.A1(pi0219), .A2(new_n29317_), .B(new_n29484_), .ZN(new_n30447_));
  NOR2_X1    g28011(.A1(new_n30446_), .A2(new_n30447_), .ZN(new_n30448_));
  NOR2_X1    g28012(.A1(new_n2628_), .A2(pi1146), .ZN(new_n30449_));
  NOR2_X1    g28013(.A1(new_n29537_), .A2(new_n30449_), .ZN(new_n30450_));
  AOI21_X1   g28014(.A1(new_n29542_), .A2(new_n29768_), .B(new_n30444_), .ZN(new_n30451_));
  INV_X1     g28015(.I(new_n30451_), .ZN(new_n30452_));
  NOR3_X1    g28016(.A1(new_n30452_), .A2(new_n29536_), .A3(new_n30450_), .ZN(new_n30453_));
  NOR3_X1    g28017(.A1(new_n30453_), .A2(new_n30445_), .A3(new_n30448_), .ZN(new_n30454_));
  NOR2_X1    g28018(.A1(new_n30454_), .A2(new_n30257_), .ZN(new_n30455_));
  NOR2_X1    g28019(.A1(new_n30455_), .A2(new_n29650_), .ZN(new_n30456_));
  INV_X1     g28020(.I(new_n29542_), .ZN(new_n30457_));
  OAI21_X1   g28021(.A1(new_n29547_), .A2(new_n30457_), .B(new_n8807_), .ZN(new_n30458_));
  NOR2_X1    g28022(.A1(new_n29770_), .A2(new_n30458_), .ZN(new_n30459_));
  NOR2_X1    g28023(.A1(new_n30459_), .A2(new_n29623_), .ZN(new_n30460_));
  OAI21_X1   g28024(.A1(new_n30454_), .A2(new_n29534_), .B(new_n30460_), .ZN(new_n30461_));
  NAND2_X1   g28025(.A1(new_n30461_), .A2(new_n30228_), .ZN(new_n30462_));
  AOI21_X1   g28026(.A1(new_n30462_), .A2(new_n30456_), .B(pi1148), .ZN(new_n30463_));
  INV_X1     g28027(.I(new_n30245_), .ZN(new_n30464_));
  NOR2_X1    g28028(.A1(new_n29529_), .A2(new_n3343_), .ZN(new_n30465_));
  NAND2_X1   g28029(.A1(new_n29609_), .A2(pi0214), .ZN(new_n30466_));
  AOI21_X1   g28030(.A1(new_n29612_), .A2(new_n30466_), .B(pi0219), .ZN(new_n30467_));
  AOI21_X1   g28031(.A1(new_n30467_), .A2(new_n29608_), .B(new_n29604_), .ZN(new_n30468_));
  NOR3_X1    g28032(.A1(new_n30464_), .A2(new_n30465_), .A3(new_n30468_), .ZN(new_n30469_));
  INV_X1     g28033(.I(new_n30447_), .ZN(new_n30470_));
  NOR2_X1    g28034(.A1(new_n29417_), .A2(pi0219), .ZN(new_n30471_));
  NOR3_X1    g28035(.A1(new_n30470_), .A2(new_n29683_), .A3(new_n30471_), .ZN(new_n30472_));
  NOR3_X1    g28036(.A1(new_n30229_), .A2(new_n29617_), .A3(new_n30472_), .ZN(new_n30473_));
  NOR3_X1    g28037(.A1(new_n30473_), .A2(new_n29650_), .A3(new_n30469_), .ZN(new_n30474_));
  NOR2_X1    g28038(.A1(new_n30230_), .A2(new_n30245_), .ZN(new_n30475_));
  AOI21_X1   g28039(.A1(new_n29053_), .A2(new_n30235_), .B(new_n29474_), .ZN(new_n30476_));
  NOR2_X1    g28040(.A1(new_n30476_), .A2(new_n29479_), .ZN(new_n30477_));
  INV_X1     g28041(.I(new_n29495_), .ZN(new_n30478_));
  OAI21_X1   g28042(.A1(new_n29054_), .A2(new_n29187_), .B(new_n29475_), .ZN(new_n30479_));
  AND2_X2    g28043(.A1(new_n30479_), .A2(new_n30478_), .Z(new_n30480_));
  OAI21_X1   g28044(.A1(new_n30480_), .A2(new_n30230_), .B(new_n30477_), .ZN(new_n30481_));
  NAND2_X1   g28045(.A1(new_n30470_), .A2(new_n29482_), .ZN(new_n30482_));
  AOI21_X1   g28046(.A1(new_n30481_), .A2(new_n30482_), .B(new_n30475_), .ZN(new_n30483_));
  OAI21_X1   g28047(.A1(new_n30483_), .A2(pi1150), .B(pi1148), .ZN(new_n30484_));
  OAI21_X1   g28048(.A1(new_n30484_), .A2(new_n30474_), .B(pi1149), .ZN(new_n30485_));
  AOI21_X1   g28049(.A1(new_n30442_), .A2(new_n30463_), .B(new_n30485_), .ZN(new_n30486_));
  NOR3_X1    g28050(.A1(new_n30227_), .A2(new_n30472_), .A3(pi1147), .ZN(new_n30487_));
  NOR2_X1    g28051(.A1(new_n30257_), .A2(new_n30447_), .ZN(new_n30488_));
  OAI22_X1   g28052(.A1(new_n30488_), .A2(new_n30487_), .B1(new_n29650_), .B2(new_n29462_), .ZN(new_n30489_));
  NOR2_X1    g28053(.A1(new_n29472_), .A2(new_n28021_), .ZN(new_n30490_));
  NOR2_X1    g28054(.A1(new_n29060_), .A2(new_n29650_), .ZN(new_n30491_));
  NOR4_X1    g28055(.A1(new_n30491_), .A2(pi0219), .A3(new_n30370_), .A4(new_n30490_), .ZN(new_n30492_));
  AOI21_X1   g28056(.A1(new_n30258_), .A2(new_n30492_), .B(pi1148), .ZN(new_n30493_));
  NAND2_X1   g28057(.A1(new_n30489_), .A2(new_n30493_), .ZN(new_n30494_));
  INV_X1     g28058(.I(new_n29599_), .ZN(new_n30495_));
  NAND2_X1   g28059(.A1(new_n30495_), .A2(new_n30470_), .ZN(new_n30496_));
  INV_X1     g28060(.I(new_n29787_), .ZN(new_n30497_));
  AOI21_X1   g28061(.A1(new_n29077_), .A2(new_n8509_), .B(pi0219), .ZN(new_n30498_));
  INV_X1     g28062(.I(new_n30498_), .ZN(new_n30499_));
  NOR2_X1    g28063(.A1(new_n29738_), .A2(new_n30499_), .ZN(new_n30500_));
  OAI21_X1   g28064(.A1(new_n29594_), .A2(new_n30497_), .B(new_n30500_), .ZN(new_n30501_));
  AOI21_X1   g28065(.A1(new_n30501_), .A2(new_n30496_), .B(new_n30464_), .ZN(new_n30502_));
  NOR2_X1    g28066(.A1(new_n29591_), .A2(new_n29446_), .ZN(new_n30503_));
  OAI21_X1   g28067(.A1(new_n29437_), .A2(pi0214), .B(pi0212), .ZN(new_n30504_));
  OAI21_X1   g28068(.A1(new_n30503_), .A2(new_n30504_), .B(new_n29442_), .ZN(new_n30505_));
  AOI21_X1   g28069(.A1(new_n30505_), .A2(new_n30496_), .B(new_n30229_), .ZN(new_n30506_));
  NOR3_X1    g28070(.A1(new_n30506_), .A2(new_n29650_), .A3(new_n30502_), .ZN(new_n30507_));
  NAND2_X1   g28071(.A1(new_n29044_), .A2(new_n3343_), .ZN(new_n30508_));
  AOI21_X1   g28072(.A1(new_n29491_), .A2(new_n30508_), .B(new_n28065_), .ZN(new_n30509_));
  OAI21_X1   g28073(.A1(new_n30509_), .A2(new_n29712_), .B(new_n8807_), .ZN(new_n30510_));
  OAI21_X1   g28074(.A1(new_n29469_), .A2(new_n29482_), .B(new_n30470_), .ZN(new_n30511_));
  AOI21_X1   g28075(.A1(new_n30510_), .A2(new_n30511_), .B(new_n30475_), .ZN(new_n30512_));
  AOI21_X1   g28076(.A1(new_n8807_), .A2(new_n29471_), .B(new_n29480_), .ZN(new_n30513_));
  OAI21_X1   g28077(.A1(new_n30513_), .A2(new_n30229_), .B(new_n29650_), .ZN(new_n30514_));
  NOR2_X1    g28078(.A1(new_n30512_), .A2(new_n30514_), .ZN(new_n30515_));
  OAI21_X1   g28079(.A1(new_n30507_), .A2(new_n30515_), .B(pi1148), .ZN(new_n30516_));
  AOI21_X1   g28080(.A1(new_n30516_), .A2(new_n30494_), .B(pi1149), .ZN(new_n30517_));
  NOR3_X1    g28081(.A1(new_n30486_), .A2(pi0213), .A3(new_n30517_), .ZN(new_n30518_));
  OAI21_X1   g28082(.A1(new_n30431_), .A2(new_n30518_), .B(pi0209), .ZN(new_n30519_));
  INV_X1     g28083(.I(new_n29365_), .ZN(new_n30520_));
  AOI21_X1   g28084(.A1(new_n30378_), .A2(new_n28057_), .B(new_n30399_), .ZN(new_n30521_));
  AOI21_X1   g28085(.A1(new_n30403_), .A2(new_n30406_), .B(new_n30521_), .ZN(new_n30522_));
  NAND3_X1   g28086(.A1(new_n30522_), .A2(new_n29680_), .A3(new_n30294_), .ZN(new_n30523_));
  AND3_X2    g28087(.A1(new_n30523_), .A2(new_n29650_), .A3(new_n30520_), .Z(new_n30524_));
  OAI21_X1   g28088(.A1(new_n30284_), .A2(new_n30285_), .B(new_n29359_), .ZN(new_n30525_));
  NOR2_X1    g28089(.A1(new_n30323_), .A2(new_n29044_), .ZN(new_n30526_));
  OAI21_X1   g28090(.A1(new_n8511_), .A2(new_n30526_), .B(new_n30288_), .ZN(new_n30527_));
  NOR4_X1    g28091(.A1(new_n30335_), .A2(new_n29044_), .A3(new_n30282_), .A4(new_n30323_), .ZN(new_n30528_));
  OAI21_X1   g28092(.A1(new_n30528_), .A2(new_n8509_), .B(new_n8807_), .ZN(new_n30529_));
  AOI21_X1   g28093(.A1(new_n8509_), .A2(new_n30527_), .B(new_n30529_), .ZN(new_n30530_));
  OAI21_X1   g28094(.A1(new_n30530_), .A2(new_n30525_), .B(new_n30524_), .ZN(new_n30531_));
  NOR3_X1    g28095(.A1(new_n30288_), .A2(new_n6165_), .A3(new_n28165_), .ZN(new_n30532_));
  NOR2_X1    g28096(.A1(pi0057), .A2(pi1147), .ZN(new_n30533_));
  NOR3_X1    g28097(.A1(new_n30280_), .A2(pi0299), .A3(new_n6165_), .ZN(new_n30534_));
  OAI21_X1   g28098(.A1(new_n30534_), .A2(new_n28095_), .B(new_n30533_), .ZN(new_n30535_));
  OAI22_X1   g28099(.A1(new_n30532_), .A2(new_n30535_), .B1(new_n2582_), .B2(new_n28165_), .ZN(new_n30536_));
  NAND2_X1   g28100(.A1(new_n28165_), .A2(new_n6165_), .ZN(new_n30537_));
  NAND3_X1   g28101(.A1(new_n30537_), .A2(new_n2582_), .A3(pi1147), .ZN(new_n30538_));
  AOI21_X1   g28102(.A1(new_n30522_), .A2(new_n5477_), .B(new_n30538_), .ZN(new_n30539_));
  OAI21_X1   g28103(.A1(new_n30536_), .A2(new_n30539_), .B(pi1150), .ZN(new_n30540_));
  NAND3_X1   g28104(.A1(new_n30531_), .A2(pi1149), .A3(new_n30540_), .ZN(new_n30541_));
  NOR2_X1    g28105(.A1(new_n30521_), .A2(new_n30295_), .ZN(new_n30542_));
  OAI21_X1   g28106(.A1(new_n30379_), .A2(new_n30315_), .B(new_n8807_), .ZN(new_n30543_));
  OAI21_X1   g28107(.A1(new_n30316_), .A2(new_n29044_), .B(pi0212), .ZN(new_n30544_));
  AOI21_X1   g28108(.A1(new_n8511_), .A2(new_n30379_), .B(new_n30544_), .ZN(new_n30545_));
  OAI21_X1   g28109(.A1(new_n30545_), .A2(new_n30543_), .B(new_n30542_), .ZN(new_n30546_));
  NAND3_X1   g28110(.A1(new_n30546_), .A2(pi1150), .A3(new_n29329_), .ZN(new_n30547_));
  NAND3_X1   g28111(.A1(new_n30288_), .A2(pi0214), .A3(new_n30526_), .ZN(new_n30548_));
  AOI21_X1   g28112(.A1(new_n30392_), .A2(new_n30548_), .B(new_n30390_), .ZN(new_n30549_));
  NOR2_X1    g28113(.A1(new_n30549_), .A2(new_n30525_), .ZN(new_n30550_));
  AOI21_X1   g28114(.A1(new_n8807_), .A2(new_n30365_), .B(new_n30525_), .ZN(new_n30551_));
  NOR3_X1    g28115(.A1(new_n30551_), .A2(pi1150), .A3(new_n29124_), .ZN(new_n30552_));
  OAI21_X1   g28116(.A1(new_n30298_), .A2(pi0212), .B(new_n8807_), .ZN(new_n30553_));
  NOR2_X1    g28117(.A1(new_n30544_), .A2(new_n30313_), .ZN(new_n30554_));
  OAI21_X1   g28118(.A1(new_n30553_), .A2(new_n30554_), .B(new_n30542_), .ZN(new_n30555_));
  AOI21_X1   g28119(.A1(new_n30552_), .A2(new_n30555_), .B(pi1149), .ZN(new_n30556_));
  OAI21_X1   g28120(.A1(new_n30550_), .A2(new_n30547_), .B(new_n30556_), .ZN(new_n30557_));
  NAND3_X1   g28121(.A1(new_n30557_), .A2(new_n30541_), .A3(pi1148), .ZN(new_n30558_));
  NOR2_X1    g28122(.A1(new_n29315_), .A2(new_n29650_), .ZN(new_n30559_));
  NOR2_X1    g28123(.A1(new_n30341_), .A2(new_n29363_), .ZN(new_n30560_));
  NOR3_X1    g28124(.A1(new_n30322_), .A2(new_n30559_), .A3(pi1147), .ZN(new_n30561_));
  OAI21_X1   g28125(.A1(new_n30560_), .A2(new_n30561_), .B(new_n6643_), .ZN(new_n30562_));
  NAND2_X1   g28126(.A1(new_n30562_), .A2(new_n29297_), .ZN(new_n30563_));
  OAI21_X1   g28127(.A1(new_n30362_), .A2(pi1147), .B(new_n12618_), .ZN(new_n30564_));
  AOI21_X1   g28128(.A1(new_n30564_), .A2(new_n30559_), .B(new_n30563_), .ZN(new_n30565_));
  NAND2_X1   g28129(.A1(new_n30323_), .A2(pi0219), .ZN(new_n30566_));
  NOR2_X1    g28130(.A1(new_n30526_), .A2(new_n8511_), .ZN(new_n30567_));
  OAI21_X1   g28131(.A1(new_n30322_), .A2(pi0214), .B(new_n8509_), .ZN(new_n30568_));
  INV_X1     g28132(.I(new_n30388_), .ZN(new_n30569_));
  OAI21_X1   g28133(.A1(new_n30569_), .A2(new_n8511_), .B(pi0212), .ZN(new_n30570_));
  NOR2_X1    g28134(.A1(new_n30526_), .A2(pi0214), .ZN(new_n30571_));
  OAI22_X1   g28135(.A1(new_n30570_), .A2(new_n30571_), .B1(new_n30567_), .B2(new_n30568_), .ZN(new_n30572_));
  OAI21_X1   g28136(.A1(new_n30572_), .A2(pi0219), .B(new_n30566_), .ZN(new_n30573_));
  NAND2_X1   g28137(.A1(new_n30373_), .A2(pi0219), .ZN(new_n30574_));
  OAI21_X1   g28138(.A1(new_n30382_), .A2(pi0219), .B(new_n30574_), .ZN(new_n30575_));
  AOI22_X1   g28139(.A1(new_n30573_), .A2(new_n29359_), .B1(new_n30294_), .B2(new_n30575_), .ZN(new_n30576_));
  NAND3_X1   g28140(.A1(new_n30576_), .A2(new_n29650_), .A3(new_n29382_), .ZN(new_n30577_));
  NAND2_X1   g28141(.A1(new_n30376_), .A2(new_n30372_), .ZN(new_n30578_));
  INV_X1     g28142(.I(new_n30380_), .ZN(new_n30579_));
  OAI21_X1   g28143(.A1(pi0214), .A2(new_n30349_), .B(new_n30579_), .ZN(new_n30580_));
  NAND3_X1   g28144(.A1(new_n30580_), .A2(new_n8807_), .A3(new_n30578_), .ZN(new_n30581_));
  AOI21_X1   g28145(.A1(new_n30581_), .A2(new_n30574_), .B(new_n29363_), .ZN(new_n30582_));
  NOR2_X1    g28146(.A1(new_n30328_), .A2(pi0214), .ZN(new_n30583_));
  OAI22_X1   g28147(.A1(new_n30570_), .A2(new_n30583_), .B1(new_n30335_), .B2(new_n30568_), .ZN(new_n30584_));
  OAI21_X1   g28148(.A1(new_n30584_), .A2(pi0219), .B(new_n30566_), .ZN(new_n30585_));
  AOI21_X1   g28149(.A1(new_n30585_), .A2(new_n29363_), .B(new_n30582_), .ZN(new_n30586_));
  NOR2_X1    g28150(.A1(new_n29125_), .A2(new_n29650_), .ZN(new_n30587_));
  OAI21_X1   g28151(.A1(new_n30586_), .A2(po1038), .B(new_n30587_), .ZN(new_n30588_));
  AOI21_X1   g28152(.A1(new_n30577_), .A2(new_n30588_), .B(new_n29297_), .ZN(new_n30589_));
  OAI21_X1   g28153(.A1(new_n30589_), .A2(new_n30565_), .B(new_n29296_), .ZN(new_n30590_));
  NAND3_X1   g28154(.A1(new_n30590_), .A2(pi0213), .A3(new_n30558_), .ZN(new_n30591_));
  NAND2_X1   g28155(.A1(new_n30411_), .A2(new_n26198_), .ZN(new_n30592_));
  NAND3_X1   g28156(.A1(new_n30591_), .A2(new_n28360_), .A3(new_n30592_), .ZN(new_n30593_));
  NAND3_X1   g28157(.A1(new_n30519_), .A2(new_n30593_), .A3(pi0230), .ZN(new_n30594_));
  OAI21_X1   g28158(.A1(pi0230), .A2(new_n4430_), .B(new_n30594_), .ZN(po0403));
  NOR2_X1    g28159(.A1(new_n30445_), .A2(new_n29623_), .ZN(new_n30596_));
  NOR2_X1    g28160(.A1(new_n30596_), .A2(new_n29365_), .ZN(new_n30597_));
  NOR2_X1    g28161(.A1(new_n29544_), .A2(new_n29625_), .ZN(new_n30598_));
  OAI21_X1   g28162(.A1(new_n30598_), .A2(new_n29623_), .B(new_n29663_), .ZN(new_n30599_));
  INV_X1     g28163(.I(new_n30599_), .ZN(new_n30600_));
  AOI21_X1   g28164(.A1(new_n30597_), .A2(new_n29035_), .B(new_n30600_), .ZN(new_n30601_));
  NAND2_X1   g28165(.A1(new_n29681_), .A2(new_n30520_), .ZN(new_n30602_));
  NOR2_X1    g28166(.A1(new_n30602_), .A2(pi1151), .ZN(new_n30603_));
  NAND2_X1   g28167(.A1(new_n29666_), .A2(pi1147), .ZN(new_n30604_));
  OAI21_X1   g28168(.A1(new_n30604_), .A2(new_n30603_), .B(pi1150), .ZN(new_n30605_));
  AOI21_X1   g28169(.A1(new_n30601_), .A2(new_n29363_), .B(new_n30605_), .ZN(new_n30606_));
  OAI21_X1   g28170(.A1(new_n29770_), .A2(new_n30458_), .B(new_n30596_), .ZN(new_n30607_));
  AND2_X2    g28171(.A1(new_n30607_), .A2(new_n29655_), .Z(new_n30608_));
  NOR2_X1    g28172(.A1(new_n30460_), .A2(new_n29328_), .ZN(new_n30609_));
  AOI21_X1   g28173(.A1(pi1151), .A2(new_n30609_), .B(new_n30608_), .ZN(new_n30610_));
  NOR2_X1    g28174(.A1(new_n29656_), .A2(new_n29684_), .ZN(new_n30611_));
  INV_X1     g28175(.I(new_n30611_), .ZN(new_n30612_));
  NOR2_X1    g28176(.A1(new_n30612_), .A2(new_n29660_), .ZN(new_n30613_));
  OAI21_X1   g28177(.A1(new_n29686_), .A2(new_n29652_), .B(pi1147), .ZN(new_n30614_));
  OAI21_X1   g28178(.A1(new_n30614_), .A2(new_n30613_), .B(new_n29650_), .ZN(new_n30615_));
  AOI21_X1   g28179(.A1(new_n30610_), .A2(new_n29363_), .B(new_n30615_), .ZN(new_n30616_));
  NOR3_X1    g28180(.A1(new_n30616_), .A2(new_n29297_), .A3(new_n30606_), .ZN(new_n30617_));
  AOI21_X1   g28181(.A1(new_n30479_), .A2(new_n29478_), .B(new_n29677_), .ZN(new_n30618_));
  NOR2_X1    g28182(.A1(new_n30618_), .A2(new_n29432_), .ZN(new_n30619_));
  INV_X1     g28183(.I(new_n30619_), .ZN(new_n30620_));
  NOR2_X1    g28184(.A1(new_n30620_), .A2(new_n29035_), .ZN(new_n30621_));
  INV_X1     g28185(.I(new_n30621_), .ZN(new_n30622_));
  AOI21_X1   g28186(.A1(new_n29482_), .A2(new_n29035_), .B(new_n29363_), .ZN(new_n30623_));
  INV_X1     g28187(.I(new_n29575_), .ZN(new_n30624_));
  NAND2_X1   g28188(.A1(new_n30624_), .A2(new_n29035_), .ZN(new_n30625_));
  NAND2_X1   g28189(.A1(new_n30625_), .A2(new_n29363_), .ZN(new_n30626_));
  NOR2_X1    g28190(.A1(new_n29503_), .A2(new_n29158_), .ZN(new_n30627_));
  NAND2_X1   g28191(.A1(new_n29776_), .A2(new_n6643_), .ZN(new_n30628_));
  OAI22_X1   g28192(.A1(new_n30628_), .A2(new_n30627_), .B1(new_n6643_), .B2(new_n29299_), .ZN(new_n30629_));
  OAI21_X1   g28193(.A1(new_n30629_), .A2(new_n30626_), .B(new_n29650_), .ZN(new_n30630_));
  AOI21_X1   g28194(.A1(new_n30622_), .A2(new_n30623_), .B(new_n30630_), .ZN(new_n30631_));
  AOI21_X1   g28195(.A1(new_n30478_), .A2(new_n8807_), .B(new_n29677_), .ZN(new_n30632_));
  OAI21_X1   g28196(.A1(new_n30632_), .A2(new_n29809_), .B(pi1147), .ZN(new_n30633_));
  NOR3_X1    g28197(.A1(new_n30618_), .A2(new_n29646_), .A3(new_n30632_), .ZN(new_n30634_));
  OAI21_X1   g28198(.A1(new_n30634_), .A2(new_n30633_), .B(pi1150), .ZN(new_n30635_));
  OAI21_X1   g28199(.A1(new_n29519_), .A2(new_n29523_), .B(new_n29645_), .ZN(new_n30636_));
  NOR2_X1    g28200(.A1(new_n29643_), .A2(pi1147), .ZN(new_n30637_));
  AOI21_X1   g28201(.A1(new_n30637_), .A2(new_n30636_), .B(new_n30635_), .ZN(new_n30638_));
  NOR3_X1    g28202(.A1(new_n30638_), .A2(pi1149), .A3(new_n30631_), .ZN(new_n30639_));
  OAI21_X1   g28203(.A1(new_n30639_), .A2(new_n30617_), .B(pi1148), .ZN(new_n30640_));
  NOR2_X1    g28204(.A1(new_n29035_), .A2(pi1147), .ZN(new_n30641_));
  AOI21_X1   g28205(.A1(new_n29461_), .A2(new_n30641_), .B(pi1150), .ZN(new_n30642_));
  NOR2_X1    g28206(.A1(new_n29482_), .A2(new_n29469_), .ZN(new_n30643_));
  OAI21_X1   g28207(.A1(new_n30643_), .A2(pi1151), .B(pi1147), .ZN(new_n30644_));
  NOR2_X1    g28208(.A1(new_n29707_), .A2(new_n29432_), .ZN(new_n30645_));
  OAI21_X1   g28209(.A1(new_n30645_), .A2(new_n30644_), .B(new_n30642_), .ZN(new_n30646_));
  NOR2_X1    g28210(.A1(new_n29477_), .A2(new_n28065_), .ZN(new_n30647_));
  NOR3_X1    g28211(.A1(new_n30647_), .A2(new_n29471_), .A3(new_n29715_), .ZN(new_n30648_));
  NOR2_X1    g28212(.A1(new_n30648_), .A2(new_n29646_), .ZN(new_n30649_));
  OAI21_X1   g28213(.A1(new_n29496_), .A2(new_n29715_), .B(new_n29382_), .ZN(new_n30650_));
  OAI21_X1   g28214(.A1(new_n30650_), .A2(pi1151), .B(pi1147), .ZN(new_n30651_));
  NOR2_X1    g28215(.A1(new_n30651_), .A2(new_n30649_), .ZN(new_n30652_));
  AOI21_X1   g28216(.A1(new_n25319_), .A2(new_n28385_), .B(new_n29035_), .ZN(new_n30653_));
  INV_X1     g28217(.I(new_n29380_), .ZN(new_n30654_));
  AOI21_X1   g28218(.A1(new_n29459_), .A2(new_n30654_), .B(pi1151), .ZN(new_n30655_));
  NOR2_X1    g28219(.A1(new_n30655_), .A2(pi1147), .ZN(new_n30656_));
  INV_X1     g28220(.I(new_n30656_), .ZN(new_n30657_));
  OAI21_X1   g28221(.A1(new_n30657_), .A2(new_n30653_), .B(pi1150), .ZN(new_n30658_));
  OAI21_X1   g28222(.A1(new_n30652_), .A2(new_n30658_), .B(new_n30646_), .ZN(new_n30659_));
  AOI21_X1   g28223(.A1(new_n30659_), .A2(new_n29297_), .B(pi1148), .ZN(new_n30660_));
  AOI21_X1   g28224(.A1(new_n29060_), .A2(new_n29683_), .B(new_n29726_), .ZN(new_n30661_));
  INV_X1     g28225(.I(new_n30661_), .ZN(new_n30662_));
  NAND2_X1   g28226(.A1(new_n30662_), .A2(new_n29655_), .ZN(new_n30663_));
  INV_X1     g28227(.I(new_n29184_), .ZN(new_n30664_));
  NOR2_X1    g28228(.A1(new_n29048_), .A2(new_n30664_), .ZN(new_n30665_));
  AOI21_X1   g28229(.A1(new_n8811_), .A2(new_n30665_), .B(new_n30661_), .ZN(new_n30666_));
  NAND2_X1   g28230(.A1(new_n30666_), .A2(new_n29651_), .ZN(new_n30667_));
  NAND3_X1   g28231(.A1(new_n30667_), .A2(new_n29363_), .A3(new_n30663_), .ZN(new_n30668_));
  NAND3_X1   g28232(.A1(new_n29720_), .A2(new_n8807_), .A3(new_n29735_), .ZN(new_n30669_));
  NAND2_X1   g28233(.A1(new_n29455_), .A2(new_n30669_), .ZN(new_n30670_));
  OAI21_X1   g28234(.A1(new_n29452_), .A2(new_n30670_), .B(new_n29655_), .ZN(new_n30671_));
  NOR2_X1    g28235(.A1(new_n29653_), .A2(new_n29363_), .ZN(new_n30672_));
  AOI21_X1   g28236(.A1(new_n30672_), .A2(new_n30671_), .B(pi1150), .ZN(new_n30673_));
  INV_X1     g28237(.I(new_n30500_), .ZN(new_n30674_));
  NOR2_X1    g28238(.A1(new_n29086_), .A2(new_n8509_), .ZN(new_n30675_));
  OAI21_X1   g28239(.A1(new_n30674_), .A2(new_n30675_), .B(new_n29455_), .ZN(new_n30676_));
  NAND2_X1   g28240(.A1(new_n30676_), .A2(new_n29663_), .ZN(new_n30677_));
  NAND2_X1   g28241(.A1(new_n30677_), .A2(pi1147), .ZN(new_n30678_));
  INV_X1     g28242(.I(new_n30678_), .ZN(new_n30679_));
  NAND2_X1   g28243(.A1(new_n30670_), .A2(new_n30520_), .ZN(new_n30680_));
  OAI21_X1   g28244(.A1(pi1151), .A2(new_n30680_), .B(new_n30679_), .ZN(new_n30681_));
  OR3_X2     g28245(.A1(new_n29740_), .A2(new_n29664_), .A3(new_n30665_), .Z(new_n30682_));
  NOR2_X1    g28246(.A1(new_n29740_), .A2(new_n29365_), .ZN(new_n30683_));
  NAND2_X1   g28247(.A1(new_n30683_), .A2(new_n29035_), .ZN(new_n30684_));
  AND2_X2    g28248(.A1(new_n30684_), .A2(new_n30682_), .Z(new_n30685_));
  AOI21_X1   g28249(.A1(new_n30685_), .A2(new_n29363_), .B(new_n29650_), .ZN(new_n30686_));
  AOI22_X1   g28250(.A1(new_n30673_), .A2(new_n30668_), .B1(new_n30681_), .B2(new_n30686_), .ZN(new_n30687_));
  OAI21_X1   g28251(.A1(new_n30687_), .A2(new_n29297_), .B(new_n30660_), .ZN(new_n30688_));
  NAND3_X1   g28252(.A1(new_n30640_), .A2(new_n30688_), .A3(pi0213), .ZN(new_n30689_));
  OR2_X2     g28253(.A1(new_n29559_), .A2(pi0213), .Z(new_n30690_));
  AOI21_X1   g28254(.A1(new_n30689_), .A2(new_n30690_), .B(pi0209), .ZN(new_n30691_));
  NOR2_X1    g28255(.A1(new_n29668_), .A2(new_n26198_), .ZN(new_n30692_));
  NOR3_X1    g28256(.A1(new_n29617_), .A2(new_n29035_), .A3(new_n29432_), .ZN(new_n30693_));
  NOR2_X1    g28257(.A1(new_n30620_), .A2(pi1151), .ZN(new_n30694_));
  NOR3_X1    g28258(.A1(new_n30694_), .A2(pi1147), .A3(new_n30693_), .ZN(new_n30695_));
  NOR2_X1    g28259(.A1(new_n29487_), .A2(new_n29328_), .ZN(new_n30696_));
  AOI21_X1   g28260(.A1(new_n30696_), .A2(new_n29035_), .B(new_n30614_), .ZN(new_n30697_));
  NOR3_X1    g28261(.A1(new_n30695_), .A2(new_n29650_), .A3(new_n30697_), .ZN(new_n30698_));
  NAND2_X1   g28262(.A1(new_n30645_), .A2(new_n29035_), .ZN(new_n30699_));
  AOI21_X1   g28263(.A1(new_n29450_), .A2(new_n29599_), .B(new_n29432_), .ZN(new_n30700_));
  NAND2_X1   g28264(.A1(new_n30700_), .A2(pi1151), .ZN(new_n30701_));
  AND3_X2    g28265(.A1(new_n30701_), .A2(new_n29363_), .A3(new_n30699_), .Z(new_n30702_));
  NOR2_X1    g28266(.A1(new_n29328_), .A2(pi1151), .ZN(new_n30703_));
  INV_X1     g28267(.I(new_n30703_), .ZN(new_n30704_));
  NOR2_X1    g28268(.A1(new_n29489_), .A2(new_n30704_), .ZN(new_n30705_));
  NOR3_X1    g28269(.A1(new_n29653_), .A2(new_n29363_), .A3(new_n30705_), .ZN(new_n30706_));
  NOR3_X1    g28270(.A1(new_n30706_), .A2(new_n30702_), .A3(pi1150), .ZN(new_n30707_));
  OAI21_X1   g28271(.A1(new_n30707_), .A2(new_n30698_), .B(pi1149), .ZN(new_n30708_));
  AOI21_X1   g28272(.A1(new_n29463_), .A2(new_n30641_), .B(pi1150), .ZN(new_n30709_));
  NAND3_X1   g28273(.A1(new_n30662_), .A2(pi1151), .A3(new_n30226_), .ZN(new_n30710_));
  NAND3_X1   g28274(.A1(new_n30710_), .A2(pi1147), .A3(new_n30612_), .ZN(new_n30711_));
  NAND2_X1   g28275(.A1(new_n30711_), .A2(new_n30709_), .ZN(new_n30712_));
  NAND3_X1   g28276(.A1(new_n30607_), .A2(pi1151), .A3(new_n30226_), .ZN(new_n30713_));
  INV_X1     g28277(.I(new_n30713_), .ZN(new_n30714_));
  NAND2_X1   g28278(.A1(new_n30435_), .A2(new_n30226_), .ZN(new_n30715_));
  OAI21_X1   g28279(.A1(new_n30715_), .A2(pi1151), .B(pi1147), .ZN(new_n30716_));
  NOR2_X1    g28280(.A1(new_n30714_), .A2(new_n30716_), .ZN(new_n30717_));
  NOR2_X1    g28281(.A1(new_n29534_), .A2(new_n29035_), .ZN(new_n30718_));
  OAI21_X1   g28282(.A1(new_n30626_), .A2(new_n30718_), .B(pi1150), .ZN(new_n30719_));
  OAI21_X1   g28283(.A1(new_n30717_), .A2(new_n30719_), .B(new_n30712_), .ZN(new_n30720_));
  AOI21_X1   g28284(.A1(new_n30720_), .A2(new_n29297_), .B(pi1148), .ZN(new_n30721_));
  NAND2_X1   g28285(.A1(new_n30597_), .A2(pi1151), .ZN(new_n30722_));
  INV_X1     g28286(.I(new_n30722_), .ZN(new_n30723_));
  NOR2_X1    g28287(.A1(new_n29511_), .A2(new_n29506_), .ZN(new_n30724_));
  OAI21_X1   g28288(.A1(new_n30432_), .A2(new_n30724_), .B(new_n30520_), .ZN(new_n30725_));
  OAI21_X1   g28289(.A1(new_n30725_), .A2(pi1151), .B(pi1147), .ZN(new_n30726_));
  NOR2_X1    g28290(.A1(new_n30723_), .A2(new_n30726_), .ZN(new_n30727_));
  NOR2_X1    g28291(.A1(new_n29381_), .A2(new_n29035_), .ZN(new_n30728_));
  OAI21_X1   g28292(.A1(new_n30451_), .A2(new_n29535_), .B(new_n30728_), .ZN(new_n30729_));
  AND2_X2    g28293(.A1(new_n30637_), .A2(new_n30729_), .Z(new_n30730_));
  NOR3_X1    g28294(.A1(new_n30730_), .A2(pi1149), .A3(new_n30727_), .ZN(new_n30731_));
  NOR4_X1    g28295(.A1(new_n29388_), .A2(pi1151), .A3(new_n29481_), .A4(new_n29528_), .ZN(new_n30732_));
  OAI21_X1   g28296(.A1(new_n30604_), .A2(new_n30732_), .B(pi1149), .ZN(new_n30733_));
  NAND2_X1   g28297(.A1(new_n29126_), .A2(new_n29035_), .ZN(new_n30734_));
  NOR3_X1    g28298(.A1(new_n30618_), .A2(new_n30632_), .A3(new_n30734_), .ZN(new_n30735_));
  NOR2_X1    g28299(.A1(new_n30468_), .A2(new_n29646_), .ZN(new_n30736_));
  NOR3_X1    g28300(.A1(new_n30735_), .A2(pi1147), .A3(new_n30736_), .ZN(new_n30737_));
  OAI21_X1   g28301(.A1(new_n30737_), .A2(new_n30733_), .B(pi1150), .ZN(new_n30738_));
  AOI21_X1   g28302(.A1(new_n29786_), .A2(new_n29787_), .B(new_n30674_), .ZN(new_n30739_));
  OAI21_X1   g28303(.A1(new_n30739_), .A2(new_n30495_), .B(new_n29126_), .ZN(new_n30740_));
  NOR2_X1    g28304(.A1(new_n30648_), .A2(new_n30734_), .ZN(new_n30741_));
  INV_X1     g28305(.I(new_n30741_), .ZN(new_n30742_));
  OAI21_X1   g28306(.A1(new_n30740_), .A2(new_n29035_), .B(new_n30742_), .ZN(new_n30743_));
  NOR2_X1    g28307(.A1(new_n30743_), .A2(pi1147), .ZN(new_n30744_));
  NOR4_X1    g28308(.A1(new_n29489_), .A2(pi1151), .A3(new_n29388_), .A4(new_n30648_), .ZN(new_n30745_));
  OAI21_X1   g28309(.A1(new_n30678_), .A2(new_n30745_), .B(pi1149), .ZN(new_n30746_));
  OR2_X2     g28310(.A1(new_n29530_), .A2(pi1151), .Z(new_n30747_));
  AOI21_X1   g28311(.A1(new_n30683_), .A2(pi1151), .B(new_n29363_), .ZN(new_n30748_));
  AOI21_X1   g28312(.A1(new_n30748_), .A2(new_n30747_), .B(pi1149), .ZN(new_n30749_));
  INV_X1     g28313(.I(new_n30728_), .ZN(new_n30750_));
  NOR2_X1    g28314(.A1(new_n29801_), .A2(new_n30664_), .ZN(new_n30751_));
  OAI21_X1   g28315(.A1(new_n30751_), .A2(new_n30750_), .B(new_n30656_), .ZN(new_n30752_));
  AOI21_X1   g28316(.A1(new_n30749_), .A2(new_n30752_), .B(pi1150), .ZN(new_n30753_));
  OAI21_X1   g28317(.A1(new_n30746_), .A2(new_n30744_), .B(new_n30753_), .ZN(new_n30754_));
  OAI21_X1   g28318(.A1(new_n30731_), .A2(new_n30738_), .B(new_n30754_), .ZN(new_n30755_));
  AOI22_X1   g28319(.A1(new_n30755_), .A2(pi1148), .B1(new_n30708_), .B2(new_n30721_), .ZN(new_n30756_));
  AOI21_X1   g28320(.A1(new_n30756_), .A2(new_n26198_), .B(new_n30692_), .ZN(new_n30757_));
  OAI21_X1   g28321(.A1(new_n30757_), .A2(new_n28360_), .B(pi0230), .ZN(new_n30758_));
  OAI22_X1   g28322(.A1(new_n30758_), .A2(new_n30691_), .B1(pi0230), .B2(new_n4339_), .ZN(po0404));
  NAND4_X1   g28323(.A1(new_n29459_), .A2(new_n30654_), .A3(pi1151), .A4(new_n28422_), .ZN(new_n30760_));
  NOR2_X1    g28324(.A1(new_n29461_), .A2(pi1151), .ZN(new_n30761_));
  OR3_X2     g28325(.A1(new_n30761_), .A2(new_n28422_), .A3(new_n30653_), .Z(new_n30762_));
  NAND3_X1   g28326(.A1(new_n30762_), .A2(new_n29650_), .A3(new_n30760_), .ZN(new_n30763_));
  NAND2_X1   g28327(.A1(new_n30683_), .A2(pi1151), .ZN(new_n30764_));
  NAND3_X1   g28328(.A1(new_n30764_), .A2(new_n30663_), .A3(new_n28422_), .ZN(new_n30765_));
  NAND2_X1   g28329(.A1(new_n30666_), .A2(new_n30703_), .ZN(new_n30766_));
  NAND3_X1   g28330(.A1(new_n30766_), .A2(pi1152), .A3(new_n30682_), .ZN(new_n30767_));
  NAND3_X1   g28331(.A1(new_n30767_), .A2(pi1150), .A3(new_n30765_), .ZN(new_n30768_));
  NAND3_X1   g28332(.A1(new_n30768_), .A2(new_n29297_), .A3(new_n30763_), .ZN(new_n30769_));
  NAND2_X1   g28333(.A1(new_n30609_), .A2(new_n29035_), .ZN(new_n30770_));
  NAND3_X1   g28334(.A1(new_n30770_), .A2(pi1152), .A3(new_n30599_), .ZN(new_n30771_));
  NOR2_X1    g28335(.A1(new_n30608_), .A2(new_n30723_), .ZN(new_n30772_));
  AOI21_X1   g28336(.A1(new_n30772_), .A2(new_n28422_), .B(new_n29650_), .ZN(new_n30773_));
  AOI21_X1   g28337(.A1(new_n30773_), .A2(new_n30771_), .B(new_n29297_), .ZN(new_n30774_));
  OAI21_X1   g28338(.A1(new_n29524_), .A2(new_n30750_), .B(new_n28422_), .ZN(new_n30775_));
  INV_X1     g28339(.I(new_n30775_), .ZN(new_n30776_));
  AOI21_X1   g28340(.A1(new_n30629_), .A2(new_n29035_), .B(new_n28422_), .ZN(new_n30777_));
  AOI22_X1   g28341(.A1(new_n30776_), .A2(new_n30625_), .B1(new_n30636_), .B2(new_n30777_), .ZN(new_n30778_));
  NAND2_X1   g28342(.A1(new_n30778_), .A2(new_n29650_), .ZN(new_n30779_));
  AOI21_X1   g28343(.A1(new_n30779_), .A2(new_n30774_), .B(pi1148), .ZN(new_n30780_));
  NOR2_X1    g28344(.A1(new_n30632_), .A2(new_n30750_), .ZN(new_n30781_));
  OAI21_X1   g28345(.A1(new_n30781_), .A2(new_n29696_), .B(new_n29650_), .ZN(new_n30782_));
  NOR3_X1    g28346(.A1(new_n30694_), .A2(new_n28422_), .A3(new_n30634_), .ZN(new_n30783_));
  NOR2_X1    g28347(.A1(new_n30783_), .A2(new_n30782_), .ZN(new_n30784_));
  NOR2_X1    g28348(.A1(new_n30602_), .A2(new_n29035_), .ZN(new_n30785_));
  OAI21_X1   g28349(.A1(new_n30612_), .A2(new_n29660_), .B(new_n28422_), .ZN(new_n30786_));
  OAI21_X1   g28350(.A1(new_n30786_), .A2(new_n30785_), .B(pi1150), .ZN(new_n30787_));
  NOR2_X1    g28351(.A1(new_n29665_), .A2(new_n28422_), .ZN(new_n30788_));
  INV_X1     g28352(.I(new_n30788_), .ZN(new_n30789_));
  AOI21_X1   g28353(.A1(new_n29685_), .A2(new_n30703_), .B(new_n30789_), .ZN(new_n30790_));
  OAI21_X1   g28354(.A1(new_n30790_), .A2(new_n30787_), .B(pi1149), .ZN(new_n30791_));
  OAI21_X1   g28355(.A1(new_n30784_), .A2(new_n30791_), .B(pi1148), .ZN(new_n30792_));
  NAND3_X1   g28356(.A1(new_n30670_), .A2(pi1151), .A3(new_n30520_), .ZN(new_n30793_));
  NAND3_X1   g28357(.A1(new_n30671_), .A2(new_n28422_), .A3(new_n30793_), .ZN(new_n30794_));
  NOR2_X1    g28358(.A1(new_n29457_), .A2(new_n30704_), .ZN(new_n30795_));
  NOR2_X1    g28359(.A1(new_n30795_), .A2(new_n28422_), .ZN(new_n30796_));
  AOI21_X1   g28360(.A1(new_n30796_), .A2(new_n30677_), .B(new_n29650_), .ZN(new_n30797_));
  INV_X1     g28361(.I(new_n30699_), .ZN(new_n30798_));
  OAI21_X1   g28362(.A1(new_n30648_), .A2(new_n29646_), .B(pi1152), .ZN(new_n30799_));
  OAI21_X1   g28363(.A1(new_n30799_), .A2(new_n30798_), .B(new_n29650_), .ZN(new_n30800_));
  NOR2_X1    g28364(.A1(new_n30643_), .A2(pi1151), .ZN(new_n30801_));
  NOR2_X1    g28365(.A1(new_n30650_), .A2(new_n29035_), .ZN(new_n30802_));
  NOR3_X1    g28366(.A1(new_n30802_), .A2(pi1152), .A3(new_n30801_), .ZN(new_n30803_));
  OAI21_X1   g28367(.A1(new_n30803_), .A2(new_n30800_), .B(new_n29297_), .ZN(new_n30804_));
  AOI21_X1   g28368(.A1(new_n30797_), .A2(new_n30794_), .B(new_n30804_), .ZN(new_n30805_));
  OAI21_X1   g28369(.A1(new_n30805_), .A2(new_n30792_), .B(pi0213), .ZN(new_n30806_));
  AOI21_X1   g28370(.A1(new_n30780_), .A2(new_n30769_), .B(new_n30806_), .ZN(new_n30807_));
  NOR3_X1    g28371(.A1(new_n30429_), .A2(pi0213), .A3(new_n30421_), .ZN(new_n30808_));
  NOR3_X1    g28372(.A1(new_n30807_), .A2(pi0209), .A3(new_n30808_), .ZN(new_n30809_));
  AOI21_X1   g28373(.A1(new_n29531_), .A2(pi1151), .B(pi1152), .ZN(new_n30810_));
  NAND2_X1   g28374(.A1(new_n29657_), .A2(new_n30810_), .ZN(new_n30811_));
  NOR2_X1    g28375(.A1(new_n30795_), .A2(new_n30789_), .ZN(new_n30812_));
  NOR2_X1    g28376(.A1(new_n30812_), .A2(new_n29650_), .ZN(new_n30813_));
  NAND3_X1   g28377(.A1(new_n29642_), .A2(pi1151), .A3(new_n28422_), .ZN(new_n30814_));
  AOI21_X1   g28378(.A1(new_n30761_), .A2(new_n29462_), .B(new_n28422_), .ZN(new_n30815_));
  AOI21_X1   g28379(.A1(new_n29648_), .A2(new_n30815_), .B(pi1150), .ZN(new_n30816_));
  AOI22_X1   g28380(.A1(new_n30813_), .A2(new_n30811_), .B1(new_n30814_), .B2(new_n30816_), .ZN(new_n30817_));
  NOR2_X1    g28381(.A1(new_n30817_), .A2(new_n26198_), .ZN(new_n30818_));
  NOR2_X1    g28382(.A1(new_n29463_), .A2(pi1151), .ZN(new_n30819_));
  NOR3_X1    g28383(.A1(new_n30819_), .A2(new_n28422_), .A3(new_n30718_), .ZN(new_n30820_));
  NOR3_X1    g28384(.A1(new_n30624_), .A2(new_n29035_), .A3(pi1152), .ZN(new_n30821_));
  NOR3_X1    g28385(.A1(new_n30821_), .A2(pi1150), .A3(new_n30820_), .ZN(new_n30822_));
  INV_X1     g28386(.I(new_n30693_), .ZN(new_n30823_));
  AOI21_X1   g28387(.A1(new_n30700_), .A2(new_n29035_), .B(new_n28422_), .ZN(new_n30824_));
  NAND3_X1   g28388(.A1(new_n30622_), .A2(new_n28422_), .A3(new_n30699_), .ZN(new_n30825_));
  NAND2_X1   g28389(.A1(new_n30825_), .A2(pi1150), .ZN(new_n30826_));
  AOI21_X1   g28390(.A1(new_n30823_), .A2(new_n30824_), .B(new_n30826_), .ZN(new_n30827_));
  OAI21_X1   g28391(.A1(new_n30827_), .A2(new_n30822_), .B(new_n29296_), .ZN(new_n30828_));
  OAI21_X1   g28392(.A1(new_n30715_), .A2(new_n29035_), .B(new_n30612_), .ZN(new_n30829_));
  NAND2_X1   g28393(.A1(new_n30829_), .A2(new_n28422_), .ZN(new_n30830_));
  NAND2_X1   g28394(.A1(new_n30713_), .A2(new_n30663_), .ZN(new_n30831_));
  AOI21_X1   g28395(.A1(new_n30831_), .A2(pi1152), .B(pi1150), .ZN(new_n30832_));
  AOI21_X1   g28396(.A1(new_n30832_), .A2(new_n30830_), .B(new_n29296_), .ZN(new_n30833_));
  NOR3_X1    g28397(.A1(new_n29487_), .A2(new_n29035_), .A3(new_n29328_), .ZN(new_n30834_));
  NOR3_X1    g28398(.A1(new_n30705_), .A2(new_n30834_), .A3(pi1152), .ZN(new_n30835_));
  INV_X1     g28399(.I(new_n30796_), .ZN(new_n30836_));
  AOI21_X1   g28400(.A1(new_n29651_), .A2(new_n29685_), .B(new_n30836_), .ZN(new_n30837_));
  OAI21_X1   g28401(.A1(new_n30837_), .A2(new_n30835_), .B(pi1150), .ZN(new_n30838_));
  AOI21_X1   g28402(.A1(new_n30838_), .A2(new_n30833_), .B(pi1149), .ZN(new_n30839_));
  NOR2_X1    g28403(.A1(new_n30751_), .A2(new_n29809_), .ZN(new_n30840_));
  NOR2_X1    g28404(.A1(new_n30840_), .A2(new_n28422_), .ZN(new_n30841_));
  AOI21_X1   g28405(.A1(new_n30841_), .A2(new_n30729_), .B(pi1150), .ZN(new_n30842_));
  OAI21_X1   g28406(.A1(new_n30775_), .A2(new_n30655_), .B(new_n30842_), .ZN(new_n30843_));
  OAI21_X1   g28407(.A1(new_n30740_), .A2(pi1151), .B(pi1152), .ZN(new_n30844_));
  NOR2_X1    g28408(.A1(new_n30634_), .A2(pi1152), .ZN(new_n30845_));
  AOI21_X1   g28409(.A1(new_n30845_), .A2(new_n30742_), .B(new_n29650_), .ZN(new_n30846_));
  OAI21_X1   g28410(.A1(new_n30736_), .A2(new_n30844_), .B(new_n30846_), .ZN(new_n30847_));
  NAND3_X1   g28411(.A1(new_n30843_), .A2(new_n29296_), .A3(new_n30847_), .ZN(new_n30848_));
  OR2_X2     g28412(.A1(new_n30725_), .A2(new_n29035_), .Z(new_n30849_));
  NAND3_X1   g28413(.A1(new_n30849_), .A2(new_n28422_), .A3(new_n30747_), .ZN(new_n30850_));
  NAND3_X1   g28414(.A1(new_n30722_), .A2(pi1152), .A3(new_n30684_), .ZN(new_n30851_));
  NAND3_X1   g28415(.A1(new_n30851_), .A2(new_n29650_), .A3(new_n30850_), .ZN(new_n30852_));
  NAND3_X1   g28416(.A1(new_n29554_), .A2(pi1151), .A3(new_n29482_), .ZN(new_n30853_));
  NOR2_X1    g28417(.A1(new_n30745_), .A2(pi1152), .ZN(new_n30854_));
  NAND2_X1   g28418(.A1(new_n30854_), .A2(new_n30853_), .ZN(new_n30855_));
  NOR2_X1    g28419(.A1(new_n29388_), .A2(pi1151), .ZN(new_n30856_));
  NAND2_X1   g28420(.A1(new_n30676_), .A2(new_n30856_), .ZN(new_n30857_));
  NAND2_X1   g28421(.A1(new_n30857_), .A2(new_n30788_), .ZN(new_n30858_));
  NAND3_X1   g28422(.A1(new_n30855_), .A2(pi1150), .A3(new_n30858_), .ZN(new_n30859_));
  NAND3_X1   g28423(.A1(new_n30859_), .A2(pi1148), .A3(new_n30852_), .ZN(new_n30860_));
  NAND2_X1   g28424(.A1(new_n30860_), .A2(new_n30848_), .ZN(new_n30861_));
  AOI22_X1   g28425(.A1(new_n30839_), .A2(new_n30828_), .B1(pi1149), .B2(new_n30861_), .ZN(new_n30862_));
  AOI21_X1   g28426(.A1(new_n30862_), .A2(new_n26198_), .B(new_n30818_), .ZN(new_n30863_));
  OAI21_X1   g28427(.A1(new_n30863_), .A2(new_n28360_), .B(pi0230), .ZN(new_n30864_));
  OAI22_X1   g28428(.A1(new_n30864_), .A2(new_n30809_), .B1(pi0230), .B2(new_n4105_), .ZN(po0405));
  OAI21_X1   g28429(.A1(new_n28500_), .A2(new_n28421_), .B(pi0213), .ZN(new_n30866_));
  OR2_X2     g28430(.A1(new_n28459_), .A2(new_n29159_), .Z(new_n30867_));
  NAND2_X1   g28431(.A1(new_n28460_), .A2(new_n29159_), .ZN(new_n30868_));
  AOI21_X1   g28432(.A1(new_n30867_), .A2(new_n30868_), .B(po1038), .ZN(new_n30869_));
  NOR3_X1    g28433(.A1(new_n30869_), .A2(pi1151), .A3(new_n29432_), .ZN(new_n30870_));
  AOI21_X1   g28434(.A1(new_n28457_), .A2(pi0219), .B(po1038), .ZN(new_n30871_));
  INV_X1     g28435(.I(new_n28447_), .ZN(new_n30872_));
  OAI21_X1   g28436(.A1(new_n30872_), .A2(new_n8511_), .B(new_n28491_), .ZN(new_n30873_));
  AOI21_X1   g28437(.A1(new_n30873_), .A2(new_n8509_), .B(pi0219), .ZN(new_n30874_));
  NOR2_X1    g28438(.A1(new_n28459_), .A2(new_n8511_), .ZN(new_n30875_));
  AOI21_X1   g28439(.A1(new_n8511_), .A2(new_n28447_), .B(new_n30875_), .ZN(new_n30876_));
  OAI21_X1   g28440(.A1(new_n30876_), .A2(new_n8509_), .B(new_n30874_), .ZN(new_n30877_));
  AOI21_X1   g28441(.A1(new_n30877_), .A2(new_n30871_), .B(new_n29646_), .ZN(new_n30878_));
  NOR3_X1    g28442(.A1(new_n30878_), .A2(new_n28422_), .A3(new_n30870_), .ZN(new_n30879_));
  OAI21_X1   g28443(.A1(new_n28384_), .A2(po1038), .B(new_n29035_), .ZN(new_n30880_));
  NAND2_X1   g28444(.A1(new_n30880_), .A2(new_n28422_), .ZN(new_n30881_));
  NAND2_X1   g28445(.A1(new_n28739_), .A2(new_n28097_), .ZN(new_n30882_));
  AOI21_X1   g28446(.A1(new_n28404_), .A2(new_n28580_), .B(new_n8522_), .ZN(new_n30883_));
  NAND2_X1   g28447(.A1(new_n28738_), .A2(new_n8521_), .ZN(new_n30884_));
  NAND2_X1   g28448(.A1(new_n30884_), .A2(new_n30883_), .ZN(new_n30885_));
  NAND2_X1   g28449(.A1(new_n30882_), .A2(new_n30885_), .ZN(new_n30886_));
  NAND2_X1   g28450(.A1(new_n28384_), .A2(new_n8513_), .ZN(new_n30887_));
  OAI21_X1   g28451(.A1(new_n8513_), .A2(new_n30886_), .B(new_n30887_), .ZN(new_n30888_));
  OAI21_X1   g28452(.A1(new_n30888_), .A2(pi0212), .B(new_n8807_), .ZN(new_n30889_));
  INV_X1     g28453(.I(new_n28530_), .ZN(new_n30890_));
  OAI21_X1   g28454(.A1(new_n8510_), .A2(new_n30886_), .B(new_n30890_), .ZN(new_n30891_));
  AOI21_X1   g28455(.A1(new_n30891_), .A2(new_n8511_), .B(new_n8509_), .ZN(new_n30892_));
  INV_X1     g28456(.I(new_n30892_), .ZN(new_n30893_));
  AOI21_X1   g28457(.A1(new_n8510_), .A2(new_n30886_), .B(new_n28526_), .ZN(new_n30894_));
  AOI21_X1   g28458(.A1(pi0214), .A2(new_n30894_), .B(new_n30893_), .ZN(new_n30895_));
  AOI21_X1   g28459(.A1(new_n28384_), .A2(pi0219), .B(po1038), .ZN(new_n30896_));
  OAI21_X1   g28460(.A1(new_n30895_), .A2(new_n30889_), .B(new_n30896_), .ZN(new_n30897_));
  AOI21_X1   g28461(.A1(new_n30897_), .A2(new_n30728_), .B(new_n30881_), .ZN(new_n30898_));
  NOR3_X1    g28462(.A1(new_n30879_), .A2(pi1150), .A3(new_n30898_), .ZN(new_n30899_));
  NAND3_X1   g28463(.A1(new_n30882_), .A2(new_n30885_), .A3(pi0214), .ZN(new_n30900_));
  AOI21_X1   g28464(.A1(new_n30892_), .A2(new_n30900_), .B(new_n30889_), .ZN(new_n30901_));
  OAI21_X1   g28465(.A1(new_n30894_), .A2(new_n28056_), .B(new_n28528_), .ZN(new_n30902_));
  OAI21_X1   g28466(.A1(new_n30902_), .A2(new_n8807_), .B(new_n6643_), .ZN(new_n30903_));
  OAI21_X1   g28467(.A1(new_n30901_), .A2(new_n30903_), .B(pi1151), .ZN(new_n30904_));
  NAND2_X1   g28468(.A1(new_n30888_), .A2(pi0212), .ZN(new_n30905_));
  NAND2_X1   g28469(.A1(new_n28384_), .A2(new_n8509_), .ZN(new_n30906_));
  AOI21_X1   g28470(.A1(new_n30905_), .A2(new_n30906_), .B(pi0219), .ZN(new_n30907_));
  NOR2_X1    g28471(.A1(new_n30903_), .A2(new_n30907_), .ZN(new_n30908_));
  OAI22_X1   g28472(.A1(new_n30904_), .A2(new_n29365_), .B1(new_n29656_), .B2(new_n30908_), .ZN(new_n30909_));
  NOR2_X1    g28473(.A1(new_n30909_), .A2(pi1152), .ZN(new_n30910_));
  NAND2_X1   g28474(.A1(new_n30872_), .A2(new_n28297_), .ZN(new_n30911_));
  NAND2_X1   g28475(.A1(new_n28457_), .A2(new_n28298_), .ZN(new_n30912_));
  AOI21_X1   g28476(.A1(new_n30911_), .A2(new_n30912_), .B(new_n8509_), .ZN(new_n30913_));
  NOR3_X1    g28477(.A1(new_n30875_), .A2(pi0212), .A3(new_n28490_), .ZN(new_n30914_));
  OAI21_X1   g28478(.A1(new_n30914_), .A2(new_n30913_), .B(new_n8807_), .ZN(new_n30915_));
  AOI21_X1   g28479(.A1(new_n30915_), .A2(new_n28464_), .B(new_n30704_), .ZN(new_n30916_));
  NAND2_X1   g28480(.A1(new_n28447_), .A2(pi0212), .ZN(new_n30917_));
  AOI21_X1   g28481(.A1(new_n30874_), .A2(new_n30917_), .B(new_n28463_), .ZN(new_n30918_));
  OAI21_X1   g28482(.A1(new_n30918_), .A2(new_n29664_), .B(pi1152), .ZN(new_n30919_));
  OAI21_X1   g28483(.A1(new_n30919_), .A2(new_n30916_), .B(pi1150), .ZN(new_n30920_));
  NOR2_X1    g28484(.A1(new_n30920_), .A2(new_n30910_), .ZN(new_n30921_));
  OAI21_X1   g28485(.A1(new_n30899_), .A2(new_n30921_), .B(new_n26198_), .ZN(new_n30922_));
  AOI21_X1   g28486(.A1(new_n30866_), .A2(new_n30922_), .B(new_n28360_), .ZN(new_n30923_));
  NOR2_X1    g28487(.A1(new_n30817_), .A2(pi0213), .ZN(new_n30924_));
  NOR2_X1    g28488(.A1(new_n28364_), .A2(new_n2628_), .ZN(new_n30925_));
  NAND2_X1   g28489(.A1(new_n30925_), .A2(new_n8811_), .ZN(new_n30926_));
  NAND2_X1   g28490(.A1(new_n30926_), .A2(new_n29014_), .ZN(new_n30927_));
  NAND3_X1   g28491(.A1(new_n30927_), .A2(new_n28365_), .A3(new_n29007_), .ZN(new_n30928_));
  INV_X1     g28492(.I(new_n30928_), .ZN(new_n30929_));
  NOR2_X1    g28493(.A1(new_n28669_), .A2(new_n28000_), .ZN(new_n30930_));
  AOI22_X1   g28494(.A1(new_n29775_), .A2(new_n8809_), .B1(new_n29503_), .B2(new_n30930_), .ZN(new_n30931_));
  NAND3_X1   g28495(.A1(new_n29774_), .A2(pi0211), .A3(new_n28580_), .ZN(new_n30932_));
  NAND2_X1   g28496(.A1(new_n29514_), .A2(new_n28395_), .ZN(new_n30933_));
  NAND3_X1   g28497(.A1(new_n30933_), .A2(new_n30932_), .A3(new_n28669_), .ZN(new_n30934_));
  NAND2_X1   g28498(.A1(new_n30931_), .A2(new_n30934_), .ZN(new_n30935_));
  AOI21_X1   g28499(.A1(new_n30935_), .A2(new_n8807_), .B(new_n29035_), .ZN(new_n30936_));
  AOI21_X1   g28500(.A1(new_n30936_), .A2(new_n29744_), .B(new_n30929_), .ZN(new_n30937_));
  NAND2_X1   g28501(.A1(new_n30661_), .A2(new_n29035_), .ZN(new_n30938_));
  NAND3_X1   g28502(.A1(new_n30938_), .A2(new_n28428_), .A3(new_n30928_), .ZN(new_n30939_));
  NOR2_X1    g28503(.A1(new_n28363_), .A2(new_n2628_), .ZN(new_n30940_));
  AOI21_X1   g28504(.A1(new_n29009_), .A2(new_n8509_), .B(pi0219), .ZN(new_n30941_));
  OAI21_X1   g28505(.A1(new_n29737_), .A2(new_n30940_), .B(new_n30941_), .ZN(new_n30942_));
  OAI21_X1   g28506(.A1(new_n29765_), .A2(new_n30925_), .B(pi0212), .ZN(new_n30943_));
  AOI21_X1   g28507(.A1(new_n29756_), .A2(pi0214), .B(new_n30943_), .ZN(new_n30944_));
  OAI21_X1   g28508(.A1(new_n30944_), .A2(new_n30942_), .B(new_n29622_), .ZN(new_n30945_));
  NOR2_X1    g28509(.A1(new_n30945_), .A2(new_n29037_), .ZN(new_n30946_));
  OAI21_X1   g28510(.A1(new_n30939_), .A2(new_n30946_), .B(new_n29650_), .ZN(new_n30947_));
  AOI21_X1   g28511(.A1(new_n28368_), .A2(new_n30937_), .B(new_n30947_), .ZN(new_n30948_));
  INV_X1     g28512(.I(new_n29679_), .ZN(new_n30949_));
  AOI21_X1   g28513(.A1(new_n30926_), .A2(new_n28425_), .B(new_n29527_), .ZN(new_n30950_));
  AOI21_X1   g28514(.A1(new_n29486_), .A2(new_n29604_), .B(new_n29035_), .ZN(new_n30951_));
  OAI21_X1   g28515(.A1(new_n30949_), .A2(new_n30950_), .B(new_n30951_), .ZN(new_n30952_));
  NOR2_X1    g28516(.A1(new_n29737_), .A2(new_n30940_), .ZN(new_n30953_));
  NOR2_X1    g28517(.A1(new_n30953_), .A2(new_n30499_), .ZN(new_n30954_));
  OAI21_X1   g28518(.A1(new_n29086_), .A2(new_n28581_), .B(pi0214), .ZN(new_n30955_));
  OAI21_X1   g28519(.A1(new_n29086_), .A2(new_n30940_), .B(new_n8511_), .ZN(new_n30956_));
  NAND3_X1   g28520(.A1(new_n30955_), .A2(new_n30956_), .A3(pi0212), .ZN(new_n30957_));
  AOI21_X1   g28521(.A1(new_n30957_), .A2(new_n30954_), .B(pi1151), .ZN(new_n30958_));
  AOI21_X1   g28522(.A1(new_n29455_), .A2(new_n30958_), .B(new_n28429_), .ZN(new_n30959_));
  AOI21_X1   g28523(.A1(new_n30959_), .A2(new_n30952_), .B(new_n29650_), .ZN(new_n30960_));
  NOR2_X1    g28524(.A1(new_n29470_), .A2(new_n8807_), .ZN(new_n30961_));
  NOR2_X1    g28525(.A1(new_n29471_), .A2(new_n30940_), .ZN(new_n30962_));
  NAND2_X1   g28526(.A1(new_n30962_), .A2(new_n8511_), .ZN(new_n30963_));
  NOR2_X1    g28527(.A1(new_n29470_), .A2(new_n29187_), .ZN(new_n30964_));
  OR3_X2     g28528(.A1(new_n30964_), .A2(new_n8511_), .A3(new_n29705_), .Z(new_n30965_));
  NAND3_X1   g28529(.A1(new_n30963_), .A2(new_n30965_), .A3(pi0212), .ZN(new_n30966_));
  NAND2_X1   g28530(.A1(new_n30962_), .A2(new_n29063_), .ZN(new_n30967_));
  NAND2_X1   g28531(.A1(new_n30967_), .A2(new_n8509_), .ZN(new_n30968_));
  AOI21_X1   g28532(.A1(new_n30966_), .A2(new_n30968_), .B(pi0219), .ZN(new_n30969_));
  NOR3_X1    g28533(.A1(new_n30969_), .A2(new_n6165_), .A3(new_n30961_), .ZN(new_n30970_));
  NAND2_X1   g28534(.A1(new_n28367_), .A2(new_n6165_), .ZN(new_n30971_));
  INV_X1     g28535(.I(new_n30971_), .ZN(new_n30972_));
  NOR4_X1    g28536(.A1(new_n30970_), .A2(pi0057), .A3(pi1151), .A4(new_n30972_), .ZN(new_n30973_));
  NAND2_X1   g28537(.A1(new_n29218_), .A2(new_n29014_), .ZN(new_n30974_));
  NAND2_X1   g28538(.A1(new_n30974_), .A2(pi0212), .ZN(new_n30975_));
  NOR3_X1    g28539(.A1(new_n29672_), .A2(pi0214), .A3(new_n30925_), .ZN(new_n30976_));
  OAI21_X1   g28540(.A1(new_n30975_), .A2(new_n30976_), .B(new_n8807_), .ZN(new_n30977_));
  NOR3_X1    g28541(.A1(new_n29672_), .A2(new_n8511_), .A3(new_n30925_), .ZN(new_n30978_));
  NOR3_X1    g28542(.A1(new_n30978_), .A2(pi0212), .A3(new_n29062_), .ZN(new_n30979_));
  NOR2_X1    g28543(.A1(new_n29055_), .A2(new_n6165_), .ZN(new_n30980_));
  OAI21_X1   g28544(.A1(new_n30977_), .A2(new_n30979_), .B(new_n30980_), .ZN(new_n30981_));
  NAND3_X1   g28545(.A1(new_n30981_), .A2(new_n2582_), .A3(new_n30971_), .ZN(new_n30982_));
  OAI22_X1   g28546(.A1(new_n30982_), .A2(new_n29035_), .B1(new_n2582_), .B2(new_n28367_), .ZN(new_n30983_));
  OAI21_X1   g28547(.A1(new_n30973_), .A2(new_n30983_), .B(new_n28422_), .ZN(new_n30984_));
  AOI21_X1   g28548(.A1(new_n30960_), .A2(new_n30984_), .B(new_n30948_), .ZN(new_n30985_));
  AOI21_X1   g28549(.A1(pi0213), .A2(new_n30985_), .B(new_n30924_), .ZN(new_n30986_));
  OAI21_X1   g28550(.A1(new_n30986_), .A2(pi0209), .B(pi0230), .ZN(new_n30987_));
  OAI22_X1   g28551(.A1(new_n30987_), .A2(new_n30923_), .B1(pi0230), .B2(new_n3865_), .ZN(po0406));
  OAI21_X1   g28552(.A1(new_n9276_), .A2(new_n2575_), .B(new_n5339_), .ZN(new_n30989_));
  NOR4_X1    g28553(.A1(new_n5337_), .A2(pi0038), .A3(new_n3465_), .A4(pi0100), .ZN(new_n30990_));
  AOI21_X1   g28554(.A1(new_n30989_), .A2(new_n3465_), .B(new_n30990_), .ZN(new_n30991_));
  NOR4_X1    g28555(.A1(new_n30991_), .A2(pi0087), .A3(pi0250), .A4(new_n7268_), .ZN(po0407));
  INV_X1     g28556(.I(pi0251), .ZN(new_n30993_));
  NOR2_X1    g28557(.A1(new_n8531_), .A2(pi0476), .ZN(new_n30994_));
  AOI21_X1   g28558(.A1(new_n8531_), .A2(pi0897), .B(new_n30994_), .ZN(new_n30995_));
  NOR2_X1    g28559(.A1(new_n30995_), .A2(pi0199), .ZN(new_n30996_));
  NOR2_X1    g28560(.A1(new_n8531_), .A2(pi1039), .ZN(new_n30997_));
  NOR2_X1    g28561(.A1(pi0200), .A2(pi1053), .ZN(new_n30998_));
  OAI21_X1   g28562(.A1(new_n30997_), .A2(new_n30998_), .B(new_n8525_), .ZN(new_n30999_));
  NAND2_X1   g28563(.A1(new_n30996_), .A2(new_n30999_), .ZN(new_n31000_));
  OAI21_X1   g28564(.A1(new_n30993_), .A2(new_n30996_), .B(new_n31000_), .ZN(po0408));
  NAND3_X1   g28565(.A1(pi0057), .A2(pi0252), .A3(pi1092), .ZN(new_n31002_));
  NAND2_X1   g28566(.A1(new_n7253_), .A2(new_n31002_), .ZN(new_n31003_));
  NOR2_X1    g28567(.A1(pi0979), .A2(pi0984), .ZN(new_n31004_));
  NAND4_X1   g28568(.A1(new_n31004_), .A2(pi0835), .A3(pi0950), .A4(pi1001), .ZN(new_n31005_));
  NOR4_X1    g28569(.A1(new_n16148_), .A2(new_n5431_), .A3(new_n8896_), .A4(new_n31005_), .ZN(new_n31006_));
  NAND3_X1   g28570(.A1(new_n27986_), .A2(new_n9149_), .A3(new_n31006_), .ZN(new_n31007_));
  NAND2_X1   g28571(.A1(new_n31007_), .A2(new_n2704_), .ZN(new_n31008_));
  NOR2_X1    g28572(.A1(new_n3040_), .A2(pi0057), .ZN(new_n31009_));
  AOI21_X1   g28573(.A1(new_n31008_), .A2(new_n31009_), .B(new_n31003_), .ZN(new_n31010_));
  NOR2_X1    g28574(.A1(new_n31005_), .A2(new_n5329_), .ZN(new_n31011_));
  AOI21_X1   g28575(.A1(new_n9149_), .A2(new_n31011_), .B(pi0252), .ZN(new_n31012_));
  NOR3_X1    g28576(.A1(new_n31012_), .A2(new_n3040_), .A3(pi1093), .ZN(new_n31013_));
  MUX2_X1    g28577(.I0(new_n5551_), .I1(new_n27903_), .S(new_n31013_), .Z(new_n31014_));
  NOR2_X1    g28578(.A1(new_n5449_), .A2(new_n9345_), .ZN(new_n31015_));
  AOI21_X1   g28579(.A1(new_n31014_), .A2(new_n5449_), .B(new_n31015_), .ZN(new_n31016_));
  NOR2_X1    g28580(.A1(new_n31016_), .A2(new_n6764_), .ZN(new_n31017_));
  NOR2_X1    g28581(.A1(new_n5427_), .A2(new_n9345_), .ZN(new_n31018_));
  AOI21_X1   g28582(.A1(new_n31014_), .A2(new_n5427_), .B(new_n31018_), .ZN(new_n31019_));
  NOR2_X1    g28583(.A1(new_n31019_), .A2(new_n5422_), .ZN(new_n31020_));
  OAI21_X1   g28584(.A1(new_n31017_), .A2(new_n31020_), .B(pi0299), .ZN(new_n31021_));
  NOR2_X1    g28585(.A1(new_n31016_), .A2(new_n5445_), .ZN(new_n31022_));
  NOR2_X1    g28586(.A1(new_n31019_), .A2(new_n5446_), .ZN(new_n31023_));
  OAI21_X1   g28587(.A1(new_n31022_), .A2(new_n31023_), .B(new_n2628_), .ZN(new_n31024_));
  NAND3_X1   g28588(.A1(new_n31021_), .A2(new_n31024_), .A3(new_n8897_), .ZN(new_n31025_));
  AOI21_X1   g28589(.A1(new_n8898_), .A2(new_n9345_), .B(new_n7253_), .ZN(new_n31026_));
  AOI21_X1   g28590(.A1(new_n31025_), .A2(new_n31026_), .B(new_n31010_), .ZN(po0409));
  NOR2_X1    g28591(.A1(new_n28722_), .A2(new_n3022_), .ZN(new_n31028_));
  NOR2_X1    g28592(.A1(pi0253), .A2(pi1091), .ZN(new_n31029_));
  NOR3_X1    g28593(.A1(new_n6643_), .A2(new_n31028_), .A3(new_n31029_), .ZN(new_n31030_));
  INV_X1     g28594(.I(new_n31030_), .ZN(new_n31031_));
  NOR2_X1    g28595(.A1(new_n3022_), .A2(pi0211), .ZN(new_n31032_));
  INV_X1     g28596(.I(new_n31032_), .ZN(new_n31033_));
  NOR2_X1    g28597(.A1(new_n31033_), .A2(pi0219), .ZN(new_n31034_));
  OAI21_X1   g28598(.A1(new_n31031_), .A2(new_n31034_), .B(pi1152), .ZN(new_n31035_));
  NOR2_X1    g28599(.A1(new_n29187_), .A2(new_n8761_), .ZN(new_n31036_));
  NOR2_X1    g28600(.A1(new_n3022_), .A2(pi1153), .ZN(new_n31037_));
  OAI22_X1   g28601(.A1(new_n31036_), .A2(new_n31037_), .B1(new_n29991_), .B2(pi1091), .ZN(new_n31038_));
  NAND2_X1   g28602(.A1(new_n28045_), .A2(new_n9183_), .ZN(new_n31039_));
  OAI22_X1   g28603(.A1(new_n31038_), .A2(new_n31039_), .B1(pi0253), .B2(pi1091), .ZN(new_n31040_));
  OAI21_X1   g28604(.A1(po1038), .A2(new_n31040_), .B(new_n31031_), .ZN(new_n31041_));
  AOI21_X1   g28605(.A1(new_n31041_), .A2(pi1151), .B(new_n31035_), .ZN(new_n31042_));
  NOR2_X1    g28606(.A1(new_n28128_), .A2(pi0299), .ZN(new_n31043_));
  NOR2_X1    g28607(.A1(new_n9219_), .A2(new_n3022_), .ZN(new_n31044_));
  AOI21_X1   g28608(.A1(new_n31043_), .A2(new_n31044_), .B(new_n29991_), .ZN(new_n31045_));
  NAND2_X1   g28609(.A1(new_n28124_), .A2(new_n29946_), .ZN(new_n31046_));
  AOI21_X1   g28610(.A1(new_n31046_), .A2(pi1153), .B(new_n28044_), .ZN(new_n31047_));
  OAI21_X1   g28611(.A1(new_n9217_), .A2(new_n3022_), .B(new_n12841_), .ZN(new_n31048_));
  NAND2_X1   g28612(.A1(new_n31047_), .A2(new_n31048_), .ZN(new_n31049_));
  NAND2_X1   g28613(.A1(new_n28978_), .A2(pi1091), .ZN(new_n31050_));
  NAND2_X1   g28614(.A1(new_n29941_), .A2(new_n28451_), .ZN(new_n31051_));
  NAND3_X1   g28615(.A1(new_n31050_), .A2(new_n8808_), .A3(new_n31051_), .ZN(new_n31052_));
  OAI21_X1   g28616(.A1(new_n28128_), .A2(pi0299), .B(pi1091), .ZN(new_n31053_));
  AOI21_X1   g28617(.A1(new_n31053_), .A2(pi0211), .B(pi0253), .ZN(new_n31054_));
  AOI22_X1   g28618(.A1(new_n31054_), .A2(new_n31052_), .B1(new_n31045_), .B2(new_n31049_), .ZN(new_n31055_));
  NOR2_X1    g28619(.A1(pi0211), .A2(pi0219), .ZN(new_n31056_));
  NOR2_X1    g28620(.A1(new_n29385_), .A2(new_n31056_), .ZN(new_n31057_));
  INV_X1     g28621(.I(new_n31057_), .ZN(new_n31058_));
  NOR2_X1    g28622(.A1(new_n28128_), .A2(new_n3022_), .ZN(new_n31059_));
  OAI21_X1   g28623(.A1(new_n31059_), .A2(new_n31029_), .B(new_n31058_), .ZN(new_n31060_));
  NAND2_X1   g28624(.A1(new_n31060_), .A2(new_n29007_), .ZN(new_n31061_));
  OAI21_X1   g28625(.A1(new_n31055_), .A2(new_n31061_), .B(new_n31042_), .ZN(new_n31062_));
  NOR2_X1    g28626(.A1(new_n31036_), .A2(new_n12841_), .ZN(new_n31063_));
  INV_X1     g28627(.I(new_n31063_), .ZN(new_n31064_));
  AOI21_X1   g28628(.A1(new_n31064_), .A2(new_n10290_), .B(new_n3022_), .ZN(new_n31065_));
  OAI21_X1   g28629(.A1(new_n31065_), .A2(pi0253), .B(new_n6643_), .ZN(new_n31066_));
  NAND2_X1   g28630(.A1(new_n29969_), .A2(new_n12841_), .ZN(new_n31067_));
  NAND2_X1   g28631(.A1(new_n29942_), .A2(pi1153), .ZN(new_n31068_));
  NAND2_X1   g28632(.A1(new_n31067_), .A2(new_n31068_), .ZN(new_n31069_));
  AOI22_X1   g28633(.A1(new_n28135_), .A2(new_n31056_), .B1(pi0211), .B2(new_n28167_), .ZN(new_n31070_));
  OAI22_X1   g28634(.A1(new_n31070_), .A2(new_n3022_), .B1(new_n28044_), .B2(new_n31069_), .ZN(new_n31071_));
  AOI21_X1   g28635(.A1(new_n31071_), .A2(pi0253), .B(new_n31066_), .ZN(new_n31072_));
  NAND2_X1   g28636(.A1(new_n12841_), .A2(pi0219), .ZN(new_n31073_));
  AOI21_X1   g28637(.A1(new_n31073_), .A2(new_n8510_), .B(new_n3022_), .ZN(new_n31074_));
  NOR3_X1    g28638(.A1(new_n6643_), .A2(new_n31029_), .A3(new_n31074_), .ZN(new_n31075_));
  NOR3_X1    g28639(.A1(new_n31072_), .A2(new_n29035_), .A3(new_n31075_), .ZN(new_n31076_));
  NOR2_X1    g28640(.A1(new_n29991_), .A2(pi1091), .ZN(new_n31077_));
  NOR4_X1    g28641(.A1(po1038), .A2(new_n10289_), .A3(new_n28151_), .A4(new_n29044_), .ZN(new_n31078_));
  AND3_X2    g28642(.A1(new_n31078_), .A2(pi1091), .A3(pi1153), .Z(new_n31079_));
  NOR2_X1    g28643(.A1(new_n31031_), .A2(new_n8807_), .ZN(new_n31080_));
  NOR4_X1    g28644(.A1(new_n31080_), .A2(pi1151), .A3(new_n31077_), .A4(new_n31079_), .ZN(new_n31081_));
  OAI21_X1   g28645(.A1(new_n31076_), .A2(new_n31081_), .B(new_n28422_), .ZN(new_n31082_));
  NAND3_X1   g28646(.A1(new_n31082_), .A2(new_n29934_), .A3(new_n31062_), .ZN(new_n31083_));
  NOR2_X1    g28647(.A1(new_n30011_), .A2(pi0219), .ZN(new_n31084_));
  INV_X1     g28648(.I(new_n31084_), .ZN(new_n31085_));
  NOR2_X1    g28649(.A1(new_n30037_), .A2(pi0211), .ZN(new_n31086_));
  INV_X1     g28650(.I(new_n30029_), .ZN(new_n31087_));
  NOR2_X1    g28651(.A1(new_n31087_), .A2(new_n8510_), .ZN(new_n31088_));
  NOR3_X1    g28652(.A1(new_n31086_), .A2(new_n31088_), .A3(new_n8807_), .ZN(new_n31089_));
  INV_X1     g28653(.I(new_n31089_), .ZN(new_n31090_));
  AOI21_X1   g28654(.A1(new_n31090_), .A2(new_n31085_), .B(pi0253), .ZN(new_n31091_));
  NOR2_X1    g28655(.A1(new_n30021_), .A2(pi0219), .ZN(new_n31092_));
  INV_X1     g28656(.I(new_n31092_), .ZN(new_n31093_));
  AOI21_X1   g28657(.A1(new_n31093_), .A2(new_n31087_), .B(new_n29991_), .ZN(new_n31094_));
  NOR4_X1    g28658(.A1(new_n31094_), .A2(new_n6643_), .A3(new_n31028_), .A4(new_n31091_), .ZN(new_n31095_));
  OAI21_X1   g28659(.A1(new_n30104_), .A2(pi1091), .B(new_n12841_), .ZN(new_n31096_));
  NOR2_X1    g28660(.A1(new_n30048_), .A2(new_n30088_), .ZN(new_n31097_));
  INV_X1     g28661(.I(new_n31097_), .ZN(new_n31098_));
  OAI21_X1   g28662(.A1(pi0219), .A2(new_n31098_), .B(new_n31096_), .ZN(new_n31099_));
  INV_X1     g28663(.I(new_n30078_), .ZN(new_n31100_));
  INV_X1     g28664(.I(new_n30081_), .ZN(new_n31101_));
  NOR2_X1    g28665(.A1(new_n30063_), .A2(new_n30088_), .ZN(new_n31102_));
  OAI21_X1   g28666(.A1(pi0211), .A2(new_n31101_), .B(new_n31102_), .ZN(new_n31103_));
  NOR3_X1    g28667(.A1(new_n31103_), .A2(new_n30072_), .A3(new_n31100_), .ZN(new_n31104_));
  NOR2_X1    g28668(.A1(new_n31104_), .A2(new_n30050_), .ZN(new_n31105_));
  INV_X1     g28669(.I(new_n31105_), .ZN(new_n31106_));
  OAI21_X1   g28670(.A1(new_n31106_), .A2(new_n31099_), .B(pi0253), .ZN(new_n31107_));
  NAND2_X1   g28671(.A1(new_n31107_), .A2(new_n6643_), .ZN(new_n31108_));
  NOR2_X1    g28672(.A1(new_n30153_), .A2(pi1153), .ZN(new_n31109_));
  NOR2_X1    g28673(.A1(new_n31109_), .A2(new_n30058_), .ZN(new_n31110_));
  NOR2_X1    g28674(.A1(new_n30150_), .A2(pi0219), .ZN(new_n31111_));
  AOI21_X1   g28675(.A1(new_n31110_), .A2(new_n31111_), .B(pi0253), .ZN(new_n31112_));
  INV_X1     g28676(.I(new_n30122_), .ZN(new_n31113_));
  NOR2_X1    g28677(.A1(new_n31113_), .A2(new_n30058_), .ZN(new_n31114_));
  NAND2_X1   g28678(.A1(new_n31114_), .A2(new_n8510_), .ZN(new_n31115_));
  NAND2_X1   g28679(.A1(new_n31115_), .A2(new_n30067_), .ZN(new_n31116_));
  AOI21_X1   g28680(.A1(new_n31116_), .A2(pi1153), .B(new_n30104_), .ZN(new_n31117_));
  NOR2_X1    g28681(.A1(new_n31117_), .A2(new_n8807_), .ZN(new_n31118_));
  NAND2_X1   g28682(.A1(new_n31118_), .A2(new_n30071_), .ZN(new_n31119_));
  AOI21_X1   g28683(.A1(new_n31119_), .A2(new_n31112_), .B(new_n31108_), .ZN(new_n31120_));
  NOR3_X1    g28684(.A1(new_n31120_), .A2(pi1151), .A3(new_n31095_), .ZN(new_n31121_));
  AOI21_X1   g28685(.A1(new_n8510_), .A2(new_n30012_), .B(new_n31093_), .ZN(new_n31122_));
  NOR2_X1    g28686(.A1(new_n31122_), .A2(pi0219), .ZN(new_n31123_));
  NAND2_X1   g28687(.A1(new_n31123_), .A2(po1038), .ZN(new_n31124_));
  NOR2_X1    g28688(.A1(new_n31124_), .A2(new_n30037_), .ZN(new_n31125_));
  NOR3_X1    g28689(.A1(new_n31125_), .A2(new_n29035_), .A3(new_n31095_), .ZN(new_n31126_));
  INV_X1     g28690(.I(new_n31126_), .ZN(new_n31127_));
  NOR2_X1    g28691(.A1(new_n31104_), .A2(new_n30054_), .ZN(new_n31128_));
  NOR2_X1    g28692(.A1(new_n31128_), .A2(new_n12841_), .ZN(new_n31129_));
  INV_X1     g28693(.I(new_n30109_), .ZN(new_n31130_));
  NOR2_X1    g28694(.A1(new_n31130_), .A2(pi1153), .ZN(new_n31131_));
  OAI21_X1   g28695(.A1(new_n31129_), .A2(new_n31131_), .B(pi0219), .ZN(new_n31132_));
  NOR2_X1    g28696(.A1(new_n31103_), .A2(new_n31093_), .ZN(new_n31133_));
  NAND2_X1   g28697(.A1(new_n30090_), .A2(pi1153), .ZN(new_n31134_));
  NAND2_X1   g28698(.A1(new_n31133_), .A2(new_n31134_), .ZN(new_n31135_));
  NAND3_X1   g28699(.A1(new_n31132_), .A2(pi0253), .A3(new_n31135_), .ZN(new_n31136_));
  AOI21_X1   g28700(.A1(new_n31115_), .A2(new_n30129_), .B(new_n31093_), .ZN(new_n31137_));
  INV_X1     g28701(.I(new_n30160_), .ZN(new_n31138_));
  NOR2_X1    g28702(.A1(new_n31138_), .A2(pi1153), .ZN(new_n31139_));
  NOR2_X1    g28703(.A1(new_n31139_), .A2(pi0219), .ZN(new_n31140_));
  OAI21_X1   g28704(.A1(new_n12841_), .A2(new_n30133_), .B(new_n31140_), .ZN(new_n31141_));
  AOI21_X1   g28705(.A1(new_n31137_), .A2(new_n31141_), .B(new_n31118_), .ZN(new_n31142_));
  OR3_X2     g28706(.A1(new_n31142_), .A2(pi0253), .A3(new_n30058_), .Z(new_n31143_));
  AOI21_X1   g28707(.A1(new_n31143_), .A2(new_n31136_), .B(po1038), .ZN(new_n31144_));
  OAI21_X1   g28708(.A1(new_n31144_), .A2(new_n31127_), .B(new_n28422_), .ZN(new_n31145_));
  NAND2_X1   g28709(.A1(new_n30073_), .A2(pi0219), .ZN(new_n31146_));
  AOI21_X1   g28710(.A1(new_n31105_), .A2(pi1153), .B(new_n31146_), .ZN(new_n31147_));
  INV_X1     g28711(.I(new_n31137_), .ZN(new_n31148_));
  NAND2_X1   g28712(.A1(new_n31098_), .A2(new_n12841_), .ZN(new_n31149_));
  AOI21_X1   g28713(.A1(new_n30138_), .A2(new_n31149_), .B(new_n31148_), .ZN(new_n31150_));
  NOR3_X1    g28714(.A1(new_n31150_), .A2(new_n29991_), .A3(new_n31147_), .ZN(new_n31151_));
  INV_X1     g28715(.I(new_n31118_), .ZN(new_n31152_));
  INV_X1     g28716(.I(new_n31103_), .ZN(new_n31153_));
  NAND4_X1   g28717(.A1(new_n31153_), .A2(new_n8807_), .A3(new_n30140_), .A4(new_n31149_), .ZN(new_n31154_));
  OAI21_X1   g28718(.A1(new_n31152_), .A2(new_n30063_), .B(new_n31154_), .ZN(new_n31155_));
  AOI21_X1   g28719(.A1(new_n31155_), .A2(new_n29991_), .B(new_n31151_), .ZN(new_n31156_));
  OAI21_X1   g28720(.A1(new_n31156_), .A2(po1038), .B(new_n29035_), .ZN(new_n31157_));
  AOI21_X1   g28721(.A1(new_n31117_), .A2(pi0219), .B(pi0253), .ZN(new_n31158_));
  OAI21_X1   g28722(.A1(new_n30129_), .A2(new_n30090_), .B(pi1153), .ZN(new_n31159_));
  NAND2_X1   g28723(.A1(new_n30150_), .A2(new_n12841_), .ZN(new_n31160_));
  NAND3_X1   g28724(.A1(new_n31159_), .A2(new_n8807_), .A3(new_n31160_), .ZN(new_n31161_));
  INV_X1     g28725(.I(new_n31104_), .ZN(new_n31162_));
  NOR2_X1    g28726(.A1(new_n30122_), .A2(pi1153), .ZN(new_n31163_));
  AOI21_X1   g28727(.A1(new_n31162_), .A2(pi1153), .B(new_n31163_), .ZN(new_n31164_));
  AOI21_X1   g28728(.A1(new_n31164_), .A2(pi0219), .B(new_n29991_), .ZN(new_n31165_));
  AOI22_X1   g28729(.A1(new_n31158_), .A2(new_n31141_), .B1(new_n31165_), .B2(new_n31161_), .ZN(new_n31166_));
  OAI21_X1   g28730(.A1(new_n31166_), .A2(po1038), .B(new_n31126_), .ZN(new_n31167_));
  INV_X1     g28731(.I(new_n31095_), .ZN(new_n31168_));
  NOR2_X1    g28732(.A1(new_n31085_), .A2(new_n31086_), .ZN(new_n31169_));
  NOR2_X1    g28733(.A1(new_n31169_), .A2(new_n31093_), .ZN(new_n31170_));
  INV_X1     g28734(.I(new_n31170_), .ZN(new_n31171_));
  NOR2_X1    g28735(.A1(new_n30037_), .A2(new_n8807_), .ZN(new_n31172_));
  NOR2_X1    g28736(.A1(new_n31172_), .A2(new_n6643_), .ZN(new_n31173_));
  NAND2_X1   g28737(.A1(new_n31171_), .A2(new_n31173_), .ZN(new_n31174_));
  OAI21_X1   g28738(.A1(new_n30037_), .A2(new_n31174_), .B(new_n31168_), .ZN(new_n31175_));
  AOI21_X1   g28739(.A1(new_n31157_), .A2(new_n31167_), .B(new_n31175_), .ZN(new_n31176_));
  OAI22_X1   g28740(.A1(new_n31145_), .A2(new_n31121_), .B1(new_n31176_), .B2(new_n28422_), .ZN(new_n31177_));
  AOI21_X1   g28741(.A1(new_n31177_), .A2(new_n29933_), .B(pi0230), .ZN(new_n31178_));
  NAND3_X1   g28742(.A1(new_n28045_), .A2(pi1151), .A3(new_n9183_), .ZN(new_n31179_));
  OAI21_X1   g28743(.A1(new_n31063_), .A2(new_n31179_), .B(new_n6643_), .ZN(new_n31180_));
  NOR3_X1    g28744(.A1(new_n28154_), .A2(new_n12841_), .A3(new_n28044_), .ZN(new_n31181_));
  NOR4_X1    g28745(.A1(new_n31181_), .A2(new_n28128_), .A3(pi1151), .A4(new_n9220_), .ZN(new_n31182_));
  AOI21_X1   g28746(.A1(new_n29035_), .A2(new_n31056_), .B(new_n28723_), .ZN(new_n31183_));
  NOR2_X1    g28747(.A1(new_n31183_), .A2(new_n28422_), .ZN(new_n31184_));
  OAI21_X1   g28748(.A1(new_n31180_), .A2(new_n31182_), .B(new_n31184_), .ZN(new_n31185_));
  OAI21_X1   g28749(.A1(new_n28170_), .A2(new_n28102_), .B(new_n8808_), .ZN(new_n31186_));
  AND2_X2    g28750(.A1(new_n31070_), .A2(new_n31186_), .Z(new_n31187_));
  OAI21_X1   g28751(.A1(new_n28723_), .A2(new_n9218_), .B(pi1151), .ZN(new_n31188_));
  AOI21_X1   g28752(.A1(new_n31187_), .A2(new_n6643_), .B(new_n31188_), .ZN(new_n31189_));
  NOR3_X1    g28753(.A1(new_n6643_), .A2(pi0211), .A3(new_n8807_), .ZN(new_n31190_));
  NOR2_X1    g28754(.A1(new_n31190_), .A2(new_n31078_), .ZN(new_n31191_));
  INV_X1     g28755(.I(new_n31191_), .ZN(new_n31192_));
  AOI21_X1   g28756(.A1(new_n31192_), .A2(pi1153), .B(pi1151), .ZN(new_n31193_));
  OAI21_X1   g28757(.A1(new_n31189_), .A2(new_n31193_), .B(new_n28422_), .ZN(new_n31194_));
  NAND2_X1   g28758(.A1(new_n31194_), .A2(new_n31185_), .ZN(new_n31195_));
  AOI22_X1   g28759(.A1(new_n31178_), .A2(new_n31083_), .B1(pi0230), .B2(new_n31195_), .ZN(po0410));
  NOR3_X1    g28760(.A1(new_n28364_), .A2(new_n3022_), .A3(new_n31058_), .ZN(new_n31197_));
  NOR2_X1    g28761(.A1(new_n29992_), .A2(pi1091), .ZN(new_n31198_));
  OAI21_X1   g28762(.A1(new_n31197_), .A2(new_n31198_), .B(po1038), .ZN(new_n31199_));
  NOR2_X1    g28763(.A1(new_n28321_), .A2(new_n3022_), .ZN(new_n31200_));
  AOI21_X1   g28764(.A1(new_n31047_), .A2(new_n31200_), .B(new_n12785_), .ZN(new_n31201_));
  AOI21_X1   g28765(.A1(new_n12841_), .A2(new_n29937_), .B(new_n28978_), .ZN(new_n31202_));
  OAI21_X1   g28766(.A1(new_n31202_), .A2(new_n28126_), .B(pi1091), .ZN(new_n31203_));
  OAI21_X1   g28767(.A1(new_n31203_), .A2(new_n31057_), .B(new_n31201_), .ZN(new_n31204_));
  NOR2_X1    g28768(.A1(new_n9218_), .A2(new_n3022_), .ZN(new_n31205_));
  NAND2_X1   g28769(.A1(new_n28533_), .A2(new_n31205_), .ZN(new_n31206_));
  NAND2_X1   g28770(.A1(new_n31206_), .A2(new_n12785_), .ZN(new_n31207_));
  NOR2_X1    g28771(.A1(new_n3022_), .A2(pi1154), .ZN(new_n31208_));
  AOI22_X1   g28772(.A1(new_n31202_), .A2(pi1091), .B1(new_n28113_), .B2(new_n31208_), .ZN(new_n31209_));
  OAI21_X1   g28773(.A1(new_n31209_), .A2(new_n9219_), .B(pi0254), .ZN(new_n31210_));
  AOI21_X1   g28774(.A1(new_n31204_), .A2(new_n31207_), .B(new_n31210_), .ZN(new_n31211_));
  AOI21_X1   g28775(.A1(new_n28452_), .A2(pi1091), .B(new_n12785_), .ZN(new_n31212_));
  NAND2_X1   g28776(.A1(new_n31212_), .A2(pi0211), .ZN(new_n31213_));
  AOI21_X1   g28777(.A1(new_n28374_), .A2(pi1091), .B(pi1154), .ZN(new_n31214_));
  INV_X1     g28778(.I(new_n31214_), .ZN(new_n31215_));
  AOI21_X1   g28779(.A1(new_n28321_), .A2(new_n31037_), .B(new_n28004_), .ZN(new_n31216_));
  NAND2_X1   g28780(.A1(new_n31050_), .A2(new_n31216_), .ZN(new_n31217_));
  NAND4_X1   g28781(.A1(new_n31213_), .A2(new_n31217_), .A3(pi0219), .A4(new_n31215_), .ZN(new_n31218_));
  NOR3_X1    g28782(.A1(new_n31212_), .A2(pi0211), .A3(new_n31214_), .ZN(new_n31219_));
  NOR2_X1    g28783(.A1(new_n29948_), .A2(new_n12841_), .ZN(new_n31220_));
  NOR2_X1    g28784(.A1(new_n31220_), .A2(pi1154), .ZN(new_n31221_));
  NOR4_X1    g28785(.A1(new_n31202_), .A2(new_n8510_), .A3(new_n3022_), .A4(new_n31221_), .ZN(new_n31222_));
  OAI21_X1   g28786(.A1(new_n31222_), .A2(new_n31219_), .B(new_n8807_), .ZN(new_n31223_));
  AOI21_X1   g28787(.A1(new_n31223_), .A2(new_n31218_), .B(pi0254), .ZN(new_n31224_));
  OAI21_X1   g28788(.A1(new_n31211_), .A2(new_n31224_), .B(new_n6643_), .ZN(new_n31225_));
  NAND3_X1   g28789(.A1(new_n31225_), .A2(new_n28422_), .A3(new_n31199_), .ZN(new_n31226_));
  INV_X1     g28790(.I(new_n31199_), .ZN(new_n31227_));
  AOI21_X1   g28791(.A1(new_n29156_), .A2(new_n31032_), .B(new_n31227_), .ZN(new_n31228_));
  OAI21_X1   g28792(.A1(new_n28176_), .A2(new_n28405_), .B(new_n28011_), .ZN(new_n31229_));
  NAND2_X1   g28793(.A1(new_n28377_), .A2(new_n12785_), .ZN(new_n31230_));
  AND3_X2    g28794(.A1(new_n31230_), .A2(new_n31229_), .A3(new_n28433_), .Z(new_n31231_));
  NOR2_X1    g28795(.A1(new_n28003_), .A2(pi0219), .ZN(new_n31232_));
  NOR3_X1    g28796(.A1(new_n31231_), .A2(new_n3022_), .A3(new_n31232_), .ZN(new_n31233_));
  NAND4_X1   g28797(.A1(new_n28391_), .A2(pi1091), .A3(new_n28136_), .A4(new_n28011_), .ZN(new_n31234_));
  NAND2_X1   g28798(.A1(new_n28388_), .A2(new_n8510_), .ZN(new_n31235_));
  NAND3_X1   g28799(.A1(new_n31067_), .A2(new_n31221_), .A3(new_n31235_), .ZN(new_n31236_));
  AOI21_X1   g28800(.A1(new_n31236_), .A2(new_n31234_), .B(pi0219), .ZN(new_n31237_));
  NOR3_X1    g28801(.A1(new_n31233_), .A2(new_n31237_), .A3(new_n29992_), .ZN(new_n31238_));
  AOI21_X1   g28802(.A1(new_n8531_), .A2(pi1154), .B(new_n9172_), .ZN(new_n31239_));
  INV_X1     g28803(.I(new_n31239_), .ZN(new_n31240_));
  NAND2_X1   g28804(.A1(new_n29188_), .A2(new_n28405_), .ZN(new_n31241_));
  AOI21_X1   g28805(.A1(new_n31240_), .A2(new_n31241_), .B(pi0219), .ZN(new_n31242_));
  NOR2_X1    g28806(.A1(new_n31036_), .A2(new_n12785_), .ZN(new_n31243_));
  NOR3_X1    g28807(.A1(new_n31243_), .A2(new_n8807_), .A3(new_n28376_), .ZN(new_n31244_));
  NOR4_X1    g28808(.A1(new_n31242_), .A2(pi0254), .A3(new_n3022_), .A4(new_n31244_), .ZN(new_n31245_));
  OAI21_X1   g28809(.A1(new_n31238_), .A2(new_n31245_), .B(new_n6643_), .ZN(new_n31246_));
  NAND3_X1   g28810(.A1(new_n31246_), .A2(pi1152), .A3(new_n31228_), .ZN(new_n31247_));
  NAND3_X1   g28811(.A1(new_n31226_), .A2(new_n29934_), .A3(new_n31247_), .ZN(new_n31248_));
  NOR2_X1    g28812(.A1(new_n6643_), .A2(new_n29991_), .ZN(new_n31249_));
  NAND2_X1   g28813(.A1(new_n28352_), .A2(pi1091), .ZN(new_n31250_));
  OAI21_X1   g28814(.A1(new_n3022_), .A2(new_n12841_), .B(new_n31169_), .ZN(new_n31251_));
  NAND4_X1   g28815(.A1(new_n31251_), .A2(new_n29992_), .A3(new_n31090_), .A4(new_n31250_), .ZN(new_n31252_));
  OAI21_X1   g28816(.A1(new_n31252_), .A2(new_n31123_), .B(pi0253), .ZN(new_n31253_));
  AOI21_X1   g28817(.A1(new_n31044_), .A2(new_n12841_), .B(new_n29992_), .ZN(new_n31254_));
  NOR2_X1    g28818(.A1(new_n30012_), .A2(pi0219), .ZN(new_n31255_));
  INV_X1     g28819(.I(new_n31255_), .ZN(new_n31256_));
  OAI21_X1   g28820(.A1(pi0211), .A2(new_n30025_), .B(new_n31172_), .ZN(new_n31257_));
  NAND4_X1   g28821(.A1(new_n31256_), .A2(new_n31250_), .A3(new_n31254_), .A4(new_n31257_), .ZN(new_n31258_));
  NOR2_X1    g28822(.A1(new_n31170_), .A2(new_n31258_), .ZN(new_n31259_));
  OAI22_X1   g28823(.A1(new_n31253_), .A2(new_n31259_), .B1(new_n31227_), .B2(new_n31249_), .ZN(new_n31260_));
  OAI21_X1   g28824(.A1(new_n31211_), .A2(new_n31224_), .B(new_n29991_), .ZN(new_n31261_));
  NOR2_X1    g28825(.A1(new_n30113_), .A2(pi1153), .ZN(new_n31262_));
  NOR2_X1    g28826(.A1(new_n30105_), .A2(new_n30053_), .ZN(new_n31263_));
  INV_X1     g28827(.I(new_n31263_), .ZN(new_n31264_));
  OAI21_X1   g28828(.A1(new_n31264_), .A2(new_n31262_), .B(new_n12785_), .ZN(new_n31265_));
  NOR2_X1    g28829(.A1(new_n30065_), .A2(new_n31130_), .ZN(new_n31266_));
  INV_X1     g28830(.I(new_n31266_), .ZN(new_n31267_));
  OAI21_X1   g28831(.A1(new_n31267_), .A2(new_n31163_), .B(new_n28003_), .ZN(new_n31268_));
  OAI21_X1   g28832(.A1(new_n30069_), .A2(new_n31163_), .B(new_n28011_), .ZN(new_n31269_));
  NAND4_X1   g28833(.A1(new_n31269_), .A2(pi0219), .A3(new_n31265_), .A4(new_n31268_), .ZN(new_n31270_));
  NAND2_X1   g28834(.A1(new_n30063_), .A2(pi1154), .ZN(new_n31271_));
  NAND2_X1   g28835(.A1(new_n31271_), .A2(new_n31101_), .ZN(new_n31272_));
  AOI21_X1   g28836(.A1(new_n31272_), .A2(new_n8510_), .B(pi0219), .ZN(new_n31273_));
  INV_X1     g28837(.I(new_n30151_), .ZN(new_n31274_));
  NOR2_X1    g28838(.A1(new_n31138_), .A2(new_n30053_), .ZN(new_n31275_));
  INV_X1     g28839(.I(new_n31275_), .ZN(new_n31276_));
  OAI22_X1   g28840(.A1(new_n12785_), .A2(new_n31274_), .B1(new_n31276_), .B2(new_n31109_), .ZN(new_n31277_));
  AOI21_X1   g28841(.A1(new_n31277_), .A2(new_n31273_), .B(pi0254), .ZN(new_n31278_));
  NAND2_X1   g28842(.A1(new_n31270_), .A2(new_n31278_), .ZN(new_n31279_));
  NAND2_X1   g28843(.A1(new_n30048_), .A2(pi1154), .ZN(new_n31280_));
  INV_X1     g28844(.I(new_n31280_), .ZN(new_n31281_));
  INV_X1     g28845(.I(new_n31115_), .ZN(new_n31282_));
  NOR2_X1    g28846(.A1(new_n31100_), .A2(pi1153), .ZN(new_n31283_));
  NOR3_X1    g28847(.A1(new_n31282_), .A2(new_n30082_), .A3(new_n31283_), .ZN(new_n31284_));
  NOR3_X1    g28848(.A1(new_n31284_), .A2(pi0219), .A3(new_n31281_), .ZN(new_n31285_));
  OAI21_X1   g28849(.A1(new_n30050_), .A2(new_n28004_), .B(pi0219), .ZN(new_n31286_));
  INV_X1     g28850(.I(new_n30072_), .ZN(new_n31287_));
  OAI21_X1   g28851(.A1(new_n31287_), .A2(new_n12841_), .B(new_n30078_), .ZN(new_n31288_));
  NOR2_X1    g28852(.A1(new_n30099_), .A2(new_n30042_), .ZN(new_n31289_));
  NAND2_X1   g28853(.A1(new_n31289_), .A2(new_n12785_), .ZN(new_n31290_));
  AOI21_X1   g28854(.A1(new_n31288_), .A2(new_n31290_), .B(new_n31286_), .ZN(new_n31291_));
  OAI21_X1   g28855(.A1(new_n31285_), .A2(new_n31291_), .B(pi0254), .ZN(new_n31292_));
  NAND3_X1   g28856(.A1(new_n31279_), .A2(pi0253), .A3(new_n31292_), .ZN(new_n31293_));
  NAND2_X1   g28857(.A1(new_n31293_), .A2(new_n31261_), .ZN(new_n31294_));
  AOI21_X1   g28858(.A1(new_n31294_), .A2(new_n6643_), .B(pi1152), .ZN(new_n31295_));
  AOI21_X1   g28859(.A1(new_n31295_), .A2(new_n31260_), .B(new_n29934_), .ZN(new_n31296_));
  INV_X1     g28860(.I(new_n28011_), .ZN(new_n31297_));
  NOR2_X1    g28861(.A1(new_n30067_), .A2(new_n12841_), .ZN(new_n31298_));
  NOR3_X1    g28862(.A1(new_n31298_), .A2(new_n31297_), .A3(new_n30096_), .ZN(new_n31299_));
  NOR2_X1    g28863(.A1(new_n31265_), .A2(new_n30106_), .ZN(new_n31300_));
  NOR2_X1    g28864(.A1(new_n31268_), .A2(new_n30057_), .ZN(new_n31301_));
  NOR4_X1    g28865(.A1(new_n31301_), .A2(new_n31299_), .A3(new_n31300_), .A4(pi0254), .ZN(new_n31302_));
  OAI21_X1   g28866(.A1(pi1153), .A2(new_n30055_), .B(new_n31162_), .ZN(new_n31303_));
  AOI21_X1   g28867(.A1(pi1153), .A2(new_n30122_), .B(new_n31131_), .ZN(new_n31304_));
  OAI21_X1   g28868(.A1(new_n31304_), .A2(pi1154), .B(pi0254), .ZN(new_n31305_));
  AOI21_X1   g28869(.A1(new_n31303_), .A2(pi1154), .B(new_n31305_), .ZN(new_n31306_));
  NOR3_X1    g28870(.A1(new_n31302_), .A2(new_n8807_), .A3(new_n31306_), .ZN(new_n31307_));
  OAI21_X1   g28871(.A1(new_n31267_), .A2(new_n12785_), .B(new_n31138_), .ZN(new_n31308_));
  NOR2_X1    g28872(.A1(new_n31101_), .A2(new_n8510_), .ZN(new_n31309_));
  OAI21_X1   g28873(.A1(new_n30058_), .A2(new_n31309_), .B(new_n12841_), .ZN(new_n31310_));
  NAND3_X1   g28874(.A1(new_n31308_), .A2(new_n29992_), .A3(new_n31310_), .ZN(new_n31311_));
  NAND4_X1   g28875(.A1(new_n31159_), .A2(pi1154), .A3(new_n30047_), .A4(new_n31153_), .ZN(new_n31312_));
  NOR4_X1    g28876(.A1(new_n31103_), .A2(new_n30065_), .A3(new_n31098_), .A4(pi1153), .ZN(new_n31313_));
  OAI21_X1   g28877(.A1(new_n31313_), .A2(new_n30149_), .B(new_n12785_), .ZN(new_n31314_));
  NAND3_X1   g28878(.A1(new_n31312_), .A2(new_n31314_), .A3(pi0254), .ZN(new_n31315_));
  AND3_X2    g28879(.A1(new_n31315_), .A2(new_n8807_), .A3(new_n31311_), .Z(new_n31316_));
  OAI21_X1   g28880(.A1(new_n31316_), .A2(new_n31307_), .B(pi0253), .ZN(new_n31317_));
  OR3_X2     g28881(.A1(new_n31238_), .A2(pi0253), .A3(new_n31245_), .Z(new_n31318_));
  NAND3_X1   g28882(.A1(new_n31317_), .A2(new_n6643_), .A3(new_n31318_), .ZN(new_n31319_));
  OAI21_X1   g28883(.A1(new_n29991_), .A2(new_n6643_), .B(new_n31228_), .ZN(new_n31320_));
  NAND3_X1   g28884(.A1(new_n31252_), .A2(pi0253), .A3(new_n31258_), .ZN(new_n31321_));
  AOI21_X1   g28885(.A1(new_n31321_), .A2(new_n31320_), .B(new_n28422_), .ZN(new_n31322_));
  NAND2_X1   g28886(.A1(new_n31319_), .A2(new_n31322_), .ZN(new_n31323_));
  AOI21_X1   g28887(.A1(new_n31296_), .A2(new_n31323_), .B(pi0230), .ZN(new_n31324_));
  AOI21_X1   g28888(.A1(new_n28468_), .A2(pi1154), .B(new_n28407_), .ZN(new_n31325_));
  NOR2_X1    g28889(.A1(new_n28044_), .A2(new_n2628_), .ZN(new_n31326_));
  AOI21_X1   g28890(.A1(new_n28452_), .A2(new_n9219_), .B(new_n31326_), .ZN(new_n31327_));
  OAI22_X1   g28891(.A1(new_n31327_), .A2(new_n28375_), .B1(new_n31325_), .B2(new_n9219_), .ZN(new_n31328_));
  NOR2_X1    g28892(.A1(new_n31328_), .A2(po1038), .ZN(new_n31329_));
  AOI21_X1   g28893(.A1(new_n28363_), .A2(new_n31057_), .B(new_n6643_), .ZN(new_n31330_));
  NOR2_X1    g28894(.A1(new_n31329_), .A2(new_n31330_), .ZN(new_n31331_));
  AOI21_X1   g28895(.A1(new_n8807_), .A2(new_n28362_), .B(new_n29232_), .ZN(new_n31332_));
  OAI21_X1   g28896(.A1(new_n31231_), .A2(new_n8807_), .B(new_n6643_), .ZN(new_n31333_));
  OAI21_X1   g28897(.A1(new_n31333_), .A2(new_n31242_), .B(pi1152), .ZN(new_n31334_));
  OAI22_X1   g28898(.A1(new_n31334_), .A2(new_n31332_), .B1(new_n31331_), .B2(pi1152), .ZN(new_n31335_));
  AOI22_X1   g28899(.A1(new_n31324_), .A2(new_n31248_), .B1(pi0230), .B2(new_n31335_), .ZN(po0411));
  INV_X1     g28900(.I(pi0255), .ZN(new_n31337_));
  INV_X1     g28901(.I(pi1036), .ZN(new_n31338_));
  NOR2_X1    g28902(.A1(pi0200), .A2(pi1049), .ZN(new_n31339_));
  AOI21_X1   g28903(.A1(pi0200), .A2(new_n31338_), .B(new_n31339_), .ZN(new_n31340_));
  NAND2_X1   g28904(.A1(new_n30996_), .A2(new_n31340_), .ZN(new_n31341_));
  OAI21_X1   g28905(.A1(new_n31337_), .A2(new_n30996_), .B(new_n31341_), .ZN(po0412));
  INV_X1     g28906(.I(pi0256), .ZN(new_n31343_));
  INV_X1     g28907(.I(pi1070), .ZN(new_n31344_));
  NOR2_X1    g28908(.A1(pi0200), .A2(pi1048), .ZN(new_n31345_));
  AOI21_X1   g28909(.A1(pi0200), .A2(new_n31344_), .B(new_n31345_), .ZN(new_n31346_));
  NAND2_X1   g28910(.A1(new_n30996_), .A2(new_n31346_), .ZN(new_n31347_));
  OAI21_X1   g28911(.A1(new_n31343_), .A2(new_n30996_), .B(new_n31347_), .ZN(po0413));
  INV_X1     g28912(.I(pi0257), .ZN(new_n31349_));
  INV_X1     g28913(.I(pi1065), .ZN(new_n31350_));
  NOR2_X1    g28914(.A1(pi0200), .A2(pi1084), .ZN(new_n31351_));
  AOI21_X1   g28915(.A1(pi0200), .A2(new_n31350_), .B(new_n31351_), .ZN(new_n31352_));
  NAND2_X1   g28916(.A1(new_n30996_), .A2(new_n31352_), .ZN(new_n31353_));
  OAI21_X1   g28917(.A1(new_n31349_), .A2(new_n30996_), .B(new_n31353_), .ZN(po0414));
  INV_X1     g28918(.I(pi0258), .ZN(new_n31355_));
  INV_X1     g28919(.I(pi1062), .ZN(new_n31356_));
  NOR2_X1    g28920(.A1(pi0200), .A2(pi1072), .ZN(new_n31357_));
  AOI21_X1   g28921(.A1(pi0200), .A2(new_n31356_), .B(new_n31357_), .ZN(new_n31358_));
  NAND2_X1   g28922(.A1(new_n30996_), .A2(new_n31358_), .ZN(new_n31359_));
  OAI21_X1   g28923(.A1(new_n31355_), .A2(new_n30996_), .B(new_n31359_), .ZN(po0415));
  INV_X1     g28924(.I(pi0259), .ZN(new_n31361_));
  INV_X1     g28925(.I(pi1069), .ZN(new_n31362_));
  NOR2_X1    g28926(.A1(pi0200), .A2(pi1059), .ZN(new_n31363_));
  AOI21_X1   g28927(.A1(pi0200), .A2(new_n31362_), .B(new_n31363_), .ZN(new_n31364_));
  NAND2_X1   g28928(.A1(new_n30996_), .A2(new_n31364_), .ZN(new_n31365_));
  OAI21_X1   g28929(.A1(new_n31361_), .A2(new_n30996_), .B(new_n31365_), .ZN(po0416));
  INV_X1     g28930(.I(pi0260), .ZN(new_n31367_));
  NOR2_X1    g28931(.A1(new_n8531_), .A2(pi1067), .ZN(new_n31368_));
  NOR2_X1    g28932(.A1(pi0200), .A2(pi1044), .ZN(new_n31369_));
  OAI21_X1   g28933(.A1(new_n31368_), .A2(new_n31369_), .B(new_n8525_), .ZN(new_n31370_));
  NAND2_X1   g28934(.A1(new_n30996_), .A2(new_n31370_), .ZN(new_n31371_));
  OAI21_X1   g28935(.A1(new_n31367_), .A2(new_n30996_), .B(new_n31371_), .ZN(po0417));
  INV_X1     g28936(.I(pi0261), .ZN(new_n31373_));
  NOR2_X1    g28937(.A1(new_n8531_), .A2(pi1040), .ZN(new_n31374_));
  NOR2_X1    g28938(.A1(pi0200), .A2(pi1037), .ZN(new_n31375_));
  OAI21_X1   g28939(.A1(new_n31374_), .A2(new_n31375_), .B(new_n8525_), .ZN(new_n31376_));
  NAND2_X1   g28940(.A1(new_n30996_), .A2(new_n31376_), .ZN(new_n31377_));
  OAI21_X1   g28941(.A1(new_n31373_), .A2(new_n30996_), .B(new_n31377_), .ZN(po0418));
  NAND2_X1   g28942(.A1(new_n3774_), .A2(new_n3041_), .ZN(new_n31379_));
  NAND2_X1   g28943(.A1(pi1093), .A2(pi1142), .ZN(new_n31380_));
  AOI21_X1   g28944(.A1(new_n31379_), .A2(new_n31380_), .B(pi0228), .ZN(new_n31381_));
  NAND2_X1   g28945(.A1(new_n3774_), .A2(pi0123), .ZN(new_n31382_));
  INV_X1     g28946(.I(pi0123), .ZN(new_n31383_));
  NAND2_X1   g28947(.A1(new_n31383_), .A2(pi1142), .ZN(new_n31384_));
  AOI21_X1   g28948(.A1(new_n31382_), .A2(new_n31384_), .B(new_n2458_), .ZN(new_n31385_));
  NOR2_X1    g28949(.A1(new_n31381_), .A2(new_n31385_), .ZN(new_n31386_));
  NOR2_X1    g28950(.A1(new_n2458_), .A2(pi0123), .ZN(new_n31387_));
  AOI21_X1   g28951(.A1(new_n2458_), .A2(pi1093), .B(new_n31387_), .ZN(new_n31388_));
  OAI21_X1   g28952(.A1(new_n28385_), .A2(new_n31388_), .B(po1038), .ZN(new_n31389_));
  OAI21_X1   g28953(.A1(new_n31388_), .A2(new_n29022_), .B(new_n2628_), .ZN(new_n31390_));
  NOR2_X1    g28954(.A1(new_n31390_), .A2(new_n31386_), .ZN(new_n31391_));
  INV_X1     g28955(.I(new_n31388_), .ZN(new_n31392_));
  NOR2_X1    g28956(.A1(new_n31392_), .A2(pi0262), .ZN(new_n31393_));
  NOR2_X1    g28957(.A1(new_n29730_), .A2(new_n31393_), .ZN(new_n31394_));
  OAI21_X1   g28958(.A1(new_n31394_), .A2(new_n2628_), .B(pi0208), .ZN(new_n31395_));
  NOR2_X1    g28959(.A1(new_n31395_), .A2(new_n31391_), .ZN(new_n31396_));
  AOI21_X1   g28960(.A1(new_n31393_), .A2(new_n8521_), .B(pi0208), .ZN(new_n31397_));
  NOR2_X1    g28961(.A1(new_n29730_), .A2(new_n31397_), .ZN(new_n31398_));
  OAI21_X1   g28962(.A1(new_n31388_), .A2(new_n8525_), .B(new_n28026_), .ZN(new_n31399_));
  AOI21_X1   g28963(.A1(new_n31394_), .A2(new_n31399_), .B(new_n31386_), .ZN(new_n31400_));
  OAI21_X1   g28964(.A1(new_n31400_), .A2(new_n31398_), .B(new_n6643_), .ZN(new_n31401_));
  OAI22_X1   g28965(.A1(new_n31401_), .A2(new_n31396_), .B1(new_n31386_), .B2(new_n31389_), .ZN(po0419));
  AOI21_X1   g28966(.A1(new_n28659_), .A2(new_n28182_), .B(pi1156), .ZN(new_n31403_));
  OR2_X2     g28967(.A1(new_n28216_), .A2(new_n28507_), .Z(new_n31404_));
  AOI21_X1   g28968(.A1(new_n29187_), .A2(pi1156), .B(new_n8807_), .ZN(new_n31405_));
  OAI21_X1   g28969(.A1(new_n31403_), .A2(new_n31404_), .B(new_n31405_), .ZN(new_n31406_));
  INV_X1     g28970(.I(new_n28477_), .ZN(new_n31407_));
  OAI21_X1   g28971(.A1(new_n28891_), .A2(new_n28181_), .B(new_n31407_), .ZN(new_n31408_));
  AOI21_X1   g28972(.A1(new_n31408_), .A2(new_n8510_), .B(pi0219), .ZN(new_n31409_));
  OAI21_X1   g28973(.A1(new_n31403_), .A2(new_n31404_), .B(new_n28282_), .ZN(new_n31410_));
  NAND2_X1   g28974(.A1(new_n31410_), .A2(pi0211), .ZN(new_n31411_));
  NAND2_X1   g28975(.A1(new_n31409_), .A2(new_n31411_), .ZN(new_n31412_));
  NAND3_X1   g28976(.A1(new_n31412_), .A2(new_n6643_), .A3(new_n31406_), .ZN(new_n31413_));
  AOI22_X1   g28977(.A1(new_n31232_), .A2(new_n28354_), .B1(new_n28353_), .B2(pi0219), .ZN(new_n31414_));
  AOI21_X1   g28978(.A1(new_n31414_), .A2(po1038), .B(new_n27999_), .ZN(new_n31415_));
  INV_X1     g28979(.I(pi0263), .ZN(new_n31416_));
  NOR2_X1    g28980(.A1(new_n8510_), .A2(new_n3022_), .ZN(new_n31417_));
  OAI21_X1   g28981(.A1(pi0199), .A2(pi1154), .B(new_n8761_), .ZN(new_n31418_));
  NAND3_X1   g28982(.A1(new_n28326_), .A2(new_n31417_), .A3(new_n31418_), .ZN(new_n31419_));
  NOR2_X1    g28983(.A1(new_n28125_), .A2(new_n3022_), .ZN(new_n31420_));
  NOR2_X1    g28984(.A1(new_n28465_), .A2(new_n12770_), .ZN(new_n31421_));
  INV_X1     g28985(.I(new_n31421_), .ZN(new_n31422_));
  AOI22_X1   g28986(.A1(new_n31422_), .A2(new_n29941_), .B1(new_n12785_), .B2(new_n31420_), .ZN(new_n31423_));
  OR2_X2     g28987(.A1(new_n31423_), .A2(pi0211), .Z(new_n31424_));
  NAND3_X1   g28988(.A1(new_n31424_), .A2(pi1156), .A3(new_n31419_), .ZN(new_n31425_));
  NOR2_X1    g28989(.A1(new_n29963_), .A2(new_n31208_), .ZN(new_n31426_));
  NOR2_X1    g28990(.A1(new_n31426_), .A2(new_n28325_), .ZN(new_n31427_));
  NAND2_X1   g28991(.A1(new_n31427_), .A2(pi0211), .ZN(new_n31428_));
  NAND3_X1   g28992(.A1(new_n28623_), .A2(new_n31407_), .A3(new_n31032_), .ZN(new_n31429_));
  NAND3_X1   g28993(.A1(new_n31428_), .A2(new_n12742_), .A3(new_n31429_), .ZN(new_n31430_));
  AOI21_X1   g28994(.A1(new_n31425_), .A2(new_n31430_), .B(pi0219), .ZN(new_n31431_));
  INV_X1     g28995(.I(new_n28017_), .ZN(new_n31432_));
  AOI21_X1   g28996(.A1(new_n31423_), .A2(new_n29979_), .B(new_n31432_), .ZN(new_n31433_));
  NOR3_X1    g28997(.A1(new_n31426_), .A2(pi1156), .A3(new_n28147_), .ZN(new_n31434_));
  AOI21_X1   g28998(.A1(new_n28146_), .A2(new_n28102_), .B(new_n12785_), .ZN(new_n31435_));
  NOR2_X1    g28999(.A1(new_n28156_), .A2(pi1154), .ZN(new_n31436_));
  NOR4_X1    g29000(.A1(new_n31436_), .A2(new_n3022_), .A3(new_n28353_), .A4(new_n31435_), .ZN(new_n31437_));
  NOR4_X1    g29001(.A1(new_n31437_), .A2(new_n8807_), .A3(new_n31433_), .A4(new_n31434_), .ZN(new_n31438_));
  OAI21_X1   g29002(.A1(new_n31431_), .A2(new_n31438_), .B(new_n31416_), .ZN(new_n31439_));
  NAND2_X1   g29003(.A1(new_n28215_), .A2(pi1154), .ZN(new_n31440_));
  AOI21_X1   g29004(.A1(new_n31440_), .A2(pi1156), .B(pi0299), .ZN(new_n31441_));
  OAI21_X1   g29005(.A1(new_n28188_), .A2(pi1154), .B(new_n29188_), .ZN(new_n31442_));
  OAI21_X1   g29006(.A1(new_n31442_), .A2(new_n31441_), .B(pi1156), .ZN(new_n31443_));
  NAND2_X1   g29007(.A1(new_n28623_), .A2(new_n31407_), .ZN(new_n31444_));
  AOI21_X1   g29008(.A1(new_n31441_), .A2(new_n31444_), .B(new_n8807_), .ZN(new_n31445_));
  NAND2_X1   g29009(.A1(new_n31443_), .A2(new_n31445_), .ZN(new_n31446_));
  INV_X1     g29010(.I(new_n28104_), .ZN(new_n31447_));
  OAI21_X1   g29011(.A1(new_n28129_), .A2(new_n8761_), .B(pi1154), .ZN(new_n31448_));
  NAND2_X1   g29012(.A1(new_n31448_), .A2(pi1156), .ZN(new_n31449_));
  AOI21_X1   g29013(.A1(new_n31436_), .A2(new_n31447_), .B(new_n31449_), .ZN(new_n31450_));
  NAND2_X1   g29014(.A1(new_n31427_), .A2(new_n12742_), .ZN(new_n31451_));
  NAND2_X1   g29015(.A1(new_n31451_), .A2(pi0211), .ZN(new_n31452_));
  OAI21_X1   g29016(.A1(new_n31450_), .A2(new_n31452_), .B(new_n31409_), .ZN(new_n31453_));
  NAND4_X1   g29017(.A1(new_n31453_), .A2(pi0263), .A3(pi1091), .A4(new_n31446_), .ZN(new_n31454_));
  AOI21_X1   g29018(.A1(new_n31439_), .A2(new_n31454_), .B(po1038), .ZN(new_n31455_));
  NOR2_X1    g29019(.A1(pi0263), .A2(pi1091), .ZN(new_n31456_));
  AOI21_X1   g29020(.A1(new_n31414_), .A2(pi1091), .B(new_n31456_), .ZN(new_n31457_));
  NOR2_X1    g29021(.A1(new_n31457_), .A2(new_n6643_), .ZN(new_n31458_));
  OAI21_X1   g29022(.A1(new_n31455_), .A2(new_n31458_), .B(new_n29934_), .ZN(new_n31459_));
  NAND2_X1   g29023(.A1(new_n31439_), .A2(new_n31454_), .ZN(new_n31460_));
  NOR2_X1    g29024(.A1(new_n31287_), .A2(new_n12770_), .ZN(new_n31461_));
  NOR2_X1    g29025(.A1(new_n31461_), .A2(new_n28353_), .ZN(new_n31462_));
  NAND2_X1   g29026(.A1(new_n30104_), .A2(new_n12785_), .ZN(new_n31463_));
  NAND2_X1   g29027(.A1(new_n31463_), .A2(new_n30055_), .ZN(new_n31464_));
  NAND2_X1   g29028(.A1(new_n31462_), .A2(new_n31464_), .ZN(new_n31465_));
  NOR3_X1    g29029(.A1(new_n31461_), .A2(new_n31100_), .A3(pi1154), .ZN(new_n31466_));
  NOR3_X1    g29030(.A1(new_n31461_), .A2(new_n31130_), .A3(new_n12785_), .ZN(new_n31467_));
  NAND2_X1   g29031(.A1(new_n31467_), .A2(new_n30047_), .ZN(new_n31468_));
  INV_X1     g29032(.I(new_n31468_), .ZN(new_n31469_));
  OAI21_X1   g29033(.A1(new_n31469_), .A2(new_n31466_), .B(new_n28017_), .ZN(new_n31470_));
  NOR2_X1    g29034(.A1(new_n30104_), .A2(pi1091), .ZN(new_n31471_));
  NOR2_X1    g29035(.A1(new_n31471_), .A2(pi1155), .ZN(new_n31472_));
  INV_X1     g29036(.I(new_n31472_), .ZN(new_n31473_));
  NAND2_X1   g29037(.A1(new_n30073_), .A2(pi1155), .ZN(new_n31474_));
  AOI21_X1   g29038(.A1(new_n31473_), .A2(new_n31474_), .B(pi1154), .ZN(new_n31475_));
  OAI21_X1   g29039(.A1(new_n31475_), .A2(new_n31467_), .B(new_n12742_), .ZN(new_n31476_));
  NAND4_X1   g29040(.A1(new_n31470_), .A2(pi0219), .A3(new_n31465_), .A4(new_n31476_), .ZN(new_n31477_));
  INV_X1     g29041(.I(new_n30141_), .ZN(new_n31478_));
  AOI21_X1   g29042(.A1(new_n30150_), .A2(pi1155), .B(new_n12785_), .ZN(new_n31479_));
  INV_X1     g29043(.I(new_n31479_), .ZN(new_n31480_));
  NOR2_X1    g29044(.A1(new_n31480_), .A2(new_n31478_), .ZN(new_n31481_));
  NAND2_X1   g29045(.A1(new_n30137_), .A2(new_n31101_), .ZN(new_n31482_));
  OAI21_X1   g29046(.A1(pi1155), .A2(new_n31100_), .B(new_n31482_), .ZN(new_n31483_));
  AOI21_X1   g29047(.A1(new_n31483_), .A2(new_n12785_), .B(new_n12742_), .ZN(new_n31484_));
  AOI21_X1   g29048(.A1(new_n30045_), .A2(new_n31481_), .B(new_n31466_), .ZN(new_n31485_));
  AOI21_X1   g29049(.A1(new_n31484_), .A2(new_n31485_), .B(pi0211), .ZN(new_n31486_));
  INV_X1     g29050(.I(new_n31475_), .ZN(new_n31487_));
  NOR2_X1    g29051(.A1(new_n30160_), .A2(pi1155), .ZN(new_n31488_));
  AOI22_X1   g29052(.A1(new_n30129_), .A2(pi1155), .B1(new_n31471_), .B2(new_n31488_), .ZN(new_n31489_));
  AOI21_X1   g29053(.A1(new_n31489_), .A2(new_n12785_), .B(pi1156), .ZN(new_n31490_));
  NAND2_X1   g29054(.A1(new_n31490_), .A2(new_n31487_), .ZN(new_n31491_));
  OAI21_X1   g29055(.A1(new_n31481_), .A2(new_n31491_), .B(new_n31486_), .ZN(new_n31492_));
  OAI21_X1   g29056(.A1(new_n30090_), .A2(new_n31480_), .B(new_n31484_), .ZN(new_n31493_));
  NAND2_X1   g29057(.A1(new_n31479_), .A2(new_n31102_), .ZN(new_n31494_));
  AOI21_X1   g29058(.A1(new_n31490_), .A2(new_n31494_), .B(new_n8510_), .ZN(new_n31495_));
  AOI21_X1   g29059(.A1(new_n31493_), .A2(new_n31495_), .B(pi0219), .ZN(new_n31496_));
  AOI21_X1   g29060(.A1(new_n31492_), .A2(new_n31496_), .B(pi0263), .ZN(new_n31497_));
  AOI21_X1   g29061(.A1(new_n31497_), .A2(new_n31477_), .B(new_n29996_), .ZN(new_n31498_));
  NOR2_X1    g29062(.A1(new_n30153_), .A2(pi1155), .ZN(new_n31499_));
  INV_X1     g29063(.I(new_n30103_), .ZN(new_n31500_));
  AOI21_X1   g29064(.A1(new_n30130_), .A2(new_n31500_), .B(new_n12770_), .ZN(new_n31501_));
  OAI21_X1   g29065(.A1(new_n31501_), .A2(new_n31499_), .B(new_n12785_), .ZN(new_n31502_));
  OAI21_X1   g29066(.A1(new_n31502_), .A2(new_n30151_), .B(pi1156), .ZN(new_n31503_));
  NOR3_X1    g29067(.A1(new_n30134_), .A2(new_n30176_), .A3(new_n12785_), .ZN(new_n31504_));
  OAI21_X1   g29068(.A1(new_n31504_), .A2(new_n31503_), .B(new_n8510_), .ZN(new_n31505_));
  NOR3_X1    g29069(.A1(new_n31504_), .A2(pi1156), .A3(new_n31281_), .ZN(new_n31506_));
  AND2_X2    g29070(.A1(new_n31506_), .A2(new_n31502_), .Z(new_n31507_));
  OAI21_X1   g29071(.A1(new_n31507_), .A2(new_n31505_), .B(new_n8807_), .ZN(new_n31508_));
  NOR2_X1    g29072(.A1(new_n30132_), .A2(new_n12770_), .ZN(new_n31509_));
  NOR2_X1    g29073(.A1(new_n30119_), .A2(pi1155), .ZN(new_n31510_));
  OAI21_X1   g29074(.A1(new_n31509_), .A2(new_n31510_), .B(pi1154), .ZN(new_n31511_));
  NOR2_X1    g29075(.A1(new_n31275_), .A2(new_n12770_), .ZN(new_n31512_));
  OAI21_X1   g29076(.A1(new_n31512_), .A2(new_n31499_), .B(new_n12785_), .ZN(new_n31513_));
  INV_X1     g29077(.I(new_n31513_), .ZN(new_n31514_));
  NAND2_X1   g29078(.A1(new_n31506_), .A2(new_n31513_), .ZN(new_n31515_));
  AOI22_X1   g29079(.A1(new_n31515_), .A2(new_n12742_), .B1(new_n31274_), .B2(new_n31514_), .ZN(new_n31516_));
  AOI21_X1   g29080(.A1(new_n31516_), .A2(new_n31511_), .B(new_n8510_), .ZN(new_n31517_));
  AOI21_X1   g29081(.A1(pi1155), .A2(new_n30104_), .B(new_n30060_), .ZN(new_n31518_));
  AOI21_X1   g29082(.A1(new_n30069_), .A2(new_n31271_), .B(new_n31518_), .ZN(new_n31519_));
  NAND2_X1   g29083(.A1(new_n31519_), .A2(new_n31500_), .ZN(new_n31520_));
  NAND2_X1   g29084(.A1(new_n31520_), .A2(new_n12742_), .ZN(new_n31521_));
  OAI21_X1   g29085(.A1(new_n31519_), .A2(new_n31432_), .B(pi0219), .ZN(new_n31522_));
  OAI21_X1   g29086(.A1(new_n31518_), .A2(new_n12785_), .B(new_n28013_), .ZN(new_n31523_));
  NAND2_X1   g29087(.A1(new_n31114_), .A2(new_n12770_), .ZN(new_n31524_));
  OAI21_X1   g29088(.A1(new_n12770_), .A2(new_n31267_), .B(new_n31524_), .ZN(new_n31525_));
  AOI21_X1   g29089(.A1(new_n31525_), .A2(new_n12785_), .B(new_n31523_), .ZN(new_n31526_));
  NOR2_X1    g29090(.A1(new_n31522_), .A2(new_n31526_), .ZN(new_n31527_));
  AOI21_X1   g29091(.A1(new_n31527_), .A2(new_n31521_), .B(new_n31416_), .ZN(new_n31528_));
  OAI21_X1   g29092(.A1(new_n31517_), .A2(new_n31508_), .B(new_n31528_), .ZN(new_n31529_));
  AOI22_X1   g29093(.A1(new_n31529_), .A2(new_n31498_), .B1(new_n29996_), .B2(new_n31460_), .ZN(new_n31530_));
  NAND3_X1   g29094(.A1(new_n28353_), .A2(pi0219), .A3(pi1091), .ZN(new_n31531_));
  AOI22_X1   g29095(.A1(new_n30020_), .A2(new_n28014_), .B1(pi1154), .B2(new_n31032_), .ZN(new_n31532_));
  NAND2_X1   g29096(.A1(new_n31084_), .A2(new_n31532_), .ZN(new_n31533_));
  NAND3_X1   g29097(.A1(new_n31090_), .A2(new_n31533_), .A3(pi0263), .ZN(new_n31534_));
  OAI21_X1   g29098(.A1(new_n31208_), .A2(pi0211), .B(new_n28354_), .ZN(new_n31535_));
  AOI21_X1   g29099(.A1(new_n30037_), .A2(pi0211), .B(new_n31535_), .ZN(new_n31536_));
  OAI21_X1   g29100(.A1(new_n31536_), .A2(new_n30011_), .B(new_n8807_), .ZN(new_n31537_));
  NAND3_X1   g29101(.A1(new_n31257_), .A2(new_n31537_), .A3(new_n31416_), .ZN(new_n31538_));
  AOI21_X1   g29102(.A1(new_n31534_), .A2(new_n31538_), .B(new_n29996_), .ZN(new_n31539_));
  OAI21_X1   g29103(.A1(new_n31457_), .A2(new_n29995_), .B(po1038), .ZN(new_n31540_));
  AOI21_X1   g29104(.A1(new_n31539_), .A2(new_n31531_), .B(new_n31540_), .ZN(new_n31541_));
  AOI21_X1   g29105(.A1(new_n31530_), .A2(new_n6643_), .B(new_n31541_), .ZN(new_n31542_));
  AOI21_X1   g29106(.A1(new_n31542_), .A2(new_n29933_), .B(pi0230), .ZN(new_n31543_));
  AOI22_X1   g29107(.A1(new_n31543_), .A2(new_n31459_), .B1(new_n31413_), .B2(new_n31415_), .ZN(po0420));
  NOR2_X1    g29108(.A1(new_n3926_), .A2(pi0199), .ZN(new_n31545_));
  NOR3_X1    g29109(.A1(new_n28797_), .A2(new_n31545_), .A3(pi0200), .ZN(new_n31546_));
  NOR3_X1    g29110(.A1(new_n25319_), .A2(new_n28029_), .A3(new_n31546_), .ZN(new_n31547_));
  AOI21_X1   g29111(.A1(new_n8510_), .A2(new_n3926_), .B(new_n28078_), .ZN(new_n31548_));
  OAI21_X1   g29112(.A1(new_n31548_), .A2(pi0219), .B(new_n30213_), .ZN(new_n31549_));
  NOR2_X1    g29113(.A1(new_n12618_), .A2(new_n31549_), .ZN(new_n31550_));
  OAI21_X1   g29114(.A1(new_n31547_), .A2(new_n31550_), .B(pi0230), .ZN(new_n31551_));
  NOR2_X1    g29115(.A1(new_n30003_), .A2(pi0264), .ZN(new_n31552_));
  AND2_X2    g29116(.A1(new_n30003_), .A2(pi0796), .Z(new_n31553_));
  OAI21_X1   g29117(.A1(new_n31553_), .A2(new_n31552_), .B(new_n3022_), .ZN(new_n31554_));
  NOR2_X1    g29118(.A1(new_n3022_), .A2(new_n3768_), .ZN(new_n31555_));
  INV_X1     g29119(.I(new_n31555_), .ZN(new_n31556_));
  NAND3_X1   g29120(.A1(new_n31554_), .A2(pi0211), .A3(new_n31556_), .ZN(new_n31557_));
  NOR2_X1    g29121(.A1(new_n3022_), .A2(new_n3926_), .ZN(new_n31558_));
  INV_X1     g29122(.I(new_n31558_), .ZN(new_n31559_));
  NAND3_X1   g29123(.A1(new_n31554_), .A2(new_n8510_), .A3(new_n31559_), .ZN(new_n31560_));
  AOI21_X1   g29124(.A1(new_n31557_), .A2(new_n31560_), .B(pi0219), .ZN(new_n31561_));
  INV_X1     g29125(.I(pi0264), .ZN(new_n31562_));
  NAND2_X1   g29126(.A1(new_n30015_), .A2(new_n31562_), .ZN(new_n31563_));
  NAND2_X1   g29127(.A1(new_n30014_), .A2(pi0796), .ZN(new_n31564_));
  AOI21_X1   g29128(.A1(new_n31563_), .A2(new_n31564_), .B(pi1091), .ZN(new_n31565_));
  OAI21_X1   g29129(.A1(new_n28068_), .A2(new_n31033_), .B(pi0219), .ZN(new_n31566_));
  NOR2_X1    g29130(.A1(new_n31565_), .A2(new_n31566_), .ZN(new_n31567_));
  NOR3_X1    g29131(.A1(new_n31561_), .A2(new_n12618_), .A3(new_n31567_), .ZN(new_n31568_));
  NAND3_X1   g29132(.A1(new_n31554_), .A2(pi0200), .A3(new_n31556_), .ZN(new_n31569_));
  NAND3_X1   g29133(.A1(new_n31554_), .A2(new_n8531_), .A3(new_n31559_), .ZN(new_n31570_));
  NAND2_X1   g29134(.A1(new_n31569_), .A2(new_n31570_), .ZN(new_n31571_));
  NOR2_X1    g29135(.A1(new_n3022_), .A2(new_n3605_), .ZN(new_n31572_));
  NAND2_X1   g29136(.A1(new_n31572_), .A2(new_n8531_), .ZN(new_n31573_));
  NAND2_X1   g29137(.A1(new_n31573_), .A2(pi0199), .ZN(new_n31574_));
  OAI21_X1   g29138(.A1(new_n31565_), .A2(new_n31574_), .B(new_n12618_), .ZN(new_n31575_));
  AOI21_X1   g29139(.A1(new_n31571_), .A2(new_n8525_), .B(new_n31575_), .ZN(new_n31576_));
  OAI21_X1   g29140(.A1(new_n31568_), .A2(new_n31576_), .B(new_n27999_), .ZN(new_n31577_));
  NAND2_X1   g29141(.A1(new_n31577_), .A2(new_n31551_), .ZN(po0421));
  AOI21_X1   g29142(.A1(new_n8510_), .A2(new_n3768_), .B(new_n28061_), .ZN(new_n31579_));
  NOR2_X1    g29143(.A1(new_n31579_), .A2(pi0219), .ZN(new_n31580_));
  NOR2_X1    g29144(.A1(new_n31580_), .A2(new_n29882_), .ZN(new_n31581_));
  INV_X1     g29145(.I(new_n29859_), .ZN(new_n31582_));
  OAI21_X1   g29146(.A1(new_n28028_), .A2(new_n31582_), .B(new_n28036_), .ZN(new_n31583_));
  AOI21_X1   g29147(.A1(new_n12618_), .A2(new_n31583_), .B(new_n27999_), .ZN(new_n31584_));
  OAI21_X1   g29148(.A1(new_n12618_), .A2(new_n31581_), .B(new_n31584_), .ZN(new_n31585_));
  NAND2_X1   g29149(.A1(new_n30004_), .A2(new_n2452_), .ZN(new_n31586_));
  NAND2_X1   g29150(.A1(new_n30003_), .A2(pi0819), .ZN(new_n31587_));
  AOI21_X1   g29151(.A1(new_n31586_), .A2(new_n31587_), .B(pi1091), .ZN(new_n31588_));
  NOR3_X1    g29152(.A1(new_n31588_), .A2(new_n8510_), .A3(new_n31572_), .ZN(new_n31589_));
  NOR3_X1    g29153(.A1(new_n31588_), .A2(pi0211), .A3(new_n31555_), .ZN(new_n31590_));
  OAI21_X1   g29154(.A1(new_n31589_), .A2(new_n31590_), .B(new_n8807_), .ZN(new_n31591_));
  NOR2_X1    g29155(.A1(new_n30014_), .A2(pi0265), .ZN(new_n31592_));
  AND2_X2    g29156(.A1(new_n30014_), .A2(pi0819), .Z(new_n31593_));
  OAI21_X1   g29157(.A1(new_n31593_), .A2(new_n31592_), .B(new_n3022_), .ZN(new_n31594_));
  OAI21_X1   g29158(.A1(new_n8807_), .A2(new_n31032_), .B(new_n29883_), .ZN(new_n31595_));
  AOI21_X1   g29159(.A1(new_n31594_), .A2(new_n31595_), .B(new_n12618_), .ZN(new_n31596_));
  NOR3_X1    g29160(.A1(new_n31588_), .A2(new_n8531_), .A3(new_n31572_), .ZN(new_n31597_));
  NOR3_X1    g29161(.A1(new_n31588_), .A2(pi0200), .A3(new_n31555_), .ZN(new_n31598_));
  OAI21_X1   g29162(.A1(new_n31597_), .A2(new_n31598_), .B(new_n8525_), .ZN(new_n31599_));
  NOR2_X1    g29163(.A1(new_n3022_), .A2(new_n2446_), .ZN(new_n31600_));
  AOI21_X1   g29164(.A1(new_n31600_), .A2(new_n8531_), .B(new_n8525_), .ZN(new_n31601_));
  AOI21_X1   g29165(.A1(new_n31594_), .A2(new_n31601_), .B(new_n25319_), .ZN(new_n31602_));
  AOI22_X1   g29166(.A1(new_n31591_), .A2(new_n31596_), .B1(new_n31599_), .B2(new_n31602_), .ZN(new_n31603_));
  OAI21_X1   g29167(.A1(new_n31603_), .A2(pi0230), .B(new_n31585_), .ZN(po0422));
  INV_X1     g29168(.I(new_n31056_), .ZN(new_n31605_));
  NAND2_X1   g29169(.A1(new_n8510_), .A2(pi1136), .ZN(new_n31606_));
  AOI22_X1   g29170(.A1(new_n31606_), .A2(pi0219), .B1(pi0211), .B2(new_n4888_), .ZN(new_n31607_));
  NAND2_X1   g29171(.A1(new_n31607_), .A2(new_n31605_), .ZN(new_n31608_));
  NAND2_X1   g29172(.A1(new_n8525_), .A2(pi1135), .ZN(new_n31609_));
  NAND2_X1   g29173(.A1(new_n31609_), .A2(pi0200), .ZN(new_n31610_));
  OAI21_X1   g29174(.A1(new_n8525_), .A2(new_n4724_), .B(new_n8531_), .ZN(new_n31611_));
  NAND3_X1   g29175(.A1(new_n31610_), .A2(new_n2628_), .A3(new_n31611_), .ZN(new_n31612_));
  OAI22_X1   g29176(.A1(new_n12618_), .A2(new_n31608_), .B1(po1038), .B2(new_n31612_), .ZN(new_n31613_));
  INV_X1     g29177(.I(pi0948), .ZN(new_n31614_));
  NOR2_X1    g29178(.A1(new_n30015_), .A2(new_n31614_), .ZN(new_n31615_));
  NOR2_X1    g29179(.A1(new_n30014_), .A2(new_n4727_), .ZN(new_n31616_));
  OAI21_X1   g29180(.A1(new_n31615_), .A2(new_n31616_), .B(new_n3022_), .ZN(new_n31617_));
  INV_X1     g29181(.I(new_n31617_), .ZN(new_n31618_));
  NOR2_X1    g29182(.A1(new_n31618_), .A2(new_n8525_), .ZN(new_n31619_));
  NOR2_X1    g29183(.A1(new_n31619_), .A2(new_n8531_), .ZN(new_n31620_));
  NOR2_X1    g29184(.A1(new_n30004_), .A2(new_n31614_), .ZN(new_n31621_));
  NOR2_X1    g29185(.A1(new_n30003_), .A2(new_n4727_), .ZN(new_n31622_));
  OAI21_X1   g29186(.A1(new_n31621_), .A2(new_n31622_), .B(new_n3022_), .ZN(new_n31623_));
  AND2_X2    g29187(.A1(new_n31623_), .A2(new_n8525_), .Z(new_n31624_));
  OAI21_X1   g29188(.A1(new_n3022_), .A2(new_n4888_), .B(new_n31624_), .ZN(new_n31625_));
  NAND2_X1   g29189(.A1(new_n31625_), .A2(new_n31620_), .ZN(new_n31626_));
  NAND2_X1   g29190(.A1(pi1091), .A2(pi1136), .ZN(new_n31627_));
  AOI21_X1   g29191(.A1(new_n31619_), .A2(new_n31627_), .B(new_n31624_), .ZN(new_n31628_));
  NAND2_X1   g29192(.A1(new_n31628_), .A2(new_n8531_), .ZN(new_n31629_));
  AOI21_X1   g29193(.A1(new_n31629_), .A2(new_n31626_), .B(new_n25319_), .ZN(new_n31630_));
  OAI21_X1   g29194(.A1(new_n31627_), .A2(pi0211), .B(pi0219), .ZN(new_n31631_));
  OAI21_X1   g29195(.A1(new_n31618_), .A2(new_n31631_), .B(new_n25319_), .ZN(new_n31632_));
  NAND2_X1   g29196(.A1(new_n31623_), .A2(new_n8807_), .ZN(new_n31633_));
  AOI21_X1   g29197(.A1(pi1135), .A2(new_n31417_), .B(new_n31633_), .ZN(new_n31634_));
  OAI21_X1   g29198(.A1(new_n31634_), .A2(new_n31632_), .B(new_n27999_), .ZN(new_n31635_));
  OAI22_X1   g29199(.A1(new_n31630_), .A2(new_n31635_), .B1(new_n27999_), .B2(new_n31613_), .ZN(new_n31636_));
  AOI21_X1   g29200(.A1(new_n8525_), .A2(pi1091), .B(new_n31628_), .ZN(new_n31637_));
  OAI21_X1   g29201(.A1(new_n31637_), .A2(pi0200), .B(new_n31626_), .ZN(new_n31638_));
  AOI21_X1   g29202(.A1(pi0211), .A2(new_n4888_), .B(new_n3022_), .ZN(new_n31639_));
  NOR2_X1    g29203(.A1(new_n31633_), .A2(new_n31639_), .ZN(new_n31640_));
  OAI21_X1   g29204(.A1(new_n31632_), .A2(new_n31640_), .B(new_n27999_), .ZN(new_n31641_));
  AOI21_X1   g29205(.A1(new_n31638_), .A2(new_n12618_), .B(new_n31641_), .ZN(new_n31642_));
  OAI21_X1   g29206(.A1(new_n8525_), .A2(pi1136), .B(new_n31610_), .ZN(new_n31643_));
  NOR2_X1    g29207(.A1(new_n12618_), .A2(new_n31607_), .ZN(new_n31644_));
  AOI21_X1   g29208(.A1(new_n12618_), .A2(new_n31643_), .B(new_n31644_), .ZN(new_n31645_));
  OAI21_X1   g29209(.A1(new_n31645_), .A2(new_n27999_), .B(pi1134), .ZN(new_n31646_));
  OAI22_X1   g29210(.A1(new_n31642_), .A2(new_n31646_), .B1(new_n31636_), .B2(pi1134), .ZN(po0423));
  AOI21_X1   g29211(.A1(new_n12785_), .A2(new_n28102_), .B(new_n28100_), .ZN(new_n31648_));
  NAND2_X1   g29212(.A1(new_n31648_), .A2(new_n28389_), .ZN(new_n31649_));
  NAND2_X1   g29213(.A1(new_n31649_), .A2(new_n8807_), .ZN(new_n31650_));
  AOI21_X1   g29214(.A1(new_n8525_), .A2(pi1154), .B(new_n8531_), .ZN(new_n31651_));
  OR3_X2     g29215(.A1(new_n28449_), .A2(new_n28291_), .A3(new_n31651_), .Z(new_n31652_));
  NAND3_X1   g29216(.A1(new_n31652_), .A2(pi0219), .A3(new_n28282_), .ZN(new_n31653_));
  AOI21_X1   g29217(.A1(new_n31650_), .A2(new_n31653_), .B(pi0211), .ZN(new_n31654_));
  OAI21_X1   g29218(.A1(new_n28448_), .A2(new_n28449_), .B(pi0219), .ZN(new_n31655_));
  INV_X1     g29219(.I(new_n29097_), .ZN(new_n31656_));
  NOR2_X1    g29220(.A1(new_n28826_), .A2(new_n12841_), .ZN(new_n31657_));
  AOI21_X1   g29221(.A1(new_n31657_), .A2(new_n12770_), .B(pi1154), .ZN(new_n31658_));
  OAI22_X1   g29222(.A1(new_n31658_), .A2(new_n28439_), .B1(new_n12770_), .B2(new_n31656_), .ZN(new_n31659_));
  AOI21_X1   g29223(.A1(new_n31659_), .A2(new_n31655_), .B(new_n8510_), .ZN(new_n31660_));
  OR3_X2     g29224(.A1(new_n31660_), .A2(po1038), .A3(new_n31654_), .Z(new_n31661_));
  NOR2_X1    g29225(.A1(new_n28005_), .A2(pi0219), .ZN(new_n31662_));
  AOI22_X1   g29226(.A1(new_n31662_), .A2(new_n31297_), .B1(new_n28726_), .B2(pi0219), .ZN(new_n31663_));
  AOI21_X1   g29227(.A1(new_n31663_), .A2(po1038), .B(new_n27999_), .ZN(new_n31664_));
  NOR2_X1    g29228(.A1(new_n3022_), .A2(pi1155), .ZN(new_n31665_));
  AOI21_X1   g29229(.A1(new_n28440_), .A2(new_n31665_), .B(new_n31297_), .ZN(new_n31666_));
  NAND3_X1   g29230(.A1(new_n31067_), .A2(pi1091), .A3(new_n31421_), .ZN(new_n31667_));
  NAND2_X1   g29231(.A1(new_n31667_), .A2(new_n31666_), .ZN(new_n31668_));
  OAI21_X1   g29232(.A1(new_n31649_), .A2(new_n3022_), .B(new_n8510_), .ZN(new_n31669_));
  NAND3_X1   g29233(.A1(new_n31668_), .A2(new_n31669_), .A3(new_n8807_), .ZN(new_n31670_));
  NAND2_X1   g29234(.A1(new_n31667_), .A2(pi1154), .ZN(new_n31671_));
  NOR3_X1    g29235(.A1(new_n28437_), .A2(pi0199), .A3(pi0299), .ZN(new_n31672_));
  AOI21_X1   g29236(.A1(new_n31665_), .A2(new_n31672_), .B(new_n31671_), .ZN(new_n31673_));
  NOR4_X1    g29237(.A1(new_n28450_), .A2(new_n12785_), .A3(new_n12770_), .A4(new_n28465_), .ZN(new_n31674_));
  OAI21_X1   g29238(.A1(new_n31673_), .A2(new_n31674_), .B(pi0211), .ZN(new_n31675_));
  INV_X1     g29239(.I(new_n31208_), .ZN(new_n31676_));
  NOR2_X1    g29240(.A1(new_n28152_), .A2(new_n31676_), .ZN(new_n31677_));
  AOI21_X1   g29241(.A1(new_n29098_), .A2(new_n31677_), .B(pi0211), .ZN(new_n31678_));
  OAI21_X1   g29242(.A1(new_n31673_), .A2(new_n12785_), .B(new_n31678_), .ZN(new_n31679_));
  NAND3_X1   g29243(.A1(new_n31675_), .A2(new_n31679_), .A3(pi0219), .ZN(new_n31680_));
  NAND2_X1   g29244(.A1(new_n29097_), .A2(pi1091), .ZN(new_n31681_));
  NOR2_X1    g29245(.A1(new_n28381_), .A2(pi1155), .ZN(new_n31682_));
  OAI21_X1   g29246(.A1(new_n31682_), .A2(new_n31681_), .B(pi0211), .ZN(new_n31683_));
  OAI21_X1   g29247(.A1(new_n31683_), .A2(pi1154), .B(new_n29990_), .ZN(new_n31684_));
  AOI21_X1   g29248(.A1(new_n31680_), .A2(new_n31670_), .B(new_n31684_), .ZN(new_n31685_));
  NOR2_X1    g29249(.A1(new_n31657_), .A2(new_n31676_), .ZN(new_n31686_));
  INV_X1     g29250(.I(new_n29938_), .ZN(new_n31687_));
  NAND2_X1   g29251(.A1(new_n31687_), .A2(new_n28284_), .ZN(new_n31688_));
  AOI21_X1   g29252(.A1(new_n31688_), .A2(new_n31686_), .B(new_n8510_), .ZN(new_n31689_));
  NAND2_X1   g29253(.A1(new_n28440_), .A2(new_n12770_), .ZN(new_n31690_));
  AOI22_X1   g29254(.A1(new_n28225_), .A2(new_n31690_), .B1(pi0219), .B2(pi0299), .ZN(new_n31691_));
  NAND2_X1   g29255(.A1(new_n28450_), .A2(pi1155), .ZN(new_n31692_));
  NAND3_X1   g29256(.A1(new_n31692_), .A2(pi1091), .A3(pi1154), .ZN(new_n31693_));
  OAI21_X1   g29257(.A1(new_n31691_), .A2(new_n31693_), .B(new_n31689_), .ZN(new_n31694_));
  NOR3_X1    g29258(.A1(new_n29100_), .A2(new_n31676_), .A3(new_n31657_), .ZN(new_n31695_));
  NOR3_X1    g29259(.A1(new_n31671_), .A2(new_n3022_), .A3(new_n31672_), .ZN(new_n31696_));
  NOR3_X1    g29260(.A1(new_n31696_), .A2(new_n8807_), .A3(new_n31695_), .ZN(new_n31697_));
  INV_X1     g29261(.I(new_n31220_), .ZN(new_n31698_));
  NAND3_X1   g29262(.A1(new_n31698_), .A2(new_n12770_), .A3(new_n31048_), .ZN(new_n31699_));
  NAND3_X1   g29263(.A1(new_n31068_), .A2(pi1155), .A3(new_n31420_), .ZN(new_n31700_));
  NAND3_X1   g29264(.A1(new_n31699_), .A2(new_n31700_), .A3(pi1154), .ZN(new_n31701_));
  NAND2_X1   g29265(.A1(new_n31687_), .A2(new_n12841_), .ZN(new_n31702_));
  NAND3_X1   g29266(.A1(new_n31702_), .A2(pi1155), .A3(new_n31068_), .ZN(new_n31703_));
  NAND2_X1   g29267(.A1(new_n31682_), .A2(pi1091), .ZN(new_n31704_));
  NAND3_X1   g29268(.A1(new_n31703_), .A2(new_n12785_), .A3(new_n31704_), .ZN(new_n31705_));
  AOI21_X1   g29269(.A1(new_n31705_), .A2(new_n31701_), .B(pi0219), .ZN(new_n31706_));
  OAI21_X1   g29270(.A1(new_n31697_), .A2(new_n31706_), .B(new_n8510_), .ZN(new_n31707_));
  AOI21_X1   g29271(.A1(new_n31707_), .A2(new_n31694_), .B(new_n29990_), .ZN(new_n31708_));
  NOR2_X1    g29272(.A1(new_n31685_), .A2(new_n31708_), .ZN(new_n31709_));
  NOR2_X1    g29273(.A1(new_n31709_), .A2(po1038), .ZN(new_n31710_));
  NOR2_X1    g29274(.A1(pi0267), .A2(pi1091), .ZN(new_n31711_));
  NOR2_X1    g29275(.A1(new_n31663_), .A2(new_n3022_), .ZN(new_n31712_));
  NOR3_X1    g29276(.A1(new_n31712_), .A2(new_n6643_), .A3(new_n31711_), .ZN(new_n31713_));
  OAI21_X1   g29277(.A1(new_n31710_), .A2(new_n31713_), .B(new_n29934_), .ZN(new_n31714_));
  INV_X1     g29278(.I(new_n31501_), .ZN(new_n31715_));
  NAND2_X1   g29279(.A1(new_n30060_), .A2(pi1153), .ZN(new_n31716_));
  AOI21_X1   g29280(.A1(new_n31274_), .A2(new_n31716_), .B(new_n12770_), .ZN(new_n31717_));
  NOR2_X1    g29281(.A1(new_n30160_), .A2(new_n12841_), .ZN(new_n31718_));
  AOI21_X1   g29282(.A1(new_n30130_), .A2(new_n31500_), .B(pi1153), .ZN(new_n31719_));
  OAI21_X1   g29283(.A1(new_n31719_), .A2(new_n31718_), .B(new_n12770_), .ZN(new_n31720_));
  AOI21_X1   g29284(.A1(new_n31715_), .A2(new_n31720_), .B(new_n31717_), .ZN(new_n31721_));
  NAND2_X1   g29285(.A1(new_n31721_), .A2(pi1154), .ZN(new_n31722_));
  NOR4_X1    g29286(.A1(new_n31718_), .A2(new_n31109_), .A3(pi1155), .A4(new_n30058_), .ZN(new_n31723_));
  NOR2_X1    g29287(.A1(new_n31717_), .A2(new_n31723_), .ZN(new_n31724_));
  AOI21_X1   g29288(.A1(new_n31724_), .A2(new_n12785_), .B(pi0211), .ZN(new_n31725_));
  AOI21_X1   g29289(.A1(new_n31722_), .A2(new_n31725_), .B(pi0267), .ZN(new_n31726_));
  NOR2_X1    g29290(.A1(new_n30107_), .A2(new_n31262_), .ZN(new_n31727_));
  NOR2_X1    g29291(.A1(new_n31727_), .A2(pi1155), .ZN(new_n31728_));
  AOI21_X1   g29292(.A1(new_n31728_), .A2(new_n31276_), .B(new_n8510_), .ZN(new_n31729_));
  NAND2_X1   g29293(.A1(new_n31160_), .A2(new_n12785_), .ZN(new_n31730_));
  AOI21_X1   g29294(.A1(new_n31730_), .A2(pi1155), .B(new_n30120_), .ZN(new_n31731_));
  OAI21_X1   g29295(.A1(new_n31102_), .A2(new_n31139_), .B(new_n30073_), .ZN(new_n31732_));
  AOI21_X1   g29296(.A1(new_n31732_), .A2(new_n30082_), .B(new_n12770_), .ZN(new_n31733_));
  AOI21_X1   g29297(.A1(new_n31733_), .A2(new_n31267_), .B(new_n12785_), .ZN(new_n31734_));
  OAI21_X1   g29298(.A1(new_n31734_), .A2(new_n31731_), .B(new_n31729_), .ZN(new_n31735_));
  AOI21_X1   g29299(.A1(new_n30072_), .A2(pi1154), .B(new_n12770_), .ZN(new_n31736_));
  OAI21_X1   g29300(.A1(new_n30130_), .A2(new_n31283_), .B(new_n31736_), .ZN(new_n31737_));
  NOR2_X1    g29301(.A1(new_n31139_), .A2(pi1154), .ZN(new_n31738_));
  AOI21_X1   g29302(.A1(new_n31738_), .A2(new_n31478_), .B(pi1155), .ZN(new_n31739_));
  AOI21_X1   g29303(.A1(new_n12841_), .A2(new_n30172_), .B(new_n30149_), .ZN(new_n31740_));
  NAND2_X1   g29304(.A1(new_n31740_), .A2(pi1154), .ZN(new_n31741_));
  NAND2_X1   g29305(.A1(new_n31739_), .A2(new_n31741_), .ZN(new_n31742_));
  NAND3_X1   g29306(.A1(new_n31742_), .A2(new_n8510_), .A3(new_n31737_), .ZN(new_n31743_));
  NAND2_X1   g29307(.A1(new_n31134_), .A2(pi1155), .ZN(new_n31744_));
  OAI21_X1   g29308(.A1(new_n31482_), .A2(new_n31744_), .B(pi1154), .ZN(new_n31745_));
  NOR3_X1    g29309(.A1(new_n30129_), .A2(pi1155), .A3(new_n31740_), .ZN(new_n31746_));
  NOR2_X1    g29310(.A1(new_n31745_), .A2(new_n31746_), .ZN(new_n31747_));
  NOR4_X1    g29311(.A1(new_n31739_), .A2(pi1154), .A3(new_n30089_), .A4(new_n31139_), .ZN(new_n31748_));
  OAI21_X1   g29312(.A1(new_n31748_), .A2(new_n31747_), .B(pi0211), .ZN(new_n31749_));
  NAND3_X1   g29313(.A1(new_n31749_), .A2(pi0267), .A3(new_n31743_), .ZN(new_n31750_));
  NAND2_X1   g29314(.A1(new_n31750_), .A2(new_n8807_), .ZN(new_n31751_));
  AOI21_X1   g29315(.A1(new_n31726_), .A2(new_n31735_), .B(new_n31751_), .ZN(new_n31752_));
  NAND2_X1   g29316(.A1(new_n31463_), .A2(new_n30072_), .ZN(new_n31753_));
  NAND4_X1   g29317(.A1(new_n31106_), .A2(pi1155), .A3(new_n31134_), .A4(new_n31753_), .ZN(new_n31754_));
  NAND3_X1   g29318(.A1(new_n31096_), .A2(new_n12785_), .A3(new_n31130_), .ZN(new_n31755_));
  NAND2_X1   g29319(.A1(new_n31732_), .A2(pi1154), .ZN(new_n31756_));
  NAND3_X1   g29320(.A1(new_n31756_), .A2(new_n12770_), .A3(new_n31755_), .ZN(new_n31757_));
  NAND3_X1   g29321(.A1(new_n31754_), .A2(pi0267), .A3(new_n31757_), .ZN(new_n31758_));
  OAI21_X1   g29322(.A1(new_n12785_), .A2(new_n31264_), .B(new_n31728_), .ZN(new_n31759_));
  INV_X1     g29323(.I(new_n31716_), .ZN(new_n31760_));
  NOR3_X1    g29324(.A1(new_n31114_), .A2(new_n31760_), .A3(new_n28726_), .ZN(new_n31761_));
  OAI21_X1   g29325(.A1(new_n12785_), .A2(new_n31267_), .B(new_n31761_), .ZN(new_n31762_));
  NOR4_X1    g29326(.A1(new_n30068_), .A2(new_n31298_), .A3(new_n12785_), .A4(new_n12770_), .ZN(new_n31763_));
  NOR3_X1    g29327(.A1(new_n31727_), .A2(new_n31289_), .A3(pi1154), .ZN(new_n31764_));
  OAI21_X1   g29328(.A1(new_n31763_), .A2(new_n31764_), .B(pi0211), .ZN(new_n31765_));
  NAND4_X1   g29329(.A1(new_n31765_), .A2(new_n29990_), .A3(new_n31759_), .A4(new_n31762_), .ZN(new_n31766_));
  AOI21_X1   g29330(.A1(new_n31766_), .A2(new_n31758_), .B(new_n8807_), .ZN(new_n31767_));
  NOR3_X1    g29331(.A1(new_n31752_), .A2(new_n29994_), .A3(new_n31767_), .ZN(new_n31768_));
  NOR3_X1    g29332(.A1(new_n31685_), .A2(new_n29993_), .A3(new_n31708_), .ZN(new_n31769_));
  OAI21_X1   g29333(.A1(new_n31768_), .A2(new_n31769_), .B(new_n6643_), .ZN(new_n31770_));
  AOI21_X1   g29334(.A1(new_n29994_), .A2(new_n31711_), .B(new_n31712_), .ZN(new_n31771_));
  NAND2_X1   g29335(.A1(new_n30022_), .A2(new_n29990_), .ZN(new_n31772_));
  OAI21_X1   g29336(.A1(new_n31772_), .A2(new_n31089_), .B(new_n29993_), .ZN(new_n31773_));
  INV_X1     g29337(.I(new_n31257_), .ZN(new_n31774_));
  NOR3_X1    g29338(.A1(new_n31774_), .A2(new_n29990_), .A3(new_n31255_), .ZN(new_n31775_));
  OAI21_X1   g29339(.A1(new_n31773_), .A2(new_n31775_), .B(new_n31771_), .ZN(new_n31776_));
  AOI21_X1   g29340(.A1(new_n31776_), .A2(po1038), .B(new_n29934_), .ZN(new_n31777_));
  AOI21_X1   g29341(.A1(new_n31770_), .A2(new_n31777_), .B(pi0230), .ZN(new_n31778_));
  AOI22_X1   g29342(.A1(new_n31778_), .A2(new_n31714_), .B1(new_n31661_), .B2(new_n31664_), .ZN(po0424));
  NOR2_X1    g29343(.A1(new_n12618_), .A2(pi0211), .ZN(new_n31780_));
  AOI21_X1   g29344(.A1(new_n6643_), .A2(new_n8761_), .B(new_n31780_), .ZN(new_n31781_));
  INV_X1     g29345(.I(new_n31781_), .ZN(new_n31782_));
  OAI21_X1   g29346(.A1(new_n31782_), .A2(pi1151), .B(pi1150), .ZN(new_n31783_));
  NOR2_X1    g29347(.A1(new_n25319_), .A2(pi0199), .ZN(new_n31784_));
  NOR2_X1    g29348(.A1(new_n31784_), .A2(new_n29459_), .ZN(new_n31785_));
  NAND2_X1   g29349(.A1(new_n31782_), .A2(pi1152), .ZN(new_n31786_));
  AOI21_X1   g29350(.A1(new_n31785_), .A2(new_n31786_), .B(new_n31783_), .ZN(new_n31787_));
  NOR2_X1    g29351(.A1(new_n12618_), .A2(new_n31058_), .ZN(new_n31788_));
  AOI21_X1   g29352(.A1(new_n12618_), .A2(new_n28153_), .B(new_n31788_), .ZN(new_n31789_));
  INV_X1     g29353(.I(new_n31789_), .ZN(new_n31790_));
  NOR3_X1    g29354(.A1(new_n31790_), .A2(new_n29035_), .A3(new_n28422_), .ZN(new_n31791_));
  NOR2_X1    g29355(.A1(new_n6643_), .A2(new_n9218_), .ZN(new_n31792_));
  AOI21_X1   g29356(.A1(new_n6643_), .A2(new_n9221_), .B(new_n31792_), .ZN(new_n31793_));
  AOI21_X1   g29357(.A1(new_n31793_), .A2(pi1151), .B(pi1152), .ZN(new_n31794_));
  NOR2_X1    g29358(.A1(new_n31192_), .A2(pi1151), .ZN(new_n31795_));
  NOR4_X1    g29359(.A1(new_n31791_), .A2(pi1150), .A3(new_n31794_), .A4(new_n31795_), .ZN(new_n31796_));
  NOR2_X1    g29360(.A1(new_n31787_), .A2(new_n31796_), .ZN(new_n31797_));
  NAND2_X1   g29361(.A1(new_n31787_), .A2(pi1152), .ZN(new_n31798_));
  AOI21_X1   g29362(.A1(new_n31798_), .A2(pi1091), .B(new_n29927_), .ZN(new_n31799_));
  INV_X1     g29363(.I(new_n31796_), .ZN(new_n31800_));
  OAI21_X1   g29364(.A1(new_n29927_), .A2(new_n28422_), .B(new_n31787_), .ZN(new_n31801_));
  AOI21_X1   g29365(.A1(new_n31801_), .A2(new_n31800_), .B(new_n3022_), .ZN(new_n31802_));
  OAI21_X1   g29366(.A1(new_n31802_), .A2(new_n31799_), .B(new_n29932_), .ZN(new_n31803_));
  INV_X1     g29367(.I(new_n31174_), .ZN(new_n31804_));
  NOR2_X1    g29368(.A1(new_n31137_), .A2(po1038), .ZN(new_n31805_));
  AOI21_X1   g29369(.A1(new_n31805_), .A2(new_n31146_), .B(new_n31804_), .ZN(new_n31806_));
  NOR2_X1    g29370(.A1(new_n31806_), .A2(new_n29035_), .ZN(new_n31807_));
  NOR2_X1    g29371(.A1(new_n31111_), .A2(po1038), .ZN(new_n31808_));
  OAI21_X1   g29372(.A1(new_n8807_), .A2(new_n31113_), .B(new_n31808_), .ZN(new_n31809_));
  NAND2_X1   g29373(.A1(new_n31256_), .A2(new_n31173_), .ZN(new_n31810_));
  NAND2_X1   g29374(.A1(new_n31809_), .A2(new_n31810_), .ZN(new_n31811_));
  INV_X1     g29375(.I(new_n31811_), .ZN(new_n31812_));
  NOR2_X1    g29376(.A1(new_n31812_), .A2(new_n30020_), .ZN(new_n31813_));
  INV_X1     g29377(.I(new_n31813_), .ZN(new_n31814_));
  NOR2_X1    g29378(.A1(new_n31814_), .A2(pi1151), .ZN(new_n31815_));
  OAI21_X1   g29379(.A1(new_n31815_), .A2(new_n31807_), .B(new_n28422_), .ZN(new_n31816_));
  NOR2_X1    g29380(.A1(new_n31774_), .A2(new_n6643_), .ZN(new_n31817_));
  NOR2_X1    g29381(.A1(new_n31105_), .A2(new_n8807_), .ZN(new_n31818_));
  OAI21_X1   g29382(.A1(new_n31818_), .A2(new_n31137_), .B(new_n30137_), .ZN(new_n31819_));
  AOI22_X1   g29383(.A1(new_n31819_), .A2(new_n6643_), .B1(new_n31171_), .B2(new_n31817_), .ZN(new_n31820_));
  INV_X1     g29384(.I(new_n31817_), .ZN(new_n31821_));
  NOR2_X1    g29385(.A1(new_n31821_), .A2(new_n31092_), .ZN(new_n31822_));
  NOR2_X1    g29386(.A1(new_n31098_), .A2(pi0219), .ZN(new_n31823_));
  NOR3_X1    g29387(.A1(new_n31818_), .A2(po1038), .A3(new_n31823_), .ZN(new_n31824_));
  OAI21_X1   g29388(.A1(new_n31824_), .A2(new_n31822_), .B(new_n29035_), .ZN(new_n31825_));
  OAI21_X1   g29389(.A1(new_n31820_), .A2(new_n29035_), .B(new_n31825_), .ZN(new_n31826_));
  AOI21_X1   g29390(.A1(new_n31826_), .A2(pi1152), .B(new_n29927_), .ZN(new_n31827_));
  AOI21_X1   g29391(.A1(new_n31816_), .A2(new_n31827_), .B(pi1150), .ZN(new_n31828_));
  NOR2_X1    g29392(.A1(new_n31089_), .A2(new_n6643_), .ZN(new_n31829_));
  INV_X1     g29393(.I(new_n31829_), .ZN(new_n31830_));
  NOR2_X1    g29394(.A1(new_n31123_), .A2(new_n31830_), .ZN(new_n31831_));
  NAND2_X1   g29395(.A1(new_n31133_), .A2(new_n30140_), .ZN(new_n31832_));
  NAND2_X1   g29396(.A1(new_n31116_), .A2(pi0219), .ZN(new_n31833_));
  OAI21_X1   g29397(.A1(new_n31833_), .A2(new_n30063_), .B(new_n31832_), .ZN(new_n31834_));
  AOI21_X1   g29398(.A1(new_n31834_), .A2(new_n6643_), .B(new_n31831_), .ZN(new_n31835_));
  NAND2_X1   g29399(.A1(new_n31835_), .A2(pi1151), .ZN(new_n31836_));
  OAI21_X1   g29400(.A1(pi0219), .A2(new_n30133_), .B(new_n31833_), .ZN(new_n31837_));
  NAND2_X1   g29401(.A1(new_n31837_), .A2(new_n6643_), .ZN(new_n31838_));
  AOI21_X1   g29402(.A1(new_n8807_), .A2(new_n30120_), .B(new_n31838_), .ZN(new_n31839_));
  NAND2_X1   g29403(.A1(new_n31839_), .A2(new_n30071_), .ZN(new_n31840_));
  NAND2_X1   g29404(.A1(new_n31829_), .A2(new_n31085_), .ZN(new_n31841_));
  NAND2_X1   g29405(.A1(new_n31840_), .A2(new_n31841_), .ZN(new_n31842_));
  INV_X1     g29406(.I(new_n31842_), .ZN(new_n31843_));
  NAND2_X1   g29407(.A1(new_n31843_), .A2(new_n29035_), .ZN(new_n31844_));
  AOI21_X1   g29408(.A1(new_n31844_), .A2(new_n31836_), .B(new_n28422_), .ZN(new_n31845_));
  NAND3_X1   g29409(.A1(new_n31087_), .A2(pi0219), .A3(po1038), .ZN(new_n31846_));
  OAI21_X1   g29410(.A1(new_n30054_), .A2(new_n31823_), .B(new_n31834_), .ZN(new_n31847_));
  NAND2_X1   g29411(.A1(new_n31847_), .A2(new_n6643_), .ZN(new_n31848_));
  NAND3_X1   g29412(.A1(new_n31848_), .A2(new_n31124_), .A3(new_n31846_), .ZN(new_n31849_));
  NAND2_X1   g29413(.A1(new_n31849_), .A2(pi1151), .ZN(new_n31850_));
  NAND2_X1   g29414(.A1(new_n31808_), .A2(new_n30115_), .ZN(new_n31851_));
  NAND3_X1   g29415(.A1(new_n31851_), .A2(new_n31085_), .A3(new_n31846_), .ZN(new_n31852_));
  NAND2_X1   g29416(.A1(new_n31852_), .A2(new_n29035_), .ZN(new_n31853_));
  AOI21_X1   g29417(.A1(new_n31850_), .A2(new_n31853_), .B(pi1152), .ZN(new_n31854_));
  OAI21_X1   g29418(.A1(new_n31845_), .A2(new_n31854_), .B(new_n29927_), .ZN(new_n31855_));
  NAND2_X1   g29419(.A1(new_n31855_), .A2(new_n31828_), .ZN(new_n31856_));
  OAI21_X1   g29420(.A1(new_n31255_), .A2(new_n31821_), .B(new_n31809_), .ZN(new_n31857_));
  NOR2_X1    g29421(.A1(new_n30016_), .A2(pi1091), .ZN(new_n31858_));
  NOR2_X1    g29422(.A1(new_n31858_), .A2(po1038), .ZN(new_n31859_));
  AOI21_X1   g29423(.A1(new_n31162_), .A2(new_n31859_), .B(new_n31857_), .ZN(new_n31860_));
  INV_X1     g29424(.I(new_n31860_), .ZN(new_n31861_));
  NOR2_X1    g29425(.A1(new_n31861_), .A2(new_n29035_), .ZN(new_n31862_));
  NOR2_X1    g29426(.A1(new_n31128_), .A2(new_n30029_), .ZN(new_n31863_));
  OAI22_X1   g29427(.A1(new_n31848_), .A2(new_n31863_), .B1(new_n31122_), .B2(new_n31821_), .ZN(new_n31864_));
  NOR2_X1    g29428(.A1(new_n31864_), .A2(pi1151), .ZN(new_n31865_));
  OAI21_X1   g29429(.A1(new_n31865_), .A2(new_n31862_), .B(pi0268), .ZN(new_n31866_));
  NOR2_X1    g29430(.A1(new_n31830_), .A2(new_n31169_), .ZN(new_n31867_));
  INV_X1     g29431(.I(new_n31867_), .ZN(new_n31868_));
  NOR2_X1    g29432(.A1(new_n31822_), .A2(new_n31868_), .ZN(new_n31869_));
  NOR2_X1    g29433(.A1(new_n31831_), .A2(new_n31869_), .ZN(new_n31870_));
  NAND2_X1   g29434(.A1(new_n31838_), .A2(new_n31870_), .ZN(new_n31871_));
  OAI21_X1   g29435(.A1(new_n30029_), .A2(new_n2628_), .B(pi0219), .ZN(new_n31872_));
  AOI21_X1   g29436(.A1(new_n31148_), .A2(new_n31872_), .B(new_n30058_), .ZN(new_n31873_));
  OAI21_X1   g29437(.A1(new_n31873_), .A2(new_n31282_), .B(new_n6643_), .ZN(new_n31874_));
  NAND2_X1   g29438(.A1(new_n31874_), .A2(new_n31868_), .ZN(new_n31875_));
  INV_X1     g29439(.I(new_n31875_), .ZN(new_n31876_));
  NAND2_X1   g29440(.A1(new_n31876_), .A2(new_n29035_), .ZN(new_n31877_));
  OAI21_X1   g29441(.A1(new_n29035_), .A2(new_n31871_), .B(new_n31877_), .ZN(new_n31878_));
  AOI21_X1   g29442(.A1(new_n31878_), .A2(new_n29927_), .B(new_n28422_), .ZN(new_n31879_));
  INV_X1     g29443(.I(new_n31869_), .ZN(new_n31880_));
  NAND3_X1   g29444(.A1(new_n31873_), .A2(new_n6643_), .A3(new_n31500_), .ZN(new_n31881_));
  NAND2_X1   g29445(.A1(new_n31881_), .A2(new_n31880_), .ZN(new_n31882_));
  INV_X1     g29446(.I(new_n31852_), .ZN(new_n31883_));
  AOI21_X1   g29447(.A1(new_n30020_), .A2(new_n31811_), .B(new_n31883_), .ZN(new_n31884_));
  NOR2_X1    g29448(.A1(new_n31884_), .A2(new_n29035_), .ZN(new_n31885_));
  AOI21_X1   g29449(.A1(new_n29035_), .A2(new_n31882_), .B(new_n31885_), .ZN(new_n31886_));
  INV_X1     g29450(.I(new_n31122_), .ZN(new_n31887_));
  NOR2_X1    g29451(.A1(new_n31834_), .A2(po1038), .ZN(new_n31888_));
  AOI22_X1   g29452(.A1(new_n31888_), .A2(new_n31162_), .B1(new_n31887_), .B2(new_n31173_), .ZN(new_n31889_));
  NAND2_X1   g29453(.A1(new_n31889_), .A2(new_n29035_), .ZN(new_n31890_));
  NAND2_X1   g29454(.A1(new_n31890_), .A2(pi0268), .ZN(new_n31891_));
  NOR2_X1    g29455(.A1(new_n31811_), .A2(new_n29035_), .ZN(new_n31892_));
  OAI22_X1   g29456(.A1(new_n31891_), .A2(new_n31892_), .B1(pi0268), .B2(new_n31886_), .ZN(new_n31893_));
  AOI22_X1   g29457(.A1(new_n31879_), .A2(new_n31866_), .B1(new_n28422_), .B2(new_n31893_), .ZN(new_n31894_));
  OAI21_X1   g29458(.A1(new_n31894_), .A2(new_n29650_), .B(new_n31856_), .ZN(new_n31895_));
  AOI21_X1   g29459(.A1(new_n31895_), .A2(new_n29931_), .B(pi0230), .ZN(new_n31896_));
  AOI22_X1   g29460(.A1(new_n31896_), .A2(new_n31803_), .B1(pi0230), .B2(new_n31797_), .ZN(po0425));
  NOR2_X1    g29461(.A1(pi0211), .A2(pi1136), .ZN(new_n31898_));
  AOI21_X1   g29462(.A1(pi0211), .A2(new_n4565_), .B(new_n31898_), .ZN(new_n31899_));
  AOI22_X1   g29463(.A1(new_n31899_), .A2(new_n8807_), .B1(pi1138), .B2(new_n8808_), .ZN(new_n31900_));
  NOR2_X1    g29464(.A1(new_n12618_), .A2(new_n31900_), .ZN(new_n31901_));
  NOR2_X1    g29465(.A1(new_n4565_), .A2(pi0199), .ZN(new_n31902_));
  NOR2_X1    g29466(.A1(new_n31902_), .A2(new_n8531_), .ZN(new_n31903_));
  NOR2_X1    g29467(.A1(new_n4724_), .A2(pi0199), .ZN(new_n31904_));
  NOR2_X1    g29468(.A1(new_n8525_), .A2(new_n4408_), .ZN(new_n31905_));
  NOR3_X1    g29469(.A1(new_n31905_), .A2(new_n31904_), .A3(pi0200), .ZN(new_n31906_));
  NOR3_X1    g29470(.A1(new_n25319_), .A2(new_n31903_), .A3(new_n31906_), .ZN(new_n31907_));
  OAI21_X1   g29471(.A1(new_n31907_), .A2(new_n31901_), .B(pi0230), .ZN(new_n31908_));
  NOR2_X1    g29472(.A1(new_n3022_), .A2(pi0200), .ZN(new_n31909_));
  INV_X1     g29473(.I(new_n31909_), .ZN(new_n31910_));
  NOR2_X1    g29474(.A1(new_n31910_), .A2(new_n4408_), .ZN(new_n31911_));
  NOR3_X1    g29475(.A1(new_n25319_), .A2(new_n8525_), .A3(new_n31911_), .ZN(new_n31912_));
  NOR2_X1    g29476(.A1(new_n12618_), .A2(new_n8807_), .ZN(new_n31913_));
  INV_X1     g29477(.I(new_n31913_), .ZN(new_n31914_));
  AOI21_X1   g29478(.A1(pi1138), .A2(new_n31032_), .B(new_n31914_), .ZN(new_n31915_));
  NOR2_X1    g29479(.A1(new_n30014_), .A2(pi0269), .ZN(new_n31916_));
  AOI21_X1   g29480(.A1(pi0817), .A2(new_n30014_), .B(new_n31916_), .ZN(new_n31917_));
  OAI22_X1   g29481(.A1(new_n31915_), .A2(new_n31912_), .B1(pi1091), .B2(new_n31917_), .ZN(new_n31918_));
  AOI21_X1   g29482(.A1(pi1091), .A2(new_n31899_), .B(new_n29460_), .ZN(new_n31919_));
  INV_X1     g29483(.I(new_n31784_), .ZN(new_n31920_));
  NAND2_X1   g29484(.A1(new_n8531_), .A2(pi1136), .ZN(new_n31921_));
  NAND2_X1   g29485(.A1(pi0200), .A2(pi1137), .ZN(new_n31922_));
  AOI21_X1   g29486(.A1(new_n31921_), .A2(new_n31922_), .B(new_n3022_), .ZN(new_n31923_));
  NOR2_X1    g29487(.A1(new_n31920_), .A2(new_n31923_), .ZN(new_n31924_));
  NOR2_X1    g29488(.A1(new_n30003_), .A2(pi0269), .ZN(new_n31925_));
  AOI21_X1   g29489(.A1(pi0817), .A2(new_n30003_), .B(new_n31925_), .ZN(new_n31926_));
  OAI22_X1   g29490(.A1(new_n31924_), .A2(new_n31919_), .B1(pi1091), .B2(new_n31926_), .ZN(new_n31927_));
  NAND3_X1   g29491(.A1(new_n31927_), .A2(new_n31918_), .A3(new_n27999_), .ZN(new_n31928_));
  NAND2_X1   g29492(.A1(new_n31928_), .A2(new_n31908_), .ZN(po0426));
  AOI21_X1   g29493(.A1(new_n8525_), .A2(pi1140), .B(new_n8531_), .ZN(new_n31930_));
  OAI21_X1   g29494(.A1(pi0199), .A2(new_n4238_), .B(new_n8531_), .ZN(new_n31931_));
  AOI21_X1   g29495(.A1(pi0199), .A2(pi1141), .B(new_n31931_), .ZN(new_n31932_));
  NOR2_X1    g29496(.A1(new_n31932_), .A2(new_n31930_), .ZN(new_n31933_));
  NOR2_X1    g29497(.A1(pi0211), .A2(pi1139), .ZN(new_n31934_));
  AOI21_X1   g29498(.A1(pi0211), .A2(new_n4083_), .B(new_n31934_), .ZN(new_n31935_));
  AOI22_X1   g29499(.A1(new_n31935_), .A2(new_n8807_), .B1(pi1141), .B2(new_n8808_), .ZN(new_n31936_));
  NOR2_X1    g29500(.A1(new_n12618_), .A2(new_n31936_), .ZN(new_n31937_));
  AOI21_X1   g29501(.A1(new_n12618_), .A2(new_n31933_), .B(new_n31937_), .ZN(new_n31938_));
  INV_X1     g29502(.I(pi0270), .ZN(new_n31939_));
  NAND2_X1   g29503(.A1(new_n30004_), .A2(new_n31939_), .ZN(new_n31940_));
  NAND2_X1   g29504(.A1(new_n30003_), .A2(pi0805), .ZN(new_n31941_));
  AOI21_X1   g29505(.A1(new_n31940_), .A2(new_n31941_), .B(pi1091), .ZN(new_n31942_));
  NAND2_X1   g29506(.A1(new_n31935_), .A2(pi1091), .ZN(new_n31943_));
  NOR2_X1    g29507(.A1(new_n8531_), .A2(new_n4083_), .ZN(new_n31944_));
  NOR2_X1    g29508(.A1(new_n4238_), .A2(pi0200), .ZN(new_n31945_));
  OAI21_X1   g29509(.A1(new_n31944_), .A2(new_n31945_), .B(pi1091), .ZN(new_n31946_));
  AOI22_X1   g29510(.A1(new_n31784_), .A2(new_n31946_), .B1(new_n29459_), .B2(new_n31943_), .ZN(new_n31947_));
  NOR2_X1    g29511(.A1(new_n31947_), .A2(new_n31942_), .ZN(new_n31948_));
  NAND2_X1   g29512(.A1(new_n30015_), .A2(new_n31939_), .ZN(new_n31949_));
  NAND2_X1   g29513(.A1(new_n30014_), .A2(pi0805), .ZN(new_n31950_));
  AOI21_X1   g29514(.A1(new_n31949_), .A2(new_n31950_), .B(pi1091), .ZN(new_n31951_));
  NAND2_X1   g29515(.A1(new_n31558_), .A2(new_n8510_), .ZN(new_n31952_));
  AOI21_X1   g29516(.A1(new_n31558_), .A2(new_n8531_), .B(new_n8525_), .ZN(new_n31953_));
  AOI22_X1   g29517(.A1(new_n31913_), .A2(new_n31952_), .B1(new_n12618_), .B2(new_n31953_), .ZN(new_n31954_));
  OAI21_X1   g29518(.A1(new_n31954_), .A2(new_n31951_), .B(new_n27999_), .ZN(new_n31955_));
  OAI22_X1   g29519(.A1(new_n31948_), .A2(new_n31955_), .B1(new_n27999_), .B2(new_n31938_), .ZN(po0427));
  AOI21_X1   g29520(.A1(new_n8510_), .A2(pi1147), .B(new_n8807_), .ZN(new_n31957_));
  NOR3_X1    g29521(.A1(new_n29417_), .A2(new_n29415_), .A3(pi0219), .ZN(new_n31958_));
  OAI21_X1   g29522(.A1(new_n31957_), .A2(new_n31958_), .B(po1038), .ZN(new_n31959_));
  OAI21_X1   g29523(.A1(new_n29396_), .A2(new_n29567_), .B(new_n8807_), .ZN(new_n31960_));
  NAND2_X1   g29524(.A1(new_n29309_), .A2(new_n28796_), .ZN(new_n31961_));
  NAND4_X1   g29525(.A1(new_n28321_), .A2(pi1147), .A3(new_n28045_), .A4(new_n29472_), .ZN(new_n31962_));
  NAND4_X1   g29526(.A1(new_n31960_), .A2(new_n6643_), .A3(new_n31962_), .A4(new_n31961_), .ZN(new_n31963_));
  AOI21_X1   g29527(.A1(new_n31963_), .A2(new_n31959_), .B(new_n27999_), .ZN(new_n31964_));
  XOR2_X1    g29528(.A1(new_n30006_), .A2(new_n30000_), .Z(new_n31965_));
  NOR2_X1    g29529(.A1(new_n3022_), .A2(new_n3343_), .ZN(new_n31966_));
  AOI21_X1   g29530(.A1(new_n31965_), .A2(new_n3022_), .B(new_n31966_), .ZN(new_n31967_));
  NOR2_X1    g29531(.A1(new_n31033_), .A2(new_n3343_), .ZN(new_n31968_));
  NOR2_X1    g29532(.A1(new_n31967_), .A2(new_n31968_), .ZN(new_n31969_));
  NAND2_X1   g29533(.A1(new_n31032_), .A2(pi1145), .ZN(new_n31970_));
  NAND2_X1   g29534(.A1(new_n31970_), .A2(new_n8807_), .ZN(new_n31971_));
  NOR2_X1    g29535(.A1(new_n30016_), .A2(pi0271), .ZN(new_n31972_));
  NOR3_X1    g29536(.A1(new_n30018_), .A2(pi1091), .A3(new_n31972_), .ZN(new_n31973_));
  OAI22_X1   g29537(.A1(new_n31969_), .A2(new_n31971_), .B1(new_n8807_), .B2(new_n31973_), .ZN(new_n31974_));
  NOR2_X1    g29538(.A1(new_n28044_), .A2(new_n3022_), .ZN(new_n31975_));
  AOI21_X1   g29539(.A1(pi1147), .A2(new_n31975_), .B(new_n12618_), .ZN(new_n31976_));
  NAND2_X1   g29540(.A1(new_n31974_), .A2(new_n31976_), .ZN(new_n31977_));
  OR2_X2     g29541(.A1(new_n31973_), .A2(new_n8525_), .Z(new_n31978_));
  NAND2_X1   g29542(.A1(new_n31967_), .A2(new_n8525_), .ZN(new_n31979_));
  AOI21_X1   g29543(.A1(new_n31979_), .A2(new_n31978_), .B(new_n8531_), .ZN(new_n31980_));
  NAND2_X1   g29544(.A1(new_n31965_), .A2(new_n3022_), .ZN(new_n31981_));
  NOR2_X1    g29545(.A1(new_n3022_), .A2(new_n3512_), .ZN(new_n31982_));
  NOR2_X1    g29546(.A1(new_n31982_), .A2(pi0199), .ZN(new_n31983_));
  NAND2_X1   g29547(.A1(new_n31981_), .A2(new_n31983_), .ZN(new_n31984_));
  NAND2_X1   g29548(.A1(pi0199), .A2(pi1091), .ZN(new_n31985_));
  OAI21_X1   g29549(.A1(new_n31985_), .A2(new_n29363_), .B(new_n8531_), .ZN(new_n31986_));
  AOI21_X1   g29550(.A1(new_n31984_), .A2(new_n31978_), .B(new_n31986_), .ZN(new_n31987_));
  OAI21_X1   g29551(.A1(new_n31980_), .A2(new_n31987_), .B(new_n12618_), .ZN(new_n31988_));
  NAND2_X1   g29552(.A1(new_n31977_), .A2(new_n31988_), .ZN(new_n31989_));
  AOI21_X1   g29553(.A1(new_n31989_), .A2(new_n27999_), .B(new_n31964_), .ZN(po0428));
  NOR2_X1    g29554(.A1(new_n10290_), .A2(po1038), .ZN(new_n31991_));
  AOI21_X1   g29555(.A1(new_n29156_), .A2(new_n8510_), .B(new_n31991_), .ZN(new_n31992_));
  NAND2_X1   g29556(.A1(new_n31992_), .A2(new_n29650_), .ZN(new_n31993_));
  AOI21_X1   g29557(.A1(new_n31782_), .A2(new_n31993_), .B(pi1149), .ZN(new_n31994_));
  INV_X1     g29558(.I(new_n31785_), .ZN(new_n31995_));
  OAI22_X1   g29559(.A1(new_n12618_), .A2(pi0211), .B1(po1038), .B2(new_n28448_), .ZN(new_n31996_));
  OAI21_X1   g29560(.A1(new_n31996_), .A2(new_n29459_), .B(pi1150), .ZN(new_n31997_));
  NAND2_X1   g29561(.A1(new_n31997_), .A2(pi1149), .ZN(new_n31998_));
  OAI21_X1   g29562(.A1(new_n31995_), .A2(new_n31998_), .B(pi1148), .ZN(new_n31999_));
  NOR2_X1    g29563(.A1(new_n31999_), .A2(new_n31994_), .ZN(new_n32000_));
  AOI21_X1   g29564(.A1(new_n31192_), .A2(pi1150), .B(pi1149), .ZN(new_n32001_));
  OR2_X2     g29565(.A1(new_n32001_), .A2(pi1148), .Z(new_n32002_));
  NAND2_X1   g29566(.A1(new_n31789_), .A2(pi1149), .ZN(new_n32003_));
  AOI22_X1   g29567(.A1(new_n31998_), .A2(new_n32003_), .B1(new_n29650_), .B2(new_n31793_), .ZN(new_n32004_));
  OAI21_X1   g29568(.A1(new_n32002_), .A2(new_n32004_), .B(pi0230), .ZN(new_n32005_));
  NOR2_X1    g29569(.A1(new_n32005_), .A2(new_n32000_), .ZN(new_n32006_));
  NOR2_X1    g29570(.A1(new_n31790_), .A2(new_n29650_), .ZN(new_n32007_));
  NOR2_X1    g29571(.A1(new_n31793_), .A2(pi1150), .ZN(new_n32008_));
  OAI21_X1   g29572(.A1(new_n32007_), .A2(new_n32008_), .B(pi1149), .ZN(new_n32009_));
  NOR2_X1    g29573(.A1(new_n32002_), .A2(new_n3022_), .ZN(new_n32010_));
  AOI21_X1   g29574(.A1(new_n32010_), .A2(new_n32009_), .B(pi0283), .ZN(new_n32011_));
  NAND2_X1   g29575(.A1(new_n32000_), .A2(pi1091), .ZN(new_n32012_));
  AOI21_X1   g29576(.A1(new_n32011_), .A2(new_n32012_), .B(pi0272), .ZN(new_n32013_));
  NOR2_X1    g29577(.A1(new_n31835_), .A2(new_n29650_), .ZN(new_n32014_));
  INV_X1     g29578(.I(new_n32014_), .ZN(new_n32015_));
  NAND4_X1   g29579(.A1(new_n31848_), .A2(new_n29650_), .A3(new_n31124_), .A4(new_n31846_), .ZN(new_n32016_));
  AOI21_X1   g29580(.A1(new_n32016_), .A2(new_n32015_), .B(new_n29297_), .ZN(new_n32017_));
  NAND2_X1   g29581(.A1(new_n31842_), .A2(pi1150), .ZN(new_n32018_));
  NAND2_X1   g29582(.A1(new_n31883_), .A2(new_n29650_), .ZN(new_n32019_));
  AOI21_X1   g29583(.A1(new_n32018_), .A2(new_n32019_), .B(pi1149), .ZN(new_n32020_));
  NOR3_X1    g29584(.A1(new_n32020_), .A2(new_n32017_), .A3(pi1148), .ZN(new_n32021_));
  NOR2_X1    g29585(.A1(new_n31871_), .A2(new_n29650_), .ZN(new_n32022_));
  AND2_X2    g29586(.A1(new_n31884_), .A2(new_n29650_), .Z(new_n32023_));
  OAI21_X1   g29587(.A1(new_n32022_), .A2(new_n32023_), .B(pi1149), .ZN(new_n32024_));
  NOR2_X1    g29588(.A1(new_n31875_), .A2(new_n29650_), .ZN(new_n32025_));
  NOR2_X1    g29589(.A1(new_n31882_), .A2(pi1150), .ZN(new_n32026_));
  OAI21_X1   g29590(.A1(new_n32025_), .A2(new_n32026_), .B(new_n29297_), .ZN(new_n32027_));
  AOI21_X1   g29591(.A1(new_n32027_), .A2(new_n32024_), .B(new_n29296_), .ZN(new_n32028_));
  OAI21_X1   g29592(.A1(new_n32021_), .A2(new_n32028_), .B(pi0283), .ZN(new_n32029_));
  AOI21_X1   g29593(.A1(new_n32029_), .A2(new_n32013_), .B(pi0230), .ZN(new_n32030_));
  NOR2_X1    g29594(.A1(new_n31824_), .A2(new_n31822_), .ZN(new_n32031_));
  NOR2_X1    g29595(.A1(new_n31813_), .A2(pi1150), .ZN(new_n32032_));
  AOI21_X1   g29596(.A1(pi1150), .A2(new_n32031_), .B(new_n32032_), .ZN(new_n32033_));
  NAND2_X1   g29597(.A1(new_n31820_), .A2(pi1150), .ZN(new_n32034_));
  AOI21_X1   g29598(.A1(new_n31806_), .A2(new_n29650_), .B(new_n29297_), .ZN(new_n32035_));
  AOI22_X1   g29599(.A1(new_n32033_), .A2(new_n29297_), .B1(new_n32035_), .B2(new_n32034_), .ZN(new_n32036_));
  OAI21_X1   g29600(.A1(new_n32036_), .A2(pi1148), .B(pi0283), .ZN(new_n32037_));
  NOR2_X1    g29601(.A1(new_n31860_), .A2(new_n29650_), .ZN(new_n32038_));
  NOR2_X1    g29602(.A1(new_n31812_), .A2(pi1150), .ZN(new_n32039_));
  OAI21_X1   g29603(.A1(new_n32038_), .A2(new_n32039_), .B(pi1149), .ZN(new_n32040_));
  AND2_X2    g29604(.A1(new_n31864_), .A2(pi1150), .Z(new_n32041_));
  NOR2_X1    g29605(.A1(new_n31889_), .A2(pi1150), .ZN(new_n32042_));
  OAI21_X1   g29606(.A1(new_n32041_), .A2(new_n32042_), .B(new_n29297_), .ZN(new_n32043_));
  AOI21_X1   g29607(.A1(new_n32043_), .A2(new_n32040_), .B(new_n29296_), .ZN(new_n32044_));
  INV_X1     g29608(.I(new_n29959_), .ZN(new_n32045_));
  AOI22_X1   g29609(.A1(new_n25319_), .A2(new_n31205_), .B1(new_n6643_), .B2(new_n32045_), .ZN(new_n32046_));
  NOR2_X1    g29610(.A1(new_n32046_), .A2(pi1150), .ZN(new_n32047_));
  NOR3_X1    g29611(.A1(new_n31790_), .A2(new_n3022_), .A3(new_n29650_), .ZN(new_n32048_));
  OAI21_X1   g29612(.A1(new_n32048_), .A2(new_n32047_), .B(pi1149), .ZN(new_n32049_));
  NAND2_X1   g29613(.A1(new_n32001_), .A2(pi1091), .ZN(new_n32050_));
  NAND3_X1   g29614(.A1(new_n32049_), .A2(new_n29296_), .A3(new_n32050_), .ZN(new_n32051_));
  NOR2_X1    g29615(.A1(new_n29297_), .A2(pi1150), .ZN(new_n32052_));
  NOR2_X1    g29616(.A1(new_n31781_), .A2(new_n32052_), .ZN(new_n32053_));
  NOR2_X1    g29617(.A1(new_n31995_), .A2(new_n32053_), .ZN(new_n32054_));
  OAI21_X1   g29618(.A1(new_n32054_), .A2(new_n31994_), .B(pi1091), .ZN(new_n32055_));
  AOI21_X1   g29619(.A1(new_n32055_), .A2(pi1148), .B(pi0283), .ZN(new_n32056_));
  AOI21_X1   g29620(.A1(new_n32056_), .A2(new_n32051_), .B(new_n29928_), .ZN(new_n32057_));
  OAI21_X1   g29621(.A1(new_n32044_), .A2(new_n32037_), .B(new_n32057_), .ZN(new_n32058_));
  AOI21_X1   g29622(.A1(new_n32030_), .A2(new_n32058_), .B(new_n32006_), .ZN(po0429));
  NOR3_X1    g29623(.A1(new_n31992_), .A2(new_n3343_), .A3(new_n30294_), .ZN(new_n32060_));
  AOI21_X1   g29624(.A1(new_n3343_), .A2(new_n8640_), .B(new_n31920_), .ZN(new_n32061_));
  AOI21_X1   g29625(.A1(new_n8510_), .A2(new_n29317_), .B(new_n29460_), .ZN(new_n32062_));
  OAI21_X1   g29626(.A1(new_n32061_), .A2(new_n32062_), .B(pi1147), .ZN(new_n32063_));
  NAND2_X1   g29627(.A1(new_n32063_), .A2(new_n29296_), .ZN(new_n32064_));
  NAND2_X1   g29628(.A1(new_n8525_), .A2(pi1147), .ZN(new_n32065_));
  AOI22_X1   g29629(.A1(new_n32065_), .A2(pi0200), .B1(new_n3343_), .B2(new_n8640_), .ZN(new_n32066_));
  AOI21_X1   g29630(.A1(new_n12618_), .A2(new_n32066_), .B(new_n29296_), .ZN(new_n32067_));
  NOR2_X1    g29631(.A1(new_n29460_), .A2(new_n29363_), .ZN(new_n32068_));
  OAI22_X1   g29632(.A1(new_n32068_), .A2(new_n31780_), .B1(pi1146), .B2(new_n31605_), .ZN(new_n32069_));
  AOI21_X1   g29633(.A1(new_n32069_), .A2(new_n32067_), .B(new_n27999_), .ZN(new_n32070_));
  OAI21_X1   g29634(.A1(new_n32064_), .A2(new_n32060_), .B(new_n32070_), .ZN(new_n32071_));
  XOR2_X1    g29635(.A1(new_n30018_), .A2(pi0273), .Z(new_n32072_));
  NAND2_X1   g29636(.A1(new_n32072_), .A2(new_n3022_), .ZN(new_n32073_));
  AOI21_X1   g29637(.A1(new_n32073_), .A2(pi0199), .B(pi0299), .ZN(new_n32074_));
  NAND2_X1   g29638(.A1(new_n31966_), .A2(new_n8531_), .ZN(new_n32075_));
  NAND2_X1   g29639(.A1(new_n30010_), .A2(new_n29999_), .ZN(new_n32076_));
  NAND3_X1   g29640(.A1(new_n30012_), .A2(new_n30019_), .A3(new_n32076_), .ZN(new_n32077_));
  NAND3_X1   g29641(.A1(new_n32077_), .A2(new_n8525_), .A3(new_n32075_), .ZN(new_n32078_));
  NAND2_X1   g29642(.A1(new_n32078_), .A2(new_n32074_), .ZN(new_n32079_));
  NOR2_X1    g29643(.A1(new_n31968_), .A2(pi0219), .ZN(new_n32080_));
  AOI22_X1   g29644(.A1(new_n32077_), .A2(new_n32080_), .B1(pi0219), .B2(new_n32073_), .ZN(new_n32081_));
  INV_X1     g29645(.I(new_n32081_), .ZN(new_n32082_));
  OAI21_X1   g29646(.A1(new_n2628_), .A2(new_n32082_), .B(new_n32079_), .ZN(new_n32083_));
  NOR2_X1    g29647(.A1(new_n31263_), .A2(new_n9220_), .ZN(new_n32084_));
  NOR2_X1    g29648(.A1(new_n32084_), .A2(new_n3022_), .ZN(new_n32085_));
  OAI21_X1   g29649(.A1(new_n32085_), .A2(new_n32083_), .B(new_n6643_), .ZN(new_n32086_));
  NAND2_X1   g29650(.A1(new_n31804_), .A2(pi1091), .ZN(new_n32087_));
  AOI21_X1   g29651(.A1(new_n32086_), .A2(new_n32087_), .B(new_n29363_), .ZN(new_n32088_));
  NOR2_X1    g29652(.A1(new_n32082_), .A2(new_n6643_), .ZN(new_n32089_));
  NAND2_X1   g29653(.A1(new_n31190_), .A2(pi1091), .ZN(new_n32090_));
  OAI21_X1   g29654(.A1(new_n32081_), .A2(new_n31975_), .B(pi0299), .ZN(new_n32091_));
  OR2_X2     g29655(.A1(new_n31980_), .A2(new_n29949_), .Z(new_n32092_));
  NAND3_X1   g29656(.A1(new_n32091_), .A2(new_n32079_), .A3(new_n32092_), .ZN(new_n32093_));
  AOI21_X1   g29657(.A1(new_n32093_), .A2(new_n6643_), .B(new_n29296_), .ZN(new_n32094_));
  NAND2_X1   g29658(.A1(new_n32083_), .A2(new_n29359_), .ZN(new_n32095_));
  AOI22_X1   g29659(.A1(new_n32094_), .A2(new_n32090_), .B1(new_n29296_), .B2(new_n32095_), .ZN(new_n32096_));
  NOR3_X1    g29660(.A1(new_n32088_), .A2(new_n32089_), .A3(new_n32096_), .ZN(new_n32097_));
  OAI21_X1   g29661(.A1(new_n32097_), .A2(pi0230), .B(new_n32071_), .ZN(po0430));
  NOR2_X1    g29662(.A1(new_n29308_), .A2(new_n28032_), .ZN(new_n32099_));
  NOR2_X1    g29663(.A1(new_n28783_), .A2(new_n28079_), .ZN(new_n32100_));
  NOR2_X1    g29664(.A1(new_n32100_), .A2(pi0219), .ZN(new_n32101_));
  NOR2_X1    g29665(.A1(new_n29567_), .A2(new_n10289_), .ZN(new_n32102_));
  OAI22_X1   g29666(.A1(new_n32102_), .A2(new_n32101_), .B1(new_n29858_), .B2(new_n32099_), .ZN(new_n32103_));
  OAI21_X1   g29667(.A1(new_n29416_), .A2(new_n32101_), .B(pi0230), .ZN(new_n32104_));
  AOI21_X1   g29668(.A1(new_n6643_), .A2(new_n32103_), .B(new_n32104_), .ZN(new_n32105_));
  INV_X1     g29669(.I(pi0274), .ZN(new_n32106_));
  NAND2_X1   g29670(.A1(new_n30004_), .A2(new_n32106_), .ZN(new_n32107_));
  NAND2_X1   g29671(.A1(new_n30003_), .A2(pi0659), .ZN(new_n32108_));
  AOI21_X1   g29672(.A1(new_n32107_), .A2(new_n32108_), .B(pi1091), .ZN(new_n32109_));
  NOR3_X1    g29673(.A1(new_n32109_), .A2(new_n8510_), .A3(new_n31600_), .ZN(new_n32110_));
  NOR3_X1    g29674(.A1(new_n32109_), .A2(pi0211), .A3(new_n31572_), .ZN(new_n32111_));
  OAI21_X1   g29675(.A1(new_n32110_), .A2(new_n32111_), .B(new_n8807_), .ZN(new_n32112_));
  NOR2_X1    g29676(.A1(new_n30014_), .A2(pi0274), .ZN(new_n32113_));
  AND2_X2    g29677(.A1(new_n30014_), .A2(pi0659), .Z(new_n32114_));
  OAI21_X1   g29678(.A1(new_n32114_), .A2(new_n32113_), .B(new_n3022_), .ZN(new_n32115_));
  NAND3_X1   g29679(.A1(new_n32115_), .A2(pi0219), .A3(new_n31970_), .ZN(new_n32116_));
  NAND3_X1   g29680(.A1(new_n32112_), .A2(new_n25319_), .A3(new_n32116_), .ZN(new_n32117_));
  NOR3_X1    g29681(.A1(new_n32109_), .A2(new_n8531_), .A3(new_n31600_), .ZN(new_n32118_));
  NOR3_X1    g29682(.A1(new_n32109_), .A2(pi0200), .A3(new_n31572_), .ZN(new_n32119_));
  OAI21_X1   g29683(.A1(new_n32118_), .A2(new_n32119_), .B(new_n8525_), .ZN(new_n32120_));
  AOI21_X1   g29684(.A1(new_n31982_), .A2(new_n8531_), .B(new_n8525_), .ZN(new_n32121_));
  AOI21_X1   g29685(.A1(new_n32115_), .A2(new_n32121_), .B(new_n25319_), .ZN(new_n32122_));
  AOI21_X1   g29686(.A1(new_n32120_), .A2(new_n32122_), .B(pi0230), .ZN(new_n32123_));
  AOI21_X1   g29687(.A1(new_n32123_), .A2(new_n32117_), .B(new_n32105_), .ZN(po0431));
  NOR2_X1    g29688(.A1(new_n31781_), .A2(new_n29035_), .ZN(new_n32125_));
  NOR3_X1    g29689(.A1(new_n31995_), .A2(new_n32125_), .A3(new_n29297_), .ZN(new_n32126_));
  AOI21_X1   g29690(.A1(new_n31781_), .A2(new_n32052_), .B(new_n32126_), .ZN(new_n32127_));
  AOI21_X1   g29691(.A1(new_n31192_), .A2(new_n29640_), .B(pi1149), .ZN(new_n32128_));
  NOR2_X1    g29692(.A1(new_n31790_), .A2(new_n29035_), .ZN(new_n32129_));
  NOR2_X1    g29693(.A1(new_n31793_), .A2(pi1151), .ZN(new_n32130_));
  OR3_X2     g29694(.A1(new_n32129_), .A2(new_n29650_), .A3(new_n32130_), .Z(new_n32131_));
  NAND2_X1   g29695(.A1(new_n32131_), .A2(new_n32128_), .ZN(new_n32132_));
  NAND2_X1   g29696(.A1(new_n32132_), .A2(new_n32127_), .ZN(new_n32133_));
  AOI21_X1   g29697(.A1(new_n31992_), .A2(new_n29035_), .B(new_n29297_), .ZN(new_n32134_));
  NAND2_X1   g29698(.A1(new_n31782_), .A2(new_n32134_), .ZN(new_n32135_));
  NOR2_X1    g29699(.A1(new_n29035_), .A2(pi1149), .ZN(new_n32136_));
  AOI21_X1   g29700(.A1(new_n31192_), .A2(new_n32136_), .B(pi1150), .ZN(new_n32137_));
  NAND2_X1   g29701(.A1(new_n32135_), .A2(new_n32137_), .ZN(new_n32138_));
  NOR3_X1    g29702(.A1(new_n31790_), .A2(pi1149), .A3(new_n29035_), .ZN(new_n32139_));
  OAI21_X1   g29703(.A1(new_n32126_), .A2(new_n32139_), .B(pi1150), .ZN(new_n32140_));
  AOI21_X1   g29704(.A1(new_n32140_), .A2(new_n32138_), .B(new_n3022_), .ZN(new_n32141_));
  NOR4_X1    g29705(.A1(new_n32046_), .A2(pi1149), .A3(new_n29650_), .A4(pi1151), .ZN(new_n32142_));
  OAI21_X1   g29706(.A1(new_n32141_), .A2(new_n32142_), .B(pi0275), .ZN(new_n32143_));
  NAND3_X1   g29707(.A1(new_n32132_), .A2(pi1091), .A3(new_n32127_), .ZN(new_n32144_));
  AOI22_X1   g29708(.A1(new_n32144_), .A2(new_n29929_), .B1(pi0272), .B2(pi0283), .ZN(new_n32145_));
  NAND2_X1   g29709(.A1(new_n32145_), .A2(new_n32143_), .ZN(new_n32146_));
  AOI21_X1   g29710(.A1(pi1150), .A2(new_n31884_), .B(new_n32026_), .ZN(new_n32147_));
  NOR2_X1    g29711(.A1(new_n32147_), .A2(pi1151), .ZN(new_n32148_));
  AOI21_X1   g29712(.A1(new_n31876_), .A2(new_n29650_), .B(new_n32022_), .ZN(new_n32149_));
  OAI21_X1   g29713(.A1(new_n32149_), .A2(new_n29035_), .B(new_n29929_), .ZN(new_n32150_));
  OAI21_X1   g29714(.A1(new_n32150_), .A2(new_n32148_), .B(pi1149), .ZN(new_n32151_));
  OAI21_X1   g29715(.A1(new_n31864_), .A2(new_n29035_), .B(new_n31890_), .ZN(new_n32152_));
  NOR2_X1    g29716(.A1(new_n31811_), .A2(pi1151), .ZN(new_n32153_));
  OAI21_X1   g29717(.A1(new_n31862_), .A2(new_n32153_), .B(pi1150), .ZN(new_n32154_));
  NAND2_X1   g29718(.A1(new_n32154_), .A2(pi0275), .ZN(new_n32155_));
  AOI21_X1   g29719(.A1(new_n32152_), .A2(new_n29650_), .B(new_n32155_), .ZN(new_n32156_));
  AOI21_X1   g29720(.A1(pi1150), .A2(new_n31806_), .B(new_n32032_), .ZN(new_n32157_));
  NOR2_X1    g29721(.A1(new_n32157_), .A2(pi1151), .ZN(new_n32158_));
  INV_X1     g29722(.I(new_n32034_), .ZN(new_n32159_));
  AOI21_X1   g29723(.A1(new_n29650_), .A2(new_n32031_), .B(new_n32159_), .ZN(new_n32160_));
  OAI21_X1   g29724(.A1(new_n32160_), .A2(new_n29035_), .B(pi0275), .ZN(new_n32161_));
  OAI21_X1   g29725(.A1(new_n32161_), .A2(new_n32158_), .B(new_n29297_), .ZN(new_n32162_));
  OAI21_X1   g29726(.A1(new_n31843_), .A2(pi1150), .B(new_n32015_), .ZN(new_n32163_));
  NAND2_X1   g29727(.A1(new_n32163_), .A2(pi1151), .ZN(new_n32164_));
  OAI21_X1   g29728(.A1(new_n31849_), .A2(new_n29650_), .B(new_n32019_), .ZN(new_n32165_));
  NAND2_X1   g29729(.A1(new_n32165_), .A2(new_n29035_), .ZN(new_n32166_));
  AOI21_X1   g29730(.A1(new_n32164_), .A2(new_n32166_), .B(pi0275), .ZN(new_n32167_));
  OAI22_X1   g29731(.A1(new_n32167_), .A2(new_n32162_), .B1(new_n32151_), .B2(new_n32156_), .ZN(new_n32168_));
  NOR3_X1    g29732(.A1(new_n32168_), .A2(new_n29928_), .A3(new_n29930_), .ZN(new_n32169_));
  NOR2_X1    g29733(.A1(new_n32169_), .A2(pi0230), .ZN(new_n32170_));
  AOI22_X1   g29734(.A1(new_n32170_), .A2(new_n32146_), .B1(pi0230), .B2(new_n32133_), .ZN(po0432));
  NOR2_X1    g29735(.A1(new_n29402_), .A2(new_n28062_), .ZN(new_n32172_));
  AOI22_X1   g29736(.A1(new_n32172_), .A2(new_n8807_), .B1(pi1146), .B2(new_n8808_), .ZN(new_n32173_));
  NOR2_X1    g29737(.A1(new_n12618_), .A2(new_n32173_), .ZN(new_n32174_));
  AOI21_X1   g29738(.A1(pi0199), .A2(new_n3343_), .B(new_n28790_), .ZN(new_n32175_));
  NOR2_X1    g29739(.A1(new_n32175_), .A2(pi0200), .ZN(new_n32176_));
  NOR2_X1    g29740(.A1(new_n32176_), .A2(new_n29300_), .ZN(new_n32177_));
  AOI21_X1   g29741(.A1(new_n12618_), .A2(new_n32177_), .B(new_n32174_), .ZN(new_n32178_));
  NAND2_X1   g29742(.A1(new_n32172_), .A2(pi1091), .ZN(new_n32179_));
  NOR2_X1    g29743(.A1(new_n8531_), .A2(new_n3512_), .ZN(new_n32180_));
  NOR2_X1    g29744(.A1(new_n2446_), .A2(pi0200), .ZN(new_n32181_));
  OAI21_X1   g29745(.A1(new_n32180_), .A2(new_n32181_), .B(pi1091), .ZN(new_n32182_));
  AOI22_X1   g29746(.A1(new_n31784_), .A2(new_n32182_), .B1(new_n29459_), .B2(new_n32179_), .ZN(new_n32183_));
  INV_X1     g29747(.I(new_n30006_), .ZN(new_n32184_));
  NOR2_X1    g29748(.A1(new_n30005_), .A2(pi0276), .ZN(new_n32185_));
  NOR3_X1    g29749(.A1(new_n32184_), .A2(pi1091), .A3(new_n32185_), .ZN(new_n32186_));
  OAI21_X1   g29750(.A1(new_n32183_), .A2(new_n32186_), .B(new_n27999_), .ZN(new_n32187_));
  NAND3_X1   g29751(.A1(new_n12618_), .A2(pi0199), .A3(new_n32075_), .ZN(new_n32188_));
  OAI21_X1   g29752(.A1(new_n3343_), .A2(new_n31033_), .B(new_n31913_), .ZN(new_n32189_));
  OAI21_X1   g29753(.A1(new_n30015_), .A2(new_n30001_), .B(new_n3293_), .ZN(new_n32190_));
  AOI22_X1   g29754(.A1(new_n32189_), .A2(new_n32188_), .B1(new_n31858_), .B2(new_n32190_), .ZN(new_n32191_));
  OAI22_X1   g29755(.A1(new_n32187_), .A2(new_n32191_), .B1(new_n27999_), .B2(new_n32178_), .ZN(po0433));
  NOR2_X1    g29756(.A1(new_n31545_), .A2(new_n8531_), .ZN(new_n32193_));
  AOI21_X1   g29757(.A1(new_n8525_), .A2(pi1140), .B(new_n28031_), .ZN(new_n32194_));
  NOR3_X1    g29758(.A1(new_n25319_), .A2(new_n32193_), .A3(new_n32194_), .ZN(new_n32195_));
  NAND2_X1   g29759(.A1(new_n3926_), .A2(pi0211), .ZN(new_n32196_));
  NAND2_X1   g29760(.A1(new_n8510_), .A2(new_n4083_), .ZN(new_n32197_));
  AOI21_X1   g29761(.A1(new_n32197_), .A2(new_n32196_), .B(pi0219), .ZN(new_n32198_));
  AOI21_X1   g29762(.A1(new_n8510_), .A2(pi1142), .B(new_n8807_), .ZN(new_n32199_));
  NOR3_X1    g29763(.A1(new_n12618_), .A2(new_n32198_), .A3(new_n32199_), .ZN(new_n32200_));
  OAI21_X1   g29764(.A1(new_n32195_), .A2(new_n32200_), .B(pi0230), .ZN(new_n32201_));
  NOR2_X1    g29765(.A1(new_n30003_), .A2(pi0277), .ZN(new_n32202_));
  AND2_X2    g29766(.A1(new_n30003_), .A2(pi0820), .Z(new_n32203_));
  OAI21_X1   g29767(.A1(new_n32203_), .A2(new_n32202_), .B(new_n3022_), .ZN(new_n32204_));
  NAND3_X1   g29768(.A1(new_n32204_), .A2(pi0211), .A3(new_n31559_), .ZN(new_n32205_));
  NOR2_X1    g29769(.A1(new_n3022_), .A2(new_n4083_), .ZN(new_n32206_));
  INV_X1     g29770(.I(new_n32206_), .ZN(new_n32207_));
  NAND3_X1   g29771(.A1(new_n32204_), .A2(new_n8510_), .A3(new_n32207_), .ZN(new_n32208_));
  AOI21_X1   g29772(.A1(new_n32205_), .A2(new_n32208_), .B(pi0219), .ZN(new_n32209_));
  OAI21_X1   g29773(.A1(new_n31556_), .A2(pi0211), .B(pi0219), .ZN(new_n32210_));
  INV_X1     g29774(.I(pi0277), .ZN(new_n32211_));
  NAND2_X1   g29775(.A1(new_n30015_), .A2(new_n32211_), .ZN(new_n32212_));
  NAND2_X1   g29776(.A1(new_n30014_), .A2(pi0820), .ZN(new_n32213_));
  AOI21_X1   g29777(.A1(new_n32212_), .A2(new_n32213_), .B(pi1091), .ZN(new_n32214_));
  NOR2_X1    g29778(.A1(new_n32214_), .A2(new_n32210_), .ZN(new_n32215_));
  NOR3_X1    g29779(.A1(new_n32209_), .A2(new_n12618_), .A3(new_n32215_), .ZN(new_n32216_));
  NAND3_X1   g29780(.A1(new_n32204_), .A2(pi0200), .A3(new_n31559_), .ZN(new_n32217_));
  NAND3_X1   g29781(.A1(new_n32204_), .A2(new_n8531_), .A3(new_n32207_), .ZN(new_n32218_));
  NAND2_X1   g29782(.A1(new_n32217_), .A2(new_n32218_), .ZN(new_n32219_));
  OAI21_X1   g29783(.A1(new_n31556_), .A2(pi0200), .B(pi0199), .ZN(new_n32220_));
  OAI21_X1   g29784(.A1(new_n32214_), .A2(new_n32220_), .B(new_n12618_), .ZN(new_n32221_));
  AOI21_X1   g29785(.A1(new_n32219_), .A2(new_n8525_), .B(new_n32221_), .ZN(new_n32222_));
  OAI21_X1   g29786(.A1(new_n32216_), .A2(new_n32222_), .B(new_n27999_), .ZN(new_n32223_));
  NAND2_X1   g29787(.A1(new_n32223_), .A2(new_n32201_), .ZN(po0434));
  INV_X1     g29788(.I(pi1132), .ZN(new_n32225_));
  NOR2_X1    g29789(.A1(new_n32225_), .A2(pi0211), .ZN(new_n32226_));
  AOI21_X1   g29790(.A1(pi0211), .A2(pi1133), .B(new_n32226_), .ZN(new_n32227_));
  NOR2_X1    g29791(.A1(new_n32227_), .A2(new_n28045_), .ZN(new_n32228_));
  INV_X1     g29792(.I(pi1133), .ZN(new_n32229_));
  NOR2_X1    g29793(.A1(new_n32229_), .A2(pi0199), .ZN(new_n32230_));
  OAI21_X1   g29794(.A1(new_n32230_), .A2(new_n8531_), .B(new_n2628_), .ZN(new_n32231_));
  AOI21_X1   g29795(.A1(new_n8525_), .A2(pi1132), .B(pi0200), .ZN(new_n32232_));
  NOR2_X1    g29796(.A1(new_n32231_), .A2(new_n32232_), .ZN(new_n32233_));
  OAI21_X1   g29797(.A1(new_n32228_), .A2(new_n32233_), .B(new_n6643_), .ZN(new_n32234_));
  NAND2_X1   g29798(.A1(new_n32234_), .A2(pi0230), .ZN(new_n32235_));
  NOR2_X1    g29799(.A1(new_n29379_), .A2(new_n32227_), .ZN(new_n32236_));
  NAND2_X1   g29800(.A1(new_n30014_), .A2(pi0976), .ZN(new_n32237_));
  NAND2_X1   g29801(.A1(new_n30015_), .A2(pi0278), .ZN(new_n32238_));
  AOI21_X1   g29802(.A1(new_n32238_), .A2(new_n32237_), .B(pi1091), .ZN(new_n32239_));
  NOR2_X1    g29803(.A1(new_n30004_), .A2(pi0976), .ZN(new_n32240_));
  NOR2_X1    g29804(.A1(new_n30003_), .A2(pi0278), .ZN(new_n32241_));
  OAI21_X1   g29805(.A1(new_n32240_), .A2(new_n32241_), .B(new_n3022_), .ZN(new_n32242_));
  AOI21_X1   g29806(.A1(new_n32227_), .A2(pi1091), .B(pi0219), .ZN(new_n32243_));
  AOI22_X1   g29807(.A1(new_n32242_), .A2(new_n32243_), .B1(new_n32239_), .B2(pi0219), .ZN(new_n32244_));
  OAI21_X1   g29808(.A1(new_n32244_), .A2(new_n6643_), .B(new_n27999_), .ZN(new_n32245_));
  NOR2_X1    g29809(.A1(new_n32244_), .A2(new_n2628_), .ZN(new_n32246_));
  NOR2_X1    g29810(.A1(new_n3022_), .A2(pi1133), .ZN(new_n32247_));
  NOR2_X1    g29811(.A1(new_n32247_), .A2(pi0199), .ZN(new_n32248_));
  AOI22_X1   g29812(.A1(new_n32242_), .A2(new_n32248_), .B1(new_n32239_), .B2(pi0199), .ZN(new_n32249_));
  AOI21_X1   g29813(.A1(new_n32249_), .A2(pi0200), .B(pi0299), .ZN(new_n32250_));
  NAND2_X1   g29814(.A1(new_n32239_), .A2(pi0199), .ZN(new_n32251_));
  NAND2_X1   g29815(.A1(new_n32225_), .A2(pi1091), .ZN(new_n32252_));
  NAND3_X1   g29816(.A1(new_n32242_), .A2(new_n8525_), .A3(new_n32252_), .ZN(new_n32253_));
  NAND3_X1   g29817(.A1(new_n32253_), .A2(new_n8531_), .A3(new_n32251_), .ZN(new_n32254_));
  AOI21_X1   g29818(.A1(new_n32250_), .A2(new_n32254_), .B(new_n32246_), .ZN(new_n32255_));
  NOR2_X1    g29819(.A1(new_n32255_), .A2(po1038), .ZN(new_n32256_));
  OAI22_X1   g29820(.A1(new_n32256_), .A2(new_n32245_), .B1(new_n32235_), .B2(new_n32236_), .ZN(new_n32257_));
  INV_X1     g29821(.I(new_n32090_), .ZN(new_n32258_));
  NAND4_X1   g29822(.A1(new_n32253_), .A2(new_n8531_), .A3(new_n32251_), .A4(new_n31985_), .ZN(new_n32259_));
  AOI21_X1   g29823(.A1(new_n32250_), .A2(new_n32259_), .B(new_n32246_), .ZN(new_n32260_));
  NAND3_X1   g29824(.A1(new_n31032_), .A2(pi0219), .A3(pi0299), .ZN(new_n32261_));
  AOI21_X1   g29825(.A1(new_n32260_), .A2(new_n32261_), .B(po1038), .ZN(new_n32262_));
  NOR3_X1    g29826(.A1(new_n32262_), .A2(new_n32258_), .A3(new_n32245_), .ZN(new_n32263_));
  AOI21_X1   g29827(.A1(new_n32225_), .A2(new_n8640_), .B(new_n32231_), .ZN(new_n32264_));
  NOR3_X1    g29828(.A1(new_n32264_), .A2(new_n32228_), .A3(new_n31326_), .ZN(new_n32265_));
  OAI21_X1   g29829(.A1(new_n32265_), .A2(po1038), .B(pi0230), .ZN(new_n32266_));
  AOI21_X1   g29830(.A1(new_n8807_), .A2(new_n32227_), .B(new_n29387_), .ZN(new_n32267_));
  OAI21_X1   g29831(.A1(new_n32267_), .A2(new_n32266_), .B(pi1134), .ZN(new_n32268_));
  OAI22_X1   g29832(.A1(pi1134), .A2(new_n32257_), .B1(new_n32263_), .B2(new_n32268_), .ZN(po0435));
  NOR2_X1    g29833(.A1(new_n28894_), .A2(new_n4888_), .ZN(new_n32270_));
  AOI21_X1   g29834(.A1(new_n8531_), .A2(new_n32229_), .B(pi0199), .ZN(new_n32271_));
  NOR3_X1    g29835(.A1(new_n25319_), .A2(new_n32270_), .A3(new_n32271_), .ZN(new_n32272_));
  NAND2_X1   g29836(.A1(new_n8510_), .A2(pi1135), .ZN(new_n32273_));
  AOI22_X1   g29837(.A1(new_n32273_), .A2(pi0219), .B1(new_n32229_), .B2(new_n31056_), .ZN(new_n32274_));
  NOR2_X1    g29838(.A1(new_n12618_), .A2(new_n32274_), .ZN(new_n32275_));
  OAI21_X1   g29839(.A1(new_n32272_), .A2(new_n32275_), .B(pi0230), .ZN(new_n32276_));
  INV_X1     g29840(.I(pi0958), .ZN(new_n32277_));
  NAND2_X1   g29841(.A1(new_n30003_), .A2(new_n32277_), .ZN(new_n32278_));
  NAND2_X1   g29842(.A1(new_n30004_), .A2(new_n4891_), .ZN(new_n32279_));
  AOI21_X1   g29843(.A1(new_n32279_), .A2(new_n32278_), .B(pi1091), .ZN(new_n32280_));
  NOR2_X1    g29844(.A1(new_n31910_), .A2(pi1133), .ZN(new_n32281_));
  NOR3_X1    g29845(.A1(new_n32280_), .A2(pi0199), .A3(new_n32281_), .ZN(new_n32282_));
  NOR2_X1    g29846(.A1(new_n30015_), .A2(new_n32277_), .ZN(new_n32283_));
  NOR2_X1    g29847(.A1(new_n30014_), .A2(new_n4891_), .ZN(new_n32284_));
  OAI21_X1   g29848(.A1(new_n32283_), .A2(new_n32284_), .B(new_n3022_), .ZN(new_n32285_));
  NAND2_X1   g29849(.A1(new_n31909_), .A2(pi1135), .ZN(new_n32286_));
  AOI21_X1   g29850(.A1(new_n32285_), .A2(new_n32286_), .B(new_n8525_), .ZN(new_n32287_));
  OAI21_X1   g29851(.A1(new_n32282_), .A2(new_n32287_), .B(new_n12618_), .ZN(new_n32288_));
  NOR3_X1    g29852(.A1(new_n32280_), .A2(new_n31417_), .A3(new_n32247_), .ZN(new_n32289_));
  AOI21_X1   g29853(.A1(new_n31032_), .A2(pi1135), .B(new_n8807_), .ZN(new_n32290_));
  AOI21_X1   g29854(.A1(new_n32285_), .A2(new_n32290_), .B(new_n12618_), .ZN(new_n32291_));
  OAI21_X1   g29855(.A1(new_n32289_), .A2(pi0219), .B(new_n32291_), .ZN(new_n32292_));
  NAND2_X1   g29856(.A1(new_n8510_), .A2(new_n32229_), .ZN(new_n32293_));
  NAND3_X1   g29857(.A1(new_n29459_), .A2(pi1091), .A3(new_n32293_), .ZN(new_n32294_));
  NAND4_X1   g29858(.A1(new_n32292_), .A2(new_n27999_), .A3(new_n32288_), .A4(new_n32294_), .ZN(new_n32295_));
  NAND3_X1   g29859(.A1(new_n32295_), .A2(pi1134), .A3(new_n32276_), .ZN(new_n32296_));
  NAND2_X1   g29860(.A1(new_n32292_), .A2(new_n27999_), .ZN(new_n32297_));
  AOI21_X1   g29861(.A1(pi0200), .A2(pi1091), .B(new_n32288_), .ZN(new_n32298_));
  NAND2_X1   g29862(.A1(pi0219), .A2(pi1135), .ZN(new_n32299_));
  NAND2_X1   g29863(.A1(new_n8807_), .A2(pi1133), .ZN(new_n32300_));
  AOI21_X1   g29864(.A1(new_n32300_), .A2(new_n32299_), .B(pi0211), .ZN(new_n32301_));
  AOI21_X1   g29865(.A1(pi0199), .A2(pi1135), .B(new_n32230_), .ZN(new_n32302_));
  NOR2_X1    g29866(.A1(new_n32302_), .A2(new_n28136_), .ZN(new_n32303_));
  AOI22_X1   g29867(.A1(new_n25319_), .A2(new_n32301_), .B1(new_n6643_), .B2(new_n32303_), .ZN(new_n32304_));
  AOI21_X1   g29868(.A1(new_n32304_), .A2(pi0230), .B(pi1134), .ZN(new_n32305_));
  OAI21_X1   g29869(.A1(new_n32298_), .A2(new_n32297_), .B(new_n32305_), .ZN(new_n32306_));
  NAND2_X1   g29870(.A1(new_n32296_), .A2(new_n32306_), .ZN(po0436));
  NAND2_X1   g29871(.A1(new_n31609_), .A2(new_n8531_), .ZN(new_n32308_));
  NOR2_X1    g29872(.A1(new_n8525_), .A2(new_n4565_), .ZN(new_n32309_));
  OAI22_X1   g29873(.A1(new_n32308_), .A2(new_n32309_), .B1(new_n8531_), .B2(new_n31904_), .ZN(new_n32310_));
  NAND2_X1   g29874(.A1(new_n12618_), .A2(new_n32310_), .ZN(new_n32311_));
  NOR2_X1    g29875(.A1(pi0211), .A2(pi1135), .ZN(new_n32312_));
  AOI21_X1   g29876(.A1(pi0211), .A2(new_n4724_), .B(new_n32312_), .ZN(new_n32313_));
  AOI22_X1   g29877(.A1(new_n32313_), .A2(new_n8807_), .B1(pi1137), .B2(new_n8808_), .ZN(new_n32314_));
  NAND2_X1   g29878(.A1(new_n25319_), .A2(new_n32314_), .ZN(new_n32315_));
  AOI21_X1   g29879(.A1(new_n32315_), .A2(new_n32311_), .B(new_n27999_), .ZN(new_n32316_));
  INV_X1     g29880(.I(pi0280), .ZN(new_n32317_));
  NAND2_X1   g29881(.A1(new_n30015_), .A2(new_n32317_), .ZN(new_n32318_));
  NAND2_X1   g29882(.A1(new_n30014_), .A2(pi0914), .ZN(new_n32319_));
  AOI21_X1   g29883(.A1(new_n32318_), .A2(new_n32319_), .B(pi1091), .ZN(new_n32320_));
  NOR2_X1    g29884(.A1(new_n31910_), .A2(new_n4565_), .ZN(new_n32321_));
  OAI21_X1   g29885(.A1(new_n32320_), .A2(new_n32321_), .B(pi0199), .ZN(new_n32322_));
  NOR2_X1    g29886(.A1(new_n30004_), .A2(pi0914), .ZN(new_n32323_));
  NOR2_X1    g29887(.A1(new_n30003_), .A2(new_n32317_), .ZN(new_n32324_));
  OAI21_X1   g29888(.A1(new_n32323_), .A2(new_n32324_), .B(new_n3022_), .ZN(new_n32325_));
  NOR2_X1    g29889(.A1(new_n8531_), .A2(pi1136), .ZN(new_n32326_));
  NOR2_X1    g29890(.A1(pi0200), .A2(pi1135), .ZN(new_n32327_));
  OAI21_X1   g29891(.A1(new_n32326_), .A2(new_n32327_), .B(pi1091), .ZN(new_n32328_));
  NAND3_X1   g29892(.A1(new_n32325_), .A2(new_n8525_), .A3(new_n32328_), .ZN(new_n32329_));
  NAND3_X1   g29893(.A1(new_n32329_), .A2(new_n32322_), .A3(new_n12618_), .ZN(new_n32330_));
  OR2_X2     g29894(.A1(new_n32313_), .A2(new_n3022_), .Z(new_n32331_));
  AOI21_X1   g29895(.A1(new_n32325_), .A2(new_n32331_), .B(pi0219), .ZN(new_n32332_));
  OAI21_X1   g29896(.A1(new_n31033_), .A2(new_n4565_), .B(pi0219), .ZN(new_n32333_));
  NOR2_X1    g29897(.A1(new_n32320_), .A2(new_n32333_), .ZN(new_n32334_));
  OAI21_X1   g29898(.A1(new_n32332_), .A2(new_n32334_), .B(new_n25319_), .ZN(new_n32335_));
  NAND2_X1   g29899(.A1(new_n32335_), .A2(new_n32330_), .ZN(new_n32336_));
  AOI21_X1   g29900(.A1(new_n32336_), .A2(new_n27999_), .B(new_n32316_), .ZN(po0437));
  NOR2_X1    g29901(.A1(pi0211), .A2(pi1137), .ZN(new_n32338_));
  AOI21_X1   g29902(.A1(pi0211), .A2(new_n4408_), .B(new_n32338_), .ZN(new_n32339_));
  AOI22_X1   g29903(.A1(new_n32339_), .A2(new_n8807_), .B1(pi1139), .B2(new_n8808_), .ZN(new_n32340_));
  NOR2_X1    g29904(.A1(new_n12618_), .A2(new_n32340_), .ZN(new_n32341_));
  NOR2_X1    g29905(.A1(new_n4408_), .A2(pi0199), .ZN(new_n32342_));
  NOR2_X1    g29906(.A1(new_n32342_), .A2(new_n8531_), .ZN(new_n32343_));
  NOR2_X1    g29907(.A1(new_n8525_), .A2(new_n4238_), .ZN(new_n32344_));
  NOR3_X1    g29908(.A1(new_n32344_), .A2(new_n31902_), .A3(pi0200), .ZN(new_n32345_));
  NOR3_X1    g29909(.A1(new_n25319_), .A2(new_n32343_), .A3(new_n32345_), .ZN(new_n32346_));
  OAI21_X1   g29910(.A1(new_n32346_), .A2(new_n32341_), .B(pi0230), .ZN(new_n32347_));
  NOR2_X1    g29911(.A1(new_n31910_), .A2(new_n4238_), .ZN(new_n32348_));
  NOR3_X1    g29912(.A1(new_n25319_), .A2(new_n8525_), .A3(new_n32348_), .ZN(new_n32349_));
  AOI21_X1   g29913(.A1(pi1139), .A2(new_n31032_), .B(new_n31914_), .ZN(new_n32350_));
  NOR2_X1    g29914(.A1(new_n30014_), .A2(pi0281), .ZN(new_n32351_));
  AOI21_X1   g29915(.A1(pi0830), .A2(new_n30014_), .B(new_n32351_), .ZN(new_n32352_));
  OAI22_X1   g29916(.A1(new_n32350_), .A2(new_n32349_), .B1(pi1091), .B2(new_n32352_), .ZN(new_n32353_));
  AOI21_X1   g29917(.A1(pi1091), .A2(new_n32339_), .B(new_n29460_), .ZN(new_n32354_));
  NAND2_X1   g29918(.A1(pi0200), .A2(pi1138), .ZN(new_n32355_));
  NAND2_X1   g29919(.A1(new_n8531_), .A2(pi1137), .ZN(new_n32356_));
  AOI21_X1   g29920(.A1(new_n32356_), .A2(new_n32355_), .B(new_n3022_), .ZN(new_n32357_));
  NOR2_X1    g29921(.A1(new_n31920_), .A2(new_n32357_), .ZN(new_n32358_));
  NOR2_X1    g29922(.A1(new_n30003_), .A2(pi0281), .ZN(new_n32359_));
  AOI21_X1   g29923(.A1(pi0830), .A2(new_n30003_), .B(new_n32359_), .ZN(new_n32360_));
  OAI22_X1   g29924(.A1(new_n32358_), .A2(new_n32354_), .B1(pi1091), .B2(new_n32360_), .ZN(new_n32361_));
  NAND3_X1   g29925(.A1(new_n32361_), .A2(new_n32353_), .A3(new_n27999_), .ZN(new_n32362_));
  NAND2_X1   g29926(.A1(new_n32362_), .A2(new_n32347_), .ZN(po0438));
  NOR2_X1    g29927(.A1(pi0211), .A2(pi1138), .ZN(new_n32364_));
  AOI21_X1   g29928(.A1(pi0211), .A2(new_n4238_), .B(new_n32364_), .ZN(new_n32365_));
  AOI22_X1   g29929(.A1(new_n32365_), .A2(new_n8807_), .B1(pi1140), .B2(new_n8808_), .ZN(new_n32366_));
  NOR2_X1    g29930(.A1(new_n12618_), .A2(new_n32366_), .ZN(new_n32367_));
  AOI21_X1   g29931(.A1(new_n8525_), .A2(pi1139), .B(new_n8531_), .ZN(new_n32368_));
  NOR2_X1    g29932(.A1(new_n8525_), .A2(new_n4083_), .ZN(new_n32369_));
  NOR3_X1    g29933(.A1(new_n32369_), .A2(new_n32342_), .A3(pi0200), .ZN(new_n32370_));
  NOR2_X1    g29934(.A1(new_n32370_), .A2(new_n32368_), .ZN(new_n32371_));
  AOI21_X1   g29935(.A1(new_n12618_), .A2(new_n32371_), .B(new_n32367_), .ZN(new_n32372_));
  NAND2_X1   g29936(.A1(new_n30014_), .A2(pi0836), .ZN(new_n32373_));
  OAI21_X1   g29937(.A1(pi0282), .A2(new_n30014_), .B(new_n32373_), .ZN(new_n32374_));
  OAI21_X1   g29938(.A1(new_n4083_), .A2(new_n31033_), .B(new_n31913_), .ZN(new_n32375_));
  AOI21_X1   g29939(.A1(new_n32206_), .A2(new_n8531_), .B(new_n8525_), .ZN(new_n32376_));
  NAND2_X1   g29940(.A1(new_n12618_), .A2(new_n32376_), .ZN(new_n32377_));
  AOI22_X1   g29941(.A1(new_n32375_), .A2(new_n32377_), .B1(new_n3022_), .B2(new_n32374_), .ZN(new_n32378_));
  INV_X1     g29942(.I(pi0282), .ZN(new_n32379_));
  NAND2_X1   g29943(.A1(new_n30004_), .A2(new_n32379_), .ZN(new_n32380_));
  NAND2_X1   g29944(.A1(new_n30003_), .A2(pi0836), .ZN(new_n32381_));
  AOI21_X1   g29945(.A1(new_n32380_), .A2(new_n32381_), .B(pi1091), .ZN(new_n32382_));
  NAND2_X1   g29946(.A1(new_n32365_), .A2(pi1091), .ZN(new_n32383_));
  NOR2_X1    g29947(.A1(new_n8531_), .A2(new_n4238_), .ZN(new_n32384_));
  NOR2_X1    g29948(.A1(new_n4408_), .A2(pi0200), .ZN(new_n32385_));
  OAI21_X1   g29949(.A1(new_n32384_), .A2(new_n32385_), .B(pi1091), .ZN(new_n32386_));
  AOI22_X1   g29950(.A1(new_n31784_), .A2(new_n32386_), .B1(new_n29459_), .B2(new_n32383_), .ZN(new_n32387_));
  OAI21_X1   g29951(.A1(new_n32387_), .A2(new_n32382_), .B(new_n27999_), .ZN(new_n32388_));
  OAI22_X1   g29952(.A1(new_n32388_), .A2(new_n32378_), .B1(new_n27999_), .B2(new_n32372_), .ZN(po0439));
  NOR2_X1    g29953(.A1(new_n31992_), .A2(new_n29363_), .ZN(new_n32390_));
  AOI21_X1   g29954(.A1(pi1149), .A2(new_n31192_), .B(new_n32390_), .ZN(new_n32391_));
  OAI21_X1   g29955(.A1(new_n32391_), .A2(pi1148), .B(pi0230), .ZN(new_n32392_));
  NOR2_X1    g29956(.A1(new_n32003_), .A2(new_n32390_), .ZN(new_n32393_));
  NOR2_X1    g29957(.A1(new_n31785_), .A2(new_n29363_), .ZN(new_n32394_));
  NOR3_X1    g29958(.A1(new_n32394_), .A2(pi1149), .A3(new_n31793_), .ZN(new_n32395_));
  NOR3_X1    g29959(.A1(new_n32395_), .A2(new_n29296_), .A3(new_n32393_), .ZN(new_n32396_));
  NOR2_X1    g29960(.A1(new_n32396_), .A2(new_n32392_), .ZN(new_n32397_));
  NOR2_X1    g29961(.A1(new_n31835_), .A2(pi1147), .ZN(new_n32398_));
  AOI21_X1   g29962(.A1(new_n31838_), .A2(new_n31870_), .B(new_n29363_), .ZN(new_n32399_));
  OAI21_X1   g29963(.A1(new_n32399_), .A2(new_n32398_), .B(pi1149), .ZN(new_n32400_));
  NOR2_X1    g29964(.A1(new_n31849_), .A2(pi1147), .ZN(new_n32401_));
  NOR2_X1    g29965(.A1(new_n31884_), .A2(new_n29363_), .ZN(new_n32402_));
  OAI21_X1   g29966(.A1(new_n32401_), .A2(new_n32402_), .B(new_n29297_), .ZN(new_n32403_));
  NAND3_X1   g29967(.A1(new_n32403_), .A2(pi1148), .A3(new_n32400_), .ZN(new_n32404_));
  NOR2_X1    g29968(.A1(new_n31843_), .A2(pi1147), .ZN(new_n32405_));
  NOR2_X1    g29969(.A1(new_n31876_), .A2(new_n29363_), .ZN(new_n32406_));
  OAI21_X1   g29970(.A1(new_n32405_), .A2(new_n32406_), .B(pi1149), .ZN(new_n32407_));
  AOI21_X1   g29971(.A1(new_n31881_), .A2(new_n31880_), .B(new_n29363_), .ZN(new_n32408_));
  NAND2_X1   g29972(.A1(new_n31883_), .A2(new_n29363_), .ZN(new_n32409_));
  INV_X1     g29973(.I(new_n32409_), .ZN(new_n32410_));
  OAI21_X1   g29974(.A1(new_n32408_), .A2(new_n32410_), .B(new_n29297_), .ZN(new_n32411_));
  NAND3_X1   g29975(.A1(new_n32407_), .A2(new_n32411_), .A3(new_n29296_), .ZN(new_n32412_));
  NAND3_X1   g29976(.A1(new_n32412_), .A2(new_n32404_), .A3(new_n29930_), .ZN(new_n32413_));
  NOR2_X1    g29977(.A1(new_n31806_), .A2(pi1147), .ZN(new_n32414_));
  NOR2_X1    g29978(.A1(new_n31812_), .A2(new_n29363_), .ZN(new_n32415_));
  OAI21_X1   g29979(.A1(new_n32414_), .A2(new_n32415_), .B(pi1148), .ZN(new_n32416_));
  NOR2_X1    g29980(.A1(new_n31889_), .A2(new_n29363_), .ZN(new_n32417_));
  NOR2_X1    g29981(.A1(new_n31814_), .A2(pi1147), .ZN(new_n32418_));
  OAI21_X1   g29982(.A1(new_n32417_), .A2(new_n32418_), .B(new_n29296_), .ZN(new_n32419_));
  AND3_X2    g29983(.A1(new_n32419_), .A2(new_n29297_), .A3(new_n32416_), .Z(new_n32420_));
  NOR2_X1    g29984(.A1(new_n32420_), .A2(new_n29930_), .ZN(new_n32421_));
  NOR2_X1    g29985(.A1(new_n32031_), .A2(pi1147), .ZN(new_n32422_));
  AOI21_X1   g29986(.A1(new_n31864_), .A2(pi1147), .B(new_n32422_), .ZN(new_n32423_));
  NAND2_X1   g29987(.A1(new_n31861_), .A2(pi1147), .ZN(new_n32424_));
  OAI21_X1   g29988(.A1(pi1147), .A2(new_n31820_), .B(new_n32424_), .ZN(new_n32425_));
  AOI21_X1   g29989(.A1(new_n32425_), .A2(pi1148), .B(new_n29297_), .ZN(new_n32426_));
  OAI21_X1   g29990(.A1(new_n32423_), .A2(pi1148), .B(new_n32426_), .ZN(new_n32427_));
  AOI21_X1   g29991(.A1(new_n32421_), .A2(new_n32427_), .B(pi0230), .ZN(new_n32428_));
  AOI21_X1   g29992(.A1(new_n32413_), .A2(new_n32428_), .B(new_n32397_), .ZN(po0440));
  NAND2_X1   g29993(.A1(new_n31392_), .A2(pi1143), .ZN(new_n32430_));
  OAI22_X1   g29994(.A1(new_n29464_), .A2(new_n32430_), .B1(pi0284), .B2(new_n31392_), .ZN(po0441));
  NOR3_X1    g29995(.A1(new_n11129_), .A2(pi0286), .A3(pi0288), .ZN(new_n32432_));
  NAND2_X1   g29996(.A1(new_n32432_), .A2(new_n6347_), .ZN(new_n32433_));
  INV_X1     g29997(.I(pi0288), .ZN(new_n32434_));
  INV_X1     g29998(.I(pi0286), .ZN(new_n32435_));
  NOR2_X1    g29999(.A1(new_n8437_), .A2(new_n2612_), .ZN(new_n32436_));
  INV_X1     g30000(.I(new_n32436_), .ZN(new_n32437_));
  NOR3_X1    g30001(.A1(new_n32437_), .A2(new_n32435_), .A3(new_n10093_), .ZN(new_n32438_));
  INV_X1     g30002(.I(new_n32438_), .ZN(new_n32439_));
  NOR3_X1    g30003(.A1(new_n32439_), .A2(new_n32434_), .A3(new_n6347_), .ZN(new_n32440_));
  NAND2_X1   g30004(.A1(new_n32440_), .A2(new_n6643_), .ZN(new_n32441_));
  NAND3_X1   g30005(.A1(new_n32441_), .A2(pi0285), .A3(new_n32433_), .ZN(new_n32442_));
  NOR4_X1    g30006(.A1(new_n32439_), .A2(pi0285), .A3(new_n32434_), .A4(new_n6347_), .ZN(new_n32443_));
  NOR3_X1    g30007(.A1(new_n32440_), .A2(new_n6346_), .A3(new_n32437_), .ZN(new_n32444_));
  OAI21_X1   g30008(.A1(new_n32444_), .A2(new_n32443_), .B(new_n6643_), .ZN(new_n32445_));
  AOI21_X1   g30009(.A1(new_n32445_), .A2(new_n32442_), .B(pi0793), .ZN(po0442));
  OAI21_X1   g30010(.A1(new_n6348_), .A2(pi0286), .B(new_n32434_), .ZN(new_n32447_));
  OAI21_X1   g30011(.A1(new_n32436_), .A2(new_n11129_), .B(pi0286), .ZN(new_n32448_));
  NOR3_X1    g30012(.A1(new_n32436_), .A2(pi0286), .A3(new_n11129_), .ZN(new_n32449_));
  INV_X1     g30013(.I(new_n32449_), .ZN(new_n32450_));
  AOI21_X1   g30014(.A1(new_n32450_), .A2(new_n32448_), .B(new_n32447_), .ZN(new_n32451_));
  AOI21_X1   g30015(.A1(new_n32436_), .A2(new_n11129_), .B(pi0286), .ZN(new_n32452_));
  NOR3_X1    g30016(.A1(new_n32438_), .A2(new_n32434_), .A3(new_n32452_), .ZN(new_n32453_));
  NOR3_X1    g30017(.A1(new_n32453_), .A2(new_n32451_), .A3(po1038), .ZN(new_n32454_));
  NOR2_X1    g30018(.A1(new_n11129_), .A2(new_n32447_), .ZN(new_n32455_));
  XOR2_X1    g30019(.A1(new_n32455_), .A2(pi0286), .Z(new_n32456_));
  NOR2_X1    g30020(.A1(new_n32456_), .A2(new_n6643_), .ZN(new_n32457_));
  NOR3_X1    g30021(.A1(new_n32454_), .A2(pi0793), .A3(new_n32457_), .ZN(po0443));
  AOI21_X1   g30022(.A1(new_n8282_), .A2(pi0457), .B(pi0332), .ZN(po0444));
  NOR2_X1    g30023(.A1(new_n32437_), .A2(po1038), .ZN(po0637));
  AOI21_X1   g30024(.A1(pi0288), .A2(new_n11129_), .B(new_n32455_), .ZN(new_n32461_));
  XOR2_X1    g30025(.A1(po0637), .A2(new_n32461_), .Z(new_n32462_));
  NOR2_X1    g30026(.A1(new_n32462_), .A2(pi0793), .ZN(po0445));
  NOR2_X1    g30027(.A1(new_n32450_), .A2(new_n6347_), .ZN(new_n32464_));
  AOI21_X1   g30028(.A1(new_n32449_), .A2(pi0285), .B(pi0289), .ZN(new_n32465_));
  OAI21_X1   g30029(.A1(new_n32464_), .A2(new_n32465_), .B(new_n32434_), .ZN(new_n32466_));
  NAND2_X1   g30030(.A1(new_n32439_), .A2(pi0289), .ZN(new_n32467_));
  NAND2_X1   g30031(.A1(new_n32438_), .A2(new_n6347_), .ZN(new_n32468_));
  NAND3_X1   g30032(.A1(new_n32467_), .A2(pi0288), .A3(new_n32468_), .ZN(new_n32469_));
  AOI21_X1   g30033(.A1(new_n32469_), .A2(new_n32466_), .B(po1038), .ZN(new_n32470_));
  NOR2_X1    g30034(.A1(new_n32433_), .A2(new_n6346_), .ZN(new_n32471_));
  OAI21_X1   g30035(.A1(new_n32432_), .A2(new_n6347_), .B(po1038), .ZN(new_n32472_));
  NOR2_X1    g30036(.A1(new_n32471_), .A2(new_n32472_), .ZN(new_n32473_));
  NOR3_X1    g30037(.A1(new_n32470_), .A2(pi0793), .A3(new_n32473_), .ZN(po0446));
  INV_X1     g30038(.I(pi1048), .ZN(new_n32475_));
  NAND2_X1   g30039(.A1(pi0290), .A2(pi0476), .ZN(new_n32476_));
  OAI21_X1   g30040(.A1(pi0476), .A2(new_n32475_), .B(new_n32476_), .ZN(po0447));
  INV_X1     g30041(.I(pi1049), .ZN(new_n32478_));
  NAND2_X1   g30042(.A1(pi0291), .A2(pi0476), .ZN(new_n32479_));
  OAI21_X1   g30043(.A1(pi0476), .A2(new_n32478_), .B(new_n32479_), .ZN(po0448));
  INV_X1     g30044(.I(pi1084), .ZN(new_n32481_));
  NAND2_X1   g30045(.A1(pi0292), .A2(pi0476), .ZN(new_n32482_));
  OAI21_X1   g30046(.A1(pi0476), .A2(new_n32481_), .B(new_n32482_), .ZN(po0449));
  INV_X1     g30047(.I(pi1059), .ZN(new_n32484_));
  NAND2_X1   g30048(.A1(pi0293), .A2(pi0476), .ZN(new_n32485_));
  OAI21_X1   g30049(.A1(pi0476), .A2(new_n32484_), .B(new_n32485_), .ZN(po0450));
  INV_X1     g30050(.I(pi1072), .ZN(new_n32487_));
  NAND2_X1   g30051(.A1(pi0294), .A2(pi0476), .ZN(new_n32488_));
  OAI21_X1   g30052(.A1(pi0476), .A2(new_n32487_), .B(new_n32488_), .ZN(po0451));
  INV_X1     g30053(.I(pi1053), .ZN(new_n32490_));
  NAND2_X1   g30054(.A1(pi0295), .A2(pi0476), .ZN(new_n32491_));
  OAI21_X1   g30055(.A1(pi0476), .A2(new_n32490_), .B(new_n32491_), .ZN(po0452));
  INV_X1     g30056(.I(pi1037), .ZN(new_n32493_));
  NAND2_X1   g30057(.A1(pi0296), .A2(pi0476), .ZN(new_n32494_));
  OAI21_X1   g30058(.A1(pi0476), .A2(new_n32493_), .B(new_n32494_), .ZN(po0453));
  INV_X1     g30059(.I(pi1044), .ZN(new_n32496_));
  NAND2_X1   g30060(.A1(pi0297), .A2(pi0476), .ZN(new_n32497_));
  OAI21_X1   g30061(.A1(pi0476), .A2(new_n32496_), .B(new_n32497_), .ZN(po0454));
  NAND2_X1   g30062(.A1(pi0298), .A2(pi0478), .ZN(new_n32499_));
  OAI21_X1   g30063(.A1(pi0478), .A2(new_n32496_), .B(new_n32499_), .ZN(po0455));
  NOR2_X1    g30064(.A1(new_n2530_), .A2(new_n5499_), .ZN(new_n32501_));
  NOR4_X1    g30065(.A1(new_n10505_), .A2(pi0054), .A3(new_n2787_), .A4(new_n8254_), .ZN(new_n32502_));
  NOR3_X1    g30066(.A1(new_n7266_), .A2(new_n2606_), .A3(new_n5792_), .ZN(new_n32503_));
  OAI21_X1   g30067(.A1(new_n32502_), .A2(new_n32501_), .B(new_n32503_), .ZN(new_n32504_));
  AOI21_X1   g30068(.A1(new_n32504_), .A2(new_n2627_), .B(new_n9097_), .ZN(po0456));
  INV_X1     g30069(.I(pi0312), .ZN(new_n32506_));
  NOR3_X1    g30070(.A1(new_n8189_), .A2(new_n2582_), .A3(pi0059), .ZN(new_n32507_));
  NAND2_X1   g30071(.A1(new_n32507_), .A2(new_n32506_), .ZN(new_n32508_));
  NOR2_X1    g30072(.A1(new_n32508_), .A2(pi0300), .ZN(new_n32509_));
  INV_X1     g30073(.I(new_n32509_), .ZN(new_n32510_));
  NAND2_X1   g30074(.A1(new_n32508_), .A2(pi0300), .ZN(new_n32511_));
  NAND3_X1   g30075(.A1(new_n32510_), .A2(new_n2602_), .A3(new_n32511_), .ZN(po0457));
  INV_X1     g30076(.I(pi0301), .ZN(new_n32513_));
  NAND2_X1   g30077(.A1(new_n32510_), .A2(new_n32513_), .ZN(new_n32514_));
  NOR2_X1    g30078(.A1(new_n32510_), .A2(new_n32513_), .ZN(new_n32515_));
  INV_X1     g30079(.I(new_n32515_), .ZN(new_n32516_));
  AOI21_X1   g30080(.A1(new_n32516_), .A2(new_n32514_), .B(pi0055), .ZN(po0458));
  NAND2_X1   g30081(.A1(new_n25319_), .A2(new_n3305_), .ZN(new_n32518_));
  OAI21_X1   g30082(.A1(pi0222), .A2(pi0223), .B(pi0937), .ZN(new_n32519_));
  NOR2_X1    g30083(.A1(new_n5217_), .A2(po1038), .ZN(new_n32520_));
  NAND2_X1   g30084(.A1(new_n3346_), .A2(pi0273), .ZN(new_n32521_));
  NAND3_X1   g30085(.A1(new_n32520_), .A2(new_n32519_), .A3(new_n32521_), .ZN(new_n32522_));
  AOI21_X1   g30086(.A1(new_n32518_), .A2(new_n32522_), .B(new_n25327_), .ZN(new_n32523_));
  INV_X1     g30087(.I(pi0937), .ZN(new_n32524_));
  NOR2_X1    g30088(.A1(new_n2559_), .A2(new_n2614_), .ZN(new_n32525_));
  NOR2_X1    g30089(.A1(new_n6762_), .A2(new_n2443_), .ZN(new_n32526_));
  AOI22_X1   g30090(.A1(new_n32526_), .A2(new_n32524_), .B1(new_n29999_), .B2(new_n32525_), .ZN(new_n32527_));
  OAI22_X1   g30091(.A1(new_n12618_), .A2(new_n32527_), .B1(new_n32522_), .B2(new_n2641_), .ZN(new_n32528_));
  INV_X1     g30092(.I(new_n32520_), .ZN(new_n32529_));
  OAI21_X1   g30093(.A1(new_n5200_), .A2(new_n12618_), .B(new_n32529_), .ZN(new_n32530_));
  NOR2_X1    g30094(.A1(new_n32530_), .A2(pi1148), .ZN(new_n32531_));
  NOR3_X1    g30095(.A1(new_n32531_), .A2(new_n32523_), .A3(new_n32528_), .ZN(po0459));
  NAND2_X1   g30096(.A1(pi0303), .A2(pi0478), .ZN(new_n32533_));
  OAI21_X1   g30097(.A1(pi0478), .A2(new_n32478_), .B(new_n32533_), .ZN(po0460));
  NAND2_X1   g30098(.A1(pi0304), .A2(pi0478), .ZN(new_n32535_));
  OAI21_X1   g30099(.A1(pi0478), .A2(new_n32475_), .B(new_n32535_), .ZN(po0461));
  NAND2_X1   g30100(.A1(pi0305), .A2(pi0478), .ZN(new_n32537_));
  OAI21_X1   g30101(.A1(pi0478), .A2(new_n32481_), .B(new_n32537_), .ZN(po0462));
  NAND2_X1   g30102(.A1(pi0306), .A2(pi0478), .ZN(new_n32539_));
  OAI21_X1   g30103(.A1(pi0478), .A2(new_n32484_), .B(new_n32539_), .ZN(po0463));
  NAND2_X1   g30104(.A1(pi0307), .A2(pi0478), .ZN(new_n32541_));
  OAI21_X1   g30105(.A1(pi0478), .A2(new_n32490_), .B(new_n32541_), .ZN(po0464));
  NAND2_X1   g30106(.A1(pi0308), .A2(pi0478), .ZN(new_n32543_));
  OAI21_X1   g30107(.A1(pi0478), .A2(new_n32493_), .B(new_n32543_), .ZN(po0465));
  NAND2_X1   g30108(.A1(pi0309), .A2(pi0478), .ZN(new_n32545_));
  OAI21_X1   g30109(.A1(pi0478), .A2(new_n32487_), .B(new_n32545_), .ZN(po0466));
  INV_X1     g30110(.I(pi0934), .ZN(new_n32547_));
  AOI22_X1   g30111(.A1(new_n3346_), .A2(new_n30000_), .B1(pi0222), .B2(new_n32547_), .ZN(new_n32548_));
  AOI22_X1   g30112(.A1(new_n25319_), .A2(new_n3305_), .B1(new_n32520_), .B2(new_n32548_), .ZN(new_n32549_));
  NOR2_X1    g30113(.A1(new_n2614_), .A2(pi0221), .ZN(new_n32550_));
  AOI22_X1   g30114(.A1(new_n2559_), .A2(pi0934), .B1(new_n32550_), .B2(pi0271), .ZN(new_n32551_));
  NOR2_X1    g30115(.A1(new_n12618_), .A2(new_n5200_), .ZN(new_n32552_));
  NAND2_X1   g30116(.A1(new_n32552_), .A2(new_n3304_), .ZN(new_n32553_));
  OAI21_X1   g30117(.A1(new_n32551_), .A2(new_n32553_), .B(new_n32549_), .ZN(new_n32554_));
  NOR2_X1    g30118(.A1(new_n32530_), .A2(new_n29363_), .ZN(new_n32555_));
  OAI21_X1   g30119(.A1(new_n32555_), .A2(new_n32554_), .B(new_n25326_), .ZN(new_n32556_));
  OAI21_X1   g30120(.A1(new_n32529_), .A2(new_n32548_), .B(pi1147), .ZN(new_n32557_));
  AOI21_X1   g30121(.A1(new_n2643_), .A2(new_n12618_), .B(new_n32557_), .ZN(new_n32558_));
  NAND2_X1   g30122(.A1(new_n32552_), .A2(new_n32551_), .ZN(new_n32559_));
  AOI22_X1   g30123(.A1(new_n32552_), .A2(new_n3304_), .B1(new_n2642_), .B2(new_n32520_), .ZN(new_n32560_));
  NOR2_X1    g30124(.A1(new_n32560_), .A2(pi1147), .ZN(new_n32561_));
  AOI22_X1   g30125(.A1(new_n32558_), .A2(new_n32559_), .B1(new_n32554_), .B2(new_n32561_), .ZN(new_n32562_));
  OAI21_X1   g30126(.A1(new_n32562_), .A2(new_n25326_), .B(new_n32556_), .ZN(po0467));
  XOR2_X1    g30127(.A1(new_n32515_), .A2(pi0311), .Z(new_n32564_));
  NOR2_X1    g30128(.A1(new_n32564_), .A2(pi0055), .ZN(po0468));
  XOR2_X1    g30129(.A1(new_n32507_), .A2(new_n32506_), .Z(new_n32566_));
  NOR2_X1    g30130(.A1(new_n32566_), .A2(pi0055), .ZN(po0469));
  NOR2_X1    g30131(.A1(new_n10531_), .A2(new_n8241_), .ZN(new_n32568_));
  NOR2_X1    g30132(.A1(new_n32568_), .A2(new_n8262_), .ZN(new_n32569_));
  NAND2_X1   g30133(.A1(new_n8414_), .A2(new_n10527_), .ZN(new_n32570_));
  NAND3_X1   g30134(.A1(new_n32569_), .A2(po1110), .A3(new_n32570_), .ZN(new_n32571_));
  OAI21_X1   g30135(.A1(pi0313), .A2(po1110), .B(new_n32571_), .ZN(po0470));
  NAND2_X1   g30136(.A1(new_n7265_), .A2(new_n5492_), .ZN(new_n32573_));
  NOR2_X1    g30137(.A1(new_n12135_), .A2(new_n2627_), .ZN(new_n32574_));
  AOI21_X1   g30138(.A1(new_n11303_), .A2(new_n2627_), .B(new_n32574_), .ZN(new_n32575_));
  OAI21_X1   g30139(.A1(new_n32575_), .A2(new_n3271_), .B(new_n12036_), .ZN(new_n32576_));
  NOR2_X1    g30140(.A1(new_n8256_), .A2(new_n2567_), .ZN(new_n32577_));
  AOI22_X1   g30141(.A1(new_n32576_), .A2(new_n32577_), .B1(new_n11172_), .B2(new_n32573_), .ZN(new_n32578_));
  NOR4_X1    g30142(.A1(new_n32578_), .A2(pi0125), .A3(pi0133), .A4(new_n11179_), .ZN(po0471));
  INV_X1     g30143(.I(po0637), .ZN(new_n32580_));
  NOR2_X1    g30144(.A1(new_n32580_), .A2(pi0340), .ZN(new_n32581_));
  NAND2_X1   g30145(.A1(new_n32581_), .A2(pi1080), .ZN(new_n32582_));
  OAI21_X1   g30146(.A1(new_n6506_), .A2(new_n32581_), .B(new_n32582_), .ZN(po0472));
  INV_X1     g30147(.I(pi0316), .ZN(new_n32584_));
  NAND2_X1   g30148(.A1(new_n32581_), .A2(pi1047), .ZN(new_n32585_));
  OAI21_X1   g30149(.A1(new_n32584_), .A2(new_n32581_), .B(new_n32585_), .ZN(po0473));
  NOR2_X1    g30150(.A1(new_n32580_), .A2(pi0330), .ZN(new_n32587_));
  NAND2_X1   g30151(.A1(new_n32587_), .A2(pi1078), .ZN(new_n32588_));
  OAI21_X1   g30152(.A1(new_n6602_), .A2(new_n32587_), .B(new_n32588_), .ZN(po0474));
  INV_X1     g30153(.I(pi1074), .ZN(new_n32590_));
  NOR2_X1    g30154(.A1(new_n32580_), .A2(pi0341), .ZN(new_n32591_));
  INV_X1     g30155(.I(new_n32591_), .ZN(new_n32592_));
  NAND2_X1   g30156(.A1(new_n32592_), .A2(pi0318), .ZN(new_n32593_));
  OAI21_X1   g30157(.A1(new_n32590_), .A2(new_n32592_), .B(new_n32593_), .ZN(po0475));
  NAND2_X1   g30158(.A1(new_n32591_), .A2(pi1072), .ZN(new_n32595_));
  OAI21_X1   g30159(.A1(new_n6389_), .A2(new_n32591_), .B(new_n32595_), .ZN(po0476));
  NAND2_X1   g30160(.A1(new_n32581_), .A2(pi1048), .ZN(new_n32597_));
  OAI21_X1   g30161(.A1(new_n6473_), .A2(new_n32581_), .B(new_n32597_), .ZN(po0477));
  INV_X1     g30162(.I(pi0321), .ZN(new_n32599_));
  NAND2_X1   g30163(.A1(new_n32581_), .A2(pi1058), .ZN(new_n32600_));
  OAI21_X1   g30164(.A1(new_n32599_), .A2(new_n32581_), .B(new_n32600_), .ZN(po0478));
  NAND2_X1   g30165(.A1(new_n32581_), .A2(pi1051), .ZN(new_n32602_));
  OAI21_X1   g30166(.A1(new_n6503_), .A2(new_n32581_), .B(new_n32602_), .ZN(po0479));
  NAND2_X1   g30167(.A1(new_n32581_), .A2(pi1065), .ZN(new_n32604_));
  OAI21_X1   g30168(.A1(new_n6451_), .A2(new_n32581_), .B(new_n32604_), .ZN(po0480));
  NAND2_X1   g30169(.A1(new_n32591_), .A2(pi1086), .ZN(new_n32606_));
  OAI21_X1   g30170(.A1(new_n6385_), .A2(new_n32591_), .B(new_n32606_), .ZN(po0481));
  INV_X1     g30171(.I(pi1063), .ZN(new_n32608_));
  NAND2_X1   g30172(.A1(new_n32592_), .A2(pi0325), .ZN(new_n32609_));
  OAI21_X1   g30173(.A1(new_n32608_), .A2(new_n32592_), .B(new_n32609_), .ZN(po0482));
  INV_X1     g30174(.I(pi0326), .ZN(new_n32611_));
  NAND2_X1   g30175(.A1(new_n32591_), .A2(pi1057), .ZN(new_n32612_));
  OAI21_X1   g30176(.A1(new_n32611_), .A2(new_n32591_), .B(new_n32612_), .ZN(po0483));
  INV_X1     g30177(.I(pi1040), .ZN(new_n32614_));
  INV_X1     g30178(.I(new_n32581_), .ZN(new_n32615_));
  NAND2_X1   g30179(.A1(new_n32615_), .A2(pi0327), .ZN(new_n32616_));
  OAI21_X1   g30180(.A1(new_n32614_), .A2(new_n32615_), .B(new_n32616_), .ZN(po0484));
  INV_X1     g30181(.I(pi0328), .ZN(new_n32618_));
  NAND2_X1   g30182(.A1(new_n32591_), .A2(pi1058), .ZN(new_n32619_));
  OAI21_X1   g30183(.A1(new_n32618_), .A2(new_n32591_), .B(new_n32619_), .ZN(po0485));
  INV_X1     g30184(.I(pi0329), .ZN(new_n32621_));
  NAND2_X1   g30185(.A1(new_n32591_), .A2(pi1043), .ZN(new_n32622_));
  OAI21_X1   g30186(.A1(new_n32621_), .A2(new_n32591_), .B(new_n32622_), .ZN(po0486));
  NOR2_X1    g30187(.A1(new_n3080_), .A2(new_n3040_), .ZN(new_n32624_));
  INV_X1     g30188(.I(new_n32624_), .ZN(new_n32625_));
  OR2_X2     g30189(.A1(po0637), .A2(pi0330), .Z(new_n32626_));
  AOI21_X1   g30190(.A1(new_n32615_), .A2(new_n32626_), .B(new_n32625_), .ZN(po0487));
  OR2_X2     g30191(.A1(po0637), .A2(pi0331), .Z(new_n32628_));
  AOI21_X1   g30192(.A1(new_n32592_), .A2(new_n32628_), .B(new_n32625_), .ZN(po0488));
  NAND2_X1   g30193(.A1(new_n8909_), .A2(new_n10355_), .ZN(new_n32630_));
  AOI21_X1   g30194(.A1(new_n32630_), .A2(new_n6676_), .B(pi0070), .ZN(new_n32631_));
  NAND2_X1   g30195(.A1(new_n7433_), .A2(pi0332), .ZN(new_n32632_));
  OAI22_X1   g30196(.A1(new_n32631_), .A2(new_n32632_), .B1(new_n8909_), .B2(new_n10356_), .ZN(new_n32633_));
  NAND2_X1   g30197(.A1(new_n8637_), .A2(pi0039), .ZN(new_n32634_));
  OAI21_X1   g30198(.A1(new_n32633_), .A2(pi0039), .B(new_n32634_), .ZN(new_n32635_));
  AOI21_X1   g30199(.A1(new_n32635_), .A2(new_n3265_), .B(new_n27962_), .ZN(po0489));
  NAND2_X1   g30200(.A1(new_n32591_), .A2(pi1040), .ZN(new_n32637_));
  OAI21_X1   g30201(.A1(new_n6422_), .A2(new_n32591_), .B(new_n32637_), .ZN(po0490));
  NAND2_X1   g30202(.A1(new_n32591_), .A2(pi1065), .ZN(new_n32639_));
  OAI21_X1   g30203(.A1(new_n7197_), .A2(new_n32591_), .B(new_n32639_), .ZN(po0491));
  NAND2_X1   g30204(.A1(new_n32592_), .A2(pi0335), .ZN(new_n32641_));
  OAI21_X1   g30205(.A1(new_n31362_), .A2(new_n32592_), .B(new_n32641_), .ZN(po0492));
  INV_X1     g30206(.I(pi0336), .ZN(new_n32643_));
  NAND2_X1   g30207(.A1(new_n32587_), .A2(pi1070), .ZN(new_n32644_));
  OAI21_X1   g30208(.A1(new_n32643_), .A2(new_n32587_), .B(new_n32644_), .ZN(po0493));
  INV_X1     g30209(.I(new_n32587_), .ZN(new_n32646_));
  NAND2_X1   g30210(.A1(new_n32646_), .A2(pi0337), .ZN(new_n32647_));
  OAI21_X1   g30211(.A1(new_n32496_), .A2(new_n32646_), .B(new_n32647_), .ZN(po0494));
  INV_X1     g30212(.I(pi0338), .ZN(new_n32649_));
  NAND2_X1   g30213(.A1(new_n32587_), .A2(pi1072), .ZN(new_n32650_));
  OAI21_X1   g30214(.A1(new_n32649_), .A2(new_n32587_), .B(new_n32650_), .ZN(po0495));
  NAND2_X1   g30215(.A1(new_n32587_), .A2(pi1086), .ZN(new_n32652_));
  NAND2_X1   g30216(.A1(new_n32646_), .A2(pi0339), .ZN(new_n32653_));
  NAND2_X1   g30217(.A1(new_n32653_), .A2(new_n32652_), .ZN(po0496));
  INV_X1     g30218(.I(pi0340), .ZN(new_n32655_));
  AOI21_X1   g30219(.A1(po1038), .A2(new_n32655_), .B(new_n32625_), .ZN(new_n32656_));
  NAND2_X1   g30220(.A1(new_n32436_), .A2(pi0331), .ZN(new_n32657_));
  OAI21_X1   g30221(.A1(new_n32655_), .A2(new_n32436_), .B(new_n32657_), .ZN(new_n32658_));
  OAI21_X1   g30222(.A1(new_n32658_), .A2(po1038), .B(new_n32656_), .ZN(po0497));
  OR2_X2     g30223(.A1(po0637), .A2(pi0341), .Z(new_n32660_));
  AOI21_X1   g30224(.A1(new_n32646_), .A2(new_n32660_), .B(new_n32625_), .ZN(po0498));
  NAND2_X1   g30225(.A1(new_n32581_), .A2(pi1049), .ZN(new_n32662_));
  OAI21_X1   g30226(.A1(new_n6469_), .A2(new_n32581_), .B(new_n32662_), .ZN(po0499));
  NAND2_X1   g30227(.A1(new_n32615_), .A2(pi0343), .ZN(new_n32664_));
  OAI21_X1   g30228(.A1(new_n31356_), .A2(new_n32615_), .B(new_n32664_), .ZN(po0500));
  NAND2_X1   g30229(.A1(new_n32581_), .A2(pi1069), .ZN(new_n32666_));
  OAI21_X1   g30230(.A1(new_n6459_), .A2(new_n32581_), .B(new_n32666_), .ZN(po0501));
  NAND2_X1   g30231(.A1(new_n32581_), .A2(pi1039), .ZN(new_n32668_));
  OAI21_X1   g30232(.A1(new_n6447_), .A2(new_n32581_), .B(new_n32668_), .ZN(po0502));
  NAND2_X1   g30233(.A1(new_n32581_), .A2(pi1067), .ZN(new_n32670_));
  OAI21_X1   g30234(.A1(new_n6448_), .A2(new_n32581_), .B(new_n32670_), .ZN(po0503));
  INV_X1     g30235(.I(pi1055), .ZN(new_n32672_));
  NAND2_X1   g30236(.A1(new_n32615_), .A2(pi0347), .ZN(new_n32673_));
  OAI21_X1   g30237(.A1(new_n32672_), .A2(new_n32615_), .B(new_n32673_), .ZN(po0504));
  INV_X1     g30238(.I(pi1087), .ZN(new_n32675_));
  NAND2_X1   g30239(.A1(new_n32615_), .A2(pi0348), .ZN(new_n32676_));
  OAI21_X1   g30240(.A1(new_n32675_), .A2(new_n32615_), .B(new_n32676_), .ZN(po0505));
  INV_X1     g30241(.I(pi0349), .ZN(new_n32678_));
  NAND2_X1   g30242(.A1(new_n32581_), .A2(pi1043), .ZN(new_n32679_));
  OAI21_X1   g30243(.A1(new_n32678_), .A2(new_n32581_), .B(new_n32679_), .ZN(po0506));
  NAND2_X1   g30244(.A1(new_n32581_), .A2(pi1035), .ZN(new_n32681_));
  OAI21_X1   g30245(.A1(new_n7086_), .A2(new_n32581_), .B(new_n32681_), .ZN(po0507));
  NAND2_X1   g30246(.A1(new_n32581_), .A2(pi1079), .ZN(new_n32683_));
  OAI21_X1   g30247(.A1(new_n6443_), .A2(new_n32581_), .B(new_n32683_), .ZN(po0508));
  INV_X1     g30248(.I(pi1078), .ZN(new_n32685_));
  NAND2_X1   g30249(.A1(new_n32615_), .A2(pi0352), .ZN(new_n32686_));
  OAI21_X1   g30250(.A1(new_n32685_), .A2(new_n32615_), .B(new_n32686_), .ZN(po0509));
  INV_X1     g30251(.I(pi0353), .ZN(new_n32688_));
  NAND2_X1   g30252(.A1(new_n32581_), .A2(pi1063), .ZN(new_n32689_));
  OAI21_X1   g30253(.A1(new_n32688_), .A2(new_n32581_), .B(new_n32689_), .ZN(po0510));
  NAND2_X1   g30254(.A1(new_n32581_), .A2(pi1045), .ZN(new_n32691_));
  OAI21_X1   g30255(.A1(new_n9784_), .A2(new_n32581_), .B(new_n32691_), .ZN(po0511));
  NAND2_X1   g30256(.A1(new_n32581_), .A2(pi1084), .ZN(new_n32693_));
  OAI21_X1   g30257(.A1(new_n6485_), .A2(new_n32581_), .B(new_n32693_), .ZN(po0512));
  NAND2_X1   g30258(.A1(new_n32581_), .A2(pi1081), .ZN(new_n32695_));
  OAI21_X1   g30259(.A1(new_n9785_), .A2(new_n32581_), .B(new_n32695_), .ZN(po0513));
  INV_X1     g30260(.I(pi1076), .ZN(new_n32697_));
  NAND2_X1   g30261(.A1(new_n32615_), .A2(pi0357), .ZN(new_n32698_));
  OAI21_X1   g30262(.A1(new_n32697_), .A2(new_n32615_), .B(new_n32698_), .ZN(po0514));
  NAND2_X1   g30263(.A1(new_n32581_), .A2(pi1071), .ZN(new_n32700_));
  NAND2_X1   g30264(.A1(new_n32615_), .A2(pi0358), .ZN(new_n32701_));
  NAND2_X1   g30265(.A1(new_n32701_), .A2(new_n32700_), .ZN(po0515));
  NAND2_X1   g30266(.A1(new_n32581_), .A2(pi1068), .ZN(new_n32703_));
  OAI21_X1   g30267(.A1(new_n6501_), .A2(new_n32581_), .B(new_n32703_), .ZN(po0516));
  NAND2_X1   g30268(.A1(new_n32581_), .A2(pi1042), .ZN(new_n32705_));
  OAI21_X1   g30269(.A1(new_n6542_), .A2(new_n32581_), .B(new_n32705_), .ZN(po0517));
  INV_X1     g30270(.I(pi0361), .ZN(new_n32707_));
  NAND2_X1   g30271(.A1(new_n32581_), .A2(pi1059), .ZN(new_n32708_));
  OAI21_X1   g30272(.A1(new_n32707_), .A2(new_n32581_), .B(new_n32708_), .ZN(po0518));
  NAND2_X1   g30273(.A1(new_n32581_), .A2(pi1070), .ZN(new_n32710_));
  OAI21_X1   g30274(.A1(new_n6461_), .A2(new_n32581_), .B(new_n32710_), .ZN(po0519));
  NAND2_X1   g30275(.A1(new_n32587_), .A2(pi1049), .ZN(new_n32712_));
  OAI21_X1   g30276(.A1(new_n6562_), .A2(new_n32587_), .B(new_n32712_), .ZN(po0520));
  NAND2_X1   g30277(.A1(new_n32646_), .A2(pi0364), .ZN(new_n32714_));
  OAI21_X1   g30278(.A1(new_n31356_), .A2(new_n32646_), .B(new_n32714_), .ZN(po0521));
  NAND2_X1   g30279(.A1(new_n32646_), .A2(pi0365), .ZN(new_n32716_));
  OAI21_X1   g30280(.A1(new_n31350_), .A2(new_n32646_), .B(new_n32716_), .ZN(po0522));
  NAND2_X1   g30281(.A1(new_n32587_), .A2(pi1069), .ZN(new_n32718_));
  OAI21_X1   g30282(.A1(new_n6577_), .A2(new_n32587_), .B(new_n32718_), .ZN(po0523));
  NAND2_X1   g30283(.A1(new_n32587_), .A2(pi1039), .ZN(new_n32720_));
  OAI21_X1   g30284(.A1(new_n6583_), .A2(new_n32587_), .B(new_n32720_), .ZN(po0524));
  INV_X1     g30285(.I(pi1067), .ZN(new_n32722_));
  NAND2_X1   g30286(.A1(new_n32646_), .A2(pi0368), .ZN(new_n32723_));
  OAI21_X1   g30287(.A1(new_n32722_), .A2(new_n32646_), .B(new_n32723_), .ZN(po0525));
  NAND2_X1   g30288(.A1(new_n32587_), .A2(pi1080), .ZN(new_n32725_));
  OAI21_X1   g30289(.A1(new_n9882_), .A2(new_n32587_), .B(new_n32725_), .ZN(po0526));
  INV_X1     g30290(.I(pi0370), .ZN(new_n32727_));
  NAND2_X1   g30291(.A1(new_n32587_), .A2(pi1055), .ZN(new_n32728_));
  OAI21_X1   g30292(.A1(new_n32727_), .A2(new_n32587_), .B(new_n32728_), .ZN(po0527));
  NAND2_X1   g30293(.A1(new_n32587_), .A2(pi1051), .ZN(new_n32730_));
  OAI21_X1   g30294(.A1(new_n7049_), .A2(new_n32587_), .B(new_n32730_), .ZN(po0528));
  NAND2_X1   g30295(.A1(new_n32587_), .A2(pi1048), .ZN(new_n32732_));
  OAI21_X1   g30296(.A1(new_n6559_), .A2(new_n32587_), .B(new_n32732_), .ZN(po0529));
  NAND2_X1   g30297(.A1(new_n32587_), .A2(pi1087), .ZN(new_n32734_));
  OAI21_X1   g30298(.A1(new_n7234_), .A2(new_n32587_), .B(new_n32734_), .ZN(po0530));
  NAND2_X1   g30299(.A1(new_n32587_), .A2(pi1035), .ZN(new_n32736_));
  OAI21_X1   g30300(.A1(new_n7051_), .A2(new_n32587_), .B(new_n32736_), .ZN(po0531));
  NAND2_X1   g30301(.A1(new_n32587_), .A2(pi1047), .ZN(new_n32738_));
  OAI21_X1   g30302(.A1(new_n7240_), .A2(new_n32587_), .B(new_n32738_), .ZN(po0532));
  INV_X1     g30303(.I(pi1079), .ZN(new_n32740_));
  NAND2_X1   g30304(.A1(new_n32646_), .A2(pi0376), .ZN(new_n32741_));
  OAI21_X1   g30305(.A1(new_n32740_), .A2(new_n32646_), .B(new_n32741_), .ZN(po0533));
  NAND2_X1   g30306(.A1(new_n32587_), .A2(pi1074), .ZN(new_n32743_));
  OAI21_X1   g30307(.A1(new_n6594_), .A2(new_n32587_), .B(new_n32743_), .ZN(po0534));
  NAND2_X1   g30308(.A1(new_n32587_), .A2(pi1063), .ZN(new_n32745_));
  OAI21_X1   g30309(.A1(new_n6599_), .A2(new_n32587_), .B(new_n32745_), .ZN(po0535));
  INV_X1     g30310(.I(pi0379), .ZN(new_n32747_));
  NAND2_X1   g30311(.A1(new_n32587_), .A2(pi1045), .ZN(new_n32748_));
  OAI21_X1   g30312(.A1(new_n32747_), .A2(new_n32587_), .B(new_n32748_), .ZN(po0536));
  INV_X1     g30313(.I(pi0380), .ZN(new_n32750_));
  NAND2_X1   g30314(.A1(new_n32587_), .A2(pi1084), .ZN(new_n32751_));
  OAI21_X1   g30315(.A1(new_n32750_), .A2(new_n32587_), .B(new_n32751_), .ZN(po0537));
  INV_X1     g30316(.I(pi1081), .ZN(new_n32753_));
  NAND2_X1   g30317(.A1(new_n32646_), .A2(pi0381), .ZN(new_n32754_));
  OAI21_X1   g30318(.A1(new_n32753_), .A2(new_n32646_), .B(new_n32754_), .ZN(po0538));
  NAND2_X1   g30319(.A1(new_n32646_), .A2(pi0382), .ZN(new_n32756_));
  OAI21_X1   g30320(.A1(new_n32697_), .A2(new_n32646_), .B(new_n32756_), .ZN(po0539));
  NAND2_X1   g30321(.A1(new_n32587_), .A2(pi1071), .ZN(new_n32758_));
  OAI21_X1   g30322(.A1(new_n6575_), .A2(new_n32587_), .B(new_n32758_), .ZN(po0540));
  NAND2_X1   g30323(.A1(new_n32587_), .A2(pi1068), .ZN(new_n32760_));
  OAI21_X1   g30324(.A1(new_n6626_), .A2(new_n32587_), .B(new_n32760_), .ZN(po0541));
  NAND2_X1   g30325(.A1(new_n32587_), .A2(pi1042), .ZN(new_n32762_));
  OAI21_X1   g30326(.A1(new_n6597_), .A2(new_n32587_), .B(new_n32762_), .ZN(po0542));
  NAND2_X1   g30327(.A1(new_n32587_), .A2(pi1059), .ZN(new_n32764_));
  OAI21_X1   g30328(.A1(new_n6557_), .A2(new_n32587_), .B(new_n32764_), .ZN(po0543));
  NAND2_X1   g30329(.A1(new_n32646_), .A2(pi0387), .ZN(new_n32766_));
  OAI21_X1   g30330(.A1(new_n32490_), .A2(new_n32646_), .B(new_n32766_), .ZN(po0544));
  NAND2_X1   g30331(.A1(new_n32646_), .A2(pi0388), .ZN(new_n32768_));
  OAI21_X1   g30332(.A1(new_n32493_), .A2(new_n32646_), .B(new_n32768_), .ZN(po0545));
  NAND2_X1   g30333(.A1(new_n32646_), .A2(pi0389), .ZN(new_n32770_));
  OAI21_X1   g30334(.A1(new_n31338_), .A2(new_n32646_), .B(new_n32770_), .ZN(po0546));
  INV_X1     g30335(.I(pi0390), .ZN(new_n32772_));
  NAND2_X1   g30336(.A1(new_n32591_), .A2(pi1049), .ZN(new_n32773_));
  OAI21_X1   g30337(.A1(new_n32772_), .A2(new_n32591_), .B(new_n32773_), .ZN(po0547));
  NAND2_X1   g30338(.A1(new_n32591_), .A2(pi1062), .ZN(new_n32775_));
  OAI21_X1   g30339(.A1(new_n9865_), .A2(new_n32591_), .B(new_n32775_), .ZN(po0548));
  NAND2_X1   g30340(.A1(new_n32591_), .A2(pi1039), .ZN(new_n32777_));
  OAI21_X1   g30341(.A1(new_n9936_), .A2(new_n32591_), .B(new_n32777_), .ZN(po0549));
  NAND2_X1   g30342(.A1(new_n32591_), .A2(pi1067), .ZN(new_n32779_));
  OAI21_X1   g30343(.A1(new_n7158_), .A2(new_n32591_), .B(new_n32779_), .ZN(po0550));
  INV_X1     g30344(.I(pi0394), .ZN(new_n32781_));
  NAND2_X1   g30345(.A1(new_n32591_), .A2(pi1080), .ZN(new_n32782_));
  OAI21_X1   g30346(.A1(new_n32781_), .A2(new_n32591_), .B(new_n32782_), .ZN(po0551));
  INV_X1     g30347(.I(pi0395), .ZN(new_n32784_));
  NAND2_X1   g30348(.A1(new_n32591_), .A2(pi1055), .ZN(new_n32785_));
  OAI21_X1   g30349(.A1(new_n32784_), .A2(new_n32591_), .B(new_n32785_), .ZN(po0552));
  NAND2_X1   g30350(.A1(new_n32591_), .A2(pi1051), .ZN(new_n32787_));
  OAI21_X1   g30351(.A1(new_n6368_), .A2(new_n32591_), .B(new_n32787_), .ZN(po0553));
  NAND2_X1   g30352(.A1(new_n32591_), .A2(pi1048), .ZN(new_n32789_));
  OAI21_X1   g30353(.A1(new_n9832_), .A2(new_n32591_), .B(new_n32789_), .ZN(po0554));
  INV_X1     g30354(.I(pi0398), .ZN(new_n32791_));
  NAND2_X1   g30355(.A1(new_n32591_), .A2(pi1087), .ZN(new_n32792_));
  OAI21_X1   g30356(.A1(new_n32791_), .A2(new_n32591_), .B(new_n32792_), .ZN(po0555));
  INV_X1     g30357(.I(pi0399), .ZN(new_n32794_));
  NAND2_X1   g30358(.A1(new_n32591_), .A2(pi1047), .ZN(new_n32795_));
  OAI21_X1   g30359(.A1(new_n32794_), .A2(new_n32591_), .B(new_n32795_), .ZN(po0556));
  INV_X1     g30360(.I(pi0400), .ZN(new_n32797_));
  NAND2_X1   g30361(.A1(new_n32591_), .A2(pi1035), .ZN(new_n32798_));
  OAI21_X1   g30362(.A1(new_n32797_), .A2(new_n32591_), .B(new_n32798_), .ZN(po0557));
  INV_X1     g30363(.I(pi0401), .ZN(new_n32800_));
  NAND2_X1   g30364(.A1(new_n32591_), .A2(pi1079), .ZN(new_n32801_));
  OAI21_X1   g30365(.A1(new_n32800_), .A2(new_n32591_), .B(new_n32801_), .ZN(po0558));
  INV_X1     g30366(.I(pi0402), .ZN(new_n32803_));
  NAND2_X1   g30367(.A1(new_n32591_), .A2(pi1078), .ZN(new_n32804_));
  OAI21_X1   g30368(.A1(new_n32803_), .A2(new_n32591_), .B(new_n32804_), .ZN(po0559));
  INV_X1     g30369(.I(pi0403), .ZN(new_n32806_));
  NAND2_X1   g30370(.A1(new_n32591_), .A2(pi1045), .ZN(new_n32807_));
  OAI21_X1   g30371(.A1(new_n32806_), .A2(new_n32591_), .B(new_n32807_), .ZN(po0560));
  NAND2_X1   g30372(.A1(new_n32591_), .A2(pi1084), .ZN(new_n32809_));
  OAI21_X1   g30373(.A1(new_n9829_), .A2(new_n32591_), .B(new_n32809_), .ZN(po0561));
  INV_X1     g30374(.I(pi0405), .ZN(new_n32811_));
  NAND2_X1   g30375(.A1(new_n32591_), .A2(pi1081), .ZN(new_n32812_));
  OAI21_X1   g30376(.A1(new_n32811_), .A2(new_n32591_), .B(new_n32812_), .ZN(po0562));
  INV_X1     g30377(.I(pi0406), .ZN(new_n32814_));
  NAND2_X1   g30378(.A1(new_n32591_), .A2(pi1076), .ZN(new_n32815_));
  OAI21_X1   g30379(.A1(new_n32814_), .A2(new_n32591_), .B(new_n32815_), .ZN(po0563));
  NAND2_X1   g30380(.A1(new_n32591_), .A2(pi1071), .ZN(new_n32817_));
  NAND2_X1   g30381(.A1(new_n32592_), .A2(pi0407), .ZN(new_n32818_));
  NAND2_X1   g30382(.A1(new_n32818_), .A2(new_n32817_), .ZN(po0564));
  NAND2_X1   g30383(.A1(new_n32591_), .A2(pi1068), .ZN(new_n32820_));
  OAI21_X1   g30384(.A1(new_n6370_), .A2(new_n32591_), .B(new_n32820_), .ZN(po0565));
  NAND2_X1   g30385(.A1(new_n32591_), .A2(pi1042), .ZN(new_n32822_));
  NAND2_X1   g30386(.A1(new_n32592_), .A2(pi0409), .ZN(new_n32823_));
  NAND2_X1   g30387(.A1(new_n32823_), .A2(new_n32822_), .ZN(po0566));
  INV_X1     g30388(.I(pi0410), .ZN(new_n32825_));
  NAND2_X1   g30389(.A1(new_n32591_), .A2(pi1059), .ZN(new_n32826_));
  OAI21_X1   g30390(.A1(new_n32825_), .A2(new_n32591_), .B(new_n32826_), .ZN(po0567));
  NAND2_X1   g30391(.A1(new_n32591_), .A2(pi1053), .ZN(new_n32828_));
  OAI21_X1   g30392(.A1(new_n6382_), .A2(new_n32591_), .B(new_n32828_), .ZN(po0568));
  NAND2_X1   g30393(.A1(new_n32592_), .A2(pi0412), .ZN(new_n32830_));
  OAI21_X1   g30394(.A1(new_n32493_), .A2(new_n32592_), .B(new_n32830_), .ZN(po0569));
  NAND2_X1   g30395(.A1(new_n32591_), .A2(pi1036), .ZN(new_n32832_));
  OAI21_X1   g30396(.A1(new_n6358_), .A2(new_n32591_), .B(new_n32832_), .ZN(po0570));
  INV_X1     g30397(.I(pi0414), .ZN(new_n32834_));
  NOR2_X1    g30398(.A1(new_n32580_), .A2(pi0331), .ZN(new_n32835_));
  NAND2_X1   g30399(.A1(new_n32835_), .A2(pi1049), .ZN(new_n32836_));
  OAI21_X1   g30400(.A1(new_n32834_), .A2(new_n32835_), .B(new_n32836_), .ZN(po0571));
  INV_X1     g30401(.I(pi0415), .ZN(new_n32838_));
  NAND2_X1   g30402(.A1(new_n32835_), .A2(pi1062), .ZN(new_n32839_));
  OAI21_X1   g30403(.A1(new_n32838_), .A2(new_n32835_), .B(new_n32839_), .ZN(po0572));
  INV_X1     g30404(.I(pi0416), .ZN(new_n32841_));
  NAND2_X1   g30405(.A1(new_n32835_), .A2(pi1069), .ZN(new_n32842_));
  OAI21_X1   g30406(.A1(new_n32841_), .A2(new_n32835_), .B(new_n32842_), .ZN(po0573));
  NAND2_X1   g30407(.A1(new_n32835_), .A2(pi1039), .ZN(new_n32844_));
  OAI21_X1   g30408(.A1(new_n6289_), .A2(new_n32835_), .B(new_n32844_), .ZN(po0574));
  NAND2_X1   g30409(.A1(new_n32835_), .A2(pi1067), .ZN(new_n32846_));
  OAI21_X1   g30410(.A1(new_n6285_), .A2(new_n32835_), .B(new_n32846_), .ZN(po0575));
  INV_X1     g30411(.I(pi0419), .ZN(new_n32848_));
  NAND2_X1   g30412(.A1(new_n32835_), .A2(pi1080), .ZN(new_n32849_));
  OAI21_X1   g30413(.A1(new_n32848_), .A2(new_n32835_), .B(new_n32849_), .ZN(po0576));
  INV_X1     g30414(.I(pi0420), .ZN(new_n32851_));
  NAND2_X1   g30415(.A1(new_n32835_), .A2(pi1055), .ZN(new_n32852_));
  OAI21_X1   g30416(.A1(new_n32851_), .A2(new_n32835_), .B(new_n32852_), .ZN(po0577));
  INV_X1     g30417(.I(pi0421), .ZN(new_n32854_));
  NAND2_X1   g30418(.A1(new_n32835_), .A2(pi1051), .ZN(new_n32855_));
  OAI21_X1   g30419(.A1(new_n32854_), .A2(new_n32835_), .B(new_n32855_), .ZN(po0578));
  INV_X1     g30420(.I(pi0422), .ZN(new_n32857_));
  NAND2_X1   g30421(.A1(new_n32835_), .A2(pi1048), .ZN(new_n32858_));
  OAI21_X1   g30422(.A1(new_n32857_), .A2(new_n32835_), .B(new_n32858_), .ZN(po0579));
  NAND2_X1   g30423(.A1(new_n32835_), .A2(pi1087), .ZN(new_n32860_));
  OAI21_X1   g30424(.A1(new_n6278_), .A2(new_n32835_), .B(new_n32860_), .ZN(po0580));
  INV_X1     g30425(.I(pi0424), .ZN(new_n32862_));
  NAND2_X1   g30426(.A1(new_n32835_), .A2(pi1047), .ZN(new_n32863_));
  OAI21_X1   g30427(.A1(new_n32862_), .A2(new_n32835_), .B(new_n32863_), .ZN(po0581));
  INV_X1     g30428(.I(pi0425), .ZN(new_n32865_));
  NAND2_X1   g30429(.A1(new_n32835_), .A2(pi1035), .ZN(new_n32866_));
  OAI21_X1   g30430(.A1(new_n32865_), .A2(new_n32835_), .B(new_n32866_), .ZN(po0582));
  INV_X1     g30431(.I(pi0426), .ZN(new_n32868_));
  NAND2_X1   g30432(.A1(new_n32835_), .A2(pi1079), .ZN(new_n32869_));
  OAI21_X1   g30433(.A1(new_n32868_), .A2(new_n32835_), .B(new_n32869_), .ZN(po0583));
  INV_X1     g30434(.I(pi0427), .ZN(new_n32871_));
  NAND2_X1   g30435(.A1(new_n32835_), .A2(pi1078), .ZN(new_n32872_));
  OAI21_X1   g30436(.A1(new_n32871_), .A2(new_n32835_), .B(new_n32872_), .ZN(po0584));
  NAND2_X1   g30437(.A1(new_n32835_), .A2(pi1045), .ZN(new_n32874_));
  OAI21_X1   g30438(.A1(new_n6333_), .A2(new_n32835_), .B(new_n32874_), .ZN(po0585));
  NAND2_X1   g30439(.A1(new_n32835_), .A2(pi1084), .ZN(new_n32876_));
  OAI21_X1   g30440(.A1(new_n10059_), .A2(new_n32835_), .B(new_n32876_), .ZN(po0586));
  NAND2_X1   g30441(.A1(new_n32835_), .A2(pi1076), .ZN(new_n32878_));
  OAI21_X1   g30442(.A1(new_n6335_), .A2(new_n32835_), .B(new_n32878_), .ZN(po0587));
  INV_X1     g30443(.I(pi0431), .ZN(new_n32880_));
  NAND2_X1   g30444(.A1(new_n32835_), .A2(pi1071), .ZN(new_n32881_));
  OAI21_X1   g30445(.A1(new_n32880_), .A2(new_n32835_), .B(new_n32881_), .ZN(po0588));
  INV_X1     g30446(.I(pi0432), .ZN(new_n32883_));
  NAND2_X1   g30447(.A1(new_n32835_), .A2(pi1068), .ZN(new_n32884_));
  OAI21_X1   g30448(.A1(new_n32883_), .A2(new_n32835_), .B(new_n32884_), .ZN(po0589));
  NAND2_X1   g30449(.A1(new_n32835_), .A2(pi1042), .ZN(new_n32886_));
  OAI21_X1   g30450(.A1(new_n6327_), .A2(new_n32835_), .B(new_n32886_), .ZN(po0590));
  NAND2_X1   g30451(.A1(new_n32835_), .A2(pi1059), .ZN(new_n32888_));
  OAI21_X1   g30452(.A1(new_n6309_), .A2(new_n32835_), .B(new_n32888_), .ZN(po0591));
  NAND2_X1   g30453(.A1(new_n32835_), .A2(pi1053), .ZN(new_n32890_));
  OAI21_X1   g30454(.A1(new_n10045_), .A2(new_n32835_), .B(new_n32890_), .ZN(po0592));
  NAND2_X1   g30455(.A1(new_n32835_), .A2(pi1037), .ZN(new_n32892_));
  OAI21_X1   g30456(.A1(new_n6306_), .A2(new_n32835_), .B(new_n32892_), .ZN(po0593));
  NAND2_X1   g30457(.A1(new_n32835_), .A2(pi1070), .ZN(new_n32894_));
  OAI21_X1   g30458(.A1(new_n6286_), .A2(new_n32835_), .B(new_n32894_), .ZN(po0594));
  NAND2_X1   g30459(.A1(new_n32835_), .A2(pi1036), .ZN(new_n32896_));
  OAI21_X1   g30460(.A1(new_n6297_), .A2(new_n32835_), .B(new_n32896_), .ZN(po0595));
  INV_X1     g30461(.I(pi1057), .ZN(new_n32898_));
  NAND2_X1   g30462(.A1(new_n32646_), .A2(pi0439), .ZN(new_n32899_));
  OAI21_X1   g30463(.A1(new_n32898_), .A2(new_n32646_), .B(new_n32899_), .ZN(po0596));
  NAND2_X1   g30464(.A1(new_n32587_), .A2(pi1043), .ZN(new_n32901_));
  OAI21_X1   g30465(.A1(new_n6622_), .A2(new_n32587_), .B(new_n32901_), .ZN(po0597));
  NAND2_X1   g30466(.A1(new_n32581_), .A2(pi1044), .ZN(new_n32903_));
  OAI21_X1   g30467(.A1(new_n6518_), .A2(new_n32581_), .B(new_n32903_), .ZN(po0598));
  NAND2_X1   g30468(.A1(new_n32587_), .A2(pi1058), .ZN(new_n32905_));
  OAI21_X1   g30469(.A1(new_n6623_), .A2(new_n32587_), .B(new_n32905_), .ZN(po0599));
  NAND2_X1   g30470(.A1(new_n32835_), .A2(pi1044), .ZN(new_n32907_));
  OAI21_X1   g30471(.A1(new_n10050_), .A2(new_n32835_), .B(new_n32907_), .ZN(po0600));
  NAND2_X1   g30472(.A1(new_n32835_), .A2(pi1072), .ZN(new_n32909_));
  OAI21_X1   g30473(.A1(new_n6891_), .A2(new_n32835_), .B(new_n32909_), .ZN(po0601));
  NAND2_X1   g30474(.A1(new_n32835_), .A2(pi1081), .ZN(new_n32911_));
  OAI21_X1   g30475(.A1(new_n6859_), .A2(new_n32835_), .B(new_n32911_), .ZN(po0602));
  NAND2_X1   g30476(.A1(new_n32835_), .A2(pi1086), .ZN(new_n32913_));
  OAI21_X1   g30477(.A1(new_n6311_), .A2(new_n32835_), .B(new_n32913_), .ZN(po0603));
  NAND2_X1   g30478(.A1(new_n32646_), .A2(pi0447), .ZN(new_n32915_));
  OAI21_X1   g30479(.A1(new_n32614_), .A2(new_n32646_), .B(new_n32915_), .ZN(po0604));
  NAND2_X1   g30480(.A1(new_n32835_), .A2(pi1074), .ZN(new_n32917_));
  OAI21_X1   g30481(.A1(new_n9760_), .A2(new_n32835_), .B(new_n32917_), .ZN(po0605));
  NAND2_X1   g30482(.A1(new_n32835_), .A2(pi1057), .ZN(new_n32919_));
  OAI21_X1   g30483(.A1(new_n6324_), .A2(new_n32835_), .B(new_n32919_), .ZN(po0606));
  NAND2_X1   g30484(.A1(new_n32615_), .A2(pi0450), .ZN(new_n32921_));
  OAI21_X1   g30485(.A1(new_n31338_), .A2(new_n32615_), .B(new_n32921_), .ZN(po0607));
  NAND2_X1   g30486(.A1(new_n32835_), .A2(pi1063), .ZN(new_n32923_));
  OAI21_X1   g30487(.A1(new_n6322_), .A2(new_n32835_), .B(new_n32923_), .ZN(po0608));
  NAND2_X1   g30488(.A1(new_n32581_), .A2(pi1053), .ZN(new_n32925_));
  OAI21_X1   g30489(.A1(new_n6487_), .A2(new_n32581_), .B(new_n32925_), .ZN(po0609));
  INV_X1     g30490(.I(pi0453), .ZN(new_n32927_));
  NAND2_X1   g30491(.A1(new_n32835_), .A2(pi1040), .ZN(new_n32928_));
  OAI21_X1   g30492(.A1(new_n32927_), .A2(new_n32835_), .B(new_n32928_), .ZN(po0610));
  INV_X1     g30493(.I(pi0454), .ZN(new_n32930_));
  NAND2_X1   g30494(.A1(new_n32835_), .A2(pi1043), .ZN(new_n32931_));
  OAI21_X1   g30495(.A1(new_n32930_), .A2(new_n32835_), .B(new_n32931_), .ZN(po0611));
  NAND2_X1   g30496(.A1(new_n32581_), .A2(pi1037), .ZN(new_n32933_));
  OAI21_X1   g30497(.A1(new_n6488_), .A2(new_n32581_), .B(new_n32933_), .ZN(po0612));
  NAND2_X1   g30498(.A1(new_n32591_), .A2(pi1044), .ZN(new_n32935_));
  OAI21_X1   g30499(.A1(new_n6386_), .A2(new_n32591_), .B(new_n32935_), .ZN(po0613));
  INV_X1     g30500(.I(pi0821), .ZN(new_n32937_));
  INV_X1     g30501(.I(pi0815), .ZN(new_n32938_));
  INV_X1     g30502(.I(pi0804), .ZN(new_n32939_));
  INV_X1     g30503(.I(pi0810), .ZN(new_n32940_));
  AOI21_X1   g30504(.A1(pi0600), .A2(new_n32940_), .B(new_n32939_), .ZN(new_n32941_));
  NAND3_X1   g30505(.A1(pi0594), .A2(pi0600), .A3(pi0990), .ZN(new_n32942_));
  INV_X1     g30506(.I(new_n32942_), .ZN(new_n32943_));
  NAND3_X1   g30507(.A1(new_n32941_), .A2(new_n32943_), .A3(new_n32938_), .ZN(new_n32944_));
  NOR2_X1    g30508(.A1(pi0804), .A2(pi0810), .ZN(new_n32945_));
  OAI21_X1   g30509(.A1(new_n32945_), .A2(pi0601), .B(new_n32938_), .ZN(new_n32946_));
  NOR2_X1    g30510(.A1(new_n32946_), .A2(new_n32941_), .ZN(new_n32947_));
  INV_X1     g30511(.I(pi0595), .ZN(new_n32948_));
  NAND2_X1   g30512(.A1(new_n32945_), .A2(new_n32948_), .ZN(new_n32949_));
  INV_X1     g30513(.I(pi0596), .ZN(new_n32950_));
  NOR2_X1    g30514(.A1(new_n32940_), .A2(pi0599), .ZN(new_n32951_));
  OAI21_X1   g30515(.A1(new_n32951_), .A2(new_n32950_), .B(pi0804), .ZN(new_n32952_));
  NAND3_X1   g30516(.A1(new_n32952_), .A2(pi0595), .A3(pi0815), .ZN(new_n32953_));
  NAND4_X1   g30517(.A1(pi0594), .A2(pi0597), .A3(pi0600), .A4(pi0601), .ZN(new_n32954_));
  AOI21_X1   g30518(.A1(new_n32953_), .A2(new_n32949_), .B(new_n32954_), .ZN(new_n32955_));
  OAI21_X1   g30519(.A1(new_n32955_), .A2(new_n32947_), .B(pi0605), .ZN(new_n32956_));
  AOI21_X1   g30520(.A1(new_n32956_), .A2(new_n32944_), .B(new_n32937_), .ZN(po0614));
  NAND2_X1   g30521(.A1(new_n32581_), .A2(pi1072), .ZN(new_n32958_));
  OAI21_X1   g30522(.A1(new_n7136_), .A2(new_n32581_), .B(new_n32958_), .ZN(po0615));
  INV_X1     g30523(.I(pi0459), .ZN(new_n32960_));
  NAND2_X1   g30524(.A1(new_n32835_), .A2(pi1058), .ZN(new_n32961_));
  OAI21_X1   g30525(.A1(new_n32960_), .A2(new_n32835_), .B(new_n32961_), .ZN(po0616));
  NAND2_X1   g30526(.A1(new_n32581_), .A2(pi1086), .ZN(new_n32963_));
  OAI21_X1   g30527(.A1(new_n6470_), .A2(new_n32581_), .B(new_n32963_), .ZN(po0617));
  NAND2_X1   g30528(.A1(new_n32615_), .A2(pi0461), .ZN(new_n32965_));
  OAI21_X1   g30529(.A1(new_n32898_), .A2(new_n32615_), .B(new_n32965_), .ZN(po0618));
  NAND2_X1   g30530(.A1(new_n32581_), .A2(pi1074), .ZN(new_n32967_));
  OAI21_X1   g30531(.A1(new_n6540_), .A2(new_n32581_), .B(new_n32967_), .ZN(po0619));
  NAND2_X1   g30532(.A1(new_n32591_), .A2(pi1070), .ZN(new_n32969_));
  OAI21_X1   g30533(.A1(new_n6356_), .A2(new_n32591_), .B(new_n32969_), .ZN(po0620));
  INV_X1     g30534(.I(pi0464), .ZN(new_n32971_));
  NAND2_X1   g30535(.A1(new_n32835_), .A2(pi1065), .ZN(new_n32972_));
  OAI21_X1   g30536(.A1(new_n32971_), .A2(new_n32835_), .B(new_n32972_), .ZN(po0621));
  NOR2_X1    g30537(.A1(new_n9190_), .A2(new_n9192_), .ZN(new_n32974_));
  NOR2_X1    g30538(.A1(new_n5270_), .A2(new_n5216_), .ZN(new_n32975_));
  INV_X1     g30539(.I(new_n32975_), .ZN(new_n32976_));
  NOR2_X1    g30540(.A1(new_n32976_), .A2(pi1157), .ZN(new_n32977_));
  NOR2_X1    g30541(.A1(new_n32975_), .A2(pi0926), .ZN(new_n32978_));
  OAI22_X1   g30542(.A1(new_n32977_), .A2(new_n32978_), .B1(pi0243), .B2(new_n32974_), .ZN(new_n32979_));
  INV_X1     g30543(.I(new_n32974_), .ZN(new_n32980_));
  OAI21_X1   g30544(.A1(new_n32980_), .A2(pi1157), .B(new_n29935_), .ZN(new_n32981_));
  NOR3_X1    g30545(.A1(pi0222), .A2(pi0223), .A3(pi0299), .ZN(new_n32982_));
  AOI21_X1   g30546(.A1(pi0299), .A2(new_n2558_), .B(new_n32982_), .ZN(new_n32983_));
  INV_X1     g30547(.I(new_n32983_), .ZN(new_n32984_));
  INV_X1     g30548(.I(pi0926), .ZN(new_n32985_));
  AOI21_X1   g30549(.A1(new_n3303_), .A2(new_n5113_), .B(new_n3337_), .ZN(new_n32986_));
  NOR4_X1    g30550(.A1(new_n32986_), .A2(pi0243), .A3(new_n32985_), .A4(new_n12965_), .ZN(new_n32987_));
  AOI21_X1   g30551(.A1(new_n32981_), .A2(new_n32984_), .B(new_n32987_), .ZN(new_n32988_));
  NAND2_X1   g30552(.A1(new_n32979_), .A2(new_n32988_), .ZN(new_n32989_));
  NAND2_X1   g30553(.A1(new_n32525_), .A2(new_n29935_), .ZN(new_n32990_));
  INV_X1     g30554(.I(new_n5200_), .ZN(new_n32991_));
  INV_X1     g30555(.I(new_n32526_), .ZN(new_n32992_));
  OAI22_X1   g30556(.A1(new_n32992_), .A2(new_n32985_), .B1(new_n12965_), .B2(new_n32991_), .ZN(new_n32993_));
  NOR2_X1    g30557(.A1(new_n32993_), .A2(new_n6643_), .ZN(new_n32994_));
  AOI22_X1   g30558(.A1(new_n32989_), .A2(new_n6643_), .B1(new_n32990_), .B2(new_n32994_), .ZN(po0622));
  INV_X1     g30559(.I(pi0943), .ZN(new_n32996_));
  NOR2_X1    g30560(.A1(new_n32974_), .A2(po1038), .ZN(new_n32997_));
  AOI21_X1   g30561(.A1(po1038), .A2(new_n32525_), .B(new_n32997_), .ZN(new_n32998_));
  NAND2_X1   g30562(.A1(new_n32998_), .A2(new_n32996_), .ZN(new_n32999_));
  NAND2_X1   g30563(.A1(new_n32560_), .A2(pi0943), .ZN(new_n33000_));
  AOI21_X1   g30564(.A1(new_n33000_), .A2(new_n32999_), .B(pi1151), .ZN(new_n33001_));
  NAND2_X1   g30565(.A1(new_n32530_), .A2(new_n32998_), .ZN(new_n33002_));
  NOR2_X1    g30566(.A1(new_n33002_), .A2(pi0943), .ZN(new_n33003_));
  OAI21_X1   g30567(.A1(new_n2644_), .A2(new_n25319_), .B(new_n32518_), .ZN(new_n33004_));
  NAND2_X1   g30568(.A1(new_n33004_), .A2(pi0943), .ZN(new_n33005_));
  NOR2_X1    g30569(.A1(po1038), .A2(new_n32983_), .ZN(new_n33006_));
  AOI21_X1   g30570(.A1(new_n2558_), .A2(po1038), .B(new_n33006_), .ZN(new_n33007_));
  OAI22_X1   g30571(.A1(new_n33005_), .A2(new_n29035_), .B1(pi0275), .B2(new_n33007_), .ZN(new_n33008_));
  NOR3_X1    g30572(.A1(new_n33008_), .A2(new_n33001_), .A3(new_n33003_), .ZN(po0623));
  INV_X1     g30573(.I(new_n31004_), .ZN(new_n33010_));
  NOR4_X1    g30574(.A1(new_n33010_), .A2(new_n2818_), .A3(pi0287), .A4(new_n9148_), .ZN(new_n33011_));
  NAND2_X1   g30575(.A1(po0950), .A2(new_n33011_), .ZN(new_n33012_));
  INV_X1     g30576(.I(new_n33011_), .ZN(new_n33013_));
  NOR3_X1    g30577(.A1(new_n8254_), .A2(new_n7293_), .A3(new_n13010_), .ZN(new_n33014_));
  NAND2_X1   g30578(.A1(new_n10486_), .A2(new_n2501_), .ZN(new_n33015_));
  NAND3_X1   g30579(.A1(new_n33015_), .A2(new_n13008_), .A3(new_n33014_), .ZN(new_n33016_));
  OAI21_X1   g30580(.A1(new_n6258_), .A2(new_n33013_), .B(new_n33016_), .ZN(new_n33017_));
  NOR2_X1    g30581(.A1(new_n33016_), .A2(new_n33013_), .ZN(new_n33018_));
  NAND2_X1   g30582(.A1(new_n33018_), .A2(new_n6259_), .ZN(new_n33019_));
  AOI21_X1   g30583(.A1(new_n33019_), .A2(new_n33017_), .B(new_n3041_), .ZN(new_n33020_));
  NAND2_X1   g30584(.A1(new_n33011_), .A2(new_n5331_), .ZN(new_n33021_));
  AOI22_X1   g30585(.A1(new_n33018_), .A2(new_n5331_), .B1(new_n33016_), .B2(new_n33021_), .ZN(new_n33022_));
  NOR2_X1    g30586(.A1(new_n33022_), .A2(pi1093), .ZN(new_n33023_));
  OAI21_X1   g30587(.A1(new_n33023_), .A2(new_n33020_), .B(new_n3022_), .ZN(new_n33024_));
  INV_X1     g30588(.I(new_n6781_), .ZN(new_n33025_));
  INV_X1     g30589(.I(new_n33018_), .ZN(new_n33026_));
  NAND2_X1   g30590(.A1(new_n33016_), .A2(new_n33013_), .ZN(new_n33027_));
  AOI21_X1   g30591(.A1(new_n33026_), .A2(new_n33027_), .B(new_n33025_), .ZN(new_n33028_));
  NOR2_X1    g30592(.A1(new_n33022_), .A2(new_n6781_), .ZN(new_n33029_));
  OAI21_X1   g30593(.A1(new_n33029_), .A2(new_n33028_), .B(pi1091), .ZN(new_n33030_));
  NAND2_X1   g30594(.A1(new_n33024_), .A2(new_n33030_), .ZN(new_n33031_));
  NOR2_X1    g30595(.A1(new_n2659_), .A2(new_n32573_), .ZN(new_n33032_));
  AOI22_X1   g30596(.A1(new_n33031_), .A2(new_n33032_), .B1(new_n8260_), .B2(new_n33012_), .ZN(po0624));
  NOR4_X1    g30597(.A1(new_n7335_), .A2(new_n3265_), .A3(pi0039), .A4(new_n8265_), .ZN(new_n33034_));
  OAI22_X1   g30598(.A1(new_n33034_), .A2(new_n10534_), .B1(new_n8281_), .B2(new_n9151_), .ZN(po0625));
  NOR2_X1    g30599(.A1(new_n32976_), .A2(pi1156), .ZN(new_n33036_));
  NOR2_X1    g30600(.A1(new_n32975_), .A2(pi0942), .ZN(new_n33037_));
  OAI22_X1   g30601(.A1(new_n33036_), .A2(new_n33037_), .B1(pi0263), .B2(new_n32974_), .ZN(new_n33038_));
  OAI21_X1   g30602(.A1(new_n32980_), .A2(pi1156), .B(new_n31416_), .ZN(new_n33039_));
  INV_X1     g30603(.I(pi0942), .ZN(new_n33040_));
  NOR4_X1    g30604(.A1(new_n32986_), .A2(pi0263), .A3(new_n33040_), .A4(new_n12742_), .ZN(new_n33041_));
  AOI21_X1   g30605(.A1(new_n33039_), .A2(new_n32984_), .B(new_n33041_), .ZN(new_n33042_));
  NAND2_X1   g30606(.A1(new_n33038_), .A2(new_n33042_), .ZN(new_n33043_));
  NAND2_X1   g30607(.A1(new_n32525_), .A2(new_n31416_), .ZN(new_n33044_));
  OAI22_X1   g30608(.A1(new_n32992_), .A2(new_n33040_), .B1(new_n12742_), .B2(new_n32991_), .ZN(new_n33045_));
  NOR2_X1    g30609(.A1(new_n33045_), .A2(new_n6643_), .ZN(new_n33046_));
  AOI22_X1   g30610(.A1(new_n33043_), .A2(new_n6643_), .B1(new_n33044_), .B2(new_n33046_), .ZN(po0626));
  NOR2_X1    g30611(.A1(new_n32976_), .A2(pi1155), .ZN(new_n33048_));
  NOR2_X1    g30612(.A1(new_n32975_), .A2(pi0925), .ZN(new_n33049_));
  OAI22_X1   g30613(.A1(new_n33048_), .A2(new_n33049_), .B1(new_n29990_), .B2(new_n32974_), .ZN(new_n33050_));
  OAI21_X1   g30614(.A1(new_n32980_), .A2(pi1155), .B(pi0267), .ZN(new_n33051_));
  INV_X1     g30615(.I(pi0925), .ZN(new_n33052_));
  NOR4_X1    g30616(.A1(new_n32986_), .A2(new_n29990_), .A3(new_n33052_), .A4(new_n12770_), .ZN(new_n33053_));
  AOI21_X1   g30617(.A1(new_n33051_), .A2(new_n32984_), .B(new_n33053_), .ZN(new_n33054_));
  NAND2_X1   g30618(.A1(new_n33050_), .A2(new_n33054_), .ZN(new_n33055_));
  NAND2_X1   g30619(.A1(new_n32525_), .A2(pi0267), .ZN(new_n33056_));
  OAI22_X1   g30620(.A1(new_n32992_), .A2(new_n33052_), .B1(new_n12770_), .B2(new_n32991_), .ZN(new_n33057_));
  NOR2_X1    g30621(.A1(new_n33057_), .A2(new_n6643_), .ZN(new_n33058_));
  AOI22_X1   g30622(.A1(new_n33055_), .A2(new_n6643_), .B1(new_n33056_), .B2(new_n33058_), .ZN(po0627));
  NOR2_X1    g30623(.A1(new_n32976_), .A2(pi1153), .ZN(new_n33060_));
  NOR2_X1    g30624(.A1(new_n32975_), .A2(pi0941), .ZN(new_n33061_));
  OAI22_X1   g30625(.A1(new_n33060_), .A2(new_n33061_), .B1(new_n29991_), .B2(new_n32974_), .ZN(new_n33062_));
  OAI21_X1   g30626(.A1(new_n32980_), .A2(pi1153), .B(pi0253), .ZN(new_n33063_));
  INV_X1     g30627(.I(pi0941), .ZN(new_n33064_));
  NOR4_X1    g30628(.A1(new_n32986_), .A2(new_n29991_), .A3(new_n33064_), .A4(new_n12841_), .ZN(new_n33065_));
  AOI21_X1   g30629(.A1(new_n33063_), .A2(new_n32984_), .B(new_n33065_), .ZN(new_n33066_));
  NAND2_X1   g30630(.A1(new_n33062_), .A2(new_n33066_), .ZN(new_n33067_));
  NAND2_X1   g30631(.A1(new_n32525_), .A2(pi0253), .ZN(new_n33068_));
  OAI22_X1   g30632(.A1(new_n32992_), .A2(new_n33064_), .B1(new_n12841_), .B2(new_n32991_), .ZN(new_n33069_));
  NOR2_X1    g30633(.A1(new_n33069_), .A2(new_n6643_), .ZN(new_n33070_));
  AOI22_X1   g30634(.A1(new_n33067_), .A2(new_n6643_), .B1(new_n33068_), .B2(new_n33070_), .ZN(po0628));
  NOR2_X1    g30635(.A1(new_n32976_), .A2(pi1154), .ZN(new_n33072_));
  NOR2_X1    g30636(.A1(new_n32975_), .A2(pi0923), .ZN(new_n33073_));
  OAI22_X1   g30637(.A1(new_n33072_), .A2(new_n33073_), .B1(new_n29992_), .B2(new_n32974_), .ZN(new_n33074_));
  OAI21_X1   g30638(.A1(new_n32980_), .A2(pi1154), .B(pi0254), .ZN(new_n33075_));
  INV_X1     g30639(.I(pi0923), .ZN(new_n33076_));
  NOR4_X1    g30640(.A1(new_n32986_), .A2(new_n29992_), .A3(new_n33076_), .A4(new_n12785_), .ZN(new_n33077_));
  AOI21_X1   g30641(.A1(new_n33075_), .A2(new_n32984_), .B(new_n33077_), .ZN(new_n33078_));
  NAND2_X1   g30642(.A1(new_n33074_), .A2(new_n33078_), .ZN(new_n33079_));
  NAND2_X1   g30643(.A1(new_n32525_), .A2(pi0254), .ZN(new_n33080_));
  OAI22_X1   g30644(.A1(new_n32992_), .A2(new_n33076_), .B1(new_n12785_), .B2(new_n32991_), .ZN(new_n33081_));
  NOR2_X1    g30645(.A1(new_n33081_), .A2(new_n6643_), .ZN(new_n33082_));
  AOI22_X1   g30646(.A1(new_n33079_), .A2(new_n6643_), .B1(new_n33080_), .B2(new_n33082_), .ZN(po0629));
  INV_X1     g30647(.I(pi0922), .ZN(new_n33084_));
  NAND2_X1   g30648(.A1(new_n32998_), .A2(new_n33084_), .ZN(new_n33085_));
  NAND2_X1   g30649(.A1(new_n32560_), .A2(pi0922), .ZN(new_n33086_));
  AOI21_X1   g30650(.A1(new_n33086_), .A2(new_n33085_), .B(pi1152), .ZN(new_n33087_));
  NOR2_X1    g30651(.A1(new_n33002_), .A2(pi0922), .ZN(new_n33088_));
  NAND2_X1   g30652(.A1(new_n33004_), .A2(pi0922), .ZN(new_n33089_));
  OAI22_X1   g30653(.A1(new_n33089_), .A2(new_n28422_), .B1(pi0268), .B2(new_n33007_), .ZN(new_n33090_));
  NOR3_X1    g30654(.A1(new_n33090_), .A2(new_n33087_), .A3(new_n33088_), .ZN(po0630));
  INV_X1     g30655(.I(pi0931), .ZN(new_n33092_));
  NAND2_X1   g30656(.A1(new_n32998_), .A2(new_n33092_), .ZN(new_n33093_));
  NAND2_X1   g30657(.A1(new_n32560_), .A2(pi0931), .ZN(new_n33094_));
  AOI21_X1   g30658(.A1(new_n33094_), .A2(new_n33093_), .B(pi1150), .ZN(new_n33095_));
  NOR2_X1    g30659(.A1(new_n33002_), .A2(pi0931), .ZN(new_n33096_));
  NAND2_X1   g30660(.A1(new_n33004_), .A2(pi0931), .ZN(new_n33097_));
  OAI22_X1   g30661(.A1(new_n33097_), .A2(new_n29650_), .B1(pi0272), .B2(new_n33007_), .ZN(new_n33098_));
  NOR3_X1    g30662(.A1(new_n33098_), .A2(new_n33095_), .A3(new_n33096_), .ZN(po0631));
  INV_X1     g30663(.I(pi0936), .ZN(new_n33100_));
  NAND2_X1   g30664(.A1(new_n32998_), .A2(new_n33100_), .ZN(new_n33101_));
  NAND2_X1   g30665(.A1(new_n32560_), .A2(pi0936), .ZN(new_n33102_));
  AOI21_X1   g30666(.A1(new_n33102_), .A2(new_n33101_), .B(pi1149), .ZN(new_n33103_));
  NOR2_X1    g30667(.A1(new_n33002_), .A2(pi0936), .ZN(new_n33104_));
  NAND2_X1   g30668(.A1(new_n33004_), .A2(pi0936), .ZN(new_n33105_));
  OAI22_X1   g30669(.A1(new_n33105_), .A2(new_n29297_), .B1(pi0283), .B2(new_n33007_), .ZN(new_n33106_));
  NOR3_X1    g30670(.A1(new_n33106_), .A2(new_n33103_), .A3(new_n33104_), .ZN(po0632));
  NOR4_X1    g30671(.A1(new_n8980_), .A2(new_n7312_), .A3(new_n9217_), .A4(new_n9220_), .ZN(new_n33108_));
  NOR3_X1    g30672(.A1(new_n10326_), .A2(new_n8246_), .A3(new_n9221_), .ZN(new_n33109_));
  OAI21_X1   g30673(.A1(new_n33109_), .A2(new_n33108_), .B(new_n2611_), .ZN(new_n33110_));
  NOR4_X1    g30674(.A1(new_n33110_), .A2(new_n2475_), .A3(new_n8254_), .A4(new_n10281_), .ZN(new_n33111_));
  NOR2_X1    g30675(.A1(new_n9221_), .A2(new_n2962_), .ZN(new_n33112_));
  NOR2_X1    g30676(.A1(new_n33111_), .A2(new_n33112_), .ZN(new_n33113_));
  NAND2_X1   g30677(.A1(po1038), .A2(pi0071), .ZN(new_n33114_));
  OAI22_X1   g30678(.A1(new_n33113_), .A2(po1038), .B1(new_n9219_), .B2(new_n33114_), .ZN(po0633));
  NAND2_X1   g30679(.A1(new_n32569_), .A2(new_n32570_), .ZN(po0634));
  NOR2_X1    g30680(.A1(new_n31992_), .A2(new_n2962_), .ZN(po0635));
  INV_X1     g30681(.I(pi0481), .ZN(new_n33118_));
  NAND2_X1   g30682(.A1(new_n25330_), .A2(pi0248), .ZN(new_n33119_));
  OAI21_X1   g30683(.A1(new_n33118_), .A2(new_n25330_), .B(new_n33119_), .ZN(po0638));
  INV_X1     g30684(.I(new_n25467_), .ZN(new_n33121_));
  NAND2_X1   g30685(.A1(new_n33121_), .A2(pi0482), .ZN(new_n33122_));
  OAI21_X1   g30686(.A1(new_n3865_), .A2(new_n33121_), .B(new_n33122_), .ZN(po0639));
  INV_X1     g30687(.I(pi0483), .ZN(new_n33124_));
  NAND2_X1   g30688(.A1(new_n25554_), .A2(pi0242), .ZN(new_n33125_));
  OAI21_X1   g30689(.A1(new_n33124_), .A2(new_n25554_), .B(new_n33125_), .ZN(po0640));
  INV_X1     g30690(.I(new_n25554_), .ZN(new_n33127_));
  NAND2_X1   g30691(.A1(new_n33127_), .A2(pi0484), .ZN(new_n33128_));
  OAI21_X1   g30692(.A1(new_n3865_), .A2(new_n33127_), .B(new_n33128_), .ZN(po0641));
  INV_X1     g30693(.I(pi0485), .ZN(new_n33130_));
  NAND2_X1   g30694(.A1(new_n26388_), .A2(pi0234), .ZN(new_n33131_));
  OAI21_X1   g30695(.A1(new_n33130_), .A2(new_n26388_), .B(new_n33131_), .ZN(po0642));
  INV_X1     g30696(.I(pi0486), .ZN(new_n33133_));
  NAND2_X1   g30697(.A1(new_n26388_), .A2(pi0244), .ZN(new_n33134_));
  OAI21_X1   g30698(.A1(new_n33133_), .A2(new_n26388_), .B(new_n33134_), .ZN(po0643));
  INV_X1     g30699(.I(pi0487), .ZN(new_n33136_));
  NAND2_X1   g30700(.A1(new_n25330_), .A2(pi0246), .ZN(new_n33137_));
  OAI21_X1   g30701(.A1(new_n33136_), .A2(new_n25330_), .B(new_n33137_), .ZN(po0644));
  NAND2_X1   g30702(.A1(new_n25330_), .A2(pi0239), .ZN(new_n33139_));
  OAI21_X1   g30703(.A1(pi0488), .A2(new_n25330_), .B(new_n33139_), .ZN(po0645));
  INV_X1     g30704(.I(pi0489), .ZN(new_n33141_));
  NAND2_X1   g30705(.A1(new_n26388_), .A2(pi0242), .ZN(new_n33142_));
  OAI21_X1   g30706(.A1(new_n33141_), .A2(new_n26388_), .B(new_n33142_), .ZN(po0646));
  NAND2_X1   g30707(.A1(new_n33127_), .A2(pi0490), .ZN(new_n33144_));
  OAI21_X1   g30708(.A1(new_n3948_), .A2(new_n33127_), .B(new_n33144_), .ZN(po0647));
  NAND2_X1   g30709(.A1(new_n33127_), .A2(pi0491), .ZN(new_n33146_));
  OAI21_X1   g30710(.A1(new_n3625_), .A2(new_n33127_), .B(new_n33146_), .ZN(po0648));
  INV_X1     g30711(.I(pi0492), .ZN(new_n33148_));
  NAND2_X1   g30712(.A1(new_n25554_), .A2(pi0240), .ZN(new_n33149_));
  OAI21_X1   g30713(.A1(new_n33148_), .A2(new_n25554_), .B(new_n33149_), .ZN(po0649));
  INV_X1     g30714(.I(pi0493), .ZN(new_n33151_));
  NAND2_X1   g30715(.A1(new_n25554_), .A2(pi0244), .ZN(new_n33152_));
  OAI21_X1   g30716(.A1(new_n33151_), .A2(new_n25554_), .B(new_n33152_), .ZN(po0650));
  NAND2_X1   g30717(.A1(new_n25554_), .A2(pi0239), .ZN(new_n33154_));
  OAI21_X1   g30718(.A1(pi0494), .A2(new_n25554_), .B(new_n33154_), .ZN(po0651));
  INV_X1     g30719(.I(pi0495), .ZN(new_n33156_));
  NAND2_X1   g30720(.A1(new_n25554_), .A2(pi0235), .ZN(new_n33157_));
  OAI21_X1   g30721(.A1(new_n33156_), .A2(new_n25554_), .B(new_n33157_), .ZN(po0652));
  INV_X1     g30722(.I(new_n25547_), .ZN(new_n33159_));
  NAND2_X1   g30723(.A1(new_n33159_), .A2(pi0496), .ZN(new_n33160_));
  OAI21_X1   g30724(.A1(new_n3865_), .A2(new_n33159_), .B(new_n33160_), .ZN(po0653));
  NAND2_X1   g30725(.A1(new_n25547_), .A2(pi0239), .ZN(new_n33162_));
  OAI21_X1   g30726(.A1(pi0497), .A2(new_n25547_), .B(new_n33162_), .ZN(po0654));
  NAND2_X1   g30727(.A1(new_n33121_), .A2(pi0498), .ZN(new_n33164_));
  OAI21_X1   g30728(.A1(new_n3625_), .A2(new_n33121_), .B(new_n33164_), .ZN(po0655));
  NAND2_X1   g30729(.A1(new_n33159_), .A2(pi0499), .ZN(new_n33166_));
  OAI21_X1   g30730(.A1(new_n4430_), .A2(new_n33159_), .B(new_n33166_), .ZN(po0656));
  NAND2_X1   g30731(.A1(new_n33159_), .A2(pi0500), .ZN(new_n33168_));
  OAI21_X1   g30732(.A1(new_n3948_), .A2(new_n33159_), .B(new_n33168_), .ZN(po0657));
  NAND2_X1   g30733(.A1(new_n33159_), .A2(pi0501), .ZN(new_n33170_));
  OAI21_X1   g30734(.A1(new_n4105_), .A2(new_n33159_), .B(new_n33170_), .ZN(po0658));
  INV_X1     g30735(.I(pi0502), .ZN(new_n33172_));
  NAND2_X1   g30736(.A1(new_n25547_), .A2(pi0247), .ZN(new_n33173_));
  OAI21_X1   g30737(.A1(new_n33172_), .A2(new_n25547_), .B(new_n33173_), .ZN(po0659));
  INV_X1     g30738(.I(pi0503), .ZN(new_n33175_));
  NAND2_X1   g30739(.A1(new_n25547_), .A2(pi0245), .ZN(new_n33176_));
  OAI21_X1   g30740(.A1(new_n33175_), .A2(new_n25547_), .B(new_n33176_), .ZN(po0660));
  INV_X1     g30741(.I(pi0504), .ZN(new_n33178_));
  NAND2_X1   g30742(.A1(new_n25475_), .A2(pi0242), .ZN(new_n33179_));
  OAI21_X1   g30743(.A1(new_n33178_), .A2(new_n25475_), .B(new_n33179_), .ZN(po0661));
  INV_X1     g30744(.I(pi0505), .ZN(new_n33181_));
  NOR2_X1    g30745(.A1(new_n25319_), .A2(new_n5488_), .ZN(new_n33182_));
  NOR2_X1    g30746(.A1(new_n5475_), .A2(new_n12618_), .ZN(new_n33183_));
  NOR2_X1    g30747(.A1(new_n33182_), .A2(new_n33183_), .ZN(new_n33184_));
  INV_X1     g30748(.I(new_n33184_), .ZN(new_n33185_));
  NAND2_X1   g30749(.A1(new_n33185_), .A2(new_n3097_), .ZN(new_n33186_));
  NOR2_X1    g30750(.A1(new_n33159_), .A2(new_n33186_), .ZN(new_n33187_));
  NOR2_X1    g30751(.A1(new_n25474_), .A2(new_n3097_), .ZN(new_n33188_));
  NAND2_X1   g30752(.A1(new_n33188_), .A2(new_n33181_), .ZN(new_n33189_));
  OAI22_X1   g30753(.A1(new_n33187_), .A2(new_n33181_), .B1(new_n25459_), .B2(new_n33189_), .ZN(po0662));
  INV_X1     g30754(.I(pi0506), .ZN(new_n33191_));
  NAND2_X1   g30755(.A1(new_n25475_), .A2(pi0241), .ZN(new_n33192_));
  OAI21_X1   g30756(.A1(new_n33191_), .A2(new_n25475_), .B(new_n33192_), .ZN(po0663));
  INV_X1     g30757(.I(pi0507), .ZN(new_n33194_));
  NAND2_X1   g30758(.A1(new_n25475_), .A2(pi0238), .ZN(new_n33195_));
  OAI21_X1   g30759(.A1(new_n33194_), .A2(new_n25475_), .B(new_n33195_), .ZN(po0664));
  INV_X1     g30760(.I(pi0508), .ZN(new_n33197_));
  NAND2_X1   g30761(.A1(new_n25475_), .A2(pi0247), .ZN(new_n33198_));
  OAI21_X1   g30762(.A1(new_n33197_), .A2(new_n25475_), .B(new_n33198_), .ZN(po0665));
  INV_X1     g30763(.I(pi0509), .ZN(new_n33200_));
  NAND2_X1   g30764(.A1(new_n25475_), .A2(pi0245), .ZN(new_n33201_));
  OAI21_X1   g30765(.A1(new_n33200_), .A2(new_n25475_), .B(new_n33201_), .ZN(po0666));
  INV_X1     g30766(.I(pi0510), .ZN(new_n33203_));
  NAND2_X1   g30767(.A1(new_n25330_), .A2(pi0242), .ZN(new_n33204_));
  OAI21_X1   g30768(.A1(new_n33203_), .A2(new_n25330_), .B(new_n33204_), .ZN(po0667));
  NOR2_X1    g30769(.A1(new_n25319_), .A2(new_n5702_), .ZN(new_n33206_));
  NOR2_X1    g30770(.A1(new_n5694_), .A2(new_n12618_), .ZN(new_n33207_));
  OR2_X2     g30771(.A1(new_n33206_), .A2(new_n33207_), .Z(new_n33208_));
  NAND2_X1   g30772(.A1(new_n33208_), .A2(new_n3097_), .ZN(new_n33209_));
  MUX2_X1    g30773(.I0(pi0511), .I1(new_n33209_), .S(new_n25330_), .Z(po0668));
  INV_X1     g30774(.I(pi0512), .ZN(new_n33211_));
  NAND2_X1   g30775(.A1(new_n25330_), .A2(pi0235), .ZN(new_n33212_));
  OAI21_X1   g30776(.A1(new_n33211_), .A2(new_n25330_), .B(new_n33212_), .ZN(po0669));
  INV_X1     g30777(.I(pi0513), .ZN(new_n33214_));
  NAND2_X1   g30778(.A1(new_n25330_), .A2(pi0244), .ZN(new_n33215_));
  OAI21_X1   g30779(.A1(new_n33214_), .A2(new_n25330_), .B(new_n33215_), .ZN(po0670));
  INV_X1     g30780(.I(pi0514), .ZN(new_n33217_));
  NAND2_X1   g30781(.A1(new_n25330_), .A2(pi0245), .ZN(new_n33218_));
  OAI21_X1   g30782(.A1(new_n33217_), .A2(new_n25330_), .B(new_n33218_), .ZN(po0671));
  INV_X1     g30783(.I(pi0515), .ZN(new_n33220_));
  NAND2_X1   g30784(.A1(new_n25330_), .A2(pi0240), .ZN(new_n33221_));
  OAI21_X1   g30785(.A1(new_n33220_), .A2(new_n25330_), .B(new_n33221_), .ZN(po0672));
  INV_X1     g30786(.I(pi0516), .ZN(new_n33223_));
  NAND2_X1   g30787(.A1(new_n25330_), .A2(pi0247), .ZN(new_n33224_));
  OAI21_X1   g30788(.A1(new_n33223_), .A2(new_n25330_), .B(new_n33224_), .ZN(po0673));
  INV_X1     g30789(.I(pi0517), .ZN(new_n33226_));
  NAND2_X1   g30790(.A1(new_n25330_), .A2(pi0238), .ZN(new_n33227_));
  OAI21_X1   g30791(.A1(new_n33226_), .A2(new_n25330_), .B(new_n33227_), .ZN(po0674));
  INV_X1     g30792(.I(pi0518), .ZN(new_n33229_));
  NOR3_X1    g30793(.A1(new_n33209_), .A2(new_n25325_), .A3(new_n25459_), .ZN(new_n33230_));
  NOR2_X1    g30794(.A1(new_n25325_), .A2(new_n3097_), .ZN(new_n33231_));
  NAND2_X1   g30795(.A1(new_n33231_), .A2(new_n33229_), .ZN(new_n33232_));
  OAI22_X1   g30796(.A1(new_n33230_), .A2(new_n33229_), .B1(new_n25459_), .B2(new_n33232_), .ZN(po0675));
  NAND2_X1   g30797(.A1(new_n25460_), .A2(pi0239), .ZN(new_n33234_));
  OAI21_X1   g30798(.A1(pi0519), .A2(new_n25460_), .B(new_n33234_), .ZN(po0676));
  INV_X1     g30799(.I(pi0520), .ZN(new_n33236_));
  NAND2_X1   g30800(.A1(new_n25460_), .A2(pi0246), .ZN(new_n33237_));
  OAI21_X1   g30801(.A1(new_n33236_), .A2(new_n25460_), .B(new_n33237_), .ZN(po0677));
  INV_X1     g30802(.I(pi0521), .ZN(new_n33239_));
  NAND2_X1   g30803(.A1(new_n25460_), .A2(pi0248), .ZN(new_n33240_));
  OAI21_X1   g30804(.A1(new_n33239_), .A2(new_n25460_), .B(new_n33240_), .ZN(po0678));
  INV_X1     g30805(.I(pi0522), .ZN(new_n33242_));
  NAND2_X1   g30806(.A1(new_n25460_), .A2(pi0238), .ZN(new_n33243_));
  OAI21_X1   g30807(.A1(new_n33242_), .A2(new_n25460_), .B(new_n33243_), .ZN(po0679));
  INV_X1     g30808(.I(pi0523), .ZN(new_n33245_));
  INV_X1     g30809(.I(new_n26407_), .ZN(new_n33246_));
  NOR2_X1    g30810(.A1(new_n33246_), .A2(new_n33209_), .ZN(new_n33247_));
  NAND2_X1   g30811(.A1(new_n33231_), .A2(new_n33245_), .ZN(new_n33248_));
  OAI22_X1   g30812(.A1(new_n33247_), .A2(new_n33245_), .B1(new_n25553_), .B2(new_n33248_), .ZN(po0680));
  NAND2_X1   g30813(.A1(new_n26407_), .A2(pi0239), .ZN(new_n33250_));
  OAI21_X1   g30814(.A1(pi0524), .A2(new_n26407_), .B(new_n33250_), .ZN(po0681));
  INV_X1     g30815(.I(pi0525), .ZN(new_n33252_));
  NAND2_X1   g30816(.A1(new_n26407_), .A2(pi0245), .ZN(new_n33253_));
  OAI21_X1   g30817(.A1(new_n33252_), .A2(new_n26407_), .B(new_n33253_), .ZN(po0682));
  NAND2_X1   g30818(.A1(new_n33246_), .A2(pi0526), .ZN(new_n33255_));
  OAI21_X1   g30819(.A1(new_n4430_), .A2(new_n33246_), .B(new_n33255_), .ZN(po0683));
  INV_X1     g30820(.I(pi0527), .ZN(new_n33257_));
  NAND2_X1   g30821(.A1(new_n26407_), .A2(pi0247), .ZN(new_n33258_));
  OAI21_X1   g30822(.A1(new_n33257_), .A2(new_n26407_), .B(new_n33258_), .ZN(po0684));
  NAND2_X1   g30823(.A1(new_n33246_), .A2(pi0528), .ZN(new_n33260_));
  OAI21_X1   g30824(.A1(new_n3865_), .A2(new_n33246_), .B(new_n33260_), .ZN(po0685));
  INV_X1     g30825(.I(pi0529), .ZN(new_n33262_));
  NAND2_X1   g30826(.A1(new_n26407_), .A2(pi0238), .ZN(new_n33263_));
  OAI21_X1   g30827(.A1(new_n33262_), .A2(new_n26407_), .B(new_n33263_), .ZN(po0686));
  INV_X1     g30828(.I(pi0530), .ZN(new_n33265_));
  NAND2_X1   g30829(.A1(new_n26407_), .A2(pi0240), .ZN(new_n33266_));
  OAI21_X1   g30830(.A1(new_n33265_), .A2(new_n26407_), .B(new_n33266_), .ZN(po0687));
  INV_X1     g30831(.I(pi0531), .ZN(new_n33268_));
  NAND2_X1   g30832(.A1(new_n25467_), .A2(pi0235), .ZN(new_n33269_));
  OAI21_X1   g30833(.A1(new_n33268_), .A2(new_n25467_), .B(new_n33269_), .ZN(po0688));
  INV_X1     g30834(.I(pi0532), .ZN(new_n33271_));
  NAND2_X1   g30835(.A1(new_n25467_), .A2(pi0247), .ZN(new_n33272_));
  OAI21_X1   g30836(.A1(new_n33271_), .A2(new_n25467_), .B(new_n33272_), .ZN(po0689));
  INV_X1     g30837(.I(pi0533), .ZN(new_n33274_));
  NAND2_X1   g30838(.A1(new_n25475_), .A2(pi0235), .ZN(new_n33275_));
  OAI21_X1   g30839(.A1(new_n33274_), .A2(new_n25475_), .B(new_n33275_), .ZN(po0690));
  NAND2_X1   g30840(.A1(new_n25475_), .A2(pi0239), .ZN(new_n33277_));
  OAI21_X1   g30841(.A1(pi0534), .A2(new_n25475_), .B(new_n33277_), .ZN(po0691));
  INV_X1     g30842(.I(pi0535), .ZN(new_n33279_));
  NAND2_X1   g30843(.A1(new_n25475_), .A2(pi0240), .ZN(new_n33280_));
  OAI21_X1   g30844(.A1(new_n33279_), .A2(new_n25475_), .B(new_n33280_), .ZN(po0692));
  INV_X1     g30845(.I(new_n25475_), .ZN(new_n33282_));
  NAND2_X1   g30846(.A1(new_n33282_), .A2(pi0536), .ZN(new_n33283_));
  OAI21_X1   g30847(.A1(new_n4430_), .A2(new_n33282_), .B(new_n33283_), .ZN(po0693));
  INV_X1     g30848(.I(pi0537), .ZN(new_n33285_));
  NAND2_X1   g30849(.A1(new_n25475_), .A2(pi0248), .ZN(new_n33286_));
  OAI21_X1   g30850(.A1(new_n33285_), .A2(new_n25475_), .B(new_n33286_), .ZN(po0694));
  INV_X1     g30851(.I(pi0538), .ZN(new_n33288_));
  NAND2_X1   g30852(.A1(new_n25475_), .A2(pi0249), .ZN(new_n33289_));
  OAI21_X1   g30853(.A1(new_n33288_), .A2(new_n25475_), .B(new_n33289_), .ZN(po0695));
  INV_X1     g30854(.I(pi0539), .ZN(new_n33291_));
  NAND2_X1   g30855(.A1(new_n25547_), .A2(pi0242), .ZN(new_n33292_));
  OAI21_X1   g30856(.A1(new_n33291_), .A2(new_n25547_), .B(new_n33292_), .ZN(po0696));
  INV_X1     g30857(.I(pi0540), .ZN(new_n33294_));
  NAND2_X1   g30858(.A1(new_n25547_), .A2(pi0235), .ZN(new_n33295_));
  OAI21_X1   g30859(.A1(new_n33294_), .A2(new_n25547_), .B(new_n33295_), .ZN(po0697));
  INV_X1     g30860(.I(pi0541), .ZN(new_n33297_));
  NAND2_X1   g30861(.A1(new_n25547_), .A2(pi0244), .ZN(new_n33298_));
  OAI21_X1   g30862(.A1(new_n33297_), .A2(new_n25547_), .B(new_n33298_), .ZN(po0698));
  INV_X1     g30863(.I(pi0542), .ZN(new_n33300_));
  NAND2_X1   g30864(.A1(new_n25547_), .A2(pi0240), .ZN(new_n33301_));
  OAI21_X1   g30865(.A1(new_n33300_), .A2(new_n25547_), .B(new_n33301_), .ZN(po0699));
  NAND2_X1   g30866(.A1(new_n33159_), .A2(pi0543), .ZN(new_n33303_));
  OAI21_X1   g30867(.A1(new_n3625_), .A2(new_n33159_), .B(new_n33303_), .ZN(po0700));
  INV_X1     g30868(.I(pi0544), .ZN(new_n33305_));
  NOR2_X1    g30869(.A1(new_n33127_), .A2(new_n33186_), .ZN(new_n33306_));
  NAND2_X1   g30870(.A1(new_n33188_), .A2(new_n33305_), .ZN(new_n33307_));
  OAI22_X1   g30871(.A1(new_n33306_), .A2(new_n33305_), .B1(new_n25553_), .B2(new_n33307_), .ZN(po0701));
  INV_X1     g30872(.I(pi0545), .ZN(new_n33309_));
  NAND2_X1   g30873(.A1(new_n25554_), .A2(pi0245), .ZN(new_n33310_));
  OAI21_X1   g30874(.A1(new_n33309_), .A2(new_n25554_), .B(new_n33310_), .ZN(po0702));
  NAND2_X1   g30875(.A1(new_n33127_), .A2(pi0546), .ZN(new_n33312_));
  OAI21_X1   g30876(.A1(new_n4430_), .A2(new_n33127_), .B(new_n33312_), .ZN(po0703));
  INV_X1     g30877(.I(pi0547), .ZN(new_n33314_));
  NAND2_X1   g30878(.A1(new_n25554_), .A2(pi0247), .ZN(new_n33315_));
  OAI21_X1   g30879(.A1(new_n33314_), .A2(new_n25554_), .B(new_n33315_), .ZN(po0704));
  NAND2_X1   g30880(.A1(new_n33127_), .A2(pi0548), .ZN(new_n33317_));
  OAI21_X1   g30881(.A1(new_n4105_), .A2(new_n33127_), .B(new_n33317_), .ZN(po0705));
  INV_X1     g30882(.I(pi0549), .ZN(new_n33319_));
  NAND2_X1   g30883(.A1(new_n26388_), .A2(pi0235), .ZN(new_n33320_));
  OAI21_X1   g30884(.A1(new_n33319_), .A2(new_n26388_), .B(new_n33320_), .ZN(po0706));
  NAND2_X1   g30885(.A1(new_n26388_), .A2(pi0239), .ZN(new_n33322_));
  OAI21_X1   g30886(.A1(pi0550), .A2(new_n26388_), .B(new_n33322_), .ZN(po0707));
  INV_X1     g30887(.I(pi0551), .ZN(new_n33324_));
  NAND2_X1   g30888(.A1(new_n26388_), .A2(pi0240), .ZN(new_n33325_));
  OAI21_X1   g30889(.A1(new_n33324_), .A2(new_n26388_), .B(new_n33325_), .ZN(po0708));
  INV_X1     g30890(.I(pi0552), .ZN(new_n33327_));
  NAND2_X1   g30891(.A1(new_n26388_), .A2(pi0247), .ZN(new_n33328_));
  OAI21_X1   g30892(.A1(new_n33327_), .A2(new_n26388_), .B(new_n33328_), .ZN(po0709));
  INV_X1     g30893(.I(pi0553), .ZN(new_n33330_));
  NAND2_X1   g30894(.A1(new_n26388_), .A2(pi0241), .ZN(new_n33331_));
  OAI21_X1   g30895(.A1(new_n33330_), .A2(new_n26388_), .B(new_n33331_), .ZN(po0710));
  INV_X1     g30896(.I(pi0554), .ZN(new_n33333_));
  NAND2_X1   g30897(.A1(new_n26388_), .A2(pi0248), .ZN(new_n33334_));
  OAI21_X1   g30898(.A1(new_n33333_), .A2(new_n26388_), .B(new_n33334_), .ZN(po0711));
  INV_X1     g30899(.I(pi0555), .ZN(new_n33336_));
  NAND2_X1   g30900(.A1(new_n26388_), .A2(pi0249), .ZN(new_n33337_));
  OAI21_X1   g30901(.A1(new_n33336_), .A2(new_n26388_), .B(new_n33337_), .ZN(po0712));
  INV_X1     g30902(.I(pi0556), .ZN(new_n33339_));
  NAND2_X1   g30903(.A1(new_n25467_), .A2(pi0242), .ZN(new_n33340_));
  OAI21_X1   g30904(.A1(new_n33339_), .A2(new_n25467_), .B(new_n33340_), .ZN(po0713));
  INV_X1     g30905(.I(pi0557), .ZN(new_n33342_));
  NOR2_X1    g30906(.A1(new_n33282_), .A2(new_n33186_), .ZN(new_n33343_));
  NAND2_X1   g30907(.A1(new_n33188_), .A2(new_n33342_), .ZN(new_n33344_));
  OAI22_X1   g30908(.A1(new_n33343_), .A2(new_n33342_), .B1(new_n25329_), .B2(new_n33344_), .ZN(po0714));
  INV_X1     g30909(.I(pi0558), .ZN(new_n33346_));
  NAND2_X1   g30910(.A1(new_n25475_), .A2(pi0244), .ZN(new_n33347_));
  OAI21_X1   g30911(.A1(new_n33346_), .A2(new_n25475_), .B(new_n33347_), .ZN(po0715));
  INV_X1     g30912(.I(pi0559), .ZN(new_n33349_));
  NAND2_X1   g30913(.A1(new_n25330_), .A2(pi0241), .ZN(new_n33350_));
  OAI21_X1   g30914(.A1(new_n33349_), .A2(new_n25330_), .B(new_n33350_), .ZN(po0716));
  INV_X1     g30915(.I(pi0560), .ZN(new_n33352_));
  NAND2_X1   g30916(.A1(new_n25467_), .A2(pi0240), .ZN(new_n33353_));
  OAI21_X1   g30917(.A1(new_n33352_), .A2(new_n25467_), .B(new_n33353_), .ZN(po0717));
  INV_X1     g30918(.I(pi0561), .ZN(new_n33355_));
  NAND2_X1   g30919(.A1(new_n25460_), .A2(pi0247), .ZN(new_n33356_));
  OAI21_X1   g30920(.A1(new_n33355_), .A2(new_n25460_), .B(new_n33356_), .ZN(po0718));
  NAND2_X1   g30921(.A1(new_n33121_), .A2(pi0562), .ZN(new_n33358_));
  OAI21_X1   g30922(.A1(new_n3948_), .A2(new_n33121_), .B(new_n33358_), .ZN(po0719));
  INV_X1     g30923(.I(pi0563), .ZN(new_n33360_));
  NAND2_X1   g30924(.A1(new_n26388_), .A2(pi0246), .ZN(new_n33361_));
  OAI21_X1   g30925(.A1(new_n33360_), .A2(new_n26388_), .B(new_n33361_), .ZN(po0720));
  INV_X1     g30926(.I(pi0564), .ZN(new_n33363_));
  NAND2_X1   g30927(.A1(new_n25467_), .A2(pi0246), .ZN(new_n33364_));
  OAI21_X1   g30928(.A1(new_n33363_), .A2(new_n25467_), .B(new_n33364_), .ZN(po0721));
  NAND2_X1   g30929(.A1(new_n33121_), .A2(pi0565), .ZN(new_n33366_));
  OAI21_X1   g30930(.A1(new_n4105_), .A2(new_n33121_), .B(new_n33366_), .ZN(po0722));
  INV_X1     g30931(.I(pi0566), .ZN(new_n33368_));
  NAND2_X1   g30932(.A1(new_n25467_), .A2(pi0244), .ZN(new_n33369_));
  OAI21_X1   g30933(.A1(new_n33368_), .A2(new_n25467_), .B(new_n33369_), .ZN(po0723));
  NOR3_X1    g30934(.A1(new_n3040_), .A2(pi0567), .A3(pi1093), .ZN(new_n33371_));
  INV_X1     g30935(.I(new_n33371_), .ZN(new_n33372_));
  NOR4_X1    g30936(.A1(new_n15241_), .A2(new_n12751_), .A3(new_n27382_), .A4(new_n15232_), .ZN(new_n33373_));
  NAND2_X1   g30937(.A1(new_n33373_), .A2(new_n15807_), .ZN(new_n33374_));
  NAND3_X1   g30938(.A1(new_n33374_), .A2(pi0789), .A3(new_n33372_), .ZN(new_n33375_));
  INV_X1     g30939(.I(new_n33375_), .ZN(new_n33376_));
  NOR3_X1    g30940(.A1(new_n33373_), .A2(pi0789), .A3(new_n33371_), .ZN(new_n33377_));
  NOR2_X1    g30941(.A1(new_n33376_), .A2(new_n33377_), .ZN(new_n33378_));
  INV_X1     g30942(.I(new_n33378_), .ZN(new_n33379_));
  NAND2_X1   g30943(.A1(new_n13510_), .A2(pi0680), .ZN(new_n33380_));
  OAI21_X1   g30944(.A1(new_n33380_), .A2(new_n14285_), .B(new_n33372_), .ZN(new_n33381_));
  INV_X1     g30945(.I(new_n33381_), .ZN(new_n33382_));
  NOR2_X1    g30946(.A1(new_n33382_), .A2(new_n14290_), .ZN(new_n33383_));
  OAI21_X1   g30947(.A1(new_n33375_), .A2(new_n12909_), .B(new_n33383_), .ZN(new_n33384_));
  AOI21_X1   g30948(.A1(new_n33379_), .A2(new_n33384_), .B(new_n14303_), .ZN(new_n33385_));
  NAND2_X1   g30949(.A1(new_n33383_), .A2(new_n12911_), .ZN(new_n33386_));
  OAI21_X1   g30950(.A1(new_n33386_), .A2(new_n12814_), .B(new_n33372_), .ZN(new_n33387_));
  NAND2_X1   g30951(.A1(new_n33387_), .A2(new_n12746_), .ZN(new_n33388_));
  OAI21_X1   g30952(.A1(new_n33386_), .A2(pi0641), .B(new_n33372_), .ZN(new_n33389_));
  AOI22_X1   g30953(.A1(new_n33378_), .A2(new_n25833_), .B1(new_n12748_), .B2(new_n33389_), .ZN(new_n33390_));
  AOI21_X1   g30954(.A1(new_n33390_), .A2(new_n33388_), .B(new_n12808_), .ZN(new_n33391_));
  OAI21_X1   g30955(.A1(new_n33391_), .A2(new_n33385_), .B(new_n15824_), .ZN(new_n33392_));
  INV_X1     g30956(.I(new_n33392_), .ZN(new_n33393_));
  NOR2_X1    g30957(.A1(new_n14292_), .A2(new_n33382_), .ZN(new_n33394_));
  INV_X1     g30958(.I(new_n33394_), .ZN(new_n33395_));
  OAI21_X1   g30959(.A1(new_n33395_), .A2(new_n12920_), .B(new_n33372_), .ZN(new_n33396_));
  NOR2_X1    g30960(.A1(new_n17504_), .A2(new_n33371_), .ZN(new_n33397_));
  AOI21_X1   g30961(.A1(new_n33379_), .A2(new_n17504_), .B(new_n33397_), .ZN(new_n33398_));
  INV_X1     g30962(.I(new_n33398_), .ZN(new_n33399_));
  OAI21_X1   g30963(.A1(new_n33399_), .A2(new_n15694_), .B(new_n12919_), .ZN(new_n33400_));
  AOI21_X1   g30964(.A1(pi1156), .A2(new_n33396_), .B(new_n33400_), .ZN(new_n33401_));
  OAI21_X1   g30965(.A1(new_n33395_), .A2(pi0628), .B(new_n33372_), .ZN(new_n33402_));
  OAI21_X1   g30966(.A1(new_n33399_), .A2(new_n15699_), .B(pi0629), .ZN(new_n33403_));
  AOI21_X1   g30967(.A1(new_n12742_), .A2(new_n33402_), .B(new_n33403_), .ZN(new_n33404_));
  NOR3_X1    g30968(.A1(new_n33401_), .A2(new_n33404_), .A3(new_n12937_), .ZN(new_n33405_));
  NOR2_X1    g30969(.A1(new_n33405_), .A2(new_n33393_), .ZN(new_n33406_));
  INV_X1     g30970(.I(new_n33406_), .ZN(new_n33407_));
  NAND2_X1   g30971(.A1(new_n33406_), .A2(pi0647), .ZN(new_n33408_));
  NOR2_X1    g30972(.A1(new_n33399_), .A2(new_n12943_), .ZN(new_n33409_));
  AOI21_X1   g30973(.A1(new_n12943_), .A2(new_n33371_), .B(new_n33409_), .ZN(new_n33410_));
  NAND2_X1   g30974(.A1(new_n33410_), .A2(new_n12741_), .ZN(new_n33411_));
  AOI21_X1   g30975(.A1(new_n33408_), .A2(new_n33411_), .B(new_n12965_), .ZN(new_n33412_));
  NOR2_X1    g30976(.A1(new_n33395_), .A2(new_n12951_), .ZN(new_n33413_));
  INV_X1     g30977(.I(new_n33413_), .ZN(new_n33414_));
  OAI21_X1   g30978(.A1(new_n33414_), .A2(pi0647), .B(new_n12965_), .ZN(new_n33415_));
  NOR2_X1    g30979(.A1(new_n33415_), .A2(new_n33371_), .ZN(new_n33416_));
  NOR3_X1    g30980(.A1(new_n33412_), .A2(new_n12981_), .A3(new_n33416_), .ZN(new_n33417_));
  NAND2_X1   g30981(.A1(new_n33410_), .A2(pi0647), .ZN(new_n33418_));
  OAI21_X1   g30982(.A1(new_n33407_), .A2(pi0647), .B(new_n33418_), .ZN(new_n33419_));
  OAI21_X1   g30983(.A1(new_n33414_), .A2(new_n12741_), .B(pi1157), .ZN(new_n33420_));
  OAI21_X1   g30984(.A1(new_n33420_), .A2(new_n33371_), .B(new_n12981_), .ZN(new_n33421_));
  AOI21_X1   g30985(.A1(new_n33419_), .A2(new_n12965_), .B(new_n33421_), .ZN(new_n33422_));
  OR3_X2     g30986(.A1(new_n33417_), .A2(new_n12972_), .A3(new_n33422_), .Z(new_n33423_));
  OAI21_X1   g30987(.A1(pi0787), .A2(new_n33407_), .B(new_n33423_), .ZN(new_n33424_));
  NOR2_X1    g30988(.A1(new_n33424_), .A2(new_n12975_), .ZN(new_n33425_));
  NOR2_X1    g30989(.A1(new_n33414_), .A2(new_n14300_), .ZN(new_n33426_));
  NOR2_X1    g30990(.A1(new_n33426_), .A2(new_n33371_), .ZN(new_n33427_));
  NOR2_X1    g30991(.A1(new_n33427_), .A2(pi0644), .ZN(new_n33428_));
  OAI21_X1   g30992(.A1(new_n33425_), .A2(new_n33428_), .B(pi0715), .ZN(new_n33429_));
  NAND2_X1   g30993(.A1(new_n33409_), .A2(new_n12985_), .ZN(new_n33430_));
  OAI21_X1   g30994(.A1(new_n33430_), .A2(new_n12975_), .B(new_n33372_), .ZN(new_n33431_));
  NAND2_X1   g30995(.A1(new_n33431_), .A2(new_n12740_), .ZN(new_n33432_));
  NAND3_X1   g30996(.A1(new_n33429_), .A2(pi1160), .A3(new_n33432_), .ZN(new_n33433_));
  OAI21_X1   g30997(.A1(new_n33430_), .A2(pi0644), .B(pi0715), .ZN(new_n33434_));
  NOR3_X1    g30998(.A1(new_n33426_), .A2(new_n12975_), .A3(new_n33371_), .ZN(new_n33435_));
  AOI21_X1   g30999(.A1(new_n33424_), .A2(new_n12975_), .B(new_n33435_), .ZN(new_n33436_));
  OAI22_X1   g31000(.A1(new_n33436_), .A2(pi0715), .B1(new_n33371_), .B2(new_n33434_), .ZN(new_n33437_));
  AOI21_X1   g31001(.A1(new_n33437_), .A2(new_n12739_), .B(new_n13000_), .ZN(new_n33438_));
  NOR2_X1    g31002(.A1(new_n33424_), .A2(pi0790), .ZN(new_n33439_));
  AOI21_X1   g31003(.A1(new_n33438_), .A2(new_n33433_), .B(new_n33439_), .ZN(new_n33440_));
  NAND2_X1   g31004(.A1(new_n27999_), .A2(pi1092), .ZN(new_n33441_));
  OAI22_X1   g31005(.A1(new_n33440_), .A2(new_n27999_), .B1(pi0567), .B2(new_n33441_), .ZN(po0724));
  INV_X1     g31006(.I(pi0568), .ZN(new_n33443_));
  NAND2_X1   g31007(.A1(new_n25467_), .A2(pi0245), .ZN(new_n33444_));
  OAI21_X1   g31008(.A1(new_n33443_), .A2(new_n25467_), .B(new_n33444_), .ZN(po0725));
  NAND2_X1   g31009(.A1(new_n25467_), .A2(pi0239), .ZN(new_n33446_));
  OAI21_X1   g31010(.A1(pi0569), .A2(new_n25467_), .B(new_n33446_), .ZN(po0726));
  NOR2_X1    g31011(.A1(new_n25466_), .A2(pi0570), .ZN(new_n33448_));
  NAND2_X1   g31012(.A1(new_n33231_), .A2(new_n33448_), .ZN(new_n33449_));
  OAI21_X1   g31013(.A1(new_n33121_), .A2(new_n33209_), .B(pi0570), .ZN(new_n33450_));
  NAND2_X1   g31014(.A1(new_n33450_), .A2(new_n33449_), .ZN(po0727));
  NAND2_X1   g31015(.A1(new_n33246_), .A2(pi0571), .ZN(new_n33452_));
  OAI21_X1   g31016(.A1(new_n3948_), .A2(new_n33246_), .B(new_n33452_), .ZN(po0728));
  INV_X1     g31017(.I(pi0572), .ZN(new_n33454_));
  NAND2_X1   g31018(.A1(new_n26407_), .A2(pi0244), .ZN(new_n33455_));
  OAI21_X1   g31019(.A1(new_n33454_), .A2(new_n26407_), .B(new_n33455_), .ZN(po0729));
  INV_X1     g31020(.I(pi0573), .ZN(new_n33457_));
  NAND2_X1   g31021(.A1(new_n26407_), .A2(pi0242), .ZN(new_n33458_));
  OAI21_X1   g31022(.A1(new_n33457_), .A2(new_n26407_), .B(new_n33458_), .ZN(po0730));
  INV_X1     g31023(.I(pi0574), .ZN(new_n33460_));
  NAND2_X1   g31024(.A1(new_n25460_), .A2(pi0241), .ZN(new_n33461_));
  OAI21_X1   g31025(.A1(new_n33460_), .A2(new_n25460_), .B(new_n33461_), .ZN(po0731));
  INV_X1     g31026(.I(pi0575), .ZN(new_n33463_));
  NAND2_X1   g31027(.A1(new_n26407_), .A2(pi0235), .ZN(new_n33464_));
  OAI21_X1   g31028(.A1(new_n33463_), .A2(new_n26407_), .B(new_n33464_), .ZN(po0732));
  NAND2_X1   g31029(.A1(new_n33246_), .A2(pi0576), .ZN(new_n33466_));
  OAI21_X1   g31030(.A1(new_n4105_), .A2(new_n33246_), .B(new_n33466_), .ZN(po0733));
  INV_X1     g31031(.I(pi0577), .ZN(new_n33468_));
  NAND2_X1   g31032(.A1(new_n26388_), .A2(pi0238), .ZN(new_n33469_));
  OAI21_X1   g31033(.A1(new_n33468_), .A2(new_n26388_), .B(new_n33469_), .ZN(po0734));
  INV_X1     g31034(.I(pi0578), .ZN(new_n33471_));
  NAND2_X1   g31035(.A1(new_n25460_), .A2(pi0249), .ZN(new_n33472_));
  OAI21_X1   g31036(.A1(new_n33471_), .A2(new_n25460_), .B(new_n33472_), .ZN(po0735));
  INV_X1     g31037(.I(pi0579), .ZN(new_n33474_));
  NAND2_X1   g31038(.A1(new_n25330_), .A2(pi0249), .ZN(new_n33475_));
  OAI21_X1   g31039(.A1(new_n33474_), .A2(new_n25330_), .B(new_n33475_), .ZN(po0736));
  INV_X1     g31040(.I(pi0580), .ZN(new_n33477_));
  NAND2_X1   g31041(.A1(new_n26388_), .A2(pi0245), .ZN(new_n33478_));
  OAI21_X1   g31042(.A1(new_n33477_), .A2(new_n26388_), .B(new_n33478_), .ZN(po0737));
  INV_X1     g31043(.I(pi0581), .ZN(new_n33480_));
  NAND2_X1   g31044(.A1(new_n25460_), .A2(pi0235), .ZN(new_n33481_));
  OAI21_X1   g31045(.A1(new_n33480_), .A2(new_n25460_), .B(new_n33481_), .ZN(po0738));
  INV_X1     g31046(.I(pi0582), .ZN(new_n33483_));
  NAND2_X1   g31047(.A1(new_n25460_), .A2(pi0240), .ZN(new_n33484_));
  OAI21_X1   g31048(.A1(new_n33483_), .A2(new_n25460_), .B(new_n33484_), .ZN(po0739));
  INV_X1     g31049(.I(pi0584), .ZN(new_n33486_));
  NAND2_X1   g31050(.A1(new_n25460_), .A2(pi0245), .ZN(new_n33487_));
  OAI21_X1   g31051(.A1(new_n33486_), .A2(new_n25460_), .B(new_n33487_), .ZN(po0741));
  INV_X1     g31052(.I(pi0585), .ZN(new_n33489_));
  NAND2_X1   g31053(.A1(new_n25460_), .A2(pi0244), .ZN(new_n33490_));
  OAI21_X1   g31054(.A1(new_n33489_), .A2(new_n25460_), .B(new_n33490_), .ZN(po0742));
  INV_X1     g31055(.I(pi0586), .ZN(new_n33492_));
  NAND2_X1   g31056(.A1(new_n25460_), .A2(pi0242), .ZN(new_n33493_));
  OAI21_X1   g31057(.A1(new_n33492_), .A2(new_n25460_), .B(new_n33493_), .ZN(po0743));
  NOR2_X1    g31058(.A1(new_n15232_), .A2(new_n25969_), .ZN(new_n33495_));
  NAND4_X1   g31059(.A1(new_n15245_), .A2(pi0230), .A3(new_n12754_), .A4(new_n33495_), .ZN(new_n33496_));
  OAI22_X1   g31060(.A1(new_n33496_), .A2(new_n22504_), .B1(pi0230), .B2(new_n5700_), .ZN(po0744));
  NOR3_X1    g31061(.A1(new_n5428_), .A2(new_n3045_), .A3(pi0123), .ZN(new_n33498_));
  NAND2_X1   g31062(.A1(new_n33498_), .A2(pi0591), .ZN(new_n33499_));
  INV_X1     g31063(.I(new_n33498_), .ZN(new_n33500_));
  NAND2_X1   g31064(.A1(new_n33500_), .A2(pi0588), .ZN(new_n33501_));
  AOI21_X1   g31065(.A1(new_n33501_), .A2(new_n33499_), .B(new_n32625_), .ZN(po0745));
  INV_X1     g31066(.I(pi0202), .ZN(new_n33503_));
  AOI21_X1   g31067(.A1(new_n33208_), .A2(new_n33503_), .B(pi0233), .ZN(new_n33504_));
  OAI21_X1   g31068(.A1(pi0205), .A2(new_n33184_), .B(new_n33504_), .ZN(new_n33505_));
  INV_X1     g31069(.I(pi0201), .ZN(new_n33506_));
  AOI21_X1   g31070(.A1(new_n33208_), .A2(new_n33506_), .B(new_n25326_), .ZN(new_n33507_));
  OAI21_X1   g31071(.A1(pi0204), .A2(new_n33184_), .B(new_n33507_), .ZN(new_n33508_));
  NAND3_X1   g31072(.A1(new_n33505_), .A2(new_n33508_), .A3(pi0237), .ZN(new_n33509_));
  INV_X1     g31073(.I(pi0203), .ZN(new_n33510_));
  AOI21_X1   g31074(.A1(new_n33208_), .A2(new_n33510_), .B(pi0233), .ZN(new_n33511_));
  OAI21_X1   g31075(.A1(pi0218), .A2(new_n33184_), .B(new_n33511_), .ZN(new_n33512_));
  INV_X1     g31076(.I(pi0220), .ZN(new_n33513_));
  AOI21_X1   g31077(.A1(new_n33208_), .A2(new_n33513_), .B(new_n25326_), .ZN(new_n33514_));
  OAI21_X1   g31078(.A1(pi0206), .A2(new_n33184_), .B(new_n33514_), .ZN(new_n33515_));
  NAND3_X1   g31079(.A1(new_n33512_), .A2(new_n33515_), .A3(new_n25327_), .ZN(new_n33516_));
  NAND2_X1   g31080(.A1(new_n33509_), .A2(new_n33516_), .ZN(po0746));
  NOR2_X1    g31081(.A1(new_n33500_), .A2(pi0588), .ZN(new_n33518_));
  NOR2_X1    g31082(.A1(new_n33498_), .A2(pi0590), .ZN(new_n33519_));
  OAI21_X1   g31083(.A1(new_n33518_), .A2(new_n33519_), .B(new_n32624_), .ZN(po0747));
  NAND2_X1   g31084(.A1(new_n33498_), .A2(pi0592), .ZN(new_n33521_));
  NAND2_X1   g31085(.A1(new_n33500_), .A2(pi0591), .ZN(new_n33522_));
  AOI21_X1   g31086(.A1(new_n33522_), .A2(new_n33521_), .B(new_n32625_), .ZN(po0748));
  NAND2_X1   g31087(.A1(new_n33498_), .A2(pi0590), .ZN(new_n33524_));
  NAND2_X1   g31088(.A1(new_n33500_), .A2(pi0592), .ZN(new_n33525_));
  AOI21_X1   g31089(.A1(new_n33525_), .A2(new_n33524_), .B(new_n32625_), .ZN(po0749));
  XNOR2_X1   g31090(.A1(pi0246), .A2(pi0487), .ZN(new_n33527_));
  XOR2_X1    g31091(.A1(pi0234), .A2(pi0511), .Z(new_n33528_));
  INV_X1     g31092(.I(new_n33528_), .ZN(new_n33529_));
  NAND3_X1   g31093(.A1(new_n33208_), .A2(new_n33527_), .A3(new_n33529_), .ZN(new_n33530_));
  XOR2_X1    g31094(.A1(pi0249), .A2(pi0579), .Z(new_n33531_));
  NOR2_X1    g31095(.A1(new_n33530_), .A2(new_n33531_), .ZN(new_n33532_));
  NOR2_X1    g31096(.A1(new_n33532_), .A2(pi0537), .ZN(new_n33533_));
  XNOR2_X1   g31097(.A1(pi0246), .A2(pi0536), .ZN(new_n33534_));
  INV_X1     g31098(.I(new_n33534_), .ZN(new_n33535_));
  XOR2_X1    g31099(.A1(pi0234), .A2(pi0557), .Z(new_n33536_));
  XOR2_X1    g31100(.A1(pi0249), .A2(pi0538), .Z(new_n33537_));
  NOR4_X1    g31101(.A1(new_n33184_), .A2(new_n33535_), .A3(new_n33536_), .A4(new_n33537_), .ZN(new_n33538_));
  INV_X1     g31102(.I(new_n33538_), .ZN(new_n33539_));
  INV_X1     g31103(.I(new_n33531_), .ZN(new_n33540_));
  NOR4_X1    g31104(.A1(new_n33184_), .A2(pi0538), .A3(new_n33535_), .A4(new_n33536_), .ZN(new_n33541_));
  AOI21_X1   g31105(.A1(new_n33541_), .A2(pi0579), .B(new_n33540_), .ZN(new_n33542_));
  OAI21_X1   g31106(.A1(new_n33542_), .A2(new_n33530_), .B(new_n33539_), .ZN(new_n33543_));
  NOR2_X1    g31107(.A1(new_n33543_), .A2(new_n33285_), .ZN(new_n33544_));
  OAI21_X1   g31108(.A1(new_n33544_), .A2(new_n33533_), .B(pi0248), .ZN(new_n33545_));
  OAI21_X1   g31109(.A1(new_n33539_), .A2(pi0537), .B(new_n4105_), .ZN(new_n33546_));
  NAND3_X1   g31110(.A1(new_n33545_), .A2(pi0481), .A3(new_n33546_), .ZN(new_n33547_));
  NOR2_X1    g31111(.A1(new_n33543_), .A2(pi0537), .ZN(new_n33548_));
  NOR2_X1    g31112(.A1(new_n33532_), .A2(new_n33285_), .ZN(new_n33549_));
  OAI21_X1   g31113(.A1(new_n33548_), .A2(new_n33549_), .B(new_n4105_), .ZN(new_n33550_));
  OAI21_X1   g31114(.A1(new_n33539_), .A2(new_n33285_), .B(pi0248), .ZN(new_n33551_));
  NAND3_X1   g31115(.A1(new_n33550_), .A2(new_n33118_), .A3(new_n33551_), .ZN(new_n33552_));
  AND2_X2    g31116(.A1(new_n33547_), .A2(new_n33552_), .Z(new_n33553_));
  NAND2_X1   g31117(.A1(new_n33553_), .A2(pi0559), .ZN(new_n33554_));
  XOR2_X1    g31118(.A1(pi0248), .A2(pi0537), .Z(new_n33555_));
  OAI21_X1   g31119(.A1(new_n33539_), .A2(new_n33555_), .B(new_n33349_), .ZN(new_n33556_));
  AOI21_X1   g31120(.A1(new_n33554_), .A2(new_n33556_), .B(new_n3948_), .ZN(new_n33557_));
  XOR2_X1    g31121(.A1(pi0248), .A2(pi0481), .Z(new_n33558_));
  NOR3_X1    g31122(.A1(new_n33530_), .A2(new_n33531_), .A3(new_n33558_), .ZN(new_n33559_));
  AOI21_X1   g31123(.A1(new_n33559_), .A2(new_n33349_), .B(pi0241), .ZN(new_n33560_));
  NOR3_X1    g31124(.A1(new_n33557_), .A2(new_n33191_), .A3(new_n33560_), .ZN(new_n33561_));
  NAND2_X1   g31125(.A1(new_n33553_), .A2(new_n33349_), .ZN(new_n33562_));
  OAI21_X1   g31126(.A1(new_n33539_), .A2(new_n33555_), .B(pi0559), .ZN(new_n33563_));
  AOI21_X1   g31127(.A1(new_n33562_), .A2(new_n33563_), .B(pi0241), .ZN(new_n33564_));
  AOI21_X1   g31128(.A1(new_n33559_), .A2(pi0559), .B(new_n3948_), .ZN(new_n33565_));
  NOR3_X1    g31129(.A1(new_n33564_), .A2(pi0506), .A3(new_n33565_), .ZN(new_n33566_));
  OR2_X2     g31130(.A1(new_n33561_), .A2(new_n33566_), .Z(new_n33567_));
  NOR2_X1    g31131(.A1(new_n33567_), .A2(new_n33220_), .ZN(new_n33568_));
  NOR2_X1    g31132(.A1(new_n33539_), .A2(new_n33555_), .ZN(new_n33569_));
  XNOR2_X1   g31133(.A1(pi0241), .A2(pi0506), .ZN(new_n33570_));
  NAND2_X1   g31134(.A1(new_n33569_), .A2(new_n33570_), .ZN(new_n33571_));
  INV_X1     g31135(.I(new_n33571_), .ZN(new_n33572_));
  NOR2_X1    g31136(.A1(new_n33572_), .A2(pi0515), .ZN(new_n33573_));
  OAI21_X1   g31137(.A1(new_n33568_), .A2(new_n33573_), .B(pi0240), .ZN(new_n33574_));
  XNOR2_X1   g31138(.A1(pi0241), .A2(pi0559), .ZN(new_n33575_));
  NAND2_X1   g31139(.A1(new_n33559_), .A2(new_n33575_), .ZN(new_n33576_));
  OAI21_X1   g31140(.A1(new_n33576_), .A2(pi0515), .B(new_n4587_), .ZN(new_n33577_));
  NAND3_X1   g31141(.A1(new_n33574_), .A2(pi0535), .A3(new_n33577_), .ZN(new_n33578_));
  NOR2_X1    g31142(.A1(new_n33567_), .A2(pi0515), .ZN(new_n33579_));
  NOR2_X1    g31143(.A1(new_n33572_), .A2(new_n33220_), .ZN(new_n33580_));
  OAI21_X1   g31144(.A1(new_n33579_), .A2(new_n33580_), .B(new_n4587_), .ZN(new_n33581_));
  OAI21_X1   g31145(.A1(new_n33576_), .A2(new_n33220_), .B(pi0240), .ZN(new_n33582_));
  NAND3_X1   g31146(.A1(new_n33581_), .A2(new_n33279_), .A3(new_n33582_), .ZN(new_n33583_));
  AND2_X2    g31147(.A1(new_n33578_), .A2(new_n33583_), .Z(new_n33584_));
  NAND2_X1   g31148(.A1(new_n33584_), .A2(pi0534), .ZN(new_n33585_));
  INV_X1     g31149(.I(pi0534), .ZN(new_n33586_));
  XOR2_X1    g31150(.A1(pi0240), .A2(pi0515), .Z(new_n33587_));
  NOR2_X1    g31151(.A1(new_n33576_), .A2(new_n33587_), .ZN(new_n33588_));
  INV_X1     g31152(.I(new_n33588_), .ZN(new_n33589_));
  NAND2_X1   g31153(.A1(new_n33589_), .A2(new_n33586_), .ZN(new_n33590_));
  NAND2_X1   g31154(.A1(new_n33585_), .A2(new_n33590_), .ZN(new_n33591_));
  XOR2_X1    g31155(.A1(pi0240), .A2(pi0535), .Z(new_n33592_));
  NOR2_X1    g31156(.A1(new_n33571_), .A2(new_n33592_), .ZN(new_n33593_));
  AOI21_X1   g31157(.A1(new_n33593_), .A2(new_n33586_), .B(new_n3476_), .ZN(new_n33594_));
  AOI21_X1   g31158(.A1(new_n33591_), .A2(new_n3476_), .B(new_n33594_), .ZN(new_n33595_));
  NAND2_X1   g31159(.A1(new_n33584_), .A2(new_n33586_), .ZN(new_n33596_));
  NAND2_X1   g31160(.A1(new_n33589_), .A2(pi0534), .ZN(new_n33597_));
  NAND2_X1   g31161(.A1(new_n33596_), .A2(new_n33597_), .ZN(new_n33598_));
  AOI21_X1   g31162(.A1(new_n33593_), .A2(pi0534), .B(pi0239), .ZN(new_n33599_));
  AOI21_X1   g31163(.A1(new_n33598_), .A2(pi0239), .B(new_n33599_), .ZN(new_n33600_));
  MUX2_X1    g31164(.I0(new_n33600_), .I1(new_n33595_), .S(pi0488), .Z(new_n33601_));
  NOR2_X1    g31165(.A1(new_n33601_), .A2(new_n33178_), .ZN(new_n33602_));
  XNOR2_X1   g31166(.A1(pi0239), .A2(pi0488), .ZN(new_n33603_));
  NOR2_X1    g31167(.A1(new_n33589_), .A2(new_n33603_), .ZN(new_n33604_));
  NOR2_X1    g31168(.A1(new_n33604_), .A2(pi0504), .ZN(new_n33605_));
  OAI21_X1   g31169(.A1(new_n33602_), .A2(new_n33605_), .B(pi0242), .ZN(new_n33606_));
  XOR2_X1    g31170(.A1(pi0239), .A2(pi0534), .Z(new_n33607_));
  NAND2_X1   g31171(.A1(new_n33593_), .A2(new_n33607_), .ZN(new_n33608_));
  OAI21_X1   g31172(.A1(new_n33608_), .A2(pi0504), .B(new_n5143_), .ZN(new_n33609_));
  NAND3_X1   g31173(.A1(new_n33606_), .A2(pi0510), .A3(new_n33609_), .ZN(new_n33610_));
  NOR2_X1    g31174(.A1(new_n33601_), .A2(pi0504), .ZN(new_n33611_));
  NOR2_X1    g31175(.A1(new_n33604_), .A2(new_n33178_), .ZN(new_n33612_));
  OAI21_X1   g31176(.A1(new_n33611_), .A2(new_n33612_), .B(new_n5143_), .ZN(new_n33613_));
  OAI21_X1   g31177(.A1(new_n33608_), .A2(new_n33178_), .B(pi0242), .ZN(new_n33614_));
  NAND3_X1   g31178(.A1(new_n33613_), .A2(new_n33203_), .A3(new_n33614_), .ZN(new_n33615_));
  AND2_X2    g31179(.A1(new_n33610_), .A2(new_n33615_), .Z(new_n33616_));
  NAND2_X1   g31180(.A1(new_n33616_), .A2(pi0533), .ZN(new_n33617_));
  INV_X1     g31181(.I(new_n33604_), .ZN(new_n33618_));
  XOR2_X1    g31182(.A1(pi0242), .A2(pi0510), .Z(new_n33619_));
  NOR2_X1    g31183(.A1(new_n33618_), .A2(new_n33619_), .ZN(new_n33620_));
  INV_X1     g31184(.I(new_n33620_), .ZN(new_n33621_));
  NAND2_X1   g31185(.A1(new_n33621_), .A2(new_n33274_), .ZN(new_n33622_));
  AOI21_X1   g31186(.A1(new_n33617_), .A2(new_n33622_), .B(new_n3479_), .ZN(new_n33623_));
  XOR2_X1    g31187(.A1(pi0242), .A2(pi0504), .Z(new_n33624_));
  NOR2_X1    g31188(.A1(new_n33608_), .A2(new_n33624_), .ZN(new_n33625_));
  AOI21_X1   g31189(.A1(new_n33625_), .A2(new_n33274_), .B(pi0235), .ZN(new_n33626_));
  NOR3_X1    g31190(.A1(new_n33623_), .A2(new_n33211_), .A3(new_n33626_), .ZN(new_n33627_));
  NAND2_X1   g31191(.A1(new_n33616_), .A2(new_n33274_), .ZN(new_n33628_));
  NAND2_X1   g31192(.A1(new_n33621_), .A2(pi0533), .ZN(new_n33629_));
  AOI21_X1   g31193(.A1(new_n33628_), .A2(new_n33629_), .B(pi0235), .ZN(new_n33630_));
  AOI21_X1   g31194(.A1(new_n33625_), .A2(pi0533), .B(new_n3479_), .ZN(new_n33631_));
  NOR3_X1    g31195(.A1(new_n33630_), .A2(pi0512), .A3(new_n33631_), .ZN(new_n33632_));
  OR2_X2     g31196(.A1(new_n33627_), .A2(new_n33632_), .Z(new_n33633_));
  NOR2_X1    g31197(.A1(new_n33633_), .A2(new_n33346_), .ZN(new_n33634_));
  XNOR2_X1   g31198(.A1(pi0235), .A2(pi0512), .ZN(new_n33635_));
  NAND2_X1   g31199(.A1(new_n33620_), .A2(new_n33635_), .ZN(new_n33636_));
  INV_X1     g31200(.I(new_n33636_), .ZN(new_n33637_));
  NOR2_X1    g31201(.A1(new_n33637_), .A2(pi0558), .ZN(new_n33638_));
  OAI21_X1   g31202(.A1(new_n33634_), .A2(new_n33638_), .B(pi0244), .ZN(new_n33639_));
  XNOR2_X1   g31203(.A1(pi0235), .A2(pi0533), .ZN(new_n33640_));
  NAND2_X1   g31204(.A1(new_n33625_), .A2(new_n33640_), .ZN(new_n33641_));
  OAI21_X1   g31205(.A1(new_n33641_), .A2(pi0558), .B(new_n5042_), .ZN(new_n33642_));
  NAND3_X1   g31206(.A1(new_n33639_), .A2(pi0513), .A3(new_n33642_), .ZN(new_n33643_));
  NOR2_X1    g31207(.A1(new_n33633_), .A2(pi0558), .ZN(new_n33644_));
  NOR2_X1    g31208(.A1(new_n33637_), .A2(new_n33346_), .ZN(new_n33645_));
  OAI21_X1   g31209(.A1(new_n33644_), .A2(new_n33645_), .B(new_n5042_), .ZN(new_n33646_));
  OAI21_X1   g31210(.A1(new_n33641_), .A2(new_n33346_), .B(pi0244), .ZN(new_n33647_));
  NAND3_X1   g31211(.A1(new_n33646_), .A2(new_n33214_), .A3(new_n33647_), .ZN(new_n33648_));
  AND2_X2    g31212(.A1(new_n33643_), .A2(new_n33648_), .Z(new_n33649_));
  NAND2_X1   g31213(.A1(new_n33649_), .A2(pi0509), .ZN(new_n33650_));
  XOR2_X1    g31214(.A1(pi0244), .A2(pi0513), .Z(new_n33651_));
  NOR2_X1    g31215(.A1(new_n33636_), .A2(new_n33651_), .ZN(new_n33652_));
  INV_X1     g31216(.I(new_n33652_), .ZN(new_n33653_));
  NAND2_X1   g31217(.A1(new_n33653_), .A2(new_n33200_), .ZN(new_n33654_));
  AOI21_X1   g31218(.A1(new_n33650_), .A2(new_n33654_), .B(new_n4881_), .ZN(new_n33655_));
  XOR2_X1    g31219(.A1(pi0244), .A2(pi0558), .Z(new_n33656_));
  NOR2_X1    g31220(.A1(new_n33641_), .A2(new_n33656_), .ZN(new_n33657_));
  AOI21_X1   g31221(.A1(new_n33657_), .A2(new_n33200_), .B(pi0245), .ZN(new_n33658_));
  NOR3_X1    g31222(.A1(new_n33655_), .A2(new_n33217_), .A3(new_n33658_), .ZN(new_n33659_));
  NAND2_X1   g31223(.A1(new_n33649_), .A2(new_n33200_), .ZN(new_n33660_));
  NAND2_X1   g31224(.A1(new_n33653_), .A2(pi0509), .ZN(new_n33661_));
  AOI21_X1   g31225(.A1(new_n33660_), .A2(new_n33661_), .B(pi0245), .ZN(new_n33662_));
  AOI21_X1   g31226(.A1(new_n33657_), .A2(pi0509), .B(new_n4881_), .ZN(new_n33663_));
  NOR3_X1    g31227(.A1(new_n33662_), .A2(pi0514), .A3(new_n33663_), .ZN(new_n33664_));
  NOR3_X1    g31228(.A1(new_n33659_), .A2(new_n33664_), .A3(new_n33197_), .ZN(new_n33665_));
  XOR2_X1    g31229(.A1(pi0245), .A2(pi0514), .Z(new_n33666_));
  NOR2_X1    g31230(.A1(new_n33653_), .A2(new_n33666_), .ZN(new_n33667_));
  NOR2_X1    g31231(.A1(new_n33667_), .A2(pi0508), .ZN(new_n33668_));
  OAI21_X1   g31232(.A1(new_n33665_), .A2(new_n33668_), .B(pi0247), .ZN(new_n33669_));
  XNOR2_X1   g31233(.A1(pi0245), .A2(pi0509), .ZN(new_n33670_));
  NAND2_X1   g31234(.A1(new_n33657_), .A2(new_n33670_), .ZN(new_n33671_));
  OAI21_X1   g31235(.A1(new_n33671_), .A2(pi0508), .B(new_n4339_), .ZN(new_n33672_));
  NAND3_X1   g31236(.A1(new_n33669_), .A2(pi0516), .A3(new_n33672_), .ZN(new_n33673_));
  NOR3_X1    g31237(.A1(new_n33659_), .A2(new_n33664_), .A3(pi0508), .ZN(new_n33674_));
  NOR2_X1    g31238(.A1(new_n33667_), .A2(new_n33197_), .ZN(new_n33675_));
  OAI21_X1   g31239(.A1(new_n33674_), .A2(new_n33675_), .B(new_n4339_), .ZN(new_n33676_));
  OAI21_X1   g31240(.A1(new_n33671_), .A2(new_n33197_), .B(pi0247), .ZN(new_n33677_));
  NAND3_X1   g31241(.A1(new_n33676_), .A2(new_n33223_), .A3(new_n33677_), .ZN(new_n33678_));
  AOI21_X1   g31242(.A1(new_n33673_), .A2(new_n33678_), .B(new_n3625_), .ZN(new_n33679_));
  XNOR2_X1   g31243(.A1(pi0247), .A2(pi0508), .ZN(new_n33680_));
  NAND3_X1   g31244(.A1(new_n33657_), .A2(new_n33670_), .A3(new_n33680_), .ZN(new_n33681_));
  AND2_X2    g31245(.A1(new_n33681_), .A2(pi0238), .Z(new_n33682_));
  XNOR2_X1   g31246(.A1(pi0247), .A2(pi0516), .ZN(new_n33683_));
  AOI21_X1   g31247(.A1(new_n33667_), .A2(new_n33683_), .B(pi0238), .ZN(new_n33684_));
  OAI21_X1   g31248(.A1(new_n33684_), .A2(new_n33682_), .B(new_n33226_), .ZN(new_n33685_));
  OAI21_X1   g31249(.A1(new_n33679_), .A2(new_n33226_), .B(new_n33685_), .ZN(new_n33686_));
  NAND2_X1   g31250(.A1(new_n33673_), .A2(new_n33678_), .ZN(new_n33687_));
  AOI21_X1   g31251(.A1(new_n33687_), .A2(new_n3625_), .B(pi0517), .ZN(new_n33688_));
  AND2_X2    g31252(.A1(new_n33681_), .A2(new_n3625_), .Z(new_n33689_));
  AOI21_X1   g31253(.A1(new_n33667_), .A2(new_n33683_), .B(new_n3625_), .ZN(new_n33690_));
  OAI21_X1   g31254(.A1(new_n33690_), .A2(new_n33689_), .B(pi0517), .ZN(new_n33691_));
  NAND2_X1   g31255(.A1(new_n33691_), .A2(new_n33194_), .ZN(new_n33692_));
  OAI22_X1   g31256(.A1(new_n33686_), .A2(new_n33194_), .B1(new_n33688_), .B2(new_n33692_), .ZN(new_n33693_));
  NAND2_X1   g31257(.A1(pi0248), .A2(pi0521), .ZN(new_n33694_));
  NAND2_X1   g31258(.A1(new_n4105_), .A2(new_n33239_), .ZN(new_n33695_));
  NAND2_X1   g31259(.A1(new_n4430_), .A2(new_n33236_), .ZN(new_n33696_));
  NAND2_X1   g31260(.A1(pi0246), .A2(pi0520), .ZN(new_n33697_));
  AOI22_X1   g31261(.A1(new_n33694_), .A2(new_n33695_), .B1(new_n33696_), .B2(new_n33697_), .ZN(new_n33698_));
  NAND2_X1   g31262(.A1(pi0249), .A2(pi0578), .ZN(new_n33699_));
  NAND2_X1   g31263(.A1(new_n3865_), .A2(new_n33471_), .ZN(new_n33700_));
  NAND2_X1   g31264(.A1(new_n3948_), .A2(new_n33460_), .ZN(new_n33701_));
  NAND2_X1   g31265(.A1(pi0241), .A2(pi0574), .ZN(new_n33702_));
  AOI22_X1   g31266(.A1(new_n33699_), .A2(new_n33700_), .B1(new_n33701_), .B2(new_n33702_), .ZN(new_n33703_));
  XNOR2_X1   g31267(.A1(pi0234), .A2(pi0518), .ZN(new_n33704_));
  NAND4_X1   g31268(.A1(new_n33208_), .A2(new_n33698_), .A3(new_n33703_), .A4(new_n33704_), .ZN(new_n33705_));
  OAI21_X1   g31269(.A1(new_n33705_), .A2(pi0582), .B(new_n4587_), .ZN(new_n33706_));
  XNOR2_X1   g31270(.A1(pi0249), .A2(pi0496), .ZN(new_n33707_));
  XNOR2_X1   g31271(.A1(pi0246), .A2(pi0499), .ZN(new_n33708_));
  XNOR2_X1   g31272(.A1(pi0248), .A2(pi0501), .ZN(new_n33709_));
  XNOR2_X1   g31273(.A1(pi0234), .A2(pi0505), .ZN(new_n33710_));
  NAND4_X1   g31274(.A1(new_n33707_), .A2(new_n33708_), .A3(new_n33709_), .A4(new_n33710_), .ZN(new_n33711_));
  XOR2_X1    g31275(.A1(pi0241), .A2(pi0500), .Z(new_n33712_));
  OR3_X2     g31276(.A1(new_n33184_), .A2(new_n33711_), .A3(new_n33712_), .Z(new_n33713_));
  NOR2_X1    g31277(.A1(new_n33713_), .A2(pi0542), .ZN(new_n33714_));
  OAI21_X1   g31278(.A1(new_n33705_), .A2(new_n33483_), .B(pi0240), .ZN(new_n33715_));
  NOR2_X1    g31279(.A1(new_n33713_), .A2(new_n33300_), .ZN(new_n33716_));
  OAI22_X1   g31280(.A1(new_n33706_), .A2(new_n33714_), .B1(new_n33715_), .B2(new_n33716_), .ZN(new_n33717_));
  NAND2_X1   g31281(.A1(new_n33717_), .A2(pi0497), .ZN(new_n33718_));
  INV_X1     g31282(.I(pi0497), .ZN(new_n33719_));
  XOR2_X1    g31283(.A1(pi0240), .A2(pi0582), .Z(new_n33720_));
  OAI21_X1   g31284(.A1(new_n33705_), .A2(new_n33720_), .B(new_n33719_), .ZN(new_n33721_));
  NAND2_X1   g31285(.A1(new_n33718_), .A2(new_n33721_), .ZN(new_n33722_));
  XOR2_X1    g31286(.A1(pi0240), .A2(pi0542), .Z(new_n33723_));
  NOR2_X1    g31287(.A1(new_n33713_), .A2(new_n33723_), .ZN(new_n33724_));
  AOI21_X1   g31288(.A1(new_n33724_), .A2(new_n33719_), .B(new_n3476_), .ZN(new_n33725_));
  AOI21_X1   g31289(.A1(new_n33722_), .A2(new_n3476_), .B(new_n33725_), .ZN(new_n33726_));
  NAND2_X1   g31290(.A1(new_n33717_), .A2(new_n33719_), .ZN(new_n33727_));
  OAI21_X1   g31291(.A1(new_n33705_), .A2(new_n33720_), .B(pi0497), .ZN(new_n33728_));
  NAND2_X1   g31292(.A1(new_n33727_), .A2(new_n33728_), .ZN(new_n33729_));
  AOI21_X1   g31293(.A1(new_n33724_), .A2(pi0497), .B(pi0239), .ZN(new_n33730_));
  AOI21_X1   g31294(.A1(new_n33729_), .A2(pi0239), .B(new_n33730_), .ZN(new_n33731_));
  MUX2_X1    g31295(.I0(new_n33731_), .I1(new_n33726_), .S(pi0519), .Z(new_n33732_));
  NOR2_X1    g31296(.A1(new_n33732_), .A2(new_n33291_), .ZN(new_n33733_));
  NOR2_X1    g31297(.A1(new_n33705_), .A2(new_n33720_), .ZN(new_n33734_));
  XOR2_X1    g31298(.A1(pi0239), .A2(pi0519), .Z(new_n33735_));
  NAND2_X1   g31299(.A1(new_n33734_), .A2(new_n33735_), .ZN(new_n33736_));
  INV_X1     g31300(.I(new_n33736_), .ZN(new_n33737_));
  NOR2_X1    g31301(.A1(new_n33737_), .A2(pi0539), .ZN(new_n33738_));
  OAI21_X1   g31302(.A1(new_n33733_), .A2(new_n33738_), .B(pi0242), .ZN(new_n33739_));
  XOR2_X1    g31303(.A1(pi0239), .A2(pi0497), .Z(new_n33740_));
  NAND2_X1   g31304(.A1(new_n33724_), .A2(new_n33740_), .ZN(new_n33741_));
  OAI21_X1   g31305(.A1(new_n33741_), .A2(pi0539), .B(new_n5143_), .ZN(new_n33742_));
  NAND3_X1   g31306(.A1(new_n33739_), .A2(pi0586), .A3(new_n33742_), .ZN(new_n33743_));
  NOR2_X1    g31307(.A1(new_n33732_), .A2(pi0539), .ZN(new_n33744_));
  NOR2_X1    g31308(.A1(new_n33737_), .A2(new_n33291_), .ZN(new_n33745_));
  OAI21_X1   g31309(.A1(new_n33744_), .A2(new_n33745_), .B(new_n5143_), .ZN(new_n33746_));
  OAI21_X1   g31310(.A1(new_n33741_), .A2(new_n33291_), .B(pi0242), .ZN(new_n33747_));
  NAND3_X1   g31311(.A1(new_n33746_), .A2(new_n33492_), .A3(new_n33747_), .ZN(new_n33748_));
  AND2_X2    g31312(.A1(new_n33743_), .A2(new_n33748_), .Z(new_n33749_));
  NAND2_X1   g31313(.A1(new_n33749_), .A2(pi0540), .ZN(new_n33750_));
  XOR2_X1    g31314(.A1(pi0242), .A2(pi0586), .Z(new_n33751_));
  NOR2_X1    g31315(.A1(new_n33736_), .A2(new_n33751_), .ZN(new_n33752_));
  INV_X1     g31316(.I(new_n33752_), .ZN(new_n33753_));
  NAND2_X1   g31317(.A1(new_n33753_), .A2(new_n33294_), .ZN(new_n33754_));
  AOI21_X1   g31318(.A1(new_n33750_), .A2(new_n33754_), .B(new_n3479_), .ZN(new_n33755_));
  XOR2_X1    g31319(.A1(pi0242), .A2(pi0539), .Z(new_n33756_));
  NOR2_X1    g31320(.A1(new_n33741_), .A2(new_n33756_), .ZN(new_n33757_));
  AOI21_X1   g31321(.A1(new_n33757_), .A2(new_n33294_), .B(pi0235), .ZN(new_n33758_));
  NOR3_X1    g31322(.A1(new_n33755_), .A2(new_n33480_), .A3(new_n33758_), .ZN(new_n33759_));
  NAND2_X1   g31323(.A1(new_n33749_), .A2(new_n33294_), .ZN(new_n33760_));
  NAND2_X1   g31324(.A1(new_n33753_), .A2(pi0540), .ZN(new_n33761_));
  AOI21_X1   g31325(.A1(new_n33760_), .A2(new_n33761_), .B(pi0235), .ZN(new_n33762_));
  AOI21_X1   g31326(.A1(new_n33757_), .A2(pi0540), .B(new_n3479_), .ZN(new_n33763_));
  NOR3_X1    g31327(.A1(new_n33762_), .A2(pi0581), .A3(new_n33763_), .ZN(new_n33764_));
  OR2_X2     g31328(.A1(new_n33759_), .A2(new_n33764_), .Z(new_n33765_));
  NOR2_X1    g31329(.A1(new_n33765_), .A2(new_n33489_), .ZN(new_n33766_));
  XNOR2_X1   g31330(.A1(pi0235), .A2(pi0540), .ZN(new_n33767_));
  NAND2_X1   g31331(.A1(new_n33757_), .A2(new_n33767_), .ZN(new_n33768_));
  INV_X1     g31332(.I(new_n33768_), .ZN(new_n33769_));
  NOR2_X1    g31333(.A1(new_n33769_), .A2(pi0585), .ZN(new_n33770_));
  OAI21_X1   g31334(.A1(new_n33766_), .A2(new_n33770_), .B(pi0244), .ZN(new_n33771_));
  XNOR2_X1   g31335(.A1(pi0235), .A2(pi0581), .ZN(new_n33772_));
  NAND2_X1   g31336(.A1(new_n33752_), .A2(new_n33772_), .ZN(new_n33773_));
  OAI21_X1   g31337(.A1(new_n33773_), .A2(pi0585), .B(new_n5042_), .ZN(new_n33774_));
  NAND3_X1   g31338(.A1(new_n33771_), .A2(pi0541), .A3(new_n33774_), .ZN(new_n33775_));
  NOR2_X1    g31339(.A1(new_n33765_), .A2(pi0585), .ZN(new_n33776_));
  NOR2_X1    g31340(.A1(new_n33769_), .A2(new_n33489_), .ZN(new_n33777_));
  OAI21_X1   g31341(.A1(new_n33776_), .A2(new_n33777_), .B(new_n5042_), .ZN(new_n33778_));
  OAI21_X1   g31342(.A1(new_n33773_), .A2(new_n33489_), .B(pi0244), .ZN(new_n33779_));
  NAND3_X1   g31343(.A1(new_n33778_), .A2(new_n33297_), .A3(new_n33779_), .ZN(new_n33780_));
  AND2_X2    g31344(.A1(new_n33775_), .A2(new_n33780_), .Z(new_n33781_));
  NAND2_X1   g31345(.A1(new_n33781_), .A2(pi0584), .ZN(new_n33782_));
  XOR2_X1    g31346(.A1(pi0244), .A2(pi0541), .Z(new_n33783_));
  NOR2_X1    g31347(.A1(new_n33768_), .A2(new_n33783_), .ZN(new_n33784_));
  INV_X1     g31348(.I(new_n33784_), .ZN(new_n33785_));
  NAND2_X1   g31349(.A1(new_n33785_), .A2(new_n33486_), .ZN(new_n33786_));
  AOI21_X1   g31350(.A1(new_n33782_), .A2(new_n33786_), .B(new_n4881_), .ZN(new_n33787_));
  XOR2_X1    g31351(.A1(pi0244), .A2(pi0585), .Z(new_n33788_));
  NOR2_X1    g31352(.A1(new_n33773_), .A2(new_n33788_), .ZN(new_n33789_));
  AOI21_X1   g31353(.A1(new_n33789_), .A2(new_n33486_), .B(pi0245), .ZN(new_n33790_));
  NOR3_X1    g31354(.A1(new_n33787_), .A2(new_n33175_), .A3(new_n33790_), .ZN(new_n33791_));
  NAND2_X1   g31355(.A1(new_n33781_), .A2(new_n33486_), .ZN(new_n33792_));
  NAND2_X1   g31356(.A1(new_n33785_), .A2(pi0584), .ZN(new_n33793_));
  AOI21_X1   g31357(.A1(new_n33792_), .A2(new_n33793_), .B(pi0245), .ZN(new_n33794_));
  AOI21_X1   g31358(.A1(new_n33789_), .A2(pi0584), .B(new_n4881_), .ZN(new_n33795_));
  NOR3_X1    g31359(.A1(new_n33794_), .A2(pi0503), .A3(new_n33795_), .ZN(new_n33796_));
  OR2_X2     g31360(.A1(new_n33791_), .A2(new_n33796_), .Z(new_n33797_));
  NAND2_X1   g31361(.A1(new_n33797_), .A2(pi0502), .ZN(new_n33798_));
  XNOR2_X1   g31362(.A1(pi0245), .A2(pi0584), .ZN(new_n33799_));
  NAND2_X1   g31363(.A1(new_n33789_), .A2(new_n33799_), .ZN(new_n33800_));
  INV_X1     g31364(.I(new_n33800_), .ZN(new_n33801_));
  NAND2_X1   g31365(.A1(new_n33801_), .A2(new_n33172_), .ZN(new_n33802_));
  AOI21_X1   g31366(.A1(new_n33798_), .A2(new_n33802_), .B(new_n33355_), .ZN(new_n33803_));
  XOR2_X1    g31367(.A1(pi0245), .A2(pi0503), .Z(new_n33804_));
  NOR2_X1    g31368(.A1(new_n33785_), .A2(new_n33804_), .ZN(new_n33805_));
  NAND3_X1   g31369(.A1(new_n33805_), .A2(pi0502), .A3(new_n33355_), .ZN(new_n33806_));
  NAND2_X1   g31370(.A1(new_n33806_), .A2(pi0247), .ZN(new_n33807_));
  NAND2_X1   g31371(.A1(new_n33801_), .A2(pi0502), .ZN(new_n33808_));
  NAND2_X1   g31372(.A1(new_n33797_), .A2(new_n33172_), .ZN(new_n33809_));
  AOI21_X1   g31373(.A1(new_n33809_), .A2(new_n33808_), .B(pi0561), .ZN(new_n33810_));
  NAND3_X1   g31374(.A1(new_n33805_), .A2(new_n33172_), .A3(pi0561), .ZN(new_n33811_));
  NAND2_X1   g31375(.A1(new_n33811_), .A2(new_n4339_), .ZN(new_n33812_));
  OAI22_X1   g31376(.A1(new_n33803_), .A2(new_n33807_), .B1(new_n33810_), .B2(new_n33812_), .ZN(new_n33813_));
  OAI21_X1   g31377(.A1(new_n33813_), .A2(new_n3625_), .B(pi0522), .ZN(new_n33814_));
  XNOR2_X1   g31378(.A1(pi0247), .A2(pi0502), .ZN(new_n33815_));
  AOI21_X1   g31379(.A1(new_n33805_), .A2(new_n33815_), .B(new_n3625_), .ZN(new_n33816_));
  XOR2_X1    g31380(.A1(pi0247), .A2(pi0561), .Z(new_n33817_));
  NOR2_X1    g31381(.A1(new_n33800_), .A2(new_n33817_), .ZN(new_n33818_));
  NOR2_X1    g31382(.A1(new_n33818_), .A2(pi0238), .ZN(new_n33819_));
  OAI21_X1   g31383(.A1(new_n33819_), .A2(new_n33816_), .B(new_n33242_), .ZN(new_n33820_));
  NAND3_X1   g31384(.A1(new_n33814_), .A2(pi0543), .A3(new_n33820_), .ZN(new_n33821_));
  OAI21_X1   g31385(.A1(new_n33813_), .A2(pi0238), .B(new_n33242_), .ZN(new_n33822_));
  NAND2_X1   g31386(.A1(new_n33805_), .A2(new_n33815_), .ZN(new_n33823_));
  NAND2_X1   g31387(.A1(new_n33823_), .A2(new_n3625_), .ZN(new_n33824_));
  OAI21_X1   g31388(.A1(new_n3625_), .A2(new_n33818_), .B(new_n33824_), .ZN(new_n33825_));
  AOI21_X1   g31389(.A1(new_n33825_), .A2(pi0522), .B(pi0543), .ZN(new_n33826_));
  NAND2_X1   g31390(.A1(new_n33822_), .A2(new_n33826_), .ZN(new_n33827_));
  NAND3_X1   g31391(.A1(new_n33821_), .A2(new_n33827_), .A3(new_n25326_), .ZN(new_n33828_));
  OAI21_X1   g31392(.A1(new_n33693_), .A2(new_n25326_), .B(new_n33828_), .ZN(new_n33829_));
  INV_X1     g31393(.I(new_n33208_), .ZN(new_n33830_));
  XNOR2_X1   g31394(.A1(pi0248), .A2(pi0576), .ZN(new_n33831_));
  XNOR2_X1   g31395(.A1(pi0246), .A2(pi0526), .ZN(new_n33832_));
  XNOR2_X1   g31396(.A1(pi0249), .A2(pi0528), .ZN(new_n33833_));
  XNOR2_X1   g31397(.A1(pi0234), .A2(pi0523), .ZN(new_n33834_));
  NAND4_X1   g31398(.A1(new_n33831_), .A2(new_n33832_), .A3(new_n33833_), .A4(new_n33834_), .ZN(new_n33835_));
  XOR2_X1    g31399(.A1(pi0241), .A2(pi0571), .Z(new_n33836_));
  NOR3_X1    g31400(.A1(new_n33830_), .A2(new_n33835_), .A3(new_n33836_), .ZN(new_n33837_));
  INV_X1     g31401(.I(new_n33837_), .ZN(new_n33838_));
  XOR2_X1    g31402(.A1(pi0248), .A2(pi0548), .Z(new_n33839_));
  XOR2_X1    g31403(.A1(pi0246), .A2(pi0546), .Z(new_n33840_));
  XOR2_X1    g31404(.A1(pi0249), .A2(pi0484), .Z(new_n33841_));
  XOR2_X1    g31405(.A1(pi0234), .A2(pi0544), .Z(new_n33842_));
  NOR4_X1    g31406(.A1(new_n33839_), .A2(new_n33840_), .A3(new_n33841_), .A4(new_n33842_), .ZN(new_n33843_));
  NAND2_X1   g31407(.A1(new_n33185_), .A2(new_n33843_), .ZN(new_n33844_));
  XOR2_X1    g31408(.A1(pi0241), .A2(pi0490), .Z(new_n33845_));
  OAI21_X1   g31409(.A1(new_n33844_), .A2(new_n33845_), .B(new_n33838_), .ZN(new_n33846_));
  XOR2_X1    g31410(.A1(pi0241), .A2(pi0490), .Z(new_n33847_));
  NOR2_X1    g31411(.A1(new_n33844_), .A2(new_n33847_), .ZN(new_n33848_));
  INV_X1     g31412(.I(new_n33848_), .ZN(new_n33849_));
  NOR2_X1    g31413(.A1(new_n33849_), .A2(pi0530), .ZN(new_n33850_));
  AOI21_X1   g31414(.A1(new_n33846_), .A2(pi0530), .B(new_n33850_), .ZN(new_n33851_));
  NOR2_X1    g31415(.A1(new_n33838_), .A2(new_n33265_), .ZN(new_n33852_));
  AOI21_X1   g31416(.A1(new_n33852_), .A2(new_n33148_), .B(new_n4587_), .ZN(new_n33853_));
  OAI21_X1   g31417(.A1(new_n33851_), .A2(new_n33148_), .B(new_n33853_), .ZN(new_n33854_));
  NOR2_X1    g31418(.A1(new_n33849_), .A2(new_n33265_), .ZN(new_n33855_));
  AOI21_X1   g31419(.A1(new_n33846_), .A2(new_n33265_), .B(new_n33855_), .ZN(new_n33856_));
  NOR2_X1    g31420(.A1(new_n33838_), .A2(new_n33148_), .ZN(new_n33857_));
  AOI21_X1   g31421(.A1(new_n33857_), .A2(new_n33265_), .B(pi0240), .ZN(new_n33858_));
  OAI21_X1   g31422(.A1(new_n33856_), .A2(pi0492), .B(new_n33858_), .ZN(new_n33859_));
  NAND2_X1   g31423(.A1(new_n33854_), .A2(new_n33859_), .ZN(new_n33860_));
  NAND2_X1   g31424(.A1(new_n33860_), .A2(pi0494), .ZN(new_n33861_));
  INV_X1     g31425(.I(pi0494), .ZN(new_n33862_));
  XOR2_X1    g31426(.A1(pi0240), .A2(pi0530), .Z(new_n33863_));
  NOR2_X1    g31427(.A1(new_n33838_), .A2(new_n33863_), .ZN(new_n33864_));
  INV_X1     g31428(.I(new_n33864_), .ZN(new_n33865_));
  NAND2_X1   g31429(.A1(new_n33865_), .A2(new_n33862_), .ZN(new_n33866_));
  NAND2_X1   g31430(.A1(new_n33861_), .A2(new_n33866_), .ZN(new_n33867_));
  XOR2_X1    g31431(.A1(pi0240), .A2(pi0492), .Z(new_n33868_));
  NOR2_X1    g31432(.A1(new_n33849_), .A2(new_n33868_), .ZN(new_n33869_));
  AOI21_X1   g31433(.A1(new_n33869_), .A2(new_n33862_), .B(new_n3476_), .ZN(new_n33870_));
  AOI21_X1   g31434(.A1(new_n33867_), .A2(new_n3476_), .B(new_n33870_), .ZN(new_n33871_));
  NAND2_X1   g31435(.A1(new_n33860_), .A2(new_n33862_), .ZN(new_n33872_));
  NAND2_X1   g31436(.A1(new_n33865_), .A2(pi0494), .ZN(new_n33873_));
  AOI21_X1   g31437(.A1(new_n33872_), .A2(new_n33873_), .B(new_n3476_), .ZN(new_n33874_));
  AOI21_X1   g31438(.A1(new_n33869_), .A2(pi0494), .B(pi0239), .ZN(new_n33875_));
  NOR3_X1    g31439(.A1(new_n33874_), .A2(pi0524), .A3(new_n33875_), .ZN(new_n33876_));
  AOI21_X1   g31440(.A1(pi0524), .A2(new_n33871_), .B(new_n33876_), .ZN(new_n33877_));
  NAND2_X1   g31441(.A1(new_n33877_), .A2(pi0483), .ZN(new_n33878_));
  XNOR2_X1   g31442(.A1(pi0239), .A2(pi0524), .ZN(new_n33879_));
  NOR2_X1    g31443(.A1(new_n33865_), .A2(new_n33879_), .ZN(new_n33880_));
  INV_X1     g31444(.I(new_n33880_), .ZN(new_n33881_));
  NAND2_X1   g31445(.A1(new_n33881_), .A2(new_n33124_), .ZN(new_n33882_));
  AOI21_X1   g31446(.A1(new_n33878_), .A2(new_n33882_), .B(new_n5143_), .ZN(new_n33883_));
  XNOR2_X1   g31447(.A1(pi0239), .A2(pi0494), .ZN(new_n33884_));
  NOR3_X1    g31448(.A1(new_n33849_), .A2(new_n33868_), .A3(new_n33884_), .ZN(new_n33885_));
  AOI21_X1   g31449(.A1(new_n33885_), .A2(new_n33124_), .B(pi0242), .ZN(new_n33886_));
  NOR3_X1    g31450(.A1(new_n33883_), .A2(new_n33457_), .A3(new_n33886_), .ZN(new_n33887_));
  NAND2_X1   g31451(.A1(new_n33877_), .A2(new_n33124_), .ZN(new_n33888_));
  NAND2_X1   g31452(.A1(new_n33881_), .A2(pi0483), .ZN(new_n33889_));
  AOI21_X1   g31453(.A1(new_n33888_), .A2(new_n33889_), .B(pi0242), .ZN(new_n33890_));
  AOI21_X1   g31454(.A1(new_n33885_), .A2(pi0483), .B(new_n5143_), .ZN(new_n33891_));
  NOR3_X1    g31455(.A1(new_n33890_), .A2(pi0573), .A3(new_n33891_), .ZN(new_n33892_));
  NOR2_X1    g31456(.A1(new_n33887_), .A2(new_n33892_), .ZN(new_n33893_));
  NAND2_X1   g31457(.A1(new_n33893_), .A2(pi0495), .ZN(new_n33894_));
  XOR2_X1    g31458(.A1(pi0242), .A2(pi0573), .Z(new_n33895_));
  NOR2_X1    g31459(.A1(new_n33881_), .A2(new_n33895_), .ZN(new_n33896_));
  INV_X1     g31460(.I(new_n33896_), .ZN(new_n33897_));
  NAND2_X1   g31461(.A1(new_n33897_), .A2(new_n33156_), .ZN(new_n33898_));
  AOI21_X1   g31462(.A1(new_n33894_), .A2(new_n33898_), .B(new_n3479_), .ZN(new_n33899_));
  XOR2_X1    g31463(.A1(pi0242), .A2(pi0483), .Z(new_n33900_));
  NOR4_X1    g31464(.A1(new_n33849_), .A2(new_n33868_), .A3(new_n33884_), .A4(new_n33900_), .ZN(new_n33901_));
  AOI21_X1   g31465(.A1(new_n33901_), .A2(new_n33156_), .B(pi0235), .ZN(new_n33902_));
  NOR3_X1    g31466(.A1(new_n33899_), .A2(new_n33463_), .A3(new_n33902_), .ZN(new_n33903_));
  NAND2_X1   g31467(.A1(new_n33893_), .A2(new_n33156_), .ZN(new_n33904_));
  NAND2_X1   g31468(.A1(new_n33897_), .A2(pi0495), .ZN(new_n33905_));
  AOI21_X1   g31469(.A1(new_n33904_), .A2(new_n33905_), .B(pi0235), .ZN(new_n33906_));
  AOI21_X1   g31470(.A1(new_n33901_), .A2(pi0495), .B(new_n3479_), .ZN(new_n33907_));
  NOR3_X1    g31471(.A1(new_n33906_), .A2(pi0575), .A3(new_n33907_), .ZN(new_n33908_));
  NOR2_X1    g31472(.A1(new_n33903_), .A2(new_n33908_), .ZN(new_n33909_));
  NAND2_X1   g31473(.A1(new_n33909_), .A2(pi0572), .ZN(new_n33910_));
  XNOR2_X1   g31474(.A1(pi0235), .A2(pi0495), .ZN(new_n33911_));
  NAND2_X1   g31475(.A1(new_n33901_), .A2(new_n33911_), .ZN(new_n33912_));
  NAND2_X1   g31476(.A1(new_n33912_), .A2(new_n33454_), .ZN(new_n33913_));
  AOI21_X1   g31477(.A1(new_n33910_), .A2(new_n33913_), .B(new_n5042_), .ZN(new_n33914_));
  XOR2_X1    g31478(.A1(pi0235), .A2(pi0575), .Z(new_n33915_));
  NOR2_X1    g31479(.A1(new_n33897_), .A2(new_n33915_), .ZN(new_n33916_));
  AOI21_X1   g31480(.A1(new_n33916_), .A2(new_n33454_), .B(pi0244), .ZN(new_n33917_));
  NOR3_X1    g31481(.A1(new_n33914_), .A2(new_n33151_), .A3(new_n33917_), .ZN(new_n33918_));
  NAND2_X1   g31482(.A1(new_n33909_), .A2(new_n33454_), .ZN(new_n33919_));
  NAND2_X1   g31483(.A1(new_n33912_), .A2(pi0572), .ZN(new_n33920_));
  AOI21_X1   g31484(.A1(new_n33919_), .A2(new_n33920_), .B(pi0244), .ZN(new_n33921_));
  AOI21_X1   g31485(.A1(new_n33916_), .A2(pi0572), .B(new_n5042_), .ZN(new_n33922_));
  NOR3_X1    g31486(.A1(new_n33921_), .A2(pi0493), .A3(new_n33922_), .ZN(new_n33923_));
  NOR2_X1    g31487(.A1(new_n33918_), .A2(new_n33923_), .ZN(new_n33924_));
  NAND2_X1   g31488(.A1(new_n33924_), .A2(pi0545), .ZN(new_n33925_));
  XOR2_X1    g31489(.A1(pi0244), .A2(pi0572), .Z(new_n33926_));
  NOR3_X1    g31490(.A1(new_n33897_), .A2(new_n33915_), .A3(new_n33926_), .ZN(new_n33927_));
  INV_X1     g31491(.I(new_n33927_), .ZN(new_n33928_));
  NAND2_X1   g31492(.A1(new_n33928_), .A2(new_n33309_), .ZN(new_n33929_));
  AOI21_X1   g31493(.A1(new_n33925_), .A2(new_n33929_), .B(new_n4881_), .ZN(new_n33930_));
  XOR2_X1    g31494(.A1(pi0244), .A2(pi0493), .Z(new_n33931_));
  NOR2_X1    g31495(.A1(new_n33912_), .A2(new_n33931_), .ZN(new_n33932_));
  AOI21_X1   g31496(.A1(new_n33932_), .A2(new_n33309_), .B(pi0245), .ZN(new_n33933_));
  NOR3_X1    g31497(.A1(new_n33930_), .A2(new_n33252_), .A3(new_n33933_), .ZN(new_n33934_));
  NAND2_X1   g31498(.A1(new_n33924_), .A2(new_n33309_), .ZN(new_n33935_));
  NAND2_X1   g31499(.A1(new_n33928_), .A2(pi0545), .ZN(new_n33936_));
  AOI21_X1   g31500(.A1(new_n33935_), .A2(new_n33936_), .B(pi0245), .ZN(new_n33937_));
  AOI21_X1   g31501(.A1(new_n33932_), .A2(pi0545), .B(new_n4881_), .ZN(new_n33938_));
  NOR3_X1    g31502(.A1(new_n33937_), .A2(pi0525), .A3(new_n33938_), .ZN(new_n33939_));
  NOR2_X1    g31503(.A1(new_n33934_), .A2(new_n33939_), .ZN(new_n33940_));
  NAND2_X1   g31504(.A1(new_n33940_), .A2(pi0547), .ZN(new_n33941_));
  XOR2_X1    g31505(.A1(pi0245), .A2(pi0525), .Z(new_n33942_));
  NOR2_X1    g31506(.A1(new_n33928_), .A2(new_n33942_), .ZN(new_n33943_));
  INV_X1     g31507(.I(new_n33943_), .ZN(new_n33944_));
  NAND2_X1   g31508(.A1(new_n33944_), .A2(new_n33314_), .ZN(new_n33945_));
  AOI21_X1   g31509(.A1(new_n33941_), .A2(new_n33945_), .B(new_n4339_), .ZN(new_n33946_));
  XOR2_X1    g31510(.A1(pi0245), .A2(pi0545), .Z(new_n33947_));
  NOR3_X1    g31511(.A1(new_n33912_), .A2(new_n33931_), .A3(new_n33947_), .ZN(new_n33948_));
  AOI21_X1   g31512(.A1(new_n33948_), .A2(new_n33314_), .B(pi0247), .ZN(new_n33949_));
  NOR3_X1    g31513(.A1(new_n33946_), .A2(new_n33257_), .A3(new_n33949_), .ZN(new_n33950_));
  NAND2_X1   g31514(.A1(new_n33940_), .A2(new_n33314_), .ZN(new_n33951_));
  NAND2_X1   g31515(.A1(new_n33944_), .A2(pi0547), .ZN(new_n33952_));
  AOI21_X1   g31516(.A1(new_n33951_), .A2(new_n33952_), .B(pi0247), .ZN(new_n33953_));
  AOI21_X1   g31517(.A1(new_n33948_), .A2(pi0547), .B(new_n4339_), .ZN(new_n33954_));
  NOR3_X1    g31518(.A1(new_n33953_), .A2(pi0527), .A3(new_n33954_), .ZN(new_n33955_));
  NOR2_X1    g31519(.A1(new_n33950_), .A2(new_n33955_), .ZN(new_n33956_));
  OAI21_X1   g31520(.A1(new_n33956_), .A2(new_n3625_), .B(pi0529), .ZN(new_n33957_));
  XNOR2_X1   g31521(.A1(pi0247), .A2(pi0547), .ZN(new_n33958_));
  AOI21_X1   g31522(.A1(new_n33948_), .A2(new_n33958_), .B(new_n3625_), .ZN(new_n33959_));
  XNOR2_X1   g31523(.A1(pi0247), .A2(pi0527), .ZN(new_n33960_));
  AOI21_X1   g31524(.A1(new_n33943_), .A2(new_n33960_), .B(pi0238), .ZN(new_n33961_));
  OAI21_X1   g31525(.A1(new_n33961_), .A2(new_n33959_), .B(new_n33262_), .ZN(new_n33962_));
  NAND3_X1   g31526(.A1(new_n33957_), .A2(pi0491), .A3(new_n33962_), .ZN(new_n33963_));
  OAI21_X1   g31527(.A1(new_n33956_), .A2(pi0238), .B(new_n33262_), .ZN(new_n33964_));
  AOI21_X1   g31528(.A1(new_n33948_), .A2(new_n33958_), .B(pi0238), .ZN(new_n33965_));
  AOI21_X1   g31529(.A1(new_n33943_), .A2(new_n33960_), .B(new_n3625_), .ZN(new_n33966_));
  OR2_X2     g31530(.A1(new_n33966_), .A2(new_n33965_), .Z(new_n33967_));
  AOI21_X1   g31531(.A1(new_n33967_), .A2(pi0529), .B(pi0491), .ZN(new_n33968_));
  NAND2_X1   g31532(.A1(new_n33964_), .A2(new_n33968_), .ZN(new_n33969_));
  NAND3_X1   g31533(.A1(new_n33963_), .A2(new_n33969_), .A3(pi0233), .ZN(new_n33970_));
  NOR2_X1    g31534(.A1(new_n3865_), .A2(new_n33336_), .ZN(new_n33971_));
  NOR2_X1    g31535(.A1(pi0249), .A2(pi0555), .ZN(new_n33972_));
  NOR2_X1    g31536(.A1(pi0241), .A2(pi0553), .ZN(new_n33973_));
  NOR2_X1    g31537(.A1(new_n3948_), .A2(new_n33330_), .ZN(new_n33974_));
  OAI22_X1   g31538(.A1(new_n33971_), .A2(new_n33972_), .B1(new_n33974_), .B2(new_n33973_), .ZN(new_n33975_));
  NOR2_X1    g31539(.A1(new_n4105_), .A2(new_n33333_), .ZN(new_n33976_));
  NOR2_X1    g31540(.A1(pi0248), .A2(pi0554), .ZN(new_n33977_));
  NOR2_X1    g31541(.A1(pi0246), .A2(pi0563), .ZN(new_n33978_));
  NOR2_X1    g31542(.A1(new_n4430_), .A2(new_n33360_), .ZN(new_n33979_));
  OAI22_X1   g31543(.A1(new_n33976_), .A2(new_n33977_), .B1(new_n33979_), .B2(new_n33978_), .ZN(new_n33980_));
  XOR2_X1    g31544(.A1(pi0240), .A2(pi0551), .Z(new_n33981_));
  XOR2_X1    g31545(.A1(pi0234), .A2(pi0485), .Z(new_n33982_));
  NOR4_X1    g31546(.A1(new_n33975_), .A2(new_n33980_), .A3(new_n33981_), .A4(new_n33982_), .ZN(new_n33983_));
  NAND2_X1   g31547(.A1(new_n33185_), .A2(new_n33983_), .ZN(new_n33984_));
  XNOR2_X1   g31548(.A1(pi0239), .A2(pi0550), .ZN(new_n33985_));
  NOR2_X1    g31549(.A1(new_n33984_), .A2(new_n33985_), .ZN(new_n33986_));
  AOI22_X1   g31550(.A1(new_n4430_), .A2(pi0564), .B1(new_n3865_), .B2(pi0482), .ZN(new_n33987_));
  OAI21_X1   g31551(.A1(new_n3865_), .A2(pi0482), .B(new_n33987_), .ZN(new_n33988_));
  XOR2_X1    g31552(.A1(pi0241), .A2(pi0562), .Z(new_n33989_));
  XOR2_X1    g31553(.A1(pi0234), .A2(pi0570), .Z(new_n33990_));
  NOR3_X1    g31554(.A1(new_n33988_), .A2(new_n33989_), .A3(new_n33990_), .ZN(new_n33991_));
  NAND2_X1   g31555(.A1(new_n33208_), .A2(new_n33991_), .ZN(new_n33992_));
  XNOR2_X1   g31556(.A1(pi0248), .A2(pi0565), .ZN(new_n33993_));
  NAND2_X1   g31557(.A1(new_n33352_), .A2(pi0240), .ZN(new_n33994_));
  AOI22_X1   g31558(.A1(new_n4587_), .A2(pi0560), .B1(new_n33363_), .B2(pi0246), .ZN(new_n33995_));
  NAND3_X1   g31559(.A1(new_n33993_), .A2(new_n33994_), .A3(new_n33995_), .ZN(new_n33996_));
  NOR2_X1    g31560(.A1(new_n33992_), .A2(new_n33996_), .ZN(new_n33997_));
  NOR2_X1    g31561(.A1(new_n3476_), .A2(pi0569), .ZN(new_n33998_));
  AOI21_X1   g31562(.A1(new_n33997_), .A2(new_n33998_), .B(new_n33986_), .ZN(new_n33999_));
  NOR2_X1    g31563(.A1(new_n33984_), .A2(pi0550), .ZN(new_n34000_));
  NOR2_X1    g31564(.A1(new_n34000_), .A2(new_n3476_), .ZN(new_n34001_));
  NAND2_X1   g31565(.A1(new_n33997_), .A2(new_n4587_), .ZN(new_n34002_));
  NAND2_X1   g31566(.A1(new_n33363_), .A2(pi0246), .ZN(new_n34003_));
  NAND4_X1   g31567(.A1(new_n33993_), .A2(pi0240), .A3(pi0560), .A4(new_n34003_), .ZN(new_n34004_));
  OAI21_X1   g31568(.A1(new_n33992_), .A2(new_n34004_), .B(new_n34002_), .ZN(new_n34005_));
  NAND2_X1   g31569(.A1(new_n34005_), .A2(pi0569), .ZN(new_n34006_));
  OAI21_X1   g31570(.A1(new_n34006_), .A2(new_n34001_), .B(new_n33999_), .ZN(new_n34007_));
  XOR2_X1    g31571(.A1(pi0239), .A2(pi0569), .Z(new_n34008_));
  NAND2_X1   g31572(.A1(new_n34005_), .A2(new_n34008_), .ZN(new_n34009_));
  NOR2_X1    g31573(.A1(new_n34009_), .A2(pi0489), .ZN(new_n34010_));
  AOI21_X1   g31574(.A1(new_n34007_), .A2(pi0489), .B(new_n34010_), .ZN(new_n34011_));
  INV_X1     g31575(.I(new_n33986_), .ZN(new_n34012_));
  NOR2_X1    g31576(.A1(new_n34012_), .A2(new_n33141_), .ZN(new_n34013_));
  AOI21_X1   g31577(.A1(new_n34013_), .A2(new_n33339_), .B(new_n5143_), .ZN(new_n34014_));
  OAI21_X1   g31578(.A1(new_n34011_), .A2(new_n33339_), .B(new_n34014_), .ZN(new_n34015_));
  NOR2_X1    g31579(.A1(new_n34009_), .A2(new_n33141_), .ZN(new_n34016_));
  AOI21_X1   g31580(.A1(new_n34007_), .A2(new_n33141_), .B(new_n34016_), .ZN(new_n34017_));
  NOR2_X1    g31581(.A1(new_n34012_), .A2(new_n33339_), .ZN(new_n34018_));
  AOI21_X1   g31582(.A1(new_n34018_), .A2(new_n33141_), .B(pi0242), .ZN(new_n34019_));
  OAI21_X1   g31583(.A1(new_n34017_), .A2(pi0556), .B(new_n34019_), .ZN(new_n34020_));
  NAND2_X1   g31584(.A1(new_n34015_), .A2(new_n34020_), .ZN(new_n34021_));
  NAND2_X1   g31585(.A1(new_n34021_), .A2(pi0549), .ZN(new_n34022_));
  XOR2_X1    g31586(.A1(pi0242), .A2(pi0556), .Z(new_n34023_));
  NOR2_X1    g31587(.A1(new_n34009_), .A2(new_n34023_), .ZN(new_n34024_));
  INV_X1     g31588(.I(new_n34024_), .ZN(new_n34025_));
  NAND2_X1   g31589(.A1(new_n34025_), .A2(new_n33319_), .ZN(new_n34026_));
  AOI21_X1   g31590(.A1(new_n34022_), .A2(new_n34026_), .B(new_n3479_), .ZN(new_n34027_));
  XOR2_X1    g31591(.A1(pi0242), .A2(pi0489), .Z(new_n34028_));
  NOR2_X1    g31592(.A1(new_n34012_), .A2(new_n34028_), .ZN(new_n34029_));
  AOI21_X1   g31593(.A1(new_n34029_), .A2(new_n33319_), .B(pi0235), .ZN(new_n34030_));
  NOR3_X1    g31594(.A1(new_n34027_), .A2(new_n33268_), .A3(new_n34030_), .ZN(new_n34031_));
  NAND2_X1   g31595(.A1(new_n34021_), .A2(new_n33319_), .ZN(new_n34032_));
  NAND2_X1   g31596(.A1(new_n34025_), .A2(pi0549), .ZN(new_n34033_));
  AOI21_X1   g31597(.A1(new_n34032_), .A2(new_n34033_), .B(pi0235), .ZN(new_n34034_));
  AOI21_X1   g31598(.A1(new_n34029_), .A2(pi0549), .B(new_n3479_), .ZN(new_n34035_));
  NOR3_X1    g31599(.A1(new_n34034_), .A2(pi0531), .A3(new_n34035_), .ZN(new_n34036_));
  NOR2_X1    g31600(.A1(new_n34031_), .A2(new_n34036_), .ZN(new_n34037_));
  NAND2_X1   g31601(.A1(new_n34037_), .A2(pi0486), .ZN(new_n34038_));
  XNOR2_X1   g31602(.A1(pi0235), .A2(pi0531), .ZN(new_n34039_));
  NAND2_X1   g31603(.A1(new_n34024_), .A2(new_n34039_), .ZN(new_n34040_));
  NAND2_X1   g31604(.A1(new_n34040_), .A2(new_n33133_), .ZN(new_n34041_));
  AOI21_X1   g31605(.A1(new_n34038_), .A2(new_n34041_), .B(new_n5042_), .ZN(new_n34042_));
  XOR2_X1    g31606(.A1(pi0235), .A2(pi0549), .Z(new_n34043_));
  NOR3_X1    g31607(.A1(new_n34012_), .A2(new_n34028_), .A3(new_n34043_), .ZN(new_n34044_));
  AOI21_X1   g31608(.A1(new_n34044_), .A2(new_n33133_), .B(pi0244), .ZN(new_n34045_));
  NOR3_X1    g31609(.A1(new_n34042_), .A2(new_n33368_), .A3(new_n34045_), .ZN(new_n34046_));
  NAND2_X1   g31610(.A1(new_n34037_), .A2(new_n33133_), .ZN(new_n34047_));
  NAND2_X1   g31611(.A1(new_n34040_), .A2(pi0486), .ZN(new_n34048_));
  AOI21_X1   g31612(.A1(new_n34047_), .A2(new_n34048_), .B(pi0244), .ZN(new_n34049_));
  AOI21_X1   g31613(.A1(new_n34044_), .A2(pi0486), .B(new_n5042_), .ZN(new_n34050_));
  NOR3_X1    g31614(.A1(new_n34049_), .A2(pi0566), .A3(new_n34050_), .ZN(new_n34051_));
  NOR2_X1    g31615(.A1(new_n34046_), .A2(new_n34051_), .ZN(new_n34052_));
  NAND2_X1   g31616(.A1(new_n34052_), .A2(pi0568), .ZN(new_n34053_));
  XOR2_X1    g31617(.A1(pi0244), .A2(pi0486), .Z(new_n34054_));
  NOR4_X1    g31618(.A1(new_n34012_), .A2(new_n34028_), .A3(new_n34043_), .A4(new_n34054_), .ZN(new_n34055_));
  INV_X1     g31619(.I(new_n34055_), .ZN(new_n34056_));
  NAND2_X1   g31620(.A1(new_n34056_), .A2(new_n33443_), .ZN(new_n34057_));
  AOI21_X1   g31621(.A1(new_n34053_), .A2(new_n34057_), .B(new_n4881_), .ZN(new_n34058_));
  XOR2_X1    g31622(.A1(pi0244), .A2(pi0566), .Z(new_n34059_));
  NOR2_X1    g31623(.A1(new_n34040_), .A2(new_n34059_), .ZN(new_n34060_));
  AOI21_X1   g31624(.A1(new_n34060_), .A2(new_n33443_), .B(pi0245), .ZN(new_n34061_));
  NOR3_X1    g31625(.A1(new_n34058_), .A2(new_n33477_), .A3(new_n34061_), .ZN(new_n34062_));
  NAND2_X1   g31626(.A1(new_n34052_), .A2(new_n33443_), .ZN(new_n34063_));
  NAND2_X1   g31627(.A1(new_n34056_), .A2(pi0568), .ZN(new_n34064_));
  AOI21_X1   g31628(.A1(new_n34063_), .A2(new_n34064_), .B(pi0245), .ZN(new_n34065_));
  AOI21_X1   g31629(.A1(new_n34060_), .A2(pi0568), .B(new_n4881_), .ZN(new_n34066_));
  NOR3_X1    g31630(.A1(new_n34065_), .A2(pi0580), .A3(new_n34066_), .ZN(new_n34067_));
  NOR2_X1    g31631(.A1(new_n34062_), .A2(new_n34067_), .ZN(new_n34068_));
  NAND2_X1   g31632(.A1(new_n34068_), .A2(pi0552), .ZN(new_n34069_));
  XNOR2_X1   g31633(.A1(pi0245), .A2(pi0568), .ZN(new_n34070_));
  NAND2_X1   g31634(.A1(new_n34060_), .A2(new_n34070_), .ZN(new_n34071_));
  NAND2_X1   g31635(.A1(new_n34071_), .A2(new_n33327_), .ZN(new_n34072_));
  AOI21_X1   g31636(.A1(new_n34069_), .A2(new_n34072_), .B(new_n4339_), .ZN(new_n34073_));
  XOR2_X1    g31637(.A1(pi0245), .A2(pi0580), .Z(new_n34074_));
  NOR2_X1    g31638(.A1(new_n34056_), .A2(new_n34074_), .ZN(new_n34075_));
  AOI21_X1   g31639(.A1(new_n34075_), .A2(new_n33327_), .B(pi0247), .ZN(new_n34076_));
  NOR3_X1    g31640(.A1(new_n34073_), .A2(new_n33271_), .A3(new_n34076_), .ZN(new_n34077_));
  NAND2_X1   g31641(.A1(new_n34068_), .A2(new_n33327_), .ZN(new_n34078_));
  NAND2_X1   g31642(.A1(new_n34071_), .A2(pi0552), .ZN(new_n34079_));
  AOI21_X1   g31643(.A1(new_n34078_), .A2(new_n34079_), .B(pi0247), .ZN(new_n34080_));
  AOI21_X1   g31644(.A1(new_n34075_), .A2(pi0552), .B(new_n4339_), .ZN(new_n34081_));
  NOR3_X1    g31645(.A1(new_n34080_), .A2(pi0532), .A3(new_n34081_), .ZN(new_n34082_));
  NOR2_X1    g31646(.A1(new_n34077_), .A2(new_n34082_), .ZN(new_n34083_));
  OAI21_X1   g31647(.A1(new_n34083_), .A2(new_n3625_), .B(pi0577), .ZN(new_n34084_));
  XOR2_X1    g31648(.A1(pi0247), .A2(pi0532), .Z(new_n34085_));
  NOR2_X1    g31649(.A1(new_n34071_), .A2(new_n34085_), .ZN(new_n34086_));
  XNOR2_X1   g31650(.A1(pi0247), .A2(pi0552), .ZN(new_n34087_));
  NAND2_X1   g31651(.A1(new_n34075_), .A2(new_n34087_), .ZN(new_n34088_));
  NAND2_X1   g31652(.A1(new_n34088_), .A2(new_n3625_), .ZN(new_n34089_));
  OAI21_X1   g31653(.A1(new_n34086_), .A2(new_n3625_), .B(new_n34089_), .ZN(new_n34090_));
  NAND2_X1   g31654(.A1(new_n34090_), .A2(new_n33468_), .ZN(new_n34091_));
  NAND3_X1   g31655(.A1(new_n34084_), .A2(pi0498), .A3(new_n34091_), .ZN(new_n34092_));
  OAI21_X1   g31656(.A1(new_n34083_), .A2(pi0238), .B(new_n33468_), .ZN(new_n34093_));
  NAND2_X1   g31657(.A1(new_n34088_), .A2(pi0238), .ZN(new_n34094_));
  OAI21_X1   g31658(.A1(new_n34086_), .A2(pi0238), .B(new_n34094_), .ZN(new_n34095_));
  AOI21_X1   g31659(.A1(new_n34095_), .A2(pi0577), .B(pi0498), .ZN(new_n34096_));
  NAND2_X1   g31660(.A1(new_n34093_), .A2(new_n34096_), .ZN(new_n34097_));
  NAND3_X1   g31661(.A1(new_n34092_), .A2(new_n34097_), .A3(new_n25326_), .ZN(new_n34098_));
  AOI21_X1   g31662(.A1(new_n33970_), .A2(new_n34098_), .B(pi0237), .ZN(new_n34099_));
  AOI21_X1   g31663(.A1(new_n33829_), .A2(pi0237), .B(new_n34099_), .ZN(po0750));
  NOR2_X1    g31664(.A1(new_n32942_), .A2(pi0806), .ZN(new_n34101_));
  NOR2_X1    g31665(.A1(pi0332), .A2(pi0806), .ZN(new_n34102_));
  NAND3_X1   g31666(.A1(new_n34102_), .A2(pi0600), .A3(pi0990), .ZN(new_n34103_));
  NAND2_X1   g31667(.A1(new_n2630_), .A2(pi0594), .ZN(new_n34104_));
  AOI21_X1   g31668(.A1(new_n34103_), .A2(new_n34104_), .B(new_n34101_), .ZN(po0751));
  INV_X1     g31669(.I(pi0605), .ZN(new_n34106_));
  NOR3_X1    g31670(.A1(new_n32954_), .A2(new_n34106_), .A3(pi0806), .ZN(new_n34107_));
  XOR2_X1    g31671(.A1(new_n34107_), .A2(new_n32948_), .Z(new_n34108_));
  NOR2_X1    g31672(.A1(new_n34108_), .A2(pi0332), .ZN(po0752));
  NAND4_X1   g31673(.A1(new_n32943_), .A2(pi0595), .A3(pi0597), .A4(new_n34102_), .ZN(new_n34110_));
  NOR2_X1    g31674(.A1(new_n34110_), .A2(new_n32950_), .ZN(new_n34111_));
  NAND2_X1   g31675(.A1(new_n2630_), .A2(pi0596), .ZN(new_n34112_));
  AOI21_X1   g31676(.A1(new_n34110_), .A2(new_n34112_), .B(new_n34111_), .ZN(po0753));
  OAI21_X1   g31677(.A1(new_n32942_), .A2(pi0806), .B(pi0597), .ZN(new_n34114_));
  INV_X1     g31678(.I(pi0597), .ZN(new_n34115_));
  NAND2_X1   g31679(.A1(new_n34101_), .A2(new_n34115_), .ZN(new_n34116_));
  AOI21_X1   g31680(.A1(new_n34116_), .A2(new_n34114_), .B(pi0332), .ZN(po0754));
  INV_X1     g31681(.I(pi0598), .ZN(new_n34118_));
  OR2_X2     g31682(.A1(po1038), .A2(pi0882), .Z(new_n34119_));
  NOR2_X1    g31683(.A1(new_n34119_), .A2(new_n5692_), .ZN(new_n34120_));
  NAND2_X1   g31684(.A1(pi0740), .A2(pi0780), .ZN(new_n34121_));
  OAI22_X1   g31685(.A1(new_n34120_), .A2(new_n34118_), .B1(new_n5409_), .B2(new_n34121_), .ZN(po0755));
  INV_X1     g31686(.I(new_n34111_), .ZN(new_n34123_));
  NAND3_X1   g31687(.A1(new_n34123_), .A2(new_n2630_), .A3(pi0599), .ZN(new_n34124_));
  OAI21_X1   g31688(.A1(pi0599), .A2(new_n34123_), .B(new_n34124_), .ZN(po0756));
  INV_X1     g31689(.I(pi0806), .ZN(new_n34126_));
  AOI21_X1   g31690(.A1(new_n34126_), .A2(pi0990), .B(pi0600), .ZN(new_n34127_));
  AND3_X2    g31691(.A1(new_n34126_), .A2(pi0600), .A3(pi0990), .Z(new_n34128_));
  NOR3_X1    g31692(.A1(new_n34128_), .A2(new_n34127_), .A3(pi0332), .ZN(po0757));
  NAND2_X1   g31693(.A1(pi0601), .A2(pi0806), .ZN(new_n34130_));
  NAND2_X1   g31694(.A1(new_n34126_), .A2(pi0989), .ZN(new_n34131_));
  AOI21_X1   g31695(.A1(new_n34131_), .A2(new_n34130_), .B(pi0332), .ZN(po0758));
  NAND2_X1   g31696(.A1(new_n12740_), .A2(pi1160), .ZN(new_n34133_));
  NAND2_X1   g31697(.A1(new_n12739_), .A2(pi0715), .ZN(new_n34134_));
  AOI21_X1   g31698(.A1(new_n34133_), .A2(new_n34134_), .B(new_n13000_), .ZN(new_n34135_));
  NOR3_X1    g31699(.A1(new_n14300_), .A2(new_n14285_), .A3(new_n34135_), .ZN(new_n34136_));
  NAND4_X1   g31700(.A1(new_n34136_), .A2(pi0230), .A3(new_n12824_), .A4(new_n12952_), .ZN(new_n34137_));
  OAI22_X1   g31701(.A1(new_n14292_), .A2(new_n34137_), .B1(pi0230), .B2(new_n5486_), .ZN(po0759));
  INV_X1     g31702(.I(pi0966), .ZN(new_n34139_));
  INV_X1     g31703(.I(pi1061), .ZN(new_n34140_));
  INV_X1     g31704(.I(pi1038), .ZN(new_n34141_));
  INV_X1     g31705(.I(pi1060), .ZN(new_n34142_));
  NOR3_X1    g31706(.A1(new_n34141_), .A2(new_n34142_), .A3(pi0980), .ZN(new_n34143_));
  NAND3_X1   g31707(.A1(new_n34143_), .A2(pi0952), .A3(new_n34140_), .ZN(new_n34144_));
  NOR3_X1    g31708(.A1(new_n34144_), .A2(new_n12738_), .A3(pi1100), .ZN(new_n34145_));
  NOR2_X1    g31709(.A1(new_n34144_), .A2(new_n12738_), .ZN(po0897));
  OAI21_X1   g31710(.A1(po0897), .A2(pi0603), .B(new_n34139_), .ZN(new_n34147_));
  NOR2_X1    g31711(.A1(pi0871), .A2(pi0872), .ZN(new_n34148_));
  OAI22_X1   g31712(.A1(new_n34147_), .A2(new_n34145_), .B1(new_n34139_), .B2(new_n34148_), .ZN(po0760));
  AND2_X2    g31713(.A1(new_n13118_), .A2(pi0823), .Z(new_n34150_));
  INV_X1     g31714(.I(pi0779), .ZN(new_n34151_));
  NAND2_X1   g31715(.A1(new_n34150_), .A2(new_n34151_), .ZN(new_n34152_));
  NAND2_X1   g31716(.A1(new_n2628_), .A2(pi0983), .ZN(new_n34153_));
  OAI21_X1   g31717(.A1(new_n34153_), .A2(new_n5473_), .B(pi0604), .ZN(new_n34154_));
  OAI21_X1   g31718(.A1(new_n34150_), .A2(new_n34154_), .B(new_n34152_), .ZN(po0761));
  NAND2_X1   g31719(.A1(new_n34106_), .A2(new_n34126_), .ZN(new_n34156_));
  NAND2_X1   g31720(.A1(pi0605), .A2(pi0806), .ZN(new_n34157_));
  AOI21_X1   g31721(.A1(new_n34156_), .A2(new_n34157_), .B(pi0332), .ZN(po0762));
  NAND2_X1   g31722(.A1(pi0837), .A2(pi0966), .ZN(new_n34159_));
  NOR2_X1    g31723(.A1(po0897), .A2(new_n25131_), .ZN(new_n34160_));
  AOI21_X1   g31724(.A1(pi1104), .A2(po0897), .B(new_n34160_), .ZN(new_n34161_));
  OAI21_X1   g31725(.A1(new_n34161_), .A2(pi0966), .B(new_n34159_), .ZN(po0763));
  NAND2_X1   g31726(.A1(po0897), .A2(pi1107), .ZN(new_n34163_));
  INV_X1     g31727(.I(po0897), .ZN(new_n34164_));
  NAND2_X1   g31728(.A1(new_n34164_), .A2(pi0607), .ZN(new_n34165_));
  AOI21_X1   g31729(.A1(new_n34165_), .A2(new_n34163_), .B(pi0966), .ZN(po0764));
  NAND2_X1   g31730(.A1(po0897), .A2(pi1116), .ZN(new_n34167_));
  NAND2_X1   g31731(.A1(new_n34164_), .A2(pi0608), .ZN(new_n34168_));
  AOI21_X1   g31732(.A1(new_n34168_), .A2(new_n34167_), .B(pi0966), .ZN(po0765));
  NAND2_X1   g31733(.A1(po0897), .A2(pi1118), .ZN(new_n34170_));
  NAND2_X1   g31734(.A1(new_n34164_), .A2(pi0609), .ZN(new_n34171_));
  AOI21_X1   g31735(.A1(new_n34171_), .A2(new_n34170_), .B(pi0966), .ZN(po0766));
  NAND2_X1   g31736(.A1(po0897), .A2(pi1113), .ZN(new_n34173_));
  NAND2_X1   g31737(.A1(new_n34164_), .A2(pi0610), .ZN(new_n34174_));
  AOI21_X1   g31738(.A1(new_n34174_), .A2(new_n34173_), .B(pi0966), .ZN(po0767));
  NAND2_X1   g31739(.A1(po0897), .A2(pi1114), .ZN(new_n34176_));
  NAND2_X1   g31740(.A1(new_n34164_), .A2(pi0611), .ZN(new_n34177_));
  AOI21_X1   g31741(.A1(new_n34177_), .A2(new_n34176_), .B(pi0966), .ZN(po0768));
  NAND2_X1   g31742(.A1(po0897), .A2(pi1111), .ZN(new_n34179_));
  NAND2_X1   g31743(.A1(new_n34164_), .A2(pi0612), .ZN(new_n34180_));
  AOI21_X1   g31744(.A1(new_n34180_), .A2(new_n34179_), .B(pi0966), .ZN(po0769));
  NAND2_X1   g31745(.A1(po0897), .A2(pi1115), .ZN(new_n34182_));
  NAND2_X1   g31746(.A1(new_n34164_), .A2(pi0613), .ZN(new_n34183_));
  AOI21_X1   g31747(.A1(new_n34183_), .A2(new_n34182_), .B(pi0966), .ZN(po0770));
  NOR2_X1    g31748(.A1(po0897), .A2(new_n5405_), .ZN(new_n34185_));
  AOI21_X1   g31749(.A1(pi1102), .A2(po0897), .B(new_n34185_), .ZN(new_n34186_));
  NAND2_X1   g31750(.A1(pi0871), .A2(pi0966), .ZN(new_n34187_));
  OAI21_X1   g31751(.A1(new_n34186_), .A2(pi0966), .B(new_n34187_), .ZN(po0771));
  NOR2_X1    g31752(.A1(new_n34119_), .A2(new_n5473_), .ZN(new_n34189_));
  NAND2_X1   g31753(.A1(pi0779), .A2(pi0797), .ZN(new_n34190_));
  OAI22_X1   g31754(.A1(new_n34189_), .A2(pi0615), .B1(new_n5403_), .B2(new_n34190_), .ZN(po0772));
  NOR2_X1    g31755(.A1(po0897), .A2(new_n13111_), .ZN(new_n34192_));
  AOI21_X1   g31756(.A1(pi1101), .A2(po0897), .B(new_n34192_), .ZN(new_n34193_));
  NAND2_X1   g31757(.A1(pi0872), .A2(pi0966), .ZN(new_n34194_));
  OAI21_X1   g31758(.A1(new_n34193_), .A2(pi0966), .B(new_n34194_), .ZN(po0773));
  NAND2_X1   g31759(.A1(pi0850), .A2(pi0966), .ZN(new_n34196_));
  NOR2_X1    g31760(.A1(po0897), .A2(new_n24970_), .ZN(new_n34197_));
  AOI21_X1   g31761(.A1(pi1105), .A2(po0897), .B(new_n34197_), .ZN(new_n34198_));
  OAI21_X1   g31762(.A1(new_n34198_), .A2(pi0966), .B(new_n34196_), .ZN(po0774));
  NAND2_X1   g31763(.A1(po0897), .A2(pi1117), .ZN(new_n34200_));
  NAND2_X1   g31764(.A1(new_n34164_), .A2(pi0618), .ZN(new_n34201_));
  AOI21_X1   g31765(.A1(new_n34201_), .A2(new_n34200_), .B(pi0966), .ZN(po0775));
  NAND2_X1   g31766(.A1(po0897), .A2(pi1122), .ZN(new_n34203_));
  NAND2_X1   g31767(.A1(new_n34164_), .A2(pi0619), .ZN(new_n34204_));
  AOI21_X1   g31768(.A1(new_n34204_), .A2(new_n34203_), .B(pi0966), .ZN(po0776));
  NAND2_X1   g31769(.A1(po0897), .A2(pi1112), .ZN(new_n34206_));
  NAND2_X1   g31770(.A1(new_n34164_), .A2(pi0620), .ZN(new_n34207_));
  AOI21_X1   g31771(.A1(new_n34207_), .A2(new_n34206_), .B(pi0966), .ZN(po0777));
  NAND2_X1   g31772(.A1(po0897), .A2(pi1108), .ZN(new_n34209_));
  NAND2_X1   g31773(.A1(new_n34164_), .A2(pi0621), .ZN(new_n34210_));
  AOI21_X1   g31774(.A1(new_n34210_), .A2(new_n34209_), .B(pi0966), .ZN(po0778));
  NAND2_X1   g31775(.A1(po0897), .A2(pi1109), .ZN(new_n34212_));
  NAND2_X1   g31776(.A1(new_n34164_), .A2(pi0622), .ZN(new_n34213_));
  AOI21_X1   g31777(.A1(new_n34213_), .A2(new_n34212_), .B(pi0966), .ZN(po0779));
  NAND2_X1   g31778(.A1(po0897), .A2(pi1106), .ZN(new_n34215_));
  NAND2_X1   g31779(.A1(new_n34164_), .A2(pi0623), .ZN(new_n34216_));
  AOI21_X1   g31780(.A1(new_n34216_), .A2(new_n34215_), .B(pi0966), .ZN(po0780));
  AND2_X2    g31781(.A1(new_n5408_), .A2(pi0831), .Z(new_n34218_));
  INV_X1     g31782(.I(pi0780), .ZN(new_n34219_));
  NAND2_X1   g31783(.A1(new_n34218_), .A2(new_n34219_), .ZN(new_n34220_));
  OAI21_X1   g31784(.A1(new_n34153_), .A2(new_n5692_), .B(pi0624), .ZN(new_n34221_));
  OAI21_X1   g31785(.A1(new_n34218_), .A2(new_n34221_), .B(new_n34220_), .ZN(po0781));
  INV_X1     g31786(.I(pi1054), .ZN(new_n34223_));
  AND3_X2    g31787(.A1(new_n34223_), .A2(pi1066), .A3(pi1088), .Z(new_n34224_));
  NOR2_X1    g31788(.A1(new_n12738_), .A2(pi0973), .ZN(new_n34225_));
  NAND2_X1   g31789(.A1(new_n34224_), .A2(new_n34225_), .ZN(new_n34226_));
  NOR2_X1    g31790(.A1(new_n34226_), .A2(pi0953), .ZN(po0954));
  NAND2_X1   g31791(.A1(po0954), .A2(pi1116), .ZN(new_n34228_));
  INV_X1     g31792(.I(po0954), .ZN(new_n34229_));
  NAND2_X1   g31793(.A1(new_n34229_), .A2(pi0625), .ZN(new_n34230_));
  AOI21_X1   g31794(.A1(new_n34230_), .A2(new_n34228_), .B(pi0962), .ZN(po0782));
  NAND2_X1   g31795(.A1(po0897), .A2(pi1121), .ZN(new_n34232_));
  NAND2_X1   g31796(.A1(new_n34164_), .A2(pi0626), .ZN(new_n34233_));
  AOI21_X1   g31797(.A1(new_n34233_), .A2(new_n34232_), .B(pi0966), .ZN(po0783));
  NAND2_X1   g31798(.A1(po0954), .A2(pi1117), .ZN(new_n34235_));
  NAND2_X1   g31799(.A1(new_n34229_), .A2(pi0627), .ZN(new_n34236_));
  AOI21_X1   g31800(.A1(new_n34236_), .A2(new_n34235_), .B(pi0962), .ZN(po0784));
  NAND2_X1   g31801(.A1(po0954), .A2(pi1119), .ZN(new_n34238_));
  NAND2_X1   g31802(.A1(new_n34229_), .A2(pi0628), .ZN(new_n34239_));
  AOI21_X1   g31803(.A1(new_n34239_), .A2(new_n34238_), .B(pi0962), .ZN(po0785));
  NAND2_X1   g31804(.A1(po0897), .A2(pi1119), .ZN(new_n34241_));
  NAND2_X1   g31805(.A1(new_n34164_), .A2(pi0629), .ZN(new_n34242_));
  AOI21_X1   g31806(.A1(new_n34242_), .A2(new_n34241_), .B(pi0966), .ZN(po0786));
  NAND2_X1   g31807(.A1(po0897), .A2(pi1120), .ZN(new_n34244_));
  NAND2_X1   g31808(.A1(new_n34164_), .A2(pi0630), .ZN(new_n34245_));
  AOI21_X1   g31809(.A1(new_n34245_), .A2(new_n34244_), .B(pi0966), .ZN(po0787));
  OR2_X2     g31810(.A1(po0954), .A2(pi0631), .Z(new_n34247_));
  NAND2_X1   g31811(.A1(po0954), .A2(pi1113), .ZN(new_n34248_));
  AOI21_X1   g31812(.A1(new_n34247_), .A2(new_n34248_), .B(pi0962), .ZN(po0788));
  OR2_X2     g31813(.A1(po0954), .A2(pi0632), .Z(new_n34250_));
  NAND2_X1   g31814(.A1(po0954), .A2(pi1115), .ZN(new_n34251_));
  AOI21_X1   g31815(.A1(new_n34250_), .A2(new_n34251_), .B(pi0962), .ZN(po0789));
  NAND2_X1   g31816(.A1(po0897), .A2(pi1110), .ZN(new_n34253_));
  NAND2_X1   g31817(.A1(new_n34164_), .A2(pi0633), .ZN(new_n34254_));
  AOI21_X1   g31818(.A1(new_n34254_), .A2(new_n34253_), .B(pi0966), .ZN(po0790));
  NAND2_X1   g31819(.A1(po0954), .A2(pi1110), .ZN(new_n34256_));
  NAND2_X1   g31820(.A1(new_n34229_), .A2(pi0634), .ZN(new_n34257_));
  AOI21_X1   g31821(.A1(new_n34257_), .A2(new_n34256_), .B(pi0962), .ZN(po0791));
  OR2_X2     g31822(.A1(po0954), .A2(pi0635), .Z(new_n34259_));
  NAND2_X1   g31823(.A1(po0954), .A2(pi1112), .ZN(new_n34260_));
  AOI21_X1   g31824(.A1(new_n34259_), .A2(new_n34260_), .B(pi0962), .ZN(po0792));
  NAND2_X1   g31825(.A1(po0897), .A2(pi1127), .ZN(new_n34262_));
  NAND2_X1   g31826(.A1(new_n34164_), .A2(pi0636), .ZN(new_n34263_));
  AOI21_X1   g31827(.A1(new_n34263_), .A2(new_n34262_), .B(pi0966), .ZN(po0793));
  NAND2_X1   g31828(.A1(po0954), .A2(pi1105), .ZN(new_n34265_));
  NAND2_X1   g31829(.A1(new_n34229_), .A2(pi0637), .ZN(new_n34266_));
  AOI21_X1   g31830(.A1(new_n34266_), .A2(new_n34265_), .B(pi0962), .ZN(po0794));
  NAND2_X1   g31831(.A1(po0954), .A2(pi1107), .ZN(new_n34268_));
  NAND2_X1   g31832(.A1(new_n34229_), .A2(pi0638), .ZN(new_n34269_));
  AOI21_X1   g31833(.A1(new_n34269_), .A2(new_n34268_), .B(pi0962), .ZN(po0795));
  NAND2_X1   g31834(.A1(po0954), .A2(pi1109), .ZN(new_n34271_));
  NAND2_X1   g31835(.A1(new_n34229_), .A2(pi0639), .ZN(new_n34272_));
  AOI21_X1   g31836(.A1(new_n34272_), .A2(new_n34271_), .B(pi0962), .ZN(po0796));
  NAND2_X1   g31837(.A1(po0897), .A2(pi1128), .ZN(new_n34274_));
  NAND2_X1   g31838(.A1(new_n34164_), .A2(pi0640), .ZN(new_n34275_));
  AOI21_X1   g31839(.A1(new_n34275_), .A2(new_n34274_), .B(pi0966), .ZN(po0797));
  NAND2_X1   g31840(.A1(po0954), .A2(pi1121), .ZN(new_n34277_));
  NAND2_X1   g31841(.A1(new_n34229_), .A2(pi0641), .ZN(new_n34278_));
  AOI21_X1   g31842(.A1(new_n34278_), .A2(new_n34277_), .B(pi0962), .ZN(po0798));
  NAND2_X1   g31843(.A1(po0897), .A2(pi1103), .ZN(new_n34280_));
  NAND2_X1   g31844(.A1(new_n34164_), .A2(pi0642), .ZN(new_n34281_));
  AOI21_X1   g31845(.A1(new_n34281_), .A2(new_n34280_), .B(pi0966), .ZN(po0799));
  NAND2_X1   g31846(.A1(po0954), .A2(pi1104), .ZN(new_n34283_));
  NAND2_X1   g31847(.A1(new_n34229_), .A2(pi0643), .ZN(new_n34284_));
  AOI21_X1   g31848(.A1(new_n34284_), .A2(new_n34283_), .B(pi0962), .ZN(po0800));
  NAND2_X1   g31849(.A1(po0897), .A2(pi1123), .ZN(new_n34286_));
  NAND2_X1   g31850(.A1(new_n34164_), .A2(pi0644), .ZN(new_n34287_));
  AOI21_X1   g31851(.A1(new_n34287_), .A2(new_n34286_), .B(pi0966), .ZN(po0801));
  NAND2_X1   g31852(.A1(po0897), .A2(pi1125), .ZN(new_n34289_));
  NAND2_X1   g31853(.A1(new_n34164_), .A2(pi0645), .ZN(new_n34290_));
  AOI21_X1   g31854(.A1(new_n34290_), .A2(new_n34289_), .B(pi0966), .ZN(po0802));
  OR2_X2     g31855(.A1(po0954), .A2(pi0646), .Z(new_n34292_));
  NAND2_X1   g31856(.A1(po0954), .A2(pi1114), .ZN(new_n34293_));
  AOI21_X1   g31857(.A1(new_n34292_), .A2(new_n34293_), .B(pi0962), .ZN(po0803));
  NAND2_X1   g31858(.A1(po0954), .A2(pi1120), .ZN(new_n34295_));
  NAND2_X1   g31859(.A1(new_n34229_), .A2(pi0647), .ZN(new_n34296_));
  AOI21_X1   g31860(.A1(new_n34296_), .A2(new_n34295_), .B(pi0962), .ZN(po0804));
  NAND2_X1   g31861(.A1(po0954), .A2(pi1122), .ZN(new_n34298_));
  NAND2_X1   g31862(.A1(new_n34229_), .A2(pi0648), .ZN(new_n34299_));
  AOI21_X1   g31863(.A1(new_n34299_), .A2(new_n34298_), .B(pi0962), .ZN(po0805));
  OR2_X2     g31864(.A1(po0954), .A2(pi0649), .Z(new_n34301_));
  NAND2_X1   g31865(.A1(po0954), .A2(pi1126), .ZN(new_n34302_));
  AOI21_X1   g31866(.A1(new_n34301_), .A2(new_n34302_), .B(pi0962), .ZN(po0806));
  OR2_X2     g31867(.A1(po0954), .A2(pi0650), .Z(new_n34304_));
  NAND2_X1   g31868(.A1(po0954), .A2(pi1127), .ZN(new_n34305_));
  AOI21_X1   g31869(.A1(new_n34304_), .A2(new_n34305_), .B(pi0962), .ZN(po0807));
  NAND2_X1   g31870(.A1(po0897), .A2(pi1130), .ZN(new_n34307_));
  NAND2_X1   g31871(.A1(new_n34164_), .A2(pi0651), .ZN(new_n34308_));
  AOI21_X1   g31872(.A1(new_n34308_), .A2(new_n34307_), .B(pi0966), .ZN(po0808));
  NAND2_X1   g31873(.A1(po0897), .A2(pi1131), .ZN(new_n34310_));
  NAND2_X1   g31874(.A1(new_n34164_), .A2(pi0652), .ZN(new_n34311_));
  AOI21_X1   g31875(.A1(new_n34311_), .A2(new_n34310_), .B(pi0966), .ZN(po0809));
  NAND2_X1   g31876(.A1(po0897), .A2(pi1129), .ZN(new_n34313_));
  NAND2_X1   g31877(.A1(new_n34164_), .A2(pi0653), .ZN(new_n34314_));
  AOI21_X1   g31878(.A1(new_n34314_), .A2(new_n34313_), .B(pi0966), .ZN(po0810));
  OR2_X2     g31879(.A1(po0954), .A2(pi0654), .Z(new_n34316_));
  NAND2_X1   g31880(.A1(po0954), .A2(pi1130), .ZN(new_n34317_));
  AOI21_X1   g31881(.A1(new_n34316_), .A2(new_n34317_), .B(pi0962), .ZN(po0811));
  OR2_X2     g31882(.A1(po0954), .A2(pi0655), .Z(new_n34319_));
  NAND2_X1   g31883(.A1(po0954), .A2(pi1124), .ZN(new_n34320_));
  AOI21_X1   g31884(.A1(new_n34319_), .A2(new_n34320_), .B(pi0962), .ZN(po0812));
  NAND2_X1   g31885(.A1(po0897), .A2(pi1126), .ZN(new_n34322_));
  NAND2_X1   g31886(.A1(new_n34164_), .A2(pi0656), .ZN(new_n34323_));
  AOI21_X1   g31887(.A1(new_n34323_), .A2(new_n34322_), .B(pi0966), .ZN(po0813));
  OR2_X2     g31888(.A1(po0954), .A2(pi0657), .Z(new_n34325_));
  NAND2_X1   g31889(.A1(po0954), .A2(pi1131), .ZN(new_n34326_));
  AOI21_X1   g31890(.A1(new_n34325_), .A2(new_n34326_), .B(pi0962), .ZN(po0814));
  NAND2_X1   g31891(.A1(po0897), .A2(pi1124), .ZN(new_n34328_));
  NAND2_X1   g31892(.A1(new_n34164_), .A2(pi0658), .ZN(new_n34329_));
  AOI21_X1   g31893(.A1(new_n34329_), .A2(new_n34328_), .B(pi0966), .ZN(po0815));
  NAND3_X1   g31894(.A1(new_n32317_), .A2(pi0266), .A3(pi0992), .ZN(new_n34331_));
  NOR3_X1    g31895(.A1(new_n34331_), .A2(pi0269), .A3(pi0281), .ZN(new_n34332_));
  NOR3_X1    g31896(.A1(pi0270), .A2(pi0277), .A3(pi0282), .ZN(new_n34333_));
  NAND3_X1   g31897(.A1(new_n34332_), .A2(new_n31562_), .A3(new_n34333_), .ZN(new_n34334_));
  NOR2_X1    g31898(.A1(new_n34334_), .A2(pi0265), .ZN(new_n34335_));
  XOR2_X1    g31899(.A1(new_n34335_), .A2(new_n32106_), .Z(po0816));
  NAND2_X1   g31900(.A1(po0954), .A2(pi1118), .ZN(new_n34337_));
  NAND2_X1   g31901(.A1(new_n34229_), .A2(pi0660), .ZN(new_n34338_));
  AOI21_X1   g31902(.A1(new_n34338_), .A2(new_n34337_), .B(pi0962), .ZN(po0817));
  NAND2_X1   g31903(.A1(po0954), .A2(pi1101), .ZN(new_n34340_));
  NAND2_X1   g31904(.A1(new_n34229_), .A2(pi0661), .ZN(new_n34341_));
  AOI21_X1   g31905(.A1(new_n34341_), .A2(new_n34340_), .B(pi0962), .ZN(po0818));
  NAND2_X1   g31906(.A1(po0954), .A2(pi1102), .ZN(new_n34343_));
  NAND2_X1   g31907(.A1(new_n34229_), .A2(pi0662), .ZN(new_n34344_));
  AOI21_X1   g31908(.A1(new_n34344_), .A2(new_n34343_), .B(pi0962), .ZN(po0819));
  OAI22_X1   g31909(.A1(new_n4888_), .A2(pi0700), .B1(pi0855), .B2(pi1136), .ZN(new_n34346_));
  NOR2_X1    g31910(.A1(pi1137), .A2(pi1138), .ZN(new_n34347_));
  INV_X1     g31911(.I(new_n34347_), .ZN(new_n34348_));
  NOR2_X1    g31912(.A1(new_n34348_), .A2(new_n5045_), .ZN(new_n34349_));
  NOR2_X1    g31913(.A1(new_n4888_), .A2(pi1136), .ZN(new_n34350_));
  INV_X1     g31914(.I(new_n34350_), .ZN(new_n34351_));
  NAND2_X1   g31915(.A1(new_n34349_), .A2(new_n34351_), .ZN(new_n34352_));
  AOI21_X1   g31916(.A1(new_n34347_), .A2(pi1135), .B(new_n4724_), .ZN(new_n34353_));
  INV_X1     g31917(.I(new_n34353_), .ZN(new_n34354_));
  NOR2_X1    g31918(.A1(new_n34354_), .A2(pi0766), .ZN(new_n34355_));
  NOR3_X1    g31919(.A1(new_n34355_), .A2(new_n34352_), .A3(new_n34346_), .ZN(new_n34356_));
  NOR2_X1    g31920(.A1(new_n34348_), .A2(pi1134), .ZN(new_n34357_));
  INV_X1     g31921(.I(new_n34357_), .ZN(new_n34358_));
  NOR2_X1    g31922(.A1(new_n24493_), .A2(new_n4724_), .ZN(new_n34359_));
  INV_X1     g31923(.I(pi0784), .ZN(new_n34360_));
  NOR2_X1    g31924(.A1(new_n34360_), .A2(pi1136), .ZN(new_n34361_));
  OAI21_X1   g31925(.A1(new_n34359_), .A2(new_n34361_), .B(pi1135), .ZN(new_n34362_));
  NOR2_X1    g31926(.A1(new_n24611_), .A2(new_n4724_), .ZN(new_n34363_));
  NOR2_X1    g31927(.A1(new_n32938_), .A2(pi1136), .ZN(new_n34364_));
  OAI21_X1   g31928(.A1(new_n34363_), .A2(new_n34364_), .B(new_n4888_), .ZN(new_n34365_));
  AOI21_X1   g31929(.A1(new_n34362_), .A2(new_n34365_), .B(new_n34358_), .ZN(new_n34366_));
  NOR3_X1    g31930(.A1(new_n34356_), .A2(new_n34366_), .A3(new_n7253_), .ZN(new_n34367_));
  NOR2_X1    g31931(.A1(pi0223), .A2(pi0224), .ZN(new_n34368_));
  INV_X1     g31932(.I(new_n34368_), .ZN(new_n34369_));
  NOR2_X1    g31933(.A1(new_n6254_), .A2(pi0592), .ZN(new_n34370_));
  NAND2_X1   g31934(.A1(new_n34370_), .A2(pi0464), .ZN(new_n34371_));
  AOI21_X1   g31935(.A1(new_n34371_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34372_));
  NOR2_X1    g31936(.A1(pi0591), .A2(pi0592), .ZN(new_n34373_));
  INV_X1     g31937(.I(new_n34373_), .ZN(new_n34374_));
  NOR2_X1    g31938(.A1(new_n34374_), .A2(new_n6352_), .ZN(new_n34375_));
  AOI21_X1   g31939(.A1(new_n34375_), .A2(pi0323), .B(pi0588), .ZN(new_n34376_));
  NOR2_X1    g31940(.A1(new_n6268_), .A2(pi0591), .ZN(new_n34377_));
  NOR2_X1    g31941(.A1(new_n6440_), .A2(pi0592), .ZN(new_n34378_));
  AOI22_X1   g31942(.A1(pi0334), .A2(new_n34378_), .B1(new_n34377_), .B2(pi0365), .ZN(new_n34379_));
  OAI21_X1   g31943(.A1(pi0590), .A2(new_n34379_), .B(new_n34376_), .ZN(new_n34380_));
  NOR2_X1    g31944(.A1(new_n31349_), .A2(pi0199), .ZN(new_n34381_));
  AOI21_X1   g31945(.A1(pi0199), .A2(pi1065), .B(new_n34381_), .ZN(new_n34382_));
  OAI21_X1   g31946(.A1(new_n34382_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34383_));
  AOI21_X1   g31947(.A1(new_n34380_), .A2(new_n34372_), .B(new_n34383_), .ZN(new_n34384_));
  NOR2_X1    g31948(.A1(new_n34384_), .A2(new_n34367_), .ZN(po0820));
  NAND2_X1   g31949(.A1(pi0199), .A2(pi1084), .ZN(new_n34386_));
  NAND2_X1   g31950(.A1(new_n8525_), .A2(pi0292), .ZN(new_n34387_));
  AOI21_X1   g31951(.A1(new_n34387_), .A2(new_n34386_), .B(new_n34368_), .ZN(new_n34388_));
  INV_X1     g31952(.I(new_n34370_), .ZN(new_n34389_));
  OAI21_X1   g31953(.A1(new_n34389_), .A2(new_n10059_), .B(pi0588), .ZN(new_n34390_));
  NAND2_X1   g31954(.A1(new_n34390_), .A2(new_n34368_), .ZN(new_n34391_));
  NOR2_X1    g31955(.A1(new_n6268_), .A2(pi0590), .ZN(new_n34392_));
  NOR2_X1    g31956(.A1(new_n34392_), .A2(pi0588), .ZN(new_n34393_));
  INV_X1     g31957(.I(new_n34393_), .ZN(new_n34394_));
  NOR3_X1    g31958(.A1(new_n9829_), .A2(new_n6440_), .A3(pi0590), .ZN(new_n34395_));
  NOR2_X1    g31959(.A1(new_n32750_), .A2(pi0591), .ZN(new_n34396_));
  OAI22_X1   g31960(.A1(new_n34394_), .A2(new_n34395_), .B1(new_n6268_), .B2(new_n34396_), .ZN(new_n34397_));
  NAND2_X1   g31961(.A1(new_n34375_), .A2(pi0355), .ZN(new_n34398_));
  AOI21_X1   g31962(.A1(new_n34397_), .A2(new_n34398_), .B(new_n34391_), .ZN(new_n34399_));
  OAI21_X1   g31963(.A1(new_n34399_), .A2(new_n34388_), .B(new_n7253_), .ZN(new_n34400_));
  NAND2_X1   g31964(.A1(new_n12764_), .A2(pi1135), .ZN(new_n34401_));
  INV_X1     g31965(.I(pi0811), .ZN(new_n34402_));
  NAND2_X1   g31966(.A1(new_n34402_), .A2(new_n4888_), .ZN(new_n34403_));
  AOI21_X1   g31967(.A1(new_n34403_), .A2(new_n34401_), .B(pi1136), .ZN(new_n34404_));
  NAND2_X1   g31968(.A1(new_n5405_), .A2(new_n4888_), .ZN(new_n34405_));
  NAND2_X1   g31969(.A1(new_n5400_), .A2(pi1135), .ZN(new_n34406_));
  AOI21_X1   g31970(.A1(new_n34405_), .A2(new_n34406_), .B(new_n4724_), .ZN(new_n34407_));
  OAI21_X1   g31971(.A1(new_n34404_), .A2(new_n34407_), .B(new_n5045_), .ZN(new_n34408_));
  NOR2_X1    g31972(.A1(new_n16845_), .A2(pi1135), .ZN(new_n34409_));
  AOI21_X1   g31973(.A1(pi0727), .A2(pi1135), .B(new_n34409_), .ZN(new_n34410_));
  NOR2_X1    g31974(.A1(pi1135), .A2(pi1136), .ZN(new_n34411_));
  AOI21_X1   g31975(.A1(new_n34411_), .A2(pi0872), .B(new_n5045_), .ZN(new_n34412_));
  OAI21_X1   g31976(.A1(new_n34410_), .A2(new_n4724_), .B(new_n34412_), .ZN(new_n34413_));
  NOR2_X1    g31977(.A1(new_n34348_), .A2(new_n7253_), .ZN(new_n34414_));
  NAND3_X1   g31978(.A1(new_n34408_), .A2(new_n34413_), .A3(new_n34414_), .ZN(new_n34415_));
  NAND2_X1   g31979(.A1(new_n34400_), .A2(new_n34415_), .ZN(po0821));
  NAND2_X1   g31980(.A1(po0954), .A2(pi1108), .ZN(new_n34417_));
  NAND2_X1   g31981(.A1(new_n34229_), .A2(pi0665), .ZN(new_n34418_));
  AOI21_X1   g31982(.A1(new_n34418_), .A2(new_n34417_), .B(pi0962), .ZN(po0822));
  OAI22_X1   g31983(.A1(new_n4888_), .A2(pi0691), .B1(pi0873), .B2(pi1136), .ZN(new_n34420_));
  NOR2_X1    g31984(.A1(new_n34354_), .A2(pi0764), .ZN(new_n34421_));
  NOR3_X1    g31985(.A1(new_n34421_), .A2(new_n34352_), .A3(new_n34420_), .ZN(new_n34422_));
  NOR2_X1    g31986(.A1(new_n25921_), .A2(new_n4888_), .ZN(new_n34423_));
  NOR2_X1    g31987(.A1(new_n25938_), .A2(pi1135), .ZN(new_n34424_));
  OAI21_X1   g31988(.A1(new_n34423_), .A2(new_n34424_), .B(pi1136), .ZN(new_n34425_));
  NOR2_X1    g31989(.A1(pi0799), .A2(pi1135), .ZN(new_n34426_));
  NOR2_X1    g31990(.A1(new_n13000_), .A2(new_n4888_), .ZN(new_n34427_));
  OAI21_X1   g31991(.A1(new_n34427_), .A2(new_n34426_), .B(new_n4724_), .ZN(new_n34428_));
  AOI21_X1   g31992(.A1(new_n34425_), .A2(new_n34428_), .B(new_n34358_), .ZN(new_n34429_));
  NOR3_X1    g31993(.A1(new_n34422_), .A2(new_n34429_), .A3(new_n7253_), .ZN(new_n34430_));
  NAND2_X1   g31994(.A1(new_n34370_), .A2(pi0443), .ZN(new_n34431_));
  AOI21_X1   g31995(.A1(new_n34431_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34432_));
  INV_X1     g31996(.I(new_n34375_), .ZN(new_n34433_));
  NOR3_X1    g31997(.A1(new_n6386_), .A2(new_n6440_), .A3(pi0590), .ZN(new_n34434_));
  NOR2_X1    g31998(.A1(new_n34394_), .A2(new_n34434_), .ZN(new_n34435_));
  AOI21_X1   g31999(.A1(pi0337), .A2(new_n6440_), .B(new_n6268_), .ZN(new_n34436_));
  OAI22_X1   g32000(.A1(new_n34435_), .A2(new_n34436_), .B1(new_n6518_), .B2(new_n34433_), .ZN(new_n34437_));
  NOR2_X1    g32001(.A1(new_n8525_), .A2(new_n32496_), .ZN(new_n34438_));
  AOI21_X1   g32002(.A1(new_n8525_), .A2(pi0297), .B(new_n34438_), .ZN(new_n34439_));
  OAI21_X1   g32003(.A1(new_n34439_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34440_));
  AOI21_X1   g32004(.A1(new_n34437_), .A2(new_n34432_), .B(new_n34440_), .ZN(new_n34441_));
  NOR2_X1    g32005(.A1(new_n34441_), .A2(new_n34430_), .ZN(po0823));
  NAND2_X1   g32006(.A1(pi0199), .A2(pi1072), .ZN(new_n34443_));
  NAND2_X1   g32007(.A1(new_n8525_), .A2(pi0294), .ZN(new_n34444_));
  AOI21_X1   g32008(.A1(new_n34444_), .A2(new_n34443_), .B(new_n34368_), .ZN(new_n34445_));
  OAI21_X1   g32009(.A1(new_n34389_), .A2(new_n6891_), .B(pi0588), .ZN(new_n34446_));
  NAND2_X1   g32010(.A1(new_n34446_), .A2(new_n34368_), .ZN(new_n34447_));
  NOR3_X1    g32011(.A1(new_n6389_), .A2(new_n6440_), .A3(pi0590), .ZN(new_n34448_));
  NOR2_X1    g32012(.A1(new_n32649_), .A2(pi0591), .ZN(new_n34449_));
  OAI22_X1   g32013(.A1(new_n34394_), .A2(new_n34448_), .B1(new_n6268_), .B2(new_n34449_), .ZN(new_n34450_));
  NAND2_X1   g32014(.A1(new_n34375_), .A2(pi0458), .ZN(new_n34451_));
  AOI21_X1   g32015(.A1(new_n34450_), .A2(new_n34451_), .B(new_n34447_), .ZN(new_n34452_));
  OAI21_X1   g32016(.A1(new_n34452_), .A2(new_n34445_), .B(new_n7253_), .ZN(new_n34453_));
  NAND2_X1   g32017(.A1(new_n5406_), .A2(pi1136), .ZN(new_n34454_));
  NAND2_X1   g32018(.A1(new_n4724_), .A2(pi0809), .ZN(new_n34455_));
  AOI21_X1   g32019(.A1(new_n34454_), .A2(new_n34455_), .B(pi1135), .ZN(new_n34456_));
  NAND2_X1   g32020(.A1(new_n5399_), .A2(pi1136), .ZN(new_n34457_));
  NAND2_X1   g32021(.A1(new_n12937_), .A2(new_n4724_), .ZN(new_n34458_));
  AOI21_X1   g32022(.A1(new_n34458_), .A2(new_n34457_), .B(new_n4888_), .ZN(new_n34459_));
  OAI21_X1   g32023(.A1(new_n34459_), .A2(new_n34456_), .B(new_n5045_), .ZN(new_n34460_));
  NOR2_X1    g32024(.A1(new_n16945_), .A2(pi1135), .ZN(new_n34461_));
  AOI21_X1   g32025(.A1(pi0699), .A2(pi1135), .B(new_n34461_), .ZN(new_n34462_));
  AOI21_X1   g32026(.A1(new_n34411_), .A2(pi0871), .B(new_n5045_), .ZN(new_n34463_));
  OAI21_X1   g32027(.A1(new_n34462_), .A2(new_n4724_), .B(new_n34463_), .ZN(new_n34464_));
  NAND3_X1   g32028(.A1(new_n34460_), .A2(new_n34464_), .A3(new_n34414_), .ZN(new_n34465_));
  NAND2_X1   g32029(.A1(new_n34453_), .A2(new_n34465_), .ZN(po0824));
  OAI22_X1   g32030(.A1(new_n4888_), .A2(pi0696), .B1(pi0837), .B2(pi1136), .ZN(new_n34467_));
  NOR2_X1    g32031(.A1(new_n34354_), .A2(pi0759), .ZN(new_n34468_));
  NOR3_X1    g32032(.A1(new_n34468_), .A2(new_n34352_), .A3(new_n34467_), .ZN(new_n34469_));
  NOR2_X1    g32033(.A1(new_n12821_), .A2(new_n4888_), .ZN(new_n34470_));
  NOR2_X1    g32034(.A1(new_n12751_), .A2(pi1135), .ZN(new_n34471_));
  OAI21_X1   g32035(.A1(new_n34470_), .A2(new_n34471_), .B(pi1136), .ZN(new_n34472_));
  NOR2_X1    g32036(.A1(new_n12758_), .A2(new_n4888_), .ZN(new_n34473_));
  INV_X1     g32037(.I(pi0981), .ZN(new_n34474_));
  NOR2_X1    g32038(.A1(new_n34474_), .A2(pi1135), .ZN(new_n34475_));
  OAI21_X1   g32039(.A1(new_n34473_), .A2(new_n34475_), .B(new_n4724_), .ZN(new_n34476_));
  AOI21_X1   g32040(.A1(new_n34472_), .A2(new_n34476_), .B(new_n34358_), .ZN(new_n34477_));
  NOR3_X1    g32041(.A1(new_n34469_), .A2(new_n34477_), .A3(new_n7253_), .ZN(new_n34478_));
  NAND2_X1   g32042(.A1(new_n34370_), .A2(pi0414), .ZN(new_n34479_));
  AOI21_X1   g32043(.A1(new_n34479_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34480_));
  NOR3_X1    g32044(.A1(new_n32772_), .A2(new_n6440_), .A3(pi0590), .ZN(new_n34481_));
  NOR2_X1    g32045(.A1(new_n34394_), .A2(new_n34481_), .ZN(new_n34482_));
  AOI21_X1   g32046(.A1(pi0363), .A2(new_n6440_), .B(new_n6268_), .ZN(new_n34483_));
  OAI22_X1   g32047(.A1(new_n34482_), .A2(new_n34483_), .B1(new_n6469_), .B2(new_n34433_), .ZN(new_n34484_));
  NOR2_X1    g32048(.A1(new_n8525_), .A2(new_n32478_), .ZN(new_n34485_));
  AOI21_X1   g32049(.A1(new_n8525_), .A2(pi0291), .B(new_n34485_), .ZN(new_n34486_));
  OAI21_X1   g32050(.A1(new_n34486_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34487_));
  AOI21_X1   g32051(.A1(new_n34484_), .A2(new_n34480_), .B(new_n34487_), .ZN(new_n34488_));
  NOR2_X1    g32052(.A1(new_n34488_), .A2(new_n34478_), .ZN(po0825));
  OR2_X2     g32053(.A1(po0954), .A2(pi0669), .Z(new_n34490_));
  NAND2_X1   g32054(.A1(po0954), .A2(pi1125), .ZN(new_n34491_));
  AOI21_X1   g32055(.A1(new_n34490_), .A2(new_n34491_), .B(pi0962), .ZN(po0826));
  OAI22_X1   g32056(.A1(new_n16263_), .A2(new_n4888_), .B1(pi0852), .B2(pi1136), .ZN(new_n34493_));
  NOR2_X1    g32057(.A1(new_n34354_), .A2(new_n16245_), .ZN(new_n34494_));
  NOR3_X1    g32058(.A1(new_n34494_), .A2(new_n34352_), .A3(new_n34493_), .ZN(new_n34495_));
  NOR2_X1    g32059(.A1(new_n26373_), .A2(pi1135), .ZN(new_n34496_));
  AOI21_X1   g32060(.A1(new_n26376_), .A2(pi1135), .B(new_n34496_), .ZN(new_n34497_));
  NAND2_X1   g32061(.A1(new_n34347_), .A2(pi1136), .ZN(new_n34498_));
  NOR3_X1    g32062(.A1(new_n34497_), .A2(pi1134), .A3(new_n34498_), .ZN(new_n34499_));
  NOR3_X1    g32063(.A1(new_n34495_), .A2(new_n7253_), .A3(new_n34499_), .ZN(new_n34500_));
  NAND2_X1   g32064(.A1(new_n34370_), .A2(pi0415), .ZN(new_n34501_));
  AOI21_X1   g32065(.A1(new_n34501_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34502_));
  AOI21_X1   g32066(.A1(new_n34375_), .A2(pi0343), .B(pi0588), .ZN(new_n34503_));
  AOI22_X1   g32067(.A1(pi0364), .A2(new_n34377_), .B1(new_n34378_), .B2(pi0391), .ZN(new_n34504_));
  OAI21_X1   g32068(.A1(pi0590), .A2(new_n34504_), .B(new_n34503_), .ZN(new_n34505_));
  NOR2_X1    g32069(.A1(new_n31355_), .A2(pi0199), .ZN(new_n34506_));
  AOI21_X1   g32070(.A1(pi0199), .A2(pi1062), .B(new_n34506_), .ZN(new_n34507_));
  OAI21_X1   g32071(.A1(new_n34507_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34508_));
  AOI21_X1   g32072(.A1(new_n34505_), .A2(new_n34502_), .B(new_n34508_), .ZN(new_n34509_));
  NOR2_X1    g32073(.A1(new_n34509_), .A2(new_n34500_), .ZN(po0827));
  OAI22_X1   g32074(.A1(new_n16499_), .A2(new_n4888_), .B1(pi0865), .B2(pi1136), .ZN(new_n34511_));
  NOR2_X1    g32075(.A1(new_n34354_), .A2(new_n16500_), .ZN(new_n34512_));
  NOR3_X1    g32076(.A1(new_n34512_), .A2(new_n34352_), .A3(new_n34511_), .ZN(new_n34513_));
  NOR2_X1    g32077(.A1(new_n4888_), .A2(pi0646), .ZN(new_n34514_));
  AOI21_X1   g32078(.A1(pi0611), .A2(new_n4888_), .B(new_n34514_), .ZN(new_n34515_));
  NOR3_X1    g32079(.A1(new_n34515_), .A2(pi1134), .A3(new_n34498_), .ZN(new_n34516_));
  NOR3_X1    g32080(.A1(new_n34513_), .A2(new_n7253_), .A3(new_n34516_), .ZN(new_n34517_));
  NAND2_X1   g32081(.A1(new_n34370_), .A2(pi0453), .ZN(new_n34518_));
  AOI21_X1   g32082(.A1(new_n34518_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34519_));
  AOI21_X1   g32083(.A1(new_n34375_), .A2(pi0327), .B(pi0588), .ZN(new_n34520_));
  AOI22_X1   g32084(.A1(pi0333), .A2(new_n34378_), .B1(new_n34377_), .B2(pi0447), .ZN(new_n34521_));
  OAI21_X1   g32085(.A1(pi0590), .A2(new_n34521_), .B(new_n34520_), .ZN(new_n34522_));
  NOR2_X1    g32086(.A1(new_n31373_), .A2(pi0199), .ZN(new_n34523_));
  AOI21_X1   g32087(.A1(pi0199), .A2(pi1040), .B(new_n34523_), .ZN(new_n34524_));
  OAI21_X1   g32088(.A1(new_n34524_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34525_));
  AOI21_X1   g32089(.A1(new_n34522_), .A2(new_n34519_), .B(new_n34525_), .ZN(new_n34526_));
  NOR2_X1    g32090(.A1(new_n34526_), .A2(new_n34517_), .ZN(po0828));
  OAI22_X1   g32091(.A1(new_n4888_), .A2(pi0736), .B1(pi0850), .B2(pi1136), .ZN(new_n34528_));
  NOR2_X1    g32092(.A1(new_n34354_), .A2(pi0758), .ZN(new_n34529_));
  NOR3_X1    g32093(.A1(new_n34529_), .A2(new_n34352_), .A3(new_n34528_), .ZN(new_n34530_));
  NOR2_X1    g32094(.A1(new_n26413_), .A2(new_n4888_), .ZN(new_n34531_));
  NOR2_X1    g32095(.A1(new_n13111_), .A2(pi1135), .ZN(new_n34532_));
  OAI21_X1   g32096(.A1(new_n34531_), .A2(new_n34532_), .B(pi1136), .ZN(new_n34533_));
  NOR2_X1    g32097(.A1(new_n12779_), .A2(new_n4888_), .ZN(new_n34534_));
  INV_X1     g32098(.I(pi0808), .ZN(new_n34535_));
  NOR2_X1    g32099(.A1(new_n34535_), .A2(pi1135), .ZN(new_n34536_));
  OAI21_X1   g32100(.A1(new_n34534_), .A2(new_n34536_), .B(new_n4724_), .ZN(new_n34537_));
  AOI21_X1   g32101(.A1(new_n34533_), .A2(new_n34537_), .B(new_n34358_), .ZN(new_n34538_));
  NOR3_X1    g32102(.A1(new_n34530_), .A2(new_n34538_), .A3(new_n7253_), .ZN(new_n34539_));
  NAND2_X1   g32103(.A1(new_n34370_), .A2(pi0422), .ZN(new_n34540_));
  AOI21_X1   g32104(.A1(new_n34540_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34541_));
  NOR3_X1    g32105(.A1(new_n9832_), .A2(new_n6440_), .A3(pi0590), .ZN(new_n34542_));
  NOR2_X1    g32106(.A1(new_n34394_), .A2(new_n34542_), .ZN(new_n34543_));
  AOI21_X1   g32107(.A1(pi0372), .A2(new_n6440_), .B(new_n6268_), .ZN(new_n34544_));
  OAI22_X1   g32108(.A1(new_n34543_), .A2(new_n34544_), .B1(new_n6473_), .B2(new_n34433_), .ZN(new_n34545_));
  NOR2_X1    g32109(.A1(new_n8525_), .A2(new_n32475_), .ZN(new_n34546_));
  AOI21_X1   g32110(.A1(new_n8525_), .A2(pi0290), .B(new_n34546_), .ZN(new_n34547_));
  OAI21_X1   g32111(.A1(new_n34547_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34548_));
  AOI21_X1   g32112(.A1(new_n34545_), .A2(new_n34541_), .B(new_n34548_), .ZN(new_n34549_));
  NOR2_X1    g32113(.A1(new_n34549_), .A2(new_n34539_), .ZN(po0829));
  OAI22_X1   g32114(.A1(new_n4888_), .A2(pi0706), .B1(pi0866), .B2(pi1136), .ZN(new_n34551_));
  NOR2_X1    g32115(.A1(new_n34354_), .A2(pi0749), .ZN(new_n34552_));
  NOR3_X1    g32116(.A1(new_n34552_), .A2(new_n34352_), .A3(new_n34551_), .ZN(new_n34553_));
  NOR2_X1    g32117(.A1(new_n24943_), .A2(new_n4888_), .ZN(new_n34554_));
  NOR2_X1    g32118(.A1(new_n24970_), .A2(pi1135), .ZN(new_n34555_));
  OAI21_X1   g32119(.A1(new_n34554_), .A2(new_n34555_), .B(pi1136), .ZN(new_n34556_));
  NOR2_X1    g32120(.A1(pi0814), .A2(pi1135), .ZN(new_n34557_));
  NOR2_X1    g32121(.A1(new_n12808_), .A2(new_n4888_), .ZN(new_n34558_));
  OAI21_X1   g32122(.A1(new_n34558_), .A2(new_n34557_), .B(new_n4724_), .ZN(new_n34559_));
  AOI21_X1   g32123(.A1(new_n34556_), .A2(new_n34559_), .B(new_n34358_), .ZN(new_n34560_));
  NOR3_X1    g32124(.A1(new_n34553_), .A2(new_n34560_), .A3(new_n7253_), .ZN(new_n34561_));
  NAND2_X1   g32125(.A1(new_n34370_), .A2(pi0435), .ZN(new_n34562_));
  AOI21_X1   g32126(.A1(new_n34562_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34563_));
  NOR3_X1    g32127(.A1(new_n6382_), .A2(new_n6440_), .A3(pi0590), .ZN(new_n34564_));
  NOR2_X1    g32128(.A1(new_n34394_), .A2(new_n34564_), .ZN(new_n34565_));
  AOI21_X1   g32129(.A1(pi0387), .A2(new_n6440_), .B(new_n6268_), .ZN(new_n34566_));
  OAI22_X1   g32130(.A1(new_n34565_), .A2(new_n34566_), .B1(new_n6487_), .B2(new_n34433_), .ZN(new_n34567_));
  NOR2_X1    g32131(.A1(new_n8525_), .A2(new_n32490_), .ZN(new_n34568_));
  AOI21_X1   g32132(.A1(new_n8525_), .A2(pi0295), .B(new_n34568_), .ZN(new_n34569_));
  OAI21_X1   g32133(.A1(new_n34569_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34570_));
  AOI21_X1   g32134(.A1(new_n34567_), .A2(new_n34563_), .B(new_n34570_), .ZN(new_n34571_));
  NOR2_X1    g32135(.A1(new_n34571_), .A2(new_n34561_), .ZN(po0830));
  NAND2_X1   g32136(.A1(pi0199), .A2(pi1070), .ZN(new_n34573_));
  NAND2_X1   g32137(.A1(new_n8525_), .A2(pi0256), .ZN(new_n34574_));
  AOI21_X1   g32138(.A1(new_n34574_), .A2(new_n34573_), .B(new_n34368_), .ZN(new_n34575_));
  OAI21_X1   g32139(.A1(new_n34389_), .A2(new_n6286_), .B(pi0588), .ZN(new_n34576_));
  NAND2_X1   g32140(.A1(new_n34576_), .A2(new_n34368_), .ZN(new_n34577_));
  AOI21_X1   g32141(.A1(new_n34375_), .A2(pi0362), .B(pi0588), .ZN(new_n34578_));
  INV_X1     g32142(.I(new_n34377_), .ZN(new_n34579_));
  INV_X1     g32143(.I(new_n34378_), .ZN(new_n34580_));
  OAI22_X1   g32144(.A1(new_n32643_), .A2(new_n34579_), .B1(new_n34580_), .B2(new_n6356_), .ZN(new_n34581_));
  NAND2_X1   g32145(.A1(new_n34581_), .A2(new_n6352_), .ZN(new_n34582_));
  AOI21_X1   g32146(.A1(new_n34578_), .A2(new_n34582_), .B(new_n34577_), .ZN(new_n34583_));
  OAI21_X1   g32147(.A1(new_n34583_), .A2(new_n34575_), .B(new_n7253_), .ZN(new_n34584_));
  INV_X1     g32148(.I(pi0783), .ZN(new_n34585_));
  NAND2_X1   g32149(.A1(new_n34585_), .A2(pi1135), .ZN(new_n34586_));
  NAND2_X1   g32150(.A1(new_n32939_), .A2(new_n4888_), .ZN(new_n34587_));
  AOI21_X1   g32151(.A1(new_n34587_), .A2(new_n34586_), .B(pi1136), .ZN(new_n34588_));
  NAND2_X1   g32152(.A1(new_n25973_), .A2(new_n4888_), .ZN(new_n34589_));
  NAND2_X1   g32153(.A1(new_n25966_), .A2(pi1135), .ZN(new_n34590_));
  AOI21_X1   g32154(.A1(new_n34589_), .A2(new_n34590_), .B(new_n4724_), .ZN(new_n34591_));
  OAI21_X1   g32155(.A1(new_n34588_), .A2(new_n34591_), .B(new_n5045_), .ZN(new_n34592_));
  NOR2_X1    g32156(.A1(new_n14304_), .A2(pi1135), .ZN(new_n34593_));
  AOI21_X1   g32157(.A1(pi0735), .A2(pi1135), .B(new_n34593_), .ZN(new_n34594_));
  AOI21_X1   g32158(.A1(new_n34411_), .A2(pi0859), .B(new_n5045_), .ZN(new_n34595_));
  OAI21_X1   g32159(.A1(new_n34594_), .A2(new_n4724_), .B(new_n34595_), .ZN(new_n34596_));
  NAND3_X1   g32160(.A1(new_n34592_), .A2(new_n34596_), .A3(new_n34414_), .ZN(new_n34597_));
  NAND2_X1   g32161(.A1(new_n34584_), .A2(new_n34597_), .ZN(po0831));
  INV_X1     g32162(.I(pi0876), .ZN(new_n34599_));
  INV_X1     g32163(.I(new_n34411_), .ZN(new_n34600_));
  NOR2_X1    g32164(.A1(new_n17036_), .A2(pi1135), .ZN(new_n34601_));
  AOI21_X1   g32165(.A1(pi0730), .A2(pi1135), .B(new_n34601_), .ZN(new_n34602_));
  OAI22_X1   g32166(.A1(new_n34602_), .A2(new_n4724_), .B1(new_n34599_), .B2(new_n34600_), .ZN(new_n34603_));
  NOR2_X1    g32167(.A1(pi0803), .A2(pi1135), .ZN(new_n34604_));
  OAI22_X1   g32168(.A1(new_n34604_), .A2(pi1136), .B1(pi0710), .B2(new_n4888_), .ZN(new_n34605_));
  NAND2_X1   g32169(.A1(new_n34350_), .A2(pi0789), .ZN(new_n34606_));
  AOI21_X1   g32170(.A1(new_n34606_), .A2(new_n34605_), .B(new_n34358_), .ZN(new_n34607_));
  NAND2_X1   g32171(.A1(new_n34353_), .A2(new_n25648_), .ZN(new_n34608_));
  AOI22_X1   g32172(.A1(new_n34607_), .A2(new_n34608_), .B1(new_n34349_), .B2(new_n34603_), .ZN(new_n34609_));
  NAND2_X1   g32173(.A1(new_n34370_), .A2(pi0436), .ZN(new_n34610_));
  AOI21_X1   g32174(.A1(new_n34610_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34611_));
  NAND3_X1   g32175(.A1(new_n6352_), .A2(pi0412), .A3(pi0591), .ZN(new_n34612_));
  NAND2_X1   g32176(.A1(new_n6440_), .A2(pi0388), .ZN(new_n34613_));
  AOI22_X1   g32177(.A1(new_n34393_), .A2(new_n34612_), .B1(new_n34613_), .B2(pi0592), .ZN(new_n34614_));
  NOR2_X1    g32178(.A1(new_n34433_), .A2(new_n6488_), .ZN(new_n34615_));
  OAI21_X1   g32179(.A1(new_n34614_), .A2(new_n34615_), .B(new_n34611_), .ZN(new_n34616_));
  NAND2_X1   g32180(.A1(new_n8525_), .A2(pi0296), .ZN(new_n34617_));
  OAI21_X1   g32181(.A1(new_n8525_), .A2(new_n32493_), .B(new_n34617_), .ZN(new_n34618_));
  AOI21_X1   g32182(.A1(new_n34618_), .A2(new_n34369_), .B(new_n10920_), .ZN(new_n34619_));
  AOI22_X1   g32183(.A1(new_n10920_), .A2(new_n34609_), .B1(new_n34616_), .B2(new_n34619_), .ZN(po0832));
  OAI22_X1   g32184(.A1(new_n4888_), .A2(pi0729), .B1(pi0881), .B2(pi1136), .ZN(new_n34621_));
  NOR2_X1    g32185(.A1(new_n34354_), .A2(pi0746), .ZN(new_n34622_));
  NOR3_X1    g32186(.A1(new_n34622_), .A2(new_n34352_), .A3(new_n34621_), .ZN(new_n34623_));
  NOR2_X1    g32187(.A1(new_n25167_), .A2(new_n4888_), .ZN(new_n34624_));
  NOR2_X1    g32188(.A1(new_n25131_), .A2(pi1135), .ZN(new_n34625_));
  OAI21_X1   g32189(.A1(new_n34624_), .A2(new_n34625_), .B(pi1136), .ZN(new_n34626_));
  NOR2_X1    g32190(.A1(pi0812), .A2(pi1135), .ZN(new_n34627_));
  NOR2_X1    g32191(.A1(new_n12972_), .A2(new_n4888_), .ZN(new_n34628_));
  OAI21_X1   g32192(.A1(new_n34628_), .A2(new_n34627_), .B(new_n4724_), .ZN(new_n34629_));
  AOI21_X1   g32193(.A1(new_n34626_), .A2(new_n34629_), .B(new_n34358_), .ZN(new_n34630_));
  NOR3_X1    g32194(.A1(new_n34623_), .A2(new_n34630_), .A3(new_n7253_), .ZN(new_n34631_));
  NAND2_X1   g32195(.A1(new_n34370_), .A2(pi0434), .ZN(new_n34632_));
  AOI21_X1   g32196(.A1(new_n34632_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34633_));
  NOR3_X1    g32197(.A1(new_n32825_), .A2(new_n6440_), .A3(pi0590), .ZN(new_n34634_));
  NOR2_X1    g32198(.A1(new_n34394_), .A2(new_n34634_), .ZN(new_n34635_));
  AOI21_X1   g32199(.A1(pi0386), .A2(new_n6440_), .B(new_n6268_), .ZN(new_n34636_));
  OAI22_X1   g32200(.A1(new_n34635_), .A2(new_n34636_), .B1(new_n32707_), .B2(new_n34433_), .ZN(new_n34637_));
  NOR2_X1    g32201(.A1(new_n8525_), .A2(new_n32484_), .ZN(new_n34638_));
  AOI21_X1   g32202(.A1(new_n8525_), .A2(pi0293), .B(new_n34638_), .ZN(new_n34639_));
  OAI21_X1   g32203(.A1(new_n34639_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34640_));
  AOI21_X1   g32204(.A1(new_n34637_), .A2(new_n34633_), .B(new_n34640_), .ZN(new_n34641_));
  NOR2_X1    g32205(.A1(new_n34641_), .A2(new_n34631_), .ZN(po0833));
  OAI22_X1   g32206(.A1(new_n16429_), .A2(new_n4888_), .B1(pi0870), .B2(pi1136), .ZN(new_n34643_));
  NOR2_X1    g32207(.A1(new_n34354_), .A2(new_n16430_), .ZN(new_n34644_));
  NOR3_X1    g32208(.A1(new_n34644_), .A2(new_n34352_), .A3(new_n34643_), .ZN(new_n34645_));
  NOR2_X1    g32209(.A1(new_n4888_), .A2(pi0635), .ZN(new_n34646_));
  AOI21_X1   g32210(.A1(pi0620), .A2(new_n4888_), .B(new_n34646_), .ZN(new_n34647_));
  NOR3_X1    g32211(.A1(new_n34647_), .A2(pi1134), .A3(new_n34498_), .ZN(new_n34648_));
  NOR3_X1    g32212(.A1(new_n34645_), .A2(new_n7253_), .A3(new_n34648_), .ZN(new_n34649_));
  NAND2_X1   g32213(.A1(new_n34370_), .A2(pi0416), .ZN(new_n34650_));
  AOI21_X1   g32214(.A1(new_n34650_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34651_));
  AOI21_X1   g32215(.A1(new_n34375_), .A2(pi0344), .B(pi0588), .ZN(new_n34652_));
  AOI22_X1   g32216(.A1(pi0335), .A2(new_n34378_), .B1(new_n34377_), .B2(pi0366), .ZN(new_n34653_));
  OAI21_X1   g32217(.A1(pi0590), .A2(new_n34653_), .B(new_n34652_), .ZN(new_n34654_));
  NOR2_X1    g32218(.A1(new_n31361_), .A2(pi0199), .ZN(new_n34655_));
  AOI21_X1   g32219(.A1(pi0199), .A2(pi1069), .B(new_n34655_), .ZN(new_n34656_));
  OAI21_X1   g32220(.A1(new_n34656_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34657_));
  AOI21_X1   g32221(.A1(new_n34654_), .A2(new_n34651_), .B(new_n34657_), .ZN(new_n34658_));
  NOR2_X1    g32222(.A1(new_n34658_), .A2(new_n34649_), .ZN(po0834));
  OAI22_X1   g32223(.A1(new_n16510_), .A2(new_n4888_), .B1(pi0856), .B2(pi1136), .ZN(new_n34660_));
  NOR2_X1    g32224(.A1(new_n34354_), .A2(new_n16512_), .ZN(new_n34661_));
  NOR3_X1    g32225(.A1(new_n34661_), .A2(new_n34352_), .A3(new_n34660_), .ZN(new_n34662_));
  NOR2_X1    g32226(.A1(new_n4888_), .A2(pi0632), .ZN(new_n34663_));
  AOI21_X1   g32227(.A1(pi0613), .A2(new_n4888_), .B(new_n34663_), .ZN(new_n34664_));
  NOR3_X1    g32228(.A1(new_n34664_), .A2(pi1134), .A3(new_n34498_), .ZN(new_n34665_));
  NOR3_X1    g32229(.A1(new_n34662_), .A2(new_n7253_), .A3(new_n34665_), .ZN(new_n34666_));
  NAND2_X1   g32230(.A1(new_n34370_), .A2(pi0418), .ZN(new_n34667_));
  AOI21_X1   g32231(.A1(new_n34667_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34668_));
  AOI21_X1   g32232(.A1(new_n34375_), .A2(pi0346), .B(pi0588), .ZN(new_n34669_));
  AOI22_X1   g32233(.A1(pi0368), .A2(new_n34377_), .B1(new_n34378_), .B2(pi0393), .ZN(new_n34670_));
  OAI21_X1   g32234(.A1(pi0590), .A2(new_n34670_), .B(new_n34669_), .ZN(new_n34671_));
  NOR2_X1    g32235(.A1(new_n31367_), .A2(pi0199), .ZN(new_n34672_));
  AOI21_X1   g32236(.A1(pi0199), .A2(pi1067), .B(new_n34672_), .ZN(new_n34673_));
  OAI21_X1   g32237(.A1(new_n34673_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34674_));
  AOI21_X1   g32238(.A1(new_n34671_), .A2(new_n34668_), .B(new_n34674_), .ZN(new_n34675_));
  NOR2_X1    g32239(.A1(new_n34675_), .A2(new_n34666_), .ZN(po0835));
  OAI22_X1   g32240(.A1(new_n4888_), .A2(pi0690), .B1(pi0874), .B2(pi1136), .ZN(new_n34677_));
  NOR2_X1    g32241(.A1(new_n34354_), .A2(pi0739), .ZN(new_n34678_));
  NOR3_X1    g32242(.A1(new_n34678_), .A2(new_n34352_), .A3(new_n34677_), .ZN(new_n34679_));
  NOR2_X1    g32243(.A1(new_n12822_), .A2(new_n4724_), .ZN(new_n34680_));
  INV_X1     g32244(.I(pi0791), .ZN(new_n34681_));
  NOR2_X1    g32245(.A1(new_n34681_), .A2(pi1136), .ZN(new_n34682_));
  OAI21_X1   g32246(.A1(new_n34680_), .A2(new_n34682_), .B(pi1135), .ZN(new_n34683_));
  NOR2_X1    g32247(.A1(new_n12752_), .A2(new_n4724_), .ZN(new_n34684_));
  NOR2_X1    g32248(.A1(new_n32940_), .A2(pi1136), .ZN(new_n34685_));
  OAI21_X1   g32249(.A1(new_n34684_), .A2(new_n34685_), .B(new_n4888_), .ZN(new_n34686_));
  AOI21_X1   g32250(.A1(new_n34683_), .A2(new_n34686_), .B(new_n34358_), .ZN(new_n34687_));
  NOR3_X1    g32251(.A1(new_n34679_), .A2(new_n34687_), .A3(new_n7253_), .ZN(new_n34688_));
  NAND2_X1   g32252(.A1(new_n34370_), .A2(pi0438), .ZN(new_n34689_));
  AOI21_X1   g32253(.A1(new_n34689_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34690_));
  AOI21_X1   g32254(.A1(new_n34375_), .A2(pi0450), .B(pi0588), .ZN(new_n34691_));
  AOI22_X1   g32255(.A1(pi0389), .A2(new_n34377_), .B1(new_n34378_), .B2(pi0413), .ZN(new_n34692_));
  OAI21_X1   g32256(.A1(pi0590), .A2(new_n34692_), .B(new_n34691_), .ZN(new_n34693_));
  NOR2_X1    g32257(.A1(new_n31337_), .A2(pi0199), .ZN(new_n34694_));
  AOI21_X1   g32258(.A1(pi0199), .A2(pi1036), .B(new_n34694_), .ZN(new_n34695_));
  OAI21_X1   g32259(.A1(new_n34695_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34696_));
  AOI21_X1   g32260(.A1(new_n34693_), .A2(new_n34690_), .B(new_n34696_), .ZN(new_n34697_));
  NOR2_X1    g32261(.A1(new_n34697_), .A2(new_n34688_), .ZN(po0836));
  NAND2_X1   g32262(.A1(po0954), .A2(pi1100), .ZN(new_n34699_));
  NAND2_X1   g32263(.A1(new_n34229_), .A2(pi0680), .ZN(new_n34700_));
  AOI21_X1   g32264(.A1(new_n34700_), .A2(new_n34699_), .B(pi0962), .ZN(po0837));
  NAND2_X1   g32265(.A1(po0954), .A2(pi1103), .ZN(new_n34702_));
  NAND2_X1   g32266(.A1(new_n34229_), .A2(pi0681), .ZN(new_n34703_));
  AOI21_X1   g32267(.A1(new_n34703_), .A2(new_n34702_), .B(pi0962), .ZN(po0838));
  OAI22_X1   g32268(.A1(new_n16459_), .A2(new_n4888_), .B1(pi0848), .B2(pi1136), .ZN(new_n34705_));
  NOR2_X1    g32269(.A1(new_n34354_), .A2(new_n16460_), .ZN(new_n34706_));
  NOR3_X1    g32270(.A1(new_n34706_), .A2(new_n34352_), .A3(new_n34705_), .ZN(new_n34707_));
  NOR2_X1    g32271(.A1(new_n4888_), .A2(pi0631), .ZN(new_n34708_));
  AOI21_X1   g32272(.A1(pi0610), .A2(new_n4888_), .B(new_n34708_), .ZN(new_n34709_));
  NOR3_X1    g32273(.A1(new_n34709_), .A2(pi1134), .A3(new_n34498_), .ZN(new_n34710_));
  NOR3_X1    g32274(.A1(new_n34707_), .A2(new_n7253_), .A3(new_n34710_), .ZN(new_n34711_));
  NAND2_X1   g32275(.A1(new_n34370_), .A2(pi0417), .ZN(new_n34712_));
  AOI21_X1   g32276(.A1(new_n34712_), .A2(pi0588), .B(new_n34369_), .ZN(new_n34713_));
  AOI21_X1   g32277(.A1(new_n34375_), .A2(pi0345), .B(pi0588), .ZN(new_n34714_));
  AOI22_X1   g32278(.A1(pi0367), .A2(new_n34377_), .B1(new_n34378_), .B2(pi0392), .ZN(new_n34715_));
  OAI21_X1   g32279(.A1(pi0590), .A2(new_n34715_), .B(new_n34714_), .ZN(new_n34716_));
  NOR2_X1    g32280(.A1(new_n30993_), .A2(pi0199), .ZN(new_n34717_));
  AOI21_X1   g32281(.A1(pi0199), .A2(pi1039), .B(new_n34717_), .ZN(new_n34718_));
  OAI21_X1   g32282(.A1(new_n34718_), .A2(new_n34368_), .B(new_n7253_), .ZN(new_n34719_));
  AOI21_X1   g32283(.A1(new_n34716_), .A2(new_n34713_), .B(new_n34719_), .ZN(new_n34720_));
  NOR2_X1    g32284(.A1(new_n34720_), .A2(new_n34711_), .ZN(po0839));
  INV_X1     g32285(.I(pi0684), .ZN(new_n34722_));
  NAND3_X1   g32286(.A1(new_n34224_), .A2(pi0953), .A3(new_n34225_), .ZN(new_n34723_));
  NAND2_X1   g32287(.A1(new_n34723_), .A2(new_n34722_), .ZN(new_n34724_));
  INV_X1     g32288(.I(new_n34723_), .ZN(po0980));
  NAND2_X1   g32289(.A1(po0980), .A2(pi1130), .ZN(new_n34726_));
  AOI21_X1   g32290(.A1(new_n34726_), .A2(new_n34724_), .B(pi0962), .ZN(po0841));
  AOI21_X1   g32291(.A1(pi0199), .A2(new_n32697_), .B(new_n34368_), .ZN(new_n34728_));
  NOR2_X1    g32292(.A1(new_n6251_), .A2(pi0590), .ZN(new_n34729_));
  NAND2_X1   g32293(.A1(new_n34729_), .A2(new_n34373_), .ZN(new_n34730_));
  NAND3_X1   g32294(.A1(new_n6352_), .A2(new_n6268_), .A3(pi0591), .ZN(new_n34731_));
  NOR2_X1    g32295(.A1(new_n6352_), .A2(pi0592), .ZN(new_n34732_));
  AOI22_X1   g32296(.A1(pi0357), .A2(new_n34732_), .B1(new_n34392_), .B2(pi0382), .ZN(new_n34733_));
  OAI22_X1   g32297(.A1(new_n34733_), .A2(pi0591), .B1(new_n32814_), .B2(new_n34731_), .ZN(new_n34734_));
  NAND2_X1   g32298(.A1(new_n34734_), .A2(new_n6251_), .ZN(new_n34735_));
  OAI21_X1   g32299(.A1(new_n6335_), .A2(new_n34730_), .B(new_n34735_), .ZN(new_n34736_));
  AOI22_X1   g32300(.A1(new_n34736_), .A2(new_n34368_), .B1(new_n31370_), .B2(new_n34728_), .ZN(new_n34737_));
  INV_X1     g32301(.I(new_n34349_), .ZN(new_n34738_));
  NOR2_X1    g32302(.A1(new_n4888_), .A2(pi0728), .ZN(new_n34739_));
  NOR2_X1    g32303(.A1(pi0744), .A2(pi1135), .ZN(new_n34740_));
  OAI21_X1   g32304(.A1(new_n34739_), .A2(new_n34740_), .B(pi1136), .ZN(new_n34741_));
  NAND2_X1   g32305(.A1(new_n34411_), .A2(pi0860), .ZN(new_n34742_));
  AOI21_X1   g32306(.A1(new_n34741_), .A2(new_n34742_), .B(new_n34738_), .ZN(new_n34743_));
  NAND2_X1   g32307(.A1(new_n4888_), .A2(pi0652), .ZN(new_n34744_));
  OAI21_X1   g32308(.A1(pi0657), .A2(new_n4888_), .B(new_n34744_), .ZN(new_n34745_));
  INV_X1     g32309(.I(pi0813), .ZN(new_n34746_));
  NOR2_X1    g32310(.A1(new_n34348_), .A2(new_n34746_), .ZN(new_n34747_));
  AOI22_X1   g32311(.A1(new_n34745_), .A2(pi1136), .B1(new_n34747_), .B2(new_n34411_), .ZN(new_n34748_));
  NOR2_X1    g32312(.A1(new_n34347_), .A2(new_n4724_), .ZN(new_n34749_));
  NOR3_X1    g32313(.A1(new_n34748_), .A2(pi1134), .A3(new_n34749_), .ZN(new_n34750_));
  NOR3_X1    g32314(.A1(new_n34750_), .A2(new_n7253_), .A3(new_n34743_), .ZN(new_n34751_));
  AOI21_X1   g32315(.A1(new_n34737_), .A2(new_n7253_), .B(new_n34751_), .ZN(po0842));
  NAND2_X1   g32316(.A1(new_n34723_), .A2(new_n16459_), .ZN(new_n34753_));
  NAND2_X1   g32317(.A1(po0980), .A2(pi1113), .ZN(new_n34754_));
  AOI21_X1   g32318(.A1(new_n34754_), .A2(new_n34753_), .B(pi0962), .ZN(po0843));
  NAND2_X1   g32319(.A1(po0980), .A2(pi1127), .ZN(new_n34756_));
  NAND2_X1   g32320(.A1(new_n34723_), .A2(pi0687), .ZN(new_n34757_));
  AOI21_X1   g32321(.A1(new_n34756_), .A2(new_n34757_), .B(pi0962), .ZN(po0844));
  NAND2_X1   g32322(.A1(new_n34723_), .A2(new_n16510_), .ZN(new_n34759_));
  NAND2_X1   g32323(.A1(po0980), .A2(pi1115), .ZN(new_n34760_));
  AOI21_X1   g32324(.A1(new_n34760_), .A2(new_n34759_), .B(pi0962), .ZN(po0845));
  NAND2_X1   g32325(.A1(new_n31340_), .A2(new_n8525_), .ZN(new_n34762_));
  NAND2_X1   g32326(.A1(pi0199), .A2(pi1079), .ZN(new_n34763_));
  AOI21_X1   g32327(.A1(new_n34762_), .A2(new_n34763_), .B(new_n34368_), .ZN(new_n34764_));
  AOI22_X1   g32328(.A1(pi0351), .A2(new_n34732_), .B1(new_n34392_), .B2(pi0376), .ZN(new_n34765_));
  OAI22_X1   g32329(.A1(new_n34765_), .A2(pi0591), .B1(new_n32800_), .B2(new_n34731_), .ZN(new_n34766_));
  NAND2_X1   g32330(.A1(new_n34766_), .A2(new_n6251_), .ZN(new_n34767_));
  OAI21_X1   g32331(.A1(new_n32868_), .A2(new_n34730_), .B(new_n34767_), .ZN(new_n34768_));
  AOI21_X1   g32332(.A1(new_n34768_), .A2(new_n34368_), .B(new_n34764_), .ZN(new_n34769_));
  OAI22_X1   g32333(.A1(new_n4888_), .A2(pi0703), .B1(pi0843), .B2(pi1136), .ZN(new_n34770_));
  NOR2_X1    g32334(.A1(new_n34354_), .A2(new_n16803_), .ZN(new_n34771_));
  NOR3_X1    g32335(.A1(new_n34771_), .A2(new_n34352_), .A3(new_n34770_), .ZN(new_n34772_));
  NOR2_X1    g32336(.A1(new_n4888_), .A2(pi0655), .ZN(new_n34773_));
  INV_X1     g32337(.I(pi0658), .ZN(new_n34774_));
  NOR2_X1    g32338(.A1(new_n34774_), .A2(pi1135), .ZN(new_n34775_));
  OAI21_X1   g32339(.A1(new_n34773_), .A2(new_n34775_), .B(pi1136), .ZN(new_n34776_));
  NAND2_X1   g32340(.A1(new_n34411_), .A2(pi0798), .ZN(new_n34777_));
  AOI21_X1   g32341(.A1(new_n34776_), .A2(new_n34777_), .B(new_n34358_), .ZN(new_n34778_));
  NOR3_X1    g32342(.A1(new_n34772_), .A2(new_n34778_), .A3(new_n7253_), .ZN(new_n34779_));
  AOI21_X1   g32343(.A1(new_n34769_), .A2(new_n7253_), .B(new_n34779_), .ZN(po0846));
  NAND2_X1   g32344(.A1(po0980), .A2(pi1108), .ZN(new_n34781_));
  NAND2_X1   g32345(.A1(new_n34723_), .A2(pi0690), .ZN(new_n34782_));
  AOI21_X1   g32346(.A1(new_n34781_), .A2(new_n34782_), .B(pi0962), .ZN(po0847));
  NAND2_X1   g32347(.A1(po0980), .A2(pi1107), .ZN(new_n34784_));
  NAND2_X1   g32348(.A1(new_n34723_), .A2(pi0691), .ZN(new_n34785_));
  AOI21_X1   g32349(.A1(new_n34784_), .A2(new_n34785_), .B(pi0962), .ZN(po0848));
  NOR2_X1    g32350(.A1(pi0770), .A2(pi1135), .ZN(new_n34787_));
  AOI21_X1   g32351(.A1(pi0726), .A2(pi1135), .B(new_n34787_), .ZN(new_n34788_));
  AOI21_X1   g32352(.A1(new_n34411_), .A2(pi0844), .B(new_n5045_), .ZN(new_n34789_));
  OAI21_X1   g32353(.A1(new_n34788_), .A2(new_n4724_), .B(new_n34789_), .ZN(new_n34790_));
  NOR2_X1    g32354(.A1(new_n4888_), .A2(pi0649), .ZN(new_n34791_));
  AOI21_X1   g32355(.A1(pi0656), .A2(new_n4888_), .B(new_n34791_), .ZN(new_n34792_));
  AOI21_X1   g32356(.A1(new_n34411_), .A2(pi0801), .B(pi1134), .ZN(new_n34793_));
  OAI21_X1   g32357(.A1(new_n34792_), .A2(new_n4724_), .B(new_n34793_), .ZN(new_n34794_));
  NAND3_X1   g32358(.A1(new_n34794_), .A2(new_n34414_), .A3(new_n34790_), .ZN(new_n34795_));
  NAND2_X1   g32359(.A1(new_n31352_), .A2(new_n8525_), .ZN(new_n34796_));
  NAND2_X1   g32360(.A1(pi0199), .A2(pi1078), .ZN(new_n34797_));
  AOI21_X1   g32361(.A1(new_n34796_), .A2(new_n34797_), .B(new_n34368_), .ZN(new_n34798_));
  AOI22_X1   g32362(.A1(pi0317), .A2(new_n34392_), .B1(new_n34732_), .B2(pi0352), .ZN(new_n34799_));
  OAI22_X1   g32363(.A1(new_n34799_), .A2(pi0591), .B1(new_n32803_), .B2(new_n34731_), .ZN(new_n34800_));
  NAND2_X1   g32364(.A1(new_n34800_), .A2(new_n6251_), .ZN(new_n34801_));
  OAI21_X1   g32365(.A1(new_n32871_), .A2(new_n34730_), .B(new_n34801_), .ZN(new_n34802_));
  AOI21_X1   g32366(.A1(new_n34802_), .A2(new_n34368_), .B(new_n34798_), .ZN(new_n34803_));
  OAI21_X1   g32367(.A1(new_n34803_), .A2(new_n10920_), .B(new_n34795_), .ZN(po0849));
  OR2_X2     g32368(.A1(po0954), .A2(pi0693), .Z(new_n34805_));
  NAND2_X1   g32369(.A1(po0954), .A2(pi1129), .ZN(new_n34806_));
  AOI21_X1   g32370(.A1(new_n34805_), .A2(new_n34806_), .B(pi0962), .ZN(po0850));
  INV_X1     g32371(.I(pi0694), .ZN(new_n34808_));
  NAND2_X1   g32372(.A1(new_n34723_), .A2(new_n34808_), .ZN(new_n34809_));
  NAND2_X1   g32373(.A1(po0980), .A2(pi1128), .ZN(new_n34810_));
  AOI21_X1   g32374(.A1(new_n34810_), .A2(new_n34809_), .B(pi0962), .ZN(po0851));
  NAND2_X1   g32375(.A1(new_n34229_), .A2(new_n26376_), .ZN(new_n34812_));
  NAND2_X1   g32376(.A1(po0954), .A2(pi1111), .ZN(new_n34813_));
  AOI21_X1   g32377(.A1(new_n34812_), .A2(new_n34813_), .B(pi0962), .ZN(po0852));
  NAND2_X1   g32378(.A1(po0980), .A2(pi1100), .ZN(new_n34815_));
  NAND2_X1   g32379(.A1(new_n34723_), .A2(pi0696), .ZN(new_n34816_));
  AOI21_X1   g32380(.A1(new_n34815_), .A2(new_n34816_), .B(pi0962), .ZN(po0853));
  INV_X1     g32381(.I(pi0697), .ZN(new_n34818_));
  NAND2_X1   g32382(.A1(new_n34723_), .A2(new_n34818_), .ZN(new_n34819_));
  NAND2_X1   g32383(.A1(po0980), .A2(pi1129), .ZN(new_n34820_));
  AOI21_X1   g32384(.A1(new_n34820_), .A2(new_n34819_), .B(pi0962), .ZN(po0854));
  NAND2_X1   g32385(.A1(new_n34723_), .A2(new_n15577_), .ZN(new_n34822_));
  NAND2_X1   g32386(.A1(po0980), .A2(pi1116), .ZN(new_n34823_));
  AOI21_X1   g32387(.A1(new_n34823_), .A2(new_n34822_), .B(pi0962), .ZN(po0855));
  NAND2_X1   g32388(.A1(po0980), .A2(pi1103), .ZN(new_n34825_));
  NAND2_X1   g32389(.A1(new_n34723_), .A2(pi0699), .ZN(new_n34826_));
  AOI21_X1   g32390(.A1(new_n34825_), .A2(new_n34826_), .B(pi0962), .ZN(po0856));
  NAND2_X1   g32391(.A1(po0980), .A2(pi1110), .ZN(new_n34828_));
  NAND2_X1   g32392(.A1(new_n34723_), .A2(pi0700), .ZN(new_n34829_));
  AOI21_X1   g32393(.A1(new_n34828_), .A2(new_n34829_), .B(pi0962), .ZN(po0857));
  NAND2_X1   g32394(.A1(new_n34723_), .A2(new_n16218_), .ZN(new_n34831_));
  NAND2_X1   g32395(.A1(po0980), .A2(pi1123), .ZN(new_n34832_));
  AOI21_X1   g32396(.A1(new_n34832_), .A2(new_n34831_), .B(pi0962), .ZN(po0858));
  NAND2_X1   g32397(.A1(new_n34723_), .A2(new_n16558_), .ZN(new_n34834_));
  NAND2_X1   g32398(.A1(po0980), .A2(pi1117), .ZN(new_n34835_));
  AOI21_X1   g32399(.A1(new_n34835_), .A2(new_n34834_), .B(pi0962), .ZN(po0859));
  NAND2_X1   g32400(.A1(po0980), .A2(pi1124), .ZN(new_n34837_));
  NAND2_X1   g32401(.A1(new_n34723_), .A2(pi0703), .ZN(new_n34838_));
  AOI21_X1   g32402(.A1(new_n34837_), .A2(new_n34838_), .B(pi0962), .ZN(po0860));
  NAND2_X1   g32403(.A1(new_n34723_), .A2(new_n16429_), .ZN(new_n34840_));
  NAND2_X1   g32404(.A1(po0980), .A2(pi1112), .ZN(new_n34841_));
  AOI21_X1   g32405(.A1(new_n34841_), .A2(new_n34840_), .B(pi0962), .ZN(po0861));
  NAND2_X1   g32406(.A1(po0980), .A2(pi1125), .ZN(new_n34843_));
  NAND2_X1   g32407(.A1(new_n34723_), .A2(pi0705), .ZN(new_n34844_));
  AOI21_X1   g32408(.A1(new_n34843_), .A2(new_n34844_), .B(pi0962), .ZN(po0862));
  NAND2_X1   g32409(.A1(po0980), .A2(pi1105), .ZN(new_n34846_));
  NAND2_X1   g32410(.A1(new_n34723_), .A2(pi0706), .ZN(new_n34847_));
  AOI21_X1   g32411(.A1(new_n34846_), .A2(new_n34847_), .B(pi0962), .ZN(po0863));
  NOR2_X1    g32412(.A1(new_n8525_), .A2(new_n32672_), .ZN(new_n34849_));
  NAND2_X1   g32413(.A1(new_n8531_), .A2(pi0304), .ZN(new_n34850_));
  OAI21_X1   g32414(.A1(new_n8531_), .A2(new_n32475_), .B(new_n34850_), .ZN(new_n34851_));
  AOI21_X1   g32415(.A1(new_n34851_), .A2(new_n8525_), .B(new_n34849_), .ZN(new_n34852_));
  NOR2_X1    g32416(.A1(new_n34389_), .A2(new_n34369_), .ZN(new_n34853_));
  INV_X1     g32417(.I(new_n34853_), .ZN(new_n34854_));
  NAND2_X1   g32418(.A1(pi0420), .A2(pi0588), .ZN(new_n34855_));
  OAI22_X1   g32419(.A1(new_n34854_), .A2(new_n34855_), .B1(new_n34368_), .B2(new_n34852_), .ZN(new_n34856_));
  OAI22_X1   g32420(.A1(new_n32727_), .A2(new_n34579_), .B1(new_n34580_), .B2(new_n32784_), .ZN(new_n34857_));
  AOI22_X1   g32421(.A1(new_n34857_), .A2(new_n6352_), .B1(pi0347), .B2(new_n34375_), .ZN(new_n34858_));
  NOR2_X1    g32422(.A1(new_n34369_), .A2(pi0588), .ZN(new_n34859_));
  INV_X1     g32423(.I(new_n34859_), .ZN(new_n34860_));
  NOR2_X1    g32424(.A1(new_n34858_), .A2(new_n34860_), .ZN(new_n34861_));
  NOR2_X1    g32425(.A1(new_n34856_), .A2(new_n34861_), .ZN(new_n34862_));
  OAI22_X1   g32426(.A1(new_n16558_), .A2(new_n4888_), .B1(pi0847), .B2(pi1136), .ZN(new_n34863_));
  NOR2_X1    g32427(.A1(new_n34354_), .A2(new_n16550_), .ZN(new_n34864_));
  NOR3_X1    g32428(.A1(new_n34864_), .A2(new_n34352_), .A3(new_n34863_), .ZN(new_n34865_));
  NOR2_X1    g32429(.A1(new_n12880_), .A2(new_n4888_), .ZN(new_n34866_));
  NOR2_X1    g32430(.A1(new_n12781_), .A2(pi1135), .ZN(new_n34867_));
  OAI21_X1   g32431(.A1(new_n34866_), .A2(new_n34867_), .B(new_n5045_), .ZN(new_n34868_));
  OAI21_X1   g32432(.A1(new_n34868_), .A2(new_n34498_), .B(new_n10920_), .ZN(new_n34869_));
  NOR2_X1    g32433(.A1(new_n34865_), .A2(new_n34869_), .ZN(new_n34870_));
  AOI21_X1   g32434(.A1(new_n34862_), .A2(new_n7253_), .B(new_n34870_), .ZN(po0864));
  NOR2_X1    g32435(.A1(new_n13829_), .A2(new_n4888_), .ZN(new_n34872_));
  NOR2_X1    g32436(.A1(new_n12766_), .A2(pi1135), .ZN(new_n34873_));
  OAI21_X1   g32437(.A1(new_n34872_), .A2(new_n34873_), .B(new_n5045_), .ZN(new_n34874_));
  OAI21_X1   g32438(.A1(new_n34874_), .A2(new_n34498_), .B(new_n10920_), .ZN(new_n34875_));
  NAND2_X1   g32439(.A1(new_n34351_), .A2(new_n34347_), .ZN(new_n34876_));
  OAI21_X1   g32440(.A1(pi0857), .A2(pi1136), .B(pi1134), .ZN(new_n34877_));
  NOR2_X1    g32441(.A1(new_n16593_), .A2(new_n4888_), .ZN(new_n34878_));
  NOR2_X1    g32442(.A1(new_n34354_), .A2(new_n16585_), .ZN(new_n34879_));
  NOR4_X1    g32443(.A1(new_n34879_), .A2(new_n34876_), .A3(new_n34877_), .A4(new_n34878_), .ZN(new_n34880_));
  NOR2_X1    g32444(.A1(new_n34880_), .A2(new_n34875_), .ZN(new_n34881_));
  NAND2_X1   g32445(.A1(new_n34375_), .A2(new_n34368_), .ZN(new_n34882_));
  OAI22_X1   g32446(.A1(new_n32618_), .A2(new_n34580_), .B1(new_n34579_), .B2(new_n6623_), .ZN(new_n34883_));
  NAND2_X1   g32447(.A1(new_n34883_), .A2(new_n34368_), .ZN(new_n34884_));
  OAI22_X1   g32448(.A1(new_n34884_), .A2(pi0590), .B1(new_n32599_), .B2(new_n34882_), .ZN(new_n34885_));
  NAND2_X1   g32449(.A1(new_n34885_), .A2(new_n6251_), .ZN(new_n34886_));
  NAND2_X1   g32450(.A1(pi0199), .A2(pi1058), .ZN(new_n34887_));
  NOR2_X1    g32451(.A1(new_n8531_), .A2(new_n32481_), .ZN(new_n34888_));
  AOI21_X1   g32452(.A1(new_n8531_), .A2(pi0305), .B(new_n34888_), .ZN(new_n34889_));
  OAI21_X1   g32453(.A1(new_n34889_), .A2(pi0199), .B(new_n34887_), .ZN(new_n34890_));
  NAND2_X1   g32454(.A1(new_n34368_), .A2(new_n34373_), .ZN(new_n34891_));
  NAND2_X1   g32455(.A1(new_n34729_), .A2(pi0459), .ZN(new_n34892_));
  OAI21_X1   g32456(.A1(new_n34892_), .A2(new_n34891_), .B(new_n7253_), .ZN(new_n34893_));
  AOI21_X1   g32457(.A1(new_n34890_), .A2(new_n34369_), .B(new_n34893_), .ZN(new_n34894_));
  AOI21_X1   g32458(.A1(new_n34886_), .A2(new_n34894_), .B(new_n34881_), .ZN(po0865));
  NAND2_X1   g32459(.A1(new_n34723_), .A2(new_n16593_), .ZN(new_n34896_));
  NAND2_X1   g32460(.A1(po0980), .A2(pi1118), .ZN(new_n34897_));
  AOI21_X1   g32461(.A1(new_n34897_), .A2(new_n34896_), .B(pi0962), .ZN(po0866));
  NAND2_X1   g32462(.A1(po0954), .A2(pi1106), .ZN(new_n34899_));
  NAND2_X1   g32463(.A1(new_n34229_), .A2(pi0710), .ZN(new_n34900_));
  AOI21_X1   g32464(.A1(new_n34900_), .A2(new_n34899_), .B(pi0962), .ZN(po0867));
  NOR2_X1    g32465(.A1(new_n8525_), .A2(new_n32675_), .ZN(new_n34902_));
  NAND2_X1   g32466(.A1(new_n8531_), .A2(pi0306), .ZN(new_n34903_));
  OAI21_X1   g32467(.A1(new_n8531_), .A2(new_n32484_), .B(new_n34903_), .ZN(new_n34904_));
  AOI21_X1   g32468(.A1(new_n34904_), .A2(new_n8525_), .B(new_n34902_), .ZN(new_n34905_));
  NAND2_X1   g32469(.A1(pi0423), .A2(pi0588), .ZN(new_n34906_));
  OAI22_X1   g32470(.A1(new_n34854_), .A2(new_n34906_), .B1(new_n34368_), .B2(new_n34905_), .ZN(new_n34907_));
  OAI22_X1   g32471(.A1(new_n7234_), .A2(new_n34579_), .B1(new_n34580_), .B2(new_n32791_), .ZN(new_n34908_));
  AOI22_X1   g32472(.A1(new_n34908_), .A2(new_n6352_), .B1(pi0348), .B2(new_n34375_), .ZN(new_n34909_));
  NOR2_X1    g32473(.A1(new_n34909_), .A2(new_n34860_), .ZN(new_n34910_));
  NOR2_X1    g32474(.A1(new_n34907_), .A2(new_n34910_), .ZN(new_n34911_));
  OAI22_X1   g32475(.A1(new_n16168_), .A2(new_n4888_), .B1(pi0858), .B2(pi1136), .ZN(new_n34912_));
  NOR2_X1    g32476(.A1(new_n34354_), .A2(new_n16169_), .ZN(new_n34913_));
  NOR3_X1    g32477(.A1(new_n34913_), .A2(new_n34352_), .A3(new_n34912_), .ZN(new_n34914_));
  NOR2_X1    g32478(.A1(new_n12741_), .A2(new_n4888_), .ZN(new_n34915_));
  NOR2_X1    g32479(.A1(new_n12981_), .A2(pi1135), .ZN(new_n34916_));
  OAI21_X1   g32480(.A1(new_n34915_), .A2(new_n34916_), .B(new_n5045_), .ZN(new_n34917_));
  OAI21_X1   g32481(.A1(new_n34917_), .A2(new_n34498_), .B(new_n10920_), .ZN(new_n34918_));
  NOR2_X1    g32482(.A1(new_n34914_), .A2(new_n34918_), .ZN(new_n34919_));
  AOI21_X1   g32483(.A1(new_n34911_), .A2(new_n7253_), .B(new_n34919_), .ZN(po0868));
  INV_X1     g32484(.I(new_n34730_), .ZN(new_n34921_));
  OAI22_X1   g32485(.A1(new_n7051_), .A2(new_n34579_), .B1(new_n34580_), .B2(new_n32797_), .ZN(new_n34922_));
  AOI22_X1   g32486(.A1(new_n34922_), .A2(new_n6352_), .B1(pi0350), .B2(new_n34375_), .ZN(new_n34923_));
  OAI21_X1   g32487(.A1(new_n34923_), .A2(pi0588), .B(new_n34368_), .ZN(new_n34924_));
  AOI21_X1   g32488(.A1(pi0425), .A2(new_n34921_), .B(new_n34924_), .ZN(new_n34925_));
  AOI22_X1   g32489(.A1(new_n28112_), .A2(pi1044), .B1(pi0199), .B2(pi1035), .ZN(new_n34926_));
  NAND2_X1   g32490(.A1(new_n34926_), .A2(new_n34369_), .ZN(new_n34927_));
  AND2_X2    g32491(.A1(new_n8640_), .A2(pi0298), .Z(new_n34928_));
  OAI21_X1   g32492(.A1(new_n34927_), .A2(new_n34928_), .B(new_n7253_), .ZN(new_n34929_));
  OAI21_X1   g32493(.A1(pi0842), .A2(pi1136), .B(pi1134), .ZN(new_n34930_));
  NOR2_X1    g32494(.A1(new_n16218_), .A2(new_n4888_), .ZN(new_n34931_));
  NOR2_X1    g32495(.A1(new_n34354_), .A2(new_n16210_), .ZN(new_n34932_));
  NOR4_X1    g32496(.A1(new_n34932_), .A2(new_n34876_), .A3(new_n34930_), .A4(new_n34931_), .ZN(new_n34933_));
  NOR2_X1    g32497(.A1(new_n12975_), .A2(pi1135), .ZN(new_n34934_));
  AOI21_X1   g32498(.A1(pi0715), .A2(pi1135), .B(new_n34934_), .ZN(new_n34935_));
  NOR3_X1    g32499(.A1(new_n34935_), .A2(pi1134), .A3(new_n34498_), .ZN(new_n34936_));
  NOR2_X1    g32500(.A1(new_n34933_), .A2(new_n34936_), .ZN(new_n34937_));
  OAI22_X1   g32501(.A1(new_n34925_), .A2(new_n34929_), .B1(new_n7253_), .B2(new_n34937_), .ZN(po0869));
  INV_X1     g32502(.I(pi1051), .ZN(new_n34939_));
  NOR2_X1    g32503(.A1(new_n8525_), .A2(new_n34939_), .ZN(new_n34940_));
  NAND2_X1   g32504(.A1(new_n8531_), .A2(pi0309), .ZN(new_n34941_));
  OAI21_X1   g32505(.A1(new_n8531_), .A2(new_n32487_), .B(new_n34941_), .ZN(new_n34942_));
  AOI21_X1   g32506(.A1(new_n34942_), .A2(new_n8525_), .B(new_n34940_), .ZN(new_n34943_));
  NAND2_X1   g32507(.A1(pi0421), .A2(pi0588), .ZN(new_n34944_));
  OAI22_X1   g32508(.A1(new_n34854_), .A2(new_n34944_), .B1(new_n34368_), .B2(new_n34943_), .ZN(new_n34945_));
  OAI22_X1   g32509(.A1(new_n7049_), .A2(new_n34579_), .B1(new_n34580_), .B2(new_n6368_), .ZN(new_n34946_));
  AOI22_X1   g32510(.A1(new_n34946_), .A2(new_n6352_), .B1(pi0322), .B2(new_n34375_), .ZN(new_n34947_));
  NOR2_X1    g32511(.A1(new_n34947_), .A2(new_n34860_), .ZN(new_n34948_));
  NOR2_X1    g32512(.A1(new_n34945_), .A2(new_n34948_), .ZN(new_n34949_));
  OAI22_X1   g32513(.A1(new_n16620_), .A2(new_n4888_), .B1(pi0854), .B2(pi1136), .ZN(new_n34950_));
  NOR2_X1    g32514(.A1(new_n34354_), .A2(new_n16621_), .ZN(new_n34951_));
  NOR3_X1    g32515(.A1(new_n34951_), .A2(new_n34352_), .A3(new_n34950_), .ZN(new_n34952_));
  NOR2_X1    g32516(.A1(new_n12920_), .A2(new_n4888_), .ZN(new_n34953_));
  NOR2_X1    g32517(.A1(new_n12919_), .A2(pi1135), .ZN(new_n34954_));
  OAI21_X1   g32518(.A1(new_n34953_), .A2(new_n34954_), .B(new_n5045_), .ZN(new_n34955_));
  OAI21_X1   g32519(.A1(new_n34955_), .A2(new_n34498_), .B(new_n10920_), .ZN(new_n34956_));
  NOR2_X1    g32520(.A1(new_n34952_), .A2(new_n34956_), .ZN(new_n34957_));
  AOI21_X1   g32521(.A1(new_n34949_), .A2(new_n7253_), .B(new_n34957_), .ZN(po0870));
  AOI21_X1   g32522(.A1(pi0199), .A2(new_n32898_), .B(new_n34368_), .ZN(new_n34959_));
  AOI22_X1   g32523(.A1(pi0439), .A2(new_n34392_), .B1(new_n34732_), .B2(pi0461), .ZN(new_n34960_));
  OAI22_X1   g32524(.A1(new_n34960_), .A2(pi0591), .B1(new_n32611_), .B2(new_n34731_), .ZN(new_n34961_));
  NAND2_X1   g32525(.A1(new_n34961_), .A2(new_n6251_), .ZN(new_n34962_));
  OAI21_X1   g32526(.A1(new_n6324_), .A2(new_n34730_), .B(new_n34962_), .ZN(new_n34963_));
  AOI22_X1   g32527(.A1(new_n34963_), .A2(new_n34368_), .B1(new_n30999_), .B2(new_n34959_), .ZN(new_n34964_));
  NOR2_X1    g32528(.A1(new_n4888_), .A2(pi0697), .ZN(new_n34965_));
  NOR2_X1    g32529(.A1(pi0762), .A2(pi1135), .ZN(new_n34966_));
  OAI21_X1   g32530(.A1(new_n34965_), .A2(new_n34966_), .B(pi1136), .ZN(new_n34967_));
  NAND2_X1   g32531(.A1(new_n34411_), .A2(pi0867), .ZN(new_n34968_));
  AOI21_X1   g32532(.A1(new_n34967_), .A2(new_n34968_), .B(new_n34738_), .ZN(new_n34969_));
  NAND2_X1   g32533(.A1(new_n4888_), .A2(pi0653), .ZN(new_n34970_));
  OAI21_X1   g32534(.A1(pi0693), .A2(new_n4888_), .B(new_n34970_), .ZN(new_n34971_));
  INV_X1     g32535(.I(pi0816), .ZN(new_n34972_));
  NOR2_X1    g32536(.A1(new_n34348_), .A2(new_n34972_), .ZN(new_n34973_));
  AOI22_X1   g32537(.A1(new_n34971_), .A2(pi1136), .B1(new_n34973_), .B2(new_n34411_), .ZN(new_n34974_));
  NOR3_X1    g32538(.A1(new_n34974_), .A2(pi1134), .A3(new_n34749_), .ZN(new_n34975_));
  NOR3_X1    g32539(.A1(new_n34975_), .A2(new_n7253_), .A3(new_n34969_), .ZN(new_n34976_));
  AOI21_X1   g32540(.A1(new_n34964_), .A2(new_n7253_), .B(new_n34976_), .ZN(po0871));
  NAND2_X1   g32541(.A1(po0954), .A2(pi1123), .ZN(new_n34978_));
  NAND2_X1   g32542(.A1(new_n34229_), .A2(pi0715), .ZN(new_n34979_));
  AOI21_X1   g32543(.A1(new_n34979_), .A2(new_n34978_), .B(pi0962), .ZN(po0872));
  NOR2_X1    g32544(.A1(new_n12814_), .A2(new_n4888_), .ZN(new_n34981_));
  NOR2_X1    g32545(.A1(new_n12747_), .A2(pi1135), .ZN(new_n34982_));
  OAI21_X1   g32546(.A1(new_n34981_), .A2(new_n34982_), .B(new_n5045_), .ZN(new_n34983_));
  OAI21_X1   g32547(.A1(new_n34983_), .A2(new_n34498_), .B(new_n10920_), .ZN(new_n34984_));
  OAI21_X1   g32548(.A1(pi0845), .A2(pi1136), .B(pi1134), .ZN(new_n34985_));
  NOR2_X1    g32549(.A1(new_n12820_), .A2(new_n4888_), .ZN(new_n34986_));
  NOR2_X1    g32550(.A1(new_n34354_), .A2(new_n12750_), .ZN(new_n34987_));
  NOR4_X1    g32551(.A1(new_n34987_), .A2(new_n34876_), .A3(new_n34985_), .A4(new_n34986_), .ZN(new_n34988_));
  NOR2_X1    g32552(.A1(new_n34988_), .A2(new_n34984_), .ZN(new_n34989_));
  OAI22_X1   g32553(.A1(new_n32621_), .A2(new_n34580_), .B1(new_n34579_), .B2(new_n6622_), .ZN(new_n34990_));
  NAND2_X1   g32554(.A1(new_n34990_), .A2(new_n34368_), .ZN(new_n34991_));
  OAI22_X1   g32555(.A1(new_n34991_), .A2(pi0590), .B1(new_n32678_), .B2(new_n34882_), .ZN(new_n34992_));
  NAND2_X1   g32556(.A1(new_n34992_), .A2(new_n6251_), .ZN(new_n34993_));
  NAND2_X1   g32557(.A1(pi0199), .A2(pi1043), .ZN(new_n34994_));
  NOR2_X1    g32558(.A1(new_n8531_), .A2(new_n32490_), .ZN(new_n34995_));
  AOI21_X1   g32559(.A1(new_n8531_), .A2(pi0307), .B(new_n34995_), .ZN(new_n34996_));
  OAI21_X1   g32560(.A1(new_n34996_), .A2(pi0199), .B(new_n34994_), .ZN(new_n34997_));
  NAND2_X1   g32561(.A1(new_n34729_), .A2(pi0454), .ZN(new_n34998_));
  OAI21_X1   g32562(.A1(new_n34998_), .A2(new_n34891_), .B(new_n7253_), .ZN(new_n34999_));
  AOI21_X1   g32563(.A1(new_n34997_), .A2(new_n34369_), .B(new_n34999_), .ZN(new_n35000_));
  AOI21_X1   g32564(.A1(new_n34993_), .A2(new_n35000_), .B(new_n34989_), .ZN(po0873));
  INV_X1     g32565(.I(pi0800), .ZN(new_n35002_));
  NOR2_X1    g32566(.A1(new_n4888_), .A2(pi0669), .ZN(new_n35003_));
  AOI21_X1   g32567(.A1(pi0645), .A2(new_n4888_), .B(new_n35003_), .ZN(new_n35004_));
  OAI22_X1   g32568(.A1(new_n35004_), .A2(new_n4724_), .B1(new_n35002_), .B2(new_n34600_), .ZN(new_n35005_));
  NOR2_X1    g32569(.A1(pi0839), .A2(pi1136), .ZN(new_n35006_));
  NOR2_X1    g32570(.A1(new_n4888_), .A2(pi0705), .ZN(new_n35007_));
  NOR4_X1    g32571(.A1(new_n34876_), .A2(new_n5045_), .A3(new_n35006_), .A4(new_n35007_), .ZN(new_n35008_));
  NAND2_X1   g32572(.A1(new_n34353_), .A2(pi0768), .ZN(new_n35009_));
  AOI22_X1   g32573(.A1(new_n35008_), .A2(new_n35009_), .B1(new_n35005_), .B2(new_n34357_), .ZN(new_n35010_));
  NAND2_X1   g32574(.A1(new_n31346_), .A2(new_n8525_), .ZN(new_n35011_));
  NAND2_X1   g32575(.A1(pi0199), .A2(pi1074), .ZN(new_n35012_));
  AOI21_X1   g32576(.A1(new_n35011_), .A2(new_n35012_), .B(new_n34368_), .ZN(new_n35013_));
  NOR3_X1    g32577(.A1(new_n34854_), .A2(new_n9760_), .A3(new_n6251_), .ZN(new_n35014_));
  NOR3_X1    g32578(.A1(new_n35014_), .A2(new_n10920_), .A3(new_n35013_), .ZN(new_n35015_));
  AOI22_X1   g32579(.A1(pi0318), .A2(new_n34378_), .B1(new_n34377_), .B2(pi0377), .ZN(new_n35016_));
  OAI22_X1   g32580(.A1(new_n34433_), .A2(new_n6540_), .B1(new_n35016_), .B2(pi0590), .ZN(new_n35017_));
  NAND2_X1   g32581(.A1(new_n35017_), .A2(new_n34859_), .ZN(new_n35018_));
  AOI22_X1   g32582(.A1(new_n35015_), .A2(new_n35018_), .B1(new_n10920_), .B2(new_n35010_), .ZN(po0874));
  NOR2_X1    g32583(.A1(new_n13521_), .A2(new_n4888_), .ZN(new_n35020_));
  NOR2_X1    g32584(.A1(new_n13560_), .A2(pi1135), .ZN(new_n35021_));
  OAI21_X1   g32585(.A1(new_n35020_), .A2(new_n35021_), .B(new_n5045_), .ZN(new_n35022_));
  OAI21_X1   g32586(.A1(new_n35022_), .A2(new_n34498_), .B(new_n10920_), .ZN(new_n35023_));
  OAI21_X1   g32587(.A1(pi0853), .A2(pi1136), .B(pi1134), .ZN(new_n35024_));
  NOR2_X1    g32588(.A1(new_n15577_), .A2(new_n4888_), .ZN(new_n35025_));
  NOR2_X1    g32589(.A1(new_n34354_), .A2(new_n15782_), .ZN(new_n35026_));
  NOR4_X1    g32590(.A1(new_n35026_), .A2(new_n34876_), .A3(new_n35024_), .A4(new_n35025_), .ZN(new_n35027_));
  NOR2_X1    g32591(.A1(new_n35027_), .A2(new_n35023_), .ZN(new_n35028_));
  OAI22_X1   g32592(.A1(new_n9882_), .A2(new_n34579_), .B1(new_n34580_), .B2(new_n32781_), .ZN(new_n35029_));
  NAND2_X1   g32593(.A1(new_n35029_), .A2(new_n34368_), .ZN(new_n35030_));
  OAI22_X1   g32594(.A1(new_n35030_), .A2(pi0590), .B1(new_n6506_), .B2(new_n34882_), .ZN(new_n35031_));
  NAND2_X1   g32595(.A1(new_n35031_), .A2(new_n6251_), .ZN(new_n35032_));
  NAND2_X1   g32596(.A1(pi0199), .A2(pi1080), .ZN(new_n35033_));
  NOR2_X1    g32597(.A1(new_n8531_), .A2(new_n32478_), .ZN(new_n35034_));
  AOI21_X1   g32598(.A1(new_n8531_), .A2(pi0303), .B(new_n35034_), .ZN(new_n35035_));
  OAI21_X1   g32599(.A1(new_n35035_), .A2(pi0199), .B(new_n35033_), .ZN(new_n35036_));
  NAND2_X1   g32600(.A1(new_n34729_), .A2(pi0419), .ZN(new_n35037_));
  OAI21_X1   g32601(.A1(new_n35037_), .A2(new_n34891_), .B(new_n7253_), .ZN(new_n35038_));
  AOI21_X1   g32602(.A1(new_n35036_), .A2(new_n34369_), .B(new_n35038_), .ZN(new_n35039_));
  AOI21_X1   g32603(.A1(new_n35032_), .A2(new_n35039_), .B(new_n35028_), .ZN(po0875));
  INV_X1     g32604(.I(pi0807), .ZN(new_n35041_));
  NOR2_X1    g32605(.A1(new_n4888_), .A2(pi0650), .ZN(new_n35042_));
  AOI21_X1   g32606(.A1(pi0636), .A2(new_n4888_), .B(new_n35042_), .ZN(new_n35043_));
  OAI22_X1   g32607(.A1(new_n35043_), .A2(new_n4724_), .B1(new_n35041_), .B2(new_n34600_), .ZN(new_n35044_));
  NOR2_X1    g32608(.A1(pi0868), .A2(pi1136), .ZN(new_n35045_));
  NOR2_X1    g32609(.A1(new_n4888_), .A2(pi0687), .ZN(new_n35046_));
  NOR4_X1    g32610(.A1(new_n34876_), .A2(new_n5045_), .A3(new_n35045_), .A4(new_n35046_), .ZN(new_n35047_));
  NAND2_X1   g32611(.A1(new_n34353_), .A2(pi0774), .ZN(new_n35048_));
  AOI22_X1   g32612(.A1(new_n35047_), .A2(new_n35048_), .B1(new_n35044_), .B2(new_n34357_), .ZN(new_n35049_));
  NAND2_X1   g32613(.A1(new_n31358_), .A2(new_n8525_), .ZN(new_n35050_));
  NAND2_X1   g32614(.A1(pi0199), .A2(pi1063), .ZN(new_n35051_));
  AOI21_X1   g32615(.A1(new_n35050_), .A2(new_n35051_), .B(new_n34368_), .ZN(new_n35052_));
  NOR3_X1    g32616(.A1(new_n34854_), .A2(new_n6322_), .A3(new_n6251_), .ZN(new_n35053_));
  NOR3_X1    g32617(.A1(new_n35053_), .A2(new_n10920_), .A3(new_n35052_), .ZN(new_n35054_));
  AOI22_X1   g32618(.A1(pi0325), .A2(new_n34378_), .B1(new_n34377_), .B2(pi0378), .ZN(new_n35055_));
  OAI22_X1   g32619(.A1(new_n34433_), .A2(new_n32688_), .B1(new_n35055_), .B2(pi0590), .ZN(new_n35056_));
  NAND2_X1   g32620(.A1(new_n35056_), .A2(new_n34859_), .ZN(new_n35057_));
  AOI22_X1   g32621(.A1(new_n35054_), .A2(new_n35057_), .B1(new_n10920_), .B2(new_n35049_), .ZN(po0876));
  AOI21_X1   g32622(.A1(pi0199), .A2(new_n32753_), .B(new_n34368_), .ZN(new_n35059_));
  AOI22_X1   g32623(.A1(pi0356), .A2(new_n34732_), .B1(new_n34392_), .B2(pi0381), .ZN(new_n35060_));
  OAI22_X1   g32624(.A1(new_n35060_), .A2(pi0591), .B1(new_n32811_), .B2(new_n34731_), .ZN(new_n35061_));
  NAND2_X1   g32625(.A1(new_n35061_), .A2(new_n6251_), .ZN(new_n35062_));
  OAI21_X1   g32626(.A1(new_n6859_), .A2(new_n34730_), .B(new_n35062_), .ZN(new_n35063_));
  AOI22_X1   g32627(.A1(new_n35063_), .A2(new_n34368_), .B1(new_n31376_), .B2(new_n35059_), .ZN(new_n35064_));
  NOR2_X1    g32628(.A1(new_n4888_), .A2(pi0684), .ZN(new_n35065_));
  NOR2_X1    g32629(.A1(pi0750), .A2(pi1135), .ZN(new_n35066_));
  OAI21_X1   g32630(.A1(new_n35065_), .A2(new_n35066_), .B(pi1136), .ZN(new_n35067_));
  NAND2_X1   g32631(.A1(new_n34411_), .A2(pi0880), .ZN(new_n35068_));
  AOI21_X1   g32632(.A1(new_n35067_), .A2(new_n35068_), .B(new_n34738_), .ZN(new_n35069_));
  NAND2_X1   g32633(.A1(new_n4888_), .A2(pi0651), .ZN(new_n35070_));
  OAI21_X1   g32634(.A1(pi0654), .A2(new_n4888_), .B(new_n35070_), .ZN(new_n35071_));
  INV_X1     g32635(.I(pi0794), .ZN(new_n35072_));
  NOR2_X1    g32636(.A1(new_n34348_), .A2(new_n35072_), .ZN(new_n35073_));
  AOI22_X1   g32637(.A1(new_n35071_), .A2(pi1136), .B1(new_n35073_), .B2(new_n34411_), .ZN(new_n35074_));
  NOR3_X1    g32638(.A1(new_n35074_), .A2(pi1134), .A3(new_n34749_), .ZN(new_n35075_));
  NOR3_X1    g32639(.A1(new_n35075_), .A2(new_n7253_), .A3(new_n35069_), .ZN(new_n35076_));
  AOI21_X1   g32640(.A1(new_n35064_), .A2(new_n7253_), .B(new_n35076_), .ZN(po0877));
  INV_X1     g32641(.I(pi0731), .ZN(new_n35078_));
  INV_X1     g32642(.I(pi0945), .ZN(new_n35079_));
  NAND2_X1   g32643(.A1(new_n35079_), .A2(pi0988), .ZN(new_n35080_));
  NOR2_X1    g32644(.A1(new_n35080_), .A2(new_n35078_), .ZN(new_n35081_));
  INV_X1     g32645(.I(new_n35081_), .ZN(new_n35082_));
  NOR2_X1    g32646(.A1(pi0775), .A2(pi0816), .ZN(new_n35083_));
  INV_X1     g32647(.I(pi0775), .ZN(new_n35084_));
  NOR2_X1    g32648(.A1(new_n35084_), .A2(new_n34972_), .ZN(new_n35085_));
  NOR2_X1    g32649(.A1(new_n35085_), .A2(new_n35083_), .ZN(new_n35086_));
  XNOR2_X1   g32650(.A1(pi0771), .A2(pi0800), .ZN(new_n35087_));
  INV_X1     g32651(.I(new_n35087_), .ZN(new_n35088_));
  INV_X1     g32652(.I(pi0747), .ZN(new_n35089_));
  XOR2_X1    g32653(.A1(pi0765), .A2(pi0798), .Z(new_n35090_));
  NOR2_X1    g32654(.A1(new_n35090_), .A2(new_n35041_), .ZN(new_n35091_));
  INV_X1     g32655(.I(new_n35091_), .ZN(new_n35092_));
  NOR2_X1    g32656(.A1(new_n35092_), .A2(new_n35089_), .ZN(new_n35093_));
  NOR3_X1    g32657(.A1(new_n35090_), .A2(pi0747), .A3(pi0807), .ZN(new_n35094_));
  NOR2_X1    g32658(.A1(new_n35093_), .A2(new_n35094_), .ZN(new_n35095_));
  NOR2_X1    g32659(.A1(pi0769), .A2(pi0794), .ZN(new_n35096_));
  INV_X1     g32660(.I(pi0769), .ZN(new_n35097_));
  NOR2_X1    g32661(.A1(new_n35097_), .A2(new_n35072_), .ZN(new_n35098_));
  NOR2_X1    g32662(.A1(new_n35098_), .A2(new_n35096_), .ZN(new_n35099_));
  NOR2_X1    g32663(.A1(new_n35095_), .A2(new_n35099_), .ZN(new_n35100_));
  INV_X1     g32664(.I(new_n35100_), .ZN(new_n35101_));
  NOR2_X1    g32665(.A1(pi0773), .A2(pi0801), .ZN(new_n35102_));
  INV_X1     g32666(.I(pi0773), .ZN(new_n35103_));
  INV_X1     g32667(.I(pi0801), .ZN(new_n35104_));
  NOR2_X1    g32668(.A1(new_n35103_), .A2(new_n35104_), .ZN(new_n35105_));
  NOR2_X1    g32669(.A1(new_n35105_), .A2(new_n35102_), .ZN(new_n35106_));
  NOR3_X1    g32670(.A1(new_n35101_), .A2(new_n35088_), .A3(new_n35106_), .ZN(new_n35107_));
  INV_X1     g32671(.I(new_n35107_), .ZN(new_n35108_));
  INV_X1     g32672(.I(pi0721), .ZN(new_n35109_));
  NOR2_X1    g32673(.A1(new_n35109_), .A2(new_n34746_), .ZN(new_n35110_));
  INV_X1     g32674(.I(new_n35110_), .ZN(new_n35111_));
  NOR2_X1    g32675(.A1(new_n35108_), .A2(new_n35111_), .ZN(new_n35112_));
  INV_X1     g32676(.I(new_n35112_), .ZN(new_n35113_));
  NOR2_X1    g32677(.A1(new_n35113_), .A2(new_n35086_), .ZN(new_n35114_));
  XNOR2_X1   g32678(.A1(pi0731), .A2(pi0795), .ZN(new_n35115_));
  NAND2_X1   g32679(.A1(new_n35114_), .A2(new_n35115_), .ZN(new_n35116_));
  NAND3_X1   g32680(.A1(new_n35116_), .A2(pi0721), .A3(new_n35082_), .ZN(new_n35117_));
  INV_X1     g32681(.I(pi0795), .ZN(new_n35118_));
  NOR2_X1    g32682(.A1(new_n35089_), .A2(new_n35103_), .ZN(new_n35119_));
  AOI21_X1   g32683(.A1(new_n35119_), .A2(pi0769), .B(new_n35109_), .ZN(new_n35120_));
  INV_X1     g32684(.I(new_n35119_), .ZN(new_n35121_));
  NOR3_X1    g32685(.A1(new_n35121_), .A2(pi0721), .A3(new_n35097_), .ZN(new_n35122_));
  OAI21_X1   g32686(.A1(new_n35122_), .A2(new_n35120_), .B(pi0775), .ZN(new_n35123_));
  NAND2_X1   g32687(.A1(new_n35084_), .A2(pi0721), .ZN(new_n35124_));
  AOI21_X1   g32688(.A1(new_n35123_), .A2(new_n35124_), .B(new_n35082_), .ZN(new_n35125_));
  NOR2_X1    g32689(.A1(new_n35092_), .A2(new_n35088_), .ZN(new_n35126_));
  NOR2_X1    g32690(.A1(pi0721), .A2(pi0813), .ZN(new_n35127_));
  NAND4_X1   g32691(.A1(new_n35126_), .A2(pi0794), .A3(pi0801), .A4(new_n35127_), .ZN(new_n35128_));
  NAND2_X1   g32692(.A1(new_n35113_), .A2(new_n35128_), .ZN(new_n35129_));
  AOI21_X1   g32693(.A1(new_n35129_), .A2(pi0816), .B(new_n35123_), .ZN(new_n35130_));
  OAI21_X1   g32694(.A1(new_n35130_), .A2(new_n35118_), .B(new_n35125_), .ZN(new_n35131_));
  OR2_X2     g32695(.A1(new_n35114_), .A2(new_n35124_), .Z(new_n35132_));
  NAND3_X1   g32696(.A1(new_n35131_), .A2(new_n35117_), .A3(new_n35132_), .ZN(po0878));
  INV_X1     g32697(.I(pi1045), .ZN(new_n35134_));
  NOR2_X1    g32698(.A1(new_n8525_), .A2(new_n35134_), .ZN(new_n35135_));
  AOI21_X1   g32699(.A1(new_n31364_), .A2(new_n8525_), .B(new_n35135_), .ZN(new_n35136_));
  NAND2_X1   g32700(.A1(pi0428), .A2(pi0588), .ZN(new_n35137_));
  OAI22_X1   g32701(.A1(new_n34854_), .A2(new_n35137_), .B1(new_n34368_), .B2(new_n35136_), .ZN(new_n35138_));
  OAI22_X1   g32702(.A1(new_n32747_), .A2(new_n34579_), .B1(new_n34580_), .B2(new_n32806_), .ZN(new_n35139_));
  AOI22_X1   g32703(.A1(new_n35139_), .A2(new_n6352_), .B1(pi0354), .B2(new_n34375_), .ZN(new_n35140_));
  NOR2_X1    g32704(.A1(new_n35140_), .A2(new_n34860_), .ZN(new_n35141_));
  OAI21_X1   g32705(.A1(new_n35138_), .A2(new_n35141_), .B(new_n7253_), .ZN(new_n35142_));
  NAND2_X1   g32706(.A1(pi1135), .A2(pi1136), .ZN(new_n35143_));
  NAND2_X1   g32707(.A1(new_n34808_), .A2(pi1134), .ZN(new_n35144_));
  INV_X1     g32708(.I(pi0732), .ZN(new_n35145_));
  NAND2_X1   g32709(.A1(new_n35145_), .A2(new_n5045_), .ZN(new_n35146_));
  AOI21_X1   g32710(.A1(new_n35146_), .A2(new_n35144_), .B(new_n35143_), .ZN(new_n35147_));
  AND2_X2    g32711(.A1(pi0851), .A2(pi1134), .Z(new_n35148_));
  NOR2_X1    g32712(.A1(new_n35118_), .A2(pi1134), .ZN(new_n35149_));
  OAI21_X1   g32713(.A1(new_n35148_), .A2(new_n35149_), .B(new_n4724_), .ZN(new_n35150_));
  NOR2_X1    g32714(.A1(new_n5045_), .A2(pi0776), .ZN(new_n35151_));
  INV_X1     g32715(.I(pi0640), .ZN(new_n35152_));
  NOR2_X1    g32716(.A1(new_n35152_), .A2(pi1134), .ZN(new_n35153_));
  OAI21_X1   g32717(.A1(new_n35151_), .A2(new_n35153_), .B(pi1136), .ZN(new_n35154_));
  AOI21_X1   g32718(.A1(new_n35150_), .A2(new_n35154_), .B(pi1135), .ZN(new_n35155_));
  OAI21_X1   g32719(.A1(new_n35155_), .A2(new_n35147_), .B(new_n34414_), .ZN(new_n35156_));
  NAND2_X1   g32720(.A1(new_n35142_), .A2(new_n35156_), .ZN(po0879));
  NAND2_X1   g32721(.A1(new_n34723_), .A2(new_n16263_), .ZN(new_n35158_));
  NAND2_X1   g32722(.A1(po0980), .A2(pi1111), .ZN(new_n35159_));
  AOI21_X1   g32723(.A1(new_n35159_), .A2(new_n35158_), .B(pi0962), .ZN(po0880));
  NAND2_X1   g32724(.A1(new_n34723_), .A2(new_n16499_), .ZN(new_n35161_));
  NAND2_X1   g32725(.A1(po0980), .A2(pi1114), .ZN(new_n35162_));
  AOI21_X1   g32726(.A1(new_n35162_), .A2(new_n35161_), .B(pi0962), .ZN(po0881));
  NAND2_X1   g32727(.A1(new_n34723_), .A2(new_n16168_), .ZN(new_n35164_));
  NAND2_X1   g32728(.A1(po0980), .A2(pi1120), .ZN(new_n35165_));
  AOI21_X1   g32729(.A1(new_n35165_), .A2(new_n35164_), .B(pi0962), .ZN(po0882));
  NAND2_X1   g32730(.A1(po0980), .A2(pi1126), .ZN(new_n35167_));
  NAND2_X1   g32731(.A1(new_n34723_), .A2(pi0726), .ZN(new_n35168_));
  AOI21_X1   g32732(.A1(new_n35167_), .A2(new_n35168_), .B(pi0962), .ZN(po0883));
  NAND2_X1   g32733(.A1(po0980), .A2(pi1102), .ZN(new_n35170_));
  NAND2_X1   g32734(.A1(new_n34723_), .A2(pi0727), .ZN(new_n35171_));
  AOI21_X1   g32735(.A1(new_n35170_), .A2(new_n35171_), .B(pi0962), .ZN(po0884));
  INV_X1     g32736(.I(pi0728), .ZN(new_n35173_));
  NAND2_X1   g32737(.A1(new_n34723_), .A2(new_n35173_), .ZN(new_n35174_));
  NAND2_X1   g32738(.A1(po0980), .A2(pi1131), .ZN(new_n35175_));
  AOI21_X1   g32739(.A1(new_n35175_), .A2(new_n35174_), .B(pi0962), .ZN(po0885));
  NAND2_X1   g32740(.A1(po0980), .A2(pi1104), .ZN(new_n35177_));
  NAND2_X1   g32741(.A1(new_n34723_), .A2(pi0729), .ZN(new_n35178_));
  AOI21_X1   g32742(.A1(new_n35177_), .A2(new_n35178_), .B(pi0962), .ZN(po0886));
  NAND2_X1   g32743(.A1(po0980), .A2(pi1106), .ZN(new_n35180_));
  NAND2_X1   g32744(.A1(new_n34723_), .A2(pi0730), .ZN(new_n35181_));
  AOI21_X1   g32745(.A1(new_n35180_), .A2(new_n35181_), .B(pi0962), .ZN(po0887));
  NOR2_X1    g32746(.A1(new_n35110_), .A2(new_n35127_), .ZN(new_n35183_));
  NOR2_X1    g32747(.A1(new_n35086_), .A2(new_n35183_), .ZN(new_n35184_));
  NOR2_X1    g32748(.A1(new_n35099_), .A2(new_n35104_), .ZN(new_n35185_));
  NAND4_X1   g32749(.A1(new_n35126_), .A2(new_n35118_), .A3(new_n35184_), .A4(new_n35185_), .ZN(new_n35186_));
  AOI21_X1   g32750(.A1(new_n35186_), .A2(new_n35119_), .B(pi0731), .ZN(new_n35187_));
  INV_X1     g32751(.I(new_n35080_), .ZN(new_n35188_));
  INV_X1     g32752(.I(new_n35086_), .ZN(new_n35189_));
  NOR2_X1    g32753(.A1(new_n35108_), .A2(new_n35183_), .ZN(new_n35190_));
  NAND3_X1   g32754(.A1(new_n35190_), .A2(pi0795), .A3(new_n35189_), .ZN(new_n35191_));
  AOI21_X1   g32755(.A1(new_n35191_), .A2(pi0731), .B(new_n35188_), .ZN(new_n35192_));
  AOI21_X1   g32756(.A1(new_n35191_), .A2(new_n35121_), .B(new_n35082_), .ZN(new_n35193_));
  NOR3_X1    g32757(.A1(new_n35192_), .A2(new_n35193_), .A3(new_n35187_), .ZN(po0888));
  NAND2_X1   g32758(.A1(new_n34229_), .A2(new_n35145_), .ZN(new_n35195_));
  NAND2_X1   g32759(.A1(po0954), .A2(pi1128), .ZN(new_n35196_));
  AOI21_X1   g32760(.A1(new_n35195_), .A2(new_n35196_), .B(pi0962), .ZN(po0889));
  NOR2_X1    g32761(.A1(new_n12895_), .A2(new_n4888_), .ZN(new_n35198_));
  NOR2_X1    g32762(.A1(new_n12793_), .A2(pi1135), .ZN(new_n35199_));
  OAI21_X1   g32763(.A1(new_n35198_), .A2(new_n35199_), .B(new_n5045_), .ZN(new_n35200_));
  OAI21_X1   g32764(.A1(new_n35200_), .A2(new_n34498_), .B(new_n10920_), .ZN(new_n35201_));
  OAI21_X1   g32765(.A1(pi0838), .A2(pi1136), .B(pi1134), .ZN(new_n35202_));
  NOR2_X1    g32766(.A1(new_n16756_), .A2(new_n4888_), .ZN(new_n35203_));
  NOR2_X1    g32767(.A1(new_n34354_), .A2(new_n16757_), .ZN(new_n35204_));
  NOR4_X1    g32768(.A1(new_n35204_), .A2(new_n34876_), .A3(new_n35202_), .A4(new_n35203_), .ZN(new_n35205_));
  NOR2_X1    g32769(.A1(new_n35205_), .A2(new_n35201_), .ZN(new_n35206_));
  OAI22_X1   g32770(.A1(new_n7240_), .A2(new_n34579_), .B1(new_n34580_), .B2(new_n32794_), .ZN(new_n35207_));
  NAND2_X1   g32771(.A1(new_n35207_), .A2(new_n34368_), .ZN(new_n35208_));
  OAI22_X1   g32772(.A1(new_n35208_), .A2(pi0590), .B1(new_n32584_), .B2(new_n34882_), .ZN(new_n35209_));
  NAND2_X1   g32773(.A1(new_n35209_), .A2(new_n6251_), .ZN(new_n35210_));
  NAND2_X1   g32774(.A1(pi0199), .A2(pi1047), .ZN(new_n35211_));
  NOR2_X1    g32775(.A1(new_n8531_), .A2(new_n32493_), .ZN(new_n35212_));
  AOI21_X1   g32776(.A1(new_n8531_), .A2(pi0308), .B(new_n35212_), .ZN(new_n35213_));
  OAI21_X1   g32777(.A1(new_n35213_), .A2(pi0199), .B(new_n35211_), .ZN(new_n35214_));
  NAND2_X1   g32778(.A1(new_n34729_), .A2(pi0424), .ZN(new_n35215_));
  OAI21_X1   g32779(.A1(new_n35215_), .A2(new_n34891_), .B(new_n7253_), .ZN(new_n35216_));
  AOI21_X1   g32780(.A1(new_n35214_), .A2(new_n34369_), .B(new_n35216_), .ZN(new_n35217_));
  AOI21_X1   g32781(.A1(new_n35210_), .A2(new_n35217_), .B(new_n35206_), .ZN(po0890));
  NAND2_X1   g32782(.A1(new_n34723_), .A2(new_n16620_), .ZN(new_n35219_));
  NAND2_X1   g32783(.A1(po0980), .A2(pi1119), .ZN(new_n35220_));
  AOI21_X1   g32784(.A1(new_n35220_), .A2(new_n35219_), .B(pi0962), .ZN(po0891));
  NAND2_X1   g32785(.A1(po0980), .A2(pi1109), .ZN(new_n35222_));
  NAND2_X1   g32786(.A1(new_n34723_), .A2(pi0735), .ZN(new_n35223_));
  AOI21_X1   g32787(.A1(new_n35222_), .A2(new_n35223_), .B(pi0962), .ZN(po0892));
  NAND2_X1   g32788(.A1(po0980), .A2(pi1101), .ZN(new_n35225_));
  NAND2_X1   g32789(.A1(new_n34723_), .A2(pi0736), .ZN(new_n35226_));
  AOI21_X1   g32790(.A1(new_n35225_), .A2(new_n35226_), .B(pi0962), .ZN(po0893));
  NAND2_X1   g32791(.A1(new_n34723_), .A2(new_n16756_), .ZN(new_n35228_));
  NAND2_X1   g32792(.A1(po0980), .A2(pi1122), .ZN(new_n35229_));
  AOI21_X1   g32793(.A1(new_n35229_), .A2(new_n35228_), .B(pi0962), .ZN(po0894));
  NAND2_X1   g32794(.A1(new_n34723_), .A2(new_n12820_), .ZN(new_n35231_));
  NAND2_X1   g32795(.A1(po0980), .A2(pi1121), .ZN(new_n35232_));
  AOI21_X1   g32796(.A1(new_n35232_), .A2(new_n35231_), .B(pi0962), .ZN(po0895));
  INV_X1     g32797(.I(new_n34143_), .ZN(new_n35234_));
  OR2_X2     g32798(.A1(pi0952), .A2(pi1061), .Z(new_n35235_));
  NOR3_X1    g32799(.A1(new_n35234_), .A2(new_n12738_), .A3(new_n35235_), .ZN(po0988));
  INV_X1     g32800(.I(po0988), .ZN(new_n35237_));
  NOR2_X1    g32801(.A1(new_n35237_), .A2(pi1108), .ZN(new_n35238_));
  NOR2_X1    g32802(.A1(po0988), .A2(pi0739), .ZN(new_n35239_));
  OAI21_X1   g32803(.A1(new_n35238_), .A2(new_n35239_), .B(new_n34139_), .ZN(po0896));
  NOR2_X1    g32804(.A1(new_n35237_), .A2(pi1114), .ZN(new_n35241_));
  NOR2_X1    g32805(.A1(po0988), .A2(new_n16500_), .ZN(new_n35242_));
  OAI21_X1   g32806(.A1(new_n35241_), .A2(new_n35242_), .B(new_n34139_), .ZN(po0898));
  NOR2_X1    g32807(.A1(new_n35237_), .A2(pi1112), .ZN(new_n35244_));
  NOR2_X1    g32808(.A1(po0988), .A2(new_n16430_), .ZN(new_n35245_));
  OAI21_X1   g32809(.A1(new_n35244_), .A2(new_n35245_), .B(new_n34139_), .ZN(po0899));
  NOR2_X1    g32810(.A1(new_n35237_), .A2(pi1109), .ZN(new_n35247_));
  NOR2_X1    g32811(.A1(po0988), .A2(pi0743), .ZN(new_n35248_));
  OAI21_X1   g32812(.A1(new_n35247_), .A2(new_n35248_), .B(new_n34139_), .ZN(po0900));
  NOR2_X1    g32813(.A1(new_n35237_), .A2(pi1131), .ZN(new_n35250_));
  INV_X1     g32814(.I(pi0744), .ZN(new_n35251_));
  NOR2_X1    g32815(.A1(po0988), .A2(new_n35251_), .ZN(new_n35252_));
  OAI21_X1   g32816(.A1(new_n35250_), .A2(new_n35252_), .B(new_n34139_), .ZN(po0901));
  NOR2_X1    g32817(.A1(new_n35237_), .A2(pi1111), .ZN(new_n35254_));
  NOR2_X1    g32818(.A1(po0988), .A2(new_n16245_), .ZN(new_n35255_));
  OAI21_X1   g32819(.A1(new_n35254_), .A2(new_n35255_), .B(new_n34139_), .ZN(po0902));
  NOR2_X1    g32820(.A1(new_n35237_), .A2(pi1104), .ZN(new_n35257_));
  NOR2_X1    g32821(.A1(po0988), .A2(pi0746), .ZN(new_n35258_));
  OAI21_X1   g32822(.A1(new_n35257_), .A2(new_n35258_), .B(new_n34139_), .ZN(po0903));
  NAND2_X1   g32823(.A1(new_n35184_), .A2(new_n35115_), .ZN(new_n35260_));
  NOR3_X1    g32824(.A1(new_n35260_), .A2(new_n35088_), .A3(new_n35099_), .ZN(new_n35261_));
  NOR2_X1    g32825(.A1(new_n35080_), .A2(new_n35103_), .ZN(new_n35262_));
  OR3_X2     g32826(.A1(new_n35092_), .A2(new_n35106_), .A3(new_n35262_), .Z(new_n35263_));
  NAND2_X1   g32827(.A1(new_n35094_), .A2(pi0801), .ZN(new_n35264_));
  NAND2_X1   g32828(.A1(new_n35263_), .A2(new_n35264_), .ZN(new_n35265_));
  XOR2_X1    g32829(.A1(new_n35262_), .A2(new_n35089_), .Z(new_n35266_));
  AOI21_X1   g32830(.A1(new_n35265_), .A2(new_n35261_), .B(new_n35266_), .ZN(po0904));
  NOR2_X1    g32831(.A1(new_n35237_), .A2(pi1106), .ZN(new_n35268_));
  NOR2_X1    g32832(.A1(po0988), .A2(pi0748), .ZN(new_n35269_));
  OAI21_X1   g32833(.A1(new_n35268_), .A2(new_n35269_), .B(new_n34139_), .ZN(po0905));
  NOR2_X1    g32834(.A1(new_n35237_), .A2(pi1105), .ZN(new_n35271_));
  NOR2_X1    g32835(.A1(po0988), .A2(pi0749), .ZN(new_n35272_));
  OAI21_X1   g32836(.A1(new_n35271_), .A2(new_n35272_), .B(new_n34139_), .ZN(po0906));
  NOR2_X1    g32837(.A1(new_n35237_), .A2(pi1130), .ZN(new_n35274_));
  INV_X1     g32838(.I(pi0750), .ZN(new_n35275_));
  NOR2_X1    g32839(.A1(po0988), .A2(new_n35275_), .ZN(new_n35276_));
  OAI21_X1   g32840(.A1(new_n35274_), .A2(new_n35276_), .B(new_n34139_), .ZN(po0907));
  NOR2_X1    g32841(.A1(new_n35237_), .A2(pi1123), .ZN(new_n35278_));
  NOR2_X1    g32842(.A1(po0988), .A2(new_n16210_), .ZN(new_n35279_));
  OAI21_X1   g32843(.A1(new_n35278_), .A2(new_n35279_), .B(new_n34139_), .ZN(po0908));
  NOR2_X1    g32844(.A1(new_n35237_), .A2(pi1124), .ZN(new_n35281_));
  NOR2_X1    g32845(.A1(po0988), .A2(new_n16803_), .ZN(new_n35282_));
  OAI21_X1   g32846(.A1(new_n35281_), .A2(new_n35282_), .B(new_n34139_), .ZN(po0909));
  NOR2_X1    g32847(.A1(new_n35237_), .A2(pi1117), .ZN(new_n35284_));
  NOR2_X1    g32848(.A1(po0988), .A2(new_n16550_), .ZN(new_n35285_));
  OAI21_X1   g32849(.A1(new_n35284_), .A2(new_n35285_), .B(new_n34139_), .ZN(po0910));
  NOR2_X1    g32850(.A1(new_n35237_), .A2(pi1118), .ZN(new_n35287_));
  NOR2_X1    g32851(.A1(po0988), .A2(new_n16585_), .ZN(new_n35288_));
  OAI21_X1   g32852(.A1(new_n35287_), .A2(new_n35288_), .B(new_n34139_), .ZN(po0911));
  NOR2_X1    g32853(.A1(new_n35237_), .A2(pi1120), .ZN(new_n35290_));
  NOR2_X1    g32854(.A1(po0988), .A2(new_n16169_), .ZN(new_n35291_));
  OAI21_X1   g32855(.A1(new_n35290_), .A2(new_n35291_), .B(new_n34139_), .ZN(po0912));
  NOR2_X1    g32856(.A1(new_n35237_), .A2(pi1119), .ZN(new_n35293_));
  NOR2_X1    g32857(.A1(po0988), .A2(new_n16621_), .ZN(new_n35294_));
  OAI21_X1   g32858(.A1(new_n35293_), .A2(new_n35294_), .B(new_n34139_), .ZN(po0913));
  NOR2_X1    g32859(.A1(new_n35237_), .A2(pi1113), .ZN(new_n35296_));
  NOR2_X1    g32860(.A1(po0988), .A2(new_n16460_), .ZN(new_n35297_));
  OAI21_X1   g32861(.A1(new_n35296_), .A2(new_n35297_), .B(new_n34139_), .ZN(po0914));
  NOR2_X1    g32862(.A1(new_n35237_), .A2(pi1101), .ZN(new_n35299_));
  NOR2_X1    g32863(.A1(po0988), .A2(pi0758), .ZN(new_n35300_));
  OAI21_X1   g32864(.A1(new_n35299_), .A2(new_n35300_), .B(new_n34139_), .ZN(po0915));
  NOR4_X1    g32865(.A1(new_n35234_), .A2(new_n12738_), .A3(pi1100), .A4(new_n35235_), .ZN(new_n35302_));
  NOR2_X1    g32866(.A1(po0988), .A2(pi0759), .ZN(new_n35303_));
  OAI21_X1   g32867(.A1(new_n35303_), .A2(new_n35302_), .B(new_n34139_), .ZN(po0916));
  NOR2_X1    g32868(.A1(new_n35237_), .A2(pi1115), .ZN(new_n35305_));
  NOR2_X1    g32869(.A1(po0988), .A2(new_n16512_), .ZN(new_n35306_));
  OAI21_X1   g32870(.A1(new_n35305_), .A2(new_n35306_), .B(new_n34139_), .ZN(po0917));
  NOR2_X1    g32871(.A1(new_n35237_), .A2(pi1121), .ZN(new_n35308_));
  NOR2_X1    g32872(.A1(po0988), .A2(new_n12750_), .ZN(new_n35309_));
  OAI21_X1   g32873(.A1(new_n35308_), .A2(new_n35309_), .B(new_n34139_), .ZN(po0918));
  NOR2_X1    g32874(.A1(new_n35237_), .A2(pi1129), .ZN(new_n35311_));
  INV_X1     g32875(.I(pi0762), .ZN(new_n35312_));
  NOR2_X1    g32876(.A1(po0988), .A2(new_n35312_), .ZN(new_n35313_));
  OAI21_X1   g32877(.A1(new_n35311_), .A2(new_n35313_), .B(new_n34139_), .ZN(po0919));
  NOR2_X1    g32878(.A1(new_n35237_), .A2(pi1103), .ZN(new_n35315_));
  NOR2_X1    g32879(.A1(po0988), .A2(pi0763), .ZN(new_n35316_));
  OAI21_X1   g32880(.A1(new_n35315_), .A2(new_n35316_), .B(new_n34139_), .ZN(po0920));
  NOR2_X1    g32881(.A1(new_n35237_), .A2(pi1107), .ZN(new_n35318_));
  NOR2_X1    g32882(.A1(po0988), .A2(pi0764), .ZN(new_n35319_));
  OAI21_X1   g32883(.A1(new_n35318_), .A2(new_n35319_), .B(new_n34139_), .ZN(po0921));
  INV_X1     g32884(.I(pi0765), .ZN(new_n35321_));
  INV_X1     g32885(.I(new_n35083_), .ZN(new_n35322_));
  NOR2_X1    g32886(.A1(new_n35101_), .A2(new_n35088_), .ZN(new_n35323_));
  INV_X1     g32887(.I(pi0771), .ZN(new_n35324_));
  NOR2_X1    g32888(.A1(new_n35324_), .A2(new_n35002_), .ZN(new_n35325_));
  NOR4_X1    g32889(.A1(new_n35093_), .A2(pi0765), .A3(new_n35098_), .A4(new_n35325_), .ZN(new_n35326_));
  NOR3_X1    g32890(.A1(new_n35326_), .A2(pi0773), .A3(pi0801), .ZN(new_n35327_));
  OAI21_X1   g32891(.A1(new_n35105_), .A2(new_n35327_), .B(new_n35323_), .ZN(new_n35328_));
  AOI21_X1   g32892(.A1(new_n35328_), .A2(new_n35109_), .B(new_n35322_), .ZN(new_n35329_));
  OAI21_X1   g32893(.A1(new_n35112_), .A2(new_n35127_), .B(new_n35329_), .ZN(new_n35330_));
  INV_X1     g32894(.I(new_n35190_), .ZN(new_n35331_));
  NOR3_X1    g32895(.A1(new_n35331_), .A2(new_n35084_), .A3(new_n34972_), .ZN(new_n35332_));
  NOR2_X1    g32896(.A1(new_n35332_), .A2(pi0765), .ZN(new_n35333_));
  AOI21_X1   g32897(.A1(new_n35333_), .A2(new_n35330_), .B(pi0795), .ZN(new_n35334_));
  NOR2_X1    g32898(.A1(new_n35334_), .A2(pi0731), .ZN(new_n35335_));
  NAND2_X1   g32899(.A1(new_n35191_), .A2(pi0731), .ZN(new_n35336_));
  OAI21_X1   g32900(.A1(new_n35334_), .A2(pi0731), .B(new_n35336_), .ZN(new_n35337_));
  AOI22_X1   g32901(.A1(new_n35337_), .A2(new_n35321_), .B1(new_n35335_), .B2(new_n35118_), .ZN(new_n35338_));
  NOR2_X1    g32902(.A1(new_n35108_), .A2(new_n35260_), .ZN(po0978));
  NAND2_X1   g32903(.A1(pi0765), .A2(pi0945), .ZN(new_n35340_));
  OAI22_X1   g32904(.A1(new_n35338_), .A2(pi0945), .B1(po0978), .B2(new_n35340_), .ZN(po0922));
  NOR2_X1    g32905(.A1(new_n35237_), .A2(pi1110), .ZN(new_n35342_));
  NOR2_X1    g32906(.A1(po0988), .A2(pi0766), .ZN(new_n35343_));
  OAI21_X1   g32907(.A1(new_n35342_), .A2(new_n35343_), .B(new_n34139_), .ZN(po0923));
  NOR2_X1    g32908(.A1(new_n35237_), .A2(pi1116), .ZN(new_n35345_));
  NOR2_X1    g32909(.A1(po0988), .A2(new_n15782_), .ZN(new_n35346_));
  OAI21_X1   g32910(.A1(new_n35345_), .A2(new_n35346_), .B(new_n34139_), .ZN(po0924));
  NOR2_X1    g32911(.A1(new_n35237_), .A2(pi1125), .ZN(new_n35348_));
  NOR2_X1    g32912(.A1(po0988), .A2(new_n16912_), .ZN(new_n35349_));
  OAI21_X1   g32913(.A1(new_n35348_), .A2(new_n35349_), .B(new_n34139_), .ZN(po0925));
  NOR4_X1    g32914(.A1(new_n35095_), .A2(new_n35072_), .A3(new_n35088_), .A4(new_n35106_), .ZN(new_n35351_));
  AND2_X2    g32915(.A1(new_n35351_), .A2(new_n35184_), .Z(new_n35352_));
  NAND2_X1   g32916(.A1(new_n35352_), .A2(new_n35115_), .ZN(new_n35353_));
  NAND2_X1   g32917(.A1(new_n35353_), .A2(pi0769), .ZN(new_n35354_));
  AOI21_X1   g32918(.A1(new_n35119_), .A2(pi0775), .B(new_n35097_), .ZN(new_n35355_));
  NOR3_X1    g32919(.A1(new_n35121_), .A2(pi0769), .A3(new_n35084_), .ZN(new_n35356_));
  OAI21_X1   g32920(.A1(new_n35356_), .A2(new_n35355_), .B(new_n35081_), .ZN(new_n35357_));
  AOI21_X1   g32921(.A1(new_n35084_), .A2(new_n35352_), .B(new_n35332_), .ZN(new_n35358_));
  NOR2_X1    g32922(.A1(new_n35358_), .A2(new_n35118_), .ZN(new_n35359_));
  OAI22_X1   g32923(.A1(new_n35359_), .A2(new_n35357_), .B1(new_n35081_), .B2(new_n35354_), .ZN(po0926));
  NOR2_X1    g32924(.A1(new_n35237_), .A2(pi1126), .ZN(new_n35361_));
  NOR2_X1    g32925(.A1(po0988), .A2(new_n16080_), .ZN(new_n35362_));
  OAI21_X1   g32926(.A1(new_n35361_), .A2(new_n35362_), .B(new_n34139_), .ZN(po0927));
  INV_X1     g32927(.I(po0978), .ZN(new_n35364_));
  NAND2_X1   g32928(.A1(new_n35364_), .A2(pi0771), .ZN(new_n35365_));
  INV_X1     g32929(.I(new_n35115_), .ZN(new_n35366_));
  NOR3_X1    g32930(.A1(new_n35329_), .A2(pi0731), .A3(new_n35085_), .ZN(new_n35367_));
  NOR2_X1    g32931(.A1(new_n35189_), .A2(new_n35078_), .ZN(new_n35368_));
  NOR4_X1    g32932(.A1(new_n35367_), .A2(new_n35366_), .A3(new_n35331_), .A4(new_n35368_), .ZN(po0963));
  NAND2_X1   g32933(.A1(new_n35079_), .A2(pi0987), .ZN(new_n35370_));
  OAI22_X1   g32934(.A1(po0963), .A2(new_n35370_), .B1(new_n35079_), .B2(new_n35365_), .ZN(po0928));
  NOR2_X1    g32935(.A1(new_n35237_), .A2(pi1102), .ZN(new_n35372_));
  NOR2_X1    g32936(.A1(po0988), .A2(pi0772), .ZN(new_n35373_));
  OAI21_X1   g32937(.A1(new_n35372_), .A2(new_n35373_), .B(new_n34139_), .ZN(po0929));
  NAND3_X1   g32938(.A1(po0963), .A2(new_n35104_), .A3(new_n35323_), .ZN(new_n35375_));
  NAND2_X1   g32939(.A1(new_n35375_), .A2(new_n35188_), .ZN(new_n35376_));
  AOI21_X1   g32940(.A1(new_n35184_), .A2(new_n35115_), .B(new_n35104_), .ZN(new_n35377_));
  OAI21_X1   g32941(.A1(new_n35108_), .A2(new_n35377_), .B(pi0773), .ZN(new_n35378_));
  AOI21_X1   g32942(.A1(new_n35376_), .A2(new_n35378_), .B(new_n35262_), .ZN(po0930));
  NOR2_X1    g32943(.A1(new_n35237_), .A2(pi1127), .ZN(new_n35380_));
  NOR2_X1    g32944(.A1(po0988), .A2(new_n14851_), .ZN(new_n35381_));
  OAI21_X1   g32945(.A1(new_n35380_), .A2(new_n35381_), .B(new_n34139_), .ZN(po0931));
  NOR2_X1    g32946(.A1(new_n35078_), .A2(pi0945), .ZN(new_n35383_));
  NOR3_X1    g32947(.A1(new_n35121_), .A2(new_n35321_), .A3(new_n35324_), .ZN(new_n35384_));
  INV_X1     g32948(.I(new_n35384_), .ZN(new_n35385_));
  AOI21_X1   g32949(.A1(new_n35191_), .A2(new_n35385_), .B(new_n35084_), .ZN(new_n35386_));
  NOR4_X1    g32950(.A1(new_n35118_), .A2(new_n35002_), .A3(new_n35104_), .A4(pi0816), .ZN(new_n35387_));
  OAI21_X1   g32951(.A1(new_n35110_), .A2(new_n35127_), .B(new_n35387_), .ZN(new_n35388_));
  OAI21_X1   g32952(.A1(new_n35101_), .A2(new_n35388_), .B(new_n35384_), .ZN(new_n35389_));
  NAND2_X1   g32953(.A1(new_n35389_), .A2(new_n35084_), .ZN(new_n35390_));
  AOI22_X1   g32954(.A1(new_n35364_), .A2(pi0775), .B1(new_n35383_), .B2(new_n35390_), .ZN(new_n35391_));
  AOI21_X1   g32955(.A1(new_n35386_), .A2(new_n35383_), .B(new_n35391_), .ZN(po0932));
  NOR2_X1    g32956(.A1(new_n35237_), .A2(pi1128), .ZN(new_n35393_));
  INV_X1     g32957(.I(pi0776), .ZN(new_n35394_));
  NOR2_X1    g32958(.A1(po0988), .A2(new_n35394_), .ZN(new_n35395_));
  OAI21_X1   g32959(.A1(new_n35393_), .A2(new_n35395_), .B(new_n34139_), .ZN(po0933));
  NOR2_X1    g32960(.A1(new_n35237_), .A2(pi1122), .ZN(new_n35397_));
  NOR2_X1    g32961(.A1(po0988), .A2(new_n16757_), .ZN(new_n35398_));
  OAI21_X1   g32962(.A1(new_n35397_), .A2(new_n35398_), .B(new_n34139_), .ZN(po0934));
  NOR2_X1    g32963(.A1(pi1046), .A2(pi1083), .ZN(new_n35400_));
  NAND4_X1   g32964(.A1(new_n35400_), .A2(pi0832), .A3(pi0956), .A4(pi1085), .ZN(new_n35401_));
  NOR2_X1    g32965(.A1(new_n35401_), .A2(pi0968), .ZN(new_n35402_));
  NAND2_X1   g32966(.A1(new_n35402_), .A2(pi1100), .ZN(new_n35403_));
  OAI21_X1   g32967(.A1(new_n12758_), .A2(new_n35402_), .B(new_n35403_), .ZN(po0935));
  OAI21_X1   g32968(.A1(new_n34119_), .A2(new_n5473_), .B(pi0779), .ZN(po0936));
  OAI21_X1   g32969(.A1(new_n34119_), .A2(new_n5692_), .B(pi0780), .ZN(po0937));
  NAND2_X1   g32970(.A1(new_n35402_), .A2(pi1101), .ZN(new_n35407_));
  OAI21_X1   g32971(.A1(new_n12779_), .A2(new_n35402_), .B(new_n35407_), .ZN(po0938));
  NAND3_X1   g32972(.A1(new_n34119_), .A2(new_n33010_), .A3(new_n34153_), .ZN(po0939));
  NAND2_X1   g32973(.A1(new_n35402_), .A2(pi1109), .ZN(new_n35410_));
  OAI21_X1   g32974(.A1(new_n34585_), .A2(new_n35402_), .B(new_n35410_), .ZN(po0940));
  NAND2_X1   g32975(.A1(new_n35402_), .A2(pi1110), .ZN(new_n35412_));
  OAI21_X1   g32976(.A1(new_n34360_), .A2(new_n35402_), .B(new_n35412_), .ZN(po0941));
  NAND2_X1   g32977(.A1(new_n35402_), .A2(pi1102), .ZN(new_n35414_));
  OAI21_X1   g32978(.A1(new_n12764_), .A2(new_n35402_), .B(new_n35414_), .ZN(po0942));
  NAND2_X1   g32979(.A1(new_n8297_), .A2(pi0954), .ZN(new_n35416_));
  OAI21_X1   g32980(.A1(pi0024), .A2(pi0954), .B(new_n35416_), .ZN(po0943));
  NAND2_X1   g32981(.A1(new_n35402_), .A2(pi1104), .ZN(new_n35418_));
  OAI21_X1   g32982(.A1(new_n12972_), .A2(new_n35402_), .B(new_n35418_), .ZN(po0944));
  NAND2_X1   g32983(.A1(new_n35402_), .A2(pi1105), .ZN(new_n35420_));
  OAI21_X1   g32984(.A1(new_n12808_), .A2(new_n35402_), .B(new_n35420_), .ZN(po0945));
  NAND2_X1   g32985(.A1(new_n35402_), .A2(pi1106), .ZN(new_n35422_));
  OAI21_X1   g32986(.A1(new_n12796_), .A2(new_n35402_), .B(new_n35422_), .ZN(po0946));
  NAND2_X1   g32987(.A1(new_n35402_), .A2(pi1107), .ZN(new_n35424_));
  OAI21_X1   g32988(.A1(new_n13000_), .A2(new_n35402_), .B(new_n35424_), .ZN(po0947));
  NAND2_X1   g32989(.A1(new_n35402_), .A2(pi1108), .ZN(new_n35426_));
  OAI21_X1   g32990(.A1(new_n34681_), .A2(new_n35402_), .B(new_n35426_), .ZN(po0948));
  NAND2_X1   g32991(.A1(new_n35402_), .A2(pi1103), .ZN(new_n35428_));
  OAI21_X1   g32992(.A1(new_n12937_), .A2(new_n35402_), .B(new_n35428_), .ZN(po0949));
  INV_X1     g32993(.I(pi0968), .ZN(new_n35430_));
  NOR2_X1    g32994(.A1(new_n35401_), .A2(new_n35430_), .ZN(new_n35431_));
  NAND2_X1   g32995(.A1(new_n35431_), .A2(pi1130), .ZN(new_n35432_));
  OAI21_X1   g32996(.A1(new_n35072_), .A2(new_n35431_), .B(new_n35432_), .ZN(po0951));
  NAND2_X1   g32997(.A1(new_n35431_), .A2(pi1128), .ZN(new_n35434_));
  OAI21_X1   g32998(.A1(new_n35118_), .A2(new_n35431_), .B(new_n35434_), .ZN(po0952));
  INV_X1     g32999(.I(pi0278), .ZN(po1130));
  NAND2_X1   g33000(.A1(new_n32317_), .A2(pi0279), .ZN(new_n35437_));
  NOR4_X1    g33001(.A1(new_n35437_), .A2(new_n4727_), .A3(pi0269), .A4(po1130), .ZN(new_n35438_));
  NAND3_X1   g33002(.A1(new_n35438_), .A2(new_n4278_), .A3(new_n34333_), .ZN(new_n35439_));
  XOR2_X1    g33003(.A1(new_n35439_), .A2(pi0264), .Z(po0953));
  INV_X1     g33004(.I(pi0798), .ZN(new_n35441_));
  NAND2_X1   g33005(.A1(new_n35431_), .A2(pi1124), .ZN(new_n35442_));
  OAI21_X1   g33006(.A1(new_n35441_), .A2(new_n35431_), .B(new_n35442_), .ZN(po0955));
  NAND2_X1   g33007(.A1(new_n35431_), .A2(pi1107), .ZN(new_n35444_));
  OAI21_X1   g33008(.A1(pi0799), .A2(new_n35431_), .B(new_n35444_), .ZN(po0956));
  NAND2_X1   g33009(.A1(new_n35431_), .A2(pi1125), .ZN(new_n35446_));
  OAI21_X1   g33010(.A1(new_n35002_), .A2(new_n35431_), .B(new_n35446_), .ZN(po0957));
  NAND2_X1   g33011(.A1(new_n35431_), .A2(pi1126), .ZN(new_n35448_));
  OAI21_X1   g33012(.A1(new_n35104_), .A2(new_n35431_), .B(new_n35448_), .ZN(po0958));
  NOR3_X1    g33013(.A1(new_n34334_), .A2(pi0265), .A3(pi0274), .ZN(po0959));
  NAND2_X1   g33014(.A1(new_n35431_), .A2(pi1106), .ZN(new_n35451_));
  OAI21_X1   g33015(.A1(pi0803), .A2(new_n35431_), .B(new_n35451_), .ZN(po0960));
  NAND2_X1   g33016(.A1(new_n35431_), .A2(pi1109), .ZN(new_n35453_));
  OAI21_X1   g33017(.A1(new_n32939_), .A2(new_n35431_), .B(new_n35453_), .ZN(po0961));
  NAND2_X1   g33018(.A1(new_n34332_), .A2(new_n32379_), .ZN(new_n35455_));
  XOR2_X1    g33019(.A1(new_n35455_), .A2(pi0270), .Z(po0962));
  NAND2_X1   g33020(.A1(new_n35431_), .A2(pi1127), .ZN(new_n35457_));
  OAI21_X1   g33021(.A1(new_n35041_), .A2(new_n35431_), .B(new_n35457_), .ZN(po0964));
  NAND2_X1   g33022(.A1(new_n35431_), .A2(pi1101), .ZN(new_n35459_));
  OAI21_X1   g33023(.A1(new_n34535_), .A2(new_n35431_), .B(new_n35459_), .ZN(po0965));
  NAND2_X1   g33024(.A1(new_n35431_), .A2(pi1103), .ZN(new_n35461_));
  OAI21_X1   g33025(.A1(pi0809), .A2(new_n35431_), .B(new_n35461_), .ZN(po0966));
  NAND2_X1   g33026(.A1(new_n35431_), .A2(pi1108), .ZN(new_n35463_));
  OAI21_X1   g33027(.A1(new_n32940_), .A2(new_n35431_), .B(new_n35463_), .ZN(po0967));
  NAND2_X1   g33028(.A1(new_n35431_), .A2(pi1102), .ZN(new_n35465_));
  OAI21_X1   g33029(.A1(new_n34402_), .A2(new_n35431_), .B(new_n35465_), .ZN(po0968));
  NAND2_X1   g33030(.A1(new_n35431_), .A2(pi1104), .ZN(new_n35467_));
  OAI21_X1   g33031(.A1(pi0812), .A2(new_n35431_), .B(new_n35467_), .ZN(po0969));
  NAND2_X1   g33032(.A1(new_n35431_), .A2(pi1131), .ZN(new_n35469_));
  OAI21_X1   g33033(.A1(new_n34746_), .A2(new_n35431_), .B(new_n35469_), .ZN(po0970));
  NAND2_X1   g33034(.A1(new_n35431_), .A2(pi1105), .ZN(new_n35471_));
  OAI21_X1   g33035(.A1(pi0814), .A2(new_n35431_), .B(new_n35471_), .ZN(po0971));
  NAND2_X1   g33036(.A1(new_n35431_), .A2(pi1110), .ZN(new_n35473_));
  OAI21_X1   g33037(.A1(new_n32938_), .A2(new_n35431_), .B(new_n35473_), .ZN(po0972));
  NAND2_X1   g33038(.A1(new_n35431_), .A2(pi1129), .ZN(new_n35475_));
  OAI21_X1   g33039(.A1(new_n34972_), .A2(new_n35431_), .B(new_n35475_), .ZN(po0973));
  XOR2_X1    g33040(.A1(new_n34331_), .A2(pi0269), .Z(po0974));
  OAI21_X1   g33041(.A1(new_n11010_), .A2(new_n10920_), .B(new_n10901_), .ZN(po0975));
  XOR2_X1    g33042(.A1(new_n34334_), .A2(pi0265), .Z(po0976));
  NOR2_X1    g33043(.A1(new_n35455_), .A2(pi0270), .ZN(new_n35480_));
  XOR2_X1    g33044(.A1(new_n35480_), .A2(new_n32211_), .Z(po0977));
  NOR2_X1    g33045(.A1(pi0811), .A2(pi0893), .ZN(po0979));
  OAI22_X1   g33046(.A1(new_n8218_), .A2(pi0982), .B1(new_n6871_), .B2(new_n10920_), .ZN(new_n35483_));
  AND2_X2    g33047(.A1(new_n35483_), .A2(new_n8913_), .Z(po0981));
  INV_X1     g33048(.I(pi0825), .ZN(po1147));
  NOR2_X1    g33049(.A1(new_n2644_), .A2(new_n31383_), .ZN(new_n35486_));
  INV_X1     g33050(.I(new_n35486_), .ZN(new_n35487_));
  OR3_X2     g33051(.A1(new_n35486_), .A2(pi1127), .A3(pi1131), .Z(new_n35488_));
  OAI21_X1   g33052(.A1(po1147), .A2(new_n35487_), .B(new_n35488_), .ZN(new_n35489_));
  XNOR2_X1   g33053(.A1(pi1124), .A2(pi1130), .ZN(new_n35490_));
  XOR2_X1    g33054(.A1(pi1125), .A2(pi1129), .Z(new_n35491_));
  XOR2_X1    g33055(.A1(pi1126), .A2(pi1128), .Z(new_n35492_));
  XNOR2_X1   g33056(.A1(new_n35491_), .A2(new_n35492_), .ZN(new_n35493_));
  XOR2_X1    g33057(.A1(new_n35493_), .A2(new_n35490_), .Z(new_n35494_));
  INV_X1     g33058(.I(new_n35494_), .ZN(new_n35495_));
  NAND3_X1   g33059(.A1(new_n35487_), .A2(pi1127), .A3(pi1131), .ZN(new_n35496_));
  NAND2_X1   g33060(.A1(new_n35495_), .A2(new_n35496_), .ZN(new_n35497_));
  NAND2_X1   g33061(.A1(new_n35486_), .A2(po1147), .ZN(new_n35498_));
  AND3_X2    g33062(.A1(new_n35496_), .A2(new_n35488_), .A3(new_n35498_), .Z(new_n35499_));
  OAI22_X1   g33063(.A1(new_n35497_), .A2(new_n35489_), .B1(new_n35495_), .B2(new_n35499_), .ZN(po0982));
  INV_X1     g33064(.I(pi0826), .ZN(po1148));
  OR3_X2     g33065(.A1(new_n35486_), .A2(pi1122), .A3(pi1123), .Z(new_n35502_));
  OAI21_X1   g33066(.A1(po1148), .A2(new_n35487_), .B(new_n35502_), .ZN(new_n35503_));
  XNOR2_X1   g33067(.A1(pi1118), .A2(pi1119), .ZN(new_n35504_));
  XOR2_X1    g33068(.A1(pi1116), .A2(pi1121), .Z(new_n35505_));
  XOR2_X1    g33069(.A1(pi1117), .A2(pi1120), .Z(new_n35506_));
  XNOR2_X1   g33070(.A1(new_n35505_), .A2(new_n35506_), .ZN(new_n35507_));
  XOR2_X1    g33071(.A1(new_n35507_), .A2(new_n35504_), .Z(new_n35508_));
  INV_X1     g33072(.I(new_n35508_), .ZN(new_n35509_));
  NAND3_X1   g33073(.A1(new_n35487_), .A2(pi1122), .A3(pi1123), .ZN(new_n35510_));
  NAND2_X1   g33074(.A1(new_n35509_), .A2(new_n35510_), .ZN(new_n35511_));
  NAND2_X1   g33075(.A1(new_n35486_), .A2(po1148), .ZN(new_n35512_));
  AND3_X2    g33076(.A1(new_n35510_), .A2(new_n35502_), .A3(new_n35512_), .Z(new_n35513_));
  OAI22_X1   g33077(.A1(new_n35511_), .A2(new_n35503_), .B1(new_n35509_), .B2(new_n35513_), .ZN(po0983));
  INV_X1     g33078(.I(pi0827), .ZN(po1178));
  OR3_X2     g33079(.A1(new_n35486_), .A2(pi1100), .A3(pi1107), .Z(new_n35516_));
  OAI21_X1   g33080(.A1(po1178), .A2(new_n35487_), .B(new_n35516_), .ZN(new_n35517_));
  XNOR2_X1   g33081(.A1(pi1103), .A2(pi1105), .ZN(new_n35518_));
  XOR2_X1    g33082(.A1(pi1101), .A2(pi1106), .Z(new_n35519_));
  XOR2_X1    g33083(.A1(pi1102), .A2(pi1104), .Z(new_n35520_));
  XNOR2_X1   g33084(.A1(new_n35519_), .A2(new_n35520_), .ZN(new_n35521_));
  XOR2_X1    g33085(.A1(new_n35521_), .A2(new_n35518_), .Z(new_n35522_));
  INV_X1     g33086(.I(new_n35522_), .ZN(new_n35523_));
  NAND3_X1   g33087(.A1(new_n35487_), .A2(pi1100), .A3(pi1107), .ZN(new_n35524_));
  NAND2_X1   g33088(.A1(new_n35523_), .A2(new_n35524_), .ZN(new_n35525_));
  NAND2_X1   g33089(.A1(new_n35486_), .A2(po1178), .ZN(new_n35526_));
  AND3_X2    g33090(.A1(new_n35524_), .A2(new_n35516_), .A3(new_n35526_), .Z(new_n35527_));
  OAI22_X1   g33091(.A1(new_n35525_), .A2(new_n35517_), .B1(new_n35523_), .B2(new_n35527_), .ZN(po0984));
  INV_X1     g33092(.I(pi0828), .ZN(po1182));
  OR3_X2     g33093(.A1(new_n35486_), .A2(pi1114), .A3(pi1115), .Z(new_n35530_));
  OAI21_X1   g33094(.A1(po1182), .A2(new_n35487_), .B(new_n35530_), .ZN(new_n35531_));
  XNOR2_X1   g33095(.A1(pi1110), .A2(pi1111), .ZN(new_n35532_));
  XOR2_X1    g33096(.A1(pi1108), .A2(pi1113), .Z(new_n35533_));
  XOR2_X1    g33097(.A1(pi1109), .A2(pi1112), .Z(new_n35534_));
  XNOR2_X1   g33098(.A1(new_n35533_), .A2(new_n35534_), .ZN(new_n35535_));
  XOR2_X1    g33099(.A1(new_n35535_), .A2(new_n35532_), .Z(new_n35536_));
  INV_X1     g33100(.I(new_n35536_), .ZN(new_n35537_));
  NAND3_X1   g33101(.A1(new_n35487_), .A2(pi1114), .A3(pi1115), .ZN(new_n35538_));
  NAND2_X1   g33102(.A1(new_n35537_), .A2(new_n35538_), .ZN(new_n35539_));
  NAND2_X1   g33103(.A1(new_n35486_), .A2(po1182), .ZN(new_n35540_));
  AND3_X2    g33104(.A1(new_n35538_), .A2(new_n35530_), .A3(new_n35540_), .Z(new_n35541_));
  OAI22_X1   g33105(.A1(new_n35539_), .A2(new_n35531_), .B1(new_n35537_), .B2(new_n35541_), .ZN(po0985));
  NAND2_X1   g33106(.A1(new_n3080_), .A2(new_n7253_), .ZN(new_n35543_));
  AOI21_X1   g33107(.A1(new_n35543_), .A2(pi0951), .B(new_n3040_), .ZN(po0986));
  XOR2_X1    g33108(.A1(new_n35438_), .A2(new_n4278_), .Z(po0987));
  NOR3_X1    g33109(.A1(new_n7261_), .A2(pi0832), .A3(new_n3022_), .ZN(po0989));
  OAI21_X1   g33110(.A1(new_n2443_), .A2(new_n3042_), .B(new_n6747_), .ZN(po0990));
  AND2_X2    g33111(.A1(new_n3042_), .A2(pi0946), .Z(po0991));
  XOR2_X1    g33112(.A1(new_n34332_), .A2(new_n32379_), .Z(po0992));
  NAND2_X1   g33113(.A1(pi0837), .A2(pi0955), .ZN(new_n35550_));
  OAI21_X1   g33114(.A1(pi0955), .A2(new_n32478_), .B(new_n35550_), .ZN(po0993));
  MUX2_X1    g33115(.I0(pi1047), .I1(pi0838), .S(pi0955), .Z(po0994));
  NAND2_X1   g33116(.A1(pi0839), .A2(pi0955), .ZN(new_n35553_));
  OAI21_X1   g33117(.A1(pi0955), .A2(new_n32590_), .B(new_n35553_), .ZN(po0995));
  NAND2_X1   g33118(.A1(new_n3043_), .A2(pi0840), .ZN(new_n35555_));
  OAI21_X1   g33119(.A1(new_n6302_), .A2(new_n3043_), .B(new_n35555_), .ZN(po0996));
  NOR2_X1    g33120(.A1(new_n7564_), .A2(pi0033), .ZN(po0997));
  MUX2_X1    g33121(.I0(pi1035), .I1(pi0842), .S(pi0955), .Z(po0998));
  NAND2_X1   g33122(.A1(pi0843), .A2(pi0955), .ZN(new_n35559_));
  OAI21_X1   g33123(.A1(pi0955), .A2(new_n32740_), .B(new_n35559_), .ZN(po0999));
  NAND2_X1   g33124(.A1(pi0844), .A2(pi0955), .ZN(new_n35561_));
  OAI21_X1   g33125(.A1(pi0955), .A2(new_n32685_), .B(new_n35561_), .ZN(po1000));
  MUX2_X1    g33126(.I0(pi1043), .I1(pi0845), .S(pi0955), .Z(po1001));
  NAND2_X1   g33127(.A1(new_n31388_), .A2(pi0846), .ZN(new_n35564_));
  OAI21_X1   g33128(.A1(new_n5045_), .A2(new_n31388_), .B(new_n35564_), .ZN(po1002));
  NAND2_X1   g33129(.A1(pi0847), .A2(pi0955), .ZN(new_n35566_));
  OAI21_X1   g33130(.A1(pi0955), .A2(new_n32672_), .B(new_n35566_), .ZN(po1003));
  MUX2_X1    g33131(.I0(pi1039), .I1(pi0848), .S(pi0955), .Z(po1004));
  NAND2_X1   g33132(.A1(new_n3043_), .A2(pi0849), .ZN(new_n35569_));
  OAI21_X1   g33133(.A1(new_n6274_), .A2(new_n3043_), .B(new_n35569_), .ZN(po1005));
  NAND2_X1   g33134(.A1(pi0850), .A2(pi0955), .ZN(new_n35571_));
  OAI21_X1   g33135(.A1(pi0955), .A2(new_n32475_), .B(new_n35571_), .ZN(po1006));
  NAND2_X1   g33136(.A1(pi0851), .A2(pi0955), .ZN(new_n35573_));
  OAI21_X1   g33137(.A1(pi0955), .A2(new_n35134_), .B(new_n35573_), .ZN(po1007));
  NAND2_X1   g33138(.A1(pi0852), .A2(pi0955), .ZN(new_n35575_));
  OAI21_X1   g33139(.A1(pi0955), .A2(new_n31356_), .B(new_n35575_), .ZN(po1008));
  MUX2_X1    g33140(.I0(pi1080), .I1(pi0853), .S(pi0955), .Z(po1009));
  NAND2_X1   g33141(.A1(pi0854), .A2(pi0955), .ZN(new_n35578_));
  OAI21_X1   g33142(.A1(pi0955), .A2(new_n34939_), .B(new_n35578_), .ZN(po1010));
  NAND2_X1   g33143(.A1(pi0855), .A2(pi0955), .ZN(new_n35580_));
  OAI21_X1   g33144(.A1(pi0955), .A2(new_n31350_), .B(new_n35580_), .ZN(po1011));
  NAND2_X1   g33145(.A1(pi0856), .A2(pi0955), .ZN(new_n35582_));
  OAI21_X1   g33146(.A1(pi0955), .A2(new_n32722_), .B(new_n35582_), .ZN(po1012));
  MUX2_X1    g33147(.I0(pi1058), .I1(pi0857), .S(pi0955), .Z(po1013));
  NAND2_X1   g33148(.A1(pi0858), .A2(pi0955), .ZN(new_n35585_));
  OAI21_X1   g33149(.A1(pi0955), .A2(new_n32675_), .B(new_n35585_), .ZN(po1014));
  NAND2_X1   g33150(.A1(pi0859), .A2(pi0955), .ZN(new_n35587_));
  OAI21_X1   g33151(.A1(pi0955), .A2(new_n31344_), .B(new_n35587_), .ZN(po1015));
  NAND2_X1   g33152(.A1(pi0860), .A2(pi0955), .ZN(new_n35589_));
  OAI21_X1   g33153(.A1(pi0955), .A2(new_n32697_), .B(new_n35589_), .ZN(po1016));
  NOR2_X1    g33154(.A1(new_n3041_), .A2(new_n3926_), .ZN(new_n35591_));
  NOR2_X1    g33155(.A1(new_n3934_), .A2(pi1093), .ZN(new_n35592_));
  OAI21_X1   g33156(.A1(new_n35591_), .A2(new_n35592_), .B(new_n2458_), .ZN(new_n35593_));
  NOR2_X1    g33157(.A1(new_n31383_), .A2(new_n3934_), .ZN(new_n35594_));
  NOR2_X1    g33158(.A1(new_n3926_), .A2(pi0123), .ZN(new_n35595_));
  OAI21_X1   g33159(.A1(new_n35594_), .A2(new_n35595_), .B(pi0228), .ZN(new_n35596_));
  NAND2_X1   g33160(.A1(new_n35593_), .A2(new_n35596_), .ZN(po1017));
  NAND2_X1   g33161(.A1(new_n31388_), .A2(pi0862), .ZN(new_n35598_));
  OAI21_X1   g33162(.A1(new_n4238_), .A2(new_n31388_), .B(new_n35598_), .ZN(po1018));
  NAND2_X1   g33163(.A1(new_n3043_), .A2(pi0863), .ZN(new_n35600_));
  OAI21_X1   g33164(.A1(new_n6380_), .A2(new_n3043_), .B(new_n35600_), .ZN(po1019));
  NAND2_X1   g33165(.A1(new_n3043_), .A2(pi0864), .ZN(new_n35602_));
  OAI21_X1   g33166(.A1(new_n6273_), .A2(new_n3043_), .B(new_n35602_), .ZN(po1020));
  NAND2_X1   g33167(.A1(pi0865), .A2(pi0955), .ZN(new_n35604_));
  OAI21_X1   g33168(.A1(pi0955), .A2(new_n32614_), .B(new_n35604_), .ZN(po1021));
  NAND2_X1   g33169(.A1(pi0866), .A2(pi0955), .ZN(new_n35606_));
  OAI21_X1   g33170(.A1(pi0955), .A2(new_n32490_), .B(new_n35606_), .ZN(po1022));
  NAND2_X1   g33171(.A1(pi0867), .A2(pi0955), .ZN(new_n35608_));
  OAI21_X1   g33172(.A1(pi0955), .A2(new_n32898_), .B(new_n35608_), .ZN(po1023));
  NAND2_X1   g33173(.A1(pi0868), .A2(pi0955), .ZN(new_n35610_));
  OAI21_X1   g33174(.A1(pi0955), .A2(new_n32608_), .B(new_n35610_), .ZN(po1024));
  NOR2_X1    g33175(.A1(new_n3041_), .A2(new_n4083_), .ZN(new_n35612_));
  NOR2_X1    g33176(.A1(new_n4091_), .A2(pi1093), .ZN(new_n35613_));
  OAI21_X1   g33177(.A1(new_n35612_), .A2(new_n35613_), .B(new_n2458_), .ZN(new_n35614_));
  NOR2_X1    g33178(.A1(new_n31383_), .A2(new_n4091_), .ZN(new_n35615_));
  NOR2_X1    g33179(.A1(new_n4083_), .A2(pi0123), .ZN(new_n35616_));
  OAI21_X1   g33180(.A1(new_n35615_), .A2(new_n35616_), .B(pi0228), .ZN(new_n35617_));
  NAND2_X1   g33181(.A1(new_n35614_), .A2(new_n35617_), .ZN(po1025));
  NAND2_X1   g33182(.A1(pi0870), .A2(pi0955), .ZN(new_n35619_));
  OAI21_X1   g33183(.A1(pi0955), .A2(new_n31362_), .B(new_n35619_), .ZN(po1026));
  NAND2_X1   g33184(.A1(pi0871), .A2(pi0955), .ZN(new_n35621_));
  OAI21_X1   g33185(.A1(pi0955), .A2(new_n32487_), .B(new_n35621_), .ZN(po1027));
  NAND2_X1   g33186(.A1(pi0872), .A2(pi0955), .ZN(new_n35623_));
  OAI21_X1   g33187(.A1(pi0955), .A2(new_n32481_), .B(new_n35623_), .ZN(po1028));
  NAND2_X1   g33188(.A1(pi0873), .A2(pi0955), .ZN(new_n35625_));
  OAI21_X1   g33189(.A1(pi0955), .A2(new_n32496_), .B(new_n35625_), .ZN(po1029));
  NAND2_X1   g33190(.A1(pi0874), .A2(pi0955), .ZN(new_n35627_));
  OAI21_X1   g33191(.A1(pi0955), .A2(new_n31338_), .B(new_n35627_), .ZN(po1030));
  NAND2_X1   g33192(.A1(new_n4729_), .A2(pi0123), .ZN(new_n35629_));
  OAI21_X1   g33193(.A1(pi0123), .A2(pi1136), .B(new_n35629_), .ZN(new_n35630_));
  NAND2_X1   g33194(.A1(pi1093), .A2(pi1136), .ZN(new_n35631_));
  AOI21_X1   g33195(.A1(new_n3041_), .A2(pi0875), .B(pi0228), .ZN(new_n35632_));
  AOI22_X1   g33196(.A1(new_n35630_), .A2(pi0228), .B1(new_n35631_), .B2(new_n35632_), .ZN(po1031));
  NAND2_X1   g33197(.A1(pi0876), .A2(pi0955), .ZN(new_n35634_));
  OAI21_X1   g33198(.A1(pi0955), .A2(new_n32493_), .B(new_n35634_), .ZN(po1032));
  NOR2_X1    g33199(.A1(new_n3041_), .A2(new_n4408_), .ZN(new_n35636_));
  NOR2_X1    g33200(.A1(new_n4416_), .A2(pi1093), .ZN(new_n35637_));
  OAI21_X1   g33201(.A1(new_n35636_), .A2(new_n35637_), .B(new_n2458_), .ZN(new_n35638_));
  NOR2_X1    g33202(.A1(new_n31383_), .A2(new_n4416_), .ZN(new_n35639_));
  NOR2_X1    g33203(.A1(new_n4408_), .A2(pi0123), .ZN(new_n35640_));
  OAI21_X1   g33204(.A1(new_n35639_), .A2(new_n35640_), .B(pi0228), .ZN(new_n35641_));
  NAND2_X1   g33205(.A1(new_n35638_), .A2(new_n35641_), .ZN(po1033));
  NOR2_X1    g33206(.A1(new_n3041_), .A2(new_n4565_), .ZN(new_n35643_));
  NOR2_X1    g33207(.A1(new_n4573_), .A2(pi1093), .ZN(new_n35644_));
  OAI21_X1   g33208(.A1(new_n35643_), .A2(new_n35644_), .B(new_n2458_), .ZN(new_n35645_));
  NOR2_X1    g33209(.A1(new_n31383_), .A2(new_n4573_), .ZN(new_n35646_));
  NOR2_X1    g33210(.A1(new_n4565_), .A2(pi0123), .ZN(new_n35647_));
  OAI21_X1   g33211(.A1(new_n35646_), .A2(new_n35647_), .B(pi0228), .ZN(new_n35648_));
  NAND2_X1   g33212(.A1(new_n35645_), .A2(new_n35648_), .ZN(po1034));
  NOR2_X1    g33213(.A1(new_n3041_), .A2(new_n4888_), .ZN(new_n35650_));
  NOR2_X1    g33214(.A1(new_n4893_), .A2(pi1093), .ZN(new_n35651_));
  OAI21_X1   g33215(.A1(new_n35650_), .A2(new_n35651_), .B(new_n2458_), .ZN(new_n35652_));
  NOR2_X1    g33216(.A1(new_n31383_), .A2(new_n4893_), .ZN(new_n35653_));
  NOR2_X1    g33217(.A1(new_n4888_), .A2(pi0123), .ZN(new_n35654_));
  OAI21_X1   g33218(.A1(new_n35653_), .A2(new_n35654_), .B(pi0228), .ZN(new_n35655_));
  NAND2_X1   g33219(.A1(new_n35652_), .A2(new_n35655_), .ZN(po1035));
  NAND2_X1   g33220(.A1(pi0880), .A2(pi0955), .ZN(new_n35657_));
  OAI21_X1   g33221(.A1(pi0955), .A2(new_n32753_), .B(new_n35657_), .ZN(po1036));
  NAND2_X1   g33222(.A1(pi0881), .A2(pi0955), .ZN(new_n35659_));
  OAI21_X1   g33223(.A1(pi0955), .A2(new_n32484_), .B(new_n35659_), .ZN(po1037));
  NAND2_X1   g33224(.A1(new_n35487_), .A2(pi1107), .ZN(new_n35661_));
  OAI21_X1   g33225(.A1(pi0883), .A2(new_n35487_), .B(new_n35661_), .ZN(po1039));
  NAND2_X1   g33226(.A1(new_n35487_), .A2(pi1124), .ZN(new_n35663_));
  OAI21_X1   g33227(.A1(pi0884), .A2(new_n35487_), .B(new_n35663_), .ZN(po1040));
  NAND2_X1   g33228(.A1(new_n35487_), .A2(pi1125), .ZN(new_n35665_));
  OAI21_X1   g33229(.A1(pi0885), .A2(new_n35487_), .B(new_n35665_), .ZN(po1041));
  NAND2_X1   g33230(.A1(new_n35487_), .A2(pi1109), .ZN(new_n35667_));
  OAI21_X1   g33231(.A1(pi0886), .A2(new_n35487_), .B(new_n35667_), .ZN(po1042));
  NAND2_X1   g33232(.A1(new_n35487_), .A2(pi1100), .ZN(new_n35669_));
  OAI21_X1   g33233(.A1(pi0887), .A2(new_n35487_), .B(new_n35669_), .ZN(po1043));
  NAND2_X1   g33234(.A1(new_n35487_), .A2(pi1120), .ZN(new_n35671_));
  OAI21_X1   g33235(.A1(pi0888), .A2(new_n35487_), .B(new_n35671_), .ZN(po1044));
  NAND2_X1   g33236(.A1(new_n35487_), .A2(pi1103), .ZN(new_n35673_));
  OAI21_X1   g33237(.A1(pi0889), .A2(new_n35487_), .B(new_n35673_), .ZN(po1045));
  NAND2_X1   g33238(.A1(new_n35487_), .A2(pi1126), .ZN(new_n35675_));
  OAI21_X1   g33239(.A1(pi0890), .A2(new_n35487_), .B(new_n35675_), .ZN(po1046));
  NAND2_X1   g33240(.A1(new_n35487_), .A2(pi1116), .ZN(new_n35677_));
  OAI21_X1   g33241(.A1(pi0891), .A2(new_n35487_), .B(new_n35677_), .ZN(po1047));
  NAND2_X1   g33242(.A1(new_n35487_), .A2(pi1101), .ZN(new_n35679_));
  OAI21_X1   g33243(.A1(pi0892), .A2(new_n35487_), .B(new_n35679_), .ZN(po1048));
  NAND2_X1   g33244(.A1(new_n35487_), .A2(pi1119), .ZN(new_n35681_));
  OAI21_X1   g33245(.A1(pi0894), .A2(new_n35487_), .B(new_n35681_), .ZN(po1050));
  NAND2_X1   g33246(.A1(new_n35487_), .A2(pi1113), .ZN(new_n35683_));
  OAI21_X1   g33247(.A1(pi0895), .A2(new_n35487_), .B(new_n35683_), .ZN(po1051));
  NAND2_X1   g33248(.A1(new_n35487_), .A2(pi1118), .ZN(new_n35685_));
  OAI21_X1   g33249(.A1(pi0896), .A2(new_n35487_), .B(new_n35685_), .ZN(po1052));
  NAND2_X1   g33250(.A1(new_n35487_), .A2(pi1129), .ZN(new_n35687_));
  OAI21_X1   g33251(.A1(pi0898), .A2(new_n35487_), .B(new_n35687_), .ZN(po1054));
  NAND2_X1   g33252(.A1(new_n35487_), .A2(pi1115), .ZN(new_n35689_));
  OAI21_X1   g33253(.A1(pi0899), .A2(new_n35487_), .B(new_n35689_), .ZN(po1055));
  NAND2_X1   g33254(.A1(new_n35487_), .A2(pi1110), .ZN(new_n35691_));
  OAI21_X1   g33255(.A1(pi0900), .A2(new_n35487_), .B(new_n35691_), .ZN(po1056));
  NAND2_X1   g33256(.A1(new_n35487_), .A2(pi1111), .ZN(new_n35693_));
  OAI21_X1   g33257(.A1(pi0902), .A2(new_n35487_), .B(new_n35693_), .ZN(po1058));
  NAND2_X1   g33258(.A1(new_n35487_), .A2(pi1121), .ZN(new_n35695_));
  OAI21_X1   g33259(.A1(pi0903), .A2(new_n35487_), .B(new_n35695_), .ZN(po1059));
  NAND2_X1   g33260(.A1(new_n35487_), .A2(pi1127), .ZN(new_n35697_));
  OAI21_X1   g33261(.A1(pi0904), .A2(new_n35487_), .B(new_n35697_), .ZN(po1060));
  NAND2_X1   g33262(.A1(new_n35487_), .A2(pi1131), .ZN(new_n35699_));
  OAI21_X1   g33263(.A1(pi0905), .A2(new_n35487_), .B(new_n35699_), .ZN(po1061));
  NAND2_X1   g33264(.A1(new_n35487_), .A2(pi1128), .ZN(new_n35701_));
  OAI21_X1   g33265(.A1(pi0906), .A2(new_n35487_), .B(new_n35701_), .ZN(po1062));
  NOR2_X1    g33266(.A1(new_n34118_), .A2(new_n5389_), .ZN(new_n35703_));
  INV_X1     g33267(.I(pi0624), .ZN(new_n35704_));
  NOR2_X1    g33268(.A1(new_n35704_), .A2(pi0979), .ZN(new_n35705_));
  OAI21_X1   g33269(.A1(new_n35703_), .A2(new_n35705_), .B(pi0782), .ZN(new_n35706_));
  INV_X1     g33270(.I(new_n35706_), .ZN(new_n35707_));
  NOR2_X1    g33271(.A1(new_n5389_), .A2(pi0615), .ZN(new_n35708_));
  INV_X1     g33272(.I(pi0604), .ZN(new_n35709_));
  NOR2_X1    g33273(.A1(new_n35709_), .A2(pi0979), .ZN(new_n35710_));
  OAI21_X1   g33274(.A1(new_n35708_), .A2(new_n35710_), .B(pi0782), .ZN(new_n35711_));
  INV_X1     g33275(.I(pi0782), .ZN(new_n35712_));
  NAND2_X1   g33276(.A1(new_n35712_), .A2(pi0907), .ZN(new_n35713_));
  AOI21_X1   g33277(.A1(new_n35711_), .A2(new_n35713_), .B(new_n35707_), .ZN(po1063));
  NAND2_X1   g33278(.A1(new_n35487_), .A2(pi1122), .ZN(new_n35715_));
  OAI21_X1   g33279(.A1(pi0908), .A2(new_n35487_), .B(new_n35715_), .ZN(po1064));
  NAND2_X1   g33280(.A1(new_n35487_), .A2(pi1105), .ZN(new_n35717_));
  OAI21_X1   g33281(.A1(pi0909), .A2(new_n35487_), .B(new_n35717_), .ZN(po1065));
  NAND2_X1   g33282(.A1(new_n35487_), .A2(pi1117), .ZN(new_n35719_));
  OAI21_X1   g33283(.A1(pi0910), .A2(new_n35487_), .B(new_n35719_), .ZN(po1066));
  NAND2_X1   g33284(.A1(new_n35487_), .A2(pi1130), .ZN(new_n35721_));
  OAI21_X1   g33285(.A1(pi0911), .A2(new_n35487_), .B(new_n35721_), .ZN(po1067));
  NAND2_X1   g33286(.A1(new_n35487_), .A2(pi1114), .ZN(new_n35723_));
  OAI21_X1   g33287(.A1(pi0912), .A2(new_n35487_), .B(new_n35723_), .ZN(po1068));
  NAND2_X1   g33288(.A1(new_n35487_), .A2(pi1106), .ZN(new_n35725_));
  OAI21_X1   g33289(.A1(pi0913), .A2(new_n35487_), .B(new_n35725_), .ZN(po1069));
  AND2_X2    g33290(.A1(pi0266), .A2(pi0992), .Z(new_n35727_));
  NAND2_X1   g33291(.A1(pi0280), .A2(pi0992), .ZN(new_n35728_));
  OAI22_X1   g33292(.A1(new_n35727_), .A2(pi0280), .B1(new_n4727_), .B2(new_n35728_), .ZN(po1070));
  NAND2_X1   g33293(.A1(new_n35487_), .A2(pi1108), .ZN(new_n35730_));
  OAI21_X1   g33294(.A1(pi0915), .A2(new_n35487_), .B(new_n35730_), .ZN(po1071));
  NAND2_X1   g33295(.A1(new_n35487_), .A2(pi1123), .ZN(new_n35732_));
  OAI21_X1   g33296(.A1(pi0916), .A2(new_n35487_), .B(new_n35732_), .ZN(po1072));
  NAND2_X1   g33297(.A1(new_n35487_), .A2(pi1112), .ZN(new_n35734_));
  OAI21_X1   g33298(.A1(pi0917), .A2(new_n35487_), .B(new_n35734_), .ZN(po1073));
  NAND2_X1   g33299(.A1(new_n35487_), .A2(pi1104), .ZN(new_n35736_));
  OAI21_X1   g33300(.A1(pi0918), .A2(new_n35487_), .B(new_n35736_), .ZN(po1074));
  NAND2_X1   g33301(.A1(new_n35487_), .A2(pi1102), .ZN(new_n35738_));
  OAI21_X1   g33302(.A1(pi0919), .A2(new_n35487_), .B(new_n35738_), .ZN(po1075));
  NAND2_X1   g33303(.A1(pi1093), .A2(pi1139), .ZN(new_n35740_));
  OAI21_X1   g33304(.A1(new_n4239_), .A2(pi1093), .B(new_n35740_), .ZN(po1076));
  INV_X1     g33305(.I(new_n35612_), .ZN(new_n35742_));
  OAI21_X1   g33306(.A1(new_n4081_), .A2(pi1093), .B(new_n35742_), .ZN(po1077));
  NAND2_X1   g33307(.A1(pi1093), .A2(pi1152), .ZN(new_n35744_));
  OAI21_X1   g33308(.A1(new_n33084_), .A2(pi1093), .B(new_n35744_), .ZN(po1078));
  NAND2_X1   g33309(.A1(pi1093), .A2(pi1154), .ZN(new_n35746_));
  OAI21_X1   g33310(.A1(new_n33076_), .A2(pi1093), .B(new_n35746_), .ZN(po1079));
  INV_X1     g33311(.I(pi0311), .ZN(new_n35748_));
  NOR4_X1    g33312(.A1(new_n32513_), .A2(new_n35748_), .A3(pi0300), .A4(pi0312), .ZN(po1080));
  NAND2_X1   g33313(.A1(pi1093), .A2(pi1155), .ZN(new_n35750_));
  OAI21_X1   g33314(.A1(new_n33052_), .A2(pi1093), .B(new_n35750_), .ZN(po1081));
  NAND2_X1   g33315(.A1(pi1093), .A2(pi1157), .ZN(new_n35752_));
  OAI21_X1   g33316(.A1(new_n32985_), .A2(pi1093), .B(new_n35752_), .ZN(po1082));
  NAND2_X1   g33317(.A1(pi1093), .A2(pi1145), .ZN(new_n35754_));
  OAI21_X1   g33318(.A1(new_n3514_), .A2(pi1093), .B(new_n35754_), .ZN(po1083));
  OAI21_X1   g33319(.A1(new_n4722_), .A2(pi1093), .B(new_n35631_), .ZN(po1084));
  NAND2_X1   g33320(.A1(pi1093), .A2(pi1144), .ZN(new_n35757_));
  OAI21_X1   g33321(.A1(new_n2442_), .A2(pi1093), .B(new_n35757_), .ZN(po1085));
  NAND2_X1   g33322(.A1(pi1093), .A2(pi1134), .ZN(new_n35759_));
  OAI21_X1   g33323(.A1(new_n5055_), .A2(pi1093), .B(new_n35759_), .ZN(po1086));
  NAND2_X1   g33324(.A1(pi1093), .A2(pi1150), .ZN(new_n35761_));
  OAI21_X1   g33325(.A1(new_n33092_), .A2(pi1093), .B(new_n35761_), .ZN(po1087));
  OAI21_X1   g33326(.A1(new_n3766_), .A2(pi1093), .B(new_n31380_), .ZN(po1088));
  INV_X1     g33327(.I(new_n35643_), .ZN(new_n35764_));
  OAI21_X1   g33328(.A1(new_n4563_), .A2(pi1093), .B(new_n35764_), .ZN(po1089));
  NAND2_X1   g33329(.A1(pi1093), .A2(pi1147), .ZN(new_n35766_));
  OAI21_X1   g33330(.A1(new_n32547_), .A2(pi1093), .B(new_n35766_), .ZN(po1090));
  INV_X1     g33331(.I(new_n35591_), .ZN(new_n35768_));
  OAI21_X1   g33332(.A1(new_n3924_), .A2(pi1093), .B(new_n35768_), .ZN(po1091));
  NAND2_X1   g33333(.A1(pi1093), .A2(pi1149), .ZN(new_n35770_));
  OAI21_X1   g33334(.A1(new_n33100_), .A2(pi1093), .B(new_n35770_), .ZN(po1092));
  NAND2_X1   g33335(.A1(pi1093), .A2(pi1148), .ZN(new_n35772_));
  OAI21_X1   g33336(.A1(new_n32524_), .A2(pi1093), .B(new_n35772_), .ZN(po1093));
  INV_X1     g33337(.I(new_n35650_), .ZN(new_n35774_));
  OAI21_X1   g33338(.A1(new_n4886_), .A2(pi1093), .B(new_n35774_), .ZN(po1094));
  NAND2_X1   g33339(.A1(pi1093), .A2(pi1146), .ZN(new_n35776_));
  OAI21_X1   g33340(.A1(new_n3341_), .A2(pi1093), .B(new_n35776_), .ZN(po1095));
  INV_X1     g33341(.I(new_n35636_), .ZN(new_n35778_));
  OAI21_X1   g33342(.A1(new_n4406_), .A2(pi1093), .B(new_n35778_), .ZN(po1096));
  NAND2_X1   g33343(.A1(pi1093), .A2(pi1153), .ZN(new_n35780_));
  OAI21_X1   g33344(.A1(new_n33064_), .A2(pi1093), .B(new_n35780_), .ZN(po1097));
  NAND2_X1   g33345(.A1(pi1093), .A2(pi1156), .ZN(new_n35782_));
  OAI21_X1   g33346(.A1(new_n33040_), .A2(pi1093), .B(new_n35782_), .ZN(po1098));
  NAND2_X1   g33347(.A1(pi1093), .A2(pi1151), .ZN(new_n35784_));
  OAI21_X1   g33348(.A1(new_n32996_), .A2(pi1093), .B(new_n35784_), .ZN(po1099));
  NAND2_X1   g33349(.A1(pi1093), .A2(pi1143), .ZN(new_n35786_));
  OAI21_X1   g33350(.A1(new_n3603_), .A2(pi1093), .B(new_n35786_), .ZN(po1100));
  NOR2_X1    g33351(.A1(new_n3043_), .A2(new_n27999_), .ZN(po1102));
  OAI21_X1   g33352(.A1(pi0782), .A2(new_n5692_), .B(new_n35706_), .ZN(po1103));
  XOR2_X1    g33353(.A1(pi0266), .A2(pi0992), .Z(po1104));
  NAND2_X1   g33354(.A1(pi0949), .A2(pi0954), .ZN(new_n35791_));
  OAI21_X1   g33355(.A1(pi0313), .A2(pi0954), .B(new_n35791_), .ZN(po1105));
  NOR3_X1    g33356(.A1(new_n6870_), .A2(new_n3044_), .A3(new_n3040_), .ZN(po1107));
  OAI21_X1   g33357(.A1(new_n3023_), .A2(new_n3040_), .B(new_n10900_), .ZN(po1112));
  NOR2_X1    g33358(.A1(new_n5930_), .A2(pi0782), .ZN(po1115));
  NOR2_X1    g33359(.A1(new_n5875_), .A2(pi0230), .ZN(po1116));
  NOR2_X1    g33360(.A1(new_n5990_), .A2(pi0782), .ZN(po1118));
  NOR2_X1    g33361(.A1(new_n5786_), .A2(pi0230), .ZN(po1122));
  NOR2_X1    g33362(.A1(new_n5995_), .A2(pi0230), .ZN(po1124));
  NOR2_X1    g33363(.A1(new_n5414_), .A2(pi0782), .ZN(po1125));
  NOR2_X1    g33364(.A1(new_n6054_), .A2(pi0230), .ZN(po1126));
  NOR2_X1    g33365(.A1(new_n5415_), .A2(pi0782), .ZN(po1127));
  NOR2_X1    g33366(.A1(new_n6115_), .A2(pi0230), .ZN(po1128));
  NOR2_X1    g33367(.A1(new_n5416_), .A2(pi0782), .ZN(po1129));
  NOR2_X1    g33368(.A1(new_n5935_), .A2(pi0230), .ZN(po1131));
  NOR2_X1    g33369(.A1(new_n6109_), .A2(pi0782), .ZN(po1132));
  NAND2_X1   g33370(.A1(new_n34118_), .A2(pi0615), .ZN(po1133));
  NOR2_X1    g33371(.A1(new_n5428_), .A2(new_n3040_), .ZN(po1135));
  NAND2_X1   g33372(.A1(new_n35709_), .A2(new_n35704_), .ZN(po1137));
  INV_X1     g33373(.I(pi0915), .ZN(po1146));
  INV_X1     g33374(.I(pi0913), .ZN(po1149));
  INV_X1     g33375(.I(pi0894), .ZN(po1150));
  INV_X1     g33376(.I(pi0905), .ZN(po1151));
  INV_X1     g33377(.I(pi0890), .ZN(po1153));
  INV_X1     g33378(.I(pi0906), .ZN(po1155));
  INV_X1     g33379(.I(pi0896), .ZN(po1156));
  INV_X1     g33380(.I(pi0909), .ZN(po1157));
  INV_X1     g33381(.I(pi0911), .ZN(po1158));
  INV_X1     g33382(.I(pi0908), .ZN(po1159));
  INV_X1     g33383(.I(pi0891), .ZN(po1160));
  INV_X1     g33384(.I(pi0902), .ZN(po1161));
  INV_X1     g33385(.I(pi0903), .ZN(po1162));
  INV_X1     g33386(.I(pi0883), .ZN(po1163));
  INV_X1     g33387(.I(pi0888), .ZN(po1164));
  INV_X1     g33388(.I(pi0919), .ZN(po1165));
  INV_X1     g33389(.I(pi0886), .ZN(po1166));
  INV_X1     g33390(.I(pi0912), .ZN(po1167));
  INV_X1     g33391(.I(pi0895), .ZN(po1168));
  INV_X1     g33392(.I(pi0916), .ZN(po1169));
  INV_X1     g33393(.I(pi0889), .ZN(po1170));
  INV_X1     g33394(.I(pi0900), .ZN(po1171));
  INV_X1     g33395(.I(pi0885), .ZN(po1172));
  INV_X1     g33396(.I(pi0904), .ZN(po1173));
  INV_X1     g33397(.I(pi0899), .ZN(po1174));
  INV_X1     g33398(.I(pi0918), .ZN(po1175));
  INV_X1     g33399(.I(pi0898), .ZN(po1176));
  INV_X1     g33400(.I(pi0917), .ZN(po1177));
  INV_X1     g33401(.I(pi0887), .ZN(po1179));
  INV_X1     g33402(.I(pi0884), .ZN(po1180));
  INV_X1     g33403(.I(pi0910), .ZN(po1181));
  INV_X1     g33404(.I(pi0892), .ZN(po1183));
  assign     po0166 = 1'b1;
  BUF_X16    g33405(.I(pi0668), .Z(po0000));
  BUF_X16    g33406(.I(pi0672), .Z(po0001));
  BUF_X16    g33407(.I(pi0664), .Z(po0002));
  BUF_X16    g33408(.I(pi0667), .Z(po0003));
  BUF_X16    g33409(.I(pi0676), .Z(po0004));
  BUF_X16    g33410(.I(pi0673), .Z(po0005));
  BUF_X16    g33411(.I(pi0675), .Z(po0006));
  BUF_X16    g33412(.I(pi0666), .Z(po0007));
  BUF_X16    g33413(.I(pi0679), .Z(po0008));
  BUF_X16    g33414(.I(pi0674), .Z(po0009));
  BUF_X16    g33415(.I(pi0663), .Z(po0010));
  BUF_X16    g33416(.I(pi0670), .Z(po0011));
  BUF_X16    g33417(.I(pi0677), .Z(po0012));
  BUF_X16    g33418(.I(pi0682), .Z(po0013));
  BUF_X16    g33419(.I(pi0671), .Z(po0014));
  BUF_X16    g33420(.I(pi0678), .Z(po0015));
  BUF_X16    g33421(.I(pi0718), .Z(po0016));
  BUF_X16    g33422(.I(pi0707), .Z(po0017));
  BUF_X16    g33423(.I(pi0708), .Z(po0018));
  BUF_X16    g33424(.I(pi0713), .Z(po0019));
  BUF_X16    g33425(.I(pi0711), .Z(po0020));
  BUF_X16    g33426(.I(pi0716), .Z(po0021));
  BUF_X16    g33427(.I(pi0733), .Z(po0022));
  BUF_X16    g33428(.I(pi0712), .Z(po0023));
  BUF_X16    g33429(.I(pi0689), .Z(po0024));
  BUF_X16    g33430(.I(pi0717), .Z(po0025));
  BUF_X16    g33431(.I(pi0692), .Z(po0026));
  BUF_X16    g33432(.I(pi0719), .Z(po0027));
  BUF_X16    g33433(.I(pi0722), .Z(po0028));
  BUF_X16    g33434(.I(pi0714), .Z(po0029));
  BUF_X16    g33435(.I(pi0720), .Z(po0030));
  BUF_X16    g33436(.I(pi0685), .Z(po0031));
  BUF_X16    g33437(.I(pi0837), .Z(po0032));
  BUF_X16    g33438(.I(pi0850), .Z(po0033));
  BUF_X16    g33439(.I(pi0872), .Z(po0034));
  BUF_X16    g33440(.I(pi0871), .Z(po0035));
  BUF_X16    g33441(.I(pi0881), .Z(po0036));
  BUF_X16    g33442(.I(pi0866), .Z(po0037));
  BUF_X16    g33443(.I(pi0876), .Z(po0038));
  BUF_X16    g33444(.I(pi0873), .Z(po0039));
  BUF_X16    g33445(.I(pi0874), .Z(po0040));
  BUF_X16    g33446(.I(pi0859), .Z(po0041));
  BUF_X16    g33447(.I(pi0855), .Z(po0042));
  BUF_X16    g33448(.I(pi0852), .Z(po0043));
  BUF_X16    g33449(.I(pi0870), .Z(po0044));
  BUF_X16    g33450(.I(pi0848), .Z(po0045));
  BUF_X16    g33451(.I(pi0865), .Z(po0046));
  BUF_X16    g33452(.I(pi0856), .Z(po0047));
  BUF_X16    g33453(.I(pi0853), .Z(po0048));
  BUF_X16    g33454(.I(pi0847), .Z(po0049));
  BUF_X16    g33455(.I(pi0857), .Z(po0050));
  BUF_X16    g33456(.I(pi0854), .Z(po0051));
  BUF_X16    g33457(.I(pi0858), .Z(po0052));
  BUF_X16    g33458(.I(pi0845), .Z(po0053));
  BUF_X16    g33459(.I(pi0838), .Z(po0054));
  BUF_X16    g33460(.I(pi0842), .Z(po0055));
  BUF_X16    g33461(.I(pi0843), .Z(po0056));
  BUF_X16    g33462(.I(pi0839), .Z(po0057));
  BUF_X16    g33463(.I(pi0844), .Z(po0058));
  BUF_X16    g33464(.I(pi0868), .Z(po0059));
  BUF_X16    g33465(.I(pi0851), .Z(po0060));
  BUF_X16    g33466(.I(pi0867), .Z(po0061));
  BUF_X16    g33467(.I(pi0880), .Z(po0062));
  BUF_X16    g33468(.I(pi0860), .Z(po0063));
  BUF_X16    g33469(.I(pi1030), .Z(po0064));
  BUF_X16    g33470(.I(pi1034), .Z(po0065));
  BUF_X16    g33471(.I(pi1015), .Z(po0066));
  BUF_X16    g33472(.I(pi1020), .Z(po0067));
  BUF_X16    g33473(.I(pi1025), .Z(po0068));
  BUF_X16    g33474(.I(pi1005), .Z(po0069));
  BUF_X16    g33475(.I(pi0996), .Z(po0070));
  BUF_X16    g33476(.I(pi1012), .Z(po0071));
  BUF_X16    g33477(.I(pi0993), .Z(po0072));
  BUF_X16    g33478(.I(pi1016), .Z(po0073));
  BUF_X16    g33479(.I(pi1021), .Z(po0074));
  BUF_X16    g33480(.I(pi1010), .Z(po0075));
  BUF_X16    g33481(.I(pi1027), .Z(po0076));
  BUF_X16    g33482(.I(pi1018), .Z(po0077));
  BUF_X16    g33483(.I(pi1017), .Z(po0078));
  BUF_X16    g33484(.I(pi1024), .Z(po0079));
  BUF_X16    g33485(.I(pi1009), .Z(po0080));
  BUF_X16    g33486(.I(pi1032), .Z(po0081));
  BUF_X16    g33487(.I(pi1003), .Z(po0082));
  BUF_X16    g33488(.I(pi0997), .Z(po0083));
  BUF_X16    g33489(.I(pi1013), .Z(po0084));
  BUF_X16    g33490(.I(pi1011), .Z(po0085));
  BUF_X16    g33491(.I(pi1008), .Z(po0086));
  BUF_X16    g33492(.I(pi1019), .Z(po0087));
  BUF_X16    g33493(.I(pi1031), .Z(po0088));
  BUF_X16    g33494(.I(pi1022), .Z(po0089));
  BUF_X16    g33495(.I(pi1000), .Z(po0090));
  BUF_X16    g33496(.I(pi1023), .Z(po0091));
  BUF_X16    g33497(.I(pi1002), .Z(po0092));
  BUF_X16    g33498(.I(pi1026), .Z(po0093));
  BUF_X16    g33499(.I(pi1006), .Z(po0094));
  BUF_X16    g33500(.I(pi0998), .Z(po0095));
  BUF_X16    g33501(.I(pi0031), .Z(po0096));
  BUF_X16    g33502(.I(pi0080), .Z(po0097));
  BUF_X16    g33503(.I(pi0893), .Z(po0098));
  BUF_X16    g33504(.I(pi0467), .Z(po0099));
  BUF_X16    g33505(.I(pi0078), .Z(po0100));
  BUF_X16    g33506(.I(pi0112), .Z(po0101));
  BUF_X16    g33507(.I(pi0013), .Z(po0102));
  BUF_X16    g33508(.I(pi0025), .Z(po0103));
  BUF_X16    g33509(.I(pi0226), .Z(po0104));
  BUF_X16    g33510(.I(pi0127), .Z(po0105));
  BUF_X16    g33511(.I(pi0822), .Z(po0106));
  BUF_X16    g33512(.I(pi0808), .Z(po0107));
  BUF_X16    g33513(.I(pi0227), .Z(po0108));
  BUF_X16    g33514(.I(pi0477), .Z(po0109));
  BUF_X16    g33515(.I(pi0834), .Z(po0110));
  BUF_X16    g33516(.I(pi0229), .Z(po0111));
  BUF_X16    g33517(.I(pi0012), .Z(po0112));
  BUF_X16    g33518(.I(pi0011), .Z(po0113));
  BUF_X16    g33519(.I(pi0010), .Z(po0114));
  BUF_X16    g33520(.I(pi0009), .Z(po0115));
  BUF_X16    g33521(.I(pi0008), .Z(po0116));
  BUF_X16    g33522(.I(pi0007), .Z(po0117));
  BUF_X16    g33523(.I(pi0006), .Z(po0118));
  BUF_X16    g33524(.I(pi0005), .Z(po0119));
  BUF_X16    g33525(.I(pi0004), .Z(po0120));
  BUF_X16    g33526(.I(pi0003), .Z(po0121));
  BUF_X16    g33527(.I(pi0000), .Z(po0122));
  BUF_X16    g33528(.I(pi0002), .Z(po0123));
  BUF_X16    g33529(.I(pi0001), .Z(po0124));
  BUF_X16    g33530(.I(pi0310), .Z(po0125));
  BUF_X16    g33531(.I(pi0302), .Z(po0126));
  BUF_X16    g33532(.I(pi0475), .Z(po0127));
  BUF_X16    g33533(.I(pi0474), .Z(po0128));
  BUF_X16    g33534(.I(pi0466), .Z(po0129));
  BUF_X16    g33535(.I(pi0473), .Z(po0130));
  BUF_X16    g33536(.I(pi0471), .Z(po0131));
  BUF_X16    g33537(.I(pi0472), .Z(po0132));
  BUF_X16    g33538(.I(pi0470), .Z(po0133));
  BUF_X16    g33539(.I(pi0469), .Z(po0134));
  BUF_X16    g33540(.I(pi0465), .Z(po0135));
  BUF_X16    g33541(.I(pi1028), .Z(po0136));
  BUF_X16    g33542(.I(pi1033), .Z(po0137));
  BUF_X16    g33543(.I(pi0995), .Z(po0138));
  BUF_X16    g33544(.I(pi0994), .Z(po0139));
  BUF_X16    g33545(.I(pi0028), .Z(po0140));
  BUF_X16    g33546(.I(pi0027), .Z(po0141));
  BUF_X16    g33547(.I(pi0026), .Z(po0142));
  BUF_X16    g33548(.I(pi0029), .Z(po0143));
  BUF_X16    g33549(.I(pi0015), .Z(po0144));
  BUF_X16    g33550(.I(pi0014), .Z(po0145));
  BUF_X16    g33551(.I(pi0021), .Z(po0146));
  BUF_X16    g33552(.I(pi0020), .Z(po0147));
  BUF_X16    g33553(.I(pi0019), .Z(po0148));
  BUF_X16    g33554(.I(pi0018), .Z(po0149));
  BUF_X16    g33555(.I(pi0017), .Z(po0150));
  BUF_X16    g33556(.I(pi0016), .Z(po0151));
  BUF_X16    g33557(.I(pi1096), .Z(po0152));
  BUF_X16    g33558(.I(pi0228), .Z(po0168));
  BUF_X16    g33559(.I(pi0022), .Z(po0169));
  BUF_X16    g33560(.I(pi1089), .Z(po0179));
  BUF_X16    g33561(.I(pi0023), .Z(po0180));
  OAI22_X1   g33562(.A1(new_n5466_), .A2(new_n3425_), .B1(new_n2582_), .B2(new_n5296_), .ZN(po0181));
  BUF_X16    g33563(.I(pi0037), .Z(po0188));
  BUF_X16    g33564(.I(pi0117), .Z(po0263));
  BUF_X16    g33565(.I(pi0131), .Z(po0285));
  BUF_X16    g33566(.I(pi0232), .Z(po0386));
  BUF_X16    g33567(.I(pi0236), .Z(po0388));
  BUF_X16    g33568(.I(pi0583), .Z(po0636));
  BUF_X16    g33569(.I(pi0067), .Z(po1053));
  BUF_X16    g33570(.I(pi1134), .Z(po1108));
  BUF_X16    g33571(.I(pi0964), .Z(po1109));
  BUF_X16    g33572(.I(pi0965), .Z(po1111));
  BUF_X16    g33573(.I(pi0991), .Z(po1113));
  BUF_X16    g33574(.I(pi0985), .Z(po1114));
  BUF_X16    g33575(.I(pi1014), .Z(po1117));
  BUF_X16    g33576(.I(pi1029), .Z(po1119));
  BUF_X16    g33577(.I(pi1004), .Z(po1120));
  BUF_X16    g33578(.I(pi1007), .Z(po1121));
  BUF_X16    g33579(.I(pi1135), .Z(po1123));
  BUF_X16    g33580(.I(pi1064), .Z(po1134));
  BUF_X16    g33581(.I(pi0299), .Z(po1136));
  BUF_X16    g33582(.I(pi1075), .Z(po1138));
  BUF_X16    g33583(.I(pi1052), .Z(po1139));
  BUF_X16    g33584(.I(pi0771), .Z(po1140));
  BUF_X16    g33585(.I(pi0765), .Z(po1141));
  BUF_X16    g33586(.I(pi0605), .Z(po1142));
  BUF_X16    g33587(.I(pi0601), .Z(po1143));
  BUF_X16    g33588(.I(pi0278), .Z(po1144));
  BUF_X16    g33589(.I(pi0279), .Z(po1145));
  BUF_X16    g33590(.I(pi1095), .Z(po1152));
  BUF_X16    g33591(.I(pi1094), .Z(po1154));
  BUF_X16    g33592(.I(pi1187), .Z(po1184));
  BUF_X16    g33593(.I(pi1172), .Z(po1185));
  BUF_X16    g33594(.I(pi1170), .Z(po1186));
  BUF_X16    g33595(.I(pi1138), .Z(po1187));
  BUF_X16    g33596(.I(pi1177), .Z(po1188));
  BUF_X16    g33597(.I(pi1178), .Z(po1189));
  BUF_X16    g33598(.I(pi0863), .Z(po1190));
  BUF_X16    g33599(.I(pi1203), .Z(po1191));
  BUF_X16    g33600(.I(pi1185), .Z(po1192));
  BUF_X16    g33601(.I(pi1171), .Z(po1193));
  BUF_X16    g33602(.I(pi1192), .Z(po1194));
  BUF_X16    g33603(.I(pi1137), .Z(po1195));
  BUF_X16    g33604(.I(pi1186), .Z(po1196));
  BUF_X16    g33605(.I(pi1165), .Z(po1197));
  BUF_X16    g33606(.I(pi1164), .Z(po1198));
  BUF_X16    g33607(.I(pi1098), .Z(po1199));
  BUF_X16    g33608(.I(pi1183), .Z(po1200));
  BUF_X16    g33609(.I(pi0230), .Z(po1201));
  BUF_X16    g33610(.I(pi1169), .Z(po1202));
  BUF_X16    g33611(.I(pi1136), .Z(po1203));
  BUF_X16    g33612(.I(pi1181), .Z(po1204));
  BUF_X16    g33613(.I(pi0849), .Z(po1205));
  BUF_X16    g33614(.I(pi1193), .Z(po1206));
  BUF_X16    g33615(.I(pi1182), .Z(po1207));
  BUF_X16    g33616(.I(pi1168), .Z(po1208));
  BUF_X16    g33617(.I(pi1175), .Z(po1209));
  BUF_X16    g33618(.I(pi1191), .Z(po1210));
  BUF_X16    g33619(.I(pi1099), .Z(po1211));
  BUF_X16    g33620(.I(pi1174), .Z(po1212));
  BUF_X16    g33621(.I(pi1179), .Z(po1213));
  BUF_X16    g33622(.I(pi1202), .Z(po1214));
  BUF_X16    g33623(.I(pi1176), .Z(po1215));
  BUF_X16    g33624(.I(pi1173), .Z(po1216));
  BUF_X16    g33625(.I(pi1201), .Z(po1217));
  BUF_X16    g33626(.I(pi1167), .Z(po1218));
  BUF_X16    g33627(.I(pi0840), .Z(po1219));
  BUF_X16    g33628(.I(pi1189), .Z(po1220));
  BUF_X16    g33629(.I(pi1195), .Z(po1221));
  BUF_X16    g33630(.I(pi0864), .Z(po1222));
  BUF_X16    g33631(.I(pi1190), .Z(po1223));
  BUF_X16    g33632(.I(pi1188), .Z(po1224));
  BUF_X16    g33633(.I(pi1180), .Z(po1225));
  BUF_X16    g33634(.I(pi1194), .Z(po1226));
  BUF_X16    g33635(.I(pi1097), .Z(po1227));
  BUF_X16    g33636(.I(pi1166), .Z(po1228));
  BUF_X16    g33637(.I(pi1200), .Z(po1229));
  BUF_X16    g33638(.I(pi1184), .Z(po1230));
endmodule


