// Benchmark "mem_ctrl" written by ABC on Mon Sep 11 23:44:13 2023

module mem_ctrl ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_,
    new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_,
    new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_,
    new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_,
    new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_,
    new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_,
    new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_,
    new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_,
    new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_,
    new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_,
    new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_,
    new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2989_, new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_,
    new_n2996_, new_n2997_, new_n2998_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3143_, new_n3146_, new_n3147_,
    new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_,
    new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_,
    new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_,
    new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_,
    new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_,
    new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_,
    new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_,
    new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_,
    new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_,
    new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_,
    new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_,
    new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_,
    new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_,
    new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_,
    new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_,
    new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_,
    new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_,
    new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_,
    new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_,
    new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_,
    new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_,
    new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_,
    new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_,
    new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_,
    new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_,
    new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_,
    new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_,
    new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_,
    new_n3377_, new_n3378_, new_n3379_, new_n3386_, new_n3391_, new_n3392_,
    new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_,
    new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_,
    new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3444_, new_n3445_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3533_, new_n3534_, new_n3535_,
    new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_,
    new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3548_,
    new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_,
    new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_,
    new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_,
    new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_,
    new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_,
    new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_,
    new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_,
    new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_,
    new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_,
    new_n3603_, new_n3604_, new_n3605_, new_n3608_, new_n3609_, new_n3610_,
    new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_,
    new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_,
    new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_,
    new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_,
    new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_,
    new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_,
    new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_,
    new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_,
    new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_,
    new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_,
    new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_,
    new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_,
    new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_,
    new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_,
    new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_,
    new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_,
    new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_,
    new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_,
    new_n3927_, new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_,
    new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_,
    new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_,
    new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_,
    new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_,
    new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_,
    new_n3971_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_,
    new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_,
    new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_,
    new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_,
    new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_,
    new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_,
    new_n4112_, new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_,
    new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_,
    new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_,
    new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_,
    new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_,
    new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_,
    new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_,
    new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_,
    new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_,
    new_n4167_, new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_,
    new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_,
    new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_,
    new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_,
    new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_,
    new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_,
    new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_,
    new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_,
    new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_,
    new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_,
    new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_,
    new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_,
    new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_,
    new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_,
    new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_,
    new_n4257_, new_n4258_, new_n4259_, new_n4261_, new_n4262_, new_n4263_,
    new_n4264_, new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_,
    new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_,
    new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_,
    new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_,
    new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_,
    new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_,
    new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_,
    new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_,
    new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_,
    new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_,
    new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4356_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4402_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_,
    new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_,
    new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_,
    new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_,
    new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_,
    new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_,
    new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_,
    new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_,
    new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_,
    new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_,
    new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_,
    new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_,
    new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_,
    new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_,
    new_n4495_, new_n4496_, new_n4497_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4543_, new_n4544_, new_n4545_,
    new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_,
    new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_,
    new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_,
    new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_,
    new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_,
    new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_,
    new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_,
    new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_,
    new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_,
    new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_,
    new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4696_,
    new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_,
    new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_,
    new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_,
    new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_,
    new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_,
    new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_,
    new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_,
    new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_,
    new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_,
    new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_,
    new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_,
    new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_,
    new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_,
    new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_,
    new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_,
    new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_,
    new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_,
    new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_,
    new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_,
    new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_,
    new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_,
    new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_,
    new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_,
    new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_,
    new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5113_, new_n5114_,
    new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_,
    new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_,
    new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_,
    new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_,
    new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_,
    new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_,
    new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_,
    new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_,
    new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_,
    new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_,
    new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5180_, new_n5181_,
    new_n5182_, new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_,
    new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_,
    new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_,
    new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_,
    new_n5207_, new_n5208_, new_n5209_, new_n5212_, new_n5213_, new_n5214_,
    new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_,
    new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_,
    new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_,
    new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_,
    new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_,
    new_n5245_, new_n5246_, new_n5247_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_,
    new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_,
    new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_,
    new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_,
    new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_,
    new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_,
    new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_,
    new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_,
    new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_,
    new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_,
    new_n5500_, new_n5501_, new_n5502_, new_n5504_, new_n5505_, new_n5506_,
    new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_,
    new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_,
    new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_,
    new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_,
    new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_,
    new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_,
    new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_,
    new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_,
    new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_,
    new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_,
    new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_,
    new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_,
    new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_,
    new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_,
    new_n5591_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5645_, new_n5646_,
    new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_,
    new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_,
    new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_,
    new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_,
    new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_,
    new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_,
    new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_,
    new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_,
    new_n5695_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_,
    new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_,
    new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_,
    new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5749_, new_n5750_,
    new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_,
    new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_,
    new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_,
    new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_,
    new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_,
    new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_,
    new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_,
    new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_,
    new_n5799_, new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5805_,
    new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_,
    new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_,
    new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_,
    new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_,
    new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_,
    new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_,
    new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_,
    new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5853_, new_n5854_,
    new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_,
    new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_,
    new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_,
    new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_,
    new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5898_,
    new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_,
    new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_,
    new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_,
    new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_,
    new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5929_,
    new_n5930_, new_n5931_, new_n5932_, new_n5934_, new_n5936_, new_n5938_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_,
    new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_,
    new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_,
    new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_,
    new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_,
    new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_,
    new_n6126_, new_n6127_, new_n6130_, new_n6131_, new_n6132_, new_n6133_,
    new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_,
    new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_,
    new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_,
    new_n6152_, new_n6153_, new_n6154_, new_n6156_, new_n6160_, new_n6180_,
    new_n6181_, new_n6182_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6202_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_,
    new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_,
    new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_,
    new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_,
    new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_,
    new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_,
    new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_,
    new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_,
    new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_,
    new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_,
    new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_,
    new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_,
    new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_,
    new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_,
    new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_,
    new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_,
    new_n6440_, new_n6441_, new_n6442_, new_n6445_, new_n6446_, new_n6448_,
    new_n6452_, new_n6453_, new_n6460_, new_n6462_, new_n6467_, new_n6468_,
    new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6481_, new_n6482_, new_n6488_,
    new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_,
    new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_,
    new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_,
    new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_,
    new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_,
    new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_,
    new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_,
    new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_,
    new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_,
    new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_,
    new_n6549_, new_n6551_, new_n6554_, new_n6556_, new_n6558_, new_n6559_,
    new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_,
    new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_,
    new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_,
    new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6591_, new_n6592_,
    new_n6593_, new_n6594_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_,
    new_n6609_, new_n6610_, new_n6611_, new_n6619_, new_n6620_, new_n6621_,
    new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_,
    new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_,
    new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_,
    new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6645_,
    new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_,
    new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_,
    new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_, new_n6663_,
    new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_,
    new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_,
    new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_,
    new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_,
    new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_,
    new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_,
    new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_, new_n6705_,
    new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_,
    new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_,
    new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_, new_n6723_,
    new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_, new_n6729_,
    new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_, new_n6735_,
    new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_, new_n6741_,
    new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_, new_n6747_,
    new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_,
    new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_, new_n6759_,
    new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_, new_n6765_,
    new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_, new_n6771_,
    new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_, new_n6777_,
    new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_, new_n6783_,
    new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_,
    new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_, new_n6795_,
    new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n6801_,
    new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_, new_n6807_,
    new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_,
    new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_, new_n6819_,
    new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_, new_n6825_,
    new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_, new_n6831_,
    new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_, new_n6837_,
    new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_, new_n6843_,
    new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6849_,
    new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_, new_n6855_,
    new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_, new_n6861_,
    new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_, new_n6867_,
    new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_, new_n6873_,
    new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_, new_n6879_,
    new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_, new_n6885_,
    new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_, new_n6891_,
    new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_, new_n6897_,
    new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_, new_n6903_,
    new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_, new_n6909_,
    new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_, new_n6915_,
    new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_, new_n6921_,
    new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_,
    new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_, new_n6933_,
    new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_, new_n6939_,
    new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_, new_n6945_,
    new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6951_, new_n6952_,
    new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_,
    new_n6959_, new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_,
    new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_,
    new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_,
    new_n6978_, new_n6979_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_,
    new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_,
    new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_,
    new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_,
    new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_,
    new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_,
    new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_,
    new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_,
    new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_,
    new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_,
    new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_,
    new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_,
    new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_,
    new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_,
    new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_,
    new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_, new_n7106_,
    new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_,
    new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_,
    new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_,
    new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_,
    new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_,
    new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_,
    new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_,
    new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_,
    new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_,
    new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_,
    new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_,
    new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_,
    new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_,
    new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_,
    new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_,
    new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_,
    new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_,
    new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_,
    new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_,
    new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_,
    new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_,
    new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_,
    new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_,
    new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_,
    new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_,
    new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_,
    new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_,
    new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_,
    new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_,
    new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_,
    new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_,
    new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_,
    new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_,
    new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_,
    new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_,
    new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_,
    new_n7323_, new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_,
    new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_,
    new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7405_, new_n7406_, new_n7409_, new_n7410_,
    new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_,
    new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7423_, new_n7424_,
    new_n7425_, new_n7426_, new_n7427_, new_n7430_, new_n7431_, new_n7440_,
    new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_,
    new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_,
    new_n7453_, new_n7454_, new_n7459_, new_n7460_, new_n7461_, new_n7462_,
    new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_, new_n7468_,
    new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_, new_n7474_,
    new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_, new_n7480_,
    new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_,
    new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_,
    new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_,
    new_n7499_, new_n7504_, new_n7505_, new_n7506_, new_n7511_, new_n7513_,
    new_n7514_, new_n7517_, new_n7518_, new_n7519_, new_n7531_, new_n7532_,
    new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_,
    new_n7556_, new_n7559_, new_n7560_, new_n7564_, new_n7565_, new_n7573_,
    new_n7593_, new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_,
    new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_,
    new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_,
    new_n7612_, new_n7615_, new_n7616_, new_n7620_, new_n7621_, new_n7622_,
    new_n7623_, new_n7624_, new_n7627_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_,
    new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_,
    new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_,
    new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_,
    new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_,
    new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_,
    new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_,
    new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_,
    new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_,
    new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7735_,
    new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_,
    new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_,
    new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_,
    new_n7754_, new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_,
    new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_,
    new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_,
    new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_,
    new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_,
    new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_,
    new_n7809_, new_n7810_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7832_, new_n7833_, new_n7834_, new_n7835_,
    new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_,
    new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_,
    new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_,
    new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_,
    new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_,
    new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_,
    new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_,
    new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_,
    new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_,
    new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_,
    new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_,
    new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_,
    new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_,
    new_n7915_, new_n7916_, new_n7918_, new_n7919_, new_n7920_, new_n7921_,
    new_n7922_, new_n7923_, new_n7924_, new_n7926_, new_n7927_, new_n7928_,
    new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_,
    new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_,
    new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_,
    new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_,
    new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_,
    new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_,
    new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_,
    new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_,
    new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_,
    new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_,
    new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_,
    new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_,
    new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_,
    new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_,
    new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_,
    new_n8019_, new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_,
    new_n8025_, new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_,
    new_n8031_, new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_,
    new_n8037_, new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_,
    new_n8043_, new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_,
    new_n8049_, new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_,
    new_n8055_, new_n8056_, new_n8057_, new_n8058_, new_n8059_, new_n8061_,
    new_n8062_, new_n8063_, new_n8064_, new_n8067_, new_n8070_, new_n8071_,
    new_n8072_, new_n8074_, new_n8075_, new_n8076_, new_n8077_, new_n8078_,
    new_n8079_, new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_,
    new_n8085_, new_n8086_, new_n8087_, new_n8088_, new_n8089_, new_n8090_,
    new_n8091_, new_n8092_, new_n8093_, new_n8094_, new_n8095_, new_n8096_,
    new_n8097_, new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_,
    new_n8103_, new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8108_,
    new_n8109_, new_n8110_, new_n8111_, new_n8112_, new_n8113_, new_n8114_,
    new_n8115_, new_n8116_, new_n8117_, new_n8118_, new_n8119_, new_n8120_,
    new_n8121_, new_n8122_, new_n8123_, new_n8124_, new_n8125_, new_n8126_,
    new_n8127_, new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_,
    new_n8133_, new_n8134_, new_n8135_, new_n8136_, new_n8137_, new_n8138_,
    new_n8139_, new_n8140_, new_n8141_, new_n8142_, new_n8143_, new_n8144_,
    new_n8145_, new_n8146_, new_n8147_, new_n8148_, new_n8149_, new_n8150_,
    new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_, new_n8156_,
    new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_, new_n8162_,
    new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_, new_n8168_,
    new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_, new_n8174_,
    new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_,
    new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_,
    new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_,
    new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_,
    new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_,
    new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_, new_n8210_,
    new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8215_, new_n8216_,
    new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_, new_n8222_,
    new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_, new_n8228_,
    new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_, new_n8234_,
    new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_, new_n8240_,
    new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_, new_n8247_,
    new_n8248_, new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_,
    new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_,
    new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_,
    new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_,
    new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_,
    new_n8278_, new_n8279_, new_n8280_, new_n8284_, new_n8287_, new_n8288_,
    new_n8289_, new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_,
    new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_,
    new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_,
    new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_,
    new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_,
    new_n8320_, new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_,
    new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_,
    new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_,
    new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_,
    new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_,
    new_n8369_, new_n8371_, new_n8373_, new_n8374_, new_n8375_, new_n8376_,
    new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_,
    new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_,
    new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_,
    new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_,
    new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_,
    new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_,
    new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8420_,
    new_n8421_, new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_,
    new_n8428_, new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8434_,
    new_n8435_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8446_, new_n8447_, new_n8448_,
    new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_,
    new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_,
    new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_,
    new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_,
    new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_,
    new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_,
    new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_,
    new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_, new_n8503_,
    new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_, new_n8509_,
    new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_, new_n8515_,
    new_n8516_, new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_,
    new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_,
    new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_,
    new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_,
    new_n8541_, new_n8542_, new_n8543_, new_n8544_, new_n8546_, new_n8547_,
    new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8557_, new_n8558_, new_n8559_, new_n8560_,
    new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_,
    new_n8567_, new_n8568_, new_n8569_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8588_,
    new_n8589_, new_n8590_, new_n8592_, new_n8593_, new_n8595_, new_n8596_,
    new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8603_,
    new_n8604_, new_n8606_, new_n8607_, new_n8609_, new_n8610_, new_n8611_,
    new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8618_, new_n8619_,
    new_n8620_, new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_,
    new_n8627_, new_n8628_, new_n8629_, new_n8631_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8637_, new_n8639_, new_n8640_, new_n8641_,
    new_n8642_, new_n8643_, new_n8644_, new_n8646_, new_n8647_, new_n8648_,
    new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_, new_n8654_,
    new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_, new_n8661_,
    new_n8662_, new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_,
    new_n8668_, new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_,
    new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_,
    new_n8681_, new_n8682_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8701_, new_n8702_, new_n8703_, new_n8705_, new_n8706_, new_n8708_,
    new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_, new_n8714_,
    new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_, new_n8720_,
    new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_, new_n8726_,
    new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_, new_n8732_,
    new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_, new_n8738_,
    new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_, new_n8744_,
    new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8750_,
    new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_,
    new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_, new_n8762_,
    new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_, new_n8768_,
    new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_, new_n8774_,
    new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_, new_n8780_,
    new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_, new_n8786_,
    new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_, new_n8792_,
    new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_, new_n8798_,
    new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_, new_n8804_,
    new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_, new_n8810_,
    new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_, new_n8816_,
    new_n8817_, new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8946_,
    new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_,
    new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_,
    new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_,
    new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_,
    new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_,
    new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_,
    new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_,
    new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_,
    new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_,
    new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_,
    new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_,
    new_n9013_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9051_, new_n9065_, new_n9106_, new_n9107_, new_n9109_,
    new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9120_,
    new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_,
    new_n9127_, new_n9128_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_,
    new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_,
    new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_,
    new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_,
    new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_,
    new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_,
    new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_,
    new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_,
    new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_,
    new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_,
    new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_,
    new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_,
    new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_,
    new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_,
    new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_,
    new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_,
    new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_,
    new_n9334_, new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_,
    new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_,
    new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_,
    new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_,
    new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_,
    new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_,
    new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_,
    new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_,
    new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_,
    new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_,
    new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_,
    new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_,
    new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_,
    new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_,
    new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_,
    new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_,
    new_n9432_, new_n9442_, new_n9443_, new_n9447_, new_n9448_, new_n9449_,
    new_n9450_, new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_,
    new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_,
    new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_,
    new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_,
    new_n9485_, new_n9486_, new_n9487_, new_n9489_, new_n9490_, new_n9491_,
    new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_,
    new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_,
    new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9641_, new_n9642_,
    new_n9643_, new_n9644_, new_n9645_, new_n9647_, new_n9648_, new_n9649_,
    new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_,
    new_n9658_, new_n9659_, new_n9660_, new_n9662_, new_n9663_, new_n9665_,
    new_n9667_, new_n9668_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9683_, new_n9684_, new_n9685_, new_n9686_,
    new_n9687_, new_n9689_, new_n9690_, new_n9692_, new_n9693_, new_n9694_,
    new_n9695_, new_n9696_, new_n9698_, new_n9699_, new_n9700_, new_n9701_,
    new_n9702_, new_n9703_, new_n9704_, new_n9706_, new_n9707_, new_n9708_,
    new_n9709_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_,
    new_n9722_, new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_,
    new_n9729_, new_n9730_, new_n9731_, new_n9733_, new_n9734_, new_n9735_,
    new_n9736_, new_n9737_, new_n9738_, new_n9740_, new_n9741_, new_n9742_,
    new_n9743_, new_n9745_, new_n9746_, new_n9747_, new_n9749_, new_n9750_,
    new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_,
    new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_,
    new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_,
    new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_,
    new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_,
    new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_,
    new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_,
    new_n9793_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9804_, new_n9805_, new_n9806_,
    new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_,
    new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_,
    new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_,
    new_n9825_, new_n9826_, new_n9827_, new_n9829_, new_n9830_, new_n9831_,
    new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_,
    new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9847_, new_n9849_,
    new_n9850_, new_n9852_, new_n9854_, new_n9855_, new_n9856_, new_n9858_,
    new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_,
    new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9893_, new_n9894_, new_n9896_, new_n9897_, new_n9898_, new_n9899_,
    new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9905_, new_n9906_,
    new_n9907_, new_n9909_, new_n9911_, new_n9912_, new_n9913_, new_n9914_,
    new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_,
    new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_,
    new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_,
    new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_,
    new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9944_, new_n9945_,
    new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_,
    new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9969_, new_n9970_,
    new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_,
    new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_,
    new_n9983_, new_n9985_, new_n9987_, new_n9988_, new_n9989_, new_n9990_,
    new_n9991_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10008_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10037_, new_n10038_, new_n10039_, new_n10040_, new_n10041_,
    new_n10042_, new_n10043_, new_n10044_, new_n10045_, new_n10046_,
    new_n10047_, new_n10048_, new_n10049_, new_n10050_, new_n10051_,
    new_n10052_, new_n10054_, new_n10055_, new_n10056_, new_n10057_,
    new_n10058_, new_n10059_, new_n10060_, new_n10061_, new_n10062_,
    new_n10063_, new_n10064_, new_n10065_, new_n10066_, new_n10067_,
    new_n10068_, new_n10069_, new_n10070_, new_n10071_, new_n10072_,
    new_n10073_, new_n10074_, new_n10075_, new_n10076_, new_n10077_,
    new_n10078_, new_n10079_, new_n10080_, new_n10081_, new_n10082_,
    new_n10083_, new_n10084_, new_n10085_, new_n10086_, new_n10088_,
    new_n10089_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10133_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10219_, new_n10220_, new_n10221_,
    new_n10222_, new_n10223_, new_n10224_, new_n10225_, new_n10226_,
    new_n10227_, new_n10228_, new_n10229_, new_n10230_, new_n10231_,
    new_n10232_, new_n10233_, new_n10234_, new_n10235_, new_n10236_,
    new_n10237_, new_n10238_, new_n10239_, new_n10240_, new_n10241_,
    new_n10242_, new_n10243_, new_n10244_, new_n10245_, new_n10246_,
    new_n10247_, new_n10248_, new_n10249_, new_n10250_, new_n10251_,
    new_n10252_, new_n10253_, new_n10255_, new_n10256_, new_n10257_,
    new_n10258_, new_n10259_, new_n10260_, new_n10261_, new_n10262_,
    new_n10263_, new_n10264_, new_n10265_, new_n10266_, new_n10267_,
    new_n10268_, new_n10269_, new_n10270_, new_n10271_, new_n10272_,
    new_n10273_, new_n10274_, new_n10275_, new_n10276_, new_n10277_,
    new_n10278_, new_n10279_, new_n10280_, new_n10281_, new_n10282_,
    new_n10283_, new_n10284_, new_n10285_, new_n10286_, new_n10287_,
    new_n10288_, new_n10289_, new_n10290_, new_n10291_, new_n10292_,
    new_n10293_, new_n10294_, new_n10295_, new_n10296_, new_n10297_,
    new_n10298_, new_n10299_, new_n10300_, new_n10301_, new_n10302_,
    new_n10303_, new_n10304_, new_n10305_, new_n10306_, new_n10307_,
    new_n10308_, new_n10309_, new_n10320_, new_n10321_, new_n10322_,
    new_n10323_, new_n10324_, new_n10325_, new_n10326_, new_n10327_,
    new_n10328_, new_n10329_, new_n10330_, new_n10331_, new_n10332_,
    new_n10333_, new_n10334_, new_n10335_, new_n10336_, new_n10337_,
    new_n10338_, new_n10339_, new_n10340_, new_n10341_, new_n10342_,
    new_n10343_, new_n10344_, new_n10345_, new_n10346_, new_n10347_,
    new_n10348_, new_n10349_, new_n10350_, new_n10351_, new_n10352_,
    new_n10353_, new_n10354_, new_n10355_, new_n10356_, new_n10357_,
    new_n10358_, new_n10359_, new_n10360_, new_n10361_, new_n10362_,
    new_n10363_, new_n10364_, new_n10365_, new_n10366_, new_n10367_,
    new_n10368_, new_n10369_, new_n10370_, new_n10371_, new_n10372_,
    new_n10373_, new_n10374_, new_n10375_, new_n10376_, new_n10377_,
    new_n10378_, new_n10379_, new_n10380_, new_n10381_, new_n10382_,
    new_n10383_, new_n10384_, new_n10385_, new_n10386_, new_n10387_,
    new_n10388_, new_n10389_, new_n10390_, new_n10391_, new_n10392_,
    new_n10393_, new_n10394_, new_n10395_, new_n10396_, new_n10397_,
    new_n10398_, new_n10399_, new_n10400_, new_n10401_, new_n10402_,
    new_n10403_, new_n10404_, new_n10405_, new_n10406_, new_n10407_,
    new_n10408_, new_n10409_, new_n10410_, new_n10411_, new_n10412_,
    new_n10413_, new_n10414_, new_n10415_, new_n10416_, new_n10417_,
    new_n10418_, new_n10419_, new_n10420_, new_n10421_, new_n10422_,
    new_n10423_, new_n10424_, new_n10425_, new_n10426_, new_n10427_,
    new_n10428_, new_n10429_, new_n10430_, new_n10431_, new_n10432_,
    new_n10433_, new_n10434_, new_n10435_, new_n10436_, new_n10437_,
    new_n10438_, new_n10439_, new_n10440_, new_n10441_, new_n10442_,
    new_n10443_, new_n10444_, new_n10445_, new_n10446_, new_n10447_,
    new_n10448_, new_n10449_, new_n10450_, new_n10451_, new_n10452_,
    new_n10453_, new_n10454_, new_n10455_, new_n10456_, new_n10457_,
    new_n10458_, new_n10459_, new_n10460_, new_n10461_, new_n10462_,
    new_n10463_, new_n10464_, new_n10465_, new_n10466_, new_n10467_,
    new_n10468_, new_n10469_, new_n10470_, new_n10471_, new_n10472_,
    new_n10473_, new_n10474_, new_n10475_, new_n10476_, new_n10477_,
    new_n10478_, new_n10479_, new_n10480_, new_n10481_, new_n10482_,
    new_n10483_, new_n10484_, new_n10485_, new_n10486_, new_n10487_,
    new_n10488_, new_n10489_, new_n10491_, new_n10492_, new_n10493_,
    new_n10494_, new_n10495_, new_n10496_, new_n10497_, new_n10498_,
    new_n10499_, new_n10500_, new_n10501_, new_n10502_, new_n10503_,
    new_n10504_, new_n10505_, new_n10506_, new_n10507_, new_n10508_,
    new_n10509_, new_n10510_, new_n10511_, new_n10512_, new_n10513_,
    new_n10514_, new_n10515_, new_n10516_, new_n10517_, new_n10518_,
    new_n10519_, new_n10520_, new_n10521_, new_n10522_, new_n10523_,
    new_n10524_, new_n10525_, new_n10526_, new_n10527_, new_n10528_,
    new_n10529_, new_n10530_, new_n10531_, new_n10532_, new_n10533_,
    new_n10534_, new_n10535_, new_n10536_, new_n10537_, new_n10538_,
    new_n10539_, new_n10540_, new_n10541_, new_n10542_, new_n10543_,
    new_n10544_, new_n10545_, new_n10546_, new_n10547_, new_n10548_,
    new_n10549_, new_n10550_, new_n10551_, new_n10552_, new_n10553_,
    new_n10554_, new_n10555_, new_n10556_, new_n10557_, new_n10558_,
    new_n10559_, new_n10560_, new_n10561_, new_n10562_, new_n10563_,
    new_n10564_, new_n10565_, new_n10566_, new_n10567_, new_n10568_,
    new_n10569_, new_n10570_, new_n10571_, new_n10572_, new_n10573_,
    new_n10574_, new_n10575_, new_n10576_, new_n10577_, new_n10578_,
    new_n10579_, new_n10580_, new_n10581_, new_n10582_, new_n10583_,
    new_n10584_, new_n10585_, new_n10586_, new_n10587_, new_n10588_,
    new_n10589_, new_n10590_, new_n10591_, new_n10592_, new_n10593_,
    new_n10594_, new_n10595_, new_n10596_, new_n10597_, new_n10598_,
    new_n10599_, new_n10600_, new_n10601_, new_n10602_, new_n10603_,
    new_n10604_, new_n10605_, new_n10606_, new_n10607_, new_n10608_,
    new_n10609_, new_n10610_, new_n10611_, new_n10612_, new_n10613_,
    new_n10614_, new_n10615_, new_n10616_, new_n10617_, new_n10618_,
    new_n10619_, new_n10620_, new_n10621_, new_n10622_, new_n10623_,
    new_n10624_, new_n10626_, new_n10627_, new_n10629_, new_n10631_,
    new_n10632_, new_n10633_, new_n10634_, new_n10635_, new_n10636_,
    new_n10637_, new_n10638_, new_n10639_, new_n10640_, new_n10641_,
    new_n10642_, new_n10643_, new_n10644_, new_n10645_, new_n10646_,
    new_n10647_, new_n10648_, new_n10649_, new_n10650_, new_n10651_,
    new_n10652_, new_n10653_, new_n10654_, new_n10655_, new_n10656_,
    new_n10657_, new_n10658_, new_n10659_, new_n10660_, new_n10661_,
    new_n10662_, new_n10663_, new_n10664_, new_n10665_, new_n10666_,
    new_n10667_, new_n10668_, new_n10669_, new_n10670_, new_n10671_,
    new_n10672_, new_n10673_, new_n10674_, new_n10675_, new_n10676_,
    new_n10677_, new_n10678_, new_n10679_, new_n10680_, new_n10681_,
    new_n10682_, new_n10683_, new_n10684_, new_n10685_, new_n10686_,
    new_n10687_, new_n10688_, new_n10689_, new_n10690_, new_n10691_,
    new_n10692_, new_n10693_, new_n10694_, new_n10695_, new_n10696_,
    new_n10697_, new_n10698_, new_n10699_, new_n10700_, new_n10701_,
    new_n10702_, new_n10703_, new_n10704_, new_n10705_, new_n10706_,
    new_n10707_, new_n10708_, new_n10709_, new_n10710_, new_n10711_,
    new_n10712_, new_n10713_, new_n10714_, new_n10715_, new_n10716_,
    new_n10717_, new_n10718_, new_n10719_, new_n10720_, new_n10721_,
    new_n10722_, new_n10723_, new_n10724_, new_n10725_, new_n10726_,
    new_n10727_, new_n10728_, new_n10729_, new_n10730_, new_n10731_,
    new_n10732_, new_n10733_, new_n10734_, new_n10735_, new_n10736_,
    new_n10737_, new_n10738_, new_n10739_, new_n10740_, new_n10741_,
    new_n10742_, new_n10743_, new_n10744_, new_n10745_, new_n10746_,
    new_n10747_, new_n10748_, new_n10749_, new_n10750_, new_n10751_,
    new_n10752_, new_n10753_, new_n10754_, new_n10755_, new_n10756_,
    new_n10757_, new_n10758_, new_n10759_, new_n10760_, new_n10761_,
    new_n10762_, new_n10763_, new_n10766_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10806_,
    new_n10807_, new_n10809_, new_n10810_, new_n10811_, new_n10812_,
    new_n10813_, new_n10814_, new_n10815_, new_n10816_, new_n10817_,
    new_n10818_, new_n10819_, new_n10820_, new_n10821_, new_n10822_,
    new_n10823_, new_n10824_, new_n10825_, new_n10826_, new_n10827_,
    new_n10828_, new_n10829_, new_n10830_, new_n10831_, new_n10832_,
    new_n10833_, new_n10834_, new_n10835_, new_n10836_, new_n10837_,
    new_n10838_, new_n10839_, new_n10840_, new_n10841_, new_n10842_,
    new_n10843_, new_n10844_, new_n10845_, new_n10846_, new_n10847_,
    new_n10850_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11102_, new_n11103_, new_n11104_, new_n11105_, new_n11106_,
    new_n11107_, new_n11108_, new_n11109_, new_n11110_, new_n11111_,
    new_n11112_, new_n11113_, new_n11114_, new_n11115_, new_n11116_,
    new_n11117_, new_n11118_, new_n11119_, new_n11120_, new_n11121_,
    new_n11122_, new_n11123_, new_n11124_, new_n11125_, new_n11127_,
    new_n11128_, new_n11129_, new_n11130_, new_n11131_, new_n11132_,
    new_n11133_, new_n11134_, new_n11135_, new_n11136_, new_n11137_,
    new_n11138_, new_n11139_, new_n11140_, new_n11141_, new_n11142_,
    new_n11143_, new_n11144_, new_n11145_, new_n11146_, new_n11147_,
    new_n11148_, new_n11149_, new_n11150_, new_n11151_, new_n11152_,
    new_n11153_, new_n11154_, new_n11155_, new_n11156_, new_n11157_,
    new_n11159_, new_n11160_, new_n11161_, new_n11162_, new_n11163_,
    new_n11164_, new_n11165_, new_n11166_, new_n11167_, new_n11168_,
    new_n11169_, new_n11170_, new_n11171_, new_n11172_, new_n11173_,
    new_n11174_, new_n11175_, new_n11176_, new_n11177_, new_n11178_,
    new_n11179_, new_n11180_, new_n11181_, new_n11182_, new_n11183_,
    new_n11184_, new_n11185_, new_n11186_, new_n11187_, new_n11188_,
    new_n11189_, new_n11190_, new_n11191_, new_n11192_, new_n11193_,
    new_n11194_, new_n11195_, new_n11196_, new_n11197_, new_n11198_,
    new_n11199_, new_n11200_, new_n11201_, new_n11202_, new_n11203_,
    new_n11204_, new_n11205_, new_n11206_, new_n11207_, new_n11208_,
    new_n11209_, new_n11210_, new_n11211_, new_n11212_, new_n11213_,
    new_n11214_, new_n11215_, new_n11216_, new_n11217_, new_n11218_,
    new_n11219_, new_n11220_, new_n11221_, new_n11222_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11275_, new_n11276_,
    new_n11277_, new_n11278_, new_n11279_, new_n11280_, new_n11281_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11292_, new_n11294_, new_n11295_, new_n11296_, new_n11297_,
    new_n11298_, new_n11299_, new_n11300_, new_n11301_, new_n11302_,
    new_n11303_, new_n11304_, new_n11305_, new_n11306_, new_n11307_,
    new_n11308_, new_n11309_, new_n11311_, new_n11312_, new_n11313_,
    new_n11314_, new_n11315_, new_n11316_, new_n11317_, new_n11318_,
    new_n11319_, new_n11320_, new_n11321_, new_n11322_, new_n11323_,
    new_n11324_, new_n11325_, new_n11329_, new_n11330_, new_n11331_,
    new_n11332_, new_n11333_, new_n11334_, new_n11335_, new_n11336_,
    new_n11337_, new_n11338_, new_n11339_, new_n11340_, new_n11341_,
    new_n11342_, new_n11343_, new_n11344_, new_n11345_, new_n11346_,
    new_n11347_, new_n11348_, new_n11349_, new_n11350_, new_n11351_,
    new_n11352_, new_n11353_, new_n11354_, new_n11355_, new_n11356_,
    new_n11357_, new_n11358_, new_n11359_, new_n11360_, new_n11361_,
    new_n11362_, new_n11363_, new_n11364_, new_n11365_, new_n11366_,
    new_n11367_, new_n11368_, new_n11369_, new_n11370_, new_n11371_,
    new_n11372_, new_n11373_, new_n11374_, new_n11375_, new_n11376_,
    new_n11377_, new_n11378_, new_n11379_, new_n11380_, new_n11381_,
    new_n11382_, new_n11383_, new_n11384_, new_n11385_, new_n11386_,
    new_n11387_, new_n11388_, new_n11389_, new_n11390_, new_n11391_,
    new_n11393_, new_n11394_, new_n11395_, new_n11396_, new_n11397_,
    new_n11399_, new_n11400_, new_n11401_, new_n11402_, new_n11403_,
    new_n11404_, new_n11405_, new_n11406_, new_n11407_, new_n11408_,
    new_n11409_, new_n11410_, new_n11411_, new_n11412_, new_n11413_,
    new_n11414_, new_n11415_, new_n11416_, new_n11417_, new_n11418_,
    new_n11419_, new_n11420_, new_n11421_, new_n11422_, new_n11423_,
    new_n11424_, new_n11425_, new_n11426_, new_n11427_, new_n11428_,
    new_n11429_, new_n11430_, new_n11431_, new_n11432_, new_n11433_,
    new_n11434_, new_n11435_, new_n11436_, new_n11437_, new_n11438_,
    new_n11439_, new_n11440_, new_n11441_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_,
    new_n11515_, new_n11516_, new_n11517_, new_n11518_, new_n11519_,
    new_n11520_, new_n11521_, new_n11522_, new_n11523_, new_n11524_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11556_,
    new_n11557_, new_n11558_, new_n11559_, new_n11560_, new_n11561_,
    new_n11562_, new_n11563_, new_n11564_, new_n11565_, new_n11567_,
    new_n11568_, new_n11569_, new_n11570_, new_n11571_, new_n11572_,
    new_n11573_, new_n11574_, new_n11575_, new_n11576_, new_n11577_,
    new_n11578_, new_n11579_, new_n11580_, new_n11581_, new_n11582_,
    new_n11583_, new_n11584_, new_n11587_, new_n11588_, new_n11589_,
    new_n11590_, new_n11591_, new_n11592_, new_n11593_, new_n11594_,
    new_n11595_, new_n11596_, new_n11597_, new_n11598_, new_n11599_,
    new_n11600_, new_n11601_, new_n11602_, new_n11603_, new_n11604_,
    new_n11605_, new_n11606_, new_n11607_, new_n11608_, new_n11609_,
    new_n11610_, new_n11611_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11667_, new_n11668_, new_n11669_, new_n11670_, new_n11671_,
    new_n11672_, new_n11673_, new_n11674_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11703_, new_n11704_, new_n11705_, new_n11716_, new_n11717_,
    new_n11718_, new_n11721_, new_n11722_, new_n11723_, new_n11724_,
    new_n11725_, new_n11726_, new_n11727_, new_n11728_, new_n11729_,
    new_n11730_, new_n11731_, new_n11732_, new_n11733_, new_n11734_,
    new_n11735_, new_n11736_, new_n11737_, new_n11738_, new_n11739_,
    new_n11740_, new_n11741_, new_n11742_, new_n11743_, new_n11744_,
    new_n11745_, new_n11747_, new_n11748_, new_n11749_, new_n11750_,
    new_n11751_, new_n11752_, new_n11753_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11762_, new_n11766_, new_n11767_, new_n11768_, new_n11769_,
    new_n11770_, new_n11771_, new_n11772_, new_n11773_, new_n11774_,
    new_n11775_, new_n11776_, new_n11777_, new_n11778_, new_n11779_,
    new_n11780_, new_n11781_, new_n11782_, new_n11783_, new_n11784_,
    new_n11785_, new_n11786_, new_n11787_, new_n11788_, new_n11789_,
    new_n11790_, new_n11791_, new_n11792_, new_n11793_, new_n11794_,
    new_n11795_, new_n11796_, new_n11797_, new_n11798_, new_n11799_,
    new_n11800_, new_n11801_, new_n11802_, new_n11803_, new_n11804_,
    new_n11805_, new_n11806_, new_n11807_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11826_,
    new_n11829_, new_n11830_, new_n11831_, new_n11832_, new_n11833_,
    new_n11834_, new_n11835_, new_n11836_, new_n11837_, new_n11838_,
    new_n11839_, new_n11840_, new_n11841_, new_n11842_, new_n11843_,
    new_n11844_, new_n11845_, new_n11846_, new_n11847_, new_n11848_,
    new_n11849_, new_n11850_, new_n11851_, new_n11852_, new_n11853_,
    new_n11854_, new_n11855_, new_n11856_, new_n11857_, new_n11858_,
    new_n11859_, new_n11860_, new_n11861_, new_n11862_, new_n11863_,
    new_n11864_, new_n11865_, new_n11867_, new_n11868_, new_n11869_,
    new_n11870_, new_n11871_, new_n11872_, new_n11873_, new_n11874_,
    new_n11875_, new_n11876_, new_n11877_, new_n11878_, new_n11879_,
    new_n11880_, new_n11881_, new_n11882_, new_n11883_, new_n11884_,
    new_n11885_, new_n11886_, new_n11887_, new_n11888_, new_n11889_,
    new_n11890_, new_n11891_, new_n11892_, new_n11893_, new_n11894_,
    new_n11895_, new_n11896_, new_n11897_, new_n11898_, new_n11899_,
    new_n11900_, new_n11901_, new_n11902_, new_n11903_, new_n11904_,
    new_n11905_, new_n11906_, new_n11907_, new_n11908_, new_n11909_,
    new_n11910_, new_n11911_, new_n11912_, new_n11913_, new_n11914_,
    new_n11915_, new_n11916_, new_n11917_, new_n11918_, new_n11919_,
    new_n11920_, new_n11921_, new_n11922_, new_n11923_, new_n11924_,
    new_n11925_, new_n11926_, new_n11927_, new_n11928_, new_n11929_,
    new_n11930_, new_n11931_, new_n11932_, new_n11933_, new_n11934_,
    new_n11935_, new_n11936_, new_n11937_, new_n11938_, new_n11939_,
    new_n11940_, new_n11941_, new_n11942_, new_n11943_, new_n11944_,
    new_n11945_, new_n11946_, new_n11947_, new_n11948_, new_n11949_,
    new_n11950_, new_n11951_, new_n11952_, new_n11953_, new_n11954_,
    new_n11955_, new_n11956_, new_n11957_, new_n11958_, new_n11959_,
    new_n11960_, new_n11961_, new_n11962_, new_n11963_, new_n11964_,
    new_n11965_, new_n11966_, new_n11967_, new_n11968_, new_n11969_,
    new_n11970_, new_n11971_, new_n11972_, new_n11973_, new_n11974_,
    new_n11975_, new_n11976_, new_n11977_, new_n11978_, new_n11979_,
    new_n11980_, new_n11981_, new_n11982_, new_n11983_, new_n11984_,
    new_n11985_, new_n11986_, new_n11987_, new_n11988_, new_n11989_,
    new_n11990_, new_n11991_, new_n11992_, new_n11993_, new_n11994_,
    new_n11995_, new_n11996_, new_n11997_, new_n11998_, new_n11999_,
    new_n12000_, new_n12001_, new_n12002_, new_n12003_, new_n12004_,
    new_n12005_, new_n12006_, new_n12007_, new_n12008_, new_n12009_,
    new_n12010_, new_n12011_, new_n12012_, new_n12013_, new_n12014_,
    new_n12015_, new_n12016_, new_n12017_, new_n12018_, new_n12019_,
    new_n12020_, new_n12021_, new_n12022_, new_n12023_, new_n12024_,
    new_n12025_, new_n12026_, new_n12027_, new_n12028_, new_n12029_,
    new_n12030_, new_n12031_, new_n12032_, new_n12033_, new_n12034_,
    new_n12035_, new_n12036_, new_n12037_, new_n12038_, new_n12039_,
    new_n12040_, new_n12041_, new_n12042_, new_n12043_, new_n12044_,
    new_n12045_, new_n12046_, new_n12047_, new_n12048_, new_n12049_,
    new_n12050_, new_n12051_, new_n12052_, new_n12053_, new_n12054_,
    new_n12055_, new_n12056_, new_n12057_, new_n12058_, new_n12059_,
    new_n12060_, new_n12061_, new_n12062_, new_n12063_, new_n12064_,
    new_n12065_, new_n12066_, new_n12067_, new_n12068_, new_n12069_,
    new_n12070_, new_n12071_, new_n12072_, new_n12073_, new_n12074_,
    new_n12075_, new_n12076_, new_n12077_, new_n12078_, new_n12079_,
    new_n12080_, new_n12081_, new_n12082_, new_n12083_, new_n12084_,
    new_n12085_, new_n12086_, new_n12087_, new_n12088_, new_n12089_,
    new_n12090_, new_n12091_, new_n12092_, new_n12093_, new_n12094_,
    new_n12095_, new_n12096_, new_n12097_, new_n12098_, new_n12099_,
    new_n12100_, new_n12101_, new_n12102_, new_n12103_, new_n12104_,
    new_n12105_, new_n12106_, new_n12107_, new_n12108_, new_n12109_,
    new_n12110_, new_n12111_, new_n12112_, new_n12113_, new_n12114_,
    new_n12115_, new_n12116_, new_n12117_, new_n12118_, new_n12119_,
    new_n12120_, new_n12121_, new_n12122_, new_n12123_, new_n12124_,
    new_n12125_, new_n12126_, new_n12127_, new_n12128_, new_n12129_,
    new_n12130_, new_n12131_, new_n12132_, new_n12133_, new_n12134_,
    new_n12135_, new_n12136_, new_n12137_, new_n12138_, new_n12139_,
    new_n12140_, new_n12141_, new_n12142_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12156_, new_n12157_, new_n12158_, new_n12159_,
    new_n12160_, new_n12161_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12171_, new_n12172_, new_n12173_, new_n12174_,
    new_n12175_, new_n12176_, new_n12177_, new_n12178_, new_n12179_,
    new_n12180_, new_n12181_, new_n12182_, new_n12183_, new_n12184_,
    new_n12185_, new_n12186_, new_n12187_, new_n12188_, new_n12189_,
    new_n12190_, new_n12191_, new_n12192_, new_n12193_, new_n12194_,
    new_n12195_, new_n12196_, new_n12197_, new_n12198_, new_n12199_,
    new_n12200_, new_n12201_, new_n12202_, new_n12203_, new_n12204_,
    new_n12205_, new_n12206_, new_n12207_, new_n12208_, new_n12209_,
    new_n12210_, new_n12211_, new_n12212_, new_n12213_, new_n12214_,
    new_n12215_, new_n12216_, new_n12217_, new_n12218_, new_n12219_,
    new_n12220_, new_n12221_, new_n12222_, new_n12223_, new_n12224_,
    new_n12225_, new_n12226_, new_n12227_, new_n12228_, new_n12229_,
    new_n12230_, new_n12231_, new_n12232_, new_n12233_, new_n12234_,
    new_n12235_, new_n12236_, new_n12237_, new_n12238_, new_n12239_,
    new_n12240_, new_n12241_, new_n12242_, new_n12243_, new_n12244_,
    new_n12245_, new_n12246_, new_n12247_, new_n12248_, new_n12249_,
    new_n12250_, new_n12251_, new_n12252_, new_n12253_, new_n12254_,
    new_n12255_, new_n12256_, new_n12257_, new_n12258_, new_n12259_,
    new_n12260_, new_n12261_, new_n12262_, new_n12263_, new_n12264_,
    new_n12265_, new_n12266_, new_n12267_, new_n12268_, new_n12269_,
    new_n12270_, new_n12271_, new_n12272_, new_n12273_, new_n12274_,
    new_n12275_, new_n12276_, new_n12277_, new_n12278_, new_n12279_,
    new_n12280_, new_n12281_, new_n12282_, new_n12283_, new_n12284_,
    new_n12285_, new_n12286_, new_n12287_, new_n12288_, new_n12289_,
    new_n12290_, new_n12291_, new_n12292_, new_n12293_, new_n12294_,
    new_n12295_, new_n12296_, new_n12297_, new_n12298_, new_n12299_,
    new_n12300_, new_n12301_, new_n12302_, new_n12303_, new_n12304_,
    new_n12305_, new_n12306_, new_n12307_, new_n12308_, new_n12309_,
    new_n12310_, new_n12311_, new_n12312_, new_n12313_, new_n12314_,
    new_n12315_, new_n12316_, new_n12317_, new_n12318_, new_n12319_,
    new_n12320_, new_n12321_, new_n12322_, new_n12323_, new_n12324_,
    new_n12325_, new_n12326_, new_n12327_, new_n12328_, new_n12329_,
    new_n12330_, new_n12331_, new_n12332_, new_n12333_, new_n12334_,
    new_n12335_, new_n12336_, new_n12337_, new_n12338_, new_n12339_,
    new_n12340_, new_n12341_, new_n12342_, new_n12343_, new_n12344_,
    new_n12345_, new_n12346_, new_n12347_, new_n12348_, new_n12349_,
    new_n12350_, new_n12351_, new_n12352_, new_n12353_, new_n12354_,
    new_n12355_, new_n12356_, new_n12357_, new_n12358_, new_n12359_,
    new_n12360_, new_n12361_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12379_,
    new_n12380_, new_n12381_, new_n12382_, new_n12383_, new_n12384_,
    new_n12385_, new_n12386_, new_n12387_, new_n12388_, new_n12389_,
    new_n12390_, new_n12391_, new_n12392_, new_n12393_, new_n12394_,
    new_n12395_, new_n12396_, new_n12397_, new_n12398_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12438_, new_n12439_,
    new_n12440_, new_n12441_, new_n12442_, new_n12443_, new_n12444_,
    new_n12445_, new_n12446_, new_n12447_, new_n12448_, new_n12449_,
    new_n12450_, new_n12451_, new_n12452_, new_n12453_, new_n12454_,
    new_n12455_, new_n12456_, new_n12457_, new_n12458_, new_n12459_,
    new_n12460_, new_n12461_, new_n12462_, new_n12463_, new_n12464_,
    new_n12465_, new_n12466_, new_n12467_, new_n12468_, new_n12469_,
    new_n12470_, new_n12471_, new_n12472_, new_n12473_, new_n12474_,
    new_n12475_, new_n12476_, new_n12477_, new_n12478_, new_n12479_,
    new_n12480_, new_n12481_, new_n12482_, new_n12483_, new_n12484_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12491_, new_n12492_, new_n12493_, new_n12494_,
    new_n12495_, new_n12496_, new_n12497_, new_n12498_, new_n12499_,
    new_n12500_, new_n12501_, new_n12502_, new_n12503_, new_n12504_,
    new_n12505_, new_n12506_, new_n12507_, new_n12508_, new_n12509_,
    new_n12510_, new_n12511_, new_n12512_, new_n12513_, new_n12514_,
    new_n12515_, new_n12516_, new_n12517_, new_n12518_, new_n12519_,
    new_n12520_, new_n12521_, new_n12522_, new_n12523_, new_n12524_,
    new_n12525_, new_n12526_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12532_, new_n12533_, new_n12534_,
    new_n12535_, new_n12536_, new_n12537_, new_n12538_, new_n12539_,
    new_n12540_, new_n12541_, new_n12542_, new_n12543_, new_n12544_,
    new_n12545_, new_n12546_, new_n12547_, new_n12548_, new_n12549_,
    new_n12550_, new_n12551_, new_n12552_, new_n12553_, new_n12554_,
    new_n12555_, new_n12556_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12806_,
    new_n12807_, new_n12808_, new_n12809_, new_n12810_, new_n12811_,
    new_n12812_, new_n12813_, new_n12814_, new_n12815_, new_n12816_,
    new_n12817_, new_n12818_, new_n12819_, new_n12820_, new_n12821_,
    new_n12822_, new_n12823_, new_n12824_, new_n12825_, new_n12826_,
    new_n12827_, new_n12828_, new_n12829_, new_n12830_, new_n12831_,
    new_n12832_, new_n12833_, new_n12834_, new_n12835_, new_n12836_,
    new_n12837_, new_n12838_, new_n12839_, new_n12840_, new_n12841_,
    new_n12842_, new_n12843_, new_n12844_, new_n12845_, new_n12846_,
    new_n12847_, new_n12848_, new_n12849_, new_n12850_, new_n12851_,
    new_n12852_, new_n12853_, new_n12854_, new_n12855_, new_n12856_,
    new_n12857_, new_n12858_, new_n12859_, new_n12860_, new_n12861_,
    new_n12862_, new_n12863_, new_n12864_, new_n12865_, new_n12866_,
    new_n12867_, new_n12868_, new_n12869_, new_n12870_, new_n12871_,
    new_n12872_, new_n12873_, new_n12874_, new_n12875_, new_n12876_,
    new_n12877_, new_n12878_, new_n12879_, new_n12880_, new_n12881_,
    new_n12882_, new_n12883_, new_n12884_, new_n12885_, new_n12886_,
    new_n12887_, new_n12888_, new_n12889_, new_n12890_, new_n12891_,
    new_n12892_, new_n12893_, new_n12894_, new_n12895_, new_n12896_,
    new_n12897_, new_n12898_, new_n12899_, new_n12900_, new_n12901_,
    new_n12902_, new_n12903_, new_n12904_, new_n12905_, new_n12906_,
    new_n12907_, new_n12908_, new_n12909_, new_n12910_, new_n12911_,
    new_n12912_, new_n12913_, new_n12914_, new_n12915_, new_n12916_,
    new_n12917_, new_n12918_, new_n12919_, new_n12920_, new_n12921_,
    new_n12922_, new_n12923_, new_n12924_, new_n12925_, new_n12926_,
    new_n12927_, new_n12928_, new_n12929_, new_n12930_, new_n12931_,
    new_n12932_, new_n12933_, new_n12934_, new_n12935_, new_n12936_,
    new_n12937_, new_n12938_, new_n12939_, new_n12940_, new_n12941_,
    new_n12942_, new_n12943_, new_n12944_, new_n12945_, new_n12946_,
    new_n12947_, new_n12948_, new_n12949_, new_n12950_, new_n12951_,
    new_n12952_, new_n12953_, new_n12954_, new_n12955_, new_n12956_,
    new_n12957_, new_n12959_, new_n12960_, new_n12961_, new_n12962_,
    new_n12963_, new_n12964_, new_n12965_, new_n12966_, new_n12967_,
    new_n12968_, new_n12969_, new_n12970_, new_n12971_, new_n12972_,
    new_n12973_, new_n12974_, new_n12975_, new_n12976_, new_n12977_,
    new_n12978_, new_n12979_, new_n12980_, new_n12981_, new_n12982_,
    new_n12983_, new_n12984_, new_n12985_, new_n12986_, new_n12987_,
    new_n12988_, new_n12989_, new_n12990_, new_n12991_, new_n12992_,
    new_n12993_, new_n12994_, new_n12995_, new_n12996_, new_n12997_,
    new_n12998_, new_n12999_, new_n13000_, new_n13001_, new_n13002_,
    new_n13003_, new_n13004_, new_n13005_, new_n13006_, new_n13007_,
    new_n13008_, new_n13009_, new_n13010_, new_n13011_, new_n13012_,
    new_n13013_, new_n13014_, new_n13015_, new_n13016_, new_n13017_,
    new_n13018_, new_n13019_, new_n13020_, new_n13021_, new_n13022_,
    new_n13023_, new_n13024_, new_n13025_, new_n13026_, new_n13027_,
    new_n13028_, new_n13029_, new_n13030_, new_n13031_, new_n13032_,
    new_n13033_, new_n13034_, new_n13035_, new_n13036_, new_n13037_,
    new_n13038_, new_n13039_, new_n13040_, new_n13041_, new_n13042_,
    new_n13043_, new_n13044_, new_n13045_, new_n13046_, new_n13047_,
    new_n13048_, new_n13049_, new_n13050_, new_n13051_, new_n13052_,
    new_n13053_, new_n13054_, new_n13055_, new_n13056_, new_n13057_,
    new_n13058_, new_n13059_, new_n13060_, new_n13061_, new_n13062_,
    new_n13063_, new_n13064_, new_n13065_, new_n13066_, new_n13067_,
    new_n13068_, new_n13069_, new_n13070_, new_n13071_, new_n13072_,
    new_n13073_, new_n13074_, new_n13075_, new_n13076_, new_n13077_,
    new_n13078_, new_n13079_, new_n13080_, new_n13081_, new_n13082_,
    new_n13083_, new_n13084_, new_n13085_, new_n13086_, new_n13087_,
    new_n13088_, new_n13089_, new_n13090_, new_n13091_, new_n13092_,
    new_n13093_, new_n13094_, new_n13095_, new_n13096_, new_n13097_,
    new_n13098_, new_n13099_, new_n13100_, new_n13101_, new_n13102_,
    new_n13103_, new_n13104_, new_n13105_, new_n13106_, new_n13107_,
    new_n13108_, new_n13109_, new_n13110_, new_n13111_, new_n13112_,
    new_n13113_, new_n13114_, new_n13115_, new_n13116_, new_n13117_,
    new_n13118_, new_n13119_, new_n13120_, new_n13121_, new_n13122_,
    new_n13123_, new_n13124_, new_n13125_, new_n13126_, new_n13127_,
    new_n13128_, new_n13129_, new_n13130_, new_n13131_, new_n13132_,
    new_n13133_, new_n13134_, new_n13135_, new_n13136_, new_n13137_,
    new_n13138_, new_n13139_, new_n13140_, new_n13141_, new_n13142_,
    new_n13143_, new_n13144_, new_n13145_, new_n13146_, new_n13147_,
    new_n13148_, new_n13149_, new_n13150_, new_n13151_, new_n13152_,
    new_n13153_, new_n13154_, new_n13155_, new_n13156_, new_n13157_,
    new_n13158_, new_n13159_, new_n13160_, new_n13161_, new_n13162_,
    new_n13163_, new_n13164_, new_n13165_, new_n13166_, new_n13167_,
    new_n13168_, new_n13169_, new_n13170_, new_n13171_, new_n13172_,
    new_n13173_, new_n13174_, new_n13175_, new_n13176_, new_n13177_,
    new_n13178_, new_n13179_, new_n13180_, new_n13181_, new_n13182_,
    new_n13183_, new_n13184_, new_n13185_, new_n13186_, new_n13187_,
    new_n13189_, new_n13190_, new_n13191_, new_n13192_, new_n13193_,
    new_n13194_, new_n13195_, new_n13196_, new_n13197_, new_n13198_,
    new_n13199_, new_n13200_, new_n13201_, new_n13202_, new_n13203_,
    new_n13204_, new_n13205_, new_n13206_, new_n13207_, new_n13208_,
    new_n13209_, new_n13210_, new_n13211_, new_n13212_, new_n13213_,
    new_n13214_, new_n13215_, new_n13216_, new_n13217_, new_n13218_,
    new_n13219_, new_n13220_, new_n13221_, new_n13222_, new_n13223_,
    new_n13224_, new_n13225_, new_n13226_, new_n13227_, new_n13228_,
    new_n13229_, new_n13230_, new_n13231_, new_n13232_, new_n13233_,
    new_n13234_, new_n13235_, new_n13236_, new_n13237_, new_n13238_,
    new_n13239_, new_n13240_, new_n13241_, new_n13242_, new_n13243_,
    new_n13244_, new_n13245_, new_n13246_, new_n13247_, new_n13248_,
    new_n13249_, new_n13250_, new_n13251_, new_n13252_, new_n13253_,
    new_n13254_, new_n13255_, new_n13256_, new_n13257_, new_n13258_,
    new_n13259_, new_n13260_, new_n13261_, new_n13262_, new_n13263_,
    new_n13264_, new_n13265_, new_n13266_, new_n13267_, new_n13268_,
    new_n13269_, new_n13270_, new_n13271_, new_n13272_, new_n13273_,
    new_n13274_, new_n13275_, new_n13276_, new_n13277_, new_n13278_,
    new_n13279_, new_n13280_, new_n13281_, new_n13282_, new_n13283_,
    new_n13284_, new_n13285_, new_n13286_, new_n13287_, new_n13288_,
    new_n13289_, new_n13290_, new_n13291_, new_n13292_, new_n13293_,
    new_n13294_, new_n13295_, new_n13296_, new_n13297_, new_n13298_,
    new_n13299_, new_n13300_, new_n13301_, new_n13302_, new_n13303_,
    new_n13304_, new_n13305_, new_n13306_, new_n13307_, new_n13308_,
    new_n13309_, new_n13310_, new_n13311_, new_n13312_, new_n13313_,
    new_n13314_, new_n13315_, new_n13316_, new_n13317_, new_n13318_,
    new_n13319_, new_n13320_, new_n13321_, new_n13322_, new_n13323_,
    new_n13324_, new_n13325_, new_n13326_, new_n13327_, new_n13328_,
    new_n13329_, new_n13330_, new_n13331_, new_n13332_, new_n13333_,
    new_n13334_, new_n13335_, new_n13336_, new_n13337_, new_n13338_,
    new_n13339_, new_n13340_, new_n13341_, new_n13342_, new_n13343_,
    new_n13344_, new_n13345_, new_n13346_, new_n13347_, new_n13348_,
    new_n13349_, new_n13350_, new_n13351_, new_n13352_, new_n13353_,
    new_n13354_, new_n13355_, new_n13356_, new_n13357_, new_n13358_,
    new_n13359_, new_n13360_, new_n13361_, new_n13362_, new_n13363_,
    new_n13364_, new_n13365_, new_n13366_, new_n13367_, new_n13368_,
    new_n13369_, new_n13370_, new_n13371_, new_n13372_, new_n13373_,
    new_n13374_, new_n13375_, new_n13376_, new_n13377_, new_n13378_,
    new_n13379_, new_n13380_, new_n13381_, new_n13382_, new_n13383_,
    new_n13384_, new_n13385_, new_n13386_, new_n13387_, new_n13388_,
    new_n13389_, new_n13390_, new_n13391_, new_n13392_, new_n13393_,
    new_n13394_, new_n13395_, new_n13396_, new_n13397_, new_n13398_,
    new_n13399_, new_n13400_, new_n13401_, new_n13402_, new_n13403_,
    new_n13404_, new_n13405_, new_n13406_, new_n13407_, new_n13408_,
    new_n13409_, new_n13410_, new_n13411_, new_n13412_, new_n13413_,
    new_n13414_, new_n13415_, new_n13416_, new_n13417_, new_n13418_,
    new_n13419_, new_n13420_, new_n13421_, new_n13422_, new_n13423_,
    new_n13424_, new_n13425_, new_n13426_, new_n13427_, new_n13428_,
    new_n13429_, new_n13430_, new_n13431_, new_n13432_, new_n13433_,
    new_n13434_, new_n13435_, new_n13436_, new_n13437_, new_n13438_,
    new_n13439_, new_n13440_, new_n13441_, new_n13442_, new_n13443_,
    new_n13444_, new_n13445_, new_n13446_, new_n13447_, new_n13448_,
    new_n13449_, new_n13450_, new_n13451_, new_n13452_, new_n13453_,
    new_n13454_, new_n13455_, new_n13456_, new_n13457_, new_n13458_,
    new_n13459_, new_n13460_, new_n13461_, new_n13462_, new_n13463_,
    new_n13464_, new_n13465_, new_n13466_, new_n13467_, new_n13468_,
    new_n13469_, new_n13470_, new_n13471_, new_n13472_, new_n13473_,
    new_n13474_, new_n13475_, new_n13476_, new_n13477_, new_n13478_,
    new_n13479_, new_n13480_, new_n13481_, new_n13482_, new_n13483_,
    new_n13484_, new_n13485_, new_n13486_, new_n13487_, new_n13488_,
    new_n13489_, new_n13490_, new_n13491_, new_n13492_, new_n13493_,
    new_n13494_, new_n13495_, new_n13496_, new_n13497_, new_n13498_,
    new_n13499_, new_n13500_, new_n13501_, new_n13502_, new_n13503_,
    new_n13504_, new_n13505_, new_n13506_, new_n13507_, new_n13508_,
    new_n13509_, new_n13510_, new_n13511_, new_n13512_, new_n13513_,
    new_n13514_, new_n13515_, new_n13516_, new_n13517_, new_n13518_,
    new_n13519_, new_n13520_, new_n13521_, new_n13522_, new_n13523_,
    new_n13524_, new_n13525_, new_n13526_, new_n13527_, new_n13528_,
    new_n13529_, new_n13530_, new_n13531_, new_n13532_, new_n13533_,
    new_n13534_, new_n13535_, new_n13536_, new_n13537_, new_n13538_,
    new_n13539_, new_n13540_, new_n13541_, new_n13542_, new_n13543_,
    new_n13544_, new_n13545_, new_n13546_, new_n13547_, new_n13548_,
    new_n13549_, new_n13550_, new_n13551_, new_n13552_, new_n13553_,
    new_n13554_, new_n13555_, new_n13556_, new_n13557_, new_n13558_,
    new_n13559_, new_n13560_, new_n13561_, new_n13562_, new_n13563_,
    new_n13564_, new_n13565_, new_n13566_, new_n13567_, new_n13568_,
    new_n13569_, new_n13570_, new_n13571_, new_n13572_, new_n13573_,
    new_n13574_, new_n13575_, new_n13576_, new_n13577_, new_n13578_,
    new_n13579_, new_n13580_, new_n13581_, new_n13582_, new_n13583_,
    new_n13584_, new_n13585_, new_n13586_, new_n13587_, new_n13588_,
    new_n13589_, new_n13590_, new_n13591_, new_n13592_, new_n13593_,
    new_n13594_, new_n13595_, new_n13596_, new_n13597_, new_n13598_,
    new_n13599_, new_n13600_, new_n13601_, new_n13602_, new_n13603_,
    new_n13604_, new_n13605_, new_n13606_, new_n13607_, new_n13608_,
    new_n13609_, new_n13610_, new_n13611_, new_n13612_, new_n13613_,
    new_n13615_, new_n13616_, new_n13617_, new_n13618_, new_n13619_,
    new_n13620_, new_n13621_, new_n13622_, new_n13623_, new_n13624_,
    new_n13625_, new_n13626_, new_n13627_, new_n13628_, new_n13629_,
    new_n13630_, new_n13631_, new_n13632_, new_n13633_, new_n13634_,
    new_n13635_, new_n13636_, new_n13637_, new_n13638_, new_n13639_,
    new_n13640_, new_n13641_, new_n13642_, new_n13643_, new_n13644_,
    new_n13645_, new_n13646_, new_n13647_, new_n13648_, new_n13649_,
    new_n13650_, new_n13651_, new_n13652_, new_n13653_, new_n13654_,
    new_n13655_, new_n13656_, new_n13657_, new_n13658_, new_n13659_,
    new_n13660_, new_n13661_, new_n13662_, new_n13663_, new_n13664_,
    new_n13665_, new_n13666_, new_n13667_, new_n13668_, new_n13669_,
    new_n13670_, new_n13671_, new_n13672_, new_n13673_, new_n13674_,
    new_n13675_, new_n13676_, new_n13677_, new_n13678_, new_n13679_,
    new_n13680_, new_n13681_, new_n13682_, new_n13683_, new_n13684_,
    new_n13685_, new_n13686_, new_n13687_, new_n13688_, new_n13689_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13750_,
    new_n13751_, new_n13752_, new_n13753_, new_n13754_, new_n13755_,
    new_n13756_, new_n13757_, new_n13758_, new_n13759_, new_n13760_,
    new_n13761_, new_n13762_, new_n13763_, new_n13764_, new_n13765_,
    new_n13766_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13831_,
    new_n13832_, new_n13833_, new_n13834_, new_n13835_, new_n13836_,
    new_n13837_, new_n13838_, new_n13839_, new_n13840_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13848_, new_n13849_, new_n13850_, new_n13851_,
    new_n13852_, new_n13853_, new_n13854_, new_n13855_, new_n13856_,
    new_n13857_, new_n13858_, new_n13859_, new_n13860_, new_n13861_,
    new_n13862_, new_n13863_, new_n13864_, new_n13865_, new_n13866_,
    new_n13867_, new_n13868_, new_n13869_, new_n13870_, new_n13871_,
    new_n13872_, new_n13873_, new_n13874_, new_n13875_, new_n13876_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13883_, new_n13884_, new_n13885_, new_n13886_,
    new_n13887_, new_n13888_, new_n13889_, new_n13890_, new_n13891_,
    new_n13892_, new_n13893_, new_n13894_, new_n13895_, new_n13896_,
    new_n13897_, new_n13898_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13952_,
    new_n13953_, new_n13954_, new_n13955_, new_n13956_, new_n13957_,
    new_n13958_, new_n13959_, new_n13960_, new_n13961_, new_n13962_,
    new_n13963_, new_n13964_, new_n13965_, new_n13966_, new_n13967_,
    new_n13968_, new_n13969_, new_n13970_, new_n13971_, new_n13972_,
    new_n13973_, new_n13974_, new_n13975_, new_n13976_, new_n13977_,
    new_n13978_, new_n13979_, new_n13980_, new_n13981_, new_n13982_,
    new_n13983_, new_n13984_, new_n13985_, new_n13986_, new_n13987_,
    new_n13988_, new_n13989_, new_n13990_, new_n13991_, new_n13992_,
    new_n13993_, new_n13994_, new_n13995_, new_n13996_, new_n13997_,
    new_n13998_, new_n13999_, new_n14000_, new_n14001_, new_n14002_,
    new_n14003_, new_n14004_, new_n14005_, new_n14006_, new_n14007_,
    new_n14008_, new_n14009_, new_n14010_, new_n14011_, new_n14012_,
    new_n14013_, new_n14014_, new_n14015_, new_n14016_, new_n14017_,
    new_n14018_, new_n14019_, new_n14020_, new_n14021_, new_n14022_,
    new_n14023_, new_n14024_, new_n14025_, new_n14026_, new_n14027_,
    new_n14028_, new_n14029_, new_n14030_, new_n14031_, new_n14032_,
    new_n14033_, new_n14034_, new_n14035_, new_n14036_, new_n14037_,
    new_n14038_, new_n14039_, new_n14040_, new_n14041_, new_n14042_,
    new_n14043_, new_n14044_, new_n14045_, new_n14046_, new_n14047_,
    new_n14048_, new_n14049_, new_n14050_, new_n14051_, new_n14052_,
    new_n14053_, new_n14054_, new_n14055_, new_n14056_, new_n14057_,
    new_n14058_, new_n14059_, new_n14060_, new_n14061_, new_n14062_,
    new_n14063_, new_n14064_, new_n14065_, new_n14066_, new_n14067_,
    new_n14068_, new_n14069_, new_n14070_, new_n14071_, new_n14072_,
    new_n14073_, new_n14074_, new_n14075_, new_n14076_, new_n14077_,
    new_n14078_, new_n14079_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14084_, new_n14085_, new_n14086_, new_n14087_,
    new_n14088_, new_n14089_, new_n14090_, new_n14091_, new_n14092_,
    new_n14093_, new_n14094_, new_n14095_, new_n14096_, new_n14097_,
    new_n14098_, new_n14099_, new_n14100_, new_n14101_, new_n14102_,
    new_n14103_, new_n14104_, new_n14105_, new_n14106_, new_n14107_,
    new_n14108_, new_n14109_, new_n14110_, new_n14111_, new_n14112_,
    new_n14113_, new_n14114_, new_n14115_, new_n14116_, new_n14117_,
    new_n14118_, new_n14119_, new_n14120_, new_n14121_, new_n14122_,
    new_n14123_, new_n14124_, new_n14125_, new_n14126_, new_n14127_,
    new_n14128_, new_n14129_, new_n14130_, new_n14131_, new_n14132_,
    new_n14133_, new_n14134_, new_n14135_, new_n14136_, new_n14137_,
    new_n14138_, new_n14139_, new_n14140_, new_n14141_, new_n14142_,
    new_n14143_, new_n14144_, new_n14145_, new_n14146_, new_n14147_,
    new_n14148_, new_n14149_, new_n14150_, new_n14151_, new_n14152_,
    new_n14153_, new_n14154_, new_n14155_, new_n14156_, new_n14157_,
    new_n14158_, new_n14159_, new_n14160_, new_n14161_, new_n14162_,
    new_n14163_, new_n14164_, new_n14165_, new_n14166_, new_n14167_,
    new_n14168_, new_n14169_, new_n14170_, new_n14171_, new_n14172_,
    new_n14173_, new_n14174_, new_n14175_, new_n14176_, new_n14177_,
    new_n14178_, new_n14179_, new_n14180_, new_n14181_, new_n14182_,
    new_n14183_, new_n14184_, new_n14185_, new_n14186_, new_n14187_,
    new_n14188_, new_n14189_, new_n14190_, new_n14191_, new_n14192_,
    new_n14193_, new_n14194_, new_n14195_, new_n14196_, new_n14197_,
    new_n14198_, new_n14199_, new_n14200_, new_n14201_, new_n14202_,
    new_n14203_, new_n14204_, new_n14205_, new_n14207_, new_n14208_,
    new_n14209_, new_n14210_, new_n14211_, new_n14212_, new_n14213_,
    new_n14214_, new_n14215_, new_n14216_, new_n14217_, new_n14218_,
    new_n14219_, new_n14220_, new_n14221_, new_n14222_, new_n14223_,
    new_n14224_, new_n14225_, new_n14226_, new_n14227_, new_n14228_,
    new_n14229_, new_n14230_, new_n14231_, new_n14232_, new_n14233_,
    new_n14234_, new_n14235_, new_n14236_, new_n14237_, new_n14238_,
    new_n14239_, new_n14240_, new_n14241_, new_n14242_, new_n14243_,
    new_n14244_, new_n14245_, new_n14246_, new_n14247_, new_n14248_,
    new_n14249_, new_n14250_, new_n14251_, new_n14252_, new_n14253_,
    new_n14254_, new_n14255_, new_n14256_, new_n14257_, new_n14258_,
    new_n14259_, new_n14260_, new_n14261_, new_n14262_, new_n14263_,
    new_n14264_, new_n14265_, new_n14266_, new_n14267_, new_n14268_,
    new_n14269_, new_n14270_, new_n14271_, new_n14272_, new_n14273_,
    new_n14274_, new_n14275_, new_n14276_, new_n14277_, new_n14278_,
    new_n14279_, new_n14280_, new_n14281_, new_n14282_, new_n14283_,
    new_n14284_, new_n14285_, new_n14286_, new_n14287_, new_n14288_,
    new_n14289_, new_n14290_, new_n14291_, new_n14292_, new_n14293_,
    new_n14294_, new_n14295_, new_n14296_, new_n14297_, new_n14298_,
    new_n14299_, new_n14300_, new_n14301_, new_n14302_, new_n14303_,
    new_n14304_, new_n14305_, new_n14306_, new_n14307_, new_n14308_,
    new_n14309_, new_n14310_, new_n14311_, new_n14312_, new_n14313_,
    new_n14314_, new_n14315_, new_n14316_, new_n14317_, new_n14318_,
    new_n14319_, new_n14320_, new_n14321_, new_n14322_, new_n14323_,
    new_n14324_, new_n14325_, new_n14326_, new_n14327_, new_n14328_,
    new_n14329_, new_n14330_, new_n14331_, new_n14332_, new_n14333_,
    new_n14334_, new_n14335_, new_n14336_, new_n14337_, new_n14338_,
    new_n14339_, new_n14340_, new_n14341_, new_n14342_, new_n14343_,
    new_n14344_, new_n14345_, new_n14346_, new_n14347_, new_n14348_,
    new_n14349_, new_n14350_, new_n14351_, new_n14352_, new_n14353_,
    new_n14354_, new_n14355_, new_n14356_, new_n14357_, new_n14358_,
    new_n14359_, new_n14360_, new_n14361_, new_n14362_, new_n14363_,
    new_n14364_, new_n14365_, new_n14366_, new_n14367_, new_n14368_,
    new_n14369_, new_n14370_, new_n14371_, new_n14372_, new_n14373_,
    new_n14374_, new_n14375_, new_n14376_, new_n14377_, new_n14378_,
    new_n14379_, new_n14380_, new_n14381_, new_n14382_, new_n14383_,
    new_n14384_, new_n14385_, new_n14386_, new_n14387_, new_n14388_,
    new_n14389_, new_n14390_, new_n14391_, new_n14392_, new_n14393_,
    new_n14394_, new_n14395_, new_n14396_, new_n14397_, new_n14398_,
    new_n14399_, new_n14400_, new_n14401_, new_n14402_, new_n14403_,
    new_n14404_, new_n14405_, new_n14406_, new_n14407_, new_n14408_,
    new_n14409_, new_n14410_, new_n14411_, new_n14412_, new_n14413_,
    new_n14414_, new_n14415_, new_n14416_, new_n14417_, new_n14418_,
    new_n14419_, new_n14420_, new_n14421_, new_n14422_, new_n14423_,
    new_n14424_, new_n14425_, new_n14426_, new_n14427_, new_n14428_,
    new_n14429_, new_n14430_, new_n14431_, new_n14432_, new_n14433_,
    new_n14434_, new_n14435_, new_n14436_, new_n14437_, new_n14438_,
    new_n14439_, new_n14440_, new_n14441_, new_n14442_, new_n14443_,
    new_n14444_, new_n14445_, new_n14446_, new_n14447_, new_n14448_,
    new_n14449_, new_n14450_, new_n14451_, new_n14452_, new_n14453_,
    new_n14454_, new_n14455_, new_n14456_, new_n14457_, new_n14458_,
    new_n14459_, new_n14460_, new_n14461_, new_n14462_, new_n14463_,
    new_n14464_, new_n14465_, new_n14466_, new_n14467_, new_n14468_,
    new_n14469_, new_n14470_, new_n14471_, new_n14472_, new_n14473_,
    new_n14474_, new_n14475_, new_n14476_, new_n14477_, new_n14478_,
    new_n14479_, new_n14480_, new_n14481_, new_n14482_, new_n14483_,
    new_n14484_, new_n14485_, new_n14486_, new_n14487_, new_n14488_,
    new_n14489_, new_n14490_, new_n14491_, new_n14492_, new_n14493_,
    new_n14494_, new_n14495_, new_n14496_, new_n14497_, new_n14498_,
    new_n14499_, new_n14500_, new_n14501_, new_n14502_, new_n14503_,
    new_n14504_, new_n14505_, new_n14506_, new_n14507_, new_n14508_,
    new_n14509_, new_n14510_, new_n14511_, new_n14512_, new_n14513_,
    new_n14514_, new_n14515_, new_n14516_, new_n14517_, new_n14518_,
    new_n14519_, new_n14520_, new_n14521_, new_n14522_, new_n14523_,
    new_n14524_, new_n14525_, new_n14526_, new_n14527_, new_n14528_,
    new_n14529_, new_n14530_, new_n14531_, new_n14532_, new_n14533_,
    new_n14534_, new_n14535_, new_n14536_, new_n14537_, new_n14538_,
    new_n14539_, new_n14540_, new_n14541_, new_n14542_, new_n14543_,
    new_n14544_, new_n14545_, new_n14546_, new_n14547_, new_n14548_,
    new_n14549_, new_n14550_, new_n14551_, new_n14552_, new_n14553_,
    new_n14554_, new_n14555_, new_n14556_, new_n14557_, new_n14558_,
    new_n14559_, new_n14560_, new_n14561_, new_n14562_, new_n14563_,
    new_n14564_, new_n14565_, new_n14566_, new_n14567_, new_n14568_,
    new_n14569_, new_n14570_, new_n14571_, new_n14572_, new_n14573_,
    new_n14574_, new_n14575_, new_n14576_, new_n14577_, new_n14578_,
    new_n14579_, new_n14580_, new_n14581_, new_n14582_, new_n14583_,
    new_n14584_, new_n14585_, new_n14586_, new_n14587_, new_n14588_,
    new_n14589_, new_n14590_, new_n14591_, new_n14592_, new_n14593_,
    new_n14594_, new_n14595_, new_n14596_, new_n14597_, new_n14598_,
    new_n14599_, new_n14600_, new_n14601_, new_n14602_, new_n14603_,
    new_n14604_, new_n14605_, new_n14606_, new_n14607_, new_n14609_,
    new_n14610_, new_n14611_, new_n14612_, new_n14613_, new_n14614_,
    new_n14615_, new_n14616_, new_n14617_, new_n14618_, new_n14619_,
    new_n14620_, new_n14621_, new_n14622_, new_n14623_, new_n14624_,
    new_n14625_, new_n14626_, new_n14627_, new_n14628_, new_n14629_,
    new_n14630_, new_n14631_, new_n14632_, new_n14633_, new_n14634_,
    new_n14635_, new_n14636_, new_n14637_, new_n14638_, new_n14639_,
    new_n14640_, new_n14641_, new_n14642_, new_n14643_, new_n14644_,
    new_n14645_, new_n14646_, new_n14647_, new_n14648_, new_n14649_,
    new_n14650_, new_n14651_, new_n14652_, new_n14653_, new_n14654_,
    new_n14655_, new_n14656_, new_n14657_, new_n14658_, new_n14659_,
    new_n14660_, new_n14661_, new_n14662_, new_n14663_, new_n14664_,
    new_n14665_, new_n14666_, new_n14667_, new_n14668_, new_n14669_,
    new_n14670_, new_n14671_, new_n14672_, new_n14673_, new_n14674_,
    new_n14675_, new_n14676_, new_n14677_, new_n14678_, new_n14679_,
    new_n14680_, new_n14681_, new_n14682_, new_n14683_, new_n14684_,
    new_n14685_, new_n14686_, new_n14687_, new_n14688_, new_n14689_,
    new_n14690_, new_n14691_, new_n14692_, new_n14693_, new_n14694_,
    new_n14695_, new_n14696_, new_n14697_, new_n14698_, new_n14699_,
    new_n14700_, new_n14701_, new_n14702_, new_n14703_, new_n14704_,
    new_n14705_, new_n14706_, new_n14707_, new_n14708_, new_n14709_,
    new_n14710_, new_n14711_, new_n14712_, new_n14714_, new_n14715_,
    new_n14716_, new_n14717_, new_n14718_, new_n14719_, new_n14720_,
    new_n14721_, new_n14722_, new_n14723_, new_n14724_, new_n14725_,
    new_n14726_, new_n14727_, new_n14728_, new_n14729_, new_n14730_,
    new_n14731_, new_n14732_, new_n14733_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14739_, new_n14740_,
    new_n14741_, new_n14742_, new_n14743_, new_n14744_, new_n14745_,
    new_n14746_, new_n14747_, new_n14748_, new_n14749_, new_n14750_,
    new_n14751_, new_n14752_, new_n14753_, new_n14754_, new_n14755_,
    new_n14756_, new_n14757_, new_n14758_, new_n14759_, new_n14760_,
    new_n14761_, new_n14762_, new_n14763_, new_n14764_, new_n14765_,
    new_n14766_, new_n14767_, new_n14768_, new_n14769_, new_n14770_,
    new_n14771_, new_n14772_, new_n14773_, new_n14774_, new_n14775_,
    new_n14776_, new_n14777_, new_n14778_, new_n14779_, new_n14780_,
    new_n14781_, new_n14782_, new_n14783_, new_n14784_, new_n14785_,
    new_n14786_, new_n14787_, new_n14788_, new_n14791_, new_n14792_,
    new_n14793_, new_n14794_, new_n14795_, new_n14796_, new_n14797_,
    new_n14798_, new_n14799_, new_n14800_, new_n14801_, new_n14802_,
    new_n14803_, new_n14804_, new_n14805_, new_n14806_, new_n14807_,
    new_n14808_, new_n14809_, new_n14810_, new_n14811_, new_n14812_,
    new_n14813_, new_n14814_, new_n14815_, new_n14816_, new_n14817_,
    new_n14818_, new_n14819_, new_n14820_, new_n14821_, new_n14822_,
    new_n14823_, new_n14824_, new_n14825_, new_n14826_, new_n14827_,
    new_n14828_, new_n14829_, new_n14830_, new_n14831_, new_n14832_,
    new_n14833_, new_n14834_, new_n14835_, new_n14836_, new_n14837_,
    new_n14838_, new_n14839_, new_n14840_, new_n14841_, new_n14844_,
    new_n14845_, new_n14846_, new_n14847_, new_n14848_, new_n14849_,
    new_n14850_, new_n14851_, new_n14852_, new_n14853_, new_n14854_,
    new_n14855_, new_n14856_, new_n14857_, new_n14858_, new_n14859_,
    new_n14860_, new_n14861_, new_n14862_, new_n14863_, new_n14864_,
    new_n14865_, new_n14866_, new_n14867_, new_n14868_, new_n14869_,
    new_n14870_, new_n14871_, new_n14872_, new_n14873_, new_n14874_,
    new_n14875_, new_n14876_, new_n14877_, new_n14878_, new_n14879_,
    new_n14880_, new_n14881_, new_n14882_, new_n14883_, new_n14884_,
    new_n14885_, new_n14886_, new_n14887_, new_n14888_, new_n14889_,
    new_n14890_, new_n14891_, new_n14892_, new_n14893_, new_n14894_,
    new_n14895_, new_n14896_, new_n14897_, new_n14898_, new_n14899_,
    new_n14900_, new_n14901_, new_n14902_, new_n14903_, new_n14904_,
    new_n14905_, new_n14906_, new_n14907_, new_n14908_, new_n14909_,
    new_n14910_, new_n14911_, new_n14912_, new_n14913_, new_n14914_,
    new_n14915_, new_n14916_, new_n14917_, new_n14918_, new_n14919_,
    new_n14920_, new_n14921_, new_n14922_, new_n14923_, new_n14924_,
    new_n14925_, new_n14926_, new_n14927_, new_n14928_, new_n14929_,
    new_n14930_, new_n14931_, new_n14932_, new_n14933_, new_n14934_,
    new_n14935_, new_n14936_, new_n14937_, new_n14938_, new_n14939_,
    new_n14940_, new_n14941_, new_n14942_, new_n14943_, new_n14944_,
    new_n14945_, new_n14946_, new_n14947_, new_n14948_, new_n14949_,
    new_n14950_, new_n14951_, new_n14952_, new_n14953_, new_n14954_,
    new_n14955_, new_n14956_, new_n14957_, new_n14958_, new_n14959_,
    new_n14960_, new_n14961_, new_n14962_, new_n14963_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14981_, new_n14982_, new_n14983_, new_n14984_, new_n14985_,
    new_n14986_, new_n14987_, new_n14988_, new_n14989_, new_n14990_,
    new_n14991_, new_n14992_, new_n14993_, new_n14994_, new_n14995_,
    new_n14996_, new_n14997_, new_n14998_, new_n14999_, new_n15000_,
    new_n15001_, new_n15002_, new_n15003_, new_n15004_, new_n15005_,
    new_n15006_, new_n15007_, new_n15008_, new_n15009_, new_n15010_,
    new_n15011_, new_n15012_, new_n15013_, new_n15014_, new_n15015_,
    new_n15016_, new_n15017_, new_n15019_, new_n15020_, new_n15021_,
    new_n15022_, new_n15023_, new_n15024_, new_n15025_, new_n15026_,
    new_n15027_, new_n15028_, new_n15029_, new_n15030_, new_n15031_,
    new_n15032_, new_n15033_, new_n15034_, new_n15035_, new_n15036_,
    new_n15037_, new_n15038_, new_n15039_, new_n15040_, new_n15041_,
    new_n15042_, new_n15043_, new_n15044_, new_n15045_, new_n15046_,
    new_n15047_, new_n15048_, new_n15049_, new_n15050_, new_n15051_,
    new_n15052_, new_n15053_, new_n15054_, new_n15055_, new_n15056_,
    new_n15057_, new_n15058_, new_n15059_, new_n15060_, new_n15061_,
    new_n15062_, new_n15063_, new_n15064_, new_n15065_, new_n15066_,
    new_n15067_, new_n15068_, new_n15069_, new_n15070_, new_n15071_,
    new_n15072_, new_n15073_, new_n15074_, new_n15075_, new_n15076_,
    new_n15077_, new_n15078_, new_n15079_, new_n15080_, new_n15081_,
    new_n15082_, new_n15083_, new_n15084_, new_n15085_, new_n15086_,
    new_n15087_, new_n15088_, new_n15089_, new_n15090_, new_n15091_,
    new_n15092_, new_n15093_, new_n15094_, new_n15095_, new_n15096_,
    new_n15097_, new_n15098_, new_n15099_, new_n15100_, new_n15101_,
    new_n15102_, new_n15103_, new_n15104_, new_n15105_, new_n15106_,
    new_n15107_, new_n15108_, new_n15109_, new_n15110_, new_n15111_,
    new_n15112_, new_n15113_, new_n15114_, new_n15115_, new_n15116_,
    new_n15117_, new_n15118_, new_n15119_, new_n15120_, new_n15121_,
    new_n15122_, new_n15123_, new_n15124_, new_n15125_, new_n15126_,
    new_n15127_, new_n15128_, new_n15129_, new_n15130_, new_n15131_,
    new_n15132_, new_n15133_, new_n15134_, new_n15135_, new_n15136_,
    new_n15137_, new_n15138_, new_n15139_, new_n15140_, new_n15141_,
    new_n15142_, new_n15143_, new_n15144_, new_n15145_, new_n15146_,
    new_n15147_, new_n15148_, new_n15149_, new_n15150_, new_n15151_,
    new_n15152_, new_n15153_, new_n15154_, new_n15155_, new_n15156_,
    new_n15157_, new_n15158_, new_n15159_, new_n15160_, new_n15161_,
    new_n15162_, new_n15163_, new_n15164_, new_n15165_, new_n15166_,
    new_n15167_, new_n15168_, new_n15169_, new_n15170_, new_n15171_,
    new_n15172_, new_n15173_, new_n15174_, new_n15175_, new_n15176_,
    new_n15177_, new_n15178_, new_n15179_, new_n15180_, new_n15181_,
    new_n15182_, new_n15183_, new_n15184_, new_n15185_, new_n15186_,
    new_n15187_, new_n15188_, new_n15189_, new_n15190_, new_n15191_,
    new_n15192_, new_n15193_, new_n15194_, new_n15195_, new_n15196_,
    new_n15197_, new_n15198_, new_n15199_, new_n15200_, new_n15201_,
    new_n15202_, new_n15203_, new_n15204_, new_n15205_, new_n15207_,
    new_n15208_, new_n15209_, new_n15210_, new_n15211_, new_n15212_,
    new_n15213_, new_n15214_, new_n15215_, new_n15216_, new_n15217_,
    new_n15218_, new_n15219_, new_n15220_, new_n15221_, new_n15222_,
    new_n15223_, new_n15224_, new_n15225_, new_n15226_, new_n15227_,
    new_n15228_, new_n15229_, new_n15230_, new_n15231_, new_n15232_,
    new_n15242_, new_n15243_, new_n15244_, new_n15245_, new_n15246_,
    new_n15247_, new_n15248_, new_n15249_, new_n15250_, new_n15251_,
    new_n15252_, new_n15253_, new_n15254_, new_n15255_, new_n15256_,
    new_n15257_, new_n15258_, new_n15259_, new_n15260_, new_n15261_,
    new_n15262_, new_n15263_, new_n15264_, new_n15265_, new_n15266_,
    new_n15267_, new_n15268_, new_n15269_, new_n15270_, new_n15271_,
    new_n15272_, new_n15273_, new_n15274_, new_n15275_, new_n15276_,
    new_n15277_, new_n15278_, new_n15279_, new_n15280_, new_n15281_,
    new_n15282_, new_n15283_, new_n15284_, new_n15285_, new_n15286_,
    new_n15287_, new_n15288_, new_n15289_, new_n15290_, new_n15291_,
    new_n15292_, new_n15293_, new_n15294_, new_n15295_, new_n15296_,
    new_n15299_, new_n15300_, new_n15301_, new_n15302_, new_n15303_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15335_, new_n15336_, new_n15337_, new_n15338_, new_n15339_,
    new_n15340_, new_n15341_, new_n15342_, new_n15343_, new_n15344_,
    new_n15345_, new_n15347_, new_n15348_, new_n15349_, new_n15350_,
    new_n15351_, new_n15352_, new_n15353_, new_n15354_, new_n15355_,
    new_n15356_, new_n15357_, new_n15358_, new_n15359_, new_n15360_,
    new_n15361_, new_n15362_, new_n15363_, new_n15364_, new_n15365_,
    new_n15366_, new_n15367_, new_n15368_, new_n15369_, new_n15370_,
    new_n15371_, new_n15372_, new_n15373_, new_n15374_, new_n15375_,
    new_n15376_, new_n15377_, new_n15378_, new_n15379_, new_n15380_,
    new_n15381_, new_n15383_, new_n15384_, new_n15385_, new_n15386_,
    new_n15387_, new_n15388_, new_n15389_, new_n15390_, new_n15391_,
    new_n15392_, new_n15393_, new_n15394_, new_n15395_, new_n15396_,
    new_n15397_, new_n15398_, new_n15399_, new_n15400_, new_n15401_,
    new_n15402_, new_n15403_, new_n15404_, new_n15405_, new_n15406_,
    new_n15407_, new_n15408_, new_n15409_, new_n15410_, new_n15411_,
    new_n15412_, new_n15413_, new_n15414_, new_n15415_, new_n15416_,
    new_n15417_, new_n15418_, new_n15419_, new_n15420_, new_n15421_,
    new_n15423_, new_n15424_, new_n15425_, new_n15426_, new_n15427_,
    new_n15428_, new_n15429_, new_n15430_, new_n15431_, new_n15432_,
    new_n15433_, new_n15434_, new_n15435_, new_n15436_, new_n15437_,
    new_n15438_, new_n15439_, new_n15440_, new_n15441_, new_n15442_,
    new_n15443_, new_n15444_, new_n15445_, new_n15446_, new_n15447_,
    new_n15448_, new_n15449_, new_n15450_, new_n15451_, new_n15452_,
    new_n15453_, new_n15454_, new_n15455_, new_n15456_, new_n15457_,
    new_n15458_, new_n15459_, new_n15460_, new_n15461_, new_n15462_,
    new_n15463_, new_n15464_, new_n15465_, new_n15466_, new_n15467_,
    new_n15469_, new_n15470_, new_n15471_, new_n15472_, new_n15473_,
    new_n15474_, new_n15475_, new_n15476_, new_n15477_, new_n15478_,
    new_n15479_, new_n15480_, new_n15481_, new_n15482_, new_n15483_,
    new_n15484_, new_n15485_, new_n15486_, new_n15487_, new_n15488_,
    new_n15489_, new_n15490_, new_n15491_, new_n15492_, new_n15493_,
    new_n15494_, new_n15495_, new_n15496_, new_n15497_, new_n15498_,
    new_n15499_, new_n15500_, new_n15501_, new_n15502_, new_n15503_,
    new_n15504_, new_n15505_, new_n15506_, new_n15507_, new_n15509_,
    new_n15510_, new_n15511_, new_n15512_, new_n15513_, new_n15514_,
    new_n15515_, new_n15516_, new_n15517_, new_n15518_, new_n15519_,
    new_n15520_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15526_, new_n15527_, new_n15528_, new_n15529_,
    new_n15530_, new_n15531_, new_n15532_, new_n15533_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15546_, new_n15547_, new_n15548_, new_n15549_, new_n15550_,
    new_n15551_, new_n15552_, new_n15553_, new_n15554_, new_n15555_,
    new_n15556_, new_n15557_, new_n15558_, new_n15559_, new_n15560_,
    new_n15561_, new_n15562_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15572_, new_n15573_, new_n15574_, new_n15576_,
    new_n15577_, new_n15578_, new_n15579_, new_n15580_, new_n15581_,
    new_n15582_, new_n15583_, new_n15584_, new_n15585_, new_n15586_,
    new_n15587_, new_n15588_, new_n15589_, new_n15590_, new_n15591_,
    new_n15592_, new_n15593_, new_n15594_, new_n15595_, new_n15596_,
    new_n15597_, new_n15598_, new_n15599_, new_n15600_, new_n15601_,
    new_n15602_, new_n15603_, new_n15604_, new_n15605_, new_n15606_,
    new_n15607_, new_n15608_, new_n15609_, new_n15610_, new_n15611_,
    new_n15612_, new_n15613_, new_n15614_, new_n15615_, new_n15616_,
    new_n15617_, new_n15618_, new_n15619_, new_n15620_, new_n15621_,
    new_n15622_, new_n15623_, new_n15624_, new_n15626_, new_n15627_,
    new_n15628_, new_n15629_, new_n15630_, new_n15631_, new_n15632_,
    new_n15633_, new_n15634_, new_n15635_, new_n15636_, new_n15637_,
    new_n15638_, new_n15639_, new_n15640_, new_n15641_, new_n15642_,
    new_n15643_, new_n15644_, new_n15645_, new_n15646_, new_n15647_,
    new_n15648_, new_n15649_, new_n15650_, new_n15651_, new_n15652_,
    new_n15653_, new_n15654_, new_n15655_, new_n15656_, new_n15657_,
    new_n15658_, new_n15659_, new_n15660_, new_n15661_, new_n15662_,
    new_n15663_, new_n15664_, new_n15665_, new_n15666_, new_n15667_,
    new_n15668_, new_n15669_, new_n15670_, new_n15671_, new_n15672_,
    new_n15673_, new_n15674_, new_n15675_, new_n15676_, new_n15677_,
    new_n15678_, new_n15679_, new_n15680_, new_n15681_, new_n15682_,
    new_n15683_, new_n15684_, new_n15685_, new_n15686_, new_n15687_,
    new_n15688_, new_n15689_, new_n15690_, new_n15691_, new_n15692_,
    new_n15693_, new_n15695_, new_n15696_, new_n15697_, new_n15698_,
    new_n15699_, new_n15700_, new_n15701_, new_n15703_, new_n15704_,
    new_n15705_, new_n15706_, new_n15707_, new_n15708_, new_n15709_,
    new_n15710_, new_n15711_, new_n15712_, new_n15713_, new_n15714_,
    new_n15715_, new_n15716_, new_n15717_, new_n15718_, new_n15719_,
    new_n15720_, new_n15721_, new_n15722_, new_n15723_, new_n15724_,
    new_n15725_, new_n15726_, new_n15727_, new_n15728_, new_n15729_,
    new_n15730_, new_n15731_, new_n15732_, new_n15733_, new_n15734_,
    new_n15735_, new_n15736_, new_n15737_, new_n15738_, new_n15739_,
    new_n15740_, new_n15741_, new_n15742_, new_n15743_, new_n15744_,
    new_n15745_, new_n15746_, new_n15747_, new_n15748_, new_n15749_,
    new_n15750_, new_n15751_, new_n15752_, new_n15753_, new_n15754_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15766_,
    new_n15767_, new_n15768_, new_n15769_, new_n15770_, new_n15771_,
    new_n15772_, new_n15773_, new_n15774_, new_n15775_, new_n15776_,
    new_n15777_, new_n15778_, new_n15779_, new_n15780_, new_n15781_,
    new_n15782_, new_n15783_, new_n15784_, new_n15785_, new_n15787_,
    new_n15788_, new_n15789_, new_n15790_, new_n15791_, new_n15792_,
    new_n15793_, new_n15794_, new_n15795_, new_n15796_, new_n15797_,
    new_n15798_, new_n15799_, new_n15800_, new_n15801_, new_n15802_,
    new_n15803_, new_n15804_, new_n15805_, new_n15806_, new_n15807_,
    new_n15808_, new_n15809_, new_n15811_, new_n15812_, new_n15813_,
    new_n15814_, new_n15815_, new_n15816_, new_n15817_, new_n15818_,
    new_n15819_, new_n15820_, new_n15821_, new_n15822_, new_n15823_,
    new_n15824_, new_n15825_, new_n15826_, new_n15827_, new_n15828_,
    new_n15830_, new_n15831_, new_n15832_, new_n15833_, new_n15834_,
    new_n15835_, new_n15836_, new_n15837_, new_n15838_, new_n15839_,
    new_n15840_, new_n15841_, new_n15842_, new_n15843_, new_n15844_,
    new_n15845_, new_n15846_, new_n15847_, new_n15848_, new_n15849_,
    new_n15850_, new_n15851_, new_n15852_, new_n15853_, new_n15854_,
    new_n15855_, new_n15856_, new_n15857_, new_n15858_, new_n15859_,
    new_n15860_, new_n15861_, new_n15862_, new_n15863_, new_n15864_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15881_, new_n15882_, new_n15883_, new_n15884_, new_n15885_,
    new_n15886_, new_n15887_, new_n15888_, new_n15889_, new_n15890_,
    new_n15891_, new_n15892_, new_n15893_, new_n15894_, new_n15896_,
    new_n15897_, new_n15898_, new_n15899_, new_n15900_, new_n15901_,
    new_n15902_, new_n15903_, new_n15904_, new_n15905_, new_n15906_,
    new_n15907_, new_n15908_, new_n15909_, new_n15910_, new_n15911_,
    new_n15912_, new_n15913_, new_n15914_, new_n15915_, new_n15916_,
    new_n15917_, new_n15918_, new_n15919_, new_n15920_, new_n15921_,
    new_n15922_, new_n15923_, new_n15924_, new_n15926_, new_n15927_,
    new_n15928_, new_n15929_, new_n15930_, new_n15931_, new_n15932_,
    new_n15933_, new_n15934_, new_n15935_, new_n15936_, new_n15937_,
    new_n15938_, new_n15939_, new_n15940_, new_n15941_, new_n15942_,
    new_n15943_, new_n15944_, new_n15945_, new_n15946_, new_n15947_,
    new_n15948_, new_n15949_, new_n15950_, new_n15951_, new_n15952_,
    new_n15953_, new_n15954_, new_n15955_, new_n15956_, new_n15957_,
    new_n15958_, new_n15960_, new_n15961_, new_n15962_, new_n15963_,
    new_n15964_, new_n15965_, new_n15966_, new_n15967_, new_n15968_,
    new_n15969_, new_n15970_, new_n15971_, new_n15972_, new_n15973_,
    new_n15974_, new_n15975_, new_n15976_, new_n15977_, new_n15978_,
    new_n15979_, new_n15980_, new_n15981_, new_n15982_, new_n15983_,
    new_n15984_, new_n15985_, new_n15986_, new_n15987_, new_n15988_,
    new_n15989_, new_n15990_, new_n15991_, new_n15992_, new_n15993_,
    new_n15994_, new_n15995_, new_n15996_, new_n15997_, new_n15998_,
    new_n15999_, new_n16000_, new_n16001_, new_n16002_, new_n16003_,
    new_n16004_, new_n16005_, new_n16006_, new_n16008_, new_n16009_,
    new_n16010_, new_n16011_, new_n16012_, new_n16013_, new_n16014_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16031_, new_n16032_, new_n16033_, new_n16034_, new_n16035_,
    new_n16036_, new_n16037_, new_n16038_, new_n16039_, new_n16040_,
    new_n16041_, new_n16042_, new_n16043_, new_n16044_, new_n16045_,
    new_n16046_, new_n16047_, new_n16049_, new_n16050_, new_n16051_,
    new_n16052_, new_n16053_, new_n16054_, new_n16055_, new_n16056_,
    new_n16057_, new_n16058_, new_n16059_, new_n16060_, new_n16061_,
    new_n16062_, new_n16063_, new_n16064_, new_n16065_, new_n16066_,
    new_n16067_, new_n16068_, new_n16069_, new_n16070_, new_n16071_,
    new_n16072_, new_n16073_, new_n16074_, new_n16075_, new_n16076_,
    new_n16077_, new_n16078_, new_n16079_, new_n16080_, new_n16081_,
    new_n16083_, new_n16084_, new_n16085_, new_n16086_, new_n16087_,
    new_n16088_, new_n16089_, new_n16091_, new_n16092_, new_n16093_,
    new_n16094_, new_n16095_, new_n16096_, new_n16097_, new_n16098_,
    new_n16099_, new_n16100_, new_n16101_, new_n16102_, new_n16103_,
    new_n16104_, new_n16105_, new_n16107_, new_n16108_, new_n16109_,
    new_n16110_, new_n16111_, new_n16112_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16128_, new_n16129_, new_n16130_, new_n16131_,
    new_n16132_, new_n16133_, new_n16134_, new_n16135_, new_n16136_,
    new_n16137_, new_n16138_, new_n16139_, new_n16140_, new_n16141_,
    new_n16142_, new_n16143_, new_n16144_, new_n16145_, new_n16146_,
    new_n16147_, new_n16148_, new_n16149_, new_n16150_, new_n16151_,
    new_n16152_, new_n16153_, new_n16154_, new_n16155_, new_n16156_,
    new_n16157_, new_n16158_, new_n16159_, new_n16160_, new_n16161_,
    new_n16162_, new_n16163_, new_n16166_, new_n16167_, new_n16168_,
    new_n16169_, new_n16170_, new_n16171_, new_n16172_, new_n16173_,
    new_n16174_, new_n16175_, new_n16176_, new_n16177_, new_n16178_,
    new_n16179_, new_n16180_, new_n16181_, new_n16182_, new_n16183_,
    new_n16184_, new_n16185_, new_n16186_, new_n16187_, new_n16188_,
    new_n16189_, new_n16190_, new_n16192_, new_n16193_, new_n16194_,
    new_n16196_, new_n16197_, new_n16198_, new_n16199_, new_n16200_,
    new_n16201_, new_n16203_, new_n16204_, new_n16205_, new_n16206_,
    new_n16207_, new_n16208_, new_n16209_, new_n16210_, new_n16211_,
    new_n16212_, new_n16213_, new_n16214_, new_n16215_, new_n16216_,
    new_n16218_, new_n16219_, new_n16220_, new_n16221_, new_n16222_,
    new_n16223_, new_n16224_, new_n16225_, new_n16226_, new_n16227_,
    new_n16228_, new_n16229_, new_n16230_, new_n16231_, new_n16232_,
    new_n16233_, new_n16234_, new_n16235_, new_n16236_, new_n16237_,
    new_n16238_, new_n16239_, new_n16240_, new_n16241_, new_n16242_,
    new_n16243_, new_n16244_, new_n16245_, new_n16246_, new_n16247_,
    new_n16248_, new_n16249_, new_n16250_, new_n16251_, new_n16252_,
    new_n16253_, new_n16254_, new_n16255_, new_n16256_, new_n16257_,
    new_n16258_, new_n16259_, new_n16260_, new_n16261_, new_n16262_,
    new_n16263_, new_n16264_, new_n16266_, new_n16267_, new_n16268_,
    new_n16269_, new_n16270_, new_n16271_, new_n16272_, new_n16273_,
    new_n16274_, new_n16275_, new_n16276_, new_n16277_, new_n16278_,
    new_n16279_, new_n16280_, new_n16281_, new_n16282_, new_n16283_,
    new_n16284_, new_n16285_, new_n16286_, new_n16287_, new_n16288_,
    new_n16289_, new_n16290_, new_n16291_, new_n16292_, new_n16293_,
    new_n16294_, new_n16295_, new_n16296_, new_n16297_, new_n16298_,
    new_n16299_, new_n16300_, new_n16301_, new_n16302_, new_n16303_,
    new_n16304_, new_n16305_, new_n16306_, new_n16307_, new_n16308_,
    new_n16309_, new_n16310_, new_n16311_, new_n16312_, new_n16314_,
    new_n16315_, new_n16316_, new_n16317_, new_n16318_, new_n16319_,
    new_n16320_, new_n16321_, new_n16322_, new_n16323_, new_n16324_,
    new_n16325_, new_n16326_, new_n16327_, new_n16328_, new_n16329_,
    new_n16330_, new_n16331_, new_n16332_, new_n16333_, new_n16334_,
    new_n16335_, new_n16336_, new_n16337_, new_n16338_, new_n16339_,
    new_n16340_, new_n16341_, new_n16342_, new_n16343_, new_n16344_,
    new_n16345_, new_n16346_, new_n16347_, new_n16348_, new_n16349_,
    new_n16350_, new_n16351_, new_n16352_, new_n16353_, new_n16354_,
    new_n16355_, new_n16356_, new_n16357_, new_n16358_, new_n16359_,
    new_n16360_, new_n16361_, new_n16362_, new_n16364_, new_n16365_,
    new_n16366_, new_n16367_, new_n16368_, new_n16369_, new_n16370_,
    new_n16371_, new_n16372_, new_n16373_, new_n16374_, new_n16375_,
    new_n16376_, new_n16377_, new_n16378_, new_n16379_, new_n16380_,
    new_n16381_, new_n16382_, new_n16383_, new_n16384_, new_n16385_,
    new_n16386_, new_n16387_, new_n16388_, new_n16389_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16395_,
    new_n16396_, new_n16397_, new_n16398_, new_n16399_, new_n16400_,
    new_n16401_, new_n16402_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16412_, new_n16413_, new_n16414_, new_n16415_, new_n16416_,
    new_n16417_, new_n16418_, new_n16419_, new_n16420_, new_n16421_,
    new_n16422_, new_n16423_, new_n16424_, new_n16425_, new_n16426_,
    new_n16427_, new_n16428_, new_n16429_, new_n16430_, new_n16431_,
    new_n16432_, new_n16433_, new_n16434_, new_n16435_, new_n16436_,
    new_n16437_, new_n16438_, new_n16439_, new_n16440_, new_n16441_,
    new_n16442_, new_n16443_, new_n16444_, new_n16445_, new_n16446_,
    new_n16447_, new_n16448_, new_n16449_, new_n16450_, new_n16451_,
    new_n16452_, new_n16453_, new_n16454_, new_n16455_, new_n16456_,
    new_n16457_, new_n16459_, new_n16460_, new_n16461_, new_n16462_,
    new_n16463_, new_n16464_, new_n16465_, new_n16466_, new_n16467_,
    new_n16468_, new_n16469_, new_n16470_, new_n16471_, new_n16472_,
    new_n16473_, new_n16474_, new_n16475_, new_n16476_, new_n16477_,
    new_n16478_, new_n16479_, new_n16480_, new_n16481_, new_n16482_,
    new_n16483_, new_n16484_, new_n16485_, new_n16486_, new_n16487_,
    new_n16488_, new_n16489_, new_n16490_, new_n16491_, new_n16492_,
    new_n16493_, new_n16494_, new_n16495_, new_n16496_, new_n16497_,
    new_n16498_, new_n16499_, new_n16500_, new_n16501_, new_n16502_,
    new_n16503_, new_n16504_, new_n16505_, new_n16506_, new_n16507_,
    new_n16508_, new_n16509_, new_n16510_, new_n16511_, new_n16512_,
    new_n16513_, new_n16514_, new_n16515_, new_n16516_, new_n16517_,
    new_n16518_, new_n16519_, new_n16520_, new_n16521_, new_n16522_,
    new_n16523_, new_n16524_, new_n16525_, new_n16526_, new_n16527_,
    new_n16528_, new_n16529_, new_n16530_, new_n16531_, new_n16532_,
    new_n16533_, new_n16534_, new_n16536_, new_n16537_, new_n16538_,
    new_n16539_, new_n16540_, new_n16541_, new_n16542_, new_n16543_,
    new_n16544_, new_n16545_, new_n16546_, new_n16547_, new_n16548_,
    new_n16549_, new_n16550_, new_n16551_, new_n16552_, new_n16553_,
    new_n16554_, new_n16555_, new_n16556_, new_n16557_, new_n16558_,
    new_n16559_, new_n16560_, new_n16561_, new_n16562_, new_n16563_,
    new_n16564_, new_n16565_, new_n16566_, new_n16567_, new_n16568_,
    new_n16569_, new_n16570_, new_n16571_, new_n16572_, new_n16573_,
    new_n16574_, new_n16575_, new_n16576_, new_n16577_, new_n16578_,
    new_n16579_, new_n16580_, new_n16581_, new_n16582_, new_n16583_,
    new_n16584_, new_n16585_, new_n16586_, new_n16587_, new_n16588_,
    new_n16589_, new_n16590_, new_n16591_, new_n16592_, new_n16593_,
    new_n16594_, new_n16595_, new_n16596_, new_n16597_, new_n16598_,
    new_n16599_, new_n16600_, new_n16601_, new_n16602_, new_n16603_,
    new_n16604_, new_n16605_, new_n16606_, new_n16607_, new_n16608_,
    new_n16609_, new_n16610_, new_n16611_, new_n16612_, new_n16613_,
    new_n16614_, new_n16615_, new_n16616_, new_n16617_, new_n16618_,
    new_n16619_, new_n16620_, new_n16621_, new_n16622_, new_n16623_,
    new_n16624_, new_n16625_, new_n16626_, new_n16627_, new_n16628_,
    new_n16629_, new_n16630_, new_n16631_, new_n16632_, new_n16633_,
    new_n16634_, new_n16635_, new_n16636_, new_n16637_, new_n16638_,
    new_n16639_, new_n16640_, new_n16641_, new_n16642_, new_n16644_,
    new_n16645_, new_n16646_, new_n16647_, new_n16648_, new_n16649_,
    new_n16650_, new_n16651_, new_n16652_, new_n16653_, new_n16654_,
    new_n16655_, new_n16656_, new_n16657_, new_n16658_, new_n16659_,
    new_n16660_, new_n16661_, new_n16662_, new_n16663_, new_n16664_,
    new_n16665_, new_n16675_, new_n16676_, new_n16677_, new_n16678_,
    new_n16679_, new_n16680_, new_n16681_, new_n16682_, new_n16683_,
    new_n16684_, new_n16685_, new_n16686_, new_n16687_, new_n16688_,
    new_n16689_, new_n16690_, new_n16691_, new_n16692_, new_n16693_,
    new_n16694_, new_n16695_, new_n16696_, new_n16697_, new_n16698_,
    new_n16699_, new_n16700_, new_n16701_, new_n16702_, new_n16703_,
    new_n16704_, new_n16705_, new_n16706_, new_n16707_, new_n16708_,
    new_n16709_, new_n16710_, new_n16711_, new_n16712_, new_n16713_,
    new_n16714_, new_n16715_, new_n16716_, new_n16717_, new_n16718_,
    new_n16719_, new_n16720_, new_n16721_, new_n16722_, new_n16723_,
    new_n16724_, new_n16725_, new_n16726_, new_n16727_, new_n16728_,
    new_n16731_, new_n16732_, new_n16733_, new_n16734_, new_n16735_,
    new_n16737_, new_n16738_, new_n16739_, new_n16740_, new_n16741_,
    new_n16742_, new_n16743_, new_n16744_, new_n16745_, new_n16746_,
    new_n16747_, new_n16748_, new_n16749_, new_n16750_, new_n16751_,
    new_n16752_, new_n16753_, new_n16754_, new_n16755_, new_n16756_,
    new_n16757_, new_n16758_, new_n16759_, new_n16760_, new_n16761_,
    new_n16762_, new_n16763_, new_n16764_, new_n16765_, new_n16766_,
    new_n16767_, new_n16768_, new_n16769_, new_n16770_, new_n16771_,
    new_n16772_, new_n16773_, new_n16774_, new_n16775_, new_n16776_,
    new_n16777_, new_n16778_, new_n16779_, new_n16780_, new_n16781_,
    new_n16782_, new_n16783_, new_n16784_, new_n16785_, new_n16786_,
    new_n16787_, new_n16788_, new_n16789_, new_n16790_, new_n16791_,
    new_n16792_, new_n16793_, new_n16794_, new_n16795_, new_n16796_,
    new_n16797_, new_n16798_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16817_, new_n16818_, new_n16819_, new_n16820_, new_n16821_,
    new_n16822_, new_n16823_, new_n16824_, new_n16825_, new_n16826_,
    new_n16827_, new_n16828_, new_n16829_, new_n16830_, new_n16831_,
    new_n16832_, new_n16833_, new_n16834_, new_n16835_, new_n16836_,
    new_n16837_, new_n16838_, new_n16839_, new_n16840_, new_n16841_,
    new_n16842_, new_n16843_, new_n16844_, new_n16845_, new_n16846_,
    new_n16847_, new_n16848_, new_n16849_, new_n16850_, new_n16851_,
    new_n16852_, new_n16853_, new_n16854_, new_n16855_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16862_, new_n16863_, new_n16864_, new_n16865_, new_n16866_,
    new_n16867_, new_n16868_, new_n16869_, new_n16870_, new_n16871_,
    new_n16872_, new_n16873_, new_n16874_, new_n16875_, new_n16876_,
    new_n16877_, new_n16878_, new_n16879_, new_n16880_, new_n16881_,
    new_n16882_, new_n16883_, new_n16884_, new_n16887_, new_n16888_,
    new_n16889_, new_n16890_, new_n16891_, new_n16892_, new_n16893_,
    new_n16894_, new_n16895_, new_n16896_, new_n16897_, new_n16898_,
    new_n16899_, new_n16900_, new_n16901_, new_n16902_, new_n16903_,
    new_n16904_, new_n16905_, new_n16906_, new_n16907_, new_n16908_,
    new_n16909_, new_n16910_, new_n16911_, new_n16912_, new_n16913_,
    new_n16914_, new_n16915_, new_n16916_, new_n16917_, new_n16918_,
    new_n16919_, new_n16920_, new_n16921_, new_n16922_, new_n16923_,
    new_n16924_, new_n16925_, new_n16926_, new_n16927_, new_n16928_,
    new_n16929_, new_n16930_, new_n16931_, new_n16932_, new_n16933_,
    new_n16934_, new_n16935_, new_n16936_, new_n16937_, new_n16938_,
    new_n16939_, new_n16940_, new_n16941_, new_n16942_, new_n16943_,
    new_n16944_, new_n16945_, new_n16946_, new_n16947_, new_n16948_,
    new_n16949_, new_n16950_, new_n16951_, new_n16952_, new_n16953_,
    new_n16954_, new_n16955_, new_n16956_, new_n16957_, new_n16958_,
    new_n16959_, new_n16960_, new_n16961_, new_n16962_, new_n16963_,
    new_n16964_, new_n16965_, new_n16966_, new_n16967_, new_n16968_,
    new_n16969_, new_n16970_, new_n16971_, new_n16972_, new_n16973_,
    new_n16974_, new_n16975_, new_n16976_, new_n16977_, new_n16978_,
    new_n16979_, new_n16980_, new_n16981_, new_n16982_, new_n16983_,
    new_n16984_, new_n16985_, new_n16986_, new_n16987_, new_n16988_,
    new_n16989_, new_n16990_, new_n16991_, new_n16992_, new_n16993_,
    new_n16994_, new_n16995_, new_n16996_, new_n16997_, new_n16998_,
    new_n16999_, new_n17000_, new_n17001_, new_n17002_, new_n17003_,
    new_n17004_, new_n17005_, new_n17006_, new_n17007_, new_n17008_,
    new_n17009_, new_n17010_, new_n17011_, new_n17012_, new_n17013_,
    new_n17014_, new_n17015_, new_n17016_, new_n17017_, new_n17018_,
    new_n17019_, new_n17020_, new_n17021_, new_n17022_, new_n17023_,
    new_n17024_, new_n17025_, new_n17026_, new_n17027_, new_n17028_,
    new_n17029_, new_n17030_, new_n17031_, new_n17032_, new_n17033_,
    new_n17034_, new_n17035_, new_n17036_, new_n17037_, new_n17038_,
    new_n17039_, new_n17040_, new_n17041_, new_n17042_, new_n17043_,
    new_n17044_, new_n17045_, new_n17046_, new_n17047_, new_n17048_,
    new_n17049_, new_n17050_, new_n17051_, new_n17052_, new_n17053_,
    new_n17054_, new_n17055_, new_n17056_, new_n17057_, new_n17058_,
    new_n17059_, new_n17060_, new_n17061_, new_n17062_, new_n17063_,
    new_n17064_, new_n17065_, new_n17066_, new_n17067_, new_n17068_,
    new_n17069_, new_n17070_, new_n17071_, new_n17072_, new_n17073_,
    new_n17074_, new_n17075_, new_n17076_, new_n17077_, new_n17078_,
    new_n17079_, new_n17081_, new_n17082_, new_n17083_, new_n17084_,
    new_n17085_, new_n17086_, new_n17087_, new_n17088_, new_n17089_,
    new_n17090_, new_n17091_, new_n17092_, new_n17093_, new_n17094_,
    new_n17095_, new_n17096_, new_n17097_, new_n17098_, new_n17099_,
    new_n17100_, new_n17101_, new_n17102_, new_n17103_, new_n17104_,
    new_n17105_, new_n17106_, new_n17107_, new_n17108_, new_n17109_,
    new_n17110_, new_n17111_, new_n17112_, new_n17113_, new_n17114_,
    new_n17115_, new_n17117_, new_n17118_, new_n17119_, new_n17120_,
    new_n17121_, new_n17122_, new_n17123_, new_n17124_, new_n17125_,
    new_n17126_, new_n17127_, new_n17128_, new_n17129_, new_n17130_,
    new_n17131_, new_n17132_, new_n17133_, new_n17134_, new_n17135_,
    new_n17136_, new_n17137_, new_n17138_, new_n17139_, new_n17140_,
    new_n17141_, new_n17142_, new_n17143_, new_n17144_, new_n17145_,
    new_n17146_, new_n17147_, new_n17148_, new_n17149_, new_n17150_,
    new_n17151_, new_n17152_, new_n17153_, new_n17154_, new_n17155_,
    new_n17156_, new_n17157_, new_n17158_, new_n17159_, new_n17160_,
    new_n17161_, new_n17162_, new_n17163_, new_n17164_, new_n17165_,
    new_n17166_, new_n17167_, new_n17168_, new_n17169_, new_n17170_,
    new_n17171_, new_n17172_, new_n17173_, new_n17174_, new_n17175_,
    new_n17176_, new_n17177_, new_n17178_, new_n17179_, new_n17180_,
    new_n17181_, new_n17182_, new_n17183_, new_n17184_, new_n17185_,
    new_n17186_, new_n17187_, new_n17188_, new_n17189_, new_n17190_,
    new_n17191_, new_n17192_, new_n17193_, new_n17194_, new_n17195_,
    new_n17196_, new_n17197_, new_n17198_, new_n17199_, new_n17200_,
    new_n17201_, new_n17202_, new_n17203_, new_n17204_, new_n17205_,
    new_n17206_, new_n17207_, new_n17208_, new_n17209_, new_n17210_,
    new_n17211_, new_n17212_, new_n17213_, new_n17214_, new_n17215_,
    new_n17216_, new_n17217_, new_n17218_, new_n17219_, new_n17220_,
    new_n17221_, new_n17222_, new_n17223_, new_n17224_, new_n17225_,
    new_n17226_, new_n17227_, new_n17228_, new_n17229_, new_n17230_,
    new_n17231_, new_n17232_, new_n17233_, new_n17234_, new_n17235_,
    new_n17236_, new_n17237_, new_n17238_, new_n17239_, new_n17240_,
    new_n17241_, new_n17242_, new_n17243_, new_n17244_, new_n17245_,
    new_n17246_, new_n17247_, new_n17248_, new_n17249_, new_n17250_,
    new_n17251_, new_n17252_, new_n17253_, new_n17254_, new_n17255_,
    new_n17256_, new_n17257_, new_n17258_, new_n17259_, new_n17260_,
    new_n17261_, new_n17262_, new_n17263_, new_n17264_, new_n17265_,
    new_n17266_, new_n17267_, new_n17268_, new_n17269_, new_n17270_,
    new_n17271_, new_n17272_, new_n17273_, new_n17274_, new_n17275_,
    new_n17276_, new_n17277_, new_n17278_, new_n17279_, new_n17280_,
    new_n17281_, new_n17282_, new_n17283_, new_n17284_, new_n17285_,
    new_n17286_, new_n17287_, new_n17288_, new_n17289_, new_n17290_,
    new_n17291_, new_n17292_, new_n17293_, new_n17294_, new_n17295_,
    new_n17296_, new_n17297_, new_n17298_, new_n17299_, new_n17300_,
    new_n17301_, new_n17302_, new_n17303_, new_n17304_, new_n17305_,
    new_n17306_, new_n17307_, new_n17308_, new_n17309_, new_n17310_,
    new_n17311_, new_n17312_, new_n17313_, new_n17314_, new_n17315_,
    new_n17316_, new_n17317_, new_n17318_, new_n17319_, new_n17320_,
    new_n17321_, new_n17322_, new_n17323_, new_n17324_, new_n17325_,
    new_n17326_, new_n17327_, new_n17328_, new_n17329_, new_n17330_,
    new_n17331_, new_n17332_, new_n17333_, new_n17334_, new_n17335_,
    new_n17336_, new_n17337_, new_n17338_, new_n17339_, new_n17340_,
    new_n17341_, new_n17342_, new_n17343_, new_n17344_, new_n17345_,
    new_n17346_, new_n17347_, new_n17348_, new_n17349_, new_n17350_,
    new_n17351_, new_n17352_, new_n17353_, new_n17354_, new_n17355_,
    new_n17356_, new_n17357_, new_n17358_, new_n17359_, new_n17360_,
    new_n17361_, new_n17362_, new_n17363_, new_n17364_, new_n17365_,
    new_n17366_, new_n17367_, new_n17368_, new_n17369_, new_n17370_,
    new_n17371_, new_n17372_, new_n17373_, new_n17374_, new_n17375_,
    new_n17376_, new_n17377_, new_n17378_, new_n17379_, new_n17381_,
    new_n17382_, new_n17383_, new_n17384_, new_n17385_, new_n17386_,
    new_n17387_, new_n17388_, new_n17389_, new_n17390_, new_n17391_,
    new_n17392_, new_n17393_, new_n17394_, new_n17395_, new_n17396_,
    new_n17397_, new_n17398_, new_n17399_, new_n17400_, new_n17401_,
    new_n17402_, new_n17403_, new_n17404_, new_n17405_, new_n17406_,
    new_n17407_, new_n17408_, new_n17409_, new_n17410_, new_n17411_,
    new_n17412_, new_n17413_, new_n17414_, new_n17415_, new_n17416_,
    new_n17417_, new_n17419_, new_n17420_, new_n17421_, new_n17422_,
    new_n17423_, new_n17424_, new_n17425_, new_n17426_, new_n17427_,
    new_n17428_, new_n17429_, new_n17430_, new_n17431_, new_n17432_,
    new_n17433_, new_n17434_, new_n17435_, new_n17436_, new_n17437_,
    new_n17438_, new_n17439_, new_n17440_, new_n17441_, new_n17442_,
    new_n17443_, new_n17444_, new_n17445_, new_n17446_, new_n17447_,
    new_n17448_, new_n17449_, new_n17450_, new_n17451_, new_n17452_,
    new_n17453_, new_n17454_, new_n17455_, new_n17456_, new_n17457_,
    new_n17458_, new_n17459_, new_n17460_, new_n17461_, new_n17462_,
    new_n17463_, new_n17464_, new_n17465_, new_n17466_, new_n17467_,
    new_n17468_, new_n17469_, new_n17470_, new_n17471_, new_n17472_,
    new_n17473_, new_n17474_, new_n17475_, new_n17476_, new_n17477_,
    new_n17478_, new_n17479_, new_n17480_, new_n17481_, new_n17482_,
    new_n17483_, new_n17484_, new_n17485_, new_n17486_, new_n17487_,
    new_n17488_, new_n17489_, new_n17490_, new_n17491_, new_n17492_,
    new_n17493_, new_n17494_, new_n17495_, new_n17496_, new_n17497_,
    new_n17498_, new_n17499_, new_n17500_, new_n17501_, new_n17502_,
    new_n17503_, new_n17504_, new_n17505_, new_n17506_, new_n17507_,
    new_n17508_, new_n17509_, new_n17510_, new_n17511_, new_n17512_,
    new_n17513_, new_n17514_, new_n17515_, new_n17516_, new_n17517_,
    new_n17518_, new_n17519_, new_n17520_, new_n17521_, new_n17522_,
    new_n17523_, new_n17524_, new_n17525_, new_n17526_, new_n17527_,
    new_n17528_, new_n17529_, new_n17530_, new_n17531_, new_n17532_,
    new_n17533_, new_n17534_, new_n17535_, new_n17536_, new_n17537_,
    new_n17538_, new_n17539_, new_n17540_, new_n17541_, new_n17542_,
    new_n17543_, new_n17544_, new_n17545_, new_n17546_, new_n17547_,
    new_n17548_, new_n17549_, new_n17550_, new_n17551_, new_n17552_,
    new_n17553_, new_n17554_, new_n17555_, new_n17556_, new_n17557_,
    new_n17558_, new_n17559_, new_n17560_, new_n17561_, new_n17562_,
    new_n17563_, new_n17564_, new_n17565_, new_n17566_, new_n17567_,
    new_n17568_, new_n17569_, new_n17570_, new_n17571_, new_n17572_,
    new_n17573_, new_n17574_, new_n17575_, new_n17576_, new_n17577_,
    new_n17578_, new_n17579_, new_n17580_, new_n17581_, new_n17582_,
    new_n17583_, new_n17584_, new_n17585_, new_n17586_, new_n17587_,
    new_n17588_, new_n17589_, new_n17590_, new_n17591_, new_n17592_,
    new_n17593_, new_n17594_, new_n17595_, new_n17596_, new_n17597_,
    new_n17598_, new_n17599_, new_n17600_, new_n17601_, new_n17602_,
    new_n17603_, new_n17604_, new_n17605_, new_n17606_, new_n17607_,
    new_n17608_, new_n17609_, new_n17610_, new_n17611_, new_n17612_,
    new_n17613_, new_n17614_, new_n17615_, new_n17616_, new_n17617_,
    new_n17618_, new_n17619_, new_n17620_, new_n17621_, new_n17622_,
    new_n17623_, new_n17624_, new_n17625_, new_n17626_, new_n17627_,
    new_n17628_, new_n17629_, new_n17630_, new_n17631_, new_n17632_,
    new_n17633_, new_n17634_, new_n17635_, new_n17636_, new_n17637_,
    new_n17638_, new_n17639_, new_n17640_, new_n17641_, new_n17642_,
    new_n17643_, new_n17644_, new_n17645_, new_n17646_, new_n17647_,
    new_n17648_, new_n17649_, new_n17650_, new_n17651_, new_n17652_,
    new_n17654_, new_n17655_, new_n17656_, new_n17657_, new_n17658_,
    new_n17659_, new_n17660_, new_n17661_, new_n17662_, new_n17663_,
    new_n17664_, new_n17665_, new_n17666_, new_n17667_, new_n17668_,
    new_n17669_, new_n17670_, new_n17671_, new_n17672_, new_n17673_,
    new_n17674_, new_n17675_, new_n17676_, new_n17677_, new_n17678_,
    new_n17679_, new_n17680_, new_n17681_, new_n17682_, new_n17683_,
    new_n17684_, new_n17685_, new_n17686_, new_n17687_, new_n17688_,
    new_n17689_, new_n17690_, new_n17692_, new_n17693_, new_n17694_,
    new_n17695_, new_n17696_, new_n17697_, new_n17698_, new_n17699_,
    new_n17700_, new_n17701_, new_n17702_, new_n17703_, new_n17704_,
    new_n17705_, new_n17706_, new_n17707_, new_n17708_, new_n17709_,
    new_n17710_, new_n17711_, new_n17712_, new_n17713_, new_n17714_,
    new_n17715_, new_n17716_, new_n17717_, new_n17718_, new_n17719_,
    new_n17720_, new_n17721_, new_n17722_, new_n17723_, new_n17724_,
    new_n17725_, new_n17726_, new_n17727_, new_n17728_, new_n17729_,
    new_n17730_, new_n17731_, new_n17732_, new_n17733_, new_n17734_,
    new_n17735_, new_n17736_, new_n17737_, new_n17738_, new_n17739_,
    new_n17740_, new_n17741_, new_n17742_, new_n17743_, new_n17744_,
    new_n17745_, new_n17746_, new_n17747_, new_n17748_, new_n17749_,
    new_n17750_, new_n17751_, new_n17752_, new_n17753_, new_n17754_,
    new_n17755_, new_n17756_, new_n17757_, new_n17758_, new_n17759_,
    new_n17760_, new_n17761_, new_n17762_, new_n17763_, new_n17764_,
    new_n17765_, new_n17766_, new_n17767_, new_n17768_, new_n17769_,
    new_n17770_, new_n17771_, new_n17772_, new_n17773_, new_n17774_,
    new_n17775_, new_n17776_, new_n17777_, new_n17778_, new_n17779_,
    new_n17780_, new_n17781_, new_n17782_, new_n17783_, new_n17784_,
    new_n17785_, new_n17786_, new_n17787_, new_n17788_, new_n17789_,
    new_n17790_, new_n17791_, new_n17792_, new_n17793_, new_n17794_,
    new_n17795_, new_n17796_, new_n17797_, new_n17798_, new_n17799_,
    new_n17800_, new_n17801_, new_n17802_, new_n17803_, new_n17804_,
    new_n17805_, new_n17806_, new_n17807_, new_n17808_, new_n17809_,
    new_n17810_, new_n17811_, new_n17813_, new_n17814_, new_n17815_,
    new_n17816_, new_n17817_, new_n17818_, new_n17819_, new_n17820_,
    new_n17821_, new_n17822_, new_n17823_, new_n17826_, new_n17827_,
    new_n17828_, new_n17829_, new_n17830_, new_n17831_, new_n17832_,
    new_n17833_, new_n17834_, new_n17835_, new_n17836_, new_n17837_,
    new_n17838_, new_n17839_, new_n17840_, new_n17841_, new_n17842_,
    new_n17843_, new_n17844_, new_n17845_, new_n17846_, new_n17847_,
    new_n17848_, new_n17849_, new_n17850_, new_n17851_, new_n17852_,
    new_n17853_, new_n17854_, new_n17855_, new_n17856_, new_n17857_,
    new_n17858_, new_n17859_, new_n17860_, new_n17861_, new_n17862_,
    new_n17863_, new_n17864_, new_n17865_, new_n17866_, new_n17867_,
    new_n17868_, new_n17869_, new_n17870_, new_n17871_, new_n17872_,
    new_n17873_, new_n17874_, new_n17875_, new_n17876_, new_n17877_,
    new_n17878_, new_n17879_, new_n17880_, new_n17881_, new_n17882_,
    new_n17883_, new_n17884_, new_n17885_, new_n17886_, new_n17887_,
    new_n17888_, new_n17889_, new_n17890_, new_n17891_, new_n17892_,
    new_n17893_, new_n17894_, new_n17895_, new_n17896_, new_n17897_,
    new_n17898_, new_n17899_, new_n17900_, new_n17901_, new_n17902_,
    new_n17903_, new_n17904_, new_n17905_, new_n17906_, new_n17907_,
    new_n17908_, new_n17909_, new_n17910_, new_n17911_, new_n17912_,
    new_n17913_, new_n17914_, new_n17915_, new_n17916_, new_n17917_,
    new_n17918_, new_n17919_, new_n17920_, new_n17921_, new_n17922_,
    new_n17923_, new_n17924_, new_n17925_, new_n17926_, new_n17927_,
    new_n17928_, new_n17929_, new_n17930_, new_n17931_, new_n17932_,
    new_n17933_, new_n17934_, new_n17935_, new_n17936_, new_n17937_,
    new_n17938_, new_n17939_, new_n17940_, new_n17941_, new_n17942_,
    new_n17943_, new_n17944_, new_n17945_, new_n17946_, new_n17947_,
    new_n17948_, new_n17949_, new_n17950_, new_n17951_, new_n17952_,
    new_n17953_, new_n17954_, new_n17955_, new_n17956_, new_n17957_,
    new_n17958_, new_n17959_, new_n17960_, new_n17961_, new_n17962_,
    new_n17963_, new_n17964_, new_n17965_, new_n17966_, new_n17967_,
    new_n17968_, new_n17969_, new_n17970_, new_n17971_, new_n17972_,
    new_n17973_, new_n17974_, new_n17975_, new_n17976_, new_n17977_,
    new_n17978_, new_n17979_, new_n17980_, new_n17981_, new_n17982_,
    new_n17983_, new_n17984_, new_n17985_, new_n17986_, new_n17987_,
    new_n17988_, new_n17989_, new_n17990_, new_n17991_, new_n17992_,
    new_n17993_, new_n17994_, new_n17995_, new_n17996_, new_n17997_,
    new_n17998_, new_n17999_, new_n18000_, new_n18001_, new_n18002_,
    new_n18003_, new_n18005_, new_n18006_, new_n18007_, new_n18008_,
    new_n18009_, new_n18010_, new_n18011_, new_n18012_, new_n18013_,
    new_n18014_, new_n18015_, new_n18016_, new_n18017_, new_n18018_,
    new_n18019_, new_n18020_, new_n18021_, new_n18022_, new_n18023_,
    new_n18024_, new_n18025_, new_n18026_, new_n18027_, new_n18028_,
    new_n18029_, new_n18030_, new_n18031_, new_n18032_, new_n18033_,
    new_n18034_, new_n18035_, new_n18036_, new_n18037_, new_n18038_,
    new_n18039_, new_n18041_, new_n18042_, new_n18043_, new_n18044_,
    new_n18045_, new_n18046_, new_n18047_, new_n18048_, new_n18049_,
    new_n18050_, new_n18051_, new_n18052_, new_n18053_, new_n18054_,
    new_n18055_, new_n18056_, new_n18057_, new_n18058_, new_n18059_,
    new_n18060_, new_n18061_, new_n18062_, new_n18063_, new_n18064_,
    new_n18065_, new_n18066_, new_n18067_, new_n18068_, new_n18069_,
    new_n18070_, new_n18071_, new_n18072_, new_n18073_, new_n18074_,
    new_n18075_, new_n18076_, new_n18077_, new_n18078_, new_n18079_,
    new_n18080_, new_n18081_, new_n18082_, new_n18083_, new_n18084_,
    new_n18085_, new_n18086_, new_n18087_, new_n18088_, new_n18089_,
    new_n18090_, new_n18091_, new_n18092_, new_n18093_, new_n18094_,
    new_n18095_, new_n18096_, new_n18097_, new_n18098_, new_n18099_,
    new_n18100_, new_n18101_, new_n18102_, new_n18103_, new_n18104_,
    new_n18105_, new_n18106_, new_n18107_, new_n18108_, new_n18109_,
    new_n18110_, new_n18111_, new_n18112_, new_n18113_, new_n18114_,
    new_n18115_, new_n18116_, new_n18117_, new_n18118_, new_n18119_,
    new_n18120_, new_n18121_, new_n18122_, new_n18123_, new_n18124_,
    new_n18125_, new_n18126_, new_n18127_, new_n18128_, new_n18129_,
    new_n18130_, new_n18131_, new_n18132_, new_n18133_, new_n18134_,
    new_n18135_, new_n18136_, new_n18137_, new_n18138_, new_n18139_,
    new_n18140_, new_n18141_, new_n18142_, new_n18143_, new_n18144_,
    new_n18145_, new_n18146_, new_n18147_, new_n18148_, new_n18149_,
    new_n18150_, new_n18151_, new_n18152_, new_n18153_, new_n18154_,
    new_n18155_, new_n18156_, new_n18157_, new_n18158_, new_n18159_,
    new_n18160_, new_n18161_, new_n18162_, new_n18163_, new_n18164_,
    new_n18165_, new_n18166_, new_n18167_, new_n18168_, new_n18169_,
    new_n18170_, new_n18171_, new_n18172_, new_n18173_, new_n18174_,
    new_n18175_, new_n18176_, new_n18177_, new_n18178_, new_n18179_,
    new_n18180_, new_n18181_, new_n18182_, new_n18183_, new_n18184_,
    new_n18185_, new_n18186_, new_n18187_, new_n18188_, new_n18189_,
    new_n18190_, new_n18191_, new_n18192_, new_n18193_, new_n18194_,
    new_n18195_, new_n18196_, new_n18197_, new_n18198_, new_n18199_,
    new_n18200_, new_n18201_, new_n18202_, new_n18203_, new_n18204_,
    new_n18205_, new_n18206_, new_n18207_, new_n18217_, new_n18218_,
    new_n18219_, new_n18220_, new_n18221_, new_n18222_, new_n18223_,
    new_n18224_, new_n18225_, new_n18226_, new_n18227_, new_n18228_,
    new_n18229_, new_n18230_, new_n18231_, new_n18232_, new_n18233_,
    new_n18234_, new_n18235_, new_n18236_, new_n18237_, new_n18238_,
    new_n18239_, new_n18240_, new_n18241_, new_n18242_, new_n18243_,
    new_n18244_, new_n18245_, new_n18246_, new_n18247_, new_n18248_,
    new_n18249_, new_n18250_, new_n18251_, new_n18252_, new_n18253_,
    new_n18254_, new_n18255_, new_n18256_, new_n18257_, new_n18258_,
    new_n18259_, new_n18260_, new_n18261_, new_n18262_, new_n18263_,
    new_n18264_, new_n18265_, new_n18266_, new_n18267_, new_n18268_,
    new_n18269_, new_n18270_, new_n18271_, new_n18272_, new_n18273_,
    new_n18274_, new_n18276_, new_n18277_, new_n18278_, new_n18279_,
    new_n18280_, new_n18281_, new_n18282_, new_n18283_, new_n18284_,
    new_n18285_, new_n18286_, new_n18287_, new_n18288_, new_n18289_,
    new_n18290_, new_n18291_, new_n18292_, new_n18293_, new_n18294_,
    new_n18295_, new_n18296_, new_n18297_, new_n18298_, new_n18299_,
    new_n18300_, new_n18301_, new_n18302_, new_n18303_, new_n18304_,
    new_n18305_, new_n18306_, new_n18307_, new_n18308_, new_n18309_,
    new_n18310_, new_n18311_, new_n18312_, new_n18314_, new_n18315_,
    new_n18316_, new_n18317_, new_n18318_, new_n18319_, new_n18320_,
    new_n18321_, new_n18322_, new_n18323_, new_n18324_, new_n18325_,
    new_n18326_, new_n18327_, new_n18328_, new_n18329_, new_n18330_,
    new_n18331_, new_n18332_, new_n18333_, new_n18334_, new_n18335_,
    new_n18336_, new_n18337_, new_n18338_, new_n18339_, new_n18340_,
    new_n18341_, new_n18342_, new_n18343_, new_n18344_, new_n18345_,
    new_n18346_, new_n18347_, new_n18348_, new_n18349_, new_n18350_,
    new_n18351_, new_n18352_, new_n18353_, new_n18354_, new_n18355_,
    new_n18356_, new_n18357_, new_n18358_, new_n18359_, new_n18360_,
    new_n18361_, new_n18362_, new_n18363_, new_n18364_, new_n18365_,
    new_n18366_, new_n18367_, new_n18368_, new_n18369_, new_n18370_,
    new_n18371_, new_n18372_, new_n18373_, new_n18374_, new_n18375_,
    new_n18376_, new_n18377_, new_n18378_, new_n18379_, new_n18380_,
    new_n18381_, new_n18382_, new_n18383_, new_n18384_, new_n18385_,
    new_n18386_, new_n18387_, new_n18388_, new_n18389_, new_n18390_,
    new_n18391_, new_n18392_, new_n18393_, new_n18394_, new_n18395_,
    new_n18396_, new_n18397_, new_n18398_, new_n18399_, new_n18400_,
    new_n18401_, new_n18402_, new_n18403_, new_n18404_, new_n18405_,
    new_n18410_, new_n18411_, new_n18412_, new_n18413_, new_n18414_,
    new_n18415_, new_n18416_, new_n18417_, new_n18418_, new_n18419_,
    new_n18420_, new_n18421_, new_n18422_, new_n18423_, new_n18424_,
    new_n18425_, new_n18427_, new_n18428_, new_n18429_, new_n18430_,
    new_n18431_, new_n18432_, new_n18433_, new_n18434_, new_n18435_,
    new_n18436_, new_n18437_, new_n18438_, new_n18439_, new_n18440_,
    new_n18441_, new_n18442_, new_n18443_, new_n18444_, new_n18445_,
    new_n18446_, new_n18447_, new_n18448_, new_n18449_, new_n18450_,
    new_n18451_, new_n18452_, new_n18453_, new_n18454_, new_n18455_,
    new_n18456_, new_n18457_, new_n18458_, new_n18459_, new_n18460_,
    new_n18461_, new_n18462_, new_n18463_, new_n18464_, new_n18465_,
    new_n18466_, new_n18467_, new_n18468_, new_n18469_, new_n18470_,
    new_n18471_, new_n18472_, new_n18473_, new_n18474_, new_n18475_,
    new_n18476_, new_n18477_, new_n18478_, new_n18479_, new_n18480_,
    new_n18481_, new_n18482_, new_n18483_, new_n18484_, new_n18485_,
    new_n18486_, new_n18487_, new_n18488_, new_n18489_, new_n18490_,
    new_n18491_, new_n18492_, new_n18493_, new_n18494_, new_n18495_,
    new_n18496_, new_n18497_, new_n18498_, new_n18499_, new_n18500_,
    new_n18501_, new_n18502_, new_n18503_, new_n18504_, new_n18505_,
    new_n18506_, new_n18507_, new_n18508_, new_n18509_, new_n18510_,
    new_n18511_, new_n18512_, new_n18513_, new_n18514_, new_n18515_,
    new_n18516_, new_n18517_, new_n18518_, new_n18519_, new_n18520_,
    new_n18521_, new_n18522_, new_n18523_, new_n18524_, new_n18525_,
    new_n18526_, new_n18527_, new_n18528_, new_n18529_, new_n18530_,
    new_n18531_, new_n18532_, new_n18533_, new_n18534_, new_n18535_,
    new_n18536_, new_n18537_, new_n18538_, new_n18539_, new_n18540_,
    new_n18541_, new_n18542_, new_n18543_, new_n18544_, new_n18545_,
    new_n18546_, new_n18547_, new_n18548_, new_n18549_, new_n18550_,
    new_n18551_, new_n18552_, new_n18553_, new_n18554_, new_n18555_,
    new_n18556_, new_n18557_, new_n18558_, new_n18559_, new_n18560_,
    new_n18561_, new_n18562_, new_n18563_, new_n18564_, new_n18565_,
    new_n18566_, new_n18567_, new_n18568_, new_n18569_, new_n18570_,
    new_n18571_, new_n18572_, new_n18573_, new_n18574_, new_n18575_,
    new_n18576_, new_n18577_, new_n18578_, new_n18579_, new_n18580_,
    new_n18581_, new_n18582_, new_n18583_, new_n18584_, new_n18585_,
    new_n18586_, new_n18587_, new_n18588_, new_n18589_, new_n18590_,
    new_n18591_, new_n18592_, new_n18594_, new_n18595_, new_n18596_,
    new_n18597_, new_n18598_, new_n18599_, new_n18600_, new_n18601_,
    new_n18602_, new_n18603_, new_n18604_, new_n18605_, new_n18606_,
    new_n18607_, new_n18608_, new_n18609_, new_n18610_, new_n18611_,
    new_n18612_, new_n18613_, new_n18614_, new_n18615_, new_n18616_,
    new_n18617_, new_n18618_, new_n18619_, new_n18620_, new_n18621_,
    new_n18622_, new_n18623_, new_n18624_, new_n18625_, new_n18626_,
    new_n18627_, new_n18628_, new_n18630_, new_n18631_, new_n18632_,
    new_n18633_, new_n18634_, new_n18635_, new_n18636_, new_n18637_,
    new_n18638_, new_n18639_, new_n18640_, new_n18641_, new_n18642_,
    new_n18643_, new_n18644_, new_n18645_, new_n18646_, new_n18647_,
    new_n18648_, new_n18649_, new_n18650_, new_n18651_, new_n18652_,
    new_n18653_, new_n18654_, new_n18655_, new_n18656_, new_n18657_,
    new_n18658_, new_n18659_, new_n18660_, new_n18661_, new_n18662_,
    new_n18663_, new_n18664_, new_n18665_, new_n18666_, new_n18667_,
    new_n18668_, new_n18669_, new_n18670_, new_n18671_, new_n18672_,
    new_n18673_, new_n18674_, new_n18675_, new_n18676_, new_n18677_,
    new_n18678_, new_n18679_, new_n18680_, new_n18681_, new_n18682_,
    new_n18683_, new_n18684_, new_n18685_, new_n18686_, new_n18687_,
    new_n18688_, new_n18689_, new_n18690_, new_n18691_, new_n18692_,
    new_n18693_, new_n18694_, new_n18695_, new_n18696_, new_n18697_,
    new_n18698_, new_n18699_, new_n18700_, new_n18701_, new_n18702_,
    new_n18703_, new_n18704_, new_n18705_, new_n18706_, new_n18707_,
    new_n18708_, new_n18709_, new_n18710_, new_n18711_, new_n18712_,
    new_n18713_, new_n18714_, new_n18715_, new_n18716_, new_n18717_,
    new_n18720_, new_n18721_, new_n18722_, new_n18723_, new_n18724_,
    new_n18725_, new_n18726_, new_n18727_, new_n18728_, new_n18729_,
    new_n18730_, new_n18731_, new_n18732_, new_n18733_, new_n18734_,
    new_n18735_, new_n18736_, new_n18737_, new_n18738_, new_n18739_,
    new_n18740_, new_n18741_, new_n18742_, new_n18743_, new_n18744_,
    new_n18745_, new_n18746_, new_n18747_, new_n18748_, new_n18749_,
    new_n18750_, new_n18751_, new_n18752_, new_n18753_, new_n18754_,
    new_n18755_, new_n18756_, new_n18757_, new_n18758_, new_n18759_,
    new_n18760_, new_n18761_, new_n18762_, new_n18763_, new_n18764_,
    new_n18765_, new_n18766_, new_n18767_, new_n18768_, new_n18769_,
    new_n18770_, new_n18771_, new_n18772_, new_n18773_, new_n18774_,
    new_n18775_, new_n18776_, new_n18777_, new_n18778_, new_n18779_,
    new_n18780_, new_n18781_, new_n18782_, new_n18783_, new_n18784_,
    new_n18785_, new_n18786_, new_n18787_, new_n18788_, new_n18789_,
    new_n18790_, new_n18791_, new_n18792_, new_n18793_, new_n18803_,
    new_n18804_, new_n18805_, new_n18806_, new_n18807_, new_n18808_,
    new_n18809_, new_n18810_, new_n18811_, new_n18812_, new_n18813_,
    new_n18814_, new_n18815_, new_n18816_, new_n18817_, new_n18818_,
    new_n18819_, new_n18820_, new_n18821_, new_n18822_, new_n18823_,
    new_n18824_, new_n18825_, new_n18826_, new_n18827_, new_n18828_,
    new_n18829_, new_n18830_, new_n18831_, new_n18832_, new_n18833_,
    new_n18834_, new_n18835_, new_n18836_, new_n18837_, new_n18838_,
    new_n18839_, new_n18840_, new_n18841_, new_n18842_, new_n18843_,
    new_n18844_, new_n18845_, new_n18846_, new_n18847_, new_n18848_,
    new_n18849_, new_n18850_, new_n18851_, new_n18852_, new_n18853_,
    new_n18854_, new_n18855_, new_n18856_, new_n18857_, new_n18858_,
    new_n18859_, new_n18860_, new_n18861_, new_n18862_, new_n18863_,
    new_n18864_, new_n18865_, new_n18866_, new_n18868_, new_n18869_,
    new_n18870_, new_n18871_, new_n18872_, new_n18873_, new_n18874_,
    new_n18875_, new_n18876_, new_n18877_, new_n18878_, new_n18879_,
    new_n18880_, new_n18881_, new_n18882_, new_n18883_, new_n18884_,
    new_n18885_, new_n18886_, new_n18887_, new_n18888_, new_n18889_,
    new_n18890_, new_n18891_, new_n18892_, new_n18893_, new_n18894_,
    new_n18895_, new_n18896_, new_n18897_, new_n18898_, new_n18899_,
    new_n18900_, new_n18901_, new_n18902_, new_n18904_, new_n18905_,
    new_n18906_, new_n18907_, new_n18908_, new_n18909_, new_n18910_,
    new_n18911_, new_n18912_, new_n18913_, new_n18914_, new_n18915_,
    new_n18916_, new_n18917_, new_n18918_, new_n18919_, new_n18920_,
    new_n18921_, new_n18922_, new_n18923_, new_n18924_, new_n18925_,
    new_n18926_, new_n18927_, new_n18928_, new_n18929_, new_n18930_,
    new_n18931_, new_n18932_, new_n18933_, new_n18934_, new_n18935_,
    new_n18936_, new_n18937_, new_n18938_, new_n18939_, new_n18940_,
    new_n18941_, new_n18942_, new_n18943_, new_n18944_, new_n18945_,
    new_n18946_, new_n18947_, new_n18948_, new_n18949_, new_n18950_,
    new_n18951_, new_n18952_, new_n18953_, new_n18954_, new_n18955_,
    new_n18956_, new_n18957_, new_n18958_, new_n18959_, new_n18960_,
    new_n18961_, new_n18962_, new_n18963_, new_n18964_, new_n18965_,
    new_n18966_, new_n18967_, new_n18968_, new_n18969_, new_n18970_,
    new_n18971_, new_n18972_, new_n18973_, new_n18974_, new_n18975_,
    new_n18976_, new_n18977_, new_n18978_, new_n18979_, new_n18980_,
    new_n18981_, new_n18982_, new_n18983_, new_n18984_, new_n18985_,
    new_n18986_, new_n18987_, new_n18988_, new_n18989_, new_n18990_,
    new_n18991_, new_n18994_, new_n18995_, new_n18996_, new_n18997_,
    new_n18998_, new_n18999_, new_n19000_, new_n19001_, new_n19002_,
    new_n19003_, new_n19004_, new_n19005_, new_n19006_, new_n19007_,
    new_n19008_, new_n19009_, new_n19010_, new_n19011_, new_n19012_,
    new_n19013_, new_n19014_, new_n19015_, new_n19016_, new_n19017_,
    new_n19018_, new_n19019_, new_n19020_, new_n19021_, new_n19022_,
    new_n19023_, new_n19024_, new_n19025_, new_n19026_, new_n19027_,
    new_n19028_, new_n19029_, new_n19030_, new_n19031_, new_n19032_,
    new_n19033_, new_n19034_, new_n19035_, new_n19036_, new_n19037_,
    new_n19038_, new_n19039_, new_n19040_, new_n19041_, new_n19042_,
    new_n19043_, new_n19044_, new_n19045_, new_n19046_, new_n19047_,
    new_n19048_, new_n19049_, new_n19050_, new_n19051_, new_n19052_,
    new_n19053_, new_n19054_, new_n19055_, new_n19056_, new_n19057_,
    new_n19058_, new_n19059_, new_n19060_, new_n19061_, new_n19062_,
    new_n19063_, new_n19064_, new_n19065_, new_n19066_, new_n19067_,
    new_n19077_, new_n19078_, new_n19079_, new_n19080_, new_n19081_,
    new_n19082_, new_n19083_, new_n19084_, new_n19085_, new_n19086_,
    new_n19087_, new_n19088_, new_n19089_, new_n19090_, new_n19091_,
    new_n19092_, new_n19093_, new_n19094_, new_n19095_, new_n19096_,
    new_n19097_, new_n19098_, new_n19099_, new_n19100_, new_n19101_,
    new_n19102_, new_n19103_, new_n19104_, new_n19105_, new_n19106_,
    new_n19107_, new_n19108_, new_n19109_, new_n19110_, new_n19111_,
    new_n19112_, new_n19113_, new_n19114_, new_n19115_, new_n19116_,
    new_n19117_, new_n19118_, new_n19119_, new_n19120_, new_n19121_,
    new_n19122_, new_n19123_, new_n19124_, new_n19125_, new_n19126_,
    new_n19127_, new_n19128_, new_n19129_, new_n19130_, new_n19131_,
    new_n19132_, new_n19133_, new_n19134_, new_n19135_, new_n19136_,
    new_n19137_, new_n19138_, new_n19139_, new_n19141_, new_n19142_,
    new_n19143_, new_n19144_, new_n19145_, new_n19146_, new_n19147_,
    new_n19148_, new_n19149_, new_n19150_, new_n19151_, new_n19152_,
    new_n19153_, new_n19154_, new_n19155_, new_n19156_, new_n19157_,
    new_n19158_, new_n19159_, new_n19160_, new_n19161_, new_n19162_,
    new_n19163_, new_n19164_, new_n19165_, new_n19166_, new_n19167_,
    new_n19168_, new_n19169_, new_n19170_, new_n19171_, new_n19172_,
    new_n19173_, new_n19174_, new_n19175_, new_n19177_, new_n19178_,
    new_n19179_, new_n19180_, new_n19181_, new_n19182_, new_n19183_,
    new_n19184_, new_n19185_, new_n19186_, new_n19187_, new_n19188_,
    new_n19189_, new_n19190_, new_n19191_, new_n19192_, new_n19193_,
    new_n19194_, new_n19195_, new_n19196_, new_n19197_, new_n19198_,
    new_n19199_, new_n19200_, new_n19201_, new_n19202_, new_n19203_,
    new_n19204_, new_n19205_, new_n19206_, new_n19207_, new_n19208_,
    new_n19209_, new_n19210_, new_n19211_, new_n19212_, new_n19213_,
    new_n19214_, new_n19215_, new_n19216_, new_n19217_, new_n19218_,
    new_n19219_, new_n19220_, new_n19221_, new_n19222_, new_n19223_,
    new_n19224_, new_n19225_, new_n19226_, new_n19227_, new_n19228_,
    new_n19229_, new_n19230_, new_n19231_, new_n19232_, new_n19233_,
    new_n19234_, new_n19235_, new_n19236_, new_n19237_, new_n19238_,
    new_n19239_, new_n19240_, new_n19241_, new_n19242_, new_n19243_,
    new_n19244_, new_n19245_, new_n19246_, new_n19247_, new_n19248_,
    new_n19249_, new_n19250_, new_n19251_, new_n19252_, new_n19253_,
    new_n19254_, new_n19255_, new_n19256_, new_n19257_, new_n19258_,
    new_n19259_, new_n19260_, new_n19261_, new_n19262_, new_n19263_,
    new_n19264_, new_n19265_, new_n19266_, new_n19267_, new_n19268_,
    new_n19269_, new_n19270_, new_n19271_, new_n19272_, new_n19273_,
    new_n19274_, new_n19275_, new_n19276_, new_n19277_, new_n19278_,
    new_n19279_, new_n19280_, new_n19281_, new_n19282_, new_n19283_,
    new_n19284_, new_n19285_, new_n19286_, new_n19287_, new_n19288_,
    new_n19289_, new_n19290_, new_n19291_, new_n19292_, new_n19293_,
    new_n19294_, new_n19295_, new_n19296_, new_n19297_, new_n19298_,
    new_n19299_, new_n19300_, new_n19301_, new_n19302_, new_n19303_,
    new_n19304_, new_n19305_, new_n19306_, new_n19307_, new_n19308_,
    new_n19309_, new_n19310_, new_n19311_, new_n19312_, new_n19313_,
    new_n19314_, new_n19315_, new_n19316_, new_n19317_, new_n19318_,
    new_n19319_, new_n19320_, new_n19321_, new_n19322_, new_n19323_,
    new_n19324_, new_n19325_, new_n19326_, new_n19327_, new_n19328_,
    new_n19329_, new_n19330_, new_n19331_, new_n19332_, new_n19333_,
    new_n19334_, new_n19335_, new_n19336_, new_n19337_, new_n19338_,
    new_n19339_, new_n19340_, new_n19341_, new_n19342_, new_n19343_,
    new_n19353_, new_n19354_, new_n19355_, new_n19356_, new_n19357_,
    new_n19358_, new_n19359_, new_n19360_, new_n19361_, new_n19362_,
    new_n19363_, new_n19364_, new_n19365_, new_n19366_, new_n19367_,
    new_n19368_, new_n19369_, new_n19370_, new_n19371_, new_n19372_,
    new_n19373_, new_n19374_, new_n19375_, new_n19376_, new_n19377_,
    new_n19378_, new_n19379_, new_n19380_, new_n19381_, new_n19382_,
    new_n19383_, new_n19384_, new_n19385_, new_n19386_, new_n19387_,
    new_n19388_, new_n19389_, new_n19390_, new_n19391_, new_n19392_,
    new_n19393_, new_n19394_, new_n19395_, new_n19396_, new_n19397_,
    new_n19398_, new_n19399_, new_n19400_, new_n19401_, new_n19402_,
    new_n19403_, new_n19404_, new_n19405_, new_n19406_, new_n19407_,
    new_n19408_, new_n19409_, new_n19410_, new_n19412_, new_n19413_,
    new_n19414_, new_n19415_, new_n19416_, new_n19417_, new_n19418_,
    new_n19419_, new_n19420_, new_n19421_, new_n19422_, new_n19423_,
    new_n19424_, new_n19425_, new_n19426_, new_n19427_, new_n19428_,
    new_n19429_, new_n19430_, new_n19431_, new_n19432_, new_n19433_,
    new_n19434_, new_n19435_, new_n19436_, new_n19437_, new_n19438_,
    new_n19439_, new_n19440_, new_n19441_, new_n19442_, new_n19443_,
    new_n19444_, new_n19445_, new_n19446_, new_n19448_, new_n19449_,
    new_n19450_, new_n19451_, new_n19452_, new_n19453_, new_n19454_,
    new_n19455_, new_n19456_, new_n19457_, new_n19458_, new_n19459_,
    new_n19460_, new_n19461_, new_n19462_, new_n19463_, new_n19464_,
    new_n19465_, new_n19466_, new_n19467_, new_n19468_, new_n19469_,
    new_n19470_, new_n19471_, new_n19472_, new_n19473_, new_n19474_,
    new_n19475_, new_n19476_, new_n19477_, new_n19478_, new_n19479_,
    new_n19480_, new_n19481_, new_n19482_, new_n19483_, new_n19484_,
    new_n19485_, new_n19486_, new_n19487_, new_n19488_, new_n19489_,
    new_n19490_, new_n19491_, new_n19492_, new_n19493_, new_n19494_,
    new_n19495_, new_n19496_, new_n19497_, new_n19498_, new_n19499_,
    new_n19500_, new_n19501_, new_n19502_, new_n19503_, new_n19504_,
    new_n19505_, new_n19506_, new_n19507_, new_n19508_, new_n19509_,
    new_n19510_, new_n19511_, new_n19512_, new_n19513_, new_n19514_,
    new_n19515_, new_n19516_, new_n19517_, new_n19518_, new_n19519_,
    new_n19520_, new_n19521_, new_n19522_, new_n19523_, new_n19524_,
    new_n19525_, new_n19526_, new_n19527_, new_n19528_, new_n19529_,
    new_n19530_, new_n19531_, new_n19532_, new_n19533_, new_n19534_,
    new_n19535_, new_n19536_, new_n19537_, new_n19538_, new_n19539_,
    new_n19540_, new_n19541_, new_n19542_, new_n19543_, new_n19544_,
    new_n19545_, new_n19546_, new_n19547_, new_n19548_, new_n19549_,
    new_n19550_, new_n19551_, new_n19552_, new_n19553_, new_n19554_,
    new_n19555_, new_n19556_, new_n19557_, new_n19558_, new_n19559_,
    new_n19560_, new_n19561_, new_n19562_, new_n19563_, new_n19564_,
    new_n19565_, new_n19566_, new_n19567_, new_n19568_, new_n19569_,
    new_n19570_, new_n19571_, new_n19572_, new_n19573_, new_n19574_,
    new_n19575_, new_n19576_, new_n19577_, new_n19578_, new_n19579_,
    new_n19580_, new_n19581_, new_n19582_, new_n19583_, new_n19584_,
    new_n19585_, new_n19586_, new_n19587_, new_n19588_, new_n19589_,
    new_n19590_, new_n19591_, new_n19592_, new_n19593_, new_n19594_,
    new_n19595_, new_n19596_, new_n19597_, new_n19598_, new_n19599_,
    new_n19600_, new_n19601_, new_n19602_, new_n19603_, new_n19604_,
    new_n19605_, new_n19606_, new_n19607_, new_n19608_, new_n19609_,
    new_n19610_, new_n19611_, new_n19612_, new_n19613_, new_n19614_,
    new_n19624_, new_n19625_, new_n19626_, new_n19627_, new_n19628_,
    new_n19629_, new_n19630_, new_n19631_, new_n19632_, new_n19633_,
    new_n19634_, new_n19635_, new_n19636_, new_n19637_, new_n19638_,
    new_n19639_, new_n19640_, new_n19641_, new_n19642_, new_n19643_,
    new_n19644_, new_n19645_, new_n19646_, new_n19647_, new_n19648_,
    new_n19649_, new_n19650_, new_n19651_, new_n19652_, new_n19653_,
    new_n19654_, new_n19655_, new_n19656_, new_n19657_, new_n19658_,
    new_n19659_, new_n19660_, new_n19661_, new_n19662_, new_n19663_,
    new_n19664_, new_n19665_, new_n19666_, new_n19667_, new_n19668_,
    new_n19669_, new_n19670_, new_n19671_, new_n19672_, new_n19673_,
    new_n19674_, new_n19675_, new_n19676_, new_n19677_, new_n19678_,
    new_n19679_, new_n19680_, new_n19681_, new_n19683_, new_n19684_,
    new_n19685_, new_n19686_, new_n19687_, new_n19688_, new_n19689_,
    new_n19690_, new_n19691_, new_n19692_, new_n19693_, new_n19694_,
    new_n19695_, new_n19696_, new_n19697_, new_n19698_, new_n19699_,
    new_n19700_, new_n19701_, new_n19702_, new_n19703_, new_n19704_,
    new_n19705_, new_n19706_, new_n19707_, new_n19708_, new_n19709_,
    new_n19710_, new_n19711_, new_n19712_, new_n19713_, new_n19714_,
    new_n19715_, new_n19716_, new_n19717_, new_n19719_, new_n19720_,
    new_n19721_, new_n19722_, new_n19723_, new_n19724_, new_n19725_,
    new_n19726_, new_n19727_, new_n19728_, new_n19729_, new_n19730_,
    new_n19731_, new_n19732_, new_n19733_, new_n19734_, new_n19735_,
    new_n19736_, new_n19737_, new_n19738_, new_n19739_, new_n19740_,
    new_n19741_, new_n19742_, new_n19743_, new_n19744_, new_n19745_,
    new_n19746_, new_n19747_, new_n19748_, new_n19749_, new_n19750_,
    new_n19751_, new_n19752_, new_n19753_, new_n19754_, new_n19755_,
    new_n19756_, new_n19757_, new_n19758_, new_n19759_, new_n19760_,
    new_n19761_, new_n19762_, new_n19763_, new_n19764_, new_n19765_,
    new_n19766_, new_n19767_, new_n19768_, new_n19769_, new_n19770_,
    new_n19771_, new_n19772_, new_n19773_, new_n19774_, new_n19775_,
    new_n19776_, new_n19777_, new_n19778_, new_n19779_, new_n19780_,
    new_n19781_, new_n19782_, new_n19783_, new_n19784_, new_n19785_,
    new_n19786_, new_n19787_, new_n19788_, new_n19789_, new_n19790_,
    new_n19791_, new_n19792_, new_n19793_, new_n19794_, new_n19795_,
    new_n19796_, new_n19797_, new_n19798_, new_n19799_, new_n19800_,
    new_n19801_, new_n19802_, new_n19803_, new_n19804_, new_n19805_,
    new_n19806_, new_n19807_, new_n19808_, new_n19809_, new_n19810_,
    new_n19811_, new_n19812_, new_n19813_, new_n19814_, new_n19815_,
    new_n19816_, new_n19817_, new_n19818_, new_n19819_, new_n19820_,
    new_n19821_, new_n19822_, new_n19823_, new_n19824_, new_n19825_,
    new_n19826_, new_n19827_, new_n19828_, new_n19829_, new_n19830_,
    new_n19831_, new_n19832_, new_n19833_, new_n19834_, new_n19835_,
    new_n19836_, new_n19837_, new_n19838_, new_n19839_, new_n19840_,
    new_n19841_, new_n19842_, new_n19843_, new_n19844_, new_n19845_,
    new_n19846_, new_n19847_, new_n19848_, new_n19849_, new_n19850_,
    new_n19851_, new_n19852_, new_n19853_, new_n19854_, new_n19855_,
    new_n19856_, new_n19857_, new_n19858_, new_n19859_, new_n19860_,
    new_n19861_, new_n19862_, new_n19863_, new_n19864_, new_n19865_,
    new_n19866_, new_n19867_, new_n19868_, new_n19869_, new_n19870_,
    new_n19871_, new_n19872_, new_n19873_, new_n19874_, new_n19875_,
    new_n19876_, new_n19877_, new_n19878_, new_n19879_, new_n19880_,
    new_n19881_, new_n19882_, new_n19883_, new_n19884_, new_n19885_,
    new_n19895_, new_n19896_, new_n19897_, new_n19898_, new_n19899_,
    new_n19900_, new_n19901_, new_n19902_, new_n19903_, new_n19904_,
    new_n19905_, new_n19906_, new_n19907_, new_n19908_, new_n19909_,
    new_n19910_, new_n19911_, new_n19912_, new_n19913_, new_n19914_,
    new_n19915_, new_n19916_, new_n19917_, new_n19918_, new_n19919_,
    new_n19920_, new_n19921_, new_n19922_, new_n19923_, new_n19924_,
    new_n19925_, new_n19926_, new_n19927_, new_n19928_, new_n19929_,
    new_n19930_, new_n19931_, new_n19932_, new_n19933_, new_n19934_,
    new_n19935_, new_n19936_, new_n19937_, new_n19938_, new_n19939_,
    new_n19940_, new_n19941_, new_n19942_, new_n19943_, new_n19944_,
    new_n19945_, new_n19946_, new_n19947_, new_n19948_, new_n19949_,
    new_n19950_, new_n19951_, new_n19952_, new_n19954_, new_n19955_,
    new_n19956_, new_n19957_, new_n19958_, new_n19959_, new_n19960_,
    new_n19961_, new_n19962_, new_n19963_, new_n19964_, new_n19965_,
    new_n19966_, new_n19967_, new_n19968_, new_n19969_, new_n19970_,
    new_n19971_, new_n19972_, new_n19973_, new_n19974_, new_n19975_,
    new_n19976_, new_n19977_, new_n19978_, new_n19979_, new_n19980_,
    new_n19981_, new_n19982_, new_n19983_, new_n19984_, new_n19985_,
    new_n19986_, new_n19987_, new_n19988_, new_n19990_, new_n19991_,
    new_n19992_, new_n19993_, new_n19994_, new_n19995_, new_n19996_,
    new_n19997_, new_n19998_, new_n19999_, new_n20000_, new_n20001_,
    new_n20002_, new_n20003_, new_n20004_, new_n20005_, new_n20006_,
    new_n20007_, new_n20008_, new_n20009_, new_n20010_, new_n20011_,
    new_n20012_, new_n20013_, new_n20014_, new_n20015_, new_n20016_,
    new_n20017_, new_n20018_, new_n20019_, new_n20020_, new_n20021_,
    new_n20022_, new_n20023_, new_n20024_, new_n20025_, new_n20026_,
    new_n20027_, new_n20028_, new_n20029_, new_n20030_, new_n20031_,
    new_n20032_, new_n20033_, new_n20034_, new_n20035_, new_n20036_,
    new_n20037_, new_n20038_, new_n20039_, new_n20040_, new_n20041_,
    new_n20042_, new_n20043_, new_n20044_, new_n20045_, new_n20046_,
    new_n20047_, new_n20048_, new_n20049_, new_n20050_, new_n20051_,
    new_n20052_, new_n20053_, new_n20054_, new_n20055_, new_n20056_,
    new_n20057_, new_n20058_, new_n20059_, new_n20060_, new_n20061_,
    new_n20062_, new_n20063_, new_n20064_, new_n20065_, new_n20066_,
    new_n20067_, new_n20068_, new_n20069_, new_n20070_, new_n20071_,
    new_n20072_, new_n20073_, new_n20074_, new_n20075_, new_n20076_,
    new_n20077_, new_n20080_, new_n20081_, new_n20082_, new_n20083_,
    new_n20084_, new_n20085_, new_n20086_, new_n20087_, new_n20088_,
    new_n20089_, new_n20090_, new_n20091_, new_n20092_, new_n20093_,
    new_n20094_, new_n20095_, new_n20096_, new_n20097_, new_n20098_,
    new_n20099_, new_n20100_, new_n20101_, new_n20102_, new_n20103_,
    new_n20104_, new_n20105_, new_n20106_, new_n20107_, new_n20108_,
    new_n20109_, new_n20110_, new_n20111_, new_n20112_, new_n20113_,
    new_n20114_, new_n20115_, new_n20116_, new_n20117_, new_n20118_,
    new_n20119_, new_n20120_, new_n20121_, new_n20122_, new_n20123_,
    new_n20124_, new_n20125_, new_n20126_, new_n20127_, new_n20128_,
    new_n20129_, new_n20130_, new_n20131_, new_n20132_, new_n20133_,
    new_n20134_, new_n20135_, new_n20136_, new_n20137_, new_n20138_,
    new_n20139_, new_n20140_, new_n20141_, new_n20142_, new_n20143_,
    new_n20144_, new_n20145_, new_n20146_, new_n20147_, new_n20148_,
    new_n20149_, new_n20150_, new_n20151_, new_n20152_, new_n20153_,
    new_n20163_, new_n20164_, new_n20165_, new_n20166_, new_n20167_,
    new_n20168_, new_n20169_, new_n20170_, new_n20171_, new_n20172_,
    new_n20173_, new_n20174_, new_n20175_, new_n20176_, new_n20177_,
    new_n20178_, new_n20179_, new_n20180_, new_n20181_, new_n20182_,
    new_n20183_, new_n20184_, new_n20185_, new_n20186_, new_n20187_,
    new_n20188_, new_n20189_, new_n20190_, new_n20191_, new_n20192_,
    new_n20193_, new_n20194_, new_n20195_, new_n20196_, new_n20197_,
    new_n20198_, new_n20199_, new_n20200_, new_n20201_, new_n20202_,
    new_n20203_, new_n20204_, new_n20205_, new_n20206_, new_n20207_,
    new_n20208_, new_n20209_, new_n20210_, new_n20211_, new_n20212_,
    new_n20213_, new_n20214_, new_n20215_, new_n20216_, new_n20217_,
    new_n20218_, new_n20219_, new_n20220_, new_n20221_, new_n20222_,
    new_n20223_, new_n20224_, new_n20225_, new_n20227_, new_n20228_,
    new_n20229_, new_n20230_, new_n20231_, new_n20232_, new_n20233_,
    new_n20234_, new_n20235_, new_n20236_, new_n20237_, new_n20238_,
    new_n20239_, new_n20240_, new_n20241_, new_n20242_, new_n20243_,
    new_n20244_, new_n20245_, new_n20246_, new_n20247_, new_n20248_,
    new_n20249_, new_n20250_, new_n20251_, new_n20252_, new_n20253_,
    new_n20254_, new_n20255_, new_n20256_, new_n20257_, new_n20258_,
    new_n20259_, new_n20260_, new_n20261_, new_n20262_, new_n20263_,
    new_n20265_, new_n20266_, new_n20267_, new_n20268_, new_n20269_,
    new_n20270_, new_n20271_, new_n20272_, new_n20273_, new_n20274_,
    new_n20275_, new_n20276_, new_n20277_, new_n20278_, new_n20279_,
    new_n20280_, new_n20281_, new_n20282_, new_n20283_, new_n20284_,
    new_n20285_, new_n20286_, new_n20287_, new_n20288_, new_n20289_,
    new_n20290_, new_n20291_, new_n20292_, new_n20293_, new_n20294_,
    new_n20295_, new_n20296_, new_n20297_, new_n20298_, new_n20299_,
    new_n20300_, new_n20301_, new_n20302_, new_n20303_, new_n20304_,
    new_n20305_, new_n20306_, new_n20307_, new_n20308_, new_n20309_,
    new_n20310_, new_n20311_, new_n20312_, new_n20313_, new_n20314_,
    new_n20315_, new_n20316_, new_n20317_, new_n20318_, new_n20319_,
    new_n20320_, new_n20321_, new_n20322_, new_n20323_, new_n20324_,
    new_n20325_, new_n20326_, new_n20327_, new_n20328_, new_n20329_,
    new_n20330_, new_n20331_, new_n20332_, new_n20333_, new_n20334_,
    new_n20335_, new_n20336_, new_n20337_, new_n20338_, new_n20339_,
    new_n20340_, new_n20341_, new_n20342_, new_n20343_, new_n20344_,
    new_n20345_, new_n20346_, new_n20347_, new_n20348_, new_n20349_,
    new_n20350_, new_n20351_, new_n20352_, new_n20353_, new_n20354_,
    new_n20355_, new_n20356_, new_n20357_, new_n20358_, new_n20359_,
    new_n20360_, new_n20361_, new_n20362_, new_n20363_, new_n20364_,
    new_n20365_, new_n20366_, new_n20367_, new_n20368_, new_n20369_,
    new_n20370_, new_n20371_, new_n20372_, new_n20373_, new_n20374_,
    new_n20375_, new_n20376_, new_n20377_, new_n20378_, new_n20379_,
    new_n20380_, new_n20381_, new_n20382_, new_n20383_, new_n20384_,
    new_n20385_, new_n20386_, new_n20387_, new_n20388_, new_n20389_,
    new_n20390_, new_n20391_, new_n20392_, new_n20393_, new_n20394_,
    new_n20395_, new_n20396_, new_n20397_, new_n20398_, new_n20399_,
    new_n20400_, new_n20401_, new_n20402_, new_n20403_, new_n20404_,
    new_n20405_, new_n20406_, new_n20407_, new_n20408_, new_n20409_,
    new_n20410_, new_n20411_, new_n20412_, new_n20413_, new_n20414_,
    new_n20415_, new_n20416_, new_n20417_, new_n20418_, new_n20419_,
    new_n20421_, new_n20422_, new_n20423_, new_n20424_, new_n20425_,
    new_n20426_, new_n20427_, new_n20428_, new_n20429_, new_n20430_,
    new_n20431_, new_n20432_, new_n20433_, new_n20434_, new_n20435_,
    new_n20436_, new_n20437_, new_n20438_, new_n20439_, new_n20440_,
    new_n20441_, new_n20442_, new_n20443_, new_n20444_, new_n20445_,
    new_n20446_, new_n20447_, new_n20448_, new_n20449_, new_n20450_,
    new_n20451_, new_n20452_, new_n20453_, new_n20454_, new_n20455_,
    new_n20456_, new_n20457_, new_n20458_, new_n20459_, new_n20460_,
    new_n20461_, new_n20462_, new_n20463_, new_n20464_, new_n20465_,
    new_n20466_, new_n20467_, new_n20468_, new_n20469_, new_n20470_,
    new_n20471_, new_n20472_, new_n20473_, new_n20474_, new_n20475_,
    new_n20476_, new_n20477_, new_n20478_, new_n20479_, new_n20480_,
    new_n20481_, new_n20482_, new_n20483_, new_n20484_, new_n20485_,
    new_n20486_, new_n20487_, new_n20488_, new_n20489_, new_n20490_,
    new_n20491_, new_n20492_, new_n20493_, new_n20494_, new_n20495_,
    new_n20496_, new_n20497_, new_n20498_, new_n20499_, new_n20500_,
    new_n20501_, new_n20502_, new_n20503_, new_n20504_, new_n20505_,
    new_n20506_, new_n20507_, new_n20508_, new_n20509_, new_n20510_,
    new_n20511_, new_n20512_, new_n20513_, new_n20514_, new_n20515_,
    new_n20516_, new_n20517_, new_n20518_, new_n20519_, new_n20520_,
    new_n20521_, new_n20522_, new_n20523_, new_n20524_, new_n20525_,
    new_n20526_, new_n20527_, new_n20528_, new_n20529_, new_n20530_,
    new_n20531_, new_n20532_, new_n20533_, new_n20534_, new_n20535_,
    new_n20536_, new_n20537_, new_n20538_, new_n20539_, new_n20540_,
    new_n20541_, new_n20542_, new_n20543_, new_n20544_, new_n20545_,
    new_n20546_, new_n20547_, new_n20548_, new_n20549_, new_n20550_,
    new_n20551_, new_n20552_, new_n20553_, new_n20554_, new_n20555_,
    new_n20556_, new_n20557_, new_n20558_, new_n20559_, new_n20560_,
    new_n20561_, new_n20562_, new_n20563_, new_n20564_, new_n20565_,
    new_n20566_, new_n20567_, new_n20568_, new_n20569_, new_n20570_,
    new_n20571_, new_n20572_, new_n20573_, new_n20574_, new_n20575_,
    new_n20576_, new_n20577_, new_n20578_, new_n20579_, new_n20580_,
    new_n20581_, new_n20582_, new_n20583_, new_n20584_, new_n20585_,
    new_n20586_, new_n20587_, new_n20588_, new_n20589_, new_n20591_,
    new_n20592_, new_n20593_, new_n20594_, new_n20595_, new_n20596_,
    new_n20597_, new_n20598_, new_n20599_, new_n20600_, new_n20601_,
    new_n20602_, new_n20603_, new_n20604_, new_n20605_, new_n20606_,
    new_n20607_, new_n20608_, new_n20609_, new_n20610_, new_n20611_,
    new_n20612_, new_n20613_, new_n20614_, new_n20615_, new_n20616_,
    new_n20617_, new_n20618_, new_n20619_, new_n20620_, new_n20621_,
    new_n20622_, new_n20623_, new_n20624_, new_n20625_, new_n20626_,
    new_n20627_, new_n20629_, new_n20630_, new_n20631_, new_n20632_,
    new_n20633_, new_n20634_, new_n20635_, new_n20636_, new_n20637_,
    new_n20638_, new_n20639_, new_n20640_, new_n20641_, new_n20642_,
    new_n20643_, new_n20644_, new_n20645_, new_n20646_, new_n20647_,
    new_n20648_, new_n20649_, new_n20650_, new_n20651_, new_n20652_,
    new_n20653_, new_n20654_, new_n20655_, new_n20656_, new_n20657_,
    new_n20658_, new_n20659_, new_n20660_, new_n20661_, new_n20662_,
    new_n20663_, new_n20664_, new_n20665_, new_n20666_, new_n20667_,
    new_n20668_, new_n20669_, new_n20670_, new_n20671_, new_n20672_,
    new_n20673_, new_n20674_, new_n20675_, new_n20676_, new_n20677_,
    new_n20678_, new_n20679_, new_n20680_, new_n20681_, new_n20682_,
    new_n20683_, new_n20684_, new_n20685_, new_n20686_, new_n20687_,
    new_n20688_, new_n20689_, new_n20690_, new_n20691_, new_n20692_,
    new_n20693_, new_n20694_, new_n20695_, new_n20696_, new_n20697_,
    new_n20698_, new_n20699_, new_n20700_, new_n20701_, new_n20702_,
    new_n20703_, new_n20704_, new_n20705_, new_n20706_, new_n20707_,
    new_n20708_, new_n20709_, new_n20710_, new_n20711_, new_n20712_,
    new_n20713_, new_n20714_, new_n20715_, new_n20716_, new_n20717_,
    new_n20718_, new_n20719_, new_n20720_, new_n20721_, new_n20722_,
    new_n20723_, new_n20724_, new_n20725_, new_n20726_, new_n20727_,
    new_n20728_, new_n20729_, new_n20730_, new_n20731_, new_n20732_,
    new_n20733_, new_n20734_, new_n20735_, new_n20736_, new_n20738_,
    new_n20739_, new_n20740_, new_n20741_, new_n20742_, new_n20743_,
    new_n20744_, new_n20745_, new_n20746_, new_n20747_, new_n20748_,
    new_n20749_, new_n20750_, new_n20751_, new_n20752_, new_n20753_,
    new_n20754_, new_n20755_, new_n20756_, new_n20757_, new_n20758_,
    new_n20759_, new_n20760_, new_n20761_, new_n20762_, new_n20763_,
    new_n20764_, new_n20765_, new_n20766_, new_n20767_, new_n20768_,
    new_n20769_, new_n20770_, new_n20771_, new_n20772_, new_n20773_,
    new_n20774_, new_n20775_, new_n20776_, new_n20777_, new_n20778_,
    new_n20779_, new_n20780_, new_n20781_, new_n20782_, new_n20783_,
    new_n20784_, new_n20785_, new_n20786_, new_n20787_, new_n20788_,
    new_n20789_, new_n20790_, new_n20791_, new_n20792_, new_n20793_,
    new_n20794_, new_n20795_, new_n20796_, new_n20797_, new_n20798_,
    new_n20799_, new_n20800_, new_n20801_, new_n20802_, new_n20803_,
    new_n20804_, new_n20805_, new_n20806_, new_n20807_, new_n20808_,
    new_n20809_, new_n20810_, new_n20811_, new_n20812_, new_n20813_,
    new_n20814_, new_n20815_, new_n20816_, new_n20817_, new_n20818_,
    new_n20819_, new_n20820_, new_n20821_, new_n20822_, new_n20823_,
    new_n20824_, new_n20825_, new_n20826_, new_n20827_, new_n20828_,
    new_n20829_, new_n20830_, new_n20831_, new_n20832_, new_n20833_,
    new_n20834_, new_n20835_, new_n20836_, new_n20837_, new_n20838_,
    new_n20839_, new_n20840_, new_n20841_, new_n20842_, new_n20843_,
    new_n20844_, new_n20845_, new_n20846_, new_n20847_, new_n20848_,
    new_n20849_, new_n20850_, new_n20851_, new_n20852_, new_n20853_,
    new_n20854_, new_n20855_, new_n20856_, new_n20857_, new_n20858_,
    new_n20859_, new_n20860_, new_n20861_, new_n20862_, new_n20863_,
    new_n20864_, new_n20865_, new_n20866_, new_n20867_, new_n20868_,
    new_n20869_, new_n20870_, new_n20871_, new_n20872_, new_n20873_,
    new_n20874_, new_n20875_, new_n20876_, new_n20877_, new_n20878_,
    new_n20879_, new_n20880_, new_n20881_, new_n20882_, new_n20883_,
    new_n20884_, new_n20885_, new_n20886_, new_n20887_, new_n20888_,
    new_n20889_, new_n20890_, new_n20891_, new_n20892_, new_n20893_,
    new_n20894_, new_n20895_, new_n20896_, new_n20897_, new_n20898_,
    new_n20899_, new_n20900_, new_n20901_, new_n20902_, new_n20903_,
    new_n20904_, new_n20905_, new_n20906_, new_n20907_, new_n20908_,
    new_n20909_, new_n20910_, new_n20911_, new_n20912_, new_n20913_,
    new_n20914_, new_n20915_, new_n20916_, new_n20917_, new_n20918_,
    new_n20919_, new_n20920_, new_n20921_, new_n20922_, new_n20923_,
    new_n20924_, new_n20925_, new_n20927_, new_n20928_, new_n20929_,
    new_n20930_, new_n20931_, new_n20932_, new_n20933_, new_n20934_,
    new_n20935_, new_n20936_, new_n20937_, new_n20938_, new_n20939_,
    new_n20940_, new_n20941_, new_n20942_, new_n20943_, new_n20944_,
    new_n20945_, new_n20946_, new_n20947_, new_n20948_, new_n20949_,
    new_n20950_, new_n20951_, new_n20952_, new_n20953_, new_n20954_,
    new_n20955_, new_n20956_, new_n20957_, new_n20958_, new_n20959_,
    new_n20960_, new_n20961_, new_n20962_, new_n20963_, new_n20965_,
    new_n20966_, new_n20967_, new_n20968_, new_n20969_, new_n20970_,
    new_n20971_, new_n20972_, new_n20973_, new_n20974_, new_n20975_,
    new_n20976_, new_n20977_, new_n20978_, new_n20979_, new_n20980_,
    new_n20981_, new_n20982_, new_n20983_, new_n20984_, new_n20985_,
    new_n20986_, new_n20987_, new_n20988_, new_n20989_, new_n20990_,
    new_n20991_, new_n20992_, new_n20993_, new_n20994_, new_n20995_,
    new_n20996_, new_n20997_, new_n20998_, new_n20999_, new_n21000_,
    new_n21001_, new_n21002_, new_n21003_, new_n21004_, new_n21005_,
    new_n21006_, new_n21007_, new_n21008_, new_n21009_, new_n21010_,
    new_n21011_, new_n21012_, new_n21013_, new_n21014_, new_n21015_,
    new_n21016_, new_n21017_, new_n21018_, new_n21019_, new_n21020_,
    new_n21021_, new_n21022_, new_n21023_, new_n21024_, new_n21025_,
    new_n21026_, new_n21027_, new_n21028_, new_n21029_, new_n21030_,
    new_n21031_, new_n21032_, new_n21033_, new_n21034_, new_n21035_,
    new_n21036_, new_n21037_, new_n21038_, new_n21039_, new_n21040_,
    new_n21041_, new_n21042_, new_n21043_, new_n21044_, new_n21045_,
    new_n21046_, new_n21047_, new_n21048_, new_n21049_, new_n21050_,
    new_n21051_, new_n21052_, new_n21053_, new_n21054_, new_n21055_,
    new_n21056_, new_n21057_, new_n21058_, new_n21059_, new_n21060_,
    new_n21061_, new_n21062_, new_n21063_, new_n21064_, new_n21065_,
    new_n21066_, new_n21067_, new_n21068_, new_n21069_, new_n21070_,
    new_n21071_, new_n21072_, new_n21073_, new_n21075_, new_n21076_,
    new_n21077_, new_n21078_, new_n21079_, new_n21080_, new_n21081_,
    new_n21082_, new_n21083_, new_n21084_, new_n21085_, new_n21086_,
    new_n21087_, new_n21088_, new_n21089_, new_n21090_, new_n21091_,
    new_n21092_, new_n21093_, new_n21094_, new_n21095_, new_n21096_,
    new_n21097_, new_n21098_, new_n21099_, new_n21100_, new_n21101_,
    new_n21102_, new_n21103_, new_n21104_, new_n21105_, new_n21106_,
    new_n21107_, new_n21108_, new_n21109_, new_n21110_, new_n21111_,
    new_n21112_, new_n21113_, new_n21114_, new_n21115_, new_n21116_,
    new_n21117_, new_n21118_, new_n21119_, new_n21120_, new_n21121_,
    new_n21122_, new_n21123_, new_n21124_, new_n21125_, new_n21126_,
    new_n21127_, new_n21128_, new_n21129_, new_n21130_, new_n21131_,
    new_n21132_, new_n21133_, new_n21134_, new_n21135_, new_n21136_,
    new_n21137_, new_n21138_, new_n21139_, new_n21140_, new_n21141_,
    new_n21142_, new_n21143_, new_n21144_, new_n21145_, new_n21146_,
    new_n21147_, new_n21148_, new_n21149_, new_n21150_, new_n21151_,
    new_n21152_, new_n21153_, new_n21154_, new_n21155_, new_n21156_,
    new_n21157_, new_n21158_, new_n21159_, new_n21160_, new_n21161_,
    new_n21162_, new_n21163_, new_n21164_, new_n21165_, new_n21166_,
    new_n21167_, new_n21168_, new_n21169_, new_n21170_, new_n21171_,
    new_n21172_, new_n21173_, new_n21174_, new_n21175_, new_n21176_,
    new_n21177_, new_n21178_, new_n21179_, new_n21180_, new_n21181_,
    new_n21182_, new_n21183_, new_n21184_, new_n21185_, new_n21186_,
    new_n21187_, new_n21188_, new_n21189_, new_n21190_, new_n21191_,
    new_n21192_, new_n21193_, new_n21194_, new_n21195_, new_n21196_,
    new_n21197_, new_n21198_, new_n21199_, new_n21200_, new_n21201_,
    new_n21202_, new_n21203_, new_n21204_, new_n21205_, new_n21206_,
    new_n21207_, new_n21208_, new_n21209_, new_n21210_, new_n21211_,
    new_n21212_, new_n21213_, new_n21214_, new_n21215_, new_n21216_,
    new_n21217_, new_n21218_, new_n21219_, new_n21220_, new_n21221_,
    new_n21222_, new_n21223_, new_n21224_, new_n21225_, new_n21226_,
    new_n21227_, new_n21228_, new_n21229_, new_n21230_, new_n21231_,
    new_n21232_, new_n21233_, new_n21234_, new_n21235_, new_n21236_,
    new_n21237_, new_n21238_, new_n21239_, new_n21240_, new_n21241_,
    new_n21242_, new_n21243_, new_n21244_, new_n21245_, new_n21246_,
    new_n21247_, new_n21248_, new_n21249_, new_n21250_, new_n21251_,
    new_n21252_, new_n21253_, new_n21254_, new_n21255_, new_n21256_,
    new_n21257_, new_n21258_, new_n21259_, new_n21260_, new_n21261_,
    new_n21262_, new_n21263_, new_n21264_, new_n21265_, new_n21266_,
    new_n21267_, new_n21268_, new_n21269_, new_n21271_, new_n21272_,
    new_n21273_, new_n21274_, new_n21275_, new_n21276_, new_n21277_,
    new_n21278_, new_n21279_, new_n21280_, new_n21281_, new_n21282_,
    new_n21283_, new_n21284_, new_n21285_, new_n21286_, new_n21287_,
    new_n21288_, new_n21289_, new_n21290_, new_n21291_, new_n21292_,
    new_n21293_, new_n21294_, new_n21295_, new_n21296_, new_n21297_,
    new_n21298_, new_n21299_, new_n21300_, new_n21301_, new_n21302_,
    new_n21303_, new_n21304_, new_n21305_, new_n21306_, new_n21307_,
    new_n21308_, new_n21309_, new_n21310_, new_n21311_, new_n21312_,
    new_n21313_, new_n21314_, new_n21315_, new_n21316_, new_n21317_,
    new_n21318_, new_n21319_, new_n21320_, new_n21321_, new_n21322_,
    new_n21323_, new_n21324_, new_n21325_, new_n21326_, new_n21327_,
    new_n21328_, new_n21329_, new_n21330_, new_n21331_, new_n21332_,
    new_n21333_, new_n21334_, new_n21335_, new_n21336_, new_n21337_,
    new_n21338_, new_n21339_, new_n21340_, new_n21341_, new_n21342_,
    new_n21343_, new_n21344_, new_n21345_, new_n21346_, new_n21347_,
    new_n21348_, new_n21349_, new_n21350_, new_n21351_, new_n21352_,
    new_n21353_, new_n21354_, new_n21355_, new_n21356_, new_n21357_,
    new_n21358_, new_n21359_, new_n21360_, new_n21361_, new_n21362_,
    new_n21363_, new_n21364_, new_n21365_, new_n21366_, new_n21367_,
    new_n21368_, new_n21369_, new_n21370_, new_n21371_, new_n21372_,
    new_n21373_, new_n21374_, new_n21375_, new_n21376_, new_n21377_,
    new_n21378_, new_n21379_, new_n21380_, new_n21381_, new_n21382_,
    new_n21383_, new_n21384_, new_n21385_, new_n21386_, new_n21387_,
    new_n21388_, new_n21389_, new_n21390_, new_n21391_, new_n21392_,
    new_n21393_, new_n21394_, new_n21395_, new_n21396_, new_n21397_,
    new_n21398_, new_n21399_, new_n21400_, new_n21401_, new_n21402_,
    new_n21403_, new_n21404_, new_n21405_, new_n21406_, new_n21407_,
    new_n21410_, new_n21411_, new_n21412_, new_n21413_, new_n21414_,
    new_n21415_, new_n21416_, new_n21417_, new_n21418_, new_n21419_,
    new_n21420_, new_n21421_, new_n21422_, new_n21423_, new_n21424_,
    new_n21425_, new_n21426_, new_n21427_, new_n21428_, new_n21429_,
    new_n21430_, new_n21431_, new_n21432_, new_n21433_, new_n21434_,
    new_n21435_, new_n21436_, new_n21437_, new_n21438_, new_n21439_,
    new_n21440_, new_n21441_, new_n21442_, new_n21443_, new_n21444_,
    new_n21445_, new_n21446_, new_n21447_, new_n21448_, new_n21449_,
    new_n21450_, new_n21451_, new_n21452_, new_n21453_, new_n21454_,
    new_n21455_, new_n21456_, new_n21457_, new_n21458_, new_n21459_,
    new_n21460_, new_n21461_, new_n21462_, new_n21463_, new_n21464_,
    new_n21465_, new_n21466_, new_n21467_, new_n21468_, new_n21469_,
    new_n21470_, new_n21471_, new_n21472_, new_n21473_, new_n21474_,
    new_n21475_, new_n21476_, new_n21477_, new_n21478_, new_n21479_,
    new_n21480_, new_n21481_, new_n21482_, new_n21483_, new_n21484_,
    new_n21485_, new_n21486_, new_n21487_, new_n21488_, new_n21489_,
    new_n21490_, new_n21491_, new_n21492_, new_n21493_, new_n21494_,
    new_n21495_, new_n21496_, new_n21497_, new_n21498_, new_n21499_,
    new_n21500_, new_n21501_, new_n21502_, new_n21503_, new_n21504_,
    new_n21505_, new_n21506_, new_n21507_, new_n21508_, new_n21509_,
    new_n21510_, new_n21511_, new_n21512_, new_n21513_, new_n21514_,
    new_n21515_, new_n21516_, new_n21517_, new_n21518_, new_n21519_,
    new_n21520_, new_n21521_, new_n21522_, new_n21523_, new_n21524_,
    new_n21525_, new_n21526_, new_n21527_, new_n21528_, new_n21529_,
    new_n21530_, new_n21531_, new_n21532_, new_n21533_, new_n21534_,
    new_n21535_, new_n21536_, new_n21537_, new_n21538_, new_n21539_,
    new_n21540_, new_n21541_, new_n21542_, new_n21543_, new_n21544_,
    new_n21545_, new_n21546_, new_n21547_, new_n21548_, new_n21549_,
    new_n21550_, new_n21551_, new_n21552_, new_n21553_, new_n21554_,
    new_n21555_, new_n21556_, new_n21557_, new_n21558_, new_n21559_,
    new_n21560_, new_n21561_, new_n21562_, new_n21563_, new_n21564_,
    new_n21565_, new_n21566_, new_n21567_, new_n21568_, new_n21569_,
    new_n21570_, new_n21571_, new_n21572_, new_n21573_, new_n21574_,
    new_n21575_, new_n21576_, new_n21577_, new_n21578_, new_n21579_,
    new_n21580_, new_n21581_, new_n21582_, new_n21583_, new_n21584_,
    new_n21585_, new_n21586_, new_n21587_, new_n21588_, new_n21589_,
    new_n21590_, new_n21591_, new_n21592_, new_n21593_, new_n21595_,
    new_n21596_, new_n21597_, new_n21598_, new_n21599_, new_n21600_,
    new_n21601_, new_n21602_, new_n21603_, new_n21604_, new_n21605_,
    new_n21606_, new_n21607_, new_n21608_, new_n21609_, new_n21610_,
    new_n21611_, new_n21612_, new_n21613_, new_n21614_, new_n21615_,
    new_n21616_, new_n21617_, new_n21618_, new_n21619_, new_n21620_,
    new_n21621_, new_n21622_, new_n21623_, new_n21624_, new_n21625_,
    new_n21626_, new_n21627_, new_n21628_, new_n21629_, new_n21631_,
    new_n21632_, new_n21633_, new_n21634_, new_n21635_, new_n21636_,
    new_n21637_, new_n21638_, new_n21639_, new_n21640_, new_n21641_,
    new_n21642_, new_n21643_, new_n21644_, new_n21645_, new_n21646_,
    new_n21647_, new_n21648_, new_n21649_, new_n21650_, new_n21651_,
    new_n21652_, new_n21653_, new_n21654_, new_n21655_, new_n21656_,
    new_n21657_, new_n21658_, new_n21659_, new_n21660_, new_n21661_,
    new_n21662_, new_n21663_, new_n21664_, new_n21665_, new_n21666_,
    new_n21667_, new_n21668_, new_n21669_, new_n21670_, new_n21671_,
    new_n21672_, new_n21673_, new_n21674_, new_n21675_, new_n21676_,
    new_n21677_, new_n21678_, new_n21679_, new_n21680_, new_n21681_,
    new_n21682_, new_n21683_, new_n21684_, new_n21685_, new_n21686_,
    new_n21687_, new_n21688_, new_n21689_, new_n21690_, new_n21691_,
    new_n21692_, new_n21693_, new_n21694_, new_n21695_, new_n21696_,
    new_n21697_, new_n21698_, new_n21699_, new_n21700_, new_n21701_,
    new_n21702_, new_n21703_, new_n21704_, new_n21705_, new_n21706_,
    new_n21707_, new_n21708_, new_n21709_, new_n21710_, new_n21711_,
    new_n21712_, new_n21713_, new_n21714_, new_n21715_, new_n21716_,
    new_n21717_, new_n21718_, new_n21719_, new_n21720_, new_n21721_,
    new_n21722_, new_n21723_, new_n21724_, new_n21725_, new_n21726_,
    new_n21727_, new_n21728_, new_n21729_, new_n21730_, new_n21731_,
    new_n21732_, new_n21733_, new_n21734_, new_n21735_, new_n21736_,
    new_n21737_, new_n21738_, new_n21739_, new_n21740_, new_n21741_,
    new_n21742_, new_n21743_, new_n21744_, new_n21745_, new_n21746_,
    new_n21747_, new_n21748_, new_n21749_, new_n21750_, new_n21751_,
    new_n21752_, new_n21753_, new_n21754_, new_n21755_, new_n21756_,
    new_n21757_, new_n21758_, new_n21759_, new_n21760_, new_n21761_,
    new_n21762_, new_n21763_, new_n21764_, new_n21765_, new_n21766_,
    new_n21767_, new_n21768_, new_n21769_, new_n21770_, new_n21771_,
    new_n21772_, new_n21773_, new_n21774_, new_n21775_, new_n21776_,
    new_n21777_, new_n21778_, new_n21779_, new_n21780_, new_n21781_,
    new_n21782_, new_n21783_, new_n21784_, new_n21785_, new_n21786_,
    new_n21787_, new_n21788_, new_n21789_, new_n21790_, new_n21791_,
    new_n21792_, new_n21793_, new_n21794_, new_n21795_, new_n21796_,
    new_n21797_, new_n21798_, new_n21799_, new_n21800_, new_n21801_,
    new_n21802_, new_n21803_, new_n21804_, new_n21805_, new_n21806_,
    new_n21807_, new_n21808_, new_n21809_, new_n21810_, new_n21811_,
    new_n21812_, new_n21813_, new_n21814_, new_n21815_, new_n21816_,
    new_n21817_, new_n21818_, new_n21819_, new_n21820_, new_n21821_,
    new_n21822_, new_n21823_, new_n21824_, new_n21825_, new_n21826_,
    new_n21827_, new_n21828_, new_n21829_, new_n21830_, new_n21831_,
    new_n21832_, new_n21833_, new_n21834_, new_n21835_, new_n21836_,
    new_n21837_, new_n21838_, new_n21839_, new_n21840_, new_n21841_,
    new_n21842_, new_n21843_, new_n21844_, new_n21845_, new_n21846_,
    new_n21847_, new_n21848_, new_n21849_, new_n21850_, new_n21851_,
    new_n21852_, new_n21853_, new_n21854_, new_n21855_, new_n21856_,
    new_n21857_, new_n21858_, new_n21859_, new_n21860_, new_n21861_,
    new_n21862_, new_n21863_, new_n21864_, new_n21865_, new_n21866_,
    new_n21867_, new_n21868_, new_n21869_, new_n21870_, new_n21871_,
    new_n21872_, new_n21873_, new_n21874_, new_n21875_, new_n21876_,
    new_n21877_, new_n21878_, new_n21879_, new_n21881_, new_n21882_,
    new_n21883_, new_n21884_, new_n21885_, new_n21886_, new_n21887_,
    new_n21888_, new_n21889_, new_n21890_, new_n21891_, new_n21892_,
    new_n21893_, new_n21894_, new_n21895_, new_n21896_, new_n21897_,
    new_n21898_, new_n21899_, new_n21900_, new_n21901_, new_n21902_,
    new_n21903_, new_n21904_, new_n21905_, new_n21906_, new_n21907_,
    new_n21908_, new_n21909_, new_n21910_, new_n21911_, new_n21912_,
    new_n21913_, new_n21914_, new_n21915_, new_n21917_, new_n21918_,
    new_n21919_, new_n21920_, new_n21921_, new_n21922_, new_n21923_,
    new_n21924_, new_n21925_, new_n21926_, new_n21927_, new_n21928_,
    new_n21929_, new_n21930_, new_n21931_, new_n21932_, new_n21933_,
    new_n21934_, new_n21935_, new_n21936_, new_n21937_, new_n21938_,
    new_n21939_, new_n21940_, new_n21941_, new_n21942_, new_n21943_,
    new_n21944_, new_n21945_, new_n21946_, new_n21947_, new_n21948_,
    new_n21949_, new_n21950_, new_n21951_, new_n21952_, new_n21953_,
    new_n21954_, new_n21955_, new_n21956_, new_n21957_, new_n21958_,
    new_n21959_, new_n21960_, new_n21961_, new_n21962_, new_n21963_,
    new_n21964_, new_n21965_, new_n21966_, new_n21967_, new_n21968_,
    new_n21969_, new_n21970_, new_n21971_, new_n21972_, new_n21973_,
    new_n21974_, new_n21975_, new_n21976_, new_n21977_, new_n21978_,
    new_n21979_, new_n21980_, new_n21981_, new_n21982_, new_n21983_,
    new_n21984_, new_n21985_, new_n21986_, new_n21987_, new_n21988_,
    new_n21989_, new_n21990_, new_n21991_, new_n21992_, new_n21993_,
    new_n21994_, new_n21995_, new_n21996_, new_n21997_, new_n21998_,
    new_n21999_, new_n22000_, new_n22001_, new_n22002_, new_n22003_,
    new_n22004_, new_n22005_, new_n22006_, new_n22007_, new_n22008_,
    new_n22009_, new_n22010_, new_n22011_, new_n22012_, new_n22013_,
    new_n22014_, new_n22015_, new_n22016_, new_n22017_, new_n22018_,
    new_n22019_, new_n22020_, new_n22021_, new_n22022_, new_n22023_,
    new_n22024_, new_n22025_, new_n22026_, new_n22027_, new_n22028_,
    new_n22029_, new_n22030_, new_n22031_, new_n22032_, new_n22033_,
    new_n22034_, new_n22035_, new_n22036_, new_n22037_, new_n22038_,
    new_n22039_, new_n22040_, new_n22041_, new_n22042_, new_n22043_,
    new_n22044_, new_n22045_, new_n22046_, new_n22047_, new_n22048_,
    new_n22049_, new_n22050_, new_n22051_, new_n22052_, new_n22053_,
    new_n22054_, new_n22055_, new_n22056_, new_n22057_, new_n22058_,
    new_n22059_, new_n22060_, new_n22061_, new_n22062_, new_n22063_,
    new_n22064_, new_n22065_, new_n22066_, new_n22067_, new_n22068_,
    new_n22069_, new_n22070_, new_n22071_, new_n22072_, new_n22073_,
    new_n22074_, new_n22075_, new_n22076_, new_n22077_, new_n22078_,
    new_n22079_, new_n22080_, new_n22081_, new_n22082_, new_n22083_,
    new_n22084_, new_n22085_, new_n22086_, new_n22087_, new_n22088_,
    new_n22089_, new_n22090_, new_n22091_, new_n22092_, new_n22093_,
    new_n22094_, new_n22095_, new_n22096_, new_n22097_, new_n22098_,
    new_n22099_, new_n22100_, new_n22101_, new_n22102_, new_n22103_,
    new_n22104_, new_n22105_, new_n22106_, new_n22107_, new_n22108_,
    new_n22109_, new_n22110_, new_n22111_, new_n22112_, new_n22113_,
    new_n22114_, new_n22115_, new_n22116_, new_n22117_, new_n22118_,
    new_n22119_, new_n22120_, new_n22121_, new_n22122_, new_n22123_,
    new_n22124_, new_n22125_, new_n22126_, new_n22127_, new_n22128_,
    new_n22129_, new_n22130_, new_n22131_, new_n22132_, new_n22133_,
    new_n22134_, new_n22135_, new_n22136_, new_n22137_, new_n22138_,
    new_n22139_, new_n22140_, new_n22141_, new_n22142_, new_n22143_,
    new_n22144_, new_n22145_, new_n22146_, new_n22147_, new_n22148_,
    new_n22149_, new_n22150_, new_n22151_, new_n22152_, new_n22153_,
    new_n22154_, new_n22155_, new_n22156_, new_n22157_, new_n22158_,
    new_n22159_, new_n22160_, new_n22161_, new_n22162_, new_n22163_,
    new_n22164_, new_n22165_, new_n22167_, new_n22168_, new_n22169_,
    new_n22170_, new_n22171_, new_n22172_, new_n22173_, new_n22174_,
    new_n22175_, new_n22176_, new_n22177_, new_n22178_, new_n22179_,
    new_n22180_, new_n22181_, new_n22182_, new_n22183_, new_n22184_,
    new_n22185_, new_n22186_, new_n22187_, new_n22188_, new_n22189_,
    new_n22190_, new_n22191_, new_n22192_, new_n22193_, new_n22194_,
    new_n22195_, new_n22196_, new_n22197_, new_n22198_, new_n22199_,
    new_n22200_, new_n22201_, new_n22203_, new_n22204_, new_n22205_,
    new_n22206_, new_n22207_, new_n22208_, new_n22209_, new_n22210_,
    new_n22211_, new_n22212_, new_n22213_, new_n22214_, new_n22215_,
    new_n22216_, new_n22217_, new_n22218_, new_n22219_, new_n22220_,
    new_n22221_, new_n22222_, new_n22223_, new_n22224_, new_n22225_,
    new_n22226_, new_n22227_, new_n22228_, new_n22229_, new_n22230_,
    new_n22231_, new_n22232_, new_n22233_, new_n22234_, new_n22235_,
    new_n22236_, new_n22237_, new_n22238_, new_n22239_, new_n22240_,
    new_n22241_, new_n22242_, new_n22243_, new_n22244_, new_n22245_,
    new_n22246_, new_n22247_, new_n22248_, new_n22249_, new_n22250_,
    new_n22251_, new_n22252_, new_n22253_, new_n22254_, new_n22255_,
    new_n22256_, new_n22257_, new_n22258_, new_n22259_, new_n22260_,
    new_n22261_, new_n22262_, new_n22263_, new_n22264_, new_n22265_,
    new_n22266_, new_n22267_, new_n22268_, new_n22269_, new_n22270_,
    new_n22271_, new_n22272_, new_n22273_, new_n22274_, new_n22275_,
    new_n22276_, new_n22277_, new_n22278_, new_n22279_, new_n22280_,
    new_n22281_, new_n22282_, new_n22283_, new_n22284_, new_n22285_,
    new_n22286_, new_n22287_, new_n22288_, new_n22289_, new_n22290_,
    new_n22291_, new_n22292_, new_n22293_, new_n22294_, new_n22295_,
    new_n22296_, new_n22297_, new_n22298_, new_n22299_, new_n22300_,
    new_n22301_, new_n22302_, new_n22303_, new_n22304_, new_n22305_,
    new_n22306_, new_n22307_, new_n22308_, new_n22309_, new_n22310_,
    new_n22311_, new_n22312_, new_n22313_, new_n22314_, new_n22315_,
    new_n22316_, new_n22317_, new_n22318_, new_n22319_, new_n22320_,
    new_n22321_, new_n22322_, new_n22323_, new_n22324_, new_n22325_,
    new_n22326_, new_n22327_, new_n22328_, new_n22329_, new_n22330_,
    new_n22331_, new_n22332_, new_n22333_, new_n22334_, new_n22335_,
    new_n22336_, new_n22337_, new_n22338_, new_n22339_, new_n22340_,
    new_n22341_, new_n22342_, new_n22343_, new_n22344_, new_n22345_,
    new_n22346_, new_n22347_, new_n22348_, new_n22349_, new_n22350_,
    new_n22351_, new_n22352_, new_n22353_, new_n22354_, new_n22355_,
    new_n22356_, new_n22357_, new_n22358_, new_n22359_, new_n22360_,
    new_n22361_, new_n22362_, new_n22363_, new_n22364_, new_n22365_,
    new_n22366_, new_n22367_, new_n22368_, new_n22369_, new_n22370_,
    new_n22371_, new_n22372_, new_n22373_, new_n22374_, new_n22375_,
    new_n22376_, new_n22377_, new_n22378_, new_n22379_, new_n22380_,
    new_n22381_, new_n22382_, new_n22383_, new_n22384_, new_n22385_,
    new_n22386_, new_n22387_, new_n22388_, new_n22389_, new_n22390_,
    new_n22391_, new_n22392_, new_n22393_, new_n22394_, new_n22395_,
    new_n22396_, new_n22397_, new_n22398_, new_n22399_, new_n22400_,
    new_n22401_, new_n22402_, new_n22403_, new_n22404_, new_n22405_,
    new_n22406_, new_n22407_, new_n22408_, new_n22409_, new_n22410_,
    new_n22411_, new_n22412_, new_n22413_, new_n22414_, new_n22415_,
    new_n22416_, new_n22417_, new_n22418_, new_n22419_, new_n22420_,
    new_n22421_, new_n22422_, new_n22423_, new_n22424_, new_n22425_,
    new_n22426_, new_n22427_, new_n22428_, new_n22429_, new_n22430_,
    new_n22431_, new_n22432_, new_n22433_, new_n22434_, new_n22435_,
    new_n22436_, new_n22437_, new_n22438_, new_n22439_, new_n22440_,
    new_n22441_, new_n22442_, new_n22443_, new_n22444_, new_n22445_,
    new_n22446_, new_n22447_, new_n22448_, new_n22449_, new_n22450_,
    new_n22451_, new_n22453_, new_n22454_, new_n22455_, new_n22456_,
    new_n22457_, new_n22458_, new_n22459_, new_n22460_, new_n22461_,
    new_n22462_, new_n22463_, new_n22464_, new_n22465_, new_n22466_,
    new_n22467_, new_n22468_, new_n22469_, new_n22470_, new_n22471_,
    new_n22472_, new_n22473_, new_n22474_, new_n22475_, new_n22476_,
    new_n22477_, new_n22478_, new_n22479_, new_n22480_, new_n22481_,
    new_n22482_, new_n22483_, new_n22484_, new_n22485_, new_n22486_,
    new_n22487_, new_n22489_, new_n22490_, new_n22491_, new_n22492_,
    new_n22493_, new_n22494_, new_n22495_, new_n22496_, new_n22497_,
    new_n22498_, new_n22499_, new_n22500_, new_n22501_, new_n22502_,
    new_n22503_, new_n22504_, new_n22505_, new_n22506_, new_n22507_,
    new_n22508_, new_n22509_, new_n22510_, new_n22511_, new_n22512_,
    new_n22513_, new_n22514_, new_n22515_, new_n22516_, new_n22517_,
    new_n22518_, new_n22519_, new_n22520_, new_n22521_, new_n22522_,
    new_n22523_, new_n22524_, new_n22525_, new_n22526_, new_n22527_,
    new_n22528_, new_n22529_, new_n22530_, new_n22531_, new_n22532_,
    new_n22533_, new_n22534_, new_n22535_, new_n22536_, new_n22537_,
    new_n22538_, new_n22539_, new_n22540_, new_n22541_, new_n22542_,
    new_n22543_, new_n22544_, new_n22545_, new_n22546_, new_n22547_,
    new_n22548_, new_n22549_, new_n22550_, new_n22551_, new_n22552_,
    new_n22553_, new_n22554_, new_n22555_, new_n22556_, new_n22557_,
    new_n22558_, new_n22559_, new_n22560_, new_n22561_, new_n22562_,
    new_n22563_, new_n22564_, new_n22565_, new_n22566_, new_n22567_,
    new_n22568_, new_n22569_, new_n22570_, new_n22571_, new_n22572_,
    new_n22573_, new_n22574_, new_n22575_, new_n22576_, new_n22577_,
    new_n22578_, new_n22579_, new_n22580_, new_n22581_, new_n22582_,
    new_n22583_, new_n22584_, new_n22585_, new_n22586_, new_n22587_,
    new_n22588_, new_n22589_, new_n22590_, new_n22591_, new_n22592_,
    new_n22593_, new_n22594_, new_n22595_, new_n22596_, new_n22597_,
    new_n22598_, new_n22599_, new_n22600_, new_n22601_, new_n22602_,
    new_n22603_, new_n22604_, new_n22605_, new_n22606_, new_n22607_,
    new_n22608_, new_n22609_, new_n22610_, new_n22611_, new_n22612_,
    new_n22613_, new_n22614_, new_n22615_, new_n22616_, new_n22617_,
    new_n22618_, new_n22619_, new_n22620_, new_n22621_, new_n22622_,
    new_n22623_, new_n22624_, new_n22625_, new_n22626_, new_n22627_,
    new_n22628_, new_n22629_, new_n22630_, new_n22631_, new_n22632_,
    new_n22633_, new_n22634_, new_n22635_, new_n22636_, new_n22637_,
    new_n22638_, new_n22639_, new_n22640_, new_n22641_, new_n22642_,
    new_n22643_, new_n22644_, new_n22645_, new_n22646_, new_n22647_,
    new_n22648_, new_n22649_, new_n22650_, new_n22651_, new_n22652_,
    new_n22653_, new_n22654_, new_n22655_, new_n22656_, new_n22657_,
    new_n22658_, new_n22659_, new_n22660_, new_n22661_, new_n22662_,
    new_n22663_, new_n22664_, new_n22665_, new_n22666_, new_n22667_,
    new_n22668_, new_n22669_, new_n22670_, new_n22671_, new_n22672_,
    new_n22673_, new_n22674_, new_n22675_, new_n22676_, new_n22677_,
    new_n22678_, new_n22679_, new_n22680_, new_n22681_, new_n22682_,
    new_n22683_, new_n22684_, new_n22685_, new_n22686_, new_n22687_,
    new_n22688_, new_n22689_, new_n22690_, new_n22691_, new_n22692_,
    new_n22693_, new_n22694_, new_n22695_, new_n22696_, new_n22697_,
    new_n22698_, new_n22699_, new_n22700_, new_n22701_, new_n22702_,
    new_n22703_, new_n22704_, new_n22705_, new_n22706_, new_n22707_,
    new_n22708_, new_n22709_, new_n22710_, new_n22711_, new_n22712_,
    new_n22713_, new_n22714_, new_n22715_, new_n22716_, new_n22717_,
    new_n22718_, new_n22719_, new_n22720_, new_n22721_, new_n22722_,
    new_n22723_, new_n22724_, new_n22725_, new_n22726_, new_n22727_,
    new_n22728_, new_n22729_, new_n22731_, new_n22732_, new_n22733_,
    new_n22734_, new_n22735_, new_n22736_, new_n22737_, new_n22738_,
    new_n22739_, new_n22740_, new_n22741_, new_n22742_, new_n22743_,
    new_n22744_, new_n22745_, new_n22746_, new_n22747_, new_n22748_,
    new_n22749_, new_n22750_, new_n22751_, new_n22752_, new_n22753_,
    new_n22754_, new_n22755_, new_n22756_, new_n22757_, new_n22758_,
    new_n22759_, new_n22760_, new_n22761_, new_n22762_, new_n22763_,
    new_n22764_, new_n22765_, new_n22766_, new_n22767_, new_n22769_,
    new_n22770_, new_n22771_, new_n22772_, new_n22773_, new_n22774_,
    new_n22775_, new_n22776_, new_n22777_, new_n22778_, new_n22779_,
    new_n22780_, new_n22781_, new_n22782_, new_n22783_, new_n22784_,
    new_n22785_, new_n22786_, new_n22787_, new_n22788_, new_n22789_,
    new_n22790_, new_n22791_, new_n22792_, new_n22793_, new_n22794_,
    new_n22795_, new_n22796_, new_n22797_, new_n22798_, new_n22799_,
    new_n22800_, new_n22801_, new_n22802_, new_n22803_, new_n22804_,
    new_n22805_, new_n22806_, new_n22807_, new_n22808_, new_n22809_,
    new_n22810_, new_n22811_, new_n22812_, new_n22813_, new_n22814_,
    new_n22815_, new_n22816_, new_n22817_, new_n22818_, new_n22819_,
    new_n22820_, new_n22821_, new_n22822_, new_n22823_, new_n22824_,
    new_n22825_, new_n22826_, new_n22827_, new_n22828_, new_n22829_,
    new_n22830_, new_n22831_, new_n22832_, new_n22833_, new_n22834_,
    new_n22835_, new_n22836_, new_n22837_, new_n22838_, new_n22839_,
    new_n22840_, new_n22841_, new_n22842_, new_n22843_, new_n22844_,
    new_n22845_, new_n22846_, new_n22847_, new_n22848_, new_n22849_,
    new_n22850_, new_n22851_, new_n22852_, new_n22853_, new_n22854_,
    new_n22855_, new_n22856_, new_n22857_, new_n22858_, new_n22859_,
    new_n22860_, new_n22861_, new_n22862_, new_n22863_, new_n22864_,
    new_n22865_, new_n22866_, new_n22867_, new_n22868_, new_n22869_,
    new_n22870_, new_n22871_, new_n22872_, new_n22873_, new_n22874_,
    new_n22875_, new_n22876_, new_n22877_, new_n22878_, new_n22879_,
    new_n22880_, new_n22881_, new_n22882_, new_n22883_, new_n22884_,
    new_n22885_, new_n22886_, new_n22887_, new_n22888_, new_n22889_,
    new_n22890_, new_n22891_, new_n22892_, new_n22893_, new_n22894_,
    new_n22895_, new_n22896_, new_n22897_, new_n22898_, new_n22899_,
    new_n22900_, new_n22901_, new_n22902_, new_n22903_, new_n22904_,
    new_n22905_, new_n22906_, new_n22907_, new_n22908_, new_n22909_,
    new_n22910_, new_n22911_, new_n22912_, new_n22913_, new_n22914_,
    new_n22915_, new_n22916_, new_n22917_, new_n22918_, new_n22919_,
    new_n22920_, new_n22921_, new_n22922_, new_n22923_, new_n22924_,
    new_n22925_, new_n22926_, new_n22927_, new_n22928_, new_n22929_,
    new_n22930_, new_n22931_, new_n22932_, new_n22933_, new_n22934_,
    new_n22935_, new_n22936_, new_n22937_, new_n22938_, new_n22939_,
    new_n22940_, new_n22941_, new_n22942_, new_n22943_, new_n22944_,
    new_n22945_, new_n22946_, new_n22947_, new_n22948_, new_n22949_,
    new_n22950_, new_n22951_, new_n22952_, new_n22953_, new_n22954_,
    new_n22955_, new_n22956_, new_n22957_, new_n22958_, new_n22959_,
    new_n22960_, new_n22961_, new_n22962_, new_n22963_, new_n22964_,
    new_n22965_, new_n22966_, new_n22967_, new_n22968_, new_n22969_,
    new_n22970_, new_n22971_, new_n22972_, new_n22973_, new_n22974_,
    new_n22975_, new_n22976_, new_n22977_, new_n22978_, new_n22979_,
    new_n22980_, new_n22981_, new_n22982_, new_n22983_, new_n22984_,
    new_n22985_, new_n22986_, new_n22987_, new_n22988_, new_n22989_,
    new_n22990_, new_n22991_, new_n22992_, new_n22993_, new_n22994_,
    new_n22995_, new_n22996_, new_n22997_, new_n22998_, new_n22999_,
    new_n23000_, new_n23001_, new_n23002_, new_n23003_, new_n23004_,
    new_n23005_, new_n23006_, new_n23007_, new_n23008_, new_n23009_,
    new_n23010_, new_n23011_, new_n23012_, new_n23013_, new_n23014_,
    new_n23015_, new_n23016_, new_n23017_, new_n23018_, new_n23019_,
    new_n23020_, new_n23021_, new_n23022_, new_n23023_, new_n23024_,
    new_n23025_, new_n23026_, new_n23027_, new_n23028_, new_n23029_,
    new_n23030_, new_n23031_, new_n23032_, new_n23033_, new_n23034_,
    new_n23035_, new_n23036_, new_n23037_, new_n23038_, new_n23039_,
    new_n23040_, new_n23041_, new_n23042_, new_n23043_, new_n23044_,
    new_n23045_, new_n23046_, new_n23047_, new_n23048_, new_n23049_,
    new_n23050_, new_n23051_, new_n23052_, new_n23053_, new_n23054_,
    new_n23055_, new_n23056_, new_n23057_, new_n23058_, new_n23059_,
    new_n23060_, new_n23061_, new_n23062_, new_n23063_, new_n23064_,
    new_n23065_, new_n23066_, new_n23068_, new_n23070_, new_n23071_,
    new_n23072_, new_n23073_, new_n23074_, new_n23075_, new_n23076_,
    new_n23077_, new_n23078_, new_n23079_, new_n23080_, new_n23081_,
    new_n23082_, new_n23083_, new_n23084_, new_n23085_, new_n23086_,
    new_n23087_, new_n23088_, new_n23089_, new_n23090_, new_n23091_,
    new_n23092_, new_n23093_, new_n23094_, new_n23095_, new_n23096_,
    new_n23098_, new_n23099_, new_n23100_, new_n23101_, new_n23102_,
    new_n23103_, new_n23104_, new_n23105_, new_n23106_, new_n23107_,
    new_n23108_, new_n23109_, new_n23110_, new_n23111_, new_n23112_,
    new_n23113_, new_n23114_, new_n23115_, new_n23116_, new_n23117_,
    new_n23118_, new_n23119_, new_n23120_, new_n23121_, new_n23122_,
    new_n23123_, new_n23124_, new_n23125_, new_n23126_, new_n23127_,
    new_n23128_, new_n23129_, new_n23130_, new_n23131_, new_n23132_,
    new_n23133_, new_n23134_, new_n23135_, new_n23136_, new_n23137_,
    new_n23138_, new_n23140_, new_n23141_, new_n23142_, new_n23143_,
    new_n23144_, new_n23145_, new_n23146_, new_n23147_, new_n23148_,
    new_n23149_, new_n23150_, new_n23151_, new_n23152_, new_n23153_,
    new_n23154_, new_n23155_, new_n23156_, new_n23157_, new_n23158_,
    new_n23159_, new_n23161_, new_n23162_, new_n23163_, new_n23164_,
    new_n23165_, new_n23166_, new_n23167_, new_n23169_, new_n23170_,
    new_n23171_, new_n23172_, new_n23173_, new_n23174_, new_n23175_,
    new_n23176_, new_n23177_, new_n23178_, new_n23179_, new_n23180_,
    new_n23181_, new_n23182_, new_n23183_, new_n23184_, new_n23185_,
    new_n23186_, new_n23187_, new_n23188_, new_n23189_, new_n23190_,
    new_n23191_, new_n23192_, new_n23193_, new_n23194_, new_n23195_,
    new_n23196_, new_n23197_, new_n23198_, new_n23199_, new_n23200_,
    new_n23201_, new_n23202_, new_n23203_, new_n23204_, new_n23205_,
    new_n23206_, new_n23207_, new_n23208_, new_n23209_, new_n23210_,
    new_n23211_, new_n23212_, new_n23213_, new_n23214_, new_n23215_,
    new_n23216_, new_n23217_, new_n23218_, new_n23219_, new_n23220_,
    new_n23221_, new_n23222_, new_n23223_, new_n23224_, new_n23225_,
    new_n23226_, new_n23227_, new_n23228_, new_n23229_, new_n23230_,
    new_n23231_, new_n23232_, new_n23233_, new_n23234_, new_n23235_,
    new_n23236_, new_n23237_, new_n23238_, new_n23239_, new_n23240_,
    new_n23241_, new_n23242_, new_n23243_, new_n23244_, new_n23245_,
    new_n23246_, new_n23247_, new_n23248_, new_n23249_, new_n23250_,
    new_n23251_, new_n23252_, new_n23253_, new_n23254_, new_n23255_,
    new_n23256_, new_n23257_, new_n23258_, new_n23259_, new_n23260_,
    new_n23261_, new_n23262_, new_n23263_, new_n23264_, new_n23265_,
    new_n23266_, new_n23267_, new_n23268_, new_n23269_, new_n23270_,
    new_n23271_, new_n23272_, new_n23273_, new_n23274_, new_n23275_,
    new_n23276_, new_n23277_, new_n23278_, new_n23279_, new_n23280_,
    new_n23281_, new_n23282_, new_n23283_, new_n23284_, new_n23285_,
    new_n23286_, new_n23287_, new_n23288_, new_n23289_, new_n23290_,
    new_n23291_, new_n23292_, new_n23293_, new_n23294_, new_n23295_,
    new_n23296_, new_n23297_, new_n23298_, new_n23299_, new_n23300_,
    new_n23301_, new_n23302_, new_n23303_, new_n23304_, new_n23305_,
    new_n23306_, new_n23307_, new_n23308_, new_n23309_, new_n23310_,
    new_n23311_, new_n23312_, new_n23313_, new_n23314_, new_n23315_,
    new_n23316_, new_n23317_, new_n23318_, new_n23319_, new_n23320_,
    new_n23321_, new_n23322_, new_n23323_, new_n23324_, new_n23325_,
    new_n23326_, new_n23327_, new_n23328_, new_n23329_, new_n23330_,
    new_n23331_, new_n23332_, new_n23333_, new_n23334_, new_n23335_,
    new_n23336_, new_n23337_, new_n23338_, new_n23339_, new_n23340_,
    new_n23341_, new_n23342_, new_n23343_, new_n23344_, new_n23345_,
    new_n23346_, new_n23347_, new_n23348_, new_n23349_, new_n23350_,
    new_n23351_, new_n23352_, new_n23353_, new_n23354_, new_n23355_,
    new_n23356_, new_n23357_, new_n23358_, new_n23359_, new_n23360_,
    new_n23361_, new_n23362_, new_n23363_, new_n23364_, new_n23365_,
    new_n23366_, new_n23367_, new_n23368_, new_n23369_, new_n23370_,
    new_n23371_, new_n23372_, new_n23373_, new_n23374_, new_n23375_,
    new_n23376_, new_n23377_, new_n23378_, new_n23379_, new_n23380_,
    new_n23381_, new_n23382_, new_n23383_, new_n23384_, new_n23385_,
    new_n23386_, new_n23387_, new_n23388_, new_n23389_, new_n23390_,
    new_n23391_, new_n23392_, new_n23393_, new_n23394_, new_n23395_,
    new_n23396_, new_n23397_, new_n23398_, new_n23399_, new_n23400_,
    new_n23401_, new_n23402_, new_n23403_, new_n23404_, new_n23405_,
    new_n23406_, new_n23407_, new_n23408_, new_n23409_, new_n23410_,
    new_n23411_, new_n23412_, new_n23413_, new_n23414_, new_n23415_,
    new_n23416_, new_n23417_, new_n23418_, new_n23419_, new_n23420_,
    new_n23421_, new_n23422_, new_n23423_, new_n23424_, new_n23425_,
    new_n23426_, new_n23429_, new_n23430_, new_n23431_, new_n23438_,
    new_n23439_, new_n23440_, new_n23441_, new_n23442_, new_n23443_,
    new_n23444_, new_n23445_, new_n23446_, new_n23447_, new_n23448_,
    new_n23449_, new_n23450_, new_n23451_, new_n23452_, new_n23453_,
    new_n23454_, new_n23455_, new_n23456_, new_n23457_, new_n23458_,
    new_n23459_, new_n23460_, new_n23461_, new_n23462_, new_n23463_,
    new_n23464_, new_n23465_, new_n23466_, new_n23467_, new_n23468_,
    new_n23469_, new_n23470_, new_n23471_, new_n23472_, new_n23473_,
    new_n23474_, new_n23475_, new_n23476_, new_n23477_, new_n23478_,
    new_n23479_, new_n23480_, new_n23481_, new_n23482_, new_n23483_,
    new_n23484_, new_n23485_, new_n23486_, new_n23487_, new_n23488_,
    new_n23489_, new_n23490_, new_n23491_, new_n23492_, new_n23493_,
    new_n23494_, new_n23495_, new_n23496_, new_n23497_, new_n23498_,
    new_n23499_, new_n23500_, new_n23501_, new_n23502_, new_n23503_,
    new_n23507_, new_n23508_, new_n23509_, new_n23510_, new_n23511_,
    new_n23512_, new_n23513_, new_n23514_, new_n23515_, new_n23516_,
    new_n23517_, new_n23518_, new_n23519_, new_n23520_, new_n23521_,
    new_n23522_, new_n23523_, new_n23524_, new_n23525_, new_n23526_,
    new_n23527_, new_n23528_, new_n23529_, new_n23530_, new_n23531_,
    new_n23532_, new_n23533_, new_n23534_, new_n23535_, new_n23536_,
    new_n23537_, new_n23538_, new_n23539_, new_n23540_, new_n23541_,
    new_n23542_, new_n23543_, new_n23544_, new_n23545_, new_n23546_,
    new_n23547_, new_n23548_, new_n23549_, new_n23550_, new_n23551_,
    new_n23552_, new_n23553_, new_n23554_, new_n23555_, new_n23556_,
    new_n23557_, new_n23558_, new_n23559_, new_n23560_, new_n23561_,
    new_n23562_, new_n23563_, new_n23564_, new_n23565_, new_n23566_,
    new_n23567_, new_n23568_, new_n23569_, new_n23570_, new_n23571_,
    new_n23572_, new_n23573_, new_n23574_, new_n23575_, new_n23576_,
    new_n23577_, new_n23578_, new_n23579_, new_n23580_, new_n23581_,
    new_n23584_, new_n23585_, new_n23586_, new_n23587_, new_n23588_,
    new_n23589_, new_n23590_, new_n23591_, new_n23592_, new_n23593_,
    new_n23594_, new_n23595_, new_n23597_, new_n23598_, new_n23599_,
    new_n23600_, new_n23601_, new_n23602_, new_n23603_, new_n23604_,
    new_n23605_, new_n23606_, new_n23607_, new_n23608_, new_n23609_,
    new_n23610_, new_n23611_, new_n23612_, new_n23613_, new_n23614_,
    new_n23615_, new_n23616_, new_n23617_, new_n23618_, new_n23619_,
    new_n23620_, new_n23621_, new_n23622_, new_n23623_, new_n23624_,
    new_n23625_, new_n23626_, new_n23627_, new_n23628_, new_n23629_,
    new_n23630_, new_n23631_, new_n23632_, new_n23633_, new_n23634_,
    new_n23635_, new_n23636_, new_n23637_, new_n23638_, new_n23639_,
    new_n23640_, new_n23641_, new_n23642_, new_n23643_, new_n23644_,
    new_n23645_, new_n23646_, new_n23647_, new_n23648_, new_n23649_,
    new_n23650_, new_n23651_, new_n23652_, new_n23653_, new_n23654_,
    new_n23655_, new_n23656_, new_n23657_, new_n23658_, new_n23659_,
    new_n23660_, new_n23661_, new_n23662_, new_n23663_, new_n23664_,
    new_n23665_, new_n23666_, new_n23667_, new_n23668_, new_n23669_,
    new_n23670_, new_n23671_, new_n23672_, new_n23673_, new_n23674_,
    new_n23675_, new_n23676_, new_n23677_, new_n23678_, new_n23679_,
    new_n23680_, new_n23681_, new_n23682_, new_n23683_, new_n23684_,
    new_n23685_, new_n23686_, new_n23687_, new_n23688_, new_n23689_,
    new_n23690_, new_n23691_, new_n23692_, new_n23693_, new_n23694_,
    new_n23695_, new_n23696_, new_n23697_, new_n23698_, new_n23699_,
    new_n23700_, new_n23701_, new_n23704_, new_n23705_, new_n23706_,
    new_n23707_, new_n23708_, new_n23709_, new_n23710_, new_n23711_,
    new_n23712_, new_n23713_, new_n23714_, new_n23715_, new_n23716_,
    new_n23717_, new_n23718_, new_n23719_, new_n23720_, new_n23721_,
    new_n23722_, new_n23723_, new_n23724_, new_n23725_, new_n23726_,
    new_n23727_, new_n23728_, new_n23729_, new_n23730_, new_n23731_,
    new_n23732_, new_n23733_, new_n23734_, new_n23735_, new_n23736_,
    new_n23737_, new_n23738_, new_n23739_, new_n23740_, new_n23741_,
    new_n23742_, new_n23743_, new_n23744_, new_n23745_, new_n23746_,
    new_n23747_, new_n23748_, new_n23749_, new_n23750_, new_n23751_,
    new_n23752_, new_n23753_, new_n23754_, new_n23755_, new_n23756_,
    new_n23757_, new_n23758_, new_n23759_, new_n23760_, new_n23761_,
    new_n23762_, new_n23763_, new_n23764_, new_n23765_, new_n23766_,
    new_n23767_, new_n23768_, new_n23769_, new_n23770_, new_n23771_,
    new_n23772_, new_n23773_, new_n23774_, new_n23775_, new_n23776_,
    new_n23777_, new_n23778_, new_n23779_, new_n23780_, new_n23781_,
    new_n23782_, new_n23783_, new_n23784_, new_n23785_, new_n23786_,
    new_n23787_, new_n23788_, new_n23789_, new_n23790_, new_n23791_,
    new_n23792_, new_n23793_, new_n23794_, new_n23795_, new_n23796_,
    new_n23797_, new_n23798_, new_n23799_, new_n23800_, new_n23801_,
    new_n23802_, new_n23803_, new_n23804_, new_n23805_, new_n23806_,
    new_n23807_, new_n23808_, new_n23809_, new_n23810_, new_n23811_,
    new_n23812_, new_n23813_, new_n23814_, new_n23815_, new_n23816_,
    new_n23817_, new_n23818_, new_n23819_, new_n23820_, new_n23821_,
    new_n23822_, new_n23823_, new_n23824_, new_n23825_, new_n23826_,
    new_n23827_, new_n23828_, new_n23829_, new_n23830_, new_n23831_,
    new_n23832_, new_n23833_, new_n23834_, new_n23835_, new_n23836_,
    new_n23837_, new_n23838_, new_n23839_, new_n23840_, new_n23841_,
    new_n23842_, new_n23843_, new_n23844_, new_n23845_, new_n23846_,
    new_n23847_, new_n23848_, new_n23849_, new_n23850_, new_n23851_,
    new_n23852_, new_n23853_, new_n23854_, new_n23855_, new_n23856_,
    new_n23857_, new_n23858_, new_n23859_, new_n23860_, new_n23861_,
    new_n23862_, new_n23863_, new_n23864_, new_n23865_, new_n23866_,
    new_n23867_, new_n23868_, new_n23869_, new_n23871_, new_n23872_,
    new_n23873_, new_n23874_, new_n23875_, new_n23876_, new_n23877_,
    new_n23878_, new_n23879_, new_n23880_, new_n23881_, new_n23882_,
    new_n23884_, new_n23885_, new_n23886_, new_n23887_, new_n23888_,
    new_n23889_, new_n23890_, new_n23891_, new_n23892_, new_n23893_,
    new_n23894_, new_n23895_, new_n23896_, new_n23897_, new_n23898_,
    new_n23899_, new_n23900_, new_n23901_, new_n23902_, new_n23903_,
    new_n23904_, new_n23905_, new_n23906_, new_n23907_, new_n23908_,
    new_n23909_, new_n23910_, new_n23911_, new_n23912_, new_n23913_,
    new_n23914_, new_n23915_, new_n23916_, new_n23917_, new_n23918_,
    new_n23919_, new_n23920_, new_n23921_, new_n23922_, new_n23923_,
    new_n23924_, new_n23925_, new_n23926_, new_n23927_, new_n23928_,
    new_n23929_, new_n23930_, new_n23931_, new_n23932_, new_n23933_,
    new_n23934_, new_n23935_, new_n23936_, new_n23937_, new_n23938_,
    new_n23939_, new_n23940_, new_n23941_, new_n23942_, new_n23943_,
    new_n23944_, new_n23945_, new_n23946_, new_n23947_, new_n23948_,
    new_n23949_, new_n23950_, new_n23951_, new_n23952_, new_n23953_,
    new_n23954_, new_n23955_, new_n23956_, new_n23957_, new_n23958_,
    new_n23959_, new_n23960_, new_n23961_, new_n23962_, new_n23963_,
    new_n23964_, new_n23965_, new_n23966_, new_n23967_, new_n23968_,
    new_n23969_, new_n23970_, new_n23971_, new_n23972_, new_n23973_,
    new_n23974_, new_n23975_, new_n23976_, new_n23977_, new_n23978_,
    new_n23979_, new_n23980_, new_n23981_, new_n23982_, new_n23983_,
    new_n23984_, new_n23985_, new_n23986_, new_n23987_, new_n23988_,
    new_n23989_, new_n23990_, new_n23991_, new_n23992_, new_n23993_,
    new_n23994_, new_n23995_, new_n23996_, new_n23997_, new_n23998_,
    new_n23999_, new_n24000_, new_n24001_, new_n24002_, new_n24003_,
    new_n24004_, new_n24005_, new_n24006_, new_n24007_, new_n24008_,
    new_n24009_, new_n24010_, new_n24011_, new_n24012_, new_n24013_,
    new_n24014_, new_n24015_, new_n24016_, new_n24017_, new_n24018_,
    new_n24019_, new_n24020_, new_n24021_, new_n24022_, new_n24023_,
    new_n24024_, new_n24025_, new_n24026_, new_n24027_, new_n24028_,
    new_n24029_, new_n24030_, new_n24031_, new_n24032_, new_n24033_,
    new_n24034_, new_n24035_, new_n24036_, new_n24037_, new_n24038_,
    new_n24039_, new_n24040_, new_n24041_, new_n24042_, new_n24043_,
    new_n24044_, new_n24045_, new_n24046_, new_n24048_, new_n24049_,
    new_n24058_, new_n24059_, new_n24060_, new_n24061_, new_n24062_,
    new_n24063_, new_n24064_, new_n24065_, new_n24066_, new_n24067_,
    new_n24068_, new_n24069_, new_n24070_, new_n24071_, new_n24072_,
    new_n24073_, new_n24074_, new_n24075_, new_n24076_, new_n24077_,
    new_n24078_, new_n24080_, new_n24081_, new_n24082_, new_n24083_,
    new_n24084_, new_n24086_, new_n24087_, new_n24088_, new_n24089_,
    new_n24090_, new_n24092_, new_n24093_, new_n24094_, new_n24095_,
    new_n24096_, new_n24097_, new_n24098_, new_n24099_, new_n24100_,
    new_n24101_, new_n24102_, new_n24103_, new_n24104_, new_n24105_,
    new_n24106_, new_n24107_, new_n24108_, new_n24109_, new_n24110_,
    new_n24111_, new_n24112_, new_n24113_, new_n24114_, new_n24115_,
    new_n24116_, new_n24118_, new_n24119_, new_n24120_, new_n24122_,
    new_n24123_, new_n24124_, new_n24125_, new_n24126_, new_n24128_,
    new_n24129_, new_n24130_, new_n24131_, new_n24132_, new_n24133_,
    new_n24134_, new_n24135_, new_n24136_, new_n24137_, new_n24138_,
    new_n24139_, new_n24140_, new_n24141_, new_n24142_, new_n24143_,
    new_n24144_, new_n24145_, new_n24146_, new_n24147_, new_n24148_,
    new_n24149_, new_n24150_, new_n24151_, new_n24152_, new_n24153_,
    new_n24154_, new_n24155_, new_n24156_, new_n24157_, new_n24158_,
    new_n24159_, new_n24160_, new_n24161_, new_n24162_, new_n24163_,
    new_n24164_, new_n24165_, new_n24166_, new_n24167_, new_n24168_,
    new_n24169_, new_n24170_, new_n24171_, new_n24172_, new_n24173_,
    new_n24174_, new_n24175_, new_n24176_, new_n24177_, new_n24178_,
    new_n24179_, new_n24180_, new_n24181_, new_n24182_, new_n24183_,
    new_n24184_, new_n24185_, new_n24186_, new_n24187_, new_n24188_,
    new_n24189_, new_n24190_, new_n24191_, new_n24192_, new_n24193_,
    new_n24194_, new_n24195_, new_n24196_, new_n24197_, new_n24198_,
    new_n24199_, new_n24200_, new_n24201_, new_n24202_, new_n24203_,
    new_n24204_, new_n24205_, new_n24206_, new_n24207_, new_n24208_,
    new_n24209_, new_n24210_, new_n24211_, new_n24212_, new_n24213_,
    new_n24214_, new_n24215_, new_n24216_, new_n24217_, new_n24218_,
    new_n24219_, new_n24220_, new_n24221_, new_n24222_, new_n24223_,
    new_n24224_, new_n24225_, new_n24226_, new_n24227_, new_n24228_,
    new_n24229_, new_n24230_, new_n24231_, new_n24232_, new_n24233_,
    new_n24234_, new_n24235_, new_n24236_, new_n24237_, new_n24238_,
    new_n24239_, new_n24240_, new_n24241_, new_n24242_, new_n24243_,
    new_n24244_, new_n24245_, new_n24246_, new_n24247_, new_n24248_,
    new_n24249_, new_n24250_, new_n24251_, new_n24252_, new_n24253_,
    new_n24254_, new_n24255_, new_n24256_, new_n24257_, new_n24258_,
    new_n24259_, new_n24260_, new_n24261_, new_n24262_, new_n24263_,
    new_n24264_, new_n24265_, new_n24266_, new_n24267_, new_n24268_,
    new_n24269_, new_n24270_, new_n24271_, new_n24272_, new_n24273_,
    new_n24274_, new_n24275_, new_n24276_, new_n24277_, new_n24278_,
    new_n24279_, new_n24280_, new_n24281_, new_n24282_, new_n24283_,
    new_n24284_, new_n24285_, new_n24286_, new_n24287_, new_n24288_,
    new_n24289_, new_n24290_, new_n24291_, new_n24292_, new_n24293_,
    new_n24294_, new_n24295_, new_n24296_, new_n24297_, new_n24298_,
    new_n24299_, new_n24300_, new_n24301_, new_n24302_, new_n24303_,
    new_n24304_, new_n24305_, new_n24306_, new_n24307_, new_n24308_,
    new_n24309_, new_n24310_, new_n24311_, new_n24312_, new_n24313_,
    new_n24314_, new_n24315_, new_n24316_, new_n24317_, new_n24318_,
    new_n24319_, new_n24320_, new_n24321_, new_n24322_, new_n24323_,
    new_n24324_, new_n24325_, new_n24326_, new_n24327_, new_n24328_,
    new_n24329_, new_n24330_, new_n24331_, new_n24332_, new_n24333_,
    new_n24334_, new_n24335_, new_n24336_, new_n24337_, new_n24338_,
    new_n24339_, new_n24340_, new_n24341_, new_n24342_, new_n24343_,
    new_n24344_, new_n24345_, new_n24346_, new_n24347_, new_n24348_,
    new_n24349_, new_n24350_, new_n24351_, new_n24352_, new_n24353_,
    new_n24354_, new_n24355_, new_n24356_, new_n24357_, new_n24358_,
    new_n24359_, new_n24360_, new_n24361_, new_n24362_, new_n24363_,
    new_n24364_, new_n24365_, new_n24366_, new_n24367_, new_n24368_,
    new_n24369_, new_n24370_, new_n24371_, new_n24372_, new_n24373_,
    new_n24374_, new_n24375_, new_n24376_, new_n24377_, new_n24378_,
    new_n24379_, new_n24380_, new_n24381_, new_n24382_, new_n24383_,
    new_n24384_, new_n24385_, new_n24386_, new_n24387_, new_n24388_,
    new_n24389_, new_n24390_, new_n24391_, new_n24392_, new_n24393_,
    new_n24394_, new_n24395_, new_n24396_, new_n24397_, new_n24398_,
    new_n24399_, new_n24400_, new_n24401_, new_n24402_, new_n24403_,
    new_n24404_, new_n24405_, new_n24406_, new_n24407_, new_n24408_,
    new_n24409_, new_n24410_, new_n24411_, new_n24412_, new_n24413_,
    new_n24414_, new_n24415_, new_n24416_, new_n24417_, new_n24418_,
    new_n24419_, new_n24420_, new_n24421_, new_n24422_, new_n24423_,
    new_n24424_, new_n24425_, new_n24426_, new_n24427_, new_n24428_,
    new_n24429_, new_n24430_, new_n24431_, new_n24432_, new_n24433_,
    new_n24434_, new_n24435_, new_n24436_, new_n24437_, new_n24438_,
    new_n24439_, new_n24440_, new_n24441_, new_n24442_, new_n24443_,
    new_n24444_, new_n24445_, new_n24446_, new_n24447_, new_n24448_,
    new_n24449_, new_n24450_, new_n24451_, new_n24452_, new_n24453_,
    new_n24454_, new_n24455_, new_n24456_, new_n24457_, new_n24458_,
    new_n24459_, new_n24460_, new_n24461_, new_n24462_, new_n24463_,
    new_n24464_, new_n24465_, new_n24466_, new_n24467_, new_n24468_,
    new_n24469_, new_n24470_, new_n24471_, new_n24472_, new_n24473_,
    new_n24474_, new_n24475_, new_n24476_, new_n24477_, new_n24478_,
    new_n24479_, new_n24480_, new_n24481_, new_n24482_, new_n24483_,
    new_n24484_, new_n24485_, new_n24486_, new_n24487_, new_n24488_,
    new_n24489_, new_n24490_, new_n24491_, new_n24493_, new_n24494_,
    new_n24495_, new_n24496_, new_n24497_, new_n24498_, new_n24499_,
    new_n24500_, new_n24501_, new_n24502_, new_n24503_, new_n24504_,
    new_n24505_, new_n24506_, new_n24507_, new_n24508_, new_n24509_,
    new_n24510_, new_n24511_, new_n24512_, new_n24513_, new_n24514_,
    new_n24515_, new_n24516_, new_n24517_, new_n24518_, new_n24519_,
    new_n24520_, new_n24521_, new_n24522_, new_n24523_, new_n24524_,
    new_n24525_, new_n24526_, new_n24527_, new_n24528_, new_n24529_,
    new_n24530_, new_n24531_, new_n24532_, new_n24533_, new_n24534_,
    new_n24535_, new_n24536_, new_n24538_, new_n24539_, new_n24540_,
    new_n24541_, new_n24542_, new_n24543_, new_n24544_, new_n24545_,
    new_n24546_, new_n24547_, new_n24548_, new_n24549_, new_n24550_,
    new_n24551_, new_n24552_, new_n24553_, new_n24554_, new_n24555_,
    new_n24556_, new_n24557_, new_n24558_, new_n24559_, new_n24560_,
    new_n24561_, new_n24562_, new_n24563_, new_n24564_, new_n24565_,
    new_n24566_, new_n24567_, new_n24568_, new_n24569_, new_n24570_,
    new_n24571_, new_n24573_, new_n24574_, new_n24575_, new_n24576_,
    new_n24577_, new_n24578_, new_n24579_, new_n24580_, new_n24581_,
    new_n24582_, new_n24583_, new_n24584_, new_n24585_, new_n24586_,
    new_n24587_, new_n24588_, new_n24589_, new_n24590_, new_n24591_,
    new_n24592_, new_n24593_, new_n24594_, new_n24595_, new_n24596_,
    new_n24597_, new_n24598_, new_n24599_, new_n24600_, new_n24601_,
    new_n24602_, new_n24603_, new_n24604_, new_n24605_, new_n24606_,
    new_n24607_, new_n24608_, new_n24609_, new_n24610_, new_n24611_,
    new_n24612_, new_n24613_, new_n24614_, new_n24615_, new_n24616_,
    new_n24617_, new_n24618_, new_n24619_, new_n24620_, new_n24621_,
    new_n24622_, new_n24623_, new_n24624_, new_n24625_, new_n24626_,
    new_n24627_, new_n24628_, new_n24629_, new_n24630_, new_n24631_,
    new_n24632_, new_n24633_, new_n24634_, new_n24635_, new_n24636_,
    new_n24637_, new_n24638_, new_n24639_, new_n24640_, new_n24641_,
    new_n24642_, new_n24643_, new_n24644_, new_n24645_, new_n24647_,
    new_n24648_, new_n24649_, new_n24650_, new_n24651_, new_n24652_,
    new_n24653_, new_n24654_, new_n24655_, new_n24656_, new_n24657_,
    new_n24658_, new_n24659_, new_n24660_, new_n24661_, new_n24662_,
    new_n24663_, new_n24664_, new_n24665_, new_n24666_, new_n24667_,
    new_n24668_, new_n24669_, new_n24670_, new_n24671_, new_n24672_,
    new_n24673_, new_n24674_, new_n24675_, new_n24676_, new_n24677_,
    new_n24678_, new_n24679_, new_n24680_, new_n24681_, new_n24682_,
    new_n24683_, new_n24684_, new_n24685_, new_n24686_, new_n24690_,
    new_n24691_, new_n24692_, new_n24701_, new_n24702_, new_n24703_,
    new_n24704_, new_n24705_, new_n24706_, new_n24707_, new_n24708_,
    new_n24709_, new_n24710_, new_n24711_, new_n24712_, new_n24713_,
    new_n24714_, new_n24715_, new_n24716_, new_n24717_, new_n24718_,
    new_n24719_, new_n24722_, new_n24723_, new_n24724_, new_n24725_,
    new_n24727_, new_n24728_, new_n24729_, new_n24730_, new_n24731_,
    new_n24732_, new_n24733_, new_n24734_, new_n24735_, new_n24736_,
    new_n24737_, new_n24738_, new_n24739_, new_n24740_, new_n24741_,
    new_n24742_, new_n24744_, new_n24745_, new_n24746_, new_n24747_,
    new_n24748_, new_n24749_, new_n24750_, new_n24751_, new_n24753_,
    new_n24754_, new_n24755_, new_n24756_, new_n24757_, new_n24758_,
    new_n24759_, new_n24760_, new_n24761_, new_n24762_, new_n24764_,
    new_n24765_, new_n24766_, new_n24767_, new_n24768_, new_n24769_,
    new_n24770_, new_n24771_, new_n24773_, new_n24774_, new_n24775_,
    new_n24776_, new_n24777_, new_n24778_, new_n24779_, new_n24780_,
    new_n24781_, new_n24782_, new_n24783_, new_n24784_, new_n24785_,
    new_n24786_, new_n24787_, new_n24788_, new_n24789_, new_n24790_,
    new_n24791_, new_n24792_, new_n24793_, new_n24794_, new_n24795_,
    new_n24796_, new_n24797_, new_n24798_, new_n24799_, new_n24800_,
    new_n24801_, new_n24802_, new_n24803_, new_n24804_, new_n24805_,
    new_n24806_, new_n24807_, new_n24808_, new_n24809_, new_n24810_,
    new_n24811_, new_n24812_, new_n24813_, new_n24814_, new_n24815_,
    new_n24816_, new_n24817_, new_n24818_, new_n24819_, new_n24822_,
    new_n24823_, new_n24824_, new_n24825_, new_n24826_, new_n24827_,
    new_n24828_, new_n24829_, new_n24830_, new_n24831_, new_n24832_,
    new_n24833_, new_n24834_, new_n24835_, new_n24836_, new_n24837_,
    new_n24838_, new_n24839_, new_n24840_, new_n24841_, new_n24842_,
    new_n24843_, new_n24844_, new_n24845_, new_n24846_, new_n24848_,
    new_n24849_, new_n24850_, new_n24851_, new_n24852_, new_n24853_,
    new_n24854_, new_n24855_, new_n24856_, new_n24857_, new_n24858_,
    new_n24859_, new_n24860_, new_n24861_, new_n24862_, new_n24863_,
    new_n24864_, new_n24865_, new_n24866_, new_n24867_, new_n24868_,
    new_n24869_, new_n24870_, new_n24871_, new_n24872_, new_n24873_,
    new_n24874_, new_n24875_, new_n24876_, new_n24877_, new_n24878_,
    new_n24879_, new_n24880_, new_n24881_, new_n24882_, new_n24883_,
    new_n24884_, new_n24885_, new_n24886_, new_n24887_, new_n24888_,
    new_n24889_, new_n24890_, new_n24891_, new_n24892_, new_n24893_,
    new_n24894_, new_n24895_, new_n24896_, new_n24897_, new_n24898_,
    new_n24899_, new_n24900_, new_n24901_, new_n24902_, new_n24903_,
    new_n24905_, new_n24906_, new_n24907_, new_n24908_, new_n24909_,
    new_n24910_, new_n24911_, new_n24912_, new_n24913_, new_n24914_,
    new_n24915_, new_n24916_, new_n24918_, new_n24919_, new_n24920_,
    new_n24921_, new_n24922_, new_n24923_, new_n24924_, new_n24925_,
    new_n24926_, new_n24927_, new_n24928_, new_n24930_, new_n24931_,
    new_n24932_, new_n24934_, new_n24935_, new_n24936_, new_n24937_,
    new_n24938_, new_n24939_, new_n24940_, new_n24941_, new_n24942_,
    new_n24943_, new_n24945_, new_n24946_, new_n24947_, new_n24948_,
    new_n24950_, new_n24951_, new_n24952_, new_n24953_, new_n24954_,
    new_n24955_, new_n24956_, new_n24957_, new_n24958_, new_n24959_,
    new_n24960_, new_n24961_, new_n24962_, new_n24963_, new_n24964_,
    new_n24965_, new_n24966_, new_n24967_, new_n24968_, new_n24969_,
    new_n24970_, new_n24971_, new_n24972_, new_n24973_, new_n24974_,
    new_n24975_, new_n24976_, new_n24977_, new_n24978_, new_n24979_,
    new_n24980_, new_n24981_, new_n24982_, new_n24983_, new_n24984_,
    new_n24985_, new_n24986_, new_n24987_, new_n24988_, new_n24989_,
    new_n24990_, new_n24991_, new_n24992_, new_n24993_, new_n24994_,
    new_n24995_, new_n24996_, new_n24997_, new_n24998_, new_n25000_,
    new_n25001_, new_n25002_, new_n25003_, new_n25004_, new_n25005_,
    new_n25006_, new_n25007_, new_n25008_, new_n25009_, new_n25010_,
    new_n25011_, new_n25012_, new_n25014_, new_n25015_, new_n25016_,
    new_n25017_, new_n25018_, new_n25019_, new_n25020_, new_n25021_,
    new_n25022_, new_n25023_, new_n25024_, new_n25025_, new_n25026_,
    new_n25027_, new_n25028_, new_n25029_, new_n25030_, new_n25031_,
    new_n25032_, new_n25033_, new_n25034_, new_n25035_, new_n25036_,
    new_n25037_, new_n25038_, new_n25039_, new_n25040_, new_n25041_,
    new_n25042_, new_n25043_, new_n25044_, new_n25045_, new_n25046_,
    new_n25047_, new_n25048_, new_n25049_, new_n25050_, new_n25051_,
    new_n25052_, new_n25053_, new_n25054_, new_n25055_, new_n25056_,
    new_n25057_, new_n25058_, new_n25059_, new_n25060_, new_n25061_,
    new_n25062_, new_n25063_, new_n25064_, new_n25065_, new_n25066_,
    new_n25067_, new_n25068_, new_n25069_, new_n25070_, new_n25071_,
    new_n25072_, new_n25073_, new_n25074_, new_n25075_, new_n25076_,
    new_n25077_, new_n25078_, new_n25079_, new_n25080_, new_n25081_,
    new_n25082_, new_n25083_, new_n25084_, new_n25085_, new_n25086_,
    new_n25087_, new_n25088_, new_n25089_, new_n25090_, new_n25091_,
    new_n25092_, new_n25093_, new_n25094_, new_n25095_, new_n25096_,
    new_n25097_, new_n25098_, new_n25099_, new_n25100_, new_n25101_,
    new_n25102_, new_n25103_, new_n25104_, new_n25105_, new_n25106_,
    new_n25107_, new_n25108_, new_n25109_, new_n25110_, new_n25111_,
    new_n25112_, new_n25113_, new_n25114_, new_n25115_, new_n25116_,
    new_n25117_, new_n25118_, new_n25119_, new_n25120_, new_n25121_,
    new_n25122_, new_n25123_, new_n25124_, new_n25125_, new_n25126_,
    new_n25127_, new_n25128_, new_n25129_, new_n25130_, new_n25131_,
    new_n25132_, new_n25133_, new_n25134_, new_n25135_, new_n25136_,
    new_n25137_, new_n25138_, new_n25139_, new_n25140_, new_n25141_,
    new_n25142_, new_n25143_, new_n25144_, new_n25145_, new_n25146_,
    new_n25147_, new_n25148_, new_n25149_, new_n25150_, new_n25151_,
    new_n25152_, new_n25153_, new_n25154_, new_n25155_, new_n25156_,
    new_n25157_, new_n25158_, new_n25159_, new_n25160_, new_n25161_,
    new_n25162_, new_n25163_, new_n25164_, new_n25165_, new_n25166_,
    new_n25167_, new_n25168_, new_n25169_, new_n25170_, new_n25171_,
    new_n25172_, new_n25173_, new_n25174_, new_n25175_, new_n25176_,
    new_n25177_, new_n25178_, new_n25179_, new_n25180_, new_n25181_,
    new_n25182_, new_n25183_, new_n25184_, new_n25185_, new_n25186_,
    new_n25187_, new_n25188_, new_n25189_, new_n25190_, new_n25191_,
    new_n25192_, new_n25193_, new_n25194_, new_n25195_, new_n25196_,
    new_n25197_, new_n25198_, new_n25199_, new_n25200_, new_n25201_,
    new_n25202_, new_n25203_, new_n25204_, new_n25205_, new_n25206_,
    new_n25207_, new_n25208_, new_n25209_, new_n25210_, new_n25211_,
    new_n25212_, new_n25213_, new_n25214_, new_n25215_, new_n25216_,
    new_n25217_, new_n25218_, new_n25219_, new_n25220_, new_n25221_,
    new_n25222_, new_n25223_, new_n25224_, new_n25225_, new_n25226_,
    new_n25227_, new_n25228_, new_n25229_, new_n25230_, new_n25231_,
    new_n25232_, new_n25233_, new_n25234_, new_n25235_, new_n25236_,
    new_n25237_, new_n25238_, new_n25239_, new_n25240_, new_n25241_,
    new_n25242_, new_n25243_, new_n25244_, new_n25245_, new_n25246_,
    new_n25247_, new_n25248_, new_n25249_, new_n25250_, new_n25251_,
    new_n25252_, new_n25253_, new_n25254_, new_n25255_, new_n25256_,
    new_n25257_, new_n25258_, new_n25259_, new_n25260_, new_n25261_,
    new_n25262_, new_n25263_, new_n25264_, new_n25265_, new_n25266_,
    new_n25267_, new_n25268_, new_n25270_, new_n25271_, new_n25272_,
    new_n25273_, new_n25274_, new_n25275_, new_n25276_, new_n25277_,
    new_n25278_, new_n25279_, new_n25280_, new_n25281_, new_n25282_,
    new_n25283_, new_n25284_, new_n25285_, new_n25286_, new_n25287_,
    new_n25288_, new_n25289_, new_n25290_, new_n25291_, new_n25292_,
    new_n25293_, new_n25294_, new_n25295_, new_n25296_, new_n25297_,
    new_n25298_, new_n25299_, new_n25300_, new_n25301_, new_n25302_,
    new_n25303_, new_n25304_, new_n25305_, new_n25306_, new_n25307_,
    new_n25308_, new_n25309_, new_n25310_, new_n25311_, new_n25312_,
    new_n25313_, new_n25314_, new_n25315_, new_n25316_, new_n25317_,
    new_n25318_, new_n25319_, new_n25320_, new_n25321_, new_n25326_,
    new_n25327_, new_n25328_, new_n25329_, new_n25330_, new_n25331_,
    new_n25332_, new_n25333_, new_n25334_, new_n25335_, new_n25336_,
    new_n25337_, new_n25338_, new_n25339_, new_n25340_, new_n25341_,
    new_n25342_, new_n25343_, new_n25344_, new_n25345_, new_n25346_,
    new_n25347_, new_n25348_, new_n25349_, new_n25350_, new_n25351_,
    new_n25352_, new_n25353_, new_n25354_, new_n25355_, new_n25356_,
    new_n25357_, new_n25358_, new_n25359_, new_n25360_, new_n25361_,
    new_n25362_, new_n25363_, new_n25364_, new_n25365_, new_n25366_,
    new_n25367_, new_n25368_, new_n25369_, new_n25370_, new_n25372_,
    new_n25373_, new_n25374_, new_n25375_, new_n25376_, new_n25377_,
    new_n25378_, new_n25379_, new_n25381_, new_n25382_, new_n25383_,
    new_n25384_, new_n25385_, new_n25386_, new_n25387_, new_n25388_,
    new_n25389_, new_n25390_, new_n25391_, new_n25392_, new_n25393_,
    new_n25394_, new_n25395_, new_n25396_, new_n25397_, new_n25398_,
    new_n25399_, new_n25400_, new_n25401_, new_n25402_, new_n25403_,
    new_n25404_, new_n25405_, new_n25406_, new_n25407_, new_n25408_,
    new_n25409_, new_n25410_, new_n25411_, new_n25412_, new_n25413_,
    new_n25414_, new_n25415_, new_n25416_, new_n25417_, new_n25418_,
    new_n25419_, new_n25420_, new_n25421_, new_n25422_, new_n25423_,
    new_n25424_, new_n25425_, new_n25426_, new_n25427_, new_n25428_,
    new_n25429_, new_n25430_, new_n25431_, new_n25432_, new_n25433_,
    new_n25434_, new_n25435_, new_n25436_, new_n25437_, new_n25438_,
    new_n25439_, new_n25440_, new_n25441_, new_n25442_, new_n25443_,
    new_n25444_, new_n25445_, new_n25446_, new_n25447_, new_n25448_,
    new_n25449_, new_n25450_, new_n25451_, new_n25452_, new_n25453_,
    new_n25454_, new_n25455_, new_n25456_, new_n25457_, new_n25458_,
    new_n25459_, new_n25460_, new_n25461_, new_n25462_, new_n25463_,
    new_n25464_, new_n25465_, new_n25466_, new_n25467_, new_n25468_,
    new_n25469_, new_n25470_, new_n25471_, new_n25472_, new_n25473_,
    new_n25474_, new_n25475_, new_n25476_, new_n25477_, new_n25478_,
    new_n25479_, new_n25480_, new_n25481_, new_n25482_, new_n25483_,
    new_n25484_, new_n25485_, new_n25486_, new_n25487_, new_n25488_,
    new_n25489_, new_n25490_, new_n25491_, new_n25492_, new_n25493_,
    new_n25494_, new_n25495_, new_n25496_, new_n25497_, new_n25498_,
    new_n25499_, new_n25500_, new_n25501_, new_n25502_, new_n25503_,
    new_n25504_, new_n25505_, new_n25506_, new_n25507_, new_n25508_,
    new_n25509_, new_n25510_, new_n25511_, new_n25512_, new_n25513_,
    new_n25514_, new_n25515_, new_n25516_, new_n25517_, new_n25518_,
    new_n25519_, new_n25520_, new_n25521_, new_n25522_, new_n25523_,
    new_n25524_, new_n25525_, new_n25526_, new_n25527_, new_n25528_,
    new_n25529_, new_n25530_, new_n25531_, new_n25532_, new_n25533_,
    new_n25534_, new_n25535_, new_n25536_, new_n25537_, new_n25538_,
    new_n25539_, new_n25540_, new_n25541_, new_n25542_, new_n25543_,
    new_n25544_, new_n25545_, new_n25546_, new_n25547_, new_n25548_,
    new_n25549_, new_n25550_, new_n25551_, new_n25552_, new_n25553_,
    new_n25554_, new_n25555_, new_n25556_, new_n25557_, new_n25558_,
    new_n25559_, new_n25560_, new_n25561_, new_n25562_, new_n25563_,
    new_n25564_, new_n25565_, new_n25566_, new_n25567_, new_n25568_,
    new_n25569_, new_n25570_, new_n25571_, new_n25572_, new_n25573_,
    new_n25574_, new_n25575_, new_n25576_, new_n25577_, new_n25578_,
    new_n25579_, new_n25580_, new_n25581_, new_n25582_, new_n25583_,
    new_n25584_, new_n25585_, new_n25586_, new_n25587_, new_n25588_,
    new_n25589_, new_n25590_, new_n25591_, new_n25592_, new_n25593_,
    new_n25594_, new_n25595_, new_n25596_, new_n25597_, new_n25598_,
    new_n25599_, new_n25600_, new_n25601_, new_n25602_, new_n25603_,
    new_n25604_, new_n25605_, new_n25606_, new_n25607_, new_n25608_,
    new_n25609_, new_n25610_, new_n25611_, new_n25612_, new_n25613_,
    new_n25614_, new_n25615_, new_n25616_, new_n25617_, new_n25618_,
    new_n25619_, new_n25620_, new_n25621_, new_n25622_, new_n25623_,
    new_n25624_, new_n25625_, new_n25626_, new_n25627_, new_n25628_,
    new_n25629_, new_n25630_, new_n25631_, new_n25632_, new_n25633_,
    new_n25634_, new_n25635_, new_n25636_, new_n25637_, new_n25638_,
    new_n25639_, new_n25640_, new_n25641_, new_n25642_, new_n25643_,
    new_n25644_, new_n25645_, new_n25646_, new_n25647_, new_n25648_,
    new_n25649_, new_n25650_, new_n25651_, new_n25652_, new_n25653_,
    new_n25654_, new_n25655_, new_n25656_, new_n25657_, new_n25658_,
    new_n25659_, new_n25660_, new_n25661_, new_n25662_, new_n25663_,
    new_n25664_, new_n25665_, new_n25666_, new_n25667_, new_n25668_,
    new_n25669_, new_n25670_, new_n25671_, new_n25672_, new_n25673_,
    new_n25674_, new_n25675_, new_n25676_, new_n25677_, new_n25678_,
    new_n25679_, new_n25680_, new_n25681_, new_n25682_, new_n25683_,
    new_n25684_, new_n25685_, new_n25686_, new_n25687_, new_n25688_,
    new_n25689_, new_n25690_, new_n25691_, new_n25692_, new_n25693_,
    new_n25694_, new_n25695_, new_n25696_, new_n25697_, new_n25698_,
    new_n25699_, new_n25700_, new_n25701_, new_n25702_, new_n25703_,
    new_n25704_, new_n25705_, new_n25706_, new_n25707_, new_n25708_,
    new_n25709_, new_n25710_, new_n25711_, new_n25712_, new_n25713_,
    new_n25714_, new_n25715_, new_n25716_, new_n25717_, new_n25718_,
    new_n25719_, new_n25720_, new_n25721_, new_n25722_, new_n25723_,
    new_n25726_, new_n25727_, new_n25728_, new_n25729_, new_n25730_,
    new_n25731_, new_n25732_, new_n25733_, new_n25735_, new_n25736_,
    new_n25737_, new_n25738_, new_n25739_, new_n25740_, new_n25741_,
    new_n25742_, new_n25743_, new_n25744_, new_n25745_, new_n25746_,
    new_n25747_, new_n25748_, new_n25749_, new_n25750_, new_n25751_,
    new_n25752_, new_n25753_, new_n25754_, new_n25755_, new_n25756_,
    new_n25757_, new_n25758_, new_n25759_, new_n25760_, new_n25761_,
    new_n25762_, new_n25763_, new_n25764_, new_n25765_, new_n25766_,
    new_n25767_, new_n25768_, new_n25769_, new_n25770_, new_n25771_,
    new_n25772_, new_n25773_, new_n25774_, new_n25775_, new_n25776_,
    new_n25777_, new_n25778_, new_n25779_, new_n25780_, new_n25781_,
    new_n25782_, new_n25783_, new_n25784_, new_n25785_, new_n25786_,
    new_n25787_, new_n25788_, new_n25789_, new_n25790_, new_n25791_,
    new_n25792_, new_n25793_, new_n25794_, new_n25795_, new_n25796_,
    new_n25797_, new_n25798_, new_n25799_, new_n25800_, new_n25801_,
    new_n25802_, new_n25803_, new_n25804_, new_n25805_, new_n25806_,
    new_n25807_, new_n25808_, new_n25809_, new_n25810_, new_n25811_,
    new_n25812_, new_n25813_, new_n25814_, new_n25815_, new_n25816_,
    new_n25817_, new_n25818_, new_n25819_, new_n25821_, new_n25822_,
    new_n25823_, new_n25824_, new_n25825_, new_n25826_, new_n25827_,
    new_n25828_, new_n25829_, new_n25830_, new_n25831_, new_n25832_,
    new_n25833_, new_n25834_, new_n25835_, new_n25836_, new_n25837_,
    new_n25838_, new_n25839_, new_n25840_, new_n25841_, new_n25842_,
    new_n25843_, new_n25844_, new_n25845_, new_n25846_, new_n25847_,
    new_n25848_, new_n25849_, new_n25850_, new_n25851_, new_n25852_,
    new_n25853_, new_n25854_, new_n25855_, new_n25856_, new_n25857_,
    new_n25858_, new_n25859_, new_n25860_, new_n25861_, new_n25862_,
    new_n25863_, new_n25864_, new_n25865_, new_n25866_, new_n25867_,
    new_n25868_, new_n25869_, new_n25870_, new_n25871_, new_n25872_,
    new_n25873_, new_n25874_, new_n25875_, new_n25876_, new_n25877_,
    new_n25878_, new_n25879_, new_n25880_, new_n25881_, new_n25882_,
    new_n25883_, new_n25884_, new_n25885_, new_n25886_, new_n25887_,
    new_n25888_, new_n25889_, new_n25890_, new_n25891_, new_n25892_,
    new_n25893_, new_n25894_, new_n25895_, new_n25896_, new_n25897_,
    new_n25898_, new_n25899_, new_n25900_, new_n25901_, new_n25902_,
    new_n25903_, new_n25904_, new_n25905_, new_n25906_, new_n25907_,
    new_n25908_, new_n25909_, new_n25910_, new_n25911_, new_n25912_,
    new_n25913_, new_n25914_, new_n25915_, new_n25916_, new_n25917_,
    new_n25918_, new_n25919_, new_n25920_, new_n25921_, new_n25922_,
    new_n25923_, new_n25924_, new_n25925_, new_n25926_, new_n25927_,
    new_n25928_, new_n25929_, new_n25930_, new_n25931_, new_n25932_,
    new_n25933_, new_n25934_, new_n25935_, new_n25936_, new_n25937_,
    new_n25938_, new_n25939_, new_n25940_, new_n25941_, new_n25942_,
    new_n25943_, new_n25944_, new_n25945_, new_n25946_, new_n25947_,
    new_n25948_, new_n25949_, new_n25950_, new_n25951_, new_n25952_,
    new_n25953_, new_n25954_, new_n25955_, new_n25956_, new_n25957_,
    new_n25958_, new_n25959_, new_n25960_, new_n25961_, new_n25962_,
    new_n25963_, new_n25964_, new_n25965_, new_n25966_, new_n25967_,
    new_n25968_, new_n25969_, new_n25970_, new_n25971_, new_n25972_,
    new_n25973_, new_n25974_, new_n25975_, new_n25976_, new_n25977_,
    new_n25978_, new_n25979_, new_n25980_, new_n25981_, new_n25982_,
    new_n25983_, new_n25984_, new_n25985_, new_n25986_, new_n25987_,
    new_n25988_, new_n25989_, new_n25990_, new_n25991_, new_n25992_,
    new_n25993_, new_n25994_, new_n25995_, new_n25996_, new_n25997_,
    new_n25998_, new_n25999_, new_n26000_, new_n26001_, new_n26002_,
    new_n26003_, new_n26004_, new_n26005_, new_n26006_, new_n26007_,
    new_n26008_, new_n26009_, new_n26010_, new_n26011_, new_n26012_,
    new_n26013_, new_n26014_, new_n26015_, new_n26016_, new_n26017_,
    new_n26018_, new_n26019_, new_n26020_, new_n26021_, new_n26022_,
    new_n26023_, new_n26024_, new_n26025_, new_n26026_, new_n26027_,
    new_n26028_, new_n26029_, new_n26030_, new_n26031_, new_n26032_,
    new_n26033_, new_n26034_, new_n26035_, new_n26036_, new_n26037_,
    new_n26038_, new_n26039_, new_n26040_, new_n26041_, new_n26042_,
    new_n26043_, new_n26044_, new_n26045_, new_n26046_, new_n26047_,
    new_n26048_, new_n26049_, new_n26050_, new_n26051_, new_n26052_,
    new_n26053_, new_n26054_, new_n26055_, new_n26056_, new_n26057_,
    new_n26058_, new_n26059_, new_n26060_, new_n26061_, new_n26062_,
    new_n26063_, new_n26064_, new_n26065_, new_n26066_, new_n26067_,
    new_n26068_, new_n26069_, new_n26070_, new_n26071_, new_n26075_,
    new_n26076_, new_n26077_, new_n26078_, new_n26079_, new_n26080_,
    new_n26081_, new_n26082_, new_n26083_, new_n26085_, new_n26086_,
    new_n26087_, new_n26088_, new_n26089_, new_n26090_, new_n26091_,
    new_n26092_, new_n26093_, new_n26094_, new_n26095_, new_n26096_,
    new_n26097_, new_n26098_, new_n26099_, new_n26100_, new_n26101_,
    new_n26102_, new_n26103_, new_n26105_, new_n26106_, new_n26107_,
    new_n26108_, new_n26109_, new_n26110_, new_n26111_, new_n26112_,
    new_n26113_, new_n26114_, new_n26115_, new_n26116_, new_n26117_,
    new_n26118_, new_n26119_, new_n26120_, new_n26121_, new_n26122_,
    new_n26123_, new_n26124_, new_n26125_, new_n26126_, new_n26127_,
    new_n26128_, new_n26129_, new_n26130_, new_n26131_, new_n26132_,
    new_n26133_, new_n26134_, new_n26135_, new_n26136_, new_n26137_,
    new_n26138_, new_n26139_, new_n26140_, new_n26141_, new_n26142_,
    new_n26143_, new_n26144_, new_n26145_, new_n26146_, new_n26147_,
    new_n26148_, new_n26149_, new_n26151_, new_n26153_, new_n26154_,
    new_n26155_, new_n26156_, new_n26157_, new_n26158_, new_n26159_,
    new_n26160_, new_n26161_, new_n26162_, new_n26163_, new_n26164_,
    new_n26165_, new_n26166_, new_n26167_, new_n26168_, new_n26169_,
    new_n26170_, new_n26171_, new_n26172_, new_n26173_, new_n26174_,
    new_n26175_, new_n26176_, new_n26177_, new_n26178_, new_n26179_,
    new_n26180_, new_n26181_, new_n26183_, new_n26184_, new_n26185_,
    new_n26186_, new_n26187_, new_n26188_, new_n26189_, new_n26190_,
    new_n26191_, new_n26192_, new_n26193_, new_n26194_, new_n26195_,
    new_n26196_, new_n26197_, new_n26198_, new_n26199_, new_n26200_,
    new_n26201_, new_n26203_, new_n26204_, new_n26205_, new_n26206_,
    new_n26207_, new_n26208_, new_n26209_, new_n26210_, new_n26212_,
    new_n26213_, new_n26214_, new_n26215_, new_n26216_, new_n26217_,
    new_n26218_, new_n26219_, new_n26220_, new_n26221_, new_n26222_,
    new_n26223_, new_n26224_, new_n26225_, new_n26226_, new_n26227_,
    new_n26228_, new_n26229_, new_n26230_, new_n26231_, new_n26232_,
    new_n26233_, new_n26234_, new_n26235_, new_n26236_, new_n26237_,
    new_n26238_, new_n26239_, new_n26240_, new_n26241_, new_n26242_,
    new_n26243_, new_n26244_, new_n26245_, new_n26246_, new_n26247_,
    new_n26248_, new_n26249_, new_n26250_, new_n26251_, new_n26252_,
    new_n26253_, new_n26254_, new_n26255_, new_n26256_, new_n26258_,
    new_n26259_, new_n26260_, new_n26261_, new_n26262_, new_n26264_,
    new_n26265_, new_n26266_, new_n26267_, new_n26268_, new_n26269_,
    new_n26270_, new_n26271_, new_n26272_, new_n26273_, new_n26274_,
    new_n26275_, new_n26276_, new_n26277_, new_n26278_, new_n26279_,
    new_n26280_, new_n26281_, new_n26282_, new_n26283_, new_n26284_,
    new_n26285_, new_n26286_, new_n26287_, new_n26288_, new_n26289_,
    new_n26290_, new_n26291_, new_n26292_, new_n26293_, new_n26294_,
    new_n26295_, new_n26296_, new_n26297_, new_n26298_, new_n26299_,
    new_n26300_, new_n26301_, new_n26302_, new_n26303_, new_n26304_,
    new_n26305_, new_n26307_, new_n26308_, new_n26309_, new_n26310_,
    new_n26311_, new_n26312_, new_n26313_, new_n26314_, new_n26315_,
    new_n26316_, new_n26317_, new_n26318_, new_n26319_, new_n26320_,
    new_n26321_, new_n26322_, new_n26323_, new_n26324_, new_n26325_,
    new_n26326_, new_n26327_, new_n26328_, new_n26329_, new_n26330_,
    new_n26331_, new_n26332_, new_n26333_, new_n26334_, new_n26335_,
    new_n26336_, new_n26337_, new_n26338_, new_n26339_, new_n26340_,
    new_n26341_, new_n26342_, new_n26343_, new_n26344_, new_n26345_,
    new_n26346_, new_n26347_, new_n26348_, new_n26349_, new_n26350_,
    new_n26351_, new_n26352_, new_n26353_, new_n26354_, new_n26355_,
    new_n26356_, new_n26357_, new_n26358_, new_n26359_, new_n26360_,
    new_n26361_, new_n26362_, new_n26363_, new_n26364_, new_n26365_,
    new_n26366_, new_n26367_, new_n26368_, new_n26369_, new_n26370_,
    new_n26371_, new_n26372_, new_n26373_, new_n26374_, new_n26375_,
    new_n26376_, new_n26377_, new_n26378_, new_n26379_, new_n26380_,
    new_n26381_, new_n26382_, new_n26383_, new_n26384_, new_n26385_,
    new_n26386_, new_n26387_, new_n26388_, new_n26389_, new_n26390_,
    new_n26391_, new_n26392_, new_n26393_, new_n26394_, new_n26395_,
    new_n26396_, new_n26397_, new_n26398_, new_n26399_, new_n26400_,
    new_n26401_, new_n26402_, new_n26403_, new_n26404_, new_n26405_,
    new_n26406_, new_n26407_, new_n26408_, new_n26409_, new_n26410_,
    new_n26411_, new_n26412_, new_n26413_, new_n26414_, new_n26415_,
    new_n26416_, new_n26417_, new_n26418_, new_n26419_, new_n26420_,
    new_n26421_, new_n26422_, new_n26423_, new_n26424_, new_n26425_,
    new_n26426_, new_n26427_, new_n26428_, new_n26429_, new_n26430_,
    new_n26431_, new_n26432_, new_n26433_, new_n26434_, new_n26435_,
    new_n26436_, new_n26437_, new_n26438_, new_n26439_, new_n26440_,
    new_n26441_, new_n26442_, new_n26443_, new_n26444_, new_n26445_,
    new_n26446_, new_n26447_, new_n26448_, new_n26449_, new_n26450_,
    new_n26451_, new_n26452_, new_n26453_, new_n26454_, new_n26455_,
    new_n26456_, new_n26457_, new_n26458_, new_n26459_, new_n26460_,
    new_n26461_, new_n26462_, new_n26463_, new_n26464_, new_n26465_,
    new_n26466_, new_n26467_, new_n26468_, new_n26469_, new_n26470_,
    new_n26471_, new_n26472_, new_n26473_, new_n26474_, new_n26475_,
    new_n26476_, new_n26477_, new_n26478_, new_n26479_, new_n26480_,
    new_n26482_, new_n26483_, new_n26484_, new_n26485_, new_n26486_,
    new_n26487_, new_n26488_, new_n26489_, new_n26490_, new_n26491_,
    new_n26492_, new_n26493_, new_n26494_, new_n26495_, new_n26496_,
    new_n26497_, new_n26498_, new_n26499_, new_n26500_, new_n26501_,
    new_n26502_, new_n26503_, new_n26504_, new_n26505_, new_n26506_,
    new_n26507_, new_n26508_, new_n26509_, new_n26510_, new_n26511_,
    new_n26512_, new_n26513_, new_n26514_, new_n26515_, new_n26516_,
    new_n26517_, new_n26518_, new_n26519_, new_n26520_, new_n26521_,
    new_n26522_, new_n26523_, new_n26524_, new_n26525_, new_n26526_,
    new_n26527_, new_n26528_, new_n26529_, new_n26530_, new_n26531_,
    new_n26532_, new_n26533_, new_n26534_, new_n26535_, new_n26536_,
    new_n26537_, new_n26538_, new_n26539_, new_n26540_, new_n26541_,
    new_n26542_, new_n26543_, new_n26544_, new_n26545_, new_n26546_,
    new_n26547_, new_n26548_, new_n26549_, new_n26550_, new_n26551_,
    new_n26552_, new_n26553_, new_n26554_, new_n26555_, new_n26556_,
    new_n26557_, new_n26558_, new_n26559_, new_n26560_, new_n26561_,
    new_n26562_, new_n26563_, new_n26564_, new_n26565_, new_n26566_,
    new_n26567_, new_n26568_, new_n26569_, new_n26570_, new_n26571_,
    new_n26572_, new_n26573_, new_n26574_, new_n26575_, new_n26576_,
    new_n26577_, new_n26578_, new_n26579_, new_n26580_, new_n26581_,
    new_n26582_, new_n26583_, new_n26584_, new_n26585_, new_n26586_,
    new_n26587_, new_n26588_, new_n26589_, new_n26590_, new_n26591_,
    new_n26592_, new_n26593_, new_n26594_, new_n26595_, new_n26596_,
    new_n26597_, new_n26598_, new_n26599_, new_n26600_, new_n26601_,
    new_n26602_, new_n26604_, new_n26605_, new_n26606_, new_n26607_,
    new_n26608_, new_n26609_, new_n26610_, new_n26611_, new_n26612_,
    new_n26613_, new_n26614_, new_n26615_, new_n26616_, new_n26617_,
    new_n26618_, new_n26619_, new_n26620_, new_n26621_, new_n26622_,
    new_n26623_, new_n26624_, new_n26625_, new_n26626_, new_n26627_,
    new_n26628_, new_n26629_, new_n26630_, new_n26631_, new_n26632_,
    new_n26633_, new_n26634_, new_n26635_, new_n26636_, new_n26637_,
    new_n26638_, new_n26639_, new_n26640_, new_n26641_, new_n26642_,
    new_n26643_, new_n26644_, new_n26645_, new_n26646_, new_n26647_,
    new_n26648_, new_n26649_, new_n26650_, new_n26651_, new_n26652_,
    new_n26653_, new_n26654_, new_n26655_, new_n26656_, new_n26657_,
    new_n26658_, new_n26659_, new_n26660_, new_n26661_, new_n26662_,
    new_n26663_, new_n26664_, new_n26665_, new_n26666_, new_n26667_,
    new_n26668_, new_n26669_, new_n26670_, new_n26671_, new_n26672_,
    new_n26673_, new_n26674_, new_n26675_, new_n26676_, new_n26677_,
    new_n26678_, new_n26679_, new_n26680_, new_n26681_, new_n26682_,
    new_n26683_, new_n26684_, new_n26685_, new_n26686_, new_n26687_,
    new_n26688_, new_n26689_, new_n26690_, new_n26691_, new_n26692_,
    new_n26693_, new_n26694_, new_n26695_, new_n26696_, new_n26697_,
    new_n26698_, new_n26699_, new_n26700_, new_n26701_, new_n26702_,
    new_n26703_, new_n26704_, new_n26705_, new_n26706_, new_n26707_,
    new_n26708_, new_n26709_, new_n26710_, new_n26711_, new_n26712_,
    new_n26713_, new_n26714_, new_n26715_, new_n26716_, new_n26717_,
    new_n26718_, new_n26719_, new_n26720_, new_n26721_, new_n26722_,
    new_n26723_, new_n26724_, new_n26725_, new_n26726_, new_n26727_,
    new_n26728_, new_n26729_, new_n26730_, new_n26731_, new_n26732_,
    new_n26733_, new_n26734_, new_n26735_, new_n26736_, new_n26737_,
    new_n26738_, new_n26739_, new_n26740_, new_n26741_, new_n26742_,
    new_n26743_, new_n26744_, new_n26745_, new_n26746_, new_n26747_,
    new_n26748_, new_n26749_, new_n26750_, new_n26751_, new_n26752_,
    new_n26753_, new_n26754_, new_n26755_, new_n26756_, new_n26757_,
    new_n26758_, new_n26759_, new_n26760_, new_n26762_, new_n26763_,
    new_n26764_, new_n26765_, new_n26766_, new_n26767_, new_n26768_,
    new_n26769_, new_n26770_, new_n26771_, new_n26772_, new_n26773_,
    new_n26774_, new_n26775_, new_n26776_, new_n26777_, new_n26778_,
    new_n26779_, new_n26780_, new_n26781_, new_n26782_, new_n26783_,
    new_n26784_, new_n26785_, new_n26786_, new_n26787_, new_n26788_,
    new_n26789_, new_n26790_, new_n26791_, new_n26792_, new_n26793_,
    new_n26794_, new_n26795_, new_n26796_, new_n26797_, new_n26798_,
    new_n26799_, new_n26800_, new_n26801_, new_n26802_, new_n26803_,
    new_n26804_, new_n26805_, new_n26806_, new_n26807_, new_n26808_,
    new_n26809_, new_n26810_, new_n26811_, new_n26812_, new_n26813_,
    new_n26814_, new_n26815_, new_n26816_, new_n26817_, new_n26818_,
    new_n26819_, new_n26820_, new_n26821_, new_n26822_, new_n26823_,
    new_n26824_, new_n26825_, new_n26827_, new_n26828_, new_n26829_,
    new_n26830_, new_n26831_, new_n26832_, new_n26833_, new_n26834_,
    new_n26835_, new_n26836_, new_n26837_, new_n26838_, new_n26839_,
    new_n26840_, new_n26841_, new_n26842_, new_n26843_, new_n26844_,
    new_n26845_, new_n26846_, new_n26847_, new_n26848_, new_n26849_,
    new_n26850_, new_n26851_, new_n26852_, new_n26853_, new_n26854_,
    new_n26855_, new_n26856_, new_n26857_, new_n26858_, new_n26859_,
    new_n26860_, new_n26861_, new_n26862_, new_n26863_, new_n26864_,
    new_n26865_, new_n26866_, new_n26867_, new_n26868_, new_n26869_,
    new_n26870_, new_n26871_, new_n26872_, new_n26873_, new_n26874_,
    new_n26875_, new_n26876_, new_n26877_, new_n26878_, new_n26879_,
    new_n26880_, new_n26881_, new_n26882_, new_n26883_, new_n26884_,
    new_n26885_, new_n26886_, new_n26887_, new_n26888_, new_n26889_,
    new_n26890_, new_n26891_, new_n26892_, new_n26893_, new_n26894_,
    new_n26895_, new_n26896_, new_n26897_, new_n26898_, new_n26899_,
    new_n26900_, new_n26901_, new_n26902_, new_n26903_, new_n26904_,
    new_n26905_, new_n26906_, new_n26907_, new_n26908_, new_n26909_,
    new_n26910_, new_n26911_, new_n26912_, new_n26913_, new_n26914_,
    new_n26915_, new_n26916_, new_n26917_, new_n26918_, new_n26919_,
    new_n26920_, new_n26921_, new_n26922_, new_n26923_, new_n26924_,
    new_n26925_, new_n26926_, new_n26927_, new_n26928_, new_n26929_,
    new_n26930_, new_n26931_, new_n26932_, new_n26933_, new_n26934_,
    new_n26935_, new_n26936_, new_n26937_, new_n26938_, new_n26939_,
    new_n26940_, new_n26941_, new_n26942_, new_n26943_, new_n26944_,
    new_n26945_, new_n26946_, new_n26947_, new_n26948_, new_n26949_,
    new_n26950_, new_n26951_, new_n26952_, new_n26953_, new_n26954_,
    new_n26955_, new_n26956_, new_n26957_, new_n26958_, new_n26959_,
    new_n26960_, new_n26961_, new_n26962_, new_n26963_, new_n26964_,
    new_n26965_, new_n26966_, new_n26967_, new_n26968_, new_n26969_,
    new_n26970_, new_n26971_, new_n26973_, new_n26974_, new_n26975_,
    new_n26976_, new_n26977_, new_n26978_, new_n26980_, new_n26981_,
    new_n26982_, new_n26983_, new_n26984_, new_n26985_, new_n26986_,
    new_n26987_, new_n26988_, new_n26989_, new_n26990_, new_n26991_,
    new_n26992_, new_n26993_, new_n26994_, new_n26995_, new_n26996_,
    new_n26997_, new_n26998_, new_n26999_, new_n27000_, new_n27001_,
    new_n27002_, new_n27003_, new_n27004_, new_n27005_, new_n27006_,
    new_n27007_, new_n27008_, new_n27009_, new_n27010_, new_n27011_,
    new_n27012_, new_n27013_, new_n27014_, new_n27015_, new_n27016_,
    new_n27017_, new_n27018_, new_n27019_, new_n27020_, new_n27021_,
    new_n27022_, new_n27023_, new_n27024_, new_n27025_, new_n27026_,
    new_n27027_, new_n27028_, new_n27029_, new_n27030_, new_n27031_,
    new_n27032_, new_n27033_, new_n27034_, new_n27035_, new_n27036_,
    new_n27037_, new_n27038_, new_n27039_, new_n27040_, new_n27041_,
    new_n27042_, new_n27043_, new_n27044_, new_n27045_, new_n27046_,
    new_n27047_, new_n27048_, new_n27049_, new_n27050_, new_n27051_,
    new_n27052_, new_n27053_, new_n27054_, new_n27055_, new_n27056_,
    new_n27057_, new_n27058_, new_n27059_, new_n27060_, new_n27061_,
    new_n27062_, new_n27063_, new_n27064_, new_n27065_, new_n27066_,
    new_n27067_, new_n27068_, new_n27069_, new_n27070_, new_n27071_,
    new_n27072_, new_n27073_, new_n27074_, new_n27075_, new_n27076_,
    new_n27077_, new_n27078_, new_n27079_, new_n27080_, new_n27081_,
    new_n27082_, new_n27083_, new_n27084_, new_n27085_, new_n27086_,
    new_n27087_, new_n27088_, new_n27089_, new_n27090_, new_n27091_,
    new_n27092_, new_n27093_, new_n27094_, new_n27095_, new_n27096_,
    new_n27097_, new_n27098_, new_n27099_, new_n27100_, new_n27101_,
    new_n27102_, new_n27103_, new_n27104_, new_n27105_, new_n27106_,
    new_n27107_, new_n27108_, new_n27109_, new_n27110_, new_n27111_,
    new_n27112_, new_n27113_, new_n27114_, new_n27115_, new_n27116_,
    new_n27117_, new_n27118_, new_n27119_, new_n27120_, new_n27121_,
    new_n27122_, new_n27123_, new_n27124_, new_n27125_, new_n27126_,
    new_n27127_, new_n27128_, new_n27129_, new_n27130_, new_n27131_,
    new_n27132_, new_n27133_, new_n27134_, new_n27135_, new_n27136_,
    new_n27137_, new_n27138_, new_n27139_, new_n27140_, new_n27142_,
    new_n27143_, new_n27144_, new_n27145_, new_n27146_, new_n27147_,
    new_n27148_, new_n27149_, new_n27150_, new_n27151_, new_n27152_,
    new_n27153_, new_n27154_, new_n27155_, new_n27156_, new_n27157_,
    new_n27158_, new_n27159_, new_n27160_, new_n27161_, new_n27162_,
    new_n27163_, new_n27164_, new_n27165_, new_n27166_, new_n27167_,
    new_n27168_, new_n27169_, new_n27170_, new_n27171_, new_n27172_,
    new_n27173_, new_n27174_, new_n27175_, new_n27176_, new_n27177_,
    new_n27178_, new_n27179_, new_n27180_, new_n27181_, new_n27182_,
    new_n27183_, new_n27184_, new_n27185_, new_n27186_, new_n27187_,
    new_n27188_, new_n27189_, new_n27190_, new_n27191_, new_n27192_,
    new_n27193_, new_n27194_, new_n27195_, new_n27196_, new_n27197_,
    new_n27198_, new_n27199_, new_n27200_, new_n27201_, new_n27202_,
    new_n27203_, new_n27204_, new_n27205_, new_n27206_, new_n27207_,
    new_n27208_, new_n27209_, new_n27210_, new_n27211_, new_n27212_,
    new_n27213_, new_n27214_, new_n27215_, new_n27216_, new_n27217_,
    new_n27218_, new_n27219_, new_n27220_, new_n27221_, new_n27222_,
    new_n27223_, new_n27224_, new_n27225_, new_n27226_, new_n27227_,
    new_n27228_, new_n27229_, new_n27230_, new_n27231_, new_n27232_,
    new_n27233_, new_n27234_, new_n27235_, new_n27236_, new_n27237_,
    new_n27238_, new_n27239_, new_n27240_, new_n27241_, new_n27242_,
    new_n27243_, new_n27244_, new_n27245_, new_n27246_, new_n27247_,
    new_n27248_, new_n27249_, new_n27250_, new_n27251_, new_n27252_,
    new_n27253_, new_n27254_, new_n27255_, new_n27256_, new_n27257_,
    new_n27258_, new_n27259_, new_n27260_, new_n27261_, new_n27262_,
    new_n27263_, new_n27264_, new_n27265_, new_n27266_, new_n27267_,
    new_n27268_, new_n27269_, new_n27270_, new_n27271_, new_n27272_,
    new_n27273_, new_n27274_, new_n27275_, new_n27276_, new_n27277_,
    new_n27278_, new_n27281_, new_n27282_, new_n27283_, new_n27284_,
    new_n27285_, new_n27286_, new_n27287_, new_n27288_, new_n27289_,
    new_n27290_, new_n27291_, new_n27292_, new_n27293_, new_n27294_,
    new_n27295_, new_n27296_, new_n27297_, new_n27298_, new_n27299_,
    new_n27300_, new_n27301_, new_n27302_, new_n27303_, new_n27304_,
    new_n27305_, new_n27306_, new_n27307_, new_n27308_, new_n27309_,
    new_n27310_, new_n27311_, new_n27312_, new_n27313_, new_n27314_,
    new_n27315_, new_n27316_, new_n27317_, new_n27318_, new_n27319_,
    new_n27320_, new_n27321_, new_n27322_, new_n27323_, new_n27324_,
    new_n27325_, new_n27326_, new_n27327_, new_n27328_, new_n27329_,
    new_n27330_, new_n27331_, new_n27332_, new_n27333_, new_n27334_,
    new_n27335_, new_n27336_, new_n27337_, new_n27338_, new_n27342_,
    new_n27343_, new_n27344_, new_n27345_, new_n27346_, new_n27347_,
    new_n27348_, new_n27349_, new_n27350_, new_n27351_, new_n27352_,
    new_n27353_, new_n27354_, new_n27355_, new_n27356_, new_n27357_,
    new_n27358_, new_n27359_, new_n27360_, new_n27361_, new_n27362_,
    new_n27363_, new_n27364_, new_n27365_, new_n27366_, new_n27367_,
    new_n27368_, new_n27369_, new_n27370_, new_n27371_, new_n27372_,
    new_n27373_, new_n27374_, new_n27375_, new_n27376_, new_n27377_,
    new_n27378_, new_n27379_, new_n27380_, new_n27381_, new_n27382_,
    new_n27383_, new_n27384_, new_n27385_, new_n27386_, new_n27387_,
    new_n27388_, new_n27389_, new_n27390_, new_n27391_, new_n27392_,
    new_n27393_, new_n27394_, new_n27395_, new_n27396_, new_n27397_,
    new_n27398_, new_n27399_, new_n27400_, new_n27401_, new_n27402_,
    new_n27403_, new_n27404_, new_n27405_, new_n27407_, new_n27408_,
    new_n27409_, new_n27410_, new_n27411_, new_n27412_, new_n27413_,
    new_n27414_, new_n27415_, new_n27416_, new_n27417_, new_n27418_,
    new_n27419_, new_n27420_, new_n27421_, new_n27422_, new_n27423_,
    new_n27424_, new_n27425_, new_n27426_, new_n27427_, new_n27428_,
    new_n27429_, new_n27430_, new_n27431_, new_n27432_, new_n27433_,
    new_n27434_, new_n27435_, new_n27436_, new_n27437_, new_n27438_,
    new_n27439_, new_n27440_, new_n27441_, new_n27442_, new_n27443_,
    new_n27444_, new_n27445_, new_n27446_, new_n27447_, new_n27448_,
    new_n27449_, new_n27450_, new_n27451_, new_n27452_, new_n27453_,
    new_n27454_, new_n27455_, new_n27456_, new_n27457_, new_n27458_,
    new_n27459_, new_n27460_, new_n27461_, new_n27462_, new_n27463_,
    new_n27464_, new_n27465_, new_n27466_, new_n27467_, new_n27468_,
    new_n27470_, new_n27471_, new_n27472_, new_n27473_, new_n27474_,
    new_n27475_, new_n27476_, new_n27477_, new_n27478_, new_n27479_,
    new_n27480_, new_n27481_, new_n27482_, new_n27483_, new_n27484_,
    new_n27485_, new_n27486_, new_n27487_, new_n27488_, new_n27489_,
    new_n27490_, new_n27491_, new_n27492_, new_n27493_, new_n27494_,
    new_n27495_, new_n27496_, new_n27497_, new_n27498_, new_n27499_,
    new_n27500_, new_n27501_, new_n27502_, new_n27503_, new_n27504_,
    new_n27505_, new_n27506_, new_n27507_, new_n27508_, new_n27509_,
    new_n27510_, new_n27511_, new_n27512_, new_n27513_, new_n27514_,
    new_n27515_, new_n27516_, new_n27517_, new_n27518_, new_n27519_,
    new_n27520_, new_n27521_, new_n27522_, new_n27523_, new_n27524_,
    new_n27525_, new_n27526_, new_n27527_, new_n27528_, new_n27529_,
    new_n27530_, new_n27531_, new_n27532_, new_n27533_, new_n27534_,
    new_n27535_, new_n27536_, new_n27537_, new_n27538_, new_n27539_,
    new_n27540_, new_n27541_, new_n27542_, new_n27543_, new_n27544_,
    new_n27545_, new_n27546_, new_n27547_, new_n27548_, new_n27549_,
    new_n27550_, new_n27551_, new_n27552_, new_n27553_, new_n27554_,
    new_n27555_, new_n27556_, new_n27557_, new_n27558_, new_n27559_,
    new_n27560_, new_n27561_, new_n27562_, new_n27563_, new_n27564_,
    new_n27565_, new_n27566_, new_n27567_, new_n27568_, new_n27569_,
    new_n27570_, new_n27571_, new_n27573_, new_n27574_, new_n27575_,
    new_n27576_, new_n27577_, new_n27578_, new_n27579_, new_n27580_,
    new_n27581_, new_n27582_, new_n27583_, new_n27584_, new_n27585_,
    new_n27586_, new_n27587_, new_n27588_, new_n27589_, new_n27590_,
    new_n27591_, new_n27592_, new_n27593_, new_n27594_, new_n27595_,
    new_n27596_, new_n27597_, new_n27598_, new_n27599_, new_n27600_,
    new_n27601_, new_n27602_, new_n27603_, new_n27604_, new_n27605_,
    new_n27606_, new_n27607_, new_n27608_, new_n27609_, new_n27610_,
    new_n27611_, new_n27612_, new_n27613_, new_n27614_, new_n27615_,
    new_n27616_, new_n27617_, new_n27618_, new_n27619_, new_n27620_,
    new_n27621_, new_n27622_, new_n27624_, new_n27625_, new_n27626_,
    new_n27627_, new_n27628_, new_n27629_, new_n27630_, new_n27631_,
    new_n27632_, new_n27633_, new_n27634_, new_n27635_, new_n27636_,
    new_n27637_, new_n27638_, new_n27639_, new_n27640_, new_n27641_,
    new_n27642_, new_n27643_, new_n27644_, new_n27645_, new_n27646_,
    new_n27647_, new_n27648_, new_n27649_, new_n27650_, new_n27651_,
    new_n27652_, new_n27653_, new_n27654_, new_n27655_, new_n27656_,
    new_n27657_, new_n27658_, new_n27659_, new_n27660_, new_n27661_,
    new_n27662_, new_n27663_, new_n27664_, new_n27665_, new_n27666_,
    new_n27667_, new_n27668_, new_n27669_, new_n27670_, new_n27671_,
    new_n27672_, new_n27673_, new_n27674_, new_n27675_, new_n27676_,
    new_n27677_, new_n27678_, new_n27679_, new_n27680_, new_n27681_,
    new_n27682_, new_n27683_, new_n27684_, new_n27685_, new_n27686_,
    new_n27687_, new_n27688_, new_n27689_, new_n27690_, new_n27691_,
    new_n27692_, new_n27693_, new_n27694_, new_n27695_, new_n27696_,
    new_n27697_, new_n27698_, new_n27699_, new_n27700_, new_n27701_,
    new_n27702_, new_n27703_, new_n27704_, new_n27705_, new_n27706_,
    new_n27707_, new_n27708_, new_n27709_, new_n27710_, new_n27711_,
    new_n27712_, new_n27713_, new_n27714_, new_n27715_, new_n27716_,
    new_n27717_, new_n27718_, new_n27719_, new_n27720_, new_n27721_,
    new_n27722_, new_n27723_, new_n27724_, new_n27725_, new_n27726_,
    new_n27727_, new_n27728_, new_n27729_, new_n27730_, new_n27731_,
    new_n27732_, new_n27733_, new_n27734_, new_n27735_, new_n27736_,
    new_n27737_, new_n27738_, new_n27739_, new_n27740_, new_n27741_,
    new_n27742_, new_n27743_, new_n27744_, new_n27745_, new_n27746_,
    new_n27747_, new_n27748_, new_n27749_, new_n27750_, new_n27751_,
    new_n27752_, new_n27753_, new_n27754_, new_n27755_, new_n27756_,
    new_n27757_, new_n27758_, new_n27759_, new_n27760_, new_n27761_,
    new_n27762_, new_n27763_, new_n27764_, new_n27765_, new_n27766_,
    new_n27767_, new_n27768_, new_n27769_, new_n27770_, new_n27771_,
    new_n27772_, new_n27773_, new_n27774_, new_n27775_, new_n27776_,
    new_n27777_, new_n27778_, new_n27779_, new_n27780_, new_n27781_,
    new_n27782_, new_n27783_, new_n27784_, new_n27785_, new_n27786_,
    new_n27787_, new_n27788_, new_n27789_, new_n27790_, new_n27791_,
    new_n27792_, new_n27793_, new_n27794_, new_n27795_, new_n27796_,
    new_n27797_, new_n27798_, new_n27799_, new_n27800_, new_n27801_,
    new_n27802_, new_n27803_, new_n27804_, new_n27805_, new_n27806_,
    new_n27807_, new_n27808_, new_n27809_, new_n27810_, new_n27811_,
    new_n27812_, new_n27813_, new_n27814_, new_n27815_, new_n27817_,
    new_n27818_, new_n27819_, new_n27820_, new_n27821_, new_n27822_,
    new_n27823_, new_n27824_, new_n27825_, new_n27826_, new_n27827_,
    new_n27828_, new_n27829_, new_n27830_, new_n27831_, new_n27832_,
    new_n27833_, new_n27835_, new_n27836_, new_n27837_, new_n27838_,
    new_n27839_, new_n27840_, new_n27841_, new_n27842_, new_n27843_,
    new_n27844_, new_n27845_, new_n27846_, new_n27847_, new_n27848_,
    new_n27849_, new_n27850_, new_n27851_, new_n27852_, new_n27853_,
    new_n27854_, new_n27855_, new_n27856_, new_n27857_, new_n27858_,
    new_n27859_, new_n27860_, new_n27861_, new_n27862_, new_n27863_,
    new_n27864_, new_n27865_, new_n27866_, new_n27867_, new_n27868_,
    new_n27869_, new_n27870_, new_n27871_, new_n27872_, new_n27873_,
    new_n27874_, new_n27875_, new_n27876_, new_n27877_, new_n27878_,
    new_n27879_, new_n27880_, new_n27881_, new_n27882_, new_n27883_,
    new_n27884_, new_n27885_, new_n27886_, new_n27887_, new_n27888_,
    new_n27889_, new_n27890_, new_n27891_, new_n27892_, new_n27893_,
    new_n27894_, new_n27895_, new_n27896_, new_n27897_, new_n27898_,
    new_n27899_, new_n27900_, new_n27901_, new_n27902_, new_n27903_,
    new_n27904_, new_n27905_, new_n27906_, new_n27907_, new_n27908_,
    new_n27909_, new_n27910_, new_n27911_, new_n27912_, new_n27913_,
    new_n27914_, new_n27915_, new_n27916_, new_n27917_, new_n27918_,
    new_n27919_, new_n27920_, new_n27921_, new_n27922_, new_n27923_,
    new_n27924_, new_n27925_, new_n27926_, new_n27927_, new_n27928_,
    new_n27929_, new_n27930_, new_n27931_, new_n27932_, new_n27933_,
    new_n27934_, new_n27935_, new_n27936_, new_n27937_, new_n27938_,
    new_n27939_, new_n27940_, new_n27941_, new_n27942_, new_n27943_,
    new_n27944_, new_n27945_, new_n27946_, new_n27947_, new_n27948_,
    new_n27949_, new_n27950_, new_n27951_, new_n27952_, new_n27953_,
    new_n27954_, new_n27955_, new_n27956_, new_n27957_, new_n27958_,
    new_n27959_, new_n27960_, new_n27961_, new_n27962_, new_n27963_,
    new_n27964_, new_n27965_, new_n27966_, new_n27967_, new_n27968_,
    new_n27969_, new_n27970_, new_n27971_, new_n27972_, new_n27973_,
    new_n27974_, new_n27975_, new_n27976_, new_n27977_, new_n27978_,
    new_n27979_, new_n27980_, new_n27981_, new_n27982_, new_n27983_,
    new_n27984_, new_n27985_, new_n27986_, new_n27987_, new_n27988_,
    new_n27989_, new_n27990_, new_n27991_, new_n27992_, new_n27993_,
    new_n27994_, new_n27995_, new_n27996_, new_n27997_, new_n27998_,
    new_n27999_, new_n28000_, new_n28001_, new_n28002_, new_n28003_,
    new_n28004_, new_n28005_, new_n28007_, new_n28008_, new_n28009_,
    new_n28010_, new_n28011_, new_n28012_, new_n28013_, new_n28014_,
    new_n28015_, new_n28016_, new_n28017_, new_n28018_, new_n28019_,
    new_n28020_, new_n28021_, new_n28022_, new_n28023_, new_n28024_,
    new_n28025_, new_n28026_, new_n28027_, new_n28028_, new_n28029_,
    new_n28030_, new_n28031_, new_n28032_, new_n28033_, new_n28034_,
    new_n28036_, new_n28037_, new_n28038_, new_n28039_, new_n28040_,
    new_n28041_, new_n28042_, new_n28043_, new_n28044_, new_n28045_,
    new_n28046_, new_n28047_, new_n28048_, new_n28049_, new_n28050_,
    new_n28051_, new_n28052_, new_n28053_, new_n28054_, new_n28055_,
    new_n28056_, new_n28057_, new_n28058_, new_n28059_, new_n28060_,
    new_n28061_, new_n28062_, new_n28063_, new_n28064_, new_n28065_,
    new_n28066_, new_n28067_, new_n28068_, new_n28069_, new_n28070_,
    new_n28071_, new_n28072_, new_n28073_, new_n28074_, new_n28075_,
    new_n28076_, new_n28077_, new_n28078_, new_n28079_, new_n28081_,
    new_n28082_, new_n28083_, new_n28084_, new_n28085_, new_n28086_,
    new_n28087_, new_n28088_, new_n28089_, new_n28090_, new_n28091_,
    new_n28092_, new_n28093_, new_n28095_, new_n28096_, new_n28097_,
    new_n28098_, new_n28099_, new_n28100_, new_n28101_, new_n28102_,
    new_n28103_, new_n28104_, new_n28105_, new_n28106_, new_n28107_,
    new_n28108_, new_n28109_, new_n28110_, new_n28111_, new_n28112_,
    new_n28113_, new_n28114_, new_n28115_, new_n28116_, new_n28117_,
    new_n28118_, new_n28119_, new_n28120_, new_n28121_, new_n28122_,
    new_n28123_, new_n28124_, new_n28125_, new_n28126_, new_n28127_,
    new_n28128_, new_n28129_, new_n28130_, new_n28131_, new_n28132_,
    new_n28133_, new_n28134_, new_n28135_, new_n28136_, new_n28137_,
    new_n28138_, new_n28139_, new_n28140_, new_n28141_, new_n28142_,
    new_n28143_, new_n28144_, new_n28145_, new_n28146_, new_n28147_,
    new_n28148_, new_n28149_, new_n28150_, new_n28151_, new_n28152_,
    new_n28153_, new_n28154_, new_n28155_, new_n28156_, new_n28157_,
    new_n28158_, new_n28159_, new_n28160_, new_n28161_, new_n28162_,
    new_n28163_, new_n28164_, new_n28165_, new_n28166_, new_n28167_,
    new_n28168_, new_n28169_, new_n28170_, new_n28171_, new_n28172_,
    new_n28173_, new_n28174_, new_n28175_, new_n28176_, new_n28177_,
    new_n28178_, new_n28179_, new_n28180_, new_n28181_, new_n28182_,
    new_n28183_, new_n28184_, new_n28185_, new_n28186_, new_n28187_,
    new_n28188_, new_n28189_, new_n28190_, new_n28191_, new_n28192_,
    new_n28193_, new_n28194_, new_n28195_, new_n28196_, new_n28197_,
    new_n28198_, new_n28199_, new_n28200_, new_n28201_, new_n28202_,
    new_n28203_, new_n28204_, new_n28205_, new_n28206_, new_n28207_,
    new_n28208_, new_n28209_, new_n28210_, new_n28211_, new_n28212_,
    new_n28213_, new_n28214_, new_n28215_, new_n28216_, new_n28217_,
    new_n28218_, new_n28219_, new_n28220_, new_n28221_, new_n28222_,
    new_n28223_, new_n28224_, new_n28225_, new_n28226_, new_n28227_,
    new_n28228_, new_n28229_, new_n28230_, new_n28231_, new_n28232_,
    new_n28233_, new_n28234_, new_n28235_, new_n28236_, new_n28237_,
    new_n28238_, new_n28239_, new_n28240_, new_n28241_, new_n28242_,
    new_n28243_, new_n28244_, new_n28245_, new_n28246_, new_n28247_,
    new_n28248_, new_n28249_, new_n28250_, new_n28251_, new_n28252_,
    new_n28253_, new_n28254_, new_n28255_, new_n28256_, new_n28257_,
    new_n28258_, new_n28259_, new_n28260_, new_n28261_, new_n28262_,
    new_n28263_, new_n28264_, new_n28265_, new_n28266_, new_n28267_,
    new_n28268_, new_n28269_, new_n28270_, new_n28271_, new_n28272_,
    new_n28273_, new_n28274_, new_n28275_, new_n28276_, new_n28277_,
    new_n28278_, new_n28279_, new_n28280_, new_n28281_, new_n28282_,
    new_n28283_, new_n28284_, new_n28285_, new_n28286_, new_n28287_,
    new_n28288_, new_n28289_, new_n28290_, new_n28291_, new_n28292_,
    new_n28293_, new_n28295_, new_n28296_, new_n28297_, new_n28298_,
    new_n28299_, new_n28300_, new_n28301_, new_n28302_, new_n28303_,
    new_n28304_, new_n28305_, new_n28306_, new_n28307_, new_n28308_,
    new_n28309_, new_n28310_, new_n28311_, new_n28312_, new_n28313_,
    new_n28314_, new_n28315_, new_n28316_, new_n28317_, new_n28318_,
    new_n28319_, new_n28320_, new_n28321_, new_n28322_, new_n28323_,
    new_n28324_, new_n28325_, new_n28326_, new_n28327_, new_n28329_,
    new_n28330_, new_n28331_, new_n28332_, new_n28333_, new_n28334_,
    new_n28335_, new_n28336_, new_n28337_, new_n28338_, new_n28339_,
    new_n28340_, new_n28341_, new_n28342_, new_n28343_, new_n28344_,
    new_n28345_, new_n28346_, new_n28347_, new_n28348_, new_n28349_,
    new_n28350_, new_n28351_, new_n28352_, new_n28353_, new_n28354_,
    new_n28355_, new_n28356_, new_n28357_, new_n28358_, new_n28359_,
    new_n28360_, new_n28361_, new_n28362_, new_n28363_, new_n28364_,
    new_n28365_, new_n28366_, new_n28367_, new_n28368_, new_n28369_,
    new_n28370_, new_n28371_, new_n28372_, new_n28373_, new_n28374_,
    new_n28375_, new_n28376_, new_n28377_, new_n28378_, new_n28379_,
    new_n28380_, new_n28381_, new_n28382_, new_n28383_, new_n28384_,
    new_n28385_, new_n28386_, new_n28387_, new_n28388_, new_n28389_,
    new_n28390_, new_n28391_, new_n28392_, new_n28393_, new_n28394_,
    new_n28395_, new_n28396_, new_n28397_, new_n28398_, new_n28399_,
    new_n28400_, new_n28401_, new_n28402_, new_n28403_, new_n28404_,
    new_n28405_, new_n28406_, new_n28407_, new_n28408_, new_n28409_,
    new_n28410_, new_n28411_, new_n28412_, new_n28413_, new_n28414_,
    new_n28415_, new_n28416_, new_n28417_, new_n28418_, new_n28419_,
    new_n28420_, new_n28421_, new_n28422_, new_n28423_, new_n28424_,
    new_n28425_, new_n28426_, new_n28427_, new_n28428_, new_n28429_,
    new_n28430_, new_n28431_, new_n28432_, new_n28433_, new_n28434_,
    new_n28437_, new_n28438_, new_n28441_, new_n28442_, new_n28443_,
    new_n28444_, new_n28445_, new_n28446_, new_n28447_, new_n28448_,
    new_n28449_, new_n28450_, new_n28451_, new_n28452_, new_n28453_,
    new_n28454_, new_n28455_, new_n28456_, new_n28457_, new_n28458_,
    new_n28459_, new_n28460_, new_n28461_, new_n28462_, new_n28463_,
    new_n28464_, new_n28465_, new_n28466_, new_n28467_, new_n28468_,
    new_n28469_, new_n28470_, new_n28471_, new_n28472_, new_n28473_,
    new_n28474_, new_n28475_, new_n28476_, new_n28477_, new_n28478_,
    new_n28479_, new_n28480_, new_n28481_, new_n28482_, new_n28483_,
    new_n28484_, new_n28485_, new_n28486_, new_n28487_, new_n28488_,
    new_n28489_, new_n28490_, new_n28491_, new_n28492_, new_n28493_,
    new_n28494_, new_n28495_, new_n28496_, new_n28497_, new_n28498_,
    new_n28499_, new_n28500_, new_n28501_, new_n28502_, new_n28503_,
    new_n28504_, new_n28505_, new_n28506_, new_n28507_, new_n28508_,
    new_n28509_, new_n28510_, new_n28511_, new_n28512_, new_n28513_,
    new_n28514_, new_n28515_, new_n28516_, new_n28518_, new_n28519_,
    new_n28520_, new_n28521_, new_n28522_, new_n28523_, new_n28524_,
    new_n28525_, new_n28526_, new_n28528_, new_n28529_, new_n28530_,
    new_n28531_, new_n28532_, new_n28533_, new_n28534_, new_n28535_,
    new_n28536_, new_n28537_, new_n28538_, new_n28539_, new_n28540_,
    new_n28541_, new_n28542_, new_n28543_, new_n28544_, new_n28545_,
    new_n28546_, new_n28547_, new_n28548_, new_n28549_, new_n28550_,
    new_n28551_, new_n28552_, new_n28553_, new_n28554_, new_n28555_,
    new_n28556_, new_n28557_, new_n28558_, new_n28559_, new_n28560_,
    new_n28561_, new_n28562_, new_n28563_, new_n28564_, new_n28565_,
    new_n28566_, new_n28567_, new_n28568_, new_n28569_, new_n28570_,
    new_n28571_, new_n28572_, new_n28573_, new_n28575_, new_n28583_,
    new_n28584_, new_n28585_, new_n28589_, new_n28590_, new_n28591_,
    new_n28592_, new_n28593_, new_n28594_, new_n28595_, new_n28596_,
    new_n28597_, new_n28598_, new_n28599_, new_n28600_, new_n28601_,
    new_n28602_, new_n28603_, new_n28604_, new_n28605_, new_n28677_,
    new_n28678_, new_n28680_, new_n28681_, new_n28682_, new_n28683_,
    new_n28684_, new_n28685_, new_n28686_, new_n28687_, new_n28688_,
    new_n28689_, new_n28690_, new_n28691_, new_n28692_, new_n28693_,
    new_n28694_, new_n28695_, new_n28696_, new_n28697_, new_n28698_,
    new_n28699_, new_n28700_, new_n28701_, new_n28702_, new_n28703_,
    new_n28704_, new_n28705_, new_n28706_, new_n28707_, new_n28708_,
    new_n28709_, new_n28710_, new_n28711_, new_n28712_, new_n28713_,
    new_n28714_, new_n28715_, new_n28716_, new_n28717_, new_n28718_,
    new_n28719_, new_n28720_, new_n28721_, new_n28722_, new_n28723_,
    new_n28724_, new_n28725_, new_n28726_, new_n28727_, new_n28728_,
    new_n28729_, new_n28730_, new_n28731_, new_n28732_, new_n28733_,
    new_n28734_, new_n28735_, new_n28736_, new_n28737_, new_n28738_,
    new_n28739_, new_n28740_, new_n28741_, new_n28742_, new_n28743_,
    new_n28744_, new_n28745_, new_n28746_, new_n28747_, new_n28748_,
    new_n28749_, new_n28750_, new_n28751_, new_n28752_, new_n28753_,
    new_n28754_, new_n28755_, new_n28756_, new_n28757_, new_n28758_,
    new_n28759_, new_n28760_, new_n28761_, new_n28762_, new_n28763_,
    new_n28764_, new_n28765_, new_n28766_, new_n28767_, new_n28768_,
    new_n28769_, new_n28770_, new_n28771_, new_n28772_, new_n28773_,
    new_n28774_, new_n28775_, new_n28776_, new_n28777_, new_n28778_,
    new_n28779_, new_n28780_, new_n28781_, new_n28782_, new_n28783_,
    new_n28784_, new_n28785_, new_n28786_, new_n28787_, new_n28788_,
    new_n28789_, new_n28790_, new_n28791_, new_n28792_, new_n28793_,
    new_n28794_, new_n28795_, new_n28796_, new_n28797_, new_n28798_,
    new_n28799_, new_n28800_, new_n28801_, new_n28802_, new_n28803_,
    new_n28804_, new_n28805_, new_n28806_, new_n28807_, new_n28808_,
    new_n28809_, new_n28810_, new_n28811_, new_n28812_, new_n28813_,
    new_n28814_, new_n28815_, new_n28816_, new_n28817_, new_n28818_,
    new_n28819_, new_n28820_, new_n28821_, new_n28822_, new_n28823_,
    new_n28824_, new_n28825_, new_n28826_, new_n28827_, new_n28828_,
    new_n28829_, new_n28830_, new_n28831_, new_n28832_, new_n28833_,
    new_n28834_, new_n28835_, new_n28837_, new_n28838_, new_n28839_,
    new_n28840_, new_n28841_, new_n28842_, new_n28843_, new_n28844_,
    new_n28845_, new_n28846_, new_n28847_, new_n28848_, new_n28849_,
    new_n28850_, new_n28851_, new_n28852_, new_n28853_, new_n28854_,
    new_n28855_, new_n28856_, new_n28857_, new_n28858_, new_n28859_,
    new_n28860_, new_n28861_, new_n28862_, new_n28863_, new_n28864_,
    new_n28865_, new_n28866_, new_n28867_, new_n28868_, new_n28869_,
    new_n28870_, new_n28871_, new_n28872_, new_n28873_, new_n28874_,
    new_n28875_, new_n28876_, new_n28877_, new_n28878_, new_n28879_,
    new_n28880_, new_n28881_, new_n28882_, new_n28883_, new_n28884_,
    new_n28885_, new_n28886_, new_n28887_, new_n28888_, new_n28889_,
    new_n28890_, new_n28891_, new_n28892_, new_n28893_, new_n28894_,
    new_n28895_, new_n28896_, new_n28897_, new_n28898_, new_n28899_,
    new_n28900_, new_n28901_, new_n28902_, new_n28903_, new_n28904_,
    new_n28905_, new_n28906_, new_n28907_, new_n28908_, new_n28909_,
    new_n28910_, new_n28911_, new_n28912_, new_n28913_, new_n28914_,
    new_n28915_, new_n28916_, new_n28917_, new_n28918_, new_n28919_,
    new_n28920_, new_n28921_, new_n28922_, new_n28923_, new_n28924_,
    new_n28925_, new_n28926_, new_n28927_, new_n28928_, new_n28929_,
    new_n28930_, new_n28931_, new_n28932_, new_n28933_, new_n28934_,
    new_n28936_, new_n28937_, new_n28938_, new_n28939_, new_n28940_,
    new_n28941_, new_n28942_, new_n28943_, new_n28944_, new_n28945_,
    new_n28946_, new_n28947_, new_n28948_, new_n28949_, new_n28950_,
    new_n28951_, new_n28952_, new_n28953_, new_n28954_, new_n28955_,
    new_n28956_, new_n28957_, new_n28958_, new_n28959_, new_n28960_,
    new_n28961_, new_n28962_, new_n28963_, new_n28964_, new_n28965_,
    new_n28966_, new_n28967_, new_n28968_, new_n28969_, new_n28970_,
    new_n28971_, new_n28972_, new_n28973_, new_n28974_, new_n28975_,
    new_n28976_, new_n28977_, new_n28978_, new_n28979_, new_n28980_,
    new_n28981_, new_n28982_, new_n28983_, new_n28984_, new_n28985_,
    new_n28986_, new_n28987_, new_n28988_, new_n28989_, new_n28990_,
    new_n28991_, new_n28992_, new_n28993_, new_n28994_, new_n28995_,
    new_n28996_, new_n28997_, new_n28998_, new_n28999_, new_n29000_,
    new_n29001_, new_n29002_, new_n29003_, new_n29004_, new_n29007_,
    new_n29008_, new_n29009_, new_n29010_, new_n29011_, new_n29012_,
    new_n29013_, new_n29015_, new_n29016_, new_n29017_, new_n29018_,
    new_n29019_, new_n29020_, new_n29021_, new_n29022_, new_n29023_,
    new_n29024_, new_n29025_, new_n29026_, new_n29027_, new_n29028_,
    new_n29029_, new_n29030_, new_n29031_, new_n29032_, new_n29033_,
    new_n29034_, new_n29035_, new_n29037_, new_n29038_, new_n29039_,
    new_n29040_, new_n29041_, new_n29042_, new_n29043_, new_n29044_,
    new_n29045_, new_n29046_, new_n29047_, new_n29048_, new_n29049_,
    new_n29050_, new_n29051_, new_n29052_, new_n29053_, new_n29054_,
    new_n29055_, new_n29056_, new_n29057_, new_n29058_, new_n29059_,
    new_n29060_, new_n29061_, new_n29062_, new_n29063_, new_n29064_,
    new_n29065_, new_n29066_, new_n29067_, new_n29068_, new_n29069_,
    new_n29070_, new_n29071_, new_n29072_, new_n29073_, new_n29074_,
    new_n29075_, new_n29076_, new_n29077_, new_n29078_, new_n29079_,
    new_n29080_, new_n29081_, new_n29082_, new_n29083_, new_n29084_,
    new_n29085_, new_n29086_, new_n29087_, new_n29088_, new_n29089_,
    new_n29090_, new_n29091_, new_n29092_, new_n29093_, new_n29094_,
    new_n29095_, new_n29096_, new_n29097_, new_n29098_, new_n29099_,
    new_n29100_, new_n29101_, new_n29102_, new_n29103_, new_n29104_,
    new_n29105_, new_n29106_, new_n29107_, new_n29108_, new_n29109_,
    new_n29110_, new_n29111_, new_n29112_, new_n29113_, new_n29114_,
    new_n29115_, new_n29116_, new_n29117_, new_n29118_, new_n29119_,
    new_n29120_, new_n29121_, new_n29122_, new_n29123_, new_n29124_,
    new_n29125_, new_n29126_, new_n29127_, new_n29128_, new_n29129_,
    new_n29130_, new_n29131_, new_n29132_, new_n29133_, new_n29134_,
    new_n29135_, new_n29136_, new_n29137_, new_n29138_, new_n29139_,
    new_n29140_, new_n29141_, new_n29142_, new_n29143_, new_n29144_,
    new_n29145_, new_n29146_, new_n29147_, new_n29148_, new_n29149_,
    new_n29150_, new_n29151_, new_n29152_, new_n29153_, new_n29154_,
    new_n29155_, new_n29156_, new_n29157_, new_n29158_, new_n29159_,
    new_n29160_, new_n29161_, new_n29162_, new_n29163_, new_n29164_,
    new_n29165_, new_n29166_, new_n29167_, new_n29168_, new_n29169_,
    new_n29170_, new_n29171_, new_n29172_, new_n29173_, new_n29174_,
    new_n29175_, new_n29176_, new_n29177_, new_n29178_, new_n29179_,
    new_n29180_, new_n29181_, new_n29182_, new_n29183_, new_n29184_,
    new_n29185_, new_n29186_, new_n29187_, new_n29188_, new_n29189_,
    new_n29190_, new_n29191_, new_n29192_, new_n29193_, new_n29194_,
    new_n29195_, new_n29196_, new_n29197_, new_n29198_, new_n29199_,
    new_n29200_, new_n29201_, new_n29202_, new_n29203_, new_n29204_,
    new_n29205_, new_n29206_, new_n29207_, new_n29208_, new_n29209_,
    new_n29210_, new_n29211_, new_n29212_, new_n29213_, new_n29214_,
    new_n29215_, new_n29216_, new_n29217_, new_n29218_, new_n29219_,
    new_n29221_, new_n29222_, new_n29223_, new_n29224_, new_n29225_,
    new_n29226_, new_n29227_, new_n29228_, new_n29229_, new_n29230_,
    new_n29231_, new_n29232_, new_n29233_, new_n29234_, new_n29235_,
    new_n29236_, new_n29237_, new_n29238_, new_n29239_, new_n29240_,
    new_n29241_, new_n29242_, new_n29243_, new_n29244_, new_n29245_,
    new_n29246_, new_n29247_, new_n29248_, new_n29249_, new_n29250_,
    new_n29251_, new_n29252_, new_n29253_, new_n29254_, new_n29255_,
    new_n29256_, new_n29257_, new_n29258_, new_n29259_, new_n29260_,
    new_n29261_, new_n29262_, new_n29263_, new_n29264_, new_n29265_,
    new_n29266_, new_n29267_, new_n29268_, new_n29269_, new_n29270_,
    new_n29271_, new_n29272_, new_n29273_, new_n29274_, new_n29275_,
    new_n29276_, new_n29277_, new_n29278_, new_n29279_, new_n29280_,
    new_n29281_, new_n29282_, new_n29283_, new_n29284_, new_n29285_,
    new_n29286_, new_n29287_, new_n29288_, new_n29289_, new_n29290_,
    new_n29291_, new_n29292_, new_n29293_, new_n29294_, new_n29295_,
    new_n29296_, new_n29297_, new_n29308_, new_n29310_, new_n29311_,
    new_n29314_, new_n29322_, new_n29323_, new_n29324_, new_n29325_,
    new_n29326_, new_n29327_, new_n29328_, new_n29329_, new_n29330_,
    new_n29331_, new_n29332_, new_n29333_, new_n29334_, new_n29335_,
    new_n29336_, new_n29337_, new_n29338_, new_n29339_, new_n29340_,
    new_n29341_, new_n29342_, new_n29343_, new_n29344_, new_n29345_,
    new_n29346_, new_n29347_, new_n29348_, new_n29349_, new_n29350_,
    new_n29351_, new_n29352_, new_n29353_, new_n29354_, new_n29355_,
    new_n29356_, new_n29357_, new_n29358_, new_n29359_, new_n29360_,
    new_n29361_, new_n29362_, new_n29363_, new_n29364_, new_n29365_,
    new_n29366_, new_n29367_, new_n29368_, new_n29369_, new_n29370_,
    new_n29371_, new_n29373_, new_n29374_, new_n29375_, new_n29376_,
    new_n29378_, new_n29379_, new_n29380_, new_n29381_, new_n29382_,
    new_n29384_, new_n29385_, new_n29386_, new_n29387_, new_n29388_,
    new_n29390_, new_n29391_, new_n29392_, new_n29393_, new_n29394_,
    new_n29396_, new_n29397_, new_n29398_, new_n29399_, new_n29400_,
    new_n29402_, new_n29403_, new_n29404_, new_n29405_, new_n29406_,
    new_n29408_, new_n29409_, new_n29410_, new_n29411_, new_n29412_,
    new_n29414_, new_n29415_, new_n29416_, new_n29417_, new_n29418_,
    new_n29419_, new_n29420_, new_n29421_, new_n29422_, new_n29423_,
    new_n29424_, new_n29425_, new_n29426_, new_n29427_, new_n29428_,
    new_n29429_, new_n29430_, new_n29431_, new_n29432_, new_n29434_,
    new_n29435_, new_n29436_, new_n29437_, new_n29438_, new_n29439_,
    new_n29440_, new_n29441_, new_n29442_, new_n29443_, new_n29444_,
    new_n29445_, new_n29446_, new_n29447_, new_n29448_, new_n29449_,
    new_n29450_, new_n29451_, new_n29452_, new_n29453_, new_n29454_,
    new_n29455_, new_n29456_, new_n29457_, new_n29458_, new_n29459_,
    new_n29460_, new_n29461_, new_n29462_, new_n29463_, new_n29464_,
    new_n29465_, new_n29466_, new_n29467_, new_n29468_, new_n29469_,
    new_n29470_, new_n29471_, new_n29472_, new_n29473_, new_n29474_,
    new_n29475_, new_n29476_, new_n29477_, new_n29478_, new_n29479_,
    new_n29480_, new_n29481_, new_n29482_, new_n29483_, new_n29484_,
    new_n29485_, new_n29486_, new_n29487_, new_n29488_, new_n29489_,
    new_n29490_, new_n29491_, new_n29492_, new_n29493_, new_n29494_,
    new_n29495_, new_n29496_, new_n29497_, new_n29498_, new_n29499_,
    new_n29500_, new_n29501_, new_n29502_, new_n29503_, new_n29504_,
    new_n29505_, new_n29506_, new_n29507_, new_n29508_, new_n29509_,
    new_n29510_, new_n29511_, new_n29512_, new_n29513_, new_n29514_,
    new_n29515_, new_n29516_, new_n29517_, new_n29518_, new_n29519_,
    new_n29520_, new_n29521_, new_n29522_, new_n29523_, new_n29524_,
    new_n29525_, new_n29526_, new_n29527_, new_n29528_, new_n29529_,
    new_n29530_, new_n29531_, new_n29532_, new_n29533_, new_n29534_,
    new_n29535_, new_n29536_, new_n29537_, new_n29538_, new_n29539_,
    new_n29540_, new_n29541_, new_n29542_, new_n29543_, new_n29544_,
    new_n29545_, new_n29546_, new_n29547_, new_n29548_, new_n29549_,
    new_n29550_, new_n29551_, new_n29552_, new_n29553_, new_n29554_,
    new_n29555_, new_n29556_, new_n29557_, new_n29558_, new_n29559_,
    new_n29560_, new_n29561_, new_n29562_, new_n29563_, new_n29564_,
    new_n29565_, new_n29566_, new_n29567_, new_n29568_, new_n29569_,
    new_n29570_, new_n29571_, new_n29573_, new_n29574_, new_n29575_,
    new_n29576_, new_n29577_, new_n29578_, new_n29579_, new_n29580_,
    new_n29581_, new_n29582_, new_n29583_, new_n29584_, new_n29585_,
    new_n29586_, new_n29587_, new_n29588_, new_n29589_, new_n29590_,
    new_n29591_, new_n29592_, new_n29593_, new_n29594_, new_n29595_,
    new_n29596_, new_n29597_, new_n29598_, new_n29599_, new_n29600_,
    new_n29601_, new_n29602_, new_n29603_, new_n29604_, new_n29605_,
    new_n29607_, new_n29608_, new_n29609_, new_n29610_, new_n29611_,
    new_n29612_, new_n29613_, new_n29614_, new_n29615_, new_n29616_,
    new_n29617_, new_n29618_, new_n29619_, new_n29620_, new_n29621_,
    new_n29622_, new_n29623_, new_n29624_, new_n29625_, new_n29626_,
    new_n29627_, new_n29628_, new_n29629_, new_n29630_, new_n29631_,
    new_n29632_, new_n29634_, new_n29635_, new_n29636_, new_n29637_,
    new_n29638_, new_n29639_, new_n29640_, new_n29641_, new_n29642_,
    new_n29643_, new_n29644_, new_n29645_, new_n29646_, new_n29647_,
    new_n29648_, new_n29649_, new_n29650_, new_n29651_, new_n29652_,
    new_n29653_, new_n29654_, new_n29655_, new_n29656_, new_n29657_,
    new_n29658_, new_n29659_, new_n29660_, new_n29661_, new_n29662_,
    new_n29663_, new_n29664_, new_n29665_, new_n29666_, new_n29667_,
    new_n29669_, new_n29670_, new_n29671_, new_n29672_, new_n29673_,
    new_n29674_, new_n29675_, new_n29676_, new_n29677_, new_n29678_,
    new_n29679_, new_n29680_, new_n29681_, new_n29682_, new_n29683_,
    new_n29684_, new_n29685_, new_n29686_, new_n29687_, new_n29688_,
    new_n29689_, new_n29690_, new_n29691_, new_n29692_, new_n29693_,
    new_n29694_, new_n29695_, new_n29696_, new_n29697_, new_n29698_,
    new_n29699_, new_n29700_, new_n29701_, new_n29702_, new_n29703_,
    new_n29704_, new_n29705_, new_n29706_, new_n29707_, new_n29708_,
    new_n29709_, new_n29710_, new_n29711_, new_n29712_, new_n29713_,
    new_n29714_, new_n29715_, new_n29716_, new_n29717_, new_n29718_,
    new_n29719_, new_n29720_, new_n29721_, new_n29722_, new_n29723_,
    new_n29724_, new_n29725_, new_n29726_, new_n29727_, new_n29728_,
    new_n29729_, new_n29730_, new_n29731_, new_n29732_, new_n29733_,
    new_n29734_, new_n29735_, new_n29736_, new_n29737_, new_n29738_,
    new_n29739_, new_n29740_, new_n29741_, new_n29742_, new_n29743_,
    new_n29744_, new_n29745_, new_n29746_, new_n29747_, new_n29748_,
    new_n29749_, new_n29750_, new_n29751_, new_n29752_, new_n29753_,
    new_n29754_, new_n29755_, new_n29756_, new_n29757_, new_n29758_,
    new_n29759_, new_n29760_, new_n29761_, new_n29762_, new_n29763_,
    new_n29764_, new_n29765_, new_n29766_, new_n29767_, new_n29768_,
    new_n29769_, new_n29770_, new_n29771_, new_n29772_, new_n29773_,
    new_n29774_, new_n29775_, new_n29776_, new_n29777_, new_n29778_,
    new_n29779_, new_n29780_, new_n29781_, new_n29782_, new_n29783_,
    new_n29784_, new_n29785_, new_n29786_, new_n29788_, new_n29789_,
    new_n29790_, new_n29791_, new_n29792_, new_n29793_, new_n29794_,
    new_n29795_, new_n29796_, new_n29797_, new_n29798_, new_n29799_,
    new_n29800_, new_n29801_, new_n29802_, new_n29803_, new_n29804_,
    new_n29805_, new_n29806_, new_n29807_, new_n29808_, new_n29809_,
    new_n29810_, new_n29811_, new_n29812_, new_n29813_, new_n29814_,
    new_n29815_, new_n29816_, new_n29817_, new_n29818_, new_n29819_,
    new_n29820_, new_n29821_, new_n29822_, new_n29823_, new_n29824_,
    new_n29825_, new_n29826_, new_n29827_, new_n29828_, new_n29829_,
    new_n29830_, new_n29831_, new_n29832_, new_n29833_, new_n29834_,
    new_n29835_, new_n29836_, new_n29837_, new_n29838_, new_n29839_,
    new_n29840_, new_n29841_, new_n29842_, new_n29843_, new_n29844_,
    new_n29845_, new_n29846_, new_n29847_, new_n29848_, new_n29849_,
    new_n29850_, new_n29851_, new_n29852_, new_n29853_, new_n29854_,
    new_n29855_, new_n29856_, new_n29857_, new_n29858_, new_n29859_,
    new_n29860_, new_n29861_, new_n29862_, new_n29863_, new_n29864_,
    new_n29865_, new_n29866_, new_n29867_, new_n29868_, new_n29869_,
    new_n29870_, new_n29871_, new_n29872_, new_n29873_, new_n29874_,
    new_n29875_, new_n29876_, new_n29877_, new_n29878_, new_n29879_,
    new_n29880_, new_n29881_, new_n29882_, new_n29883_, new_n29884_,
    new_n29885_, new_n29886_, new_n29887_, new_n29888_, new_n29889_,
    new_n29890_, new_n29891_, new_n29892_, new_n29893_, new_n29894_,
    new_n29895_, new_n29896_, new_n29897_, new_n29898_, new_n29899_,
    new_n29900_, new_n29902_, new_n29903_, new_n29904_, new_n29905_,
    new_n29906_, new_n29907_, new_n29908_, new_n29909_, new_n29910_,
    new_n29911_, new_n29912_, new_n29913_, new_n29914_, new_n29915_,
    new_n29916_, new_n29917_, new_n29918_, new_n29919_, new_n29920_,
    new_n29921_, new_n29922_, new_n29923_, new_n29924_, new_n29925_,
    new_n29926_, new_n29927_, new_n29929_, new_n29930_, new_n29931_,
    new_n29932_, new_n29933_, new_n29934_, new_n29935_, new_n29936_,
    new_n29937_, new_n29938_, new_n29939_, new_n29940_, new_n29941_,
    new_n29942_, new_n29943_, new_n29944_, new_n29945_, new_n29946_,
    new_n29947_, new_n29948_, new_n29949_, new_n29950_, new_n29951_,
    new_n29952_, new_n29954_, new_n29955_, new_n29956_, new_n29957_,
    new_n29958_, new_n29959_, new_n29960_, new_n29961_, new_n29962_,
    new_n29963_, new_n29964_, new_n29965_, new_n29966_, new_n29967_,
    new_n29968_, new_n29969_, new_n29970_, new_n29971_, new_n29972_,
    new_n29973_, new_n29974_, new_n29975_, new_n29977_, new_n29978_,
    new_n29979_, new_n29980_, new_n29981_, new_n29982_, new_n29983_,
    new_n29984_, new_n29985_, new_n29986_, new_n29987_, new_n29988_,
    new_n29989_, new_n29990_, new_n29991_, new_n29992_, new_n29993_,
    new_n29994_, new_n29995_, new_n29996_, new_n29997_, new_n29998_,
    new_n29999_, new_n30000_, new_n30001_, new_n30002_, new_n30003_,
    new_n30004_, new_n30008_, new_n30009_, new_n30010_, new_n30011_,
    new_n30012_, new_n30013_, new_n30014_, new_n30015_, new_n30016_,
    new_n30017_, new_n30018_, new_n30019_, new_n30020_, new_n30021_,
    new_n30022_, new_n30023_, new_n30024_, new_n30025_, new_n30026_,
    new_n30027_, new_n30028_, new_n30029_, new_n30030_, new_n30031_,
    new_n30032_, new_n30033_, new_n30034_, new_n30035_, new_n30036_,
    new_n30037_, new_n30038_, new_n30040_, new_n30041_, new_n30042_,
    new_n30043_, new_n30044_, new_n30045_, new_n30046_, new_n30047_,
    new_n30048_, new_n30049_, new_n30050_, new_n30051_, new_n30052_,
    new_n30053_, new_n30054_, new_n30055_, new_n30056_, new_n30057_,
    new_n30058_, new_n30059_, new_n30060_, new_n30061_, new_n30062_,
    new_n30063_, new_n30064_, new_n30065_, new_n30066_, new_n30067_,
    new_n30068_, new_n30069_, new_n30070_, new_n30071_, new_n30072_,
    new_n30073_, new_n30074_, new_n30075_, new_n30076_, new_n30077_,
    new_n30078_, new_n30079_, new_n30080_, new_n30081_, new_n30083_,
    new_n30084_, new_n30085_, new_n30086_, new_n30087_, new_n30088_,
    new_n30089_, new_n30090_, new_n30091_, new_n30092_, new_n30093_,
    new_n30094_, new_n30095_, new_n30096_, new_n30097_, new_n30098_,
    new_n30099_, new_n30100_, new_n30101_, new_n30102_, new_n30103_,
    new_n30104_, new_n30105_, new_n30106_, new_n30107_, new_n30108_,
    new_n30109_, new_n30110_, new_n30111_, new_n30112_, new_n30113_,
    new_n30115_, new_n30116_, new_n30117_, new_n30118_, new_n30119_,
    new_n30120_, new_n30121_, new_n30122_, new_n30123_, new_n30124_,
    new_n30125_, new_n30126_, new_n30127_, new_n30128_, new_n30129_,
    new_n30130_, new_n30131_, new_n30132_, new_n30133_, new_n30134_,
    new_n30135_, new_n30136_, new_n30137_, new_n30138_, new_n30139_,
    new_n30140_, new_n30141_, new_n30142_, new_n30143_, new_n30144_,
    new_n30145_, new_n30146_, new_n30147_, new_n30148_, new_n30149_,
    new_n30150_, new_n30151_, new_n30152_, new_n30153_, new_n30154_,
    new_n30155_, new_n30156_, new_n30158_, new_n30159_, new_n30160_,
    new_n30161_, new_n30162_, new_n30163_, new_n30164_, new_n30165_,
    new_n30166_, new_n30167_, new_n30168_, new_n30169_, new_n30170_,
    new_n30171_, new_n30172_, new_n30173_, new_n30174_, new_n30175_,
    new_n30176_, new_n30178_, new_n30179_, new_n30180_, new_n30181_,
    new_n30182_, new_n30183_, new_n30184_, new_n30185_, new_n30186_,
    new_n30187_, new_n30188_, new_n30189_, new_n30190_, new_n30191_,
    new_n30192_, new_n30193_, new_n30194_, new_n30195_, new_n30196_,
    new_n30197_, new_n30198_, new_n30199_, new_n30200_, new_n30201_,
    new_n30202_, new_n30203_, new_n30204_, new_n30205_, new_n30206_,
    new_n30207_, new_n30209_, new_n30211_, new_n30212_, new_n30213_,
    new_n30214_, new_n30215_, new_n30216_, new_n30217_, new_n30218_,
    new_n30219_, new_n30220_, new_n30221_, new_n30222_, new_n30223_,
    new_n30224_, new_n30225_, new_n30226_, new_n30227_, new_n30228_,
    new_n30229_, new_n30230_, new_n30231_, new_n30232_, new_n30233_,
    new_n30234_, new_n30235_, new_n30236_, new_n30237_, new_n30238_,
    new_n30239_, new_n30240_, new_n30241_, new_n30242_, new_n30243_,
    new_n30244_, new_n30245_, new_n30246_, new_n30247_, new_n30248_,
    new_n30249_, new_n30252_, new_n30253_, new_n30254_, new_n30255_,
    new_n30256_, new_n30257_, new_n30258_, new_n30259_, new_n30260_,
    new_n30261_, new_n30262_, new_n30263_, new_n30264_, new_n30265_,
    new_n30266_, new_n30267_, new_n30268_, new_n30269_, new_n30270_,
    new_n30271_, new_n30272_, new_n30273_, new_n30274_, new_n30275_,
    new_n30276_, new_n30277_, new_n30278_, new_n30279_, new_n30281_,
    new_n30282_, new_n30283_, new_n30284_, new_n30285_, new_n30286_,
    new_n30287_, new_n30288_, new_n30289_, new_n30290_, new_n30291_,
    new_n30292_, new_n30293_, new_n30294_, new_n30295_, new_n30296_,
    new_n30297_, new_n30298_, new_n30299_, new_n30300_, new_n30301_,
    new_n30302_, new_n30303_, new_n30304_, new_n30307_, new_n30308_,
    new_n30309_, new_n30310_, new_n30311_, new_n30312_, new_n30313_,
    new_n30314_, new_n30315_, new_n30316_, new_n30317_, new_n30318_,
    new_n30319_, new_n30320_, new_n30321_, new_n30322_, new_n30323_,
    new_n30324_, new_n30325_, new_n30326_, new_n30327_, new_n30328_,
    new_n30329_, new_n30330_, new_n30331_, new_n30332_, new_n30333_,
    new_n30334_, new_n30335_, new_n30338_, new_n30339_, new_n30340_,
    new_n30341_, new_n30342_, new_n30343_, new_n30344_, new_n30345_,
    new_n30346_, new_n30347_, new_n30348_, new_n30349_, new_n30350_,
    new_n30351_, new_n30352_, new_n30353_, new_n30355_, new_n30356_,
    new_n30357_, new_n30358_, new_n30359_, new_n30360_, new_n30361_,
    new_n30362_, new_n30363_, new_n30364_, new_n30365_, new_n30368_,
    new_n30369_, new_n30371_, new_n30373_, new_n30374_, new_n30375_,
    new_n30376_, new_n30377_, new_n30378_, new_n30379_, new_n30380_,
    new_n30381_, new_n30382_, new_n30383_, new_n30384_, new_n30385_,
    new_n30387_, new_n30388_, new_n30390_, new_n30391_, new_n30393_,
    new_n30394_, new_n30396_, new_n30397_, new_n30399_, new_n30400_,
    new_n30402_, new_n30403_, new_n30405_, new_n30406_, new_n30408_,
    new_n30409_, new_n30411_, new_n30413_, new_n30414_, new_n30415_,
    new_n30416_, new_n30417_, new_n30419_, new_n30420_, new_n30421_,
    new_n30423_, new_n30424_, new_n30425_, new_n30426_, new_n30427_,
    new_n30429_, new_n30430_, new_n30431_, new_n30432_, new_n30433_,
    new_n30434_, new_n30435_, new_n30436_, new_n30437_, new_n30438_,
    new_n30439_, new_n30440_, new_n30441_, new_n30442_, new_n30443_,
    new_n30444_, new_n30445_, new_n30447_, new_n30449_, new_n30451_,
    new_n30453_, new_n30455_, new_n30457_, new_n30459_, new_n30461_,
    new_n30462_, new_n30463_, new_n30464_, new_n30465_, new_n30466_,
    new_n30467_, new_n30468_, new_n30469_, new_n30470_, new_n30471_,
    new_n30472_, new_n30473_, new_n30474_, new_n30475_, new_n30476_,
    new_n30478_, new_n30479_, new_n30481_, new_n30482_, new_n30484_,
    new_n30485_, new_n30486_, new_n30487_, new_n30490_, new_n30491_,
    new_n30492_, new_n30493_, new_n30494_, new_n30495_, new_n30497_,
    new_n30498_, new_n30499_, new_n30500_, new_n30502_, new_n30503_,
    new_n30505_, new_n30506_, new_n30507_, new_n30509_, new_n30510_,
    new_n30511_, new_n30512_, new_n30514_, new_n30516_, new_n30518_,
    new_n30519_, new_n30521_, new_n30522_, new_n30524_, new_n30526_,
    new_n30527_, new_n30529_, new_n30530_, new_n30532_, new_n30533_,
    new_n30535_, new_n30537_, new_n30539_, new_n30540_, new_n30542_,
    new_n30543_, new_n30544_, new_n30545_, new_n30547_, new_n30548_,
    new_n30549_, new_n30550_, new_n30551_, new_n30557_, new_n30559_,
    new_n30561_, new_n30563_, new_n30565_, new_n30566_, new_n30568_,
    new_n30569_, new_n30571_, new_n30572_, new_n30574_, new_n30576_,
    new_n30577_, new_n30578_, new_n30580_, new_n30582_, new_n30584_,
    new_n30586_, new_n30588_, new_n30590_, new_n30592_, new_n30593_,
    new_n30595_, new_n30596_, new_n30598_, new_n30600_, new_n30601_,
    new_n30603_, new_n30604_, new_n30606_, new_n30607_, new_n30609_,
    new_n30611_, new_n30612_, new_n30614_, new_n30616_, new_n30617_,
    new_n30619_, new_n30620_, new_n30622_, new_n30623_, new_n30625_,
    new_n30626_, new_n30628_, new_n30629_, new_n30631_, new_n30633_,
    new_n30635_, new_n30637_, new_n30638_, new_n30640_, new_n30642_,
    new_n30644_, new_n30645_, new_n30647_, new_n30649_, new_n30651_,
    new_n30653_, new_n30655_, new_n30657_, new_n30659_, new_n30661_,
    new_n30663_, new_n30665_, new_n30667_, new_n30669_, new_n30670_,
    new_n30672_, new_n30673_, new_n30675_, new_n30677_, new_n30679_,
    new_n30681_, new_n30683_, new_n30685_, new_n30687_, new_n30689_,
    new_n30690_, new_n30692_, new_n30694_, new_n30696_, new_n30698_,
    new_n30700_, new_n30702_, new_n30704_, new_n30706_, new_n30708_,
    new_n30710_, new_n30712_, new_n30714_, new_n30716_, new_n30718_,
    new_n30720_, new_n30722_, new_n30724_, new_n30726_, new_n30728_,
    new_n30730_, new_n30732_, new_n30734_, new_n30736_, new_n30738_,
    new_n30740_, new_n30742_, new_n30743_, new_n30745_, new_n30747_,
    new_n30749_, new_n30751_, new_n30753_, new_n30755_, new_n30757_,
    new_n30759_, new_n30761_, new_n30763_, new_n30765_, new_n30767_,
    new_n30769_, new_n30771_, new_n30773_, new_n30775_, new_n30777_,
    new_n30779_, new_n30781_, new_n30783_, new_n30785_, new_n30787_,
    new_n30789_, new_n30791_, new_n30793_, new_n30795_, new_n30797_,
    new_n30799_, new_n30801_, new_n30803_, new_n30805_, new_n30807_,
    new_n30809_, new_n30811_, new_n30813_, new_n30815_, new_n30817_,
    new_n30819_, new_n30821_, new_n30823_, new_n30825_, new_n30827_,
    new_n30829_, new_n30830_, new_n30831_, new_n30832_, new_n30833_,
    new_n30834_, new_n30835_, new_n30836_, new_n30837_, new_n30838_,
    new_n30839_, new_n30840_, new_n30841_, new_n30842_, new_n30843_,
    new_n30844_, new_n30845_, new_n30846_, new_n30847_, new_n30848_,
    new_n30849_, new_n30851_, new_n30853_, new_n30855_, new_n30857_,
    new_n30859_, new_n30861_, new_n30863_, new_n30866_, new_n30867_,
    new_n30868_, new_n30869_, new_n30870_, new_n30871_, new_n30872_,
    new_n30873_, new_n30874_, new_n30875_, new_n30876_, new_n30877_,
    new_n30878_, new_n30879_, new_n30880_, new_n30881_, new_n30883_,
    new_n30884_, new_n30885_, new_n30886_, new_n30887_, new_n30888_,
    new_n30889_, new_n30890_, new_n30891_, new_n30892_, new_n30893_,
    new_n30894_, new_n30895_, new_n30896_, new_n30897_, new_n30898_,
    new_n30899_, new_n30900_, new_n30902_, new_n30903_, new_n30909_,
    new_n30910_, new_n30911_, new_n30912_, new_n30913_, new_n30914_,
    new_n30916_, new_n30917_, new_n30918_, new_n30919_, new_n30920_,
    new_n30921_, new_n30923_, new_n30924_, new_n30925_, new_n30926_,
    new_n30927_, new_n30928_, new_n30930_, new_n30931_, new_n30932_,
    new_n30933_, new_n30934_, new_n30935_, new_n30936_, new_n30938_,
    new_n30941_, new_n30942_, new_n30944_, new_n30945_, new_n30947_,
    new_n30948_, new_n30950_, new_n30951_, new_n30953_, new_n30954_,
    new_n30956_, new_n30957_, new_n30959_, new_n30960_, new_n30962_,
    new_n30964_, new_n30965_, new_n30967_, new_n30968_, new_n30970_,
    new_n30971_, new_n30973_, new_n30974_, new_n30976_, new_n30977_,
    new_n30979_, new_n30981_, new_n30982_, new_n30984_, new_n30985_,
    new_n30987_, new_n30989_, new_n30990_, new_n30992_, new_n30993_,
    new_n30995_, new_n30996_, new_n30998_, new_n30999_, new_n31001_,
    new_n31002_, new_n31004_, new_n31005_, new_n31007_, new_n31008_,
    new_n31010_, new_n31011_, new_n31012_, new_n31013_, new_n31014_,
    new_n31015_, new_n31016_, new_n31017_, new_n31018_, new_n31020_,
    new_n31021_, new_n31023_, new_n31024_, new_n31026_, new_n31027_,
    new_n31029_, new_n31030_, new_n31032_, new_n31033_, new_n31035_,
    new_n31036_, new_n31037_, new_n31038_, new_n31039_, new_n31041_,
    new_n31042_, new_n31044_, new_n31045_, new_n31047_, new_n31048_,
    new_n31050_, new_n31051_, new_n31053_, new_n31054_, new_n31056_,
    new_n31057_, new_n31059_, new_n31060_, new_n31061_, new_n31062_,
    new_n31064_, new_n31066_, new_n31067_, new_n31069_, new_n31070_,
    new_n31072_, new_n31073_, new_n31075_, new_n31076_, new_n31077_,
    new_n31079_, new_n31081_, new_n31082_, new_n31084_, new_n31085_,
    new_n31087_, new_n31088_, new_n31090_, new_n31091_, new_n31093_,
    new_n31094_, new_n31096_, new_n31097_, new_n31099_, new_n31100_,
    new_n31102_, new_n31103_, new_n31105_, new_n31106_, new_n31108_,
    new_n31110_, new_n31111_, new_n31113_, new_n31114_, new_n31116_,
    new_n31117_, new_n31119_, new_n31120_, new_n31122_, new_n31123_,
    new_n31125_, new_n31126_, new_n31128_, new_n31129_, new_n31131_,
    new_n31132_, new_n31134_, new_n31135_, new_n31137_, new_n31138_,
    new_n31139_, new_n31141_, new_n31142_, new_n31144_, new_n31145_,
    new_n31147_, new_n31148_, new_n31150_, new_n31151_, new_n31153_,
    new_n31154_, new_n31156_, new_n31158_, new_n31159_, new_n31161_,
    new_n31162_, new_n31164_, new_n31165_, new_n31167_, new_n31168_,
    new_n31170_, new_n31171_, new_n31173_, new_n31174_, new_n31176_,
    new_n31177_, new_n31178_, new_n31180_, new_n31181_, new_n31183_,
    new_n31184_, new_n31186_, new_n31187_, new_n31189_, new_n31190_,
    new_n31192_, new_n31193_, new_n31195_, new_n31196_, new_n31198_,
    new_n31199_, new_n31201_, new_n31202_, new_n31204_, new_n31205_,
    new_n31207_, new_n31208_, new_n31209_, new_n31210_, new_n31211_,
    new_n31212_, new_n31213_, new_n31214_, new_n31215_, new_n31216_,
    new_n31217_, new_n31218_, new_n31219_, new_n31220_, new_n31221_,
    new_n31222_, new_n31223_, new_n31224_, new_n31225_, new_n31226_,
    new_n31227_, new_n31228_, new_n31229_, new_n31230_, new_n31231_,
    new_n31232_, new_n31233_, new_n31234_, new_n31235_, new_n31236_,
    new_n31237_, new_n31238_, new_n31239_, new_n31240_, new_n31241_,
    new_n31242_, new_n31243_, new_n31244_, new_n31245_, new_n31246_,
    new_n31247_, new_n31248_, new_n31249_, new_n31250_, new_n31251_,
    new_n31252_, new_n31253_, new_n31254_, new_n31255_, new_n31256_,
    new_n31257_, new_n31258_, new_n31259_, new_n31260_, new_n31261_,
    new_n31262_, new_n31263_, new_n31264_, new_n31265_, new_n31266_,
    new_n31267_, new_n31268_, new_n31269_, new_n31270_, new_n31271_,
    new_n31272_, new_n31273_, new_n31274_, new_n31275_, new_n31276_,
    new_n31277_, new_n31278_, new_n31279_, new_n31280_, new_n31281_,
    new_n31282_, new_n31284_, new_n31285_, new_n31287_, new_n31289_,
    new_n31290_, new_n31291_, new_n31293_, new_n31294_, new_n31296_,
    new_n31297_, new_n31299_, new_n31300_, new_n31302_, new_n31303_,
    new_n31305_, new_n31306_, new_n31308_, new_n31309_, new_n31311_,
    new_n31312_, new_n31314_, new_n31315_, new_n31317_, new_n31318_,
    new_n31320_, new_n31321_, new_n31323_, new_n31324_, new_n31326_,
    new_n31327_, new_n31329_, new_n31330_, new_n31332_, new_n31333_,
    new_n31335_, new_n31336_, new_n31338_, new_n31339_, new_n31341_,
    new_n31342_, new_n31343_, new_n31344_, new_n31346_, new_n31347_,
    new_n31348_, new_n31349_, new_n31350_, new_n31351_, new_n31352_,
    new_n31353_, new_n31354_, new_n31355_, new_n31356_, new_n31357_,
    new_n31359_, new_n31361_, new_n31362_, new_n31364_, new_n31365_,
    new_n31367_, new_n31368_, new_n31369_, new_n31370_, new_n31371_,
    new_n31372_, new_n31373_, new_n31374_, new_n31375_, new_n31376_,
    new_n31377_, new_n31378_, new_n31379_, new_n31380_, new_n31381_,
    new_n31382_, new_n31383_, new_n31384_, new_n31385_, new_n31386_,
    new_n31387_, new_n31388_, new_n31389_, new_n31390_, new_n31391_,
    new_n31392_, new_n31393_, new_n31394_, new_n31395_, new_n31396_,
    new_n31397_, new_n31398_, new_n31399_, new_n31400_, new_n31401_,
    new_n31402_, new_n31403_, new_n31404_, new_n31405_, new_n31406_,
    new_n31407_, new_n31408_, new_n31409_, new_n31410_, new_n31411_,
    new_n31412_, new_n31413_, new_n31414_, new_n31415_, new_n31416_,
    new_n31417_, new_n31418_, new_n31419_, new_n31420_, new_n31421_,
    new_n31422_, new_n31423_, new_n31424_, new_n31425_, new_n31426_,
    new_n31427_, new_n31428_, new_n31429_, new_n31430_, new_n31431_,
    new_n31432_, new_n31433_, new_n31434_, new_n31435_, new_n31436_,
    new_n31437_, new_n31438_, new_n31439_, new_n31440_, new_n31441_,
    new_n31442_, new_n31443_, new_n31444_, new_n31445_, new_n31446_,
    new_n31447_, new_n31448_, new_n31449_, new_n31450_, new_n31451_,
    new_n31452_, new_n31453_, new_n31454_, new_n31455_, new_n31456_,
    new_n31457_, new_n31458_, new_n31459_, new_n31460_, new_n31461_,
    new_n31462_, new_n31463_, new_n31464_, new_n31465_, new_n31466_,
    new_n31467_, new_n31468_, new_n31469_, new_n31470_, new_n31471_,
    new_n31472_, new_n31473_, new_n31474_, new_n31475_, new_n31476_,
    new_n31477_, new_n31478_, new_n31479_, new_n31480_, new_n31481_,
    new_n31482_, new_n31483_, new_n31484_, new_n31485_, new_n31486_,
    new_n31487_, new_n31488_, new_n31489_, new_n31490_, new_n31491_,
    new_n31492_, new_n31493_, new_n31494_, new_n31495_, new_n31496_,
    new_n31497_, new_n31498_, new_n31499_, new_n31500_, new_n31501_,
    new_n31502_, new_n31503_, new_n31504_, new_n31505_, new_n31506_,
    new_n31507_, new_n31508_, new_n31509_, new_n31510_, new_n31511_,
    new_n31512_, new_n31513_, new_n31514_, new_n31515_, new_n31516_,
    new_n31517_, new_n31518_, new_n31519_, new_n31520_, new_n31521_,
    new_n31522_, new_n31523_, new_n31524_, new_n31525_, new_n31526_,
    new_n31527_, new_n31528_, new_n31529_, new_n31530_, new_n31531_,
    new_n31532_, new_n31533_, new_n31534_, new_n31535_, new_n31536_,
    new_n31537_, new_n31538_, new_n31539_, new_n31540_, new_n31541_,
    new_n31542_, new_n31543_, new_n31544_, new_n31545_, new_n31546_,
    new_n31547_, new_n31548_, new_n31549_, new_n31550_, new_n31551_,
    new_n31552_, new_n31553_, new_n31554_, new_n31555_, new_n31556_,
    new_n31557_, new_n31558_, new_n31559_, new_n31560_, new_n31561_,
    new_n31562_, new_n31563_, new_n31564_, new_n31565_, new_n31566_,
    new_n31567_, new_n31568_, new_n31569_, new_n31570_, new_n31571_,
    new_n31572_, new_n31573_, new_n31574_, new_n31575_, new_n31576_,
    new_n31577_, new_n31578_, new_n31579_, new_n31580_, new_n31581_,
    new_n31582_, new_n31583_, new_n31584_, new_n31585_, new_n31586_,
    new_n31587_, new_n31588_, new_n31589_, new_n31590_, new_n31591_,
    new_n31592_, new_n31593_, new_n31594_, new_n31595_, new_n31596_,
    new_n31597_, new_n31598_, new_n31599_, new_n31600_, new_n31601_,
    new_n31602_, new_n31603_, new_n31604_, new_n31605_, new_n31606_,
    new_n31607_, new_n31608_, new_n31609_, new_n31610_, new_n31611_,
    new_n31612_, new_n31613_, new_n31614_, new_n31615_, new_n31616_,
    new_n31617_, new_n31618_, new_n31619_, new_n31620_, new_n31621_,
    new_n31622_, new_n31623_, new_n31624_, new_n31625_, new_n31626_,
    new_n31627_, new_n31628_, new_n31629_, new_n31630_, new_n31631_,
    new_n31632_, new_n31633_, new_n31634_, new_n31635_, new_n31636_,
    new_n31637_, new_n31638_, new_n31639_, new_n31640_, new_n31641_,
    new_n31642_, new_n31643_, new_n31644_, new_n31645_, new_n31646_,
    new_n31647_, new_n31648_, new_n31649_, new_n31650_, new_n31651_,
    new_n31652_, new_n31653_, new_n31654_, new_n31655_, new_n31656_,
    new_n31657_, new_n31658_, new_n31659_, new_n31660_, new_n31661_,
    new_n31662_, new_n31663_, new_n31664_, new_n31665_, new_n31666_,
    new_n31667_, new_n31668_, new_n31669_, new_n31670_, new_n31671_,
    new_n31672_, new_n31673_, new_n31674_, new_n31675_, new_n31676_,
    new_n31677_, new_n31678_, new_n31679_, new_n31680_, new_n31681_,
    new_n31682_, new_n31683_, new_n31684_, new_n31685_, new_n31686_,
    new_n31687_, new_n31688_, new_n31689_, new_n31690_, new_n31691_,
    new_n31692_, new_n31693_, new_n31694_, new_n31695_, new_n31696_,
    new_n31697_, new_n31698_, new_n31699_, new_n31700_, new_n31701_,
    new_n31702_, new_n31703_, new_n31704_, new_n31705_, new_n31706_,
    new_n31707_, new_n31708_, new_n31709_, new_n31710_, new_n31711_,
    new_n31712_, new_n31713_, new_n31714_, new_n31715_, new_n31716_,
    new_n31717_, new_n31718_, new_n31719_, new_n31720_, new_n31721_,
    new_n31722_, new_n31723_, new_n31724_, new_n31725_, new_n31726_,
    new_n31727_, new_n31728_, new_n31729_, new_n31730_, new_n31731_,
    new_n31732_, new_n31733_, new_n31734_, new_n31735_, new_n31736_,
    new_n31737_, new_n31738_, new_n31739_, new_n31740_, new_n31741_,
    new_n31742_, new_n31743_, new_n31744_, new_n31745_, new_n31746_,
    new_n31747_, new_n31748_, new_n31749_, new_n31750_, new_n31751_,
    new_n31752_, new_n31753_, new_n31754_, new_n31755_, new_n31756_,
    new_n31757_, new_n31758_, new_n31759_, new_n31760_, new_n31761_,
    new_n31762_, new_n31763_, new_n31764_, new_n31765_, new_n31766_,
    new_n31767_, new_n31768_, new_n31769_, new_n31770_, new_n31771_,
    new_n31772_, new_n31773_, new_n31774_, new_n31775_, new_n31776_,
    new_n31777_, new_n31778_, new_n31779_, new_n31780_, new_n31781_,
    new_n31782_, new_n31783_, new_n31784_, new_n31785_, new_n31786_,
    new_n31787_, new_n31788_, new_n31789_, new_n31790_, new_n31791_,
    new_n31792_, new_n31793_, new_n31794_, new_n31795_, new_n31796_,
    new_n31797_, new_n31798_, new_n31799_, new_n31800_, new_n31801_,
    new_n31802_, new_n31803_, new_n31804_, new_n31805_, new_n31806_,
    new_n31807_, new_n31808_, new_n31809_, new_n31810_, new_n31811_,
    new_n31812_, new_n31813_, new_n31814_, new_n31815_, new_n31816_,
    new_n31817_, new_n31818_, new_n31819_, new_n31820_, new_n31821_,
    new_n31822_, new_n31823_, new_n31824_, new_n31825_, new_n31826_,
    new_n31827_, new_n31828_, new_n31829_, new_n31830_, new_n31831_,
    new_n31832_, new_n31833_, new_n31834_, new_n31835_, new_n31836_,
    new_n31837_, new_n31838_, new_n31839_, new_n31840_, new_n31841_,
    new_n31842_, new_n31843_, new_n31844_, new_n31845_, new_n31846_,
    new_n31847_, new_n31848_, new_n31849_, new_n31850_, new_n31851_,
    new_n31852_, new_n31853_, new_n31854_, new_n31855_, new_n31856_,
    new_n31857_, new_n31858_, new_n31859_, new_n31860_, new_n31861_,
    new_n31862_, new_n31863_, new_n31864_, new_n31865_, new_n31866_,
    new_n31867_, new_n31868_, new_n31869_, new_n31870_, new_n31871_,
    new_n31872_, new_n31873_, new_n31874_, new_n31875_, new_n31876_,
    new_n31877_, new_n31878_, new_n31879_, new_n31880_, new_n31881_,
    new_n31882_, new_n31883_, new_n31884_, new_n31885_, new_n31886_,
    new_n31887_, new_n31888_, new_n31889_, new_n31890_, new_n31891_,
    new_n31892_, new_n31893_, new_n31894_, new_n31895_, new_n31896_,
    new_n31897_, new_n31898_, new_n31899_, new_n31900_, new_n31901_,
    new_n31902_, new_n31903_, new_n31904_, new_n31905_, new_n31906_,
    new_n31907_, new_n31908_, new_n31909_, new_n31910_, new_n31911_,
    new_n31912_, new_n31913_, new_n31914_, new_n31915_, new_n31916_,
    new_n31917_, new_n31918_, new_n31919_, new_n31920_, new_n31921_,
    new_n31922_, new_n31923_, new_n31924_, new_n31925_, new_n31926_,
    new_n31927_, new_n31928_, new_n31929_, new_n31930_, new_n31931_,
    new_n31932_, new_n31933_, new_n31934_, new_n31935_, new_n31936_,
    new_n31937_, new_n31938_, new_n31940_, new_n31941_, new_n31942_,
    new_n31943_, new_n31944_, new_n31945_, new_n31946_, new_n31948_,
    new_n31949_, new_n31950_, new_n31952_, new_n31953_, new_n31954_,
    new_n31955_, new_n31956_, new_n31957_, new_n31959_, new_n31961_,
    new_n31962_, new_n31963_, new_n31964_, new_n31967_, new_n31968_,
    new_n31970_, new_n31971_, new_n31973_, new_n31974_, new_n31975_,
    new_n31976_, new_n31978_, new_n31979_, new_n31980_, new_n31981_,
    new_n31982_, new_n31983_, new_n31984_, new_n31985_, new_n31986_,
    new_n31987_, new_n31988_, new_n31989_, new_n31991_, new_n31992_,
    new_n31993_, new_n31995_, new_n31996_, new_n31998_, new_n31999_,
    new_n32000_, new_n32001_, new_n32003_, new_n32005_, new_n32007_,
    new_n32010_, new_n32011_, new_n32013_, new_n32014_, new_n32016_,
    new_n32018_, new_n32019_, new_n32021_, new_n32022_, new_n32023_,
    new_n32025_, new_n32026_, new_n32027_, new_n32029_, new_n32030_,
    new_n32031_, new_n32033_, new_n32034_, new_n32035_, new_n32036_,
    new_n32038_, new_n32040_, new_n32042_, new_n32043_, new_n32045_,
    new_n32047_, new_n32049_, new_n32051_, new_n32052_, new_n32054_,
    new_n32055_, new_n32056_, new_n32057_, new_n32058_, new_n32059_,
    new_n32060_, new_n32062_, new_n32064_, new_n32066_, new_n32068_,
    new_n32070_, new_n32072_, new_n32073_, new_n32075_, new_n32077_,
    new_n32078_, new_n32079_, new_n32081_, new_n32083_, new_n32085_,
    new_n32086_, new_n32087_, new_n32089_, new_n32090_, new_n32092_,
    new_n32094_, new_n32096_, new_n32098_, new_n32099_, new_n32101_,
    new_n32103_, new_n32105_, new_n32107_, new_n32109_, new_n32110_,
    new_n32112_, new_n32113_, new_n32114_, new_n32116_, new_n32118_,
    new_n32120_, new_n32121_, new_n32122_, new_n32124_, new_n32125_,
    new_n32126_, new_n32128_, new_n32129_, new_n32131_, new_n32132_,
    new_n32134_, new_n32135_, new_n32137_, new_n32138_, new_n32139_,
    new_n32141_, new_n32142_, new_n32143_, new_n32145_, new_n32146_,
    new_n32148_, new_n32149_, new_n32150_, new_n32152_, new_n32153_,
    new_n32155_, new_n32156_, new_n32157_, new_n32158_, new_n32159_,
    new_n32160_, new_n32162_, new_n32164_, new_n32166_, new_n32168_,
    new_n32169_, new_n32170_, new_n32171_, new_n32172_, new_n32173_,
    new_n32174_, new_n32175_, new_n32176_, new_n32177_, new_n32178_,
    new_n32179_, new_n32180_, new_n32181_, new_n32182_, new_n32183_,
    new_n32184_, new_n32185_, new_n32186_, new_n32187_, new_n32188_,
    new_n32189_, new_n32190_, new_n32191_, new_n32192_, new_n32193_,
    new_n32194_, new_n32195_, new_n32196_, new_n32197_, new_n32198_,
    new_n32199_, new_n32200_, new_n32201_, new_n32202_, new_n32203_,
    new_n32204_, new_n32205_, new_n32208_, new_n32209_, new_n32210_,
    new_n32211_, new_n32212_, new_n32213_, new_n32214_, new_n32215_,
    new_n32216_, new_n32217_, new_n32218_, new_n32219_, new_n32220_,
    new_n32221_, new_n32222_, new_n32223_, new_n32224_, new_n32225_,
    new_n32226_, new_n32227_, new_n32228_, new_n32230_, new_n32232_,
    new_n32233_, new_n32235_, new_n32236_, new_n32237_, new_n32238_,
    new_n32239_, new_n32240_, new_n32241_, new_n32242_, new_n32243_,
    new_n32244_, new_n32245_, new_n32246_, new_n32247_, new_n32248_,
    new_n32249_, new_n32252_, new_n32253_, new_n32254_, new_n32255_,
    new_n32256_, new_n32257_, new_n32258_, new_n32259_, new_n32260_,
    new_n32261_, new_n32262_, new_n32263_, new_n32264_, new_n32265_,
    new_n32266_, new_n32267_, new_n32268_, new_n32270_, new_n32271_,
    new_n32272_, new_n32273_, new_n32274_, new_n32275_, new_n32276_,
    new_n32277_, new_n32278_, new_n32279_, new_n32280_, new_n32281_,
    new_n32282_, new_n32283_, new_n32284_, new_n32285_, new_n32286_,
    new_n32287_, new_n32288_, new_n32290_, new_n32291_, new_n32292_,
    new_n32294_, new_n32295_, new_n32296_, new_n32297_, new_n32298_,
    new_n32299_, new_n32300_, new_n32301_, new_n32302_, new_n32303_,
    new_n32304_, new_n32305_, new_n32306_, new_n32307_, new_n32308_,
    new_n32309_, new_n32311_, new_n32312_, new_n32313_, new_n32314_,
    new_n32315_, new_n32316_, new_n32317_, new_n32318_, new_n32319_,
    new_n32320_, new_n32321_, new_n32322_, new_n32323_, new_n32324_,
    new_n32325_, new_n32327_, new_n32328_, new_n32329_, new_n32330_,
    new_n32331_, new_n32332_, new_n32333_, new_n32334_, new_n32335_,
    new_n32336_, new_n32337_, new_n32338_, new_n32339_, new_n32340_,
    new_n32341_, new_n32342_, new_n32343_, new_n32344_, new_n32345_,
    new_n32347_, new_n32348_, new_n32350_, new_n32351_, new_n32352_,
    new_n32353_, new_n32354_, new_n32355_, new_n32356_, new_n32357_,
    new_n32358_, new_n32359_, new_n32360_, new_n32361_, new_n32362_,
    new_n32363_, new_n32364_, new_n32366_, new_n32368_, new_n32369_,
    new_n32370_, new_n32371_, new_n32372_, new_n32373_, new_n32374_,
    new_n32375_, new_n32376_, new_n32377_, new_n32378_, new_n32379_,
    new_n32380_, new_n32381_, new_n32382_, new_n32383_, new_n32384_,
    new_n32386_, new_n32387_, new_n32388_, new_n32389_, new_n32390_,
    new_n32391_, new_n32392_, new_n32393_, new_n32394_, new_n32395_,
    new_n32396_, new_n32397_, new_n32398_, new_n32399_, new_n32400_,
    new_n32401_, new_n32402_, new_n32403_, new_n32404_, new_n32405_,
    new_n32406_, new_n32408_, new_n32409_, new_n32411_, new_n32412_,
    new_n32413_, new_n32414_, new_n32415_, new_n32416_, new_n32417_,
    new_n32418_, new_n32419_, new_n32420_, new_n32421_, new_n32422_,
    new_n32423_, new_n32424_, new_n32425_, new_n32427_, new_n32428_,
    new_n32429_, new_n32430_, new_n32431_, new_n32432_, new_n32433_,
    new_n32434_, new_n32435_, new_n32436_, new_n32437_, new_n32438_,
    new_n32439_, new_n32440_, new_n32441_, new_n32442_, new_n32444_,
    new_n32445_, new_n32446_, new_n32447_, new_n32448_, new_n32449_,
    new_n32450_, new_n32451_, new_n32452_, new_n32453_, new_n32454_,
    new_n32455_, new_n32456_, new_n32457_, new_n32458_, new_n32460_,
    new_n32461_, new_n32462_, new_n32463_, new_n32464_, new_n32465_,
    new_n32466_, new_n32467_, new_n32468_, new_n32469_, new_n32470_,
    new_n32471_, new_n32472_, new_n32473_, new_n32474_, new_n32475_,
    new_n32476_, new_n32477_, new_n32478_, new_n32479_, new_n32481_,
    new_n32483_, new_n32485_, new_n32486_, new_n32487_, new_n32488_,
    new_n32489_, new_n32490_, new_n32491_, new_n32492_, new_n32493_,
    new_n32494_, new_n32495_, new_n32496_, new_n32497_, new_n32498_,
    new_n32499_, new_n32501_, new_n32502_, new_n32504_, new_n32507_,
    new_n32508_, new_n32510_, new_n32512_, new_n32513_, new_n32516_,
    new_n32518_, new_n32520_, new_n32521_, new_n32522_, new_n32523_,
    new_n32524_, new_n32525_, new_n32526_, new_n32527_, new_n32528_,
    new_n32529_, new_n32530_, new_n32531_, new_n32532_, new_n32533_,
    new_n32534_, new_n32535_, new_n32536_, new_n32538_, new_n32539_,
    new_n32540_, new_n32542_, new_n32543_, new_n32544_, new_n32546_,
    new_n32547_, new_n32548_, new_n32550_, new_n32552_, new_n32553_,
    new_n32555_, new_n32556_, new_n32557_, new_n32559_, new_n32561_,
    new_n32563_, new_n32564_, new_n32565_, new_n32567_, new_n32568_,
    new_n32569_, new_n32571_, new_n32573_, new_n32574_, new_n32576_,
    new_n32578_, new_n32581_, new_n32582_, new_n32583_, new_n32584_,
    new_n32585_, new_n32586_, new_n32587_, new_n32588_, new_n32589_,
    new_n32590_, new_n32591_, new_n32592_, new_n32593_, new_n32594_,
    new_n32595_, new_n32596_, new_n32597_, new_n32598_, new_n32599_,
    new_n32600_, new_n32601_, new_n32602_, new_n32603_, new_n32604_,
    new_n32606_, new_n32607_, new_n32608_, new_n32610_, new_n32613_,
    new_n32614_, new_n32615_, new_n32616_, new_n32617_, new_n32618_,
    new_n32619_, new_n32620_, new_n32621_, new_n32622_, new_n32623_,
    new_n32624_, new_n32625_, new_n32626_, new_n32627_, new_n32628_,
    new_n32629_, new_n32630_, new_n32631_, new_n32632_, new_n32636_,
    new_n32638_, new_n32639_, new_n32640_, new_n32641_, new_n32642_,
    new_n32643_, new_n32644_, new_n32645_, new_n32646_, new_n32647_,
    new_n32648_, new_n32649_, new_n32650_, new_n32651_, new_n32652_,
    new_n32653_, new_n32654_, new_n32655_, new_n32657_, new_n32658_,
    new_n32659_, new_n32660_, new_n32661_, new_n32662_, new_n32663_,
    new_n32664_, new_n32665_, new_n32666_, new_n32667_, new_n32668_,
    new_n32669_, new_n32670_, new_n32671_, new_n32672_, new_n32673_,
    new_n32674_, new_n32675_, new_n32677_, new_n32678_, new_n32679_,
    new_n32680_, new_n32681_, new_n32682_, new_n32683_, new_n32684_,
    new_n32685_, new_n32686_, new_n32687_, new_n32688_, new_n32689_,
    new_n32690_, new_n32691_, new_n32692_, new_n32693_, new_n32694_,
    new_n32695_, new_n32697_, new_n32698_, new_n32699_, new_n32700_,
    new_n32701_, new_n32702_, new_n32703_, new_n32704_, new_n32705_,
    new_n32706_, new_n32707_, new_n32708_, new_n32709_, new_n32710_,
    new_n32711_, new_n32712_, new_n32713_, new_n32714_, new_n32717_,
    new_n32718_, new_n32719_, new_n32720_, new_n32721_, new_n32722_,
    new_n32723_, new_n32724_, new_n32725_, new_n32726_, new_n32727_,
    new_n32728_, new_n32729_, new_n32730_, new_n32731_, new_n32732_,
    new_n32733_, new_n32734_, new_n32735_, new_n32736_, new_n32737_,
    new_n32738_, new_n32739_, new_n32740_, new_n32741_, new_n32742_,
    new_n32743_, new_n32744_, new_n32745_, new_n32746_, new_n32747_,
    new_n32748_, new_n32749_, new_n32750_, new_n32751_, new_n32752_,
    new_n32753_, new_n32754_, new_n32755_, new_n32756_, new_n32757_,
    new_n32758_, new_n32759_, new_n32760_, new_n32761_, new_n32762_,
    new_n32763_, new_n32764_, new_n32766_, new_n32767_, new_n32768_,
    new_n32769_, new_n32770_, new_n32771_, new_n32772_, new_n32773_,
    new_n32774_, new_n32775_, new_n32776_, new_n32777_, new_n32778_,
    new_n32779_, new_n32780_, new_n32781_, new_n32782_, new_n32783_,
    new_n32784_, new_n32785_, new_n32786_, new_n32787_, new_n32788_,
    new_n32790_, new_n32791_, new_n32793_, new_n32794_, new_n32796_,
    new_n32797_, new_n32798_, new_n32800_, new_n32802_, new_n32804_,
    new_n32805_, new_n32807_, new_n32809_, new_n32811_, new_n32812_,
    new_n32813_, new_n32814_, new_n32815_, new_n32816_, new_n32817_,
    new_n32818_, new_n32819_, new_n32820_, new_n32821_, new_n32822_,
    new_n32823_, new_n32827_, new_n32828_, new_n32830_, new_n32831_,
    new_n32832_, new_n32833_, new_n32834_, new_n32835_, new_n32836_,
    new_n32837_, new_n32838_, new_n32839_, new_n32840_, new_n32841_,
    new_n32842_, new_n32843_, new_n32844_, new_n32845_, new_n32846_,
    new_n32847_, new_n32848_, new_n32850_, new_n32851_, new_n32852_,
    new_n32854_, new_n32856_, new_n32858_, new_n32859_, new_n32860_,
    new_n32862_, new_n32863_, new_n32864_, new_n32866_, new_n32868_,
    new_n32869_, new_n32870_, new_n32871_, new_n32873_, new_n32875_,
    new_n32877_, new_n32878_, new_n32879_, new_n32881_, new_n32882_,
    new_n32884_, new_n32886_, new_n32887_, new_n32889_, new_n32890_,
    new_n32891_, new_n32892_, new_n32893_, new_n32894_, new_n32895_,
    new_n32896_, new_n32897_, new_n32898_, new_n32900_, new_n32901_,
    new_n32902_, new_n32904_, new_n32905_, new_n32907_, new_n32908_,
    new_n32910_, new_n32912_, new_n32914_, new_n32916_, new_n32918_,
    new_n32920_, new_n32922_, new_n32924_, new_n32925_, new_n32926_,
    new_n32928_, new_n32929_, new_n32931_, new_n32933_, new_n32935_,
    new_n32936_, new_n32938_, new_n32939_, new_n32940_, new_n32942_,
    new_n32943_, new_n32944_, new_n32948_, new_n32949_, new_n32950_,
    new_n32952_, new_n32954_, new_n32956_, new_n32957_, new_n32958_,
    new_n32959_, new_n32960_, new_n32961_, new_n32962_, new_n32963_,
    new_n32964_, new_n32965_, new_n32966_, new_n32967_, new_n32969_,
    new_n32971_, new_n32972_, new_n32973_, new_n32974_, new_n32975_,
    new_n32976_, new_n32977_, new_n32978_, new_n32979_, new_n32980_,
    new_n32981_, new_n32982_, new_n32983_, new_n32985_, new_n32987_,
    new_n32988_, new_n32989_, new_n32991_, new_n32992_, new_n32993_,
    new_n32994_, new_n32996_, new_n32998_, new_n32999_, new_n33000_,
    new_n33001_, new_n33002_, new_n33003_, new_n33004_, new_n33005_,
    new_n33006_, new_n33008_, new_n33010_, new_n33012_, new_n33013_,
    new_n33014_, new_n33015_, new_n33019_, new_n33022_, new_n33023_,
    new_n33025_, new_n33026_, new_n33028_, new_n33030_, new_n33032_,
    new_n33034_, new_n33036_, new_n33038_, new_n33040_, new_n33041_,
    new_n33043_, new_n33046_, new_n33047_, new_n33048_, new_n33050_,
    new_n33052_, new_n33053_, new_n33054_, new_n33056_, new_n33058_,
    new_n33060_, new_n33061_, new_n33063_, new_n33066_, new_n33068_,
    new_n33070_, new_n33071_, new_n33072_, new_n33073_, new_n33075_,
    new_n33077_, new_n33078_, new_n33080_, new_n33082_, new_n33084_,
    new_n33085_, new_n33087_, new_n33089_, new_n33091_, new_n33093_,
    new_n33095_, new_n33099_, new_n33100_, new_n33102_, new_n33105_,
    new_n33106_, new_n33109_, new_n33110_, new_n33111_, new_n33112_,
    new_n33113_, new_n33114_, new_n33115_, new_n33116_, new_n33117_,
    new_n33118_, new_n33119_, new_n33120_, new_n33121_, new_n33122_,
    new_n33123_, new_n33124_, new_n33125_, new_n33126_, new_n33127_,
    new_n33130_, new_n33131_, new_n33132_, new_n33133_, new_n33134_,
    new_n33135_, new_n33136_, new_n33137_, new_n33138_, new_n33139_,
    new_n33140_, new_n33141_, new_n33142_, new_n33143_, new_n33144_,
    new_n33145_, new_n33148_, new_n33149_, new_n33150_, new_n33151_,
    new_n33152_, new_n33153_, new_n33154_, new_n33155_, new_n33156_,
    new_n33157_, new_n33158_, new_n33159_, new_n33160_, new_n33161_,
    new_n33162_, new_n33163_, new_n33164_, new_n33167_, new_n33168_,
    new_n33169_, new_n33170_, new_n33171_, new_n33172_, new_n33173_,
    new_n33174_, new_n33175_, new_n33176_, new_n33177_, new_n33178_,
    new_n33179_, new_n33180_, new_n33181_, new_n33182_, new_n33186_,
    new_n33191_, new_n33193_, new_n33195_, new_n33197_, new_n33200_,
    new_n33202_, new_n33204_, new_n33206_, new_n33208_, new_n33210_,
    new_n33212_, new_n33214_, new_n33216_, new_n33218_, new_n33220_,
    new_n33222_, new_n33224_, new_n33226_, new_n33228_, new_n33230_,
    new_n33232_, new_n33234_, new_n33236_, new_n33238_, new_n33239_,
    new_n33240_, new_n33242_, new_n33244_, new_n33246_, new_n33248_,
    new_n33250_, new_n33252_, new_n33254_, new_n33256_, new_n33257_,
    new_n33258_, new_n33260_, new_n33262_, new_n33264_, new_n33266_,
    new_n33268_, new_n33270_, new_n33271_, new_n33272_, new_n33273_,
    new_n33275_, new_n33277_, new_n33278_, new_n33279_, new_n33281_,
    new_n33282_, new_n33283_, new_n33285_, new_n33286_, new_n33287_,
    new_n33289_, new_n33291_, new_n33294_, new_n33297_, new_n33300_,
    new_n33303_, new_n33306_, new_n33309_, new_n33312_, new_n33315_,
    new_n33318_, new_n33321_, new_n33324_, new_n33327_, new_n33330_,
    new_n33333_, new_n33336_, new_n33339_, new_n33342_, new_n33345_,
    new_n33348_, new_n33351_, new_n33354_, new_n33356_, new_n33357_,
    new_n33358_, new_n33359_, new_n33360_, new_n33361_, new_n33362_,
    new_n33363_, new_n33364_, new_n33367_, new_n33370_, new_n33373_,
    new_n33376_, new_n33379_, new_n33382_, new_n33384_, new_n33387_,
    new_n33390_, new_n33393_, new_n33396_, new_n33399_, new_n33401_,
    new_n33403_, new_n33405_, new_n33407_, new_n33410_, new_n33412_,
    new_n33414_, new_n33416_, new_n33418_, new_n33420_, new_n33422_,
    new_n33424_, new_n33426_, new_n33428_, new_n33430_, new_n33432_,
    new_n33434_, new_n33436_, new_n33438_, new_n33440_, new_n33442_,
    new_n33444_, new_n33446_, new_n33448_, new_n33451_, new_n33454_;
  INV_X1     g00000(.I(pi0137), .ZN(new_n2436_));
  INV_X1     g00001(.I(pi0095), .ZN(new_n2437_));
  NOR2_X1    g00002(.A1(new_n2437_), .A2(pi0479), .ZN(new_n2438_));
  AOI21_X1   g00003(.A1(new_n2438_), .A2(pi0234), .B(pi0332), .ZN(new_n2439_));
  INV_X1     g00004(.I(pi0234), .ZN(new_n2440_));
  INV_X1     g00005(.I(pi0081), .ZN(new_n2441_));
  NOR4_X1    g00006(.A1(pi0061), .A2(pi0076), .A3(pi0085), .A4(pi0106), .ZN(new_n2442_));
  OR3_X2     g00007(.A1(pi0048), .A2(pi0049), .A3(pi0089), .Z(new_n2443_));
  NOR3_X1    g00008(.A1(pi0082), .A2(pi0084), .A3(pi0111), .ZN(new_n2444_));
  NOR2_X1    g00009(.A1(pi0036), .A2(pi0068), .ZN(new_n2445_));
  NOR2_X1    g00010(.A1(pi0045), .A2(pi0104), .ZN(new_n2446_));
  NAND3_X1   g00011(.A1(new_n2444_), .A2(new_n2445_), .A3(new_n2446_), .ZN(new_n2447_));
  NOR3_X1    g00012(.A1(new_n2447_), .A2(new_n2442_), .A3(new_n2443_), .ZN(new_n2448_));
  NOR2_X1    g00013(.A1(pi0083), .A2(pi0103), .ZN(new_n2449_));
  NOR2_X1    g00014(.A1(pi0066), .A2(pi0073), .ZN(new_n2450_));
  NOR2_X1    g00015(.A1(pi0067), .A2(pi0069), .ZN(new_n2451_));
  NAND3_X1   g00016(.A1(new_n2449_), .A2(new_n2450_), .A3(new_n2451_), .ZN(new_n2452_));
  INV_X1     g00017(.I(new_n2452_), .ZN(new_n2453_));
  INV_X1     g00018(.I(pi0064), .ZN(new_n2454_));
  NOR2_X1    g00019(.A1(pi0063), .A2(pi0107), .ZN(new_n2455_));
  NOR2_X1    g00020(.A1(pi0065), .A2(pi0071), .ZN(new_n2456_));
  NAND3_X1   g00021(.A1(new_n2455_), .A2(new_n2456_), .A3(new_n2454_), .ZN(new_n2457_));
  INV_X1     g00022(.I(new_n2457_), .ZN(new_n2458_));
  NAND4_X1   g00023(.A1(new_n2448_), .A2(new_n2441_), .A3(new_n2453_), .A4(new_n2458_), .ZN(new_n2459_));
  INV_X1     g00024(.I(pi0050), .ZN(new_n2460_));
  INV_X1     g00025(.I(pi0077), .ZN(new_n2461_));
  INV_X1     g00026(.I(pi0102), .ZN(new_n2462_));
  NOR2_X1    g00027(.A1(pi0088), .A2(pi0098), .ZN(new_n2463_));
  NAND4_X1   g00028(.A1(new_n2463_), .A2(new_n2460_), .A3(new_n2461_), .A4(new_n2462_), .ZN(new_n2464_));
  INV_X1     g00029(.I(pi0046), .ZN(new_n2465_));
  INV_X1     g00030(.I(pi0094), .ZN(new_n2466_));
  NOR3_X1    g00031(.A1(pi0053), .A2(pi0060), .A3(pi0086), .ZN(new_n2467_));
  NOR2_X1    g00032(.A1(pi0097), .A2(pi0108), .ZN(new_n2468_));
  NAND4_X1   g00033(.A1(new_n2467_), .A2(new_n2465_), .A3(new_n2468_), .A4(new_n2466_), .ZN(new_n2469_));
  INV_X1     g00034(.I(pi0109), .ZN(new_n2470_));
  INV_X1     g00035(.I(pi0110), .ZN(new_n2471_));
  NAND2_X1   g00036(.A1(new_n2470_), .A2(new_n2471_), .ZN(new_n2472_));
  NOR2_X1    g00037(.A1(pi0047), .A2(pi0091), .ZN(new_n2473_));
  INV_X1     g00038(.I(new_n2473_), .ZN(new_n2474_));
  NOR4_X1    g00039(.A1(new_n2469_), .A2(new_n2464_), .A3(new_n2472_), .A4(new_n2474_), .ZN(new_n2475_));
  INV_X1     g00040(.I(new_n2475_), .ZN(new_n2476_));
  NOR2_X1    g00041(.A1(pi0035), .A2(pi0093), .ZN(new_n2477_));
  INV_X1     g00042(.I(new_n2477_), .ZN(new_n2478_));
  NOR2_X1    g00043(.A1(pi0058), .A2(pi0090), .ZN(new_n2479_));
  INV_X1     g00044(.I(new_n2479_), .ZN(new_n2480_));
  NOR3_X1    g00045(.A1(new_n2478_), .A2(new_n2480_), .A3(pi0070), .ZN(new_n2481_));
  INV_X1     g00046(.I(new_n2481_), .ZN(new_n2482_));
  NOR2_X1    g00047(.A1(pi0040), .A2(pi0072), .ZN(new_n2483_));
  NOR2_X1    g00048(.A1(pi0032), .A2(pi0095), .ZN(new_n2484_));
  NAND2_X1   g00049(.A1(new_n2483_), .A2(new_n2484_), .ZN(new_n2485_));
  NOR2_X1    g00050(.A1(pi0051), .A2(pi0096), .ZN(new_n2486_));
  INV_X1     g00051(.I(new_n2486_), .ZN(new_n2487_));
  NOR2_X1    g00052(.A1(new_n2485_), .A2(new_n2487_), .ZN(new_n2488_));
  INV_X1     g00053(.I(new_n2488_), .ZN(new_n2489_));
  NOR4_X1    g00054(.A1(new_n2459_), .A2(new_n2476_), .A3(new_n2482_), .A4(new_n2489_), .ZN(new_n2490_));
  INV_X1     g00055(.I(new_n2490_), .ZN(new_n2491_));
  INV_X1     g00056(.I(pi0061), .ZN(new_n2492_));
  INV_X1     g00057(.I(pi0076), .ZN(new_n2493_));
  NAND2_X1   g00058(.A1(new_n2492_), .A2(new_n2493_), .ZN(new_n2494_));
  INV_X1     g00059(.I(pi0085), .ZN(new_n2495_));
  INV_X1     g00060(.I(pi0106), .ZN(new_n2496_));
  NAND2_X1   g00061(.A1(new_n2495_), .A2(new_n2496_), .ZN(new_n2497_));
  NOR3_X1    g00062(.A1(pi0048), .A2(pi0049), .A3(pi0089), .ZN(new_n2498_));
  OAI21_X1   g00063(.A1(new_n2494_), .A2(new_n2497_), .B(new_n2498_), .ZN(new_n2499_));
  NOR4_X1    g00064(.A1(new_n2499_), .A2(new_n2447_), .A3(new_n2452_), .A4(new_n2457_), .ZN(new_n2500_));
  NAND3_X1   g00065(.A1(new_n2500_), .A2(new_n2441_), .A3(new_n2475_), .ZN(new_n2501_));
  NOR2_X1    g00066(.A1(pi0072), .A2(pi0096), .ZN(new_n2502_));
  INV_X1     g00067(.I(new_n2502_), .ZN(new_n2503_));
  NOR2_X1    g00068(.A1(pi0051), .A2(pi0070), .ZN(new_n2504_));
  INV_X1     g00069(.I(new_n2504_), .ZN(new_n2505_));
  NOR2_X1    g00070(.A1(new_n2503_), .A2(new_n2505_), .ZN(new_n2506_));
  INV_X1     g00071(.I(new_n2506_), .ZN(new_n2507_));
  NOR2_X1    g00072(.A1(new_n2478_), .A2(new_n2480_), .ZN(new_n2508_));
  INV_X1     g00073(.I(new_n2508_), .ZN(new_n2509_));
  NOR3_X1    g00074(.A1(new_n2501_), .A2(new_n2507_), .A3(new_n2509_), .ZN(new_n2510_));
  INV_X1     g00075(.I(new_n2510_), .ZN(new_n2511_));
  NOR2_X1    g00076(.A1(pi0032), .A2(pi0040), .ZN(new_n2512_));
  INV_X1     g00077(.I(new_n2512_), .ZN(new_n2513_));
  NOR2_X1    g00078(.A1(new_n2513_), .A2(pi0095), .ZN(new_n2514_));
  INV_X1     g00079(.I(new_n2514_), .ZN(new_n2515_));
  NOR2_X1    g00080(.A1(new_n2511_), .A2(new_n2515_), .ZN(new_n2516_));
  NOR2_X1    g00081(.A1(new_n2516_), .A2(new_n2438_), .ZN(new_n2517_));
  MUX2_X1    g00082(.I0(new_n2517_), .I1(new_n2491_), .S(new_n2440_), .Z(new_n2518_));
  INV_X1     g00083(.I(new_n2518_), .ZN(new_n2519_));
  OAI21_X1   g00084(.A1(new_n2519_), .A2(new_n2436_), .B(new_n2439_), .ZN(new_n2520_));
  INV_X1     g00085(.I(new_n2520_), .ZN(new_n2521_));
  INV_X1     g00086(.I(pi0105), .ZN(new_n2522_));
  INV_X1     g00087(.I(pi0228), .ZN(new_n2523_));
  NOR2_X1    g00088(.A1(new_n2522_), .A2(new_n2523_), .ZN(new_n2524_));
  INV_X1     g00089(.I(new_n2524_), .ZN(new_n2525_));
  INV_X1     g00090(.I(pi0153), .ZN(new_n2526_));
  NOR2_X1    g00091(.A1(new_n2526_), .A2(pi0332), .ZN(new_n2527_));
  AOI21_X1   g00092(.A1(new_n2525_), .A2(new_n2527_), .B(pi0216), .ZN(new_n2528_));
  INV_X1     g00093(.I(new_n2528_), .ZN(new_n2529_));
  NOR2_X1    g00094(.A1(pi0215), .A2(pi0221), .ZN(new_n2530_));
  INV_X1     g00095(.I(new_n2530_), .ZN(new_n2531_));
  NOR3_X1    g00096(.A1(new_n2521_), .A2(new_n2529_), .A3(new_n2531_), .ZN(new_n2532_));
  NOR2_X1    g00097(.A1(pi0056), .A2(pi0062), .ZN(new_n2533_));
  NOR2_X1    g00098(.A1(pi0075), .A2(pi0087), .ZN(new_n2534_));
  INV_X1     g00099(.I(new_n2534_), .ZN(new_n2535_));
  NOR2_X1    g00100(.A1(new_n2535_), .A2(pi0092), .ZN(new_n2536_));
  INV_X1     g00101(.I(new_n2536_), .ZN(new_n2537_));
  NOR2_X1    g00102(.A1(pi0054), .A2(pi0074), .ZN(new_n2538_));
  INV_X1     g00103(.I(new_n2538_), .ZN(new_n2539_));
  NOR2_X1    g00104(.A1(new_n2537_), .A2(new_n2539_), .ZN(new_n2540_));
  INV_X1     g00105(.I(new_n2540_), .ZN(new_n2541_));
  NOR2_X1    g00106(.A1(new_n2541_), .A2(pi0055), .ZN(new_n2542_));
  INV_X1     g00107(.I(new_n2542_), .ZN(new_n2543_));
  NOR2_X1    g00108(.A1(pi0038), .A2(pi0039), .ZN(new_n2544_));
  INV_X1     g00109(.I(new_n2544_), .ZN(new_n2545_));
  NOR2_X1    g00110(.A1(new_n2545_), .A2(pi0100), .ZN(new_n2546_));
  INV_X1     g00111(.I(new_n2546_), .ZN(new_n2547_));
  NOR2_X1    g00112(.A1(new_n2543_), .A2(new_n2547_), .ZN(new_n2548_));
  AND3_X2    g00113(.A1(new_n2532_), .A2(new_n2533_), .A3(new_n2548_), .Z(new_n2549_));
  INV_X1     g00114(.I(pi0221), .ZN(new_n2550_));
  INV_X1     g00115(.I(pi0929), .ZN(new_n2551_));
  INV_X1     g00116(.I(pi1144), .ZN(new_n2552_));
  INV_X1     g00117(.I(pi0833), .ZN(new_n2553_));
  NOR2_X1    g00118(.A1(new_n2553_), .A2(pi0216), .ZN(new_n2554_));
  INV_X1     g00119(.I(new_n2554_), .ZN(new_n2555_));
  AOI21_X1   g00120(.A1(new_n2555_), .A2(new_n2552_), .B(new_n2551_), .ZN(new_n2556_));
  NOR3_X1    g00121(.A1(new_n2554_), .A2(pi0929), .A3(new_n2552_), .ZN(new_n2557_));
  NOR3_X1    g00122(.A1(new_n2556_), .A2(pi0332), .A3(new_n2557_), .ZN(new_n2558_));
  NOR2_X1    g00123(.A1(new_n2558_), .A2(new_n2550_), .ZN(new_n2559_));
  INV_X1     g00124(.I(new_n2559_), .ZN(new_n2560_));
  AOI21_X1   g00125(.A1(new_n2439_), .A2(new_n2524_), .B(new_n2529_), .ZN(new_n2561_));
  INV_X1     g00126(.I(pi0216), .ZN(new_n2562_));
  INV_X1     g00127(.I(pi0332), .ZN(new_n2563_));
  AOI21_X1   g00128(.A1(pi0265), .A2(new_n2563_), .B(new_n2562_), .ZN(new_n2564_));
  NOR4_X1    g00129(.A1(new_n2560_), .A2(new_n2531_), .A3(new_n2561_), .A4(new_n2564_), .ZN(new_n2565_));
  INV_X1     g00130(.I(pi0215), .ZN(new_n2566_));
  NOR2_X1    g00131(.A1(pi0332), .A2(pi1144), .ZN(new_n2567_));
  INV_X1     g00132(.I(new_n2567_), .ZN(new_n2568_));
  NOR2_X1    g00133(.A1(new_n2568_), .A2(new_n2566_), .ZN(new_n2569_));
  NOR2_X1    g00134(.A1(new_n2565_), .A2(new_n2569_), .ZN(new_n2570_));
  NOR2_X1    g00135(.A1(pi0057), .A2(pi0059), .ZN(new_n2571_));
  NAND3_X1   g00136(.A1(new_n2549_), .A2(new_n2570_), .A3(new_n2571_), .ZN(new_n2572_));
  INV_X1     g00137(.I(new_n2564_), .ZN(new_n2573_));
  NOR2_X1    g00138(.A1(pi0152), .A2(pi0161), .ZN(new_n2574_));
  INV_X1     g00139(.I(new_n2574_), .ZN(new_n2575_));
  NOR2_X1    g00140(.A1(new_n2575_), .A2(pi0166), .ZN(new_n2576_));
  NOR2_X1    g00141(.A1(new_n2576_), .A2(pi0146), .ZN(new_n2577_));
  NOR2_X1    g00142(.A1(new_n2577_), .A2(pi0210), .ZN(new_n2578_));
  INV_X1     g00143(.I(new_n2578_), .ZN(new_n2579_));
  AOI21_X1   g00144(.A1(pi0095), .A2(pi0234), .B(pi0137), .ZN(new_n2580_));
  AOI21_X1   g00145(.A1(new_n2579_), .A2(new_n2580_), .B(pi0332), .ZN(new_n2581_));
  NAND2_X1   g00146(.A1(new_n2518_), .A2(new_n2581_), .ZN(new_n2582_));
  NOR2_X1    g00147(.A1(new_n2522_), .A2(pi0228), .ZN(new_n2583_));
  AND2_X2    g00148(.A1(new_n2582_), .A2(new_n2583_), .Z(new_n2584_));
  OAI21_X1   g00149(.A1(new_n2584_), .A2(new_n2529_), .B(new_n2573_), .ZN(new_n2585_));
  NAND2_X1   g00150(.A1(new_n2585_), .A2(new_n2550_), .ZN(new_n2586_));
  INV_X1     g00151(.I(pi0299), .ZN(new_n2587_));
  INV_X1     g00152(.I(pi0222), .ZN(new_n2588_));
  NOR2_X1    g00153(.A1(new_n2553_), .A2(pi0224), .ZN(new_n2589_));
  NOR2_X1    g00154(.A1(new_n2589_), .A2(new_n2588_), .ZN(new_n2590_));
  NOR2_X1    g00155(.A1(new_n2590_), .A2(pi0223), .ZN(new_n2591_));
  INV_X1     g00156(.I(new_n2591_), .ZN(new_n2592_));
  INV_X1     g00157(.I(new_n2589_), .ZN(new_n2593_));
  OAI21_X1   g00158(.A1(pi0332), .A2(pi0929), .B(new_n2593_), .ZN(new_n2594_));
  INV_X1     g00159(.I(pi0224), .ZN(new_n2595_));
  NAND3_X1   g00160(.A1(new_n2595_), .A2(new_n2563_), .A3(pi0265), .ZN(new_n2596_));
  NOR2_X1    g00161(.A1(pi0222), .A2(pi0223), .ZN(new_n2597_));
  INV_X1     g00162(.I(new_n2597_), .ZN(new_n2598_));
  NOR2_X1    g00163(.A1(new_n2568_), .A2(new_n2598_), .ZN(new_n2599_));
  NAND4_X1   g00164(.A1(new_n2592_), .A2(new_n2594_), .A3(new_n2596_), .A4(new_n2599_), .ZN(new_n2600_));
  INV_X1     g00165(.I(pi0198), .ZN(new_n2601_));
  AOI21_X1   g00166(.A1(new_n2601_), .A2(pi0142), .B(pi0137), .ZN(new_n2602_));
  NOR3_X1    g00167(.A1(new_n2519_), .A2(new_n2439_), .A3(new_n2602_), .ZN(new_n2603_));
  INV_X1     g00168(.I(pi0223), .ZN(new_n2604_));
  NOR3_X1    g00169(.A1(pi0144), .A2(pi0174), .A3(pi0189), .ZN(new_n2605_));
  INV_X1     g00170(.I(new_n2605_), .ZN(new_n2606_));
  INV_X1     g00171(.I(new_n2517_), .ZN(new_n2607_));
  NOR2_X1    g00172(.A1(new_n2440_), .A2(pi0332), .ZN(new_n2608_));
  NOR2_X1    g00173(.A1(pi0095), .A2(pi0137), .ZN(new_n2609_));
  AOI21_X1   g00174(.A1(pi0198), .A2(new_n2609_), .B(new_n2608_), .ZN(new_n2610_));
  NOR2_X1    g00175(.A1(pi0234), .A2(pi0332), .ZN(new_n2611_));
  NOR4_X1    g00176(.A1(new_n2490_), .A2(pi0137), .A3(new_n2601_), .A4(new_n2611_), .ZN(new_n2612_));
  AOI21_X1   g00177(.A1(new_n2607_), .A2(new_n2610_), .B(new_n2612_), .ZN(new_n2613_));
  NOR2_X1    g00178(.A1(pi0222), .A2(pi0224), .ZN(new_n2614_));
  NAND4_X1   g00179(.A1(new_n2613_), .A2(new_n2604_), .A3(new_n2606_), .A4(new_n2614_), .ZN(new_n2615_));
  OAI21_X1   g00180(.A1(new_n2603_), .A2(new_n2615_), .B(new_n2600_), .ZN(new_n2616_));
  NAND2_X1   g00181(.A1(new_n2616_), .A2(new_n2587_), .ZN(new_n2617_));
  NAND2_X1   g00182(.A1(new_n2558_), .A2(pi0221), .ZN(new_n2618_));
  NAND2_X1   g00183(.A1(new_n2618_), .A2(new_n2566_), .ZN(new_n2619_));
  INV_X1     g00184(.I(new_n2619_), .ZN(new_n2620_));
  NOR2_X1    g00185(.A1(pi0038), .A2(pi0100), .ZN(new_n2621_));
  INV_X1     g00186(.I(new_n2621_), .ZN(new_n2622_));
  NOR2_X1    g00187(.A1(pi0039), .A2(pi0087), .ZN(new_n2623_));
  INV_X1     g00188(.I(new_n2623_), .ZN(new_n2624_));
  NOR2_X1    g00189(.A1(new_n2622_), .A2(new_n2624_), .ZN(new_n2625_));
  NOR4_X1    g00190(.A1(new_n2625_), .A2(new_n2566_), .A3(pi0299), .A4(new_n2568_), .ZN(new_n2626_));
  NAND4_X1   g00191(.A1(new_n2586_), .A2(new_n2617_), .A3(new_n2620_), .A4(new_n2626_), .ZN(new_n2627_));
  INV_X1     g00192(.I(pi0075), .ZN(new_n2628_));
  INV_X1     g00193(.I(new_n2625_), .ZN(new_n2629_));
  NOR2_X1    g00194(.A1(new_n2629_), .A2(new_n2628_), .ZN(new_n2630_));
  INV_X1     g00195(.I(pi0210), .ZN(new_n2631_));
  INV_X1     g00196(.I(pi0032), .ZN(new_n2632_));
  INV_X1     g00197(.I(new_n2483_), .ZN(new_n2633_));
  NOR2_X1    g00198(.A1(new_n2464_), .A2(pi0081), .ZN(new_n2634_));
  NAND2_X1   g00199(.A1(new_n2500_), .A2(new_n2634_), .ZN(new_n2635_));
  NOR2_X1    g00200(.A1(new_n2635_), .A2(new_n2469_), .ZN(new_n2636_));
  INV_X1     g00201(.I(new_n2636_), .ZN(new_n2637_));
  NOR2_X1    g00202(.A1(pi0058), .A2(pi0091), .ZN(new_n2638_));
  NOR3_X1    g00203(.A1(pi0047), .A2(pi0109), .A3(pi0110), .ZN(new_n2639_));
  NAND2_X1   g00204(.A1(new_n2639_), .A2(new_n2638_), .ZN(new_n2640_));
  NOR2_X1    g00205(.A1(new_n2637_), .A2(new_n2640_), .ZN(new_n2641_));
  INV_X1     g00206(.I(new_n2641_), .ZN(new_n2642_));
  NOR2_X1    g00207(.A1(pi0070), .A2(pi0096), .ZN(new_n2643_));
  INV_X1     g00208(.I(new_n2643_), .ZN(new_n2644_));
  NOR2_X1    g00209(.A1(pi0035), .A2(pi0051), .ZN(new_n2645_));
  INV_X1     g00210(.I(new_n2645_), .ZN(new_n2646_));
  NOR2_X1    g00211(.A1(new_n2644_), .A2(new_n2646_), .ZN(new_n2647_));
  INV_X1     g00212(.I(new_n2647_), .ZN(new_n2648_));
  NOR2_X1    g00213(.A1(pi0090), .A2(pi0093), .ZN(new_n2649_));
  INV_X1     g00214(.I(new_n2649_), .ZN(new_n2650_));
  NOR2_X1    g00215(.A1(new_n2648_), .A2(new_n2650_), .ZN(new_n2651_));
  INV_X1     g00216(.I(new_n2651_), .ZN(new_n2652_));
  NOR2_X1    g00217(.A1(new_n2642_), .A2(new_n2652_), .ZN(new_n2653_));
  INV_X1     g00218(.I(new_n2653_), .ZN(new_n2654_));
  NOR2_X1    g00219(.A1(new_n2654_), .A2(new_n2633_), .ZN(new_n2655_));
  AOI21_X1   g00220(.A1(new_n2655_), .A2(pi0225), .B(new_n2632_), .ZN(new_n2656_));
  INV_X1     g00221(.I(new_n2656_), .ZN(new_n2657_));
  INV_X1     g00222(.I(pi0051), .ZN(new_n2658_));
  INV_X1     g00223(.I(pi0096), .ZN(new_n2659_));
  INV_X1     g00224(.I(pi0091), .ZN(new_n2660_));
  INV_X1     g00225(.I(pi0047), .ZN(new_n2661_));
  NOR2_X1    g00226(.A1(new_n2469_), .A2(new_n2472_), .ZN(new_n2662_));
  NAND2_X1   g00227(.A1(new_n2662_), .A2(new_n2661_), .ZN(new_n2663_));
  NOR2_X1    g00228(.A1(new_n2635_), .A2(new_n2663_), .ZN(new_n2664_));
  NOR2_X1    g00229(.A1(new_n2646_), .A2(pi0070), .ZN(new_n2665_));
  NOR2_X1    g00230(.A1(new_n2480_), .A2(pi0093), .ZN(new_n2666_));
  NAND4_X1   g00231(.A1(new_n2664_), .A2(new_n2660_), .A3(new_n2665_), .A4(new_n2666_), .ZN(new_n2667_));
  NOR2_X1    g00232(.A1(new_n2667_), .A2(new_n2659_), .ZN(new_n2668_));
  NOR2_X1    g00233(.A1(new_n2501_), .A2(new_n2480_), .ZN(new_n2669_));
  INV_X1     g00234(.I(new_n2669_), .ZN(new_n2670_));
  NOR2_X1    g00235(.A1(new_n2670_), .A2(new_n2478_), .ZN(new_n2671_));
  NAND4_X1   g00236(.A1(new_n2668_), .A2(new_n2671_), .A3(new_n2658_), .A4(new_n2483_), .ZN(new_n2672_));
  NOR3_X1    g00237(.A1(new_n2459_), .A2(new_n2476_), .A3(new_n2482_), .ZN(new_n2673_));
  NOR2_X1    g00238(.A1(new_n2673_), .A2(new_n2658_), .ZN(new_n2674_));
  NOR2_X1    g00239(.A1(new_n2674_), .A2(pi0096), .ZN(new_n2675_));
  INV_X1     g00240(.I(new_n2675_), .ZN(new_n2676_));
  NOR2_X1    g00241(.A1(pi0047), .A2(pi0110), .ZN(new_n2677_));
  INV_X1     g00242(.I(new_n2677_), .ZN(new_n2678_));
  NOR2_X1    g00243(.A1(new_n2636_), .A2(new_n2470_), .ZN(new_n2679_));
  INV_X1     g00244(.I(pi0097), .ZN(new_n2680_));
  NAND4_X1   g00245(.A1(new_n2500_), .A2(new_n2441_), .A3(new_n2462_), .A4(new_n2463_), .ZN(new_n2681_));
  NOR2_X1    g00246(.A1(pi0086), .A2(pi0094), .ZN(new_n2682_));
  INV_X1     g00247(.I(new_n2682_), .ZN(new_n2683_));
  NOR3_X1    g00248(.A1(pi0050), .A2(pi0053), .A3(pi0060), .ZN(new_n2684_));
  NAND2_X1   g00249(.A1(new_n2684_), .A2(new_n2461_), .ZN(new_n2685_));
  NOR2_X1    g00250(.A1(new_n2685_), .A2(new_n2683_), .ZN(new_n2686_));
  INV_X1     g00251(.I(new_n2686_), .ZN(new_n2687_));
  NOR2_X1    g00252(.A1(new_n2681_), .A2(new_n2687_), .ZN(new_n2688_));
  NOR2_X1    g00253(.A1(new_n2688_), .A2(new_n2680_), .ZN(new_n2689_));
  INV_X1     g00254(.I(new_n2689_), .ZN(new_n2690_));
  INV_X1     g00255(.I(pi0086), .ZN(new_n2691_));
  INV_X1     g00256(.I(pi0053), .ZN(new_n2692_));
  NOR2_X1    g00257(.A1(new_n2635_), .A2(pi0060), .ZN(new_n2693_));
  NOR2_X1    g00258(.A1(new_n2693_), .A2(new_n2692_), .ZN(new_n2694_));
  INV_X1     g00259(.I(new_n2635_), .ZN(new_n2695_));
  AOI21_X1   g00260(.A1(new_n2695_), .A2(pi0060), .B(pi0053), .ZN(new_n2696_));
  INV_X1     g00261(.I(new_n2696_), .ZN(new_n2697_));
  NAND2_X1   g00262(.A1(new_n2463_), .A2(new_n2461_), .ZN(new_n2698_));
  NAND3_X1   g00263(.A1(new_n2448_), .A2(new_n2453_), .A3(new_n2458_), .ZN(new_n2699_));
  NOR2_X1    g00264(.A1(pi0081), .A2(pi0102), .ZN(new_n2700_));
  INV_X1     g00265(.I(new_n2700_), .ZN(new_n2701_));
  NOR2_X1    g00266(.A1(new_n2699_), .A2(new_n2701_), .ZN(new_n2702_));
  INV_X1     g00267(.I(new_n2702_), .ZN(new_n2703_));
  NOR2_X1    g00268(.A1(new_n2703_), .A2(new_n2698_), .ZN(new_n2704_));
  INV_X1     g00269(.I(new_n2704_), .ZN(new_n2705_));
  AOI21_X1   g00270(.A1(new_n2705_), .A2(pi0050), .B(pi0060), .ZN(new_n2706_));
  NOR2_X1    g00271(.A1(new_n2681_), .A2(new_n2461_), .ZN(new_n2707_));
  NOR2_X1    g00272(.A1(new_n2707_), .A2(pi0050), .ZN(new_n2708_));
  INV_X1     g00273(.I(new_n2708_), .ZN(new_n2709_));
  INV_X1     g00274(.I(pi0088), .ZN(new_n2710_));
  OAI21_X1   g00275(.A1(new_n2702_), .A2(new_n2710_), .B(pi0098), .ZN(new_n2711_));
  NAND2_X1   g00276(.A1(new_n2711_), .A2(new_n2461_), .ZN(new_n2712_));
  INV_X1     g00277(.I(new_n2712_), .ZN(new_n2713_));
  NOR2_X1    g00278(.A1(new_n2441_), .A2(new_n2462_), .ZN(new_n2714_));
  OAI21_X1   g00279(.A1(new_n2699_), .A2(new_n2714_), .B(new_n2701_), .ZN(new_n2715_));
  NOR2_X1    g00280(.A1(new_n2443_), .A2(new_n2442_), .ZN(new_n2716_));
  OR3_X2     g00281(.A1(pi0082), .A2(pi0084), .A3(pi0111), .Z(new_n2717_));
  OR2_X2     g00282(.A1(pi0036), .A2(pi0068), .Z(new_n2718_));
  OR2_X2     g00283(.A1(pi0045), .A2(pi0104), .Z(new_n2719_));
  NOR3_X1    g00284(.A1(new_n2717_), .A2(new_n2718_), .A3(new_n2719_), .ZN(new_n2720_));
  NAND2_X1   g00285(.A1(new_n2720_), .A2(new_n2716_), .ZN(new_n2721_));
  NOR2_X1    g00286(.A1(new_n2721_), .A2(new_n2452_), .ZN(new_n2722_));
  INV_X1     g00287(.I(new_n2722_), .ZN(new_n2723_));
  INV_X1     g00288(.I(new_n2456_), .ZN(new_n2724_));
  NOR2_X1    g00289(.A1(new_n2723_), .A2(new_n2724_), .ZN(new_n2725_));
  AOI21_X1   g00290(.A1(new_n2725_), .A2(new_n2455_), .B(new_n2454_), .ZN(new_n2726_));
  INV_X1     g00291(.I(new_n2726_), .ZN(new_n2727_));
  INV_X1     g00292(.I(pi0073), .ZN(new_n2728_));
  NOR2_X1    g00293(.A1(new_n2499_), .A2(new_n2719_), .ZN(new_n2729_));
  NOR2_X1    g00294(.A1(new_n2729_), .A2(new_n2728_), .ZN(new_n2730_));
  INV_X1     g00295(.I(pi0066), .ZN(new_n2731_));
  INV_X1     g00296(.I(pi0045), .ZN(new_n2732_));
  NOR3_X1    g00297(.A1(new_n2499_), .A2(new_n2732_), .A3(pi0104), .ZN(new_n2733_));
  INV_X1     g00298(.I(pi0048), .ZN(new_n2734_));
  NAND2_X1   g00299(.A1(pi0085), .A2(pi0106), .ZN(new_n2735_));
  NAND4_X1   g00300(.A1(new_n2497_), .A2(new_n2492_), .A3(new_n2493_), .A4(new_n2735_), .ZN(new_n2736_));
  INV_X1     g00301(.I(new_n2497_), .ZN(new_n2737_));
  XOR2_X1    g00302(.A1(pi0061), .A2(pi0076), .Z(new_n2738_));
  NAND2_X1   g00303(.A1(new_n2735_), .A2(new_n2492_), .ZN(new_n2739_));
  AOI21_X1   g00304(.A1(new_n2737_), .A2(new_n2739_), .B(new_n2738_), .ZN(new_n2740_));
  NAND3_X1   g00305(.A1(new_n2740_), .A2(new_n2734_), .A3(new_n2736_), .ZN(new_n2741_));
  AOI21_X1   g00306(.A1(new_n2741_), .A2(new_n2442_), .B(pi0049), .ZN(new_n2742_));
  XNOR2_X1   g00307(.A1(new_n2742_), .A2(pi0089), .ZN(new_n2743_));
  NOR2_X1    g00308(.A1(new_n2442_), .A2(pi0048), .ZN(new_n2744_));
  INV_X1     g00309(.I(new_n2744_), .ZN(new_n2745_));
  NAND2_X1   g00310(.A1(new_n2743_), .A2(new_n2745_), .ZN(new_n2746_));
  INV_X1     g00311(.I(pi0104), .ZN(new_n2747_));
  XOR2_X1    g00312(.A1(new_n2716_), .A2(new_n2747_), .Z(new_n2748_));
  NAND2_X1   g00313(.A1(new_n2748_), .A2(new_n2732_), .ZN(new_n2749_));
  AOI21_X1   g00314(.A1(new_n2742_), .A2(pi0089), .B(new_n2749_), .ZN(new_n2750_));
  AOI21_X1   g00315(.A1(new_n2746_), .A2(new_n2750_), .B(new_n2733_), .ZN(new_n2751_));
  NOR2_X1    g00316(.A1(new_n2751_), .A2(new_n2728_), .ZN(new_n2752_));
  XOR2_X1    g00317(.A1(new_n2752_), .A2(new_n2729_), .Z(new_n2753_));
  NAND2_X1   g00318(.A1(new_n2753_), .A2(new_n2731_), .ZN(new_n2754_));
  NAND2_X1   g00319(.A1(new_n2754_), .A2(new_n2730_), .ZN(new_n2755_));
  NOR2_X1    g00320(.A1(new_n2754_), .A2(new_n2730_), .ZN(new_n2756_));
  INV_X1     g00321(.I(pi0068), .ZN(new_n2757_));
  INV_X1     g00322(.I(new_n2450_), .ZN(new_n2758_));
  INV_X1     g00323(.I(new_n2729_), .ZN(new_n2759_));
  NOR3_X1    g00324(.A1(new_n2759_), .A2(pi0084), .A3(new_n2758_), .ZN(new_n2760_));
  OAI21_X1   g00325(.A1(new_n2760_), .A2(new_n2757_), .B(pi0111), .ZN(new_n2761_));
  NOR2_X1    g00326(.A1(new_n2759_), .A2(new_n2758_), .ZN(new_n2762_));
  NAND2_X1   g00327(.A1(new_n2762_), .A2(pi0084), .ZN(new_n2763_));
  NOR2_X1    g00328(.A1(pi0068), .A2(pi0111), .ZN(new_n2764_));
  NAND3_X1   g00329(.A1(new_n2760_), .A2(pi0082), .A3(new_n2764_), .ZN(new_n2765_));
  INV_X1     g00330(.I(pi0084), .ZN(new_n2766_));
  INV_X1     g00331(.I(pi0036), .ZN(new_n2767_));
  INV_X1     g00332(.I(pi0067), .ZN(new_n2768_));
  NAND2_X1   g00333(.A1(new_n2767_), .A2(new_n2768_), .ZN(new_n2769_));
  INV_X1     g00334(.I(new_n2769_), .ZN(new_n2770_));
  NOR4_X1    g00335(.A1(new_n2770_), .A2(pi0082), .A3(new_n2766_), .A4(new_n2764_), .ZN(new_n2771_));
  NAND4_X1   g00336(.A1(new_n2761_), .A2(new_n2765_), .A3(new_n2763_), .A4(new_n2771_), .ZN(new_n2772_));
  NOR2_X1    g00337(.A1(new_n2756_), .A2(new_n2772_), .ZN(new_n2773_));
  NAND2_X1   g00338(.A1(new_n2773_), .A2(new_n2755_), .ZN(new_n2774_));
  NOR2_X1    g00339(.A1(pi0082), .A2(pi0111), .ZN(new_n2775_));
  INV_X1     g00340(.I(new_n2760_), .ZN(new_n2776_));
  NOR2_X1    g00341(.A1(new_n2776_), .A2(pi0068), .ZN(new_n2777_));
  AOI21_X1   g00342(.A1(new_n2777_), .A2(new_n2775_), .B(new_n2767_), .ZN(new_n2778_));
  NOR2_X1    g00343(.A1(new_n2721_), .A2(new_n2758_), .ZN(new_n2779_));
  INV_X1     g00344(.I(new_n2779_), .ZN(new_n2780_));
  AOI21_X1   g00345(.A1(pi0067), .A2(new_n2780_), .B(new_n2778_), .ZN(new_n2781_));
  NAND2_X1   g00346(.A1(new_n2774_), .A2(new_n2781_), .ZN(new_n2782_));
  INV_X1     g00347(.I(pi0069), .ZN(new_n2783_));
  INV_X1     g00348(.I(pi0083), .ZN(new_n2784_));
  NAND2_X1   g00349(.A1(new_n2783_), .A2(new_n2784_), .ZN(new_n2785_));
  INV_X1     g00350(.I(new_n2451_), .ZN(new_n2786_));
  NOR2_X1    g00351(.A1(new_n2780_), .A2(new_n2786_), .ZN(new_n2787_));
  INV_X1     g00352(.I(new_n2787_), .ZN(new_n2788_));
  AOI21_X1   g00353(.A1(new_n2788_), .A2(pi0083), .B(pi0103), .ZN(new_n2789_));
  INV_X1     g00354(.I(new_n2789_), .ZN(new_n2790_));
  AOI21_X1   g00355(.A1(new_n2790_), .A2(new_n2787_), .B(new_n2785_), .ZN(new_n2791_));
  NAND2_X1   g00356(.A1(new_n2782_), .A2(new_n2791_), .ZN(new_n2792_));
  AOI21_X1   g00357(.A1(new_n2723_), .A2(pi0071), .B(pi0065), .ZN(new_n2793_));
  INV_X1     g00358(.I(new_n2793_), .ZN(new_n2794_));
  INV_X1     g00359(.I(pi0103), .ZN(new_n2795_));
  NOR4_X1    g00360(.A1(new_n2780_), .A2(pi0067), .A3(new_n2795_), .A4(new_n2785_), .ZN(new_n2796_));
  NOR3_X1    g00361(.A1(new_n2794_), .A2(pi0071), .A3(new_n2796_), .ZN(new_n2797_));
  AOI21_X1   g00362(.A1(new_n2792_), .A2(new_n2797_), .B(pi0107), .ZN(new_n2798_));
  INV_X1     g00363(.I(pi0063), .ZN(new_n2799_));
  INV_X1     g00364(.I(pi0107), .ZN(new_n2800_));
  OAI21_X1   g00365(.A1(new_n2725_), .A2(new_n2800_), .B(new_n2799_), .ZN(new_n2801_));
  NOR4_X1    g00366(.A1(new_n2723_), .A2(new_n2799_), .A3(pi0107), .A4(new_n2724_), .ZN(new_n2802_));
  OR3_X2     g00367(.A1(new_n2801_), .A2(pi0064), .A3(new_n2802_), .Z(new_n2803_));
  OAI21_X1   g00368(.A1(new_n2798_), .A2(new_n2803_), .B(new_n2727_), .ZN(new_n2804_));
  INV_X1     g00369(.I(new_n2804_), .ZN(new_n2805_));
  INV_X1     g00370(.I(pi0065), .ZN(new_n2806_));
  NOR3_X1    g00371(.A1(new_n2723_), .A2(new_n2806_), .A3(pi0071), .ZN(new_n2807_));
  INV_X1     g00372(.I(new_n2807_), .ZN(new_n2808_));
  NAND3_X1   g00373(.A1(new_n2798_), .A2(new_n2801_), .A3(new_n2808_), .ZN(new_n2809_));
  NOR2_X1    g00374(.A1(new_n2700_), .A2(pi0064), .ZN(new_n2810_));
  NAND4_X1   g00375(.A1(new_n2805_), .A2(new_n2727_), .A3(new_n2809_), .A4(new_n2810_), .ZN(new_n2811_));
  NAND2_X1   g00376(.A1(new_n2811_), .A2(new_n2715_), .ZN(new_n2812_));
  AOI21_X1   g00377(.A1(new_n2812_), .A2(new_n2463_), .B(new_n2713_), .ZN(new_n2813_));
  OAI21_X1   g00378(.A1(new_n2813_), .A2(new_n2709_), .B(new_n2706_), .ZN(new_n2814_));
  INV_X1     g00379(.I(new_n2814_), .ZN(new_n2815_));
  NOR2_X1    g00380(.A1(new_n2815_), .A2(new_n2697_), .ZN(new_n2816_));
  OAI21_X1   g00381(.A1(new_n2816_), .A2(new_n2694_), .B(new_n2691_), .ZN(new_n2817_));
  AND2_X2    g00382(.A1(new_n2704_), .A2(new_n2684_), .Z(new_n2818_));
  INV_X1     g00383(.I(new_n2818_), .ZN(new_n2819_));
  NOR3_X1    g00384(.A1(new_n2819_), .A2(pi0086), .A3(new_n2466_), .ZN(new_n2820_));
  NOR2_X1    g00385(.A1(new_n2820_), .A2(pi0097), .ZN(new_n2821_));
  AOI21_X1   g00386(.A1(new_n2819_), .A2(pi0086), .B(pi0094), .ZN(new_n2822_));
  INV_X1     g00387(.I(new_n2822_), .ZN(new_n2823_));
  NOR2_X1    g00388(.A1(new_n2821_), .A2(new_n2823_), .ZN(new_n2824_));
  NAND2_X1   g00389(.A1(new_n2817_), .A2(new_n2824_), .ZN(new_n2825_));
  NAND2_X1   g00390(.A1(new_n2825_), .A2(new_n2690_), .ZN(new_n2826_));
  INV_X1     g00391(.I(new_n2688_), .ZN(new_n2827_));
  NOR2_X1    g00392(.A1(new_n2827_), .A2(pi0097), .ZN(new_n2828_));
  NOR2_X1    g00393(.A1(new_n2465_), .A2(pi0108), .ZN(new_n2829_));
  NAND2_X1   g00394(.A1(new_n2826_), .A2(new_n2829_), .ZN(new_n2830_));
  INV_X1     g00395(.I(new_n2468_), .ZN(new_n2831_));
  NOR3_X1    g00396(.A1(new_n2827_), .A2(new_n2465_), .A3(new_n2831_), .ZN(new_n2832_));
  NOR2_X1    g00397(.A1(new_n2832_), .A2(pi0109), .ZN(new_n2833_));
  AOI21_X1   g00398(.A1(new_n2830_), .A2(new_n2833_), .B(new_n2679_), .ZN(new_n2834_));
  AOI21_X1   g00399(.A1(new_n2636_), .A2(new_n2470_), .B(new_n2471_), .ZN(new_n2835_));
  NOR2_X1    g00400(.A1(new_n2664_), .A2(pi0091), .ZN(new_n2836_));
  NOR2_X1    g00401(.A1(new_n2835_), .A2(new_n2836_), .ZN(new_n2837_));
  INV_X1     g00402(.I(new_n2837_), .ZN(new_n2838_));
  INV_X1     g00403(.I(pi0090), .ZN(new_n2839_));
  NOR2_X1    g00404(.A1(new_n2641_), .A2(new_n2839_), .ZN(new_n2840_));
  INV_X1     g00405(.I(pi0093), .ZN(new_n2841_));
  OAI21_X1   g00406(.A1(new_n2501_), .A2(pi0058), .B(new_n2841_), .ZN(new_n2842_));
  INV_X1     g00407(.I(new_n2664_), .ZN(new_n2843_));
  NOR2_X1    g00408(.A1(new_n2843_), .A2(new_n2660_), .ZN(new_n2844_));
  NOR2_X1    g00409(.A1(new_n2844_), .A2(new_n2480_), .ZN(new_n2845_));
  NOR4_X1    g00410(.A1(new_n2838_), .A2(new_n2840_), .A3(new_n2845_), .A4(new_n2842_), .ZN(new_n2846_));
  OAI21_X1   g00411(.A1(new_n2834_), .A2(new_n2678_), .B(new_n2846_), .ZN(new_n2847_));
  AOI21_X1   g00412(.A1(new_n2669_), .A2(pi0093), .B(pi0035), .ZN(new_n2848_));
  INV_X1     g00413(.I(pi0070), .ZN(new_n2849_));
  INV_X1     g00414(.I(pi0225), .ZN(new_n2850_));
  NOR2_X1    g00415(.A1(new_n2670_), .A2(pi0093), .ZN(new_n2851_));
  INV_X1     g00416(.I(new_n2851_), .ZN(new_n2852_));
  OAI21_X1   g00417(.A1(new_n2852_), .A2(new_n2850_), .B(pi0035), .ZN(new_n2853_));
  NAND2_X1   g00418(.A1(new_n2853_), .A2(new_n2849_), .ZN(new_n2854_));
  AOI21_X1   g00419(.A1(new_n2847_), .A2(new_n2848_), .B(new_n2854_), .ZN(new_n2855_));
  NOR2_X1    g00420(.A1(new_n2855_), .A2(pi0051), .ZN(new_n2856_));
  NOR2_X1    g00421(.A1(new_n2856_), .A2(new_n2676_), .ZN(new_n2857_));
  NAND2_X1   g00422(.A1(new_n2510_), .A2(pi0040), .ZN(new_n2858_));
  INV_X1     g00423(.I(new_n2858_), .ZN(new_n2859_));
  NOR2_X1    g00424(.A1(new_n2859_), .A2(pi0032), .ZN(new_n2860_));
  INV_X1     g00425(.I(pi0072), .ZN(new_n2861_));
  NOR2_X1    g00426(.A1(new_n2653_), .A2(new_n2861_), .ZN(new_n2862_));
  NOR2_X1    g00427(.A1(new_n2862_), .A2(pi0040), .ZN(new_n2863_));
  INV_X1     g00428(.I(new_n2863_), .ZN(new_n2864_));
  NOR2_X1    g00429(.A1(new_n2864_), .A2(new_n2860_), .ZN(new_n2865_));
  OAI21_X1   g00430(.A1(new_n2857_), .A2(pi0072), .B(new_n2865_), .ZN(new_n2866_));
  INV_X1     g00431(.I(new_n2866_), .ZN(new_n2867_));
  NAND2_X1   g00432(.A1(new_n2867_), .A2(new_n2672_), .ZN(new_n2868_));
  AOI21_X1   g00433(.A1(new_n2868_), .A2(new_n2657_), .B(pi0095), .ZN(new_n2869_));
  INV_X1     g00434(.I(pi0479), .ZN(new_n2870_));
  AOI21_X1   g00435(.A1(new_n2510_), .A2(new_n2512_), .B(new_n2437_), .ZN(new_n2871_));
  INV_X1     g00436(.I(new_n2871_), .ZN(new_n2872_));
  NOR2_X1    g00437(.A1(new_n2872_), .A2(new_n2870_), .ZN(new_n2873_));
  NOR3_X1    g00438(.A1(new_n2869_), .A2(new_n2436_), .A3(new_n2873_), .ZN(new_n2874_));
  AOI21_X1   g00439(.A1(new_n2667_), .A2(pi0096), .B(new_n2633_), .ZN(new_n2875_));
  INV_X1     g00440(.I(pi0035), .ZN(new_n2876_));
  NOR2_X1    g00441(.A1(new_n2876_), .A2(pi0225), .ZN(new_n2877_));
  AOI21_X1   g00442(.A1(new_n2851_), .A2(new_n2877_), .B(pi0070), .ZN(new_n2878_));
  NOR2_X1    g00443(.A1(new_n2878_), .A2(pi0051), .ZN(new_n2879_));
  INV_X1     g00444(.I(new_n2879_), .ZN(new_n2880_));
  AOI21_X1   g00445(.A1(pi0035), .A2(new_n2852_), .B(new_n2880_), .ZN(new_n2881_));
  INV_X1     g00446(.I(new_n2881_), .ZN(new_n2882_));
  NOR2_X1    g00447(.A1(new_n2694_), .A2(new_n2683_), .ZN(new_n2883_));
  INV_X1     g00448(.I(new_n2883_), .ZN(new_n2884_));
  NOR2_X1    g00449(.A1(pi0046), .A2(pi0109), .ZN(new_n2885_));
  INV_X1     g00450(.I(new_n2885_), .ZN(new_n2886_));
  NOR2_X1    g00451(.A1(new_n2886_), .A2(pi0110), .ZN(new_n2887_));
  NAND3_X1   g00452(.A1(new_n2887_), .A2(new_n2468_), .A3(new_n2473_), .ZN(new_n2888_));
  NOR2_X1    g00453(.A1(new_n2888_), .A2(pi0058), .ZN(new_n2889_));
  INV_X1     g00454(.I(new_n2889_), .ZN(new_n2890_));
  NOR4_X1    g00455(.A1(new_n2884_), .A2(new_n2650_), .A3(new_n2696_), .A4(new_n2890_), .ZN(new_n2891_));
  NOR2_X1    g00456(.A1(new_n2891_), .A2(pi0035), .ZN(new_n2892_));
  NOR2_X1    g00457(.A1(new_n2882_), .A2(new_n2892_), .ZN(new_n2893_));
  NOR2_X1    g00458(.A1(new_n2893_), .A2(pi0096), .ZN(new_n2894_));
  INV_X1     g00459(.I(new_n2894_), .ZN(new_n2895_));
  AOI21_X1   g00460(.A1(new_n2895_), .A2(new_n2875_), .B(pi0032), .ZN(new_n2896_));
  OAI21_X1   g00461(.A1(new_n2896_), .A2(new_n2656_), .B(new_n2437_), .ZN(new_n2897_));
  OAI21_X1   g00462(.A1(new_n2437_), .A2(new_n2870_), .B(new_n2897_), .ZN(new_n2898_));
  NOR2_X1    g00463(.A1(new_n2898_), .A2(pi0137), .ZN(new_n2899_));
  NOR2_X1    g00464(.A1(new_n2874_), .A2(new_n2899_), .ZN(new_n2900_));
  NOR2_X1    g00465(.A1(new_n2900_), .A2(new_n2631_), .ZN(new_n2901_));
  INV_X1     g00466(.I(pi0841), .ZN(new_n2902_));
  NOR2_X1    g00467(.A1(new_n2852_), .A2(new_n2902_), .ZN(new_n2903_));
  INV_X1     g00468(.I(new_n2903_), .ZN(new_n2904_));
  NOR3_X1    g00469(.A1(new_n2904_), .A2(pi0051), .A3(pi0072), .ZN(new_n2905_));
  NOR2_X1    g00470(.A1(pi0035), .A2(pi0040), .ZN(new_n2906_));
  INV_X1     g00471(.I(new_n2906_), .ZN(new_n2907_));
  NOR3_X1    g00472(.A1(new_n2644_), .A2(new_n2907_), .A3(new_n2850_), .ZN(new_n2908_));
  AOI21_X1   g00473(.A1(new_n2905_), .A2(new_n2908_), .B(new_n2632_), .ZN(new_n2909_));
  INV_X1     g00474(.I(new_n2909_), .ZN(new_n2910_));
  AOI21_X1   g00475(.A1(new_n2868_), .A2(new_n2910_), .B(pi0095), .ZN(new_n2911_));
  OAI21_X1   g00476(.A1(new_n2911_), .A2(new_n2873_), .B(pi0137), .ZN(new_n2912_));
  NOR2_X1    g00477(.A1(new_n2896_), .A2(new_n2909_), .ZN(new_n2913_));
  NOR2_X1    g00478(.A1(new_n2913_), .A2(pi0095), .ZN(new_n2914_));
  AOI21_X1   g00479(.A1(pi0095), .A2(pi0479), .B(new_n2914_), .ZN(new_n2915_));
  NAND2_X1   g00480(.A1(new_n2915_), .A2(new_n2436_), .ZN(new_n2916_));
  NAND2_X1   g00481(.A1(new_n2912_), .A2(new_n2916_), .ZN(new_n2917_));
  INV_X1     g00482(.I(pi1091), .ZN(new_n2918_));
  INV_X1     g00483(.I(pi0957), .ZN(new_n2919_));
  NOR2_X1    g00484(.A1(new_n2919_), .A2(pi0833), .ZN(new_n2920_));
  NOR2_X1    g00485(.A1(new_n2920_), .A2(new_n2918_), .ZN(new_n2921_));
  INV_X1     g00486(.I(new_n2921_), .ZN(new_n2922_));
  INV_X1     g00487(.I(pi1092), .ZN(new_n2923_));
  INV_X1     g00488(.I(pi1093), .ZN(new_n2924_));
  NOR2_X1    g00489(.A1(new_n2923_), .A2(new_n2924_), .ZN(new_n2925_));
  INV_X1     g00490(.I(new_n2925_), .ZN(new_n2926_));
  INV_X1     g00491(.I(pi0829), .ZN(new_n2927_));
  INV_X1     g00492(.I(pi0950), .ZN(new_n2928_));
  NOR2_X1    g00493(.A1(new_n2927_), .A2(new_n2928_), .ZN(new_n2929_));
  INV_X1     g00494(.I(new_n2929_), .ZN(new_n2930_));
  NOR2_X1    g00495(.A1(new_n2926_), .A2(new_n2930_), .ZN(new_n2931_));
  INV_X1     g00496(.I(new_n2931_), .ZN(new_n2932_));
  OAI21_X1   g00497(.A1(new_n2884_), .A2(new_n2696_), .B(new_n2680_), .ZN(new_n2933_));
  NOR3_X1    g00498(.A1(new_n2689_), .A2(pi0108), .A3(pi0110), .ZN(new_n2934_));
  NOR2_X1    g00499(.A1(new_n2474_), .A2(new_n2886_), .ZN(new_n2935_));
  INV_X1     g00500(.I(new_n2935_), .ZN(new_n2936_));
  NAND4_X1   g00501(.A1(new_n2933_), .A2(new_n2666_), .A3(new_n2934_), .A4(new_n2936_), .ZN(new_n2937_));
  NAND2_X1   g00502(.A1(new_n2937_), .A2(new_n2876_), .ZN(new_n2938_));
  OAI21_X1   g00503(.A1(new_n2882_), .A2(new_n2938_), .B(new_n2659_), .ZN(new_n2939_));
  NAND2_X1   g00504(.A1(new_n2939_), .A2(new_n2875_), .ZN(new_n2940_));
  NAND2_X1   g00505(.A1(new_n2940_), .A2(new_n2632_), .ZN(new_n2941_));
  NAND2_X1   g00506(.A1(new_n2941_), .A2(new_n2910_), .ZN(new_n2942_));
  MUX2_X1    g00507(.I0(new_n2942_), .I1(pi0479), .S(pi0095), .Z(new_n2943_));
  NOR2_X1    g00508(.A1(new_n2943_), .A2(new_n2932_), .ZN(new_n2944_));
  OAI21_X1   g00509(.A1(new_n2915_), .A2(new_n2931_), .B(new_n2436_), .ZN(new_n2945_));
  NOR2_X1    g00510(.A1(new_n2945_), .A2(new_n2944_), .ZN(new_n2946_));
  NAND2_X1   g00511(.A1(new_n2912_), .A2(new_n2946_), .ZN(new_n2947_));
  MUX2_X1    g00512(.I0(new_n2947_), .I1(new_n2917_), .S(new_n2922_), .Z(new_n2948_));
  AOI21_X1   g00513(.A1(new_n2948_), .A2(new_n2631_), .B(new_n2901_), .ZN(new_n2949_));
  NOR2_X1    g00514(.A1(new_n2871_), .A2(new_n2438_), .ZN(new_n2950_));
  NAND2_X1   g00515(.A1(new_n2866_), .A2(new_n2910_), .ZN(new_n2951_));
  NAND2_X1   g00516(.A1(new_n2951_), .A2(new_n2437_), .ZN(new_n2952_));
  AOI21_X1   g00517(.A1(new_n2952_), .A2(new_n2950_), .B(new_n2436_), .ZN(new_n2953_));
  INV_X1     g00518(.I(new_n2953_), .ZN(new_n2954_));
  NAND2_X1   g00519(.A1(pi0950), .A2(pi1092), .ZN(new_n2955_));
  NOR2_X1    g00520(.A1(new_n2955_), .A2(new_n2927_), .ZN(new_n2956_));
  INV_X1     g00521(.I(new_n2956_), .ZN(new_n2957_));
  INV_X1     g00522(.I(new_n2920_), .ZN(new_n2958_));
  NOR2_X1    g00523(.A1(new_n2918_), .A2(new_n2924_), .ZN(new_n2959_));
  NAND2_X1   g00524(.A1(new_n2958_), .A2(new_n2959_), .ZN(new_n2960_));
  NOR3_X1    g00525(.A1(new_n2938_), .A2(new_n2957_), .A3(new_n2960_), .ZN(new_n2961_));
  NOR2_X1    g00526(.A1(new_n2503_), .A2(pi0040), .ZN(new_n2962_));
  INV_X1     g00527(.I(new_n2962_), .ZN(new_n2963_));
  NOR2_X1    g00528(.A1(new_n2932_), .A2(new_n2922_), .ZN(new_n2964_));
  NOR2_X1    g00529(.A1(new_n2892_), .A2(new_n2964_), .ZN(new_n2965_));
  NOR4_X1    g00530(.A1(new_n2961_), .A2(new_n2882_), .A3(new_n2963_), .A4(new_n2965_), .ZN(new_n2966_));
  NAND2_X1   g00531(.A1(new_n2632_), .A2(new_n2437_), .ZN(new_n2967_));
  OAI21_X1   g00532(.A1(new_n2966_), .A2(new_n2967_), .B(new_n2436_), .ZN(new_n2968_));
  NAND2_X1   g00533(.A1(new_n2954_), .A2(new_n2968_), .ZN(new_n2969_));
  NAND2_X1   g00534(.A1(new_n2893_), .A2(new_n2962_), .ZN(new_n2970_));
  NAND2_X1   g00535(.A1(new_n2970_), .A2(new_n2632_), .ZN(new_n2971_));
  NOR2_X1    g00536(.A1(new_n2656_), .A2(pi0095), .ZN(new_n2972_));
  AOI21_X1   g00537(.A1(new_n2971_), .A2(new_n2972_), .B(pi0137), .ZN(new_n2973_));
  INV_X1     g00538(.I(new_n2438_), .ZN(new_n2974_));
  NOR2_X1    g00539(.A1(new_n2974_), .A2(pi0095), .ZN(new_n2975_));
  OAI21_X1   g00540(.A1(new_n2867_), .A2(new_n2656_), .B(new_n2975_), .ZN(new_n2976_));
  AOI21_X1   g00541(.A1(new_n2976_), .A2(pi0137), .B(new_n2973_), .ZN(new_n2977_));
  NAND2_X1   g00542(.A1(new_n2977_), .A2(pi0210), .ZN(new_n2978_));
  OAI21_X1   g00543(.A1(new_n2969_), .A2(pi0210), .B(new_n2978_), .ZN(new_n2979_));
  INV_X1     g00544(.I(new_n2979_), .ZN(new_n2980_));
  AOI21_X1   g00545(.A1(new_n2440_), .A2(new_n2980_), .B(new_n2949_), .ZN(new_n2981_));
  NAND3_X1   g00546(.A1(new_n2949_), .A2(new_n2440_), .A3(new_n2979_), .ZN(new_n2982_));
  NAND2_X1   g00547(.A1(new_n2982_), .A2(new_n2563_), .ZN(new_n2983_));
  OAI21_X1   g00548(.A1(new_n2983_), .A2(new_n2981_), .B(new_n2576_), .ZN(new_n2984_));
  INV_X1     g00549(.I(new_n2576_), .ZN(new_n2985_));
  INV_X1     g00550(.I(new_n2608_), .ZN(new_n2986_));
  INV_X1     g00551(.I(new_n2900_), .ZN(new_n2989_));
  NAND2_X1   g00552(.A1(new_n2986_), .A2(pi0146), .ZN(new_n2991_));
  INV_X1     g00553(.I(new_n2611_), .ZN(new_n2992_));
  NOR2_X1    g00554(.A1(new_n2909_), .A2(pi0095), .ZN(new_n2993_));
  INV_X1     g00555(.I(new_n2993_), .ZN(new_n2994_));
  INV_X1     g00556(.I(new_n2971_), .ZN(new_n2995_));
  NOR2_X1    g00557(.A1(new_n2995_), .A2(new_n2994_), .ZN(new_n2996_));
  INV_X1     g00558(.I(new_n2996_), .ZN(new_n2997_));
  NAND2_X1   g00559(.A1(new_n2997_), .A2(new_n2436_), .ZN(new_n2998_));
  NAND3_X1   g00560(.A1(new_n2979_), .A2(pi0146), .A3(new_n2992_), .ZN(new_n3003_));
  OAI21_X1   g00561(.A1(new_n2949_), .A2(new_n2991_), .B(new_n3003_), .ZN(new_n3004_));
  AOI21_X1   g00562(.A1(new_n3004_), .A2(new_n2985_), .B(new_n2522_), .ZN(new_n3005_));
  OAI21_X1   g00563(.A1(new_n2527_), .A2(pi0105), .B(new_n2523_), .ZN(new_n3006_));
  AOI21_X1   g00564(.A1(new_n2984_), .A2(new_n3005_), .B(new_n3006_), .ZN(new_n3007_));
  INV_X1     g00565(.I(new_n2865_), .ZN(new_n3008_));
  NOR3_X1    g00566(.A1(new_n2636_), .A2(new_n2470_), .A3(new_n2677_), .ZN(new_n3009_));
  NAND2_X1   g00567(.A1(new_n2830_), .A2(new_n3009_), .ZN(new_n3010_));
  NAND2_X1   g00568(.A1(new_n3010_), .A2(new_n2846_), .ZN(new_n3011_));
  NAND2_X1   g00569(.A1(new_n3011_), .A2(new_n2848_), .ZN(new_n3012_));
  INV_X1     g00570(.I(new_n3012_), .ZN(new_n3013_));
  OAI21_X1   g00571(.A1(new_n3013_), .A2(new_n2854_), .B(new_n2658_), .ZN(new_n3014_));
  AOI21_X1   g00572(.A1(new_n3014_), .A2(new_n2675_), .B(pi0072), .ZN(new_n3015_));
  NOR2_X1    g00573(.A1(new_n3015_), .A2(new_n3008_), .ZN(new_n3016_));
  AND2_X2    g00574(.A1(new_n3016_), .A2(new_n2672_), .Z(new_n3017_));
  OAI21_X1   g00575(.A1(new_n3017_), .A2(new_n2909_), .B(new_n2437_), .ZN(new_n3018_));
  AOI21_X1   g00576(.A1(new_n3018_), .A2(new_n2872_), .B(new_n2436_), .ZN(new_n3019_));
  NOR4_X1    g00577(.A1(new_n2871_), .A2(new_n2577_), .A3(new_n2922_), .A4(new_n2932_), .ZN(new_n3020_));
  NOR3_X1    g00578(.A1(new_n2871_), .A2(new_n2577_), .A3(new_n2922_), .ZN(new_n3021_));
  AOI22_X1   g00579(.A1(new_n2915_), .A2(new_n3020_), .B1(new_n2944_), .B2(new_n3021_), .ZN(new_n3022_));
  OAI21_X1   g00580(.A1(new_n3022_), .A2(pi0137), .B(new_n2631_), .ZN(new_n3023_));
  OAI21_X1   g00581(.A1(new_n3015_), .A2(new_n3008_), .B(new_n2910_), .ZN(new_n3024_));
  INV_X1     g00582(.I(new_n2577_), .ZN(new_n3025_));
  NOR2_X1    g00583(.A1(new_n2998_), .A2(new_n3025_), .ZN(new_n3026_));
  AOI21_X1   g00584(.A1(new_n2631_), .A2(new_n2440_), .B(new_n3025_), .ZN(new_n3027_));
  NAND2_X1   g00585(.A1(new_n2968_), .A2(new_n3027_), .ZN(new_n3028_));
  OAI21_X1   g00586(.A1(new_n3026_), .A2(new_n3028_), .B(pi0137), .ZN(new_n3029_));
  AOI21_X1   g00587(.A1(new_n3024_), .A2(new_n2975_), .B(new_n3029_), .ZN(new_n3030_));
  NOR2_X1    g00588(.A1(new_n3016_), .A2(new_n2656_), .ZN(new_n3031_));
  INV_X1     g00589(.I(new_n2950_), .ZN(new_n3032_));
  INV_X1     g00590(.I(new_n2973_), .ZN(new_n3033_));
  NAND4_X1   g00591(.A1(new_n3033_), .A2(new_n2631_), .A3(new_n2609_), .A4(new_n3032_), .ZN(new_n3034_));
  OAI21_X1   g00592(.A1(new_n3031_), .A2(new_n3034_), .B(pi0234), .ZN(new_n3035_));
  NOR2_X1    g00593(.A1(new_n3035_), .A2(new_n3030_), .ZN(new_n3036_));
  OAI21_X1   g00594(.A1(new_n3019_), .A2(new_n3023_), .B(new_n3036_), .ZN(new_n3037_));
  NOR2_X1    g00595(.A1(new_n3017_), .A2(new_n2656_), .ZN(new_n3038_));
  NAND2_X1   g00596(.A1(new_n2437_), .A2(new_n2436_), .ZN(new_n3039_));
  NOR2_X1    g00597(.A1(new_n2871_), .A2(pi0137), .ZN(new_n3040_));
  INV_X1     g00598(.I(new_n3040_), .ZN(new_n3041_));
  NAND2_X1   g00599(.A1(pi0210), .A2(pi0234), .ZN(new_n3042_));
  AOI21_X1   g00600(.A1(new_n2898_), .A2(new_n3041_), .B(new_n3042_), .ZN(new_n3043_));
  OAI21_X1   g00601(.A1(new_n3038_), .A2(new_n3039_), .B(new_n3043_), .ZN(new_n3044_));
  NAND2_X1   g00602(.A1(new_n3037_), .A2(new_n3044_), .ZN(new_n3045_));
  NOR2_X1    g00603(.A1(pi0032), .A2(pi0225), .ZN(new_n3046_));
  AOI21_X1   g00604(.A1(new_n2655_), .A2(new_n3046_), .B(pi0095), .ZN(new_n3047_));
  INV_X1     g00605(.I(new_n3047_), .ZN(new_n3048_));
  INV_X1     g00606(.I(new_n3009_), .ZN(new_n3049_));
  INV_X1     g00607(.I(new_n2829_), .ZN(new_n3050_));
  AOI21_X1   g00608(.A1(new_n2815_), .A2(new_n2692_), .B(pi0086), .ZN(new_n3051_));
  OAI21_X1   g00609(.A1(new_n3051_), .A2(new_n2823_), .B(new_n2821_), .ZN(new_n3052_));
  AOI21_X1   g00610(.A1(new_n3052_), .A2(new_n2690_), .B(new_n3050_), .ZN(new_n3053_));
  AOI21_X1   g00611(.A1(pi0058), .A2(new_n2501_), .B(new_n2840_), .ZN(new_n3054_));
  NOR3_X1    g00612(.A1(new_n3054_), .A2(new_n2838_), .A3(new_n2845_), .ZN(new_n3055_));
  OAI21_X1   g00613(.A1(new_n3053_), .A2(new_n3049_), .B(new_n3055_), .ZN(new_n3056_));
  MUX2_X1    g00614(.I0(new_n3056_), .I1(new_n2670_), .S(pi0093), .Z(new_n3057_));
  NOR2_X1    g00615(.A1(new_n3057_), .A2(pi0035), .ZN(new_n3058_));
  NOR2_X1    g00616(.A1(new_n2671_), .A2(new_n2849_), .ZN(new_n3059_));
  INV_X1     g00617(.I(new_n3059_), .ZN(new_n3060_));
  NAND4_X1   g00618(.A1(new_n3058_), .A2(new_n2676_), .A3(new_n2880_), .A4(new_n3060_), .ZN(new_n3061_));
  AOI21_X1   g00619(.A1(new_n3061_), .A2(new_n2861_), .B(new_n3008_), .ZN(new_n3062_));
  NOR2_X1    g00620(.A1(new_n3032_), .A2(pi0137), .ZN(new_n3063_));
  OAI21_X1   g00621(.A1(new_n3062_), .A2(new_n3048_), .B(new_n3063_), .ZN(new_n3064_));
  NOR2_X1    g00622(.A1(new_n3059_), .A2(new_n2487_), .ZN(new_n3065_));
  INV_X1     g00623(.I(new_n3065_), .ZN(new_n3066_));
  NAND2_X1   g00624(.A1(new_n2878_), .A2(new_n2483_), .ZN(new_n3067_));
  OAI21_X1   g00625(.A1(new_n3066_), .A2(new_n3067_), .B(new_n2632_), .ZN(new_n3068_));
  NOR4_X1    g00626(.A1(new_n3047_), .A2(new_n2436_), .A3(pi0210), .A4(new_n3068_), .ZN(new_n3069_));
  AOI21_X1   g00627(.A1(new_n3064_), .A2(new_n3069_), .B(new_n2986_), .ZN(new_n3070_));
  INV_X1     g00628(.I(new_n3070_), .ZN(new_n3071_));
  NOR2_X1    g00629(.A1(pi0146), .A2(pi0210), .ZN(new_n3072_));
  NOR4_X1    g00630(.A1(new_n2655_), .A2(pi0032), .A3(new_n2850_), .A4(new_n2902_), .ZN(new_n3073_));
  NOR2_X1    g00631(.A1(new_n3073_), .A2(pi0095), .ZN(new_n3074_));
  INV_X1     g00632(.I(new_n3074_), .ZN(new_n3075_));
  OAI21_X1   g00633(.A1(new_n3075_), .A2(new_n3068_), .B(pi0137), .ZN(new_n3076_));
  INV_X1     g00634(.I(new_n2975_), .ZN(new_n3077_));
  NOR2_X1    g00635(.A1(new_n3062_), .A2(new_n3073_), .ZN(new_n3078_));
  OAI21_X1   g00636(.A1(new_n3078_), .A2(new_n3077_), .B(new_n2436_), .ZN(new_n3079_));
  NAND2_X1   g00637(.A1(new_n3079_), .A2(new_n3076_), .ZN(new_n3080_));
  AOI21_X1   g00638(.A1(new_n3072_), .A2(new_n3080_), .B(new_n3071_), .ZN(new_n3081_));
  INV_X1     g00639(.I(new_n2964_), .ZN(new_n3082_));
  NAND2_X1   g00640(.A1(new_n3062_), .A2(new_n3082_), .ZN(new_n3083_));
  AOI21_X1   g00641(.A1(new_n3052_), .A2(new_n2680_), .B(new_n3050_), .ZN(new_n3084_));
  OAI21_X1   g00642(.A1(new_n3084_), .A2(new_n3049_), .B(new_n3055_), .ZN(new_n3085_));
  MUX2_X1    g00643(.I0(new_n3085_), .I1(new_n2670_), .S(pi0093), .Z(new_n3086_));
  NAND2_X1   g00644(.A1(new_n2676_), .A2(new_n2876_), .ZN(new_n3087_));
  NOR4_X1    g00645(.A1(new_n3086_), .A2(new_n2879_), .A3(new_n3059_), .A4(new_n3087_), .ZN(new_n3088_));
  NOR2_X1    g00646(.A1(new_n3088_), .A2(pi0072), .ZN(new_n3089_));
  INV_X1     g00647(.I(new_n3089_), .ZN(new_n3090_));
  INV_X1     g00648(.I(new_n2860_), .ZN(new_n3091_));
  NOR2_X1    g00649(.A1(new_n3091_), .A2(new_n3082_), .ZN(new_n3092_));
  NOR2_X1    g00650(.A1(new_n2864_), .A2(new_n3092_), .ZN(new_n3093_));
  AOI21_X1   g00651(.A1(new_n3090_), .A2(new_n3093_), .B(new_n3075_), .ZN(new_n3094_));
  AOI21_X1   g00652(.A1(new_n3083_), .A2(new_n3094_), .B(new_n3032_), .ZN(new_n3095_));
  OAI21_X1   g00653(.A1(new_n3095_), .A2(pi0137), .B(new_n3076_), .ZN(new_n3096_));
  NAND2_X1   g00654(.A1(new_n3096_), .A2(new_n2631_), .ZN(new_n3097_));
  NAND2_X1   g00655(.A1(new_n3097_), .A2(pi0146), .ZN(new_n3098_));
  OAI21_X1   g00656(.A1(new_n3098_), .A2(new_n3081_), .B(new_n2985_), .ZN(new_n3099_));
  NAND3_X1   g00657(.A1(new_n2510_), .A2(new_n2438_), .A3(new_n2512_), .ZN(new_n3100_));
  NAND3_X1   g00658(.A1(new_n2668_), .A2(new_n2861_), .A3(new_n2512_), .ZN(new_n3101_));
  NAND2_X1   g00659(.A1(new_n3068_), .A2(new_n3101_), .ZN(new_n3102_));
  NAND2_X1   g00660(.A1(new_n3048_), .A2(new_n3102_), .ZN(new_n3103_));
  AOI21_X1   g00661(.A1(new_n3103_), .A2(new_n3100_), .B(new_n2436_), .ZN(new_n3104_));
  NOR2_X1    g00662(.A1(new_n2668_), .A2(pi0072), .ZN(new_n3105_));
  INV_X1     g00663(.I(new_n3105_), .ZN(new_n3106_));
  NOR3_X1    g00664(.A1(new_n2863_), .A2(new_n2860_), .A3(new_n3106_), .ZN(new_n3107_));
  NAND2_X1   g00665(.A1(new_n3061_), .A2(new_n3107_), .ZN(new_n3108_));
  AOI21_X1   g00666(.A1(new_n3108_), .A2(new_n3047_), .B(new_n3041_), .ZN(new_n3109_));
  NOR2_X1    g00667(.A1(new_n2611_), .A2(pi0210), .ZN(new_n3110_));
  OAI21_X1   g00668(.A1(new_n3109_), .A2(new_n3104_), .B(new_n3110_), .ZN(new_n3111_));
  NOR2_X1    g00669(.A1(new_n3108_), .A2(new_n2964_), .ZN(new_n3112_));
  OR3_X2     g00670(.A1(new_n2863_), .A2(new_n3092_), .A3(new_n3106_), .Z(new_n3113_));
  OAI21_X1   g00671(.A1(new_n3088_), .A2(new_n3113_), .B(new_n3074_), .ZN(new_n3114_));
  OAI21_X1   g00672(.A1(new_n3112_), .A2(new_n3114_), .B(new_n2872_), .ZN(new_n3115_));
  NAND2_X1   g00673(.A1(new_n3100_), .A2(pi0137), .ZN(new_n3116_));
  AOI21_X1   g00674(.A1(new_n3074_), .A2(new_n3102_), .B(new_n3116_), .ZN(new_n3117_));
  NOR2_X1    g00675(.A1(new_n3117_), .A2(pi0137), .ZN(new_n3118_));
  AOI21_X1   g00676(.A1(new_n3115_), .A2(new_n3118_), .B(pi0210), .ZN(new_n3119_));
  OAI21_X1   g00677(.A1(new_n3119_), .A2(new_n3111_), .B(new_n2576_), .ZN(new_n3120_));
  NAND4_X1   g00678(.A1(new_n3120_), .A2(new_n2631_), .A3(new_n3070_), .A4(new_n3096_), .ZN(new_n3121_));
  INV_X1     g00679(.I(new_n3073_), .ZN(new_n3122_));
  NAND2_X1   g00680(.A1(new_n3108_), .A2(new_n3122_), .ZN(new_n3123_));
  AOI21_X1   g00681(.A1(new_n3123_), .A2(new_n2437_), .B(new_n3041_), .ZN(new_n3124_));
  OAI21_X1   g00682(.A1(new_n3124_), .A2(new_n3117_), .B(new_n3072_), .ZN(new_n3125_));
  NAND4_X1   g00683(.A1(new_n3119_), .A2(new_n3125_), .A3(pi0146), .A4(new_n3111_), .ZN(new_n3126_));
  NAND4_X1   g00684(.A1(new_n3099_), .A2(new_n2526_), .A3(new_n3121_), .A4(new_n3126_), .ZN(new_n3127_));
  AOI22_X1   g00685(.A1(new_n3045_), .A2(new_n2527_), .B1(new_n3127_), .B2(new_n2523_), .ZN(new_n3128_));
  OAI21_X1   g00686(.A1(new_n3007_), .A2(new_n3128_), .B(new_n2562_), .ZN(new_n3129_));
  NOR3_X1    g00687(.A1(new_n2560_), .A2(pi0221), .A3(new_n2564_), .ZN(new_n3130_));
  AOI21_X1   g00688(.A1(new_n3129_), .A2(new_n3130_), .B(pi0215), .ZN(new_n3131_));
  NOR2_X1    g00689(.A1(new_n2606_), .A2(pi0223), .ZN(new_n3132_));
  NAND2_X1   g00690(.A1(new_n2989_), .A2(pi0198), .ZN(new_n3133_));
  NAND2_X1   g00691(.A1(new_n2948_), .A2(new_n2601_), .ZN(new_n3134_));
  NAND2_X1   g00692(.A1(new_n3134_), .A2(new_n3133_), .ZN(new_n3135_));
  NAND2_X1   g00693(.A1(new_n2977_), .A2(pi0198), .ZN(new_n3136_));
  OAI21_X1   g00694(.A1(new_n2969_), .A2(pi0198), .B(new_n3136_), .ZN(new_n3137_));
  OAI21_X1   g00695(.A1(pi0234), .A2(new_n3137_), .B(new_n3135_), .ZN(new_n3138_));
  NAND4_X1   g00696(.A1(new_n3134_), .A2(new_n2440_), .A3(new_n3133_), .A4(new_n3137_), .ZN(new_n3139_));
  NAND4_X1   g00697(.A1(new_n3138_), .A2(new_n2563_), .A3(new_n3132_), .A4(new_n3139_), .ZN(new_n3140_));
  NAND3_X1   g00698(.A1(new_n3137_), .A2(pi0142), .A3(new_n2992_), .ZN(new_n3143_));
  NAND3_X1   g00699(.A1(new_n3135_), .A2(pi0142), .A3(new_n2986_), .ZN(new_n3146_));
  NOR2_X1    g00700(.A1(new_n2605_), .A2(pi0223), .ZN(new_n3147_));
  NAND4_X1   g00701(.A1(new_n3140_), .A2(new_n3143_), .A3(new_n3146_), .A4(new_n3147_), .ZN(new_n3148_));
  NAND2_X1   g00702(.A1(new_n2600_), .A2(new_n2587_), .ZN(new_n3149_));
  AOI21_X1   g00703(.A1(new_n3148_), .A2(new_n2614_), .B(new_n3149_), .ZN(new_n3150_));
  NOR2_X1    g00704(.A1(new_n2567_), .A2(new_n2566_), .ZN(new_n3151_));
  NOR2_X1    g00705(.A1(new_n3151_), .A2(new_n2587_), .ZN(new_n3152_));
  OAI21_X1   g00706(.A1(new_n3150_), .A2(pi0039), .B(new_n3152_), .ZN(new_n3153_));
  INV_X1     g00707(.I(pi0039), .ZN(new_n3154_));
  INV_X1     g00708(.I(new_n2614_), .ZN(new_n3155_));
  NOR2_X1    g00709(.A1(new_n3155_), .A2(pi0223), .ZN(new_n3156_));
  NAND2_X1   g00710(.A1(new_n2520_), .A2(new_n3156_), .ZN(new_n3157_));
  AOI21_X1   g00711(.A1(new_n3157_), .A2(new_n2600_), .B(pi0299), .ZN(new_n3158_));
  NAND2_X1   g00712(.A1(new_n2527_), .A2(new_n2522_), .ZN(new_n3159_));
  NAND2_X1   g00713(.A1(new_n2521_), .A2(pi0105), .ZN(new_n3160_));
  AOI21_X1   g00714(.A1(new_n3160_), .A2(new_n3159_), .B(new_n2523_), .ZN(new_n3161_));
  INV_X1     g00715(.I(new_n2516_), .ZN(new_n3162_));
  NOR4_X1    g00716(.A1(new_n3162_), .A2(pi0137), .A3(pi0153), .A4(pi0332), .ZN(new_n3163_));
  INV_X1     g00717(.I(new_n2527_), .ZN(new_n3164_));
  AOI21_X1   g00718(.A1(new_n2490_), .A2(pi0137), .B(new_n3164_), .ZN(new_n3165_));
  OAI21_X1   g00719(.A1(new_n3163_), .A2(new_n3165_), .B(new_n2523_), .ZN(new_n3166_));
  NAND2_X1   g00720(.A1(new_n3166_), .A2(new_n2562_), .ZN(new_n3167_));
  OAI21_X1   g00721(.A1(new_n3161_), .A2(new_n3167_), .B(new_n2573_), .ZN(new_n3168_));
  NAND4_X1   g00722(.A1(new_n3168_), .A2(new_n2550_), .A3(new_n2569_), .A4(new_n2620_), .ZN(new_n3169_));
  AOI21_X1   g00723(.A1(new_n3169_), .A2(pi0299), .B(new_n3158_), .ZN(new_n3170_));
  NOR2_X1    g00724(.A1(new_n3170_), .A2(new_n3154_), .ZN(new_n3171_));
  INV_X1     g00725(.I(pi0038), .ZN(new_n3172_));
  INV_X1     g00726(.I(pi0100), .ZN(new_n3173_));
  NOR3_X1    g00727(.A1(new_n2532_), .A2(pi0299), .A3(new_n2570_), .ZN(new_n3174_));
  NOR3_X1    g00728(.A1(new_n3174_), .A2(pi0039), .A3(new_n3158_), .ZN(new_n3175_));
  OAI21_X1   g00729(.A1(new_n3175_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n3176_));
  INV_X1     g00730(.I(pi0087), .ZN(new_n3177_));
  INV_X1     g00731(.I(new_n2584_), .ZN(new_n3178_));
  OAI21_X1   g00732(.A1(new_n2631_), .A2(pi0252), .B(new_n3025_), .ZN(new_n3179_));
  NAND4_X1   g00733(.A1(new_n2490_), .A2(pi0137), .A3(new_n3164_), .A4(new_n2577_), .ZN(new_n3180_));
  INV_X1     g00734(.I(pi0252), .ZN(new_n3181_));
  OAI21_X1   g00735(.A1(new_n2436_), .A2(pi0210), .B(new_n3181_), .ZN(new_n3182_));
  OAI21_X1   g00736(.A1(new_n2577_), .A2(new_n3182_), .B(new_n2563_), .ZN(new_n3183_));
  NOR2_X1    g00737(.A1(new_n3162_), .A2(new_n3183_), .ZN(new_n3184_));
  AOI22_X1   g00738(.A1(new_n3163_), .A2(new_n3179_), .B1(new_n3180_), .B2(new_n3184_), .ZN(new_n3185_));
  OAI21_X1   g00739(.A1(new_n3185_), .A2(pi0228), .B(new_n2562_), .ZN(new_n3186_));
  NAND2_X1   g00740(.A1(new_n3178_), .A2(new_n3186_), .ZN(new_n3187_));
  AOI21_X1   g00741(.A1(new_n3187_), .A2(new_n2573_), .B(pi0221), .ZN(new_n3188_));
  NOR2_X1    g00742(.A1(new_n2544_), .A2(pi0299), .ZN(new_n3189_));
  NAND4_X1   g00743(.A1(new_n2617_), .A2(new_n2569_), .A3(new_n2620_), .A4(new_n3189_), .ZN(new_n3190_));
  NOR2_X1    g00744(.A1(new_n2545_), .A2(new_n3173_), .ZN(new_n3191_));
  OAI21_X1   g00745(.A1(new_n3188_), .A2(new_n3190_), .B(new_n3191_), .ZN(new_n3192_));
  NAND2_X1   g00746(.A1(new_n3192_), .A2(new_n3177_), .ZN(new_n3193_));
  NAND3_X1   g00747(.A1(new_n3193_), .A2(new_n3176_), .A3(new_n3172_), .ZN(new_n3194_));
  NOR2_X1    g00748(.A1(new_n3171_), .A2(new_n3194_), .ZN(new_n3195_));
  OAI21_X1   g00749(.A1(new_n3153_), .A2(new_n3131_), .B(new_n3195_), .ZN(new_n3196_));
  NOR2_X1    g00750(.A1(new_n2622_), .A2(pi0039), .ZN(new_n3197_));
  INV_X1     g00751(.I(new_n3197_), .ZN(new_n3198_));
  OR2_X2     g00752(.A1(new_n3170_), .A2(new_n3198_), .Z(new_n3199_));
  AOI21_X1   g00753(.A1(new_n3199_), .A2(pi0087), .B(pi0075), .ZN(new_n3200_));
  AOI22_X1   g00754(.A1(new_n3196_), .A2(new_n3200_), .B1(new_n2627_), .B2(new_n2630_), .ZN(new_n3201_));
  INV_X1     g00755(.I(pi0074), .ZN(new_n3202_));
  INV_X1     g00756(.I(pi0092), .ZN(new_n3203_));
  NOR3_X1    g00757(.A1(new_n3199_), .A2(new_n3203_), .A3(new_n2535_), .ZN(new_n3204_));
  NOR2_X1    g00758(.A1(pi0087), .A2(pi0100), .ZN(new_n3205_));
  INV_X1     g00759(.I(new_n3205_), .ZN(new_n3206_));
  NOR2_X1    g00760(.A1(new_n3206_), .A2(pi0038), .ZN(new_n3207_));
  INV_X1     g00761(.I(new_n3207_), .ZN(new_n3208_));
  NOR2_X1    g00762(.A1(pi0075), .A2(pi0092), .ZN(new_n3209_));
  NAND2_X1   g00763(.A1(new_n3209_), .A2(new_n3154_), .ZN(new_n3210_));
  NOR4_X1    g00764(.A1(new_n3174_), .A2(new_n3158_), .A3(new_n3208_), .A4(new_n3210_), .ZN(new_n3211_));
  NOR3_X1    g00765(.A1(new_n3204_), .A2(pi0054), .A3(new_n3202_), .ZN(new_n3212_));
  OAI21_X1   g00766(.A1(new_n3201_), .A2(pi0092), .B(new_n3212_), .ZN(new_n3213_));
  INV_X1     g00767(.I(pi0054), .ZN(new_n3214_));
  NOR2_X1    g00768(.A1(new_n3211_), .A2(new_n3214_), .ZN(new_n3215_));
  AOI21_X1   g00769(.A1(new_n3215_), .A2(new_n3202_), .B(pi0055), .ZN(new_n3216_));
  INV_X1     g00770(.I(new_n2570_), .ZN(new_n3217_));
  NOR2_X1    g00771(.A1(new_n3217_), .A2(new_n2548_), .ZN(new_n3218_));
  AOI21_X1   g00772(.A1(new_n3169_), .A2(new_n2548_), .B(new_n3218_), .ZN(new_n3219_));
  AND2_X2    g00773(.A1(new_n3219_), .A2(pi0056), .Z(new_n3220_));
  OAI21_X1   g00774(.A1(new_n2527_), .A2(pi0105), .B(pi0228), .ZN(new_n3221_));
  NAND3_X1   g00775(.A1(new_n3221_), .A2(new_n2522_), .A3(new_n2563_), .ZN(new_n3222_));
  NOR2_X1    g00776(.A1(new_n3164_), .A2(pi0228), .ZN(new_n3223_));
  AOI21_X1   g00777(.A1(new_n2491_), .A2(new_n3223_), .B(pi0216), .ZN(new_n3224_));
  OAI21_X1   g00778(.A1(new_n2518_), .A2(new_n3222_), .B(new_n3224_), .ZN(new_n3225_));
  AOI21_X1   g00779(.A1(new_n3225_), .A2(new_n2573_), .B(new_n2550_), .ZN(new_n3226_));
  INV_X1     g00780(.I(pi0055), .ZN(new_n3227_));
  INV_X1     g00781(.I(new_n3209_), .ZN(new_n3228_));
  NOR2_X1    g00782(.A1(new_n2539_), .A2(new_n3228_), .ZN(new_n3229_));
  INV_X1     g00783(.I(new_n3229_), .ZN(new_n3230_));
  NOR2_X1    g00784(.A1(new_n3230_), .A2(new_n3206_), .ZN(new_n3231_));
  INV_X1     g00785(.I(new_n3231_), .ZN(new_n3232_));
  NOR2_X1    g00786(.A1(new_n3232_), .A2(new_n2545_), .ZN(new_n3233_));
  INV_X1     g00787(.I(new_n3233_), .ZN(new_n3234_));
  AOI21_X1   g00788(.A1(new_n3217_), .A2(new_n3234_), .B(new_n3227_), .ZN(new_n3235_));
  OR3_X2     g00789(.A1(new_n3234_), .A2(pi0215), .A3(new_n3151_), .Z(new_n3236_));
  NOR4_X1    g00790(.A1(new_n3226_), .A2(new_n2559_), .A3(new_n3235_), .A4(new_n3236_), .ZN(new_n3237_));
  OAI22_X1   g00791(.A1(new_n3220_), .A2(pi0062), .B1(pi0056), .B2(new_n3237_), .ZN(new_n3238_));
  AOI21_X1   g00792(.A1(new_n3213_), .A2(new_n3216_), .B(new_n3238_), .ZN(new_n3239_));
  INV_X1     g00793(.I(pi0062), .ZN(new_n3240_));
  MUX2_X1    g00794(.I0(new_n3219_), .I1(new_n3217_), .S(pi0056), .Z(new_n3241_));
  NOR2_X1    g00795(.A1(pi0057), .A2(pi0059), .ZN(new_n3242_));
  OAI21_X1   g00796(.A1(new_n3241_), .A2(new_n3240_), .B(new_n3242_), .ZN(new_n3243_));
  OAI21_X1   g00797(.A1(new_n3239_), .A2(new_n3243_), .B(new_n2572_), .ZN(po0153));
  NOR2_X1    g00798(.A1(new_n2491_), .A2(pi0252), .ZN(new_n3245_));
  NOR2_X1    g00799(.A1(pi0161), .A2(pi0166), .ZN(new_n3246_));
  INV_X1     g00800(.I(new_n3246_), .ZN(new_n3247_));
  NOR3_X1    g00801(.A1(new_n2491_), .A2(pi0146), .A3(new_n3181_), .ZN(new_n3248_));
  NAND2_X1   g00802(.A1(new_n3248_), .A2(new_n3247_), .ZN(new_n3249_));
  INV_X1     g00803(.I(pi0152), .ZN(new_n3250_));
  OAI21_X1   g00804(.A1(new_n3249_), .A2(new_n3245_), .B(new_n3250_), .ZN(new_n3251_));
  AOI21_X1   g00805(.A1(new_n3245_), .A2(new_n3249_), .B(new_n3251_), .ZN(new_n3252_));
  AOI21_X1   g00806(.A1(pi0146), .A2(pi0252), .B(new_n2491_), .ZN(new_n3253_));
  NOR2_X1    g00807(.A1(new_n3253_), .A2(new_n3250_), .ZN(new_n3254_));
  INV_X1     g00808(.I(new_n3254_), .ZN(new_n3255_));
  NAND2_X1   g00809(.A1(new_n3252_), .A2(new_n3255_), .ZN(new_n3256_));
  INV_X1     g00810(.I(new_n3256_), .ZN(new_n3257_));
  INV_X1     g00811(.I(pi1146), .ZN(new_n3258_));
  NOR2_X1    g00812(.A1(new_n2566_), .A2(new_n3258_), .ZN(new_n3259_));
  INV_X1     g00813(.I(new_n3259_), .ZN(new_n3260_));
  INV_X1     g00814(.I(pi0939), .ZN(new_n3261_));
  NOR3_X1    g00815(.A1(new_n2555_), .A2(new_n3261_), .A3(pi1146), .ZN(new_n3262_));
  AOI21_X1   g00816(.A1(new_n2554_), .A2(new_n3261_), .B(new_n3258_), .ZN(new_n3263_));
  OAI21_X1   g00817(.A1(new_n3262_), .A2(new_n3263_), .B(pi0221), .ZN(new_n3264_));
  NAND2_X1   g00818(.A1(new_n3264_), .A2(new_n3260_), .ZN(new_n3265_));
  INV_X1     g00819(.I(new_n3265_), .ZN(new_n3266_));
  NAND2_X1   g00820(.A1(new_n3172_), .A2(new_n2562_), .ZN(new_n3267_));
  NOR2_X1    g00821(.A1(new_n3267_), .A2(pi0228), .ZN(new_n3268_));
  NOR3_X1    g00822(.A1(new_n2587_), .A2(pi0039), .A3(pi0154), .ZN(new_n3269_));
  NAND4_X1   g00823(.A1(new_n3257_), .A2(new_n3266_), .A3(new_n3268_), .A4(new_n3269_), .ZN(new_n3270_));
  INV_X1     g00824(.I(pi0154), .ZN(new_n3271_));
  INV_X1     g00825(.I(pi0276), .ZN(new_n3272_));
  NOR3_X1    g00826(.A1(new_n2525_), .A2(pi0216), .A3(new_n3272_), .ZN(new_n3273_));
  AOI21_X1   g00827(.A1(new_n2525_), .A2(new_n2562_), .B(pi0276), .ZN(new_n3274_));
  NOR3_X1    g00828(.A1(new_n3273_), .A2(new_n3274_), .A3(pi0221), .ZN(new_n3275_));
  AOI21_X1   g00829(.A1(new_n3275_), .A2(new_n3264_), .B(pi0215), .ZN(new_n3276_));
  NOR2_X1    g00830(.A1(new_n3276_), .A2(new_n3259_), .ZN(new_n3277_));
  NOR2_X1    g00831(.A1(new_n2562_), .A2(pi0221), .ZN(new_n3278_));
  NAND2_X1   g00832(.A1(new_n3278_), .A2(pi0276), .ZN(new_n3279_));
  AOI21_X1   g00833(.A1(new_n3264_), .A2(new_n3279_), .B(pi0215), .ZN(new_n3280_));
  AOI21_X1   g00834(.A1(pi0215), .A2(new_n3258_), .B(new_n3280_), .ZN(new_n3281_));
  NOR2_X1    g00835(.A1(new_n2525_), .A2(new_n2974_), .ZN(new_n3282_));
  INV_X1     g00836(.I(new_n3282_), .ZN(new_n3283_));
  NOR2_X1    g00837(.A1(pi0216), .A2(pi0221), .ZN(new_n3284_));
  INV_X1     g00838(.I(new_n3284_), .ZN(new_n3285_));
  NOR2_X1    g00839(.A1(new_n3285_), .A2(pi0215), .ZN(new_n3286_));
  INV_X1     g00840(.I(new_n3286_), .ZN(new_n3287_));
  NOR2_X1    g00841(.A1(new_n3283_), .A2(new_n3287_), .ZN(new_n3288_));
  NOR2_X1    g00842(.A1(new_n3281_), .A2(new_n3288_), .ZN(new_n3289_));
  AOI21_X1   g00843(.A1(pi0154), .A2(new_n2566_), .B(new_n3289_), .ZN(new_n3290_));
  AOI21_X1   g00844(.A1(new_n3271_), .A2(new_n3277_), .B(new_n3290_), .ZN(new_n3291_));
  INV_X1     g00845(.I(new_n3291_), .ZN(new_n3292_));
  NOR2_X1    g00846(.A1(pi0223), .A2(pi0299), .ZN(new_n3293_));
  INV_X1     g00847(.I(new_n3293_), .ZN(new_n3294_));
  NOR2_X1    g00848(.A1(new_n3155_), .A2(new_n3294_), .ZN(new_n3295_));
  INV_X1     g00849(.I(new_n3295_), .ZN(new_n3296_));
  NOR2_X1    g00850(.A1(new_n3296_), .A2(new_n2974_), .ZN(new_n3297_));
  MUX2_X1    g00851(.I0(pi1146), .I1(pi0939), .S(new_n2589_), .Z(new_n3298_));
  NOR2_X1    g00852(.A1(new_n2595_), .A2(pi0222), .ZN(new_n3299_));
  INV_X1     g00853(.I(new_n3299_), .ZN(new_n3300_));
  NOR2_X1    g00854(.A1(pi0223), .A2(pi0299), .ZN(new_n3301_));
  OAI21_X1   g00855(.A1(new_n3300_), .A2(new_n3272_), .B(new_n3301_), .ZN(new_n3302_));
  AOI21_X1   g00856(.A1(new_n3298_), .A2(pi0222), .B(new_n3302_), .ZN(new_n3303_));
  INV_X1     g00857(.I(new_n3303_), .ZN(new_n3304_));
  NOR2_X1    g00858(.A1(new_n3304_), .A2(new_n3297_), .ZN(new_n3305_));
  OAI21_X1   g00859(.A1(new_n3292_), .A2(pi0299), .B(new_n3305_), .ZN(new_n3306_));
  OAI21_X1   g00860(.A1(new_n3306_), .A2(new_n2621_), .B(pi0100), .ZN(new_n3307_));
  NOR2_X1    g00861(.A1(new_n3270_), .A2(new_n3307_), .ZN(new_n3308_));
  INV_X1     g00862(.I(new_n3306_), .ZN(new_n3309_));
  NOR2_X1    g00863(.A1(new_n2491_), .A2(pi0228), .ZN(new_n3310_));
  INV_X1     g00864(.I(new_n3310_), .ZN(new_n3311_));
  NOR3_X1    g00865(.A1(new_n3311_), .A2(pi0216), .A3(new_n3265_), .ZN(new_n3312_));
  OAI21_X1   g00866(.A1(new_n3271_), .A2(new_n3289_), .B(new_n3312_), .ZN(new_n3313_));
  NAND2_X1   g00867(.A1(new_n3292_), .A2(new_n3313_), .ZN(new_n3314_));
  INV_X1     g00868(.I(new_n3314_), .ZN(new_n3315_));
  NOR2_X1    g00869(.A1(new_n3315_), .A2(new_n2587_), .ZN(new_n3316_));
  NAND4_X1   g00870(.A1(new_n3316_), .A2(new_n3177_), .A3(new_n3197_), .A4(new_n3309_), .ZN(new_n3317_));
  NAND2_X1   g00871(.A1(new_n3317_), .A2(new_n2628_), .ZN(new_n3318_));
  NOR2_X1    g00872(.A1(new_n2621_), .A2(new_n3154_), .ZN(new_n3319_));
  OAI21_X1   g00873(.A1(new_n3316_), .A2(new_n3306_), .B(new_n3319_), .ZN(new_n3320_));
  NAND3_X1   g00874(.A1(new_n3318_), .A2(new_n3177_), .A3(new_n3320_), .ZN(new_n3321_));
  NOR2_X1    g00875(.A1(new_n2547_), .A2(new_n2535_), .ZN(new_n3322_));
  INV_X1     g00876(.I(new_n3322_), .ZN(new_n3323_));
  NOR2_X1    g00877(.A1(new_n3323_), .A2(pi0092), .ZN(new_n3324_));
  INV_X1     g00878(.I(new_n3324_), .ZN(new_n3325_));
  NOR4_X1    g00879(.A1(new_n3315_), .A2(new_n2587_), .A3(new_n3306_), .A4(new_n3325_), .ZN(new_n3326_));
  AOI21_X1   g00880(.A1(new_n3306_), .A2(new_n2539_), .B(pi0055), .ZN(new_n3327_));
  NOR2_X1    g00881(.A1(new_n3309_), .A2(new_n2628_), .ZN(new_n3328_));
  NOR2_X1    g00882(.A1(new_n2539_), .A2(pi0092), .ZN(new_n3329_));
  INV_X1     g00883(.I(new_n3329_), .ZN(new_n3330_));
  NOR4_X1    g00884(.A1(new_n3326_), .A2(new_n3328_), .A3(new_n3327_), .A4(new_n3330_), .ZN(new_n3331_));
  OAI21_X1   g00885(.A1(new_n3321_), .A2(new_n3308_), .B(new_n3331_), .ZN(new_n3332_));
  NOR2_X1    g00886(.A1(new_n3234_), .A2(pi0055), .ZN(new_n3333_));
  NAND2_X1   g00887(.A1(new_n3315_), .A2(new_n3333_), .ZN(new_n3334_));
  INV_X1     g00888(.I(pi0056), .ZN(new_n3335_));
  INV_X1     g00889(.I(new_n2548_), .ZN(new_n3336_));
  AOI21_X1   g00890(.A1(new_n3292_), .A2(new_n3336_), .B(new_n3335_), .ZN(new_n3337_));
  NAND2_X1   g00891(.A1(new_n3292_), .A2(new_n3333_), .ZN(new_n3338_));
  OAI21_X1   g00892(.A1(new_n3338_), .A2(new_n3313_), .B(new_n2533_), .ZN(new_n3339_));
  AOI21_X1   g00893(.A1(new_n3334_), .A2(new_n3337_), .B(new_n3339_), .ZN(new_n3340_));
  NOR2_X1    g00894(.A1(new_n2543_), .A2(pi0056), .ZN(new_n3341_));
  INV_X1     g00895(.I(new_n3341_), .ZN(new_n3342_));
  NOR2_X1    g00896(.A1(new_n3342_), .A2(new_n2547_), .ZN(new_n3343_));
  NOR4_X1    g00897(.A1(new_n3334_), .A2(pi0056), .A3(new_n3291_), .A4(new_n3343_), .ZN(new_n3344_));
  OAI21_X1   g00898(.A1(new_n3344_), .A2(new_n3240_), .B(new_n2571_), .ZN(new_n3345_));
  AOI21_X1   g00899(.A1(new_n3332_), .A2(new_n3340_), .B(new_n3345_), .ZN(new_n3346_));
  OAI21_X1   g00900(.A1(new_n3292_), .A2(new_n2571_), .B(pi0239), .ZN(new_n3347_));
  INV_X1     g00901(.I(new_n3312_), .ZN(new_n3348_));
  NOR3_X1    g00902(.A1(new_n3276_), .A2(new_n2587_), .A3(new_n3259_), .ZN(new_n3349_));
  NAND2_X1   g00903(.A1(new_n3348_), .A2(new_n3349_), .ZN(new_n3350_));
  NAND2_X1   g00904(.A1(new_n3350_), .A2(new_n3303_), .ZN(new_n3351_));
  NAND2_X1   g00905(.A1(new_n3281_), .A2(pi0299), .ZN(new_n3352_));
  NAND2_X1   g00906(.A1(new_n3352_), .A2(new_n3303_), .ZN(new_n3353_));
  NAND2_X1   g00907(.A1(new_n3353_), .A2(pi0154), .ZN(new_n3354_));
  NAND2_X1   g00908(.A1(new_n3354_), .A2(new_n3197_), .ZN(new_n3355_));
  AOI21_X1   g00909(.A1(new_n3351_), .A2(new_n3271_), .B(new_n3355_), .ZN(new_n3356_));
  NOR2_X1    g00910(.A1(new_n3277_), .A2(pi0154), .ZN(new_n3357_));
  NOR2_X1    g00911(.A1(new_n3281_), .A2(new_n3271_), .ZN(new_n3358_));
  NOR2_X1    g00912(.A1(new_n3358_), .A2(new_n3357_), .ZN(new_n3359_));
  AOI21_X1   g00913(.A1(new_n3359_), .A2(pi0299), .B(new_n3304_), .ZN(new_n3360_));
  AOI21_X1   g00914(.A1(new_n3360_), .A2(new_n3323_), .B(new_n2537_), .ZN(new_n3361_));
  NAND2_X1   g00915(.A1(new_n3356_), .A2(new_n3361_), .ZN(new_n3362_));
  INV_X1     g00916(.I(new_n2655_), .ZN(new_n3363_));
  INV_X1     g00917(.I(pi0040), .ZN(new_n3364_));
  NOR2_X1    g00918(.A1(new_n2510_), .A2(new_n3364_), .ZN(new_n3365_));
  AOI21_X1   g00919(.A1(new_n3363_), .A2(pi0032), .B(new_n3365_), .ZN(new_n3366_));
  INV_X1     g00920(.I(new_n3366_), .ZN(new_n3367_));
  INV_X1     g00921(.I(new_n2862_), .ZN(new_n3368_));
  NOR2_X1    g00922(.A1(new_n3012_), .A2(pi0070), .ZN(new_n3369_));
  OAI21_X1   g00923(.A1(new_n2876_), .A2(new_n2851_), .B(new_n3060_), .ZN(new_n3370_));
  OAI21_X1   g00924(.A1(new_n3369_), .A2(new_n3370_), .B(new_n2658_), .ZN(new_n3371_));
  NAND2_X1   g00925(.A1(new_n3371_), .A2(new_n2675_), .ZN(new_n3372_));
  NAND2_X1   g00926(.A1(new_n3372_), .A2(new_n3105_), .ZN(new_n3373_));
  AOI21_X1   g00927(.A1(new_n3373_), .A2(new_n3368_), .B(new_n2513_), .ZN(new_n3374_));
  OAI21_X1   g00928(.A1(new_n3374_), .A2(new_n3367_), .B(new_n2437_), .ZN(new_n3375_));
  NAND2_X1   g00929(.A1(new_n3375_), .A2(new_n2872_), .ZN(new_n3376_));
  INV_X1     g00930(.I(new_n3376_), .ZN(new_n3377_));
  NOR2_X1    g00931(.A1(new_n2491_), .A2(new_n3154_), .ZN(new_n3378_));
  AOI21_X1   g00932(.A1(new_n3377_), .A2(new_n3154_), .B(new_n3378_), .ZN(new_n3379_));
  INV_X1     g00933(.I(new_n3360_), .ZN(new_n3386_));
  NAND3_X1   g00934(.A1(new_n3360_), .A2(pi0075), .A3(pi0092), .ZN(new_n3391_));
  OAI21_X1   g00935(.A1(new_n3386_), .A2(new_n2538_), .B(new_n3227_), .ZN(new_n3392_));
  OAI21_X1   g00936(.A1(new_n3281_), .A2(pi0154), .B(new_n3233_), .ZN(new_n3393_));
  OAI21_X1   g00937(.A1(new_n3348_), .A2(new_n3393_), .B(new_n3359_), .ZN(new_n3394_));
  NAND2_X1   g00938(.A1(new_n3394_), .A2(new_n3227_), .ZN(new_n3395_));
  NAND4_X1   g00939(.A1(new_n3395_), .A2(new_n3335_), .A3(new_n2539_), .A4(new_n3392_), .ZN(new_n3396_));
  AOI21_X1   g00940(.A1(new_n3362_), .A2(new_n3391_), .B(new_n3396_), .ZN(new_n3397_));
  NAND2_X1   g00941(.A1(new_n3359_), .A2(new_n3333_), .ZN(new_n3398_));
  NAND4_X1   g00942(.A1(new_n3348_), .A2(pi0154), .A3(new_n3281_), .A4(new_n3398_), .ZN(new_n3399_));
  INV_X1     g00943(.I(new_n3343_), .ZN(new_n3400_));
  AOI21_X1   g00944(.A1(new_n3400_), .A2(new_n3359_), .B(pi0062), .ZN(new_n3401_));
  NAND2_X1   g00945(.A1(new_n3399_), .A2(new_n3401_), .ZN(new_n3402_));
  AOI21_X1   g00946(.A1(new_n3359_), .A2(new_n3336_), .B(new_n3335_), .ZN(new_n3403_));
  NAND2_X1   g00947(.A1(new_n3399_), .A2(new_n3403_), .ZN(new_n3404_));
  INV_X1     g00948(.I(new_n2571_), .ZN(new_n3405_));
  NOR2_X1    g00949(.A1(new_n3405_), .A2(pi0062), .ZN(new_n3406_));
  NAND3_X1   g00950(.A1(new_n3402_), .A2(new_n3404_), .A3(new_n3406_), .ZN(new_n3407_));
  NOR2_X1    g00951(.A1(new_n3397_), .A2(new_n3407_), .ZN(new_n3408_));
  INV_X1     g00952(.I(pi0239), .ZN(new_n3409_));
  OAI21_X1   g00953(.A1(new_n3359_), .A2(new_n2571_), .B(new_n3409_), .ZN(new_n3410_));
  OAI22_X1   g00954(.A1(new_n3346_), .A2(new_n3347_), .B1(new_n3408_), .B2(new_n3410_), .ZN(po0154));
  INV_X1     g00955(.I(pi0927), .ZN(new_n3412_));
  NOR3_X1    g00956(.A1(new_n2555_), .A2(new_n3412_), .A3(pi1145), .ZN(new_n3413_));
  INV_X1     g00957(.I(pi1145), .ZN(new_n3414_));
  AOI21_X1   g00958(.A1(new_n2554_), .A2(new_n3412_), .B(new_n3414_), .ZN(new_n3415_));
  OAI21_X1   g00959(.A1(new_n3413_), .A2(new_n3415_), .B(pi0221), .ZN(new_n3416_));
  INV_X1     g00960(.I(pi0151), .ZN(new_n3417_));
  INV_X1     g00961(.I(new_n2485_), .ZN(new_n3418_));
  NAND2_X1   g00962(.A1(new_n2668_), .A2(new_n3418_), .ZN(new_n3419_));
  INV_X1     g00963(.I(new_n3419_), .ZN(new_n3420_));
  NOR2_X1    g00964(.A1(new_n3420_), .A2(new_n2438_), .ZN(new_n3421_));
  INV_X1     g00965(.I(new_n3421_), .ZN(new_n3422_));
  NOR2_X1    g00966(.A1(new_n3422_), .A2(new_n2522_), .ZN(new_n3423_));
  NAND4_X1   g00967(.A1(new_n3372_), .A2(pi0072), .A3(new_n2513_), .A4(new_n2654_), .ZN(new_n3424_));
  AOI21_X1   g00968(.A1(new_n3424_), .A2(new_n3366_), .B(pi0095), .ZN(new_n3425_));
  NOR2_X1    g00969(.A1(new_n3425_), .A2(new_n3032_), .ZN(new_n3426_));
  MUX2_X1    g00970(.I0(new_n3426_), .I1(new_n3423_), .S(pi0228), .Z(new_n3427_));
  NOR2_X1    g00971(.A1(new_n3421_), .A2(new_n2871_), .ZN(new_n3428_));
  NOR2_X1    g00972(.A1(new_n3421_), .A2(new_n2522_), .ZN(new_n3429_));
  INV_X1     g00973(.I(new_n3429_), .ZN(new_n3430_));
  NOR2_X1    g00974(.A1(new_n3430_), .A2(new_n2523_), .ZN(new_n3431_));
  AOI21_X1   g00975(.A1(new_n2523_), .A2(new_n3428_), .B(new_n3431_), .ZN(new_n3432_));
  NOR2_X1    g00976(.A1(new_n3432_), .A2(new_n3417_), .ZN(new_n3433_));
  INV_X1     g00977(.I(pi0274), .ZN(new_n3434_));
  NOR2_X1    g00978(.A1(new_n2562_), .A2(new_n3434_), .ZN(new_n3435_));
  NOR2_X1    g00979(.A1(new_n3435_), .A2(pi0221), .ZN(new_n3436_));
  INV_X1     g00980(.I(new_n3436_), .ZN(new_n3437_));
  NOR3_X1    g00981(.A1(new_n3433_), .A2(pi0216), .A3(new_n3437_), .ZN(new_n3438_));
  OAI21_X1   g00982(.A1(new_n3427_), .A2(new_n3417_), .B(new_n3438_), .ZN(new_n3439_));
  NAND2_X1   g00983(.A1(new_n3439_), .A2(new_n3416_), .ZN(new_n3440_));
  MUX2_X1    g00984(.I0(new_n3440_), .I1(pi1145), .S(pi0215), .Z(new_n3441_));
  NOR2_X1    g00985(.A1(new_n3441_), .A2(new_n2587_), .ZN(new_n3442_));
  XNOR2_X1   g00986(.A1(pi0927), .A2(pi1145), .ZN(new_n3444_));
  NOR2_X1    g00987(.A1(new_n3444_), .A2(new_n2593_), .ZN(new_n3445_));
  NAND3_X1   g00988(.A1(pi0223), .A2(pi0299), .A3(pi1145), .ZN(new_n3447_));
  NAND2_X1   g00989(.A1(new_n3447_), .A2(new_n3154_), .ZN(new_n3448_));
  NAND2_X1   g00990(.A1(new_n3445_), .A2(new_n3414_), .ZN(new_n3449_));
  OAI21_X1   g00991(.A1(new_n2593_), .A2(pi0927), .B(pi1145), .ZN(new_n3450_));
  NAND2_X1   g00992(.A1(new_n3449_), .A2(new_n3450_), .ZN(new_n3451_));
  NAND2_X1   g00993(.A1(new_n2588_), .A2(new_n3434_), .ZN(new_n3452_));
  AOI22_X1   g00994(.A1(new_n3451_), .A2(pi0222), .B1(new_n2595_), .B2(new_n3452_), .ZN(new_n3453_));
  NOR3_X1    g00995(.A1(new_n3453_), .A2(pi0223), .A3(new_n3414_), .ZN(new_n3454_));
  AOI21_X1   g00996(.A1(new_n3453_), .A2(new_n2604_), .B(pi1145), .ZN(new_n3455_));
  NOR3_X1    g00997(.A1(new_n3454_), .A2(new_n3455_), .A3(pi0299), .ZN(new_n3456_));
  INV_X1     g00998(.I(new_n3456_), .ZN(new_n3457_));
  NOR2_X1    g00999(.A1(new_n3457_), .A2(new_n3297_), .ZN(new_n3458_));
  NOR2_X1    g01000(.A1(new_n2566_), .A2(new_n3414_), .ZN(new_n3459_));
  NAND2_X1   g01001(.A1(new_n3310_), .A2(new_n3417_), .ZN(new_n3460_));
  NOR2_X1    g01002(.A1(new_n2525_), .A2(new_n2438_), .ZN(new_n3461_));
  AOI21_X1   g01003(.A1(pi0151), .A2(new_n2525_), .B(new_n3461_), .ZN(new_n3462_));
  AOI21_X1   g01004(.A1(new_n3460_), .A2(new_n3462_), .B(pi0216), .ZN(new_n3463_));
  OAI21_X1   g01005(.A1(new_n3463_), .A2(new_n3437_), .B(new_n3416_), .ZN(new_n3464_));
  AOI21_X1   g01006(.A1(new_n3464_), .A2(new_n2566_), .B(new_n3459_), .ZN(new_n3465_));
  INV_X1     g01007(.I(new_n3465_), .ZN(new_n3466_));
  OAI21_X1   g01008(.A1(new_n3466_), .A2(new_n2587_), .B(new_n3458_), .ZN(new_n3467_));
  AOI21_X1   g01009(.A1(new_n3467_), .A2(pi0039), .B(pi0038), .ZN(new_n3468_));
  OAI21_X1   g01010(.A1(new_n3442_), .A2(new_n3448_), .B(new_n3468_), .ZN(new_n3469_));
  NOR2_X1    g01011(.A1(new_n3256_), .A2(pi0228), .ZN(new_n3470_));
  NOR2_X1    g01012(.A1(new_n3470_), .A2(new_n3461_), .ZN(new_n3471_));
  INV_X1     g01013(.I(new_n3471_), .ZN(new_n3472_));
  OR3_X2     g01014(.A1(new_n3463_), .A2(pi0151), .A3(new_n3436_), .Z(new_n3473_));
  OAI21_X1   g01015(.A1(new_n3472_), .A2(new_n3473_), .B(new_n3416_), .ZN(new_n3474_));
  AOI21_X1   g01016(.A1(new_n3474_), .A2(new_n2566_), .B(new_n3459_), .ZN(new_n3475_));
  INV_X1     g01017(.I(new_n3458_), .ZN(new_n3476_));
  NOR2_X1    g01018(.A1(new_n3476_), .A2(new_n2545_), .ZN(new_n3477_));
  OAI21_X1   g01019(.A1(new_n3475_), .A2(pi0299), .B(new_n3477_), .ZN(new_n3478_));
  INV_X1     g01020(.I(new_n3435_), .ZN(new_n3479_));
  NOR2_X1    g01021(.A1(new_n2550_), .A2(pi0216), .ZN(new_n3480_));
  OAI21_X1   g01022(.A1(new_n2524_), .A2(pi0151), .B(new_n3480_), .ZN(new_n3481_));
  AOI21_X1   g01023(.A1(new_n3416_), .A2(new_n3481_), .B(pi0215), .ZN(new_n3482_));
  NOR2_X1    g01024(.A1(new_n3482_), .A2(new_n3459_), .ZN(new_n3483_));
  INV_X1     g01025(.I(new_n3483_), .ZN(new_n3484_));
  NOR2_X1    g01026(.A1(new_n3283_), .A2(new_n2531_), .ZN(new_n3485_));
  NOR3_X1    g01027(.A1(new_n3484_), .A2(new_n3479_), .A3(new_n3485_), .ZN(new_n3486_));
  INV_X1     g01028(.I(new_n3486_), .ZN(new_n3487_));
  AOI21_X1   g01029(.A1(pi0299), .A2(new_n3487_), .B(new_n3476_), .ZN(new_n3488_));
  AOI21_X1   g01030(.A1(new_n3488_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n3489_));
  INV_X1     g01031(.I(new_n3488_), .ZN(new_n3490_));
  OAI21_X1   g01032(.A1(new_n3490_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n3491_));
  AOI21_X1   g01033(.A1(new_n3478_), .A2(new_n3489_), .B(new_n3491_), .ZN(new_n3492_));
  AOI21_X1   g01034(.A1(new_n3469_), .A2(new_n3492_), .B(pi0087), .ZN(new_n3493_));
  NOR2_X1    g01035(.A1(new_n3488_), .A2(new_n3197_), .ZN(new_n3494_));
  AOI21_X1   g01036(.A1(new_n3467_), .A2(new_n3197_), .B(new_n3494_), .ZN(new_n3495_));
  NOR2_X1    g01037(.A1(new_n3495_), .A2(new_n3177_), .ZN(new_n3496_));
  OAI21_X1   g01038(.A1(new_n3493_), .A2(pi0075), .B(new_n3496_), .ZN(new_n3497_));
  NOR4_X1    g01039(.A1(new_n3495_), .A2(pi0092), .A3(new_n2535_), .A4(new_n3488_), .ZN(new_n3498_));
  AOI21_X1   g01040(.A1(new_n3488_), .A2(new_n2539_), .B(pi0055), .ZN(new_n3499_));
  NOR2_X1    g01041(.A1(new_n3490_), .A2(new_n2628_), .ZN(new_n3500_));
  NOR4_X1    g01042(.A1(new_n3498_), .A2(new_n3330_), .A3(new_n3499_), .A4(new_n3500_), .ZN(new_n3501_));
  MUX2_X1    g01043(.I0(new_n3465_), .I1(new_n3487_), .S(new_n3336_), .Z(new_n3502_));
  INV_X1     g01044(.I(new_n2533_), .ZN(new_n3503_));
  NAND2_X1   g01045(.A1(new_n3465_), .A2(new_n3233_), .ZN(new_n3504_));
  AOI21_X1   g01046(.A1(new_n3487_), .A2(new_n3234_), .B(pi0055), .ZN(new_n3505_));
  AOI21_X1   g01047(.A1(new_n3504_), .A2(new_n3505_), .B(new_n3503_), .ZN(new_n3506_));
  OAI21_X1   g01048(.A1(new_n3335_), .A2(new_n3502_), .B(new_n3506_), .ZN(new_n3507_));
  AOI21_X1   g01049(.A1(new_n3497_), .A2(new_n3501_), .B(new_n3507_), .ZN(new_n3508_));
  NOR2_X1    g01050(.A1(new_n3466_), .A2(new_n3400_), .ZN(new_n3509_));
  OAI21_X1   g01051(.A1(new_n3343_), .A2(new_n3486_), .B(new_n3240_), .ZN(new_n3510_));
  INV_X1     g01052(.I(pi0235), .ZN(new_n3511_));
  NOR2_X1    g01053(.A1(new_n3405_), .A2(new_n3511_), .ZN(new_n3512_));
  OAI21_X1   g01054(.A1(new_n3509_), .A2(new_n3510_), .B(new_n3512_), .ZN(new_n3513_));
  NOR2_X1    g01055(.A1(new_n3435_), .A2(new_n3511_), .ZN(new_n3514_));
  AOI21_X1   g01056(.A1(new_n3485_), .A2(new_n3514_), .B(new_n2571_), .ZN(new_n3515_));
  OAI21_X1   g01057(.A1(new_n2566_), .A2(new_n3414_), .B(new_n3416_), .ZN(new_n3516_));
  NOR3_X1    g01058(.A1(new_n3311_), .A2(pi0216), .A3(new_n3516_), .ZN(new_n3517_));
  INV_X1     g01059(.I(new_n3517_), .ZN(new_n3518_));
  NOR2_X1    g01060(.A1(new_n3484_), .A2(new_n2587_), .ZN(new_n3519_));
  NOR4_X1    g01061(.A1(new_n3518_), .A2(new_n2546_), .A3(new_n3457_), .A4(new_n3519_), .ZN(new_n3520_));
  NOR2_X1    g01062(.A1(new_n3457_), .A2(new_n3519_), .ZN(new_n3521_));
  AOI21_X1   g01063(.A1(new_n3521_), .A2(new_n3323_), .B(new_n2537_), .ZN(new_n3522_));
  INV_X1     g01064(.I(new_n3521_), .ZN(new_n3523_));
  INV_X1     g01065(.I(new_n3379_), .ZN(new_n3524_));
  NOR3_X1    g01066(.A1(new_n3523_), .A2(new_n2628_), .A3(new_n3203_), .ZN(new_n3533_));
  AOI21_X1   g01067(.A1(new_n3522_), .A2(new_n3520_), .B(new_n3533_), .ZN(new_n3534_));
  OAI21_X1   g01068(.A1(new_n3521_), .A2(pi0055), .B(new_n2539_), .ZN(new_n3535_));
  NOR3_X1    g01069(.A1(new_n3484_), .A2(pi0055), .A3(new_n3234_), .ZN(new_n3536_));
  AOI21_X1   g01070(.A1(new_n3517_), .A2(new_n3536_), .B(pi0056), .ZN(new_n3537_));
  OAI21_X1   g01071(.A1(new_n3534_), .A2(new_n3535_), .B(new_n3537_), .ZN(new_n3538_));
  NOR2_X1    g01072(.A1(new_n3518_), .A2(new_n3336_), .ZN(new_n3539_));
  NAND3_X1   g01073(.A1(new_n3539_), .A2(new_n2533_), .A3(new_n3483_), .ZN(new_n3540_));
  NOR2_X1    g01074(.A1(new_n3405_), .A2(pi0235), .ZN(new_n3541_));
  INV_X1     g01075(.I(new_n3539_), .ZN(new_n3542_));
  NAND2_X1   g01076(.A1(new_n3542_), .A2(new_n3483_), .ZN(new_n3543_));
  NAND2_X1   g01077(.A1(new_n3543_), .A2(pi0056), .ZN(new_n3544_));
  AOI22_X1   g01078(.A1(new_n3544_), .A2(new_n3240_), .B1(new_n3540_), .B2(new_n3541_), .ZN(new_n3545_));
  AOI22_X1   g01079(.A1(new_n3545_), .A2(new_n3538_), .B1(new_n3484_), .B2(new_n3515_), .ZN(new_n3546_));
  OAI21_X1   g01080(.A1(new_n3508_), .A2(new_n3513_), .B(new_n3546_), .ZN(po0155));
  INV_X1     g01081(.I(pi1143), .ZN(new_n3548_));
  INV_X1     g01082(.I(pi0944), .ZN(new_n3549_));
  NOR3_X1    g01083(.A1(new_n2555_), .A2(new_n3549_), .A3(pi1143), .ZN(new_n3550_));
  AOI21_X1   g01084(.A1(new_n2554_), .A2(new_n3549_), .B(new_n3548_), .ZN(new_n3551_));
  OAI21_X1   g01085(.A1(new_n3550_), .A2(new_n3551_), .B(pi0221), .ZN(new_n3552_));
  NAND2_X1   g01086(.A1(pi0216), .A2(pi0264), .ZN(new_n3553_));
  NAND2_X1   g01087(.A1(new_n3553_), .A2(new_n2550_), .ZN(new_n3554_));
  XOR2_X1    g01088(.A1(pi0146), .A2(pi0284), .Z(new_n3555_));
  AOI21_X1   g01089(.A1(new_n3377_), .A2(pi0146), .B(new_n3555_), .ZN(new_n3556_));
  NOR2_X1    g01090(.A1(new_n3428_), .A2(pi0284), .ZN(new_n3557_));
  OAI22_X1   g01091(.A1(new_n3556_), .A2(new_n3557_), .B1(pi0146), .B2(new_n3426_), .ZN(new_n3558_));
  NOR2_X1    g01092(.A1(new_n3421_), .A2(new_n2525_), .ZN(new_n3559_));
  INV_X1     g01093(.I(pi0146), .ZN(new_n3560_));
  INV_X1     g01094(.I(pi0284), .ZN(new_n3561_));
  NOR2_X1    g01095(.A1(new_n2438_), .A2(new_n3561_), .ZN(new_n3562_));
  NAND4_X1   g01096(.A1(new_n3562_), .A2(pi0105), .A3(new_n3560_), .A4(new_n2523_), .ZN(new_n3563_));
  INV_X1     g01097(.I(new_n3563_), .ZN(new_n3564_));
  NOR3_X1    g01098(.A1(new_n3559_), .A2(pi0228), .A3(new_n3564_), .ZN(new_n3565_));
  AOI21_X1   g01099(.A1(new_n3558_), .A2(new_n3565_), .B(pi0216), .ZN(new_n3566_));
  OAI21_X1   g01100(.A1(new_n3566_), .A2(new_n3554_), .B(new_n3552_), .ZN(new_n3567_));
  OAI21_X1   g01101(.A1(new_n3567_), .A2(pi0215), .B(new_n3548_), .ZN(new_n3568_));
  NAND3_X1   g01102(.A1(new_n3567_), .A2(new_n2566_), .A3(pi1143), .ZN(new_n3569_));
  AOI21_X1   g01103(.A1(new_n3568_), .A2(new_n3569_), .B(new_n2587_), .ZN(new_n3570_));
  NAND3_X1   g01104(.A1(new_n2589_), .A2(pi0944), .A3(new_n3548_), .ZN(new_n3571_));
  OAI21_X1   g01105(.A1(new_n2593_), .A2(pi0944), .B(pi1143), .ZN(new_n3572_));
  AOI21_X1   g01106(.A1(new_n3572_), .A2(new_n3571_), .B(new_n2588_), .ZN(new_n3573_));
  INV_X1     g01107(.I(new_n3573_), .ZN(new_n3574_));
  AOI21_X1   g01108(.A1(pi0224), .A2(pi0264), .B(pi0222), .ZN(new_n3575_));
  INV_X1     g01109(.I(new_n3575_), .ZN(new_n3576_));
  AOI21_X1   g01110(.A1(new_n3421_), .A2(new_n3561_), .B(pi0224), .ZN(new_n3577_));
  OAI21_X1   g01111(.A1(new_n3577_), .A2(new_n3576_), .B(new_n3574_), .ZN(new_n3578_));
  OAI21_X1   g01112(.A1(new_n2604_), .A2(new_n3548_), .B(new_n2587_), .ZN(new_n3579_));
  NAND3_X1   g01113(.A1(new_n3578_), .A2(new_n3422_), .A3(new_n3575_), .ZN(new_n3580_));
  NOR2_X1    g01114(.A1(pi0223), .A2(pi0299), .ZN(new_n3581_));
  AOI21_X1   g01115(.A1(new_n3580_), .A2(new_n3581_), .B(pi0039), .ZN(new_n3582_));
  OR3_X2     g01116(.A1(new_n3582_), .A2(new_n3578_), .A3(new_n3579_), .Z(new_n3583_));
  NAND3_X1   g01117(.A1(new_n3562_), .A2(new_n2595_), .A3(new_n3576_), .ZN(new_n3584_));
  NAND2_X1   g01118(.A1(new_n3574_), .A2(new_n3584_), .ZN(new_n3585_));
  NAND3_X1   g01119(.A1(new_n3585_), .A2(new_n2604_), .A3(pi1143), .ZN(new_n3586_));
  OAI21_X1   g01120(.A1(new_n3585_), .A2(pi0223), .B(new_n3548_), .ZN(new_n3587_));
  NAND3_X1   g01121(.A1(new_n3587_), .A2(new_n3586_), .A3(new_n2587_), .ZN(new_n3588_));
  INV_X1     g01122(.I(new_n3588_), .ZN(new_n3589_));
  INV_X1     g01123(.I(new_n3156_), .ZN(new_n3590_));
  NOR2_X1    g01124(.A1(new_n3590_), .A2(new_n2974_), .ZN(new_n3591_));
  NOR2_X1    g01125(.A1(new_n3589_), .A2(new_n3591_), .ZN(new_n3592_));
  NOR2_X1    g01126(.A1(new_n2566_), .A2(new_n3548_), .ZN(new_n3593_));
  INV_X1     g01127(.I(new_n3554_), .ZN(new_n3594_));
  NOR2_X1    g01128(.A1(new_n3564_), .A2(new_n3282_), .ZN(new_n3595_));
  INV_X1     g01129(.I(new_n3595_), .ZN(new_n3596_));
  NOR3_X1    g01130(.A1(new_n2490_), .A2(new_n3560_), .A3(new_n3561_), .ZN(new_n3597_));
  AOI21_X1   g01131(.A1(new_n2491_), .A2(new_n3560_), .B(pi0284), .ZN(new_n3598_));
  NOR3_X1    g01132(.A1(new_n3598_), .A2(pi0228), .A3(new_n3597_), .ZN(new_n3599_));
  INV_X1     g01133(.I(new_n3599_), .ZN(new_n3600_));
  OAI21_X1   g01134(.A1(new_n3600_), .A2(new_n3596_), .B(new_n2562_), .ZN(new_n3601_));
  NAND2_X1   g01135(.A1(new_n3601_), .A2(new_n3594_), .ZN(new_n3602_));
  AOI21_X1   g01136(.A1(new_n3602_), .A2(new_n3552_), .B(pi0215), .ZN(new_n3603_));
  NOR2_X1    g01137(.A1(new_n3603_), .A2(new_n3593_), .ZN(new_n3604_));
  AOI21_X1   g01138(.A1(new_n3604_), .A2(pi0299), .B(new_n3592_), .ZN(new_n3605_));
  INV_X1     g01139(.I(new_n3245_), .ZN(new_n3608_));
  NOR2_X1    g01140(.A1(new_n3608_), .A2(pi0146), .ZN(new_n3609_));
  NOR4_X1    g01141(.A1(new_n2490_), .A2(new_n3181_), .A3(pi0284), .A4(new_n2985_), .ZN(new_n3610_));
  AOI21_X1   g01142(.A1(new_n3560_), .A2(new_n2523_), .B(new_n3596_), .ZN(new_n3617_));
  OAI21_X1   g01143(.A1(new_n3617_), .A2(pi0216), .B(new_n3594_), .ZN(new_n3618_));
  AOI21_X1   g01144(.A1(new_n3618_), .A2(new_n3552_), .B(pi0215), .ZN(new_n3619_));
  NOR2_X1    g01145(.A1(new_n3619_), .A2(new_n3593_), .ZN(new_n3620_));
  AOI21_X1   g01146(.A1(new_n3620_), .A2(pi0299), .B(new_n3592_), .ZN(new_n3621_));
  NAND2_X1   g01147(.A1(new_n3172_), .A2(new_n3173_), .ZN(new_n3622_));
  AOI21_X1   g01148(.A1(new_n3605_), .A2(new_n3154_), .B(new_n3622_), .ZN(new_n3623_));
  OAI21_X1   g01149(.A1(new_n3570_), .A2(new_n3583_), .B(new_n3623_), .ZN(new_n3624_));
  AOI21_X1   g01150(.A1(new_n3624_), .A2(new_n3177_), .B(pi0075), .ZN(new_n3625_));
  INV_X1     g01151(.I(new_n3621_), .ZN(new_n3626_));
  NOR2_X1    g01152(.A1(new_n3605_), .A2(new_n3198_), .ZN(new_n3627_));
  AOI21_X1   g01153(.A1(new_n3198_), .A2(new_n3626_), .B(new_n3627_), .ZN(new_n3628_));
  OR2_X2     g01154(.A1(new_n3628_), .A2(new_n3177_), .Z(new_n3629_));
  NOR4_X1    g01155(.A1(new_n3628_), .A2(pi0092), .A3(new_n2535_), .A4(new_n3621_), .ZN(new_n3630_));
  AOI21_X1   g01156(.A1(new_n3621_), .A2(new_n2539_), .B(pi0055), .ZN(new_n3631_));
  NOR2_X1    g01157(.A1(new_n3626_), .A2(new_n2628_), .ZN(new_n3632_));
  NOR4_X1    g01158(.A1(new_n3630_), .A2(new_n3330_), .A3(new_n3631_), .A4(new_n3632_), .ZN(new_n3633_));
  OAI21_X1   g01159(.A1(new_n3625_), .A2(new_n3629_), .B(new_n3633_), .ZN(new_n3634_));
  INV_X1     g01160(.I(new_n3604_), .ZN(new_n3635_));
  INV_X1     g01161(.I(new_n3620_), .ZN(new_n3636_));
  MUX2_X1    g01162(.I0(new_n3635_), .I1(new_n3636_), .S(new_n3336_), .Z(new_n3637_));
  NOR2_X1    g01163(.A1(new_n3635_), .A2(new_n3234_), .ZN(new_n3638_));
  OAI21_X1   g01164(.A1(new_n3636_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n3639_));
  OAI21_X1   g01165(.A1(new_n3638_), .A2(new_n3639_), .B(new_n2533_), .ZN(new_n3640_));
  AOI21_X1   g01166(.A1(pi0056), .A2(new_n3637_), .B(new_n3640_), .ZN(new_n3641_));
  NOR2_X1    g01167(.A1(new_n3635_), .A2(new_n3400_), .ZN(new_n3642_));
  OAI21_X1   g01168(.A1(new_n3636_), .A2(new_n3343_), .B(new_n3240_), .ZN(new_n3643_));
  NOR2_X1    g01169(.A1(new_n3405_), .A2(pi0238), .ZN(new_n3644_));
  OAI21_X1   g01170(.A1(new_n3642_), .A2(new_n3643_), .B(new_n3644_), .ZN(new_n3645_));
  AOI21_X1   g01171(.A1(new_n3634_), .A2(new_n3641_), .B(new_n3645_), .ZN(new_n3646_));
  INV_X1     g01172(.I(pi0238), .ZN(new_n3647_));
  NAND2_X1   g01173(.A1(new_n3485_), .A2(new_n3553_), .ZN(new_n3648_));
  NOR4_X1    g01174(.A1(new_n3636_), .A2(new_n3647_), .A3(new_n2571_), .A4(new_n3648_), .ZN(new_n3649_));
  NAND2_X1   g01175(.A1(new_n3430_), .A2(new_n3564_), .ZN(new_n3650_));
  INV_X1     g01176(.I(new_n3426_), .ZN(new_n3651_));
  NOR4_X1    g01177(.A1(new_n3651_), .A2(new_n3560_), .A3(pi0284), .A4(new_n3428_), .ZN(new_n3652_));
  NOR3_X1    g01178(.A1(new_n3377_), .A2(pi0146), .A3(pi0284), .ZN(new_n3653_));
  OAI21_X1   g01179(.A1(new_n3653_), .A2(new_n3652_), .B(new_n2523_), .ZN(new_n3654_));
  AOI21_X1   g01180(.A1(new_n3654_), .A2(new_n3650_), .B(pi0216), .ZN(new_n3655_));
  OAI21_X1   g01181(.A1(new_n3655_), .A2(new_n3554_), .B(new_n3552_), .ZN(new_n3656_));
  OAI21_X1   g01182(.A1(new_n3656_), .A2(pi0215), .B(new_n3548_), .ZN(new_n3657_));
  NAND3_X1   g01183(.A1(new_n3656_), .A2(new_n2566_), .A3(pi1143), .ZN(new_n3658_));
  AOI21_X1   g01184(.A1(new_n3657_), .A2(new_n3658_), .B(new_n2587_), .ZN(new_n3659_));
  NOR2_X1    g01185(.A1(new_n2550_), .A2(pi0216), .ZN(new_n3660_));
  OAI21_X1   g01186(.A1(new_n3600_), .A2(new_n3564_), .B(new_n3660_), .ZN(new_n3661_));
  NAND2_X1   g01187(.A1(new_n3661_), .A2(new_n3552_), .ZN(new_n3662_));
  AOI21_X1   g01188(.A1(new_n3662_), .A2(new_n2566_), .B(new_n3593_), .ZN(new_n3663_));
  AOI21_X1   g01189(.A1(new_n3663_), .A2(pi0299), .B(new_n3588_), .ZN(new_n3664_));
  OAI21_X1   g01190(.A1(new_n3664_), .A2(new_n3154_), .B(new_n3172_), .ZN(new_n3665_));
  NAND2_X1   g01191(.A1(new_n3636_), .A2(new_n3648_), .ZN(new_n3666_));
  AOI21_X1   g01192(.A1(new_n3666_), .A2(pi0299), .B(new_n3588_), .ZN(new_n3667_));
  INV_X1     g01193(.I(new_n3667_), .ZN(new_n3668_));
  OAI21_X1   g01194(.A1(new_n3668_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n3669_));
  NAND3_X1   g01195(.A1(new_n3582_), .A2(new_n3669_), .A3(new_n3665_), .ZN(new_n3670_));
  INV_X1     g01196(.I(new_n3189_), .ZN(new_n3671_));
  INV_X1     g01197(.I(new_n3660_), .ZN(new_n3672_));
  NOR4_X1    g01198(.A1(new_n3609_), .A2(pi0228), .A3(new_n3564_), .A4(new_n3610_), .ZN(new_n3673_));
  OAI21_X1   g01199(.A1(new_n3673_), .A2(new_n3672_), .B(new_n3552_), .ZN(new_n3674_));
  AOI21_X1   g01200(.A1(new_n3674_), .A2(new_n2566_), .B(new_n3593_), .ZN(new_n3675_));
  NOR3_X1    g01201(.A1(new_n3675_), .A2(new_n3671_), .A3(new_n3588_), .ZN(new_n3676_));
  OAI21_X1   g01202(.A1(new_n3668_), .A2(new_n2544_), .B(pi0100), .ZN(new_n3677_));
  OAI22_X1   g01203(.A1(new_n3659_), .A2(new_n3670_), .B1(new_n3676_), .B2(new_n3677_), .ZN(new_n3678_));
  AOI21_X1   g01204(.A1(new_n3678_), .A2(new_n3177_), .B(pi0075), .ZN(new_n3679_));
  NOR2_X1    g01205(.A1(new_n3664_), .A2(new_n3198_), .ZN(new_n3680_));
  AOI21_X1   g01206(.A1(new_n3198_), .A2(new_n3668_), .B(new_n3680_), .ZN(new_n3681_));
  OR2_X2     g01207(.A1(new_n3681_), .A2(new_n3177_), .Z(new_n3682_));
  NOR4_X1    g01208(.A1(new_n3681_), .A2(pi0092), .A3(new_n2535_), .A4(new_n3667_), .ZN(new_n3683_));
  AOI21_X1   g01209(.A1(new_n3667_), .A2(new_n2539_), .B(pi0055), .ZN(new_n3684_));
  NOR2_X1    g01210(.A1(new_n3668_), .A2(new_n2628_), .ZN(new_n3685_));
  NOR4_X1    g01211(.A1(new_n3683_), .A2(new_n3330_), .A3(new_n3684_), .A4(new_n3685_), .ZN(new_n3686_));
  OAI21_X1   g01212(.A1(new_n3679_), .A2(new_n3682_), .B(new_n3686_), .ZN(new_n3687_));
  INV_X1     g01213(.I(new_n3663_), .ZN(new_n3688_));
  INV_X1     g01214(.I(new_n3666_), .ZN(new_n3689_));
  MUX2_X1    g01215(.I0(new_n3688_), .I1(new_n3689_), .S(new_n3336_), .Z(new_n3690_));
  NOR2_X1    g01216(.A1(new_n3688_), .A2(new_n3234_), .ZN(new_n3691_));
  OAI21_X1   g01217(.A1(new_n3689_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n3692_));
  OAI21_X1   g01218(.A1(new_n3691_), .A2(new_n3692_), .B(new_n2533_), .ZN(new_n3693_));
  AOI21_X1   g01219(.A1(pi0056), .A2(new_n3690_), .B(new_n3693_), .ZN(new_n3694_));
  AOI21_X1   g01220(.A1(new_n3666_), .A2(new_n3400_), .B(pi0062), .ZN(new_n3695_));
  OAI21_X1   g01221(.A1(new_n3688_), .A2(new_n3400_), .B(new_n3695_), .ZN(new_n3696_));
  NAND3_X1   g01222(.A1(new_n3696_), .A2(pi0238), .A3(new_n2571_), .ZN(new_n3697_));
  AOI21_X1   g01223(.A1(new_n3687_), .A2(new_n3694_), .B(new_n3697_), .ZN(new_n3698_));
  NOR3_X1    g01224(.A1(new_n3698_), .A2(new_n3646_), .A3(new_n3649_), .ZN(po0156));
  INV_X1     g01225(.I(pi1142), .ZN(new_n3700_));
  INV_X1     g01226(.I(pi0932), .ZN(new_n3701_));
  NOR3_X1    g01227(.A1(new_n2555_), .A2(new_n3701_), .A3(pi1142), .ZN(new_n3702_));
  AOI21_X1   g01228(.A1(new_n2554_), .A2(new_n3701_), .B(new_n3700_), .ZN(new_n3703_));
  OAI21_X1   g01229(.A1(new_n3702_), .A2(new_n3703_), .B(pi0221), .ZN(new_n3704_));
  INV_X1     g01230(.I(new_n3704_), .ZN(new_n3705_));
  AOI21_X1   g01231(.A1(pi0216), .A2(pi0277), .B(pi0221), .ZN(new_n3706_));
  INV_X1     g01232(.I(pi0172), .ZN(new_n3707_));
  OAI21_X1   g01233(.A1(new_n3376_), .A2(new_n3428_), .B(pi0262), .ZN(new_n3708_));
  NOR2_X1    g01234(.A1(new_n3708_), .A2(new_n3707_), .ZN(new_n3709_));
  AOI21_X1   g01235(.A1(new_n3426_), .A2(pi0262), .B(pi0172), .ZN(new_n3710_));
  OAI21_X1   g01236(.A1(new_n3707_), .A2(pi0105), .B(pi0228), .ZN(new_n3711_));
  INV_X1     g01237(.I(pi0262), .ZN(new_n3712_));
  NOR2_X1    g01238(.A1(new_n2438_), .A2(new_n3712_), .ZN(new_n3713_));
  NAND4_X1   g01239(.A1(new_n3419_), .A2(pi0105), .A3(new_n3711_), .A4(new_n3713_), .ZN(new_n3714_));
  AOI21_X1   g01240(.A1(new_n3714_), .A2(new_n2562_), .B(pi0228), .ZN(new_n3715_));
  OAI21_X1   g01241(.A1(new_n3709_), .A2(new_n3710_), .B(new_n3715_), .ZN(new_n3716_));
  AOI21_X1   g01242(.A1(new_n3716_), .A2(new_n3706_), .B(new_n3705_), .ZN(new_n3717_));
  OAI21_X1   g01243(.A1(new_n3717_), .A2(pi0215), .B(new_n3700_), .ZN(new_n3718_));
  NAND3_X1   g01244(.A1(new_n3717_), .A2(new_n2566_), .A3(pi1142), .ZN(new_n3719_));
  AOI21_X1   g01245(.A1(new_n3718_), .A2(new_n3719_), .B(new_n2587_), .ZN(new_n3720_));
  NAND3_X1   g01246(.A1(new_n2589_), .A2(pi0932), .A3(new_n3700_), .ZN(new_n3721_));
  OAI21_X1   g01247(.A1(new_n2593_), .A2(pi0932), .B(pi1142), .ZN(new_n3722_));
  AOI21_X1   g01248(.A1(new_n3722_), .A2(new_n3721_), .B(new_n2588_), .ZN(new_n3723_));
  INV_X1     g01249(.I(new_n3713_), .ZN(new_n3724_));
  AOI21_X1   g01250(.A1(pi0224), .A2(pi0277), .B(pi0222), .ZN(new_n3725_));
  NOR3_X1    g01251(.A1(new_n3724_), .A2(pi0224), .A3(new_n3725_), .ZN(new_n3726_));
  OR2_X2     g01252(.A1(new_n3723_), .A2(new_n3726_), .Z(new_n3727_));
  NAND3_X1   g01253(.A1(new_n3727_), .A2(new_n2604_), .A3(pi1142), .ZN(new_n3728_));
  OAI21_X1   g01254(.A1(new_n3727_), .A2(pi0223), .B(new_n3700_), .ZN(new_n3729_));
  NAND3_X1   g01255(.A1(new_n3729_), .A2(new_n3728_), .A3(new_n2587_), .ZN(new_n3730_));
  NOR2_X1    g01256(.A1(new_n2566_), .A2(new_n3700_), .ZN(new_n3731_));
  MUX2_X1    g01257(.I0(new_n3724_), .I1(new_n3707_), .S(new_n2522_), .Z(new_n3732_));
  NOR2_X1    g01258(.A1(new_n3732_), .A2(new_n2523_), .ZN(new_n3733_));
  OAI21_X1   g01259(.A1(new_n2491_), .A2(pi0262), .B(new_n2523_), .ZN(new_n3734_));
  AOI21_X1   g01260(.A1(new_n3707_), .A2(new_n2491_), .B(new_n3734_), .ZN(new_n3735_));
  NOR2_X1    g01261(.A1(new_n2550_), .A2(pi0216), .ZN(new_n3736_));
  OAI21_X1   g01262(.A1(new_n3735_), .A2(new_n3733_), .B(new_n3736_), .ZN(new_n3737_));
  AOI21_X1   g01263(.A1(new_n3737_), .A2(new_n3704_), .B(pi0215), .ZN(new_n3738_));
  NOR2_X1    g01264(.A1(new_n3738_), .A2(new_n3731_), .ZN(new_n3739_));
  AOI21_X1   g01265(.A1(new_n3739_), .A2(pi0299), .B(new_n3730_), .ZN(new_n3740_));
  OAI21_X1   g01266(.A1(new_n3740_), .A2(new_n3154_), .B(new_n3172_), .ZN(new_n3741_));
  AOI21_X1   g01267(.A1(pi0172), .A2(new_n2523_), .B(new_n3733_), .ZN(new_n3742_));
  OAI21_X1   g01268(.A1(new_n3742_), .A2(pi0216), .B(new_n3706_), .ZN(new_n3743_));
  AOI21_X1   g01269(.A1(new_n3743_), .A2(new_n3704_), .B(pi0215), .ZN(new_n3744_));
  NOR2_X1    g01270(.A1(new_n3744_), .A2(new_n3731_), .ZN(new_n3745_));
  AOI21_X1   g01271(.A1(new_n3745_), .A2(pi0299), .B(new_n3730_), .ZN(new_n3746_));
  INV_X1     g01272(.I(new_n3746_), .ZN(new_n3747_));
  OAI21_X1   g01273(.A1(new_n3747_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n3748_));
  OAI21_X1   g01274(.A1(new_n3422_), .A2(pi0262), .B(new_n2595_), .ZN(new_n3749_));
  AOI21_X1   g01275(.A1(new_n3749_), .A2(new_n3725_), .B(new_n3723_), .ZN(new_n3750_));
  NAND2_X1   g01276(.A1(new_n3422_), .A2(new_n3725_), .ZN(new_n3751_));
  NOR2_X1    g01277(.A1(pi0223), .A2(pi0299), .ZN(new_n3752_));
  OAI21_X1   g01278(.A1(new_n3750_), .A2(new_n3751_), .B(new_n3752_), .ZN(new_n3753_));
  NAND4_X1   g01279(.A1(new_n3753_), .A2(new_n3741_), .A3(new_n3154_), .A4(new_n3748_), .ZN(new_n3754_));
  OAI21_X1   g01280(.A1(new_n3256_), .A2(pi0262), .B(new_n2523_), .ZN(new_n3755_));
  AOI21_X1   g01281(.A1(new_n3707_), .A2(new_n3256_), .B(new_n3755_), .ZN(new_n3756_));
  OAI21_X1   g01282(.A1(new_n3756_), .A2(new_n3733_), .B(new_n3736_), .ZN(new_n3757_));
  NAND2_X1   g01283(.A1(new_n3757_), .A2(new_n3704_), .ZN(new_n3758_));
  AOI21_X1   g01284(.A1(new_n3758_), .A2(new_n2566_), .B(new_n3731_), .ZN(new_n3759_));
  NOR3_X1    g01285(.A1(new_n3759_), .A2(new_n3671_), .A3(new_n3730_), .ZN(new_n3760_));
  OAI21_X1   g01286(.A1(new_n3747_), .A2(new_n2544_), .B(pi0100), .ZN(new_n3761_));
  OAI22_X1   g01287(.A1(new_n3720_), .A2(new_n3754_), .B1(new_n3760_), .B2(new_n3761_), .ZN(new_n3762_));
  AOI21_X1   g01288(.A1(new_n3762_), .A2(new_n3177_), .B(pi0075), .ZN(new_n3763_));
  NOR2_X1    g01289(.A1(new_n3740_), .A2(new_n3198_), .ZN(new_n3764_));
  AOI21_X1   g01290(.A1(new_n3198_), .A2(new_n3747_), .B(new_n3764_), .ZN(new_n3765_));
  OR2_X2     g01291(.A1(new_n3765_), .A2(new_n3177_), .Z(new_n3766_));
  NOR4_X1    g01292(.A1(new_n3765_), .A2(pi0092), .A3(new_n2535_), .A4(new_n3746_), .ZN(new_n3767_));
  AOI21_X1   g01293(.A1(new_n3746_), .A2(new_n2539_), .B(pi0055), .ZN(new_n3768_));
  NOR2_X1    g01294(.A1(new_n3747_), .A2(new_n2628_), .ZN(new_n3769_));
  NOR4_X1    g01295(.A1(new_n3767_), .A2(new_n3330_), .A3(new_n3768_), .A4(new_n3769_), .ZN(new_n3770_));
  OAI21_X1   g01296(.A1(new_n3763_), .A2(new_n3766_), .B(new_n3770_), .ZN(new_n3771_));
  INV_X1     g01297(.I(new_n3739_), .ZN(new_n3772_));
  INV_X1     g01298(.I(new_n3745_), .ZN(new_n3773_));
  MUX2_X1    g01299(.I0(new_n3772_), .I1(new_n3773_), .S(new_n3336_), .Z(new_n3774_));
  NOR2_X1    g01300(.A1(new_n3772_), .A2(new_n3234_), .ZN(new_n3775_));
  OAI21_X1   g01301(.A1(new_n3773_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n3776_));
  OAI21_X1   g01302(.A1(new_n3775_), .A2(new_n3776_), .B(new_n2533_), .ZN(new_n3777_));
  AOI21_X1   g01303(.A1(pi0056), .A2(new_n3774_), .B(new_n3777_), .ZN(new_n3778_));
  NOR2_X1    g01304(.A1(new_n3772_), .A2(new_n3400_), .ZN(new_n3779_));
  OAI21_X1   g01305(.A1(new_n3773_), .A2(new_n3343_), .B(new_n3240_), .ZN(new_n3780_));
  OAI21_X1   g01306(.A1(new_n3779_), .A2(new_n3780_), .B(new_n2571_), .ZN(new_n3781_));
  AOI21_X1   g01307(.A1(new_n3771_), .A2(new_n3778_), .B(new_n3781_), .ZN(new_n3782_));
  OAI21_X1   g01308(.A1(new_n3745_), .A2(new_n2571_), .B(pi0249), .ZN(new_n3783_));
  NAND2_X1   g01309(.A1(pi0223), .A2(pi1142), .ZN(new_n3784_));
  NAND2_X1   g01310(.A1(new_n3753_), .A2(new_n3154_), .ZN(new_n3785_));
  NAND4_X1   g01311(.A1(new_n3785_), .A2(new_n2587_), .A3(new_n3750_), .A4(new_n3784_), .ZN(new_n3794_));
  OAI21_X1   g01312(.A1(new_n3732_), .A2(new_n2523_), .B(new_n3283_), .ZN(new_n3795_));
  OAI21_X1   g01313(.A1(new_n3756_), .A2(new_n3795_), .B(new_n2562_), .ZN(new_n3796_));
  NAND2_X1   g01314(.A1(new_n3796_), .A2(new_n3706_), .ZN(new_n3797_));
  AOI21_X1   g01315(.A1(new_n3797_), .A2(new_n3704_), .B(pi0215), .ZN(new_n3798_));
  INV_X1     g01316(.I(new_n3730_), .ZN(new_n3799_));
  NOR2_X1    g01317(.A1(new_n3799_), .A2(new_n3591_), .ZN(new_n3800_));
  NOR2_X1    g01318(.A1(new_n3800_), .A2(new_n3671_), .ZN(new_n3801_));
  OAI21_X1   g01319(.A1(new_n3798_), .A2(new_n3731_), .B(new_n3801_), .ZN(new_n3802_));
  NOR2_X1    g01320(.A1(new_n3773_), .A2(new_n3288_), .ZN(new_n3803_));
  AOI21_X1   g01321(.A1(new_n3803_), .A2(pi0299), .B(new_n3800_), .ZN(new_n3804_));
  AOI21_X1   g01322(.A1(new_n3804_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n3805_));
  INV_X1     g01323(.I(new_n3731_), .ZN(new_n3806_));
  OAI21_X1   g01324(.A1(new_n3735_), .A2(new_n3795_), .B(new_n2562_), .ZN(new_n3807_));
  AOI21_X1   g01325(.A1(new_n3807_), .A2(new_n3706_), .B(new_n3705_), .ZN(new_n3808_));
  OAI21_X1   g01326(.A1(new_n3808_), .A2(pi0215), .B(new_n3806_), .ZN(new_n3809_));
  OAI22_X1   g01327(.A1(new_n3809_), .A2(new_n2587_), .B1(new_n3591_), .B2(new_n3799_), .ZN(new_n3810_));
  NOR2_X1    g01328(.A1(pi0038), .A2(pi0100), .ZN(new_n3811_));
  OAI21_X1   g01329(.A1(new_n3810_), .A2(pi0039), .B(new_n3811_), .ZN(new_n3812_));
  AOI21_X1   g01330(.A1(new_n3802_), .A2(new_n3805_), .B(new_n3812_), .ZN(new_n3813_));
  AOI21_X1   g01331(.A1(new_n3813_), .A2(new_n3794_), .B(pi0087), .ZN(new_n3814_));
  NOR2_X1    g01332(.A1(new_n3804_), .A2(new_n3197_), .ZN(new_n3815_));
  AOI21_X1   g01333(.A1(new_n3197_), .A2(new_n3810_), .B(new_n3815_), .ZN(new_n3816_));
  NOR2_X1    g01334(.A1(new_n3816_), .A2(new_n3177_), .ZN(new_n3817_));
  OAI21_X1   g01335(.A1(new_n3814_), .A2(pi0075), .B(new_n3817_), .ZN(new_n3818_));
  NOR4_X1    g01336(.A1(new_n3816_), .A2(pi0092), .A3(new_n2535_), .A4(new_n3804_), .ZN(new_n3819_));
  AOI21_X1   g01337(.A1(new_n3804_), .A2(new_n2539_), .B(pi0055), .ZN(new_n3820_));
  AND2_X2    g01338(.A1(new_n3804_), .A2(pi0075), .Z(new_n3821_));
  NOR4_X1    g01339(.A1(new_n3819_), .A2(new_n3330_), .A3(new_n3820_), .A4(new_n3821_), .ZN(new_n3822_));
  INV_X1     g01340(.I(new_n3803_), .ZN(new_n3823_));
  NAND4_X1   g01341(.A1(new_n3823_), .A2(new_n3335_), .A3(new_n2548_), .A4(new_n3809_), .ZN(new_n3824_));
  NAND2_X1   g01342(.A1(new_n3824_), .A2(new_n2533_), .ZN(new_n3825_));
  AOI21_X1   g01343(.A1(new_n3818_), .A2(new_n3822_), .B(new_n3825_), .ZN(new_n3826_));
  NOR2_X1    g01344(.A1(new_n3826_), .A2(new_n3405_), .ZN(new_n3827_));
  INV_X1     g01345(.I(pi0249), .ZN(new_n3828_));
  OAI21_X1   g01346(.A1(new_n3803_), .A2(new_n2571_), .B(new_n3828_), .ZN(new_n3829_));
  OAI22_X1   g01347(.A1(new_n3782_), .A2(new_n3783_), .B1(new_n3827_), .B2(new_n3829_), .ZN(po0157));
  INV_X1     g01348(.I(pi1141), .ZN(new_n3831_));
  INV_X1     g01349(.I(pi0935), .ZN(new_n3832_));
  NOR3_X1    g01350(.A1(new_n2555_), .A2(new_n3832_), .A3(pi1141), .ZN(new_n3833_));
  AOI21_X1   g01351(.A1(new_n2554_), .A2(new_n3832_), .B(new_n3831_), .ZN(new_n3834_));
  OAI21_X1   g01352(.A1(new_n3833_), .A2(new_n3834_), .B(pi0221), .ZN(new_n3835_));
  INV_X1     g01353(.I(new_n3835_), .ZN(new_n3836_));
  AOI21_X1   g01354(.A1(pi0216), .A2(pi0270), .B(pi0221), .ZN(new_n3837_));
  MUX2_X1    g01355(.I0(new_n3428_), .I1(new_n3377_), .S(pi0861), .Z(new_n3838_));
  INV_X1     g01356(.I(pi0861), .ZN(new_n3839_));
  AOI21_X1   g01357(.A1(new_n3426_), .A2(new_n3839_), .B(pi0171), .ZN(new_n3840_));
  AOI21_X1   g01358(.A1(new_n3838_), .A2(pi0171), .B(new_n3840_), .ZN(new_n3841_));
  INV_X1     g01359(.I(pi0171), .ZN(new_n3842_));
  NOR2_X1    g01360(.A1(new_n2438_), .A2(new_n3839_), .ZN(new_n3843_));
  NAND4_X1   g01361(.A1(new_n3843_), .A2(pi0105), .A3(new_n3842_), .A4(new_n2523_), .ZN(new_n3844_));
  INV_X1     g01362(.I(new_n3844_), .ZN(new_n3845_));
  NOR2_X1    g01363(.A1(new_n3845_), .A2(pi0216), .ZN(new_n3846_));
  INV_X1     g01364(.I(new_n3846_), .ZN(new_n3847_));
  NOR2_X1    g01365(.A1(new_n3559_), .A2(new_n3847_), .ZN(new_n3848_));
  OAI21_X1   g01366(.A1(new_n3841_), .A2(pi0228), .B(new_n3848_), .ZN(new_n3849_));
  AOI21_X1   g01367(.A1(new_n3849_), .A2(new_n3837_), .B(new_n3836_), .ZN(new_n3850_));
  MUX2_X1    g01368(.I0(new_n3850_), .I1(new_n3831_), .S(pi0215), .Z(new_n3851_));
  NAND3_X1   g01369(.A1(new_n2589_), .A2(pi0935), .A3(new_n3831_), .ZN(new_n3852_));
  OAI21_X1   g01370(.A1(new_n2593_), .A2(pi0935), .B(pi1141), .ZN(new_n3853_));
  AOI21_X1   g01371(.A1(new_n3853_), .A2(new_n3852_), .B(new_n2588_), .ZN(new_n3854_));
  INV_X1     g01372(.I(new_n3854_), .ZN(new_n3855_));
  AOI21_X1   g01373(.A1(pi0224), .A2(pi0270), .B(pi0222), .ZN(new_n3856_));
  OAI21_X1   g01374(.A1(new_n3843_), .A2(pi0224), .B(new_n3856_), .ZN(new_n3857_));
  NAND2_X1   g01375(.A1(new_n3855_), .A2(new_n3857_), .ZN(new_n3858_));
  NAND3_X1   g01376(.A1(new_n3858_), .A2(new_n2604_), .A3(pi1141), .ZN(new_n3859_));
  OAI21_X1   g01377(.A1(new_n3858_), .A2(pi0223), .B(new_n3831_), .ZN(new_n3860_));
  NAND3_X1   g01378(.A1(new_n3860_), .A2(new_n3859_), .A3(new_n2587_), .ZN(new_n3861_));
  NOR2_X1    g01379(.A1(new_n3861_), .A2(new_n3297_), .ZN(new_n3862_));
  INV_X1     g01380(.I(new_n3862_), .ZN(new_n3863_));
  NOR2_X1    g01381(.A1(new_n2566_), .A2(new_n3831_), .ZN(new_n3864_));
  NOR3_X1    g01382(.A1(new_n2490_), .A2(new_n3842_), .A3(new_n3839_), .ZN(new_n3865_));
  AOI21_X1   g01383(.A1(new_n2491_), .A2(new_n3842_), .B(pi0861), .ZN(new_n3866_));
  NOR4_X1    g01384(.A1(new_n3866_), .A2(pi0228), .A3(new_n3282_), .A4(new_n3865_), .ZN(new_n3867_));
  NOR2_X1    g01385(.A1(new_n3846_), .A2(new_n3837_), .ZN(new_n3868_));
  INV_X1     g01386(.I(new_n3868_), .ZN(new_n3869_));
  OAI21_X1   g01387(.A1(new_n3867_), .A2(new_n3869_), .B(new_n3835_), .ZN(new_n3870_));
  AOI21_X1   g01388(.A1(new_n3870_), .A2(new_n2566_), .B(new_n3864_), .ZN(new_n3871_));
  AOI21_X1   g01389(.A1(new_n3871_), .A2(pi0299), .B(new_n3863_), .ZN(new_n3872_));
  OAI21_X1   g01390(.A1(new_n3872_), .A2(new_n3154_), .B(new_n3172_), .ZN(new_n3873_));
  OAI21_X1   g01391(.A1(new_n3422_), .A2(new_n3839_), .B(new_n2595_), .ZN(new_n3874_));
  AOI21_X1   g01392(.A1(new_n3874_), .A2(new_n3856_), .B(new_n3854_), .ZN(new_n3875_));
  NAND2_X1   g01393(.A1(new_n3422_), .A2(new_n3856_), .ZN(new_n3876_));
  NOR2_X1    g01394(.A1(pi0223), .A2(pi0299), .ZN(new_n3877_));
  OAI21_X1   g01395(.A1(new_n3875_), .A2(new_n3876_), .B(new_n3877_), .ZN(new_n3878_));
  INV_X1     g01396(.I(new_n3864_), .ZN(new_n3879_));
  AOI21_X1   g01397(.A1(new_n3842_), .A2(new_n2523_), .B(new_n3837_), .ZN(new_n3880_));
  NAND2_X1   g01398(.A1(new_n3846_), .A2(new_n3880_), .ZN(new_n3881_));
  NAND2_X1   g01399(.A1(new_n3881_), .A2(new_n3835_), .ZN(new_n3882_));
  NAND2_X1   g01400(.A1(new_n3882_), .A2(new_n2566_), .ZN(new_n3883_));
  NAND2_X1   g01401(.A1(new_n3883_), .A2(new_n3879_), .ZN(new_n3884_));
  INV_X1     g01402(.I(new_n3884_), .ZN(new_n3885_));
  INV_X1     g01403(.I(new_n3485_), .ZN(new_n3886_));
  AOI21_X1   g01404(.A1(pi0216), .A2(pi0270), .B(new_n3886_), .ZN(new_n3887_));
  NOR2_X1    g01405(.A1(new_n3885_), .A2(new_n3887_), .ZN(new_n3888_));
  INV_X1     g01406(.I(new_n3888_), .ZN(new_n3889_));
  AOI21_X1   g01407(.A1(new_n3889_), .A2(pi0299), .B(new_n3863_), .ZN(new_n3890_));
  INV_X1     g01408(.I(new_n3890_), .ZN(new_n3891_));
  OAI21_X1   g01409(.A1(new_n3891_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n3892_));
  NAND4_X1   g01410(.A1(new_n3878_), .A2(new_n3154_), .A3(new_n3873_), .A4(new_n3892_), .ZN(new_n3893_));
  AOI21_X1   g01411(.A1(new_n3851_), .A2(pi0299), .B(new_n3893_), .ZN(new_n3894_));
  NOR3_X1    g01412(.A1(new_n3257_), .A2(new_n3842_), .A3(new_n3839_), .ZN(new_n3895_));
  AOI21_X1   g01413(.A1(new_n3256_), .A2(new_n3842_), .B(pi0861), .ZN(new_n3896_));
  NOR3_X1    g01414(.A1(new_n3895_), .A2(pi0228), .A3(new_n3896_), .ZN(new_n3897_));
  NAND2_X1   g01415(.A1(new_n3897_), .A2(new_n3283_), .ZN(new_n3898_));
  AOI21_X1   g01416(.A1(new_n3898_), .A2(new_n3868_), .B(new_n3836_), .ZN(new_n3899_));
  OAI21_X1   g01417(.A1(new_n3899_), .A2(pi0215), .B(new_n3879_), .ZN(new_n3900_));
  NAND2_X1   g01418(.A1(new_n3900_), .A2(new_n2587_), .ZN(new_n3901_));
  NOR2_X1    g01419(.A1(new_n3863_), .A2(new_n2545_), .ZN(new_n3902_));
  OAI21_X1   g01420(.A1(new_n3891_), .A2(new_n2544_), .B(pi0100), .ZN(new_n3903_));
  AOI21_X1   g01421(.A1(new_n3901_), .A2(new_n3902_), .B(new_n3903_), .ZN(new_n3904_));
  OAI21_X1   g01422(.A1(new_n3894_), .A2(new_n3904_), .B(new_n3177_), .ZN(new_n3905_));
  NAND2_X1   g01423(.A1(new_n3891_), .A2(new_n3198_), .ZN(new_n3906_));
  OAI21_X1   g01424(.A1(new_n3198_), .A2(new_n3872_), .B(new_n3906_), .ZN(new_n3907_));
  NAND2_X1   g01425(.A1(new_n3907_), .A2(pi0087), .ZN(new_n3908_));
  AOI21_X1   g01426(.A1(new_n3905_), .A2(new_n2628_), .B(new_n3908_), .ZN(new_n3909_));
  NAND4_X1   g01427(.A1(new_n3907_), .A2(new_n3203_), .A3(new_n2534_), .A4(new_n3891_), .ZN(new_n3910_));
  OAI21_X1   g01428(.A1(new_n3891_), .A2(new_n2538_), .B(new_n3227_), .ZN(new_n3911_));
  NAND2_X1   g01429(.A1(new_n3890_), .A2(pi0075), .ZN(new_n3912_));
  NAND4_X1   g01430(.A1(new_n3910_), .A2(new_n3329_), .A3(new_n3911_), .A4(new_n3912_), .ZN(new_n3913_));
  INV_X1     g01431(.I(new_n3871_), .ZN(new_n3914_));
  MUX2_X1    g01432(.I0(new_n3914_), .I1(new_n3888_), .S(new_n3336_), .Z(new_n3915_));
  NOR2_X1    g01433(.A1(new_n3914_), .A2(new_n3234_), .ZN(new_n3916_));
  OAI21_X1   g01434(.A1(new_n3888_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n3917_));
  OAI21_X1   g01435(.A1(new_n3916_), .A2(new_n3917_), .B(new_n2533_), .ZN(new_n3918_));
  AOI21_X1   g01436(.A1(pi0056), .A2(new_n3915_), .B(new_n3918_), .ZN(new_n3919_));
  OAI21_X1   g01437(.A1(new_n3909_), .A2(new_n3913_), .B(new_n3919_), .ZN(new_n3920_));
  NAND2_X1   g01438(.A1(new_n3871_), .A2(new_n3343_), .ZN(new_n3921_));
  AOI21_X1   g01439(.A1(new_n3889_), .A2(new_n3400_), .B(pi0062), .ZN(new_n3922_));
  NAND2_X1   g01440(.A1(new_n2571_), .A2(pi0241), .ZN(new_n3923_));
  AOI21_X1   g01441(.A1(new_n3922_), .A2(new_n3921_), .B(new_n3923_), .ZN(new_n3924_));
  NAND4_X1   g01442(.A1(new_n3885_), .A2(pi0241), .A3(new_n3405_), .A4(new_n3887_), .ZN(new_n3925_));
  NAND2_X1   g01443(.A1(pi0223), .A2(pi1141), .ZN(new_n3926_));
  NAND2_X1   g01444(.A1(new_n3878_), .A2(new_n3154_), .ZN(new_n3927_));
  NAND4_X1   g01445(.A1(new_n3927_), .A2(new_n2587_), .A3(new_n3875_), .A4(new_n3926_), .ZN(new_n3936_));
  NOR2_X1    g01446(.A1(new_n3847_), .A2(new_n3837_), .ZN(new_n3937_));
  AOI21_X1   g01447(.A1(new_n3897_), .A2(new_n3937_), .B(new_n3836_), .ZN(new_n3938_));
  MUX2_X1    g01448(.I0(new_n3938_), .I1(new_n3831_), .S(new_n2566_), .Z(new_n3939_));
  NOR2_X1    g01449(.A1(new_n3861_), .A2(new_n2545_), .ZN(new_n3940_));
  OAI21_X1   g01450(.A1(new_n3939_), .A2(pi0299), .B(new_n3940_), .ZN(new_n3941_));
  AOI21_X1   g01451(.A1(new_n3885_), .A2(pi0299), .B(new_n3861_), .ZN(new_n3942_));
  AOI21_X1   g01452(.A1(new_n3942_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n3943_));
  NOR3_X1    g01453(.A1(new_n3866_), .A2(pi0228), .A3(new_n3865_), .ZN(new_n3944_));
  NAND2_X1   g01454(.A1(new_n3944_), .A2(new_n3937_), .ZN(new_n3945_));
  AOI21_X1   g01455(.A1(new_n3945_), .A2(new_n3835_), .B(pi0215), .ZN(new_n3946_));
  AOI21_X1   g01456(.A1(pi0215), .A2(new_n3831_), .B(new_n3946_), .ZN(new_n3947_));
  NAND3_X1   g01457(.A1(new_n3860_), .A2(new_n3859_), .A3(new_n2587_), .ZN(new_n3948_));
  NOR2_X1    g01458(.A1(pi0038), .A2(pi0100), .ZN(new_n3949_));
  OAI21_X1   g01459(.A1(new_n3948_), .A2(pi0039), .B(new_n3949_), .ZN(new_n3950_));
  AOI21_X1   g01460(.A1(new_n3941_), .A2(new_n3943_), .B(new_n3950_), .ZN(new_n3951_));
  AOI21_X1   g01461(.A1(new_n3951_), .A2(new_n3936_), .B(pi0087), .ZN(new_n3952_));
  NOR2_X1    g01462(.A1(new_n3942_), .A2(new_n3197_), .ZN(new_n3953_));
  AOI21_X1   g01463(.A1(new_n3197_), .A2(new_n3948_), .B(new_n3953_), .ZN(new_n3954_));
  NOR2_X1    g01464(.A1(new_n3954_), .A2(new_n3177_), .ZN(new_n3955_));
  OAI21_X1   g01465(.A1(new_n3952_), .A2(pi0075), .B(new_n3955_), .ZN(new_n3956_));
  NOR4_X1    g01466(.A1(new_n3954_), .A2(pi0092), .A3(new_n2535_), .A4(new_n3942_), .ZN(new_n3957_));
  AOI21_X1   g01467(.A1(new_n3942_), .A2(new_n2539_), .B(pi0055), .ZN(new_n3958_));
  AND2_X2    g01468(.A1(new_n3942_), .A2(pi0075), .Z(new_n3959_));
  NOR4_X1    g01469(.A1(new_n3957_), .A2(new_n3330_), .A3(new_n3958_), .A4(new_n3959_), .ZN(new_n3960_));
  MUX2_X1    g01470(.I0(new_n3947_), .I1(new_n3885_), .S(new_n3336_), .Z(new_n3961_));
  NAND2_X1   g01471(.A1(new_n3947_), .A2(new_n3233_), .ZN(new_n3962_));
  AOI21_X1   g01472(.A1(new_n3885_), .A2(new_n3234_), .B(pi0055), .ZN(new_n3963_));
  AOI21_X1   g01473(.A1(new_n3962_), .A2(new_n3963_), .B(new_n3503_), .ZN(new_n3964_));
  OAI21_X1   g01474(.A1(new_n3335_), .A2(new_n3961_), .B(new_n3964_), .ZN(new_n3965_));
  AOI21_X1   g01475(.A1(new_n3956_), .A2(new_n3960_), .B(new_n3965_), .ZN(new_n3966_));
  AND2_X2    g01476(.A1(new_n3947_), .A2(new_n3343_), .Z(new_n3967_));
  OAI21_X1   g01477(.A1(new_n3343_), .A2(new_n3884_), .B(new_n3240_), .ZN(new_n3968_));
  NOR2_X1    g01478(.A1(new_n3405_), .A2(pi0241), .ZN(new_n3969_));
  OAI21_X1   g01479(.A1(new_n3967_), .A2(new_n3968_), .B(new_n3969_), .ZN(new_n3970_));
  OAI21_X1   g01480(.A1(new_n3966_), .A2(new_n3970_), .B(new_n3925_), .ZN(new_n3971_));
  AOI21_X1   g01481(.A1(new_n3920_), .A2(new_n3924_), .B(new_n3971_), .ZN(po0158));
  INV_X1     g01482(.I(pi1140), .ZN(new_n3973_));
  INV_X1     g01483(.I(pi0921), .ZN(new_n3974_));
  NOR3_X1    g01484(.A1(new_n2555_), .A2(new_n3974_), .A3(pi1140), .ZN(new_n3975_));
  AOI21_X1   g01485(.A1(new_n2554_), .A2(new_n3974_), .B(new_n3973_), .ZN(new_n3976_));
  OAI21_X1   g01486(.A1(new_n3975_), .A2(new_n3976_), .B(pi0221), .ZN(new_n3977_));
  INV_X1     g01487(.I(new_n3977_), .ZN(new_n3978_));
  AOI21_X1   g01488(.A1(pi0216), .A2(pi0282), .B(pi0221), .ZN(new_n3979_));
  MUX2_X1    g01489(.I0(new_n3428_), .I1(new_n3377_), .S(pi0869), .Z(new_n3980_));
  INV_X1     g01490(.I(pi0869), .ZN(new_n3981_));
  AOI21_X1   g01491(.A1(new_n3426_), .A2(new_n3981_), .B(pi0170), .ZN(new_n3982_));
  AOI21_X1   g01492(.A1(new_n3980_), .A2(pi0170), .B(new_n3982_), .ZN(new_n3983_));
  INV_X1     g01493(.I(pi0170), .ZN(new_n3984_));
  NOR2_X1    g01494(.A1(new_n2438_), .A2(new_n3981_), .ZN(new_n3985_));
  NAND4_X1   g01495(.A1(new_n3985_), .A2(pi0105), .A3(new_n3984_), .A4(new_n2523_), .ZN(new_n3986_));
  INV_X1     g01496(.I(new_n3986_), .ZN(new_n3987_));
  NOR2_X1    g01497(.A1(new_n3987_), .A2(pi0216), .ZN(new_n3988_));
  INV_X1     g01498(.I(new_n3988_), .ZN(new_n3989_));
  NOR2_X1    g01499(.A1(new_n3559_), .A2(new_n3989_), .ZN(new_n3990_));
  OAI21_X1   g01500(.A1(new_n3983_), .A2(pi0228), .B(new_n3990_), .ZN(new_n3991_));
  AOI21_X1   g01501(.A1(new_n3991_), .A2(new_n3979_), .B(new_n3978_), .ZN(new_n3992_));
  MUX2_X1    g01502(.I0(new_n3992_), .I1(new_n3973_), .S(pi0215), .Z(new_n3993_));
  NAND3_X1   g01503(.A1(new_n2589_), .A2(pi0921), .A3(new_n3973_), .ZN(new_n3994_));
  OAI21_X1   g01504(.A1(new_n2593_), .A2(pi0921), .B(pi1140), .ZN(new_n3995_));
  AOI21_X1   g01505(.A1(new_n3995_), .A2(new_n3994_), .B(new_n2588_), .ZN(new_n3996_));
  INV_X1     g01506(.I(new_n3996_), .ZN(new_n3997_));
  AOI21_X1   g01507(.A1(pi0224), .A2(pi0282), .B(pi0222), .ZN(new_n3998_));
  OAI21_X1   g01508(.A1(new_n3985_), .A2(pi0224), .B(new_n3998_), .ZN(new_n3999_));
  NAND2_X1   g01509(.A1(new_n3997_), .A2(new_n3999_), .ZN(new_n4000_));
  NAND3_X1   g01510(.A1(new_n4000_), .A2(new_n2604_), .A3(pi1140), .ZN(new_n4001_));
  OAI21_X1   g01511(.A1(new_n4000_), .A2(pi0223), .B(new_n3973_), .ZN(new_n4002_));
  NAND3_X1   g01512(.A1(new_n4002_), .A2(new_n4001_), .A3(new_n2587_), .ZN(new_n4003_));
  NOR2_X1    g01513(.A1(new_n4003_), .A2(new_n3297_), .ZN(new_n4004_));
  INV_X1     g01514(.I(new_n4004_), .ZN(new_n4005_));
  NOR2_X1    g01515(.A1(new_n2566_), .A2(new_n3973_), .ZN(new_n4006_));
  NOR3_X1    g01516(.A1(new_n2490_), .A2(new_n3984_), .A3(new_n3981_), .ZN(new_n4007_));
  AOI21_X1   g01517(.A1(new_n2491_), .A2(new_n3984_), .B(pi0869), .ZN(new_n4008_));
  NOR4_X1    g01518(.A1(new_n4008_), .A2(pi0228), .A3(new_n3282_), .A4(new_n4007_), .ZN(new_n4009_));
  NOR2_X1    g01519(.A1(new_n3988_), .A2(new_n3979_), .ZN(new_n4010_));
  INV_X1     g01520(.I(new_n4010_), .ZN(new_n4011_));
  OAI21_X1   g01521(.A1(new_n4009_), .A2(new_n4011_), .B(new_n3977_), .ZN(new_n4012_));
  AOI21_X1   g01522(.A1(new_n4012_), .A2(new_n2566_), .B(new_n4006_), .ZN(new_n4013_));
  AOI21_X1   g01523(.A1(new_n4013_), .A2(pi0299), .B(new_n4005_), .ZN(new_n4014_));
  OAI21_X1   g01524(.A1(new_n4014_), .A2(new_n3154_), .B(new_n3172_), .ZN(new_n4015_));
  OAI21_X1   g01525(.A1(new_n3422_), .A2(new_n3981_), .B(new_n2595_), .ZN(new_n4016_));
  AOI21_X1   g01526(.A1(new_n4016_), .A2(new_n3998_), .B(new_n3996_), .ZN(new_n4017_));
  NAND2_X1   g01527(.A1(new_n3422_), .A2(new_n3998_), .ZN(new_n4018_));
  NOR2_X1    g01528(.A1(pi0223), .A2(pi0299), .ZN(new_n4019_));
  OAI21_X1   g01529(.A1(new_n4017_), .A2(new_n4018_), .B(new_n4019_), .ZN(new_n4020_));
  INV_X1     g01530(.I(new_n4006_), .ZN(new_n4021_));
  AOI21_X1   g01531(.A1(new_n3984_), .A2(new_n2523_), .B(new_n3979_), .ZN(new_n4022_));
  NAND2_X1   g01532(.A1(new_n3988_), .A2(new_n4022_), .ZN(new_n4023_));
  NAND2_X1   g01533(.A1(new_n4023_), .A2(new_n3977_), .ZN(new_n4024_));
  NAND2_X1   g01534(.A1(new_n4024_), .A2(new_n2566_), .ZN(new_n4025_));
  NAND2_X1   g01535(.A1(new_n4025_), .A2(new_n4021_), .ZN(new_n4026_));
  INV_X1     g01536(.I(new_n4026_), .ZN(new_n4027_));
  AOI21_X1   g01537(.A1(pi0216), .A2(pi0282), .B(new_n3886_), .ZN(new_n4028_));
  NOR2_X1    g01538(.A1(new_n4027_), .A2(new_n4028_), .ZN(new_n4029_));
  INV_X1     g01539(.I(new_n4029_), .ZN(new_n4030_));
  AOI21_X1   g01540(.A1(new_n4030_), .A2(pi0299), .B(new_n4005_), .ZN(new_n4031_));
  INV_X1     g01541(.I(new_n4031_), .ZN(new_n4032_));
  OAI21_X1   g01542(.A1(new_n4032_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n4033_));
  NAND4_X1   g01543(.A1(new_n4020_), .A2(new_n3154_), .A3(new_n4015_), .A4(new_n4033_), .ZN(new_n4034_));
  AOI21_X1   g01544(.A1(new_n3993_), .A2(pi0299), .B(new_n4034_), .ZN(new_n4035_));
  NOR3_X1    g01545(.A1(new_n3257_), .A2(new_n3984_), .A3(new_n3981_), .ZN(new_n4036_));
  AOI21_X1   g01546(.A1(new_n3256_), .A2(new_n3984_), .B(pi0869), .ZN(new_n4037_));
  NOR3_X1    g01547(.A1(new_n4036_), .A2(pi0228), .A3(new_n4037_), .ZN(new_n4038_));
  NAND2_X1   g01548(.A1(new_n4038_), .A2(new_n3283_), .ZN(new_n4039_));
  AOI21_X1   g01549(.A1(new_n4039_), .A2(new_n4010_), .B(new_n3978_), .ZN(new_n4040_));
  OAI21_X1   g01550(.A1(new_n4040_), .A2(pi0215), .B(new_n4021_), .ZN(new_n4041_));
  NAND2_X1   g01551(.A1(new_n4041_), .A2(new_n2587_), .ZN(new_n4042_));
  NOR2_X1    g01552(.A1(new_n4005_), .A2(new_n2545_), .ZN(new_n4043_));
  OAI21_X1   g01553(.A1(new_n4032_), .A2(new_n2544_), .B(pi0100), .ZN(new_n4044_));
  AOI21_X1   g01554(.A1(new_n4042_), .A2(new_n4043_), .B(new_n4044_), .ZN(new_n4045_));
  OAI21_X1   g01555(.A1(new_n4035_), .A2(new_n4045_), .B(new_n3177_), .ZN(new_n4046_));
  NAND2_X1   g01556(.A1(new_n4032_), .A2(new_n3198_), .ZN(new_n4047_));
  OAI21_X1   g01557(.A1(new_n3198_), .A2(new_n4014_), .B(new_n4047_), .ZN(new_n4048_));
  NAND2_X1   g01558(.A1(new_n4048_), .A2(pi0087), .ZN(new_n4049_));
  AOI21_X1   g01559(.A1(new_n4046_), .A2(new_n2628_), .B(new_n4049_), .ZN(new_n4050_));
  NAND4_X1   g01560(.A1(new_n4048_), .A2(new_n3203_), .A3(new_n2534_), .A4(new_n4032_), .ZN(new_n4051_));
  OAI21_X1   g01561(.A1(new_n4032_), .A2(new_n2538_), .B(new_n3227_), .ZN(new_n4052_));
  NAND2_X1   g01562(.A1(new_n4031_), .A2(pi0075), .ZN(new_n4053_));
  NAND4_X1   g01563(.A1(new_n4051_), .A2(new_n3329_), .A3(new_n4052_), .A4(new_n4053_), .ZN(new_n4054_));
  INV_X1     g01564(.I(new_n4013_), .ZN(new_n4055_));
  MUX2_X1    g01565(.I0(new_n4055_), .I1(new_n4029_), .S(new_n3336_), .Z(new_n4056_));
  NOR2_X1    g01566(.A1(new_n4055_), .A2(new_n3234_), .ZN(new_n4057_));
  OAI21_X1   g01567(.A1(new_n4029_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n4058_));
  OAI21_X1   g01568(.A1(new_n4057_), .A2(new_n4058_), .B(new_n2533_), .ZN(new_n4059_));
  AOI21_X1   g01569(.A1(pi0056), .A2(new_n4056_), .B(new_n4059_), .ZN(new_n4060_));
  OAI21_X1   g01570(.A1(new_n4050_), .A2(new_n4054_), .B(new_n4060_), .ZN(new_n4061_));
  NAND2_X1   g01571(.A1(new_n4013_), .A2(new_n3343_), .ZN(new_n4062_));
  AOI21_X1   g01572(.A1(new_n4030_), .A2(new_n3400_), .B(pi0062), .ZN(new_n4063_));
  NAND2_X1   g01573(.A1(new_n2571_), .A2(pi0248), .ZN(new_n4064_));
  AOI21_X1   g01574(.A1(new_n4063_), .A2(new_n4062_), .B(new_n4064_), .ZN(new_n4065_));
  NAND4_X1   g01575(.A1(new_n4027_), .A2(pi0248), .A3(new_n3405_), .A4(new_n4028_), .ZN(new_n4066_));
  NAND2_X1   g01576(.A1(pi0223), .A2(pi1140), .ZN(new_n4067_));
  NAND2_X1   g01577(.A1(new_n4020_), .A2(new_n3154_), .ZN(new_n4068_));
  NAND4_X1   g01578(.A1(new_n4068_), .A2(new_n2587_), .A3(new_n4017_), .A4(new_n4067_), .ZN(new_n4077_));
  NOR2_X1    g01579(.A1(new_n3989_), .A2(new_n3979_), .ZN(new_n4078_));
  AOI21_X1   g01580(.A1(new_n4038_), .A2(new_n4078_), .B(new_n3978_), .ZN(new_n4079_));
  MUX2_X1    g01581(.I0(new_n4079_), .I1(new_n3973_), .S(new_n2566_), .Z(new_n4080_));
  NOR2_X1    g01582(.A1(new_n4003_), .A2(new_n2545_), .ZN(new_n4081_));
  OAI21_X1   g01583(.A1(new_n4080_), .A2(pi0299), .B(new_n4081_), .ZN(new_n4082_));
  AOI21_X1   g01584(.A1(new_n4027_), .A2(pi0299), .B(new_n4003_), .ZN(new_n4083_));
  AOI21_X1   g01585(.A1(new_n4083_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4084_));
  NOR3_X1    g01586(.A1(new_n4008_), .A2(pi0228), .A3(new_n4007_), .ZN(new_n4085_));
  NAND2_X1   g01587(.A1(new_n4085_), .A2(new_n4078_), .ZN(new_n4086_));
  AOI21_X1   g01588(.A1(new_n4086_), .A2(new_n3977_), .B(pi0215), .ZN(new_n4087_));
  AOI21_X1   g01589(.A1(pi0215), .A2(new_n3973_), .B(new_n4087_), .ZN(new_n4088_));
  NAND3_X1   g01590(.A1(new_n4002_), .A2(new_n4001_), .A3(new_n2587_), .ZN(new_n4089_));
  NOR2_X1    g01591(.A1(pi0038), .A2(pi0100), .ZN(new_n4090_));
  OAI21_X1   g01592(.A1(new_n4089_), .A2(pi0039), .B(new_n4090_), .ZN(new_n4091_));
  AOI21_X1   g01593(.A1(new_n4082_), .A2(new_n4084_), .B(new_n4091_), .ZN(new_n4092_));
  AOI21_X1   g01594(.A1(new_n4092_), .A2(new_n4077_), .B(pi0087), .ZN(new_n4093_));
  NOR2_X1    g01595(.A1(new_n4083_), .A2(new_n3197_), .ZN(new_n4094_));
  AOI21_X1   g01596(.A1(new_n3197_), .A2(new_n4089_), .B(new_n4094_), .ZN(new_n4095_));
  NOR2_X1    g01597(.A1(new_n4095_), .A2(new_n3177_), .ZN(new_n4096_));
  OAI21_X1   g01598(.A1(new_n4093_), .A2(pi0075), .B(new_n4096_), .ZN(new_n4097_));
  NOR4_X1    g01599(.A1(new_n4095_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4083_), .ZN(new_n4098_));
  AOI21_X1   g01600(.A1(new_n4083_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4099_));
  AND2_X2    g01601(.A1(new_n4083_), .A2(pi0075), .Z(new_n4100_));
  NOR4_X1    g01602(.A1(new_n4098_), .A2(new_n3330_), .A3(new_n4099_), .A4(new_n4100_), .ZN(new_n4101_));
  MUX2_X1    g01603(.I0(new_n4088_), .I1(new_n4027_), .S(new_n3336_), .Z(new_n4102_));
  NAND2_X1   g01604(.A1(new_n4088_), .A2(new_n3233_), .ZN(new_n4103_));
  AOI21_X1   g01605(.A1(new_n4027_), .A2(new_n3234_), .B(pi0055), .ZN(new_n4104_));
  AOI21_X1   g01606(.A1(new_n4103_), .A2(new_n4104_), .B(new_n3503_), .ZN(new_n4105_));
  OAI21_X1   g01607(.A1(new_n3335_), .A2(new_n4102_), .B(new_n4105_), .ZN(new_n4106_));
  AOI21_X1   g01608(.A1(new_n4097_), .A2(new_n4101_), .B(new_n4106_), .ZN(new_n4107_));
  AND2_X2    g01609(.A1(new_n4088_), .A2(new_n3343_), .Z(new_n4108_));
  OAI21_X1   g01610(.A1(new_n3343_), .A2(new_n4026_), .B(new_n3240_), .ZN(new_n4109_));
  NOR2_X1    g01611(.A1(new_n3405_), .A2(pi0248), .ZN(new_n4110_));
  OAI21_X1   g01612(.A1(new_n4108_), .A2(new_n4109_), .B(new_n4110_), .ZN(new_n4111_));
  OAI21_X1   g01613(.A1(new_n4107_), .A2(new_n4111_), .B(new_n4066_), .ZN(new_n4112_));
  AOI21_X1   g01614(.A1(new_n4061_), .A2(new_n4065_), .B(new_n4112_), .ZN(po0159));
  INV_X1     g01615(.I(pi0862), .ZN(new_n4114_));
  INV_X1     g01616(.I(pi1139), .ZN(new_n4115_));
  NAND3_X1   g01617(.A1(new_n2589_), .A2(pi0920), .A3(new_n4115_), .ZN(new_n4116_));
  OAI21_X1   g01618(.A1(new_n2593_), .A2(pi0920), .B(pi1139), .ZN(new_n4117_));
  AOI21_X1   g01619(.A1(new_n4117_), .A2(new_n4116_), .B(new_n2588_), .ZN(new_n4118_));
  INV_X1     g01620(.I(pi0281), .ZN(new_n4119_));
  NOR2_X1    g01621(.A1(new_n2595_), .A2(new_n4119_), .ZN(new_n4120_));
  OAI21_X1   g01622(.A1(new_n4120_), .A2(pi0222), .B(new_n2604_), .ZN(new_n4121_));
  OAI22_X1   g01623(.A1(new_n4118_), .A2(new_n4121_), .B1(new_n2604_), .B2(pi1139), .ZN(new_n4122_));
  NOR2_X1    g01624(.A1(new_n4122_), .A2(pi0299), .ZN(new_n4123_));
  INV_X1     g01625(.I(new_n4123_), .ZN(new_n4124_));
  NOR2_X1    g01626(.A1(new_n2604_), .A2(new_n4115_), .ZN(new_n4125_));
  NOR3_X1    g01627(.A1(new_n4118_), .A2(pi0224), .A3(new_n4125_), .ZN(new_n4126_));
  INV_X1     g01628(.I(new_n4126_), .ZN(new_n4127_));
  NAND3_X1   g01629(.A1(new_n4124_), .A2(new_n4114_), .A3(new_n4127_), .ZN(new_n4128_));
  NOR2_X1    g01630(.A1(new_n3422_), .A2(new_n4128_), .ZN(new_n4129_));
  INV_X1     g01631(.I(pi0148), .ZN(new_n4130_));
  NOR2_X1    g01632(.A1(new_n4130_), .A2(pi0215), .ZN(new_n4131_));
  OAI21_X1   g01633(.A1(pi0833), .A2(pi1139), .B(pi0920), .ZN(new_n4132_));
  NOR3_X1    g01634(.A1(new_n4115_), .A2(pi0833), .A3(pi0920), .ZN(new_n4133_));
  INV_X1     g01635(.I(new_n4133_), .ZN(new_n4134_));
  NOR2_X1    g01636(.A1(new_n2550_), .A2(pi0216), .ZN(new_n4135_));
  AND3_X2    g01637(.A1(new_n4134_), .A2(new_n4132_), .A3(new_n4135_), .Z(new_n4136_));
  INV_X1     g01638(.I(new_n4136_), .ZN(new_n4137_));
  AOI21_X1   g01639(.A1(pi0216), .A2(new_n4115_), .B(new_n4137_), .ZN(new_n4138_));
  NOR2_X1    g01640(.A1(new_n2523_), .A2(pi0105), .ZN(new_n4139_));
  AOI21_X1   g01641(.A1(new_n3376_), .A2(new_n2523_), .B(new_n4139_), .ZN(new_n4140_));
  NOR3_X1    g01642(.A1(new_n4140_), .A2(pi0862), .A3(new_n3432_), .ZN(new_n4141_));
  INV_X1     g01643(.I(new_n4140_), .ZN(new_n4142_));
  AOI21_X1   g01644(.A1(new_n4114_), .A2(new_n3432_), .B(new_n4142_), .ZN(new_n4143_));
  AOI21_X1   g01645(.A1(pi0216), .A2(pi0281), .B(pi0221), .ZN(new_n4144_));
  INV_X1     g01646(.I(new_n4144_), .ZN(new_n4145_));
  NOR4_X1    g01647(.A1(new_n4143_), .A2(pi0216), .A3(new_n4141_), .A4(new_n4145_), .ZN(new_n4146_));
  OAI21_X1   g01648(.A1(new_n4146_), .A2(new_n4138_), .B(new_n4131_), .ZN(new_n4147_));
  NOR2_X1    g01649(.A1(pi0148), .A2(pi0215), .ZN(new_n4148_));
  INV_X1     g01650(.I(new_n4148_), .ZN(new_n4149_));
  INV_X1     g01651(.I(new_n4138_), .ZN(new_n4150_));
  NOR3_X1    g01652(.A1(new_n4144_), .A2(pi0216), .A3(pi0862), .ZN(new_n4151_));
  INV_X1     g01653(.I(new_n4151_), .ZN(new_n4152_));
  OAI21_X1   g01654(.A1(new_n3427_), .A2(new_n4152_), .B(new_n4150_), .ZN(new_n4153_));
  NOR2_X1    g01655(.A1(new_n4153_), .A2(new_n4149_), .ZN(new_n4154_));
  NOR2_X1    g01656(.A1(new_n2566_), .A2(new_n4115_), .ZN(new_n4155_));
  NOR3_X1    g01657(.A1(new_n4154_), .A2(pi0299), .A3(new_n4155_), .ZN(new_n4156_));
  AOI21_X1   g01658(.A1(new_n4147_), .A2(new_n4156_), .B(new_n4129_), .ZN(new_n4157_));
  INV_X1     g01659(.I(new_n3297_), .ZN(new_n4158_));
  NAND2_X1   g01660(.A1(new_n4128_), .A2(new_n4158_), .ZN(new_n4159_));
  INV_X1     g01661(.I(new_n4155_), .ZN(new_n4160_));
  NOR2_X1    g01662(.A1(new_n3310_), .A2(new_n3461_), .ZN(new_n4161_));
  OAI21_X1   g01663(.A1(new_n4161_), .A2(new_n4152_), .B(new_n4150_), .ZN(new_n4162_));
  INV_X1     g01664(.I(new_n4162_), .ZN(new_n4163_));
  NOR2_X1    g01665(.A1(new_n4136_), .A2(pi0216), .ZN(new_n4164_));
  INV_X1     g01666(.I(new_n4164_), .ZN(new_n4165_));
  NOR3_X1    g01667(.A1(new_n3310_), .A2(new_n3461_), .A3(new_n4165_), .ZN(new_n4166_));
  OAI22_X1   g01668(.A1(new_n4162_), .A2(new_n4166_), .B1(new_n4130_), .B2(pi0215), .ZN(new_n4167_));
  NAND2_X1   g01669(.A1(new_n2525_), .A2(pi0148), .ZN(new_n4168_));
  OAI21_X1   g01670(.A1(new_n4165_), .A2(new_n4168_), .B(new_n2566_), .ZN(new_n4169_));
  AOI22_X1   g01671(.A1(new_n4167_), .A2(new_n4160_), .B1(new_n4163_), .B2(new_n4169_), .ZN(new_n4170_));
  OAI21_X1   g01672(.A1(new_n4170_), .A2(new_n2587_), .B(new_n4159_), .ZN(new_n4171_));
  MUX2_X1    g01673(.I0(new_n4171_), .I1(new_n4157_), .S(new_n3154_), .Z(new_n4172_));
  AOI21_X1   g01674(.A1(new_n3471_), .A2(new_n4144_), .B(new_n4163_), .ZN(new_n4173_));
  NOR2_X1    g01675(.A1(new_n4173_), .A2(new_n4149_), .ZN(new_n4174_));
  INV_X1     g01676(.I(new_n3470_), .ZN(new_n4175_));
  NOR4_X1    g01677(.A1(new_n4162_), .A2(pi0216), .A3(new_n2524_), .A4(new_n4138_), .ZN(new_n4176_));
  AOI21_X1   g01678(.A1(new_n4175_), .A2(new_n4176_), .B(new_n4131_), .ZN(new_n4177_));
  OAI21_X1   g01679(.A1(new_n4177_), .A2(new_n4155_), .B(new_n2587_), .ZN(new_n4178_));
  INV_X1     g01680(.I(new_n4159_), .ZN(new_n4179_));
  NOR2_X1    g01681(.A1(new_n4179_), .A2(new_n2545_), .ZN(new_n4180_));
  OAI21_X1   g01682(.A1(new_n4174_), .A2(new_n4178_), .B(new_n4180_), .ZN(new_n4181_));
  NOR3_X1    g01683(.A1(new_n4152_), .A2(new_n2438_), .A3(new_n2525_), .ZN(new_n4182_));
  OAI21_X1   g01684(.A1(new_n4138_), .A2(new_n4182_), .B(new_n4169_), .ZN(new_n4183_));
  NAND2_X1   g01685(.A1(new_n4183_), .A2(new_n4160_), .ZN(new_n4184_));
  INV_X1     g01686(.I(new_n4184_), .ZN(new_n4185_));
  AOI21_X1   g01687(.A1(new_n4185_), .A2(pi0299), .B(new_n4179_), .ZN(new_n4186_));
  AOI21_X1   g01688(.A1(new_n4186_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4187_));
  INV_X1     g01689(.I(new_n4186_), .ZN(new_n4188_));
  OAI21_X1   g01690(.A1(new_n4188_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n4189_));
  AOI21_X1   g01691(.A1(new_n4181_), .A2(new_n4187_), .B(new_n4189_), .ZN(new_n4190_));
  OAI21_X1   g01692(.A1(new_n4172_), .A2(pi0038), .B(new_n4190_), .ZN(new_n4191_));
  AOI21_X1   g01693(.A1(new_n4191_), .A2(new_n3177_), .B(pi0075), .ZN(new_n4192_));
  NOR2_X1    g01694(.A1(new_n4186_), .A2(new_n3197_), .ZN(new_n4193_));
  AOI21_X1   g01695(.A1(new_n4171_), .A2(new_n3197_), .B(new_n4193_), .ZN(new_n4194_));
  OR2_X2     g01696(.A1(new_n4194_), .A2(new_n3177_), .Z(new_n4195_));
  NOR4_X1    g01697(.A1(new_n4194_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4186_), .ZN(new_n4196_));
  AOI21_X1   g01698(.A1(new_n4186_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4197_));
  NOR2_X1    g01699(.A1(new_n4188_), .A2(new_n2628_), .ZN(new_n4198_));
  NOR4_X1    g01700(.A1(new_n4196_), .A2(new_n3330_), .A3(new_n4197_), .A4(new_n4198_), .ZN(new_n4199_));
  OAI21_X1   g01701(.A1(new_n4192_), .A2(new_n4195_), .B(new_n4199_), .ZN(new_n4200_));
  MUX2_X1    g01702(.I0(new_n4170_), .I1(new_n4184_), .S(new_n3336_), .Z(new_n4201_));
  NOR2_X1    g01703(.A1(new_n4170_), .A2(new_n3234_), .ZN(new_n4202_));
  OAI21_X1   g01704(.A1(new_n4184_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n4203_));
  OAI21_X1   g01705(.A1(new_n4202_), .A2(new_n4203_), .B(new_n2533_), .ZN(new_n4204_));
  AOI21_X1   g01706(.A1(pi0056), .A2(new_n4201_), .B(new_n4204_), .ZN(new_n4205_));
  NOR2_X1    g01707(.A1(new_n4170_), .A2(new_n3400_), .ZN(new_n4206_));
  OAI21_X1   g01708(.A1(new_n3343_), .A2(new_n4184_), .B(new_n3240_), .ZN(new_n4207_));
  OAI21_X1   g01709(.A1(new_n4206_), .A2(new_n4207_), .B(new_n2571_), .ZN(new_n4208_));
  AOI21_X1   g01710(.A1(new_n4200_), .A2(new_n4205_), .B(new_n4208_), .ZN(new_n4209_));
  OAI21_X1   g01711(.A1(new_n4185_), .A2(new_n2571_), .B(pi0247), .ZN(new_n4210_));
  NOR3_X1    g01712(.A1(new_n4140_), .A2(pi0862), .A3(new_n3432_), .ZN(new_n4211_));
  OAI21_X1   g01713(.A1(new_n4142_), .A2(pi0862), .B(new_n3432_), .ZN(new_n4212_));
  NAND3_X1   g01714(.A1(new_n4212_), .A2(new_n2562_), .A3(new_n4144_), .ZN(new_n4213_));
  OAI21_X1   g01715(.A1(new_n4213_), .A2(new_n4211_), .B(new_n4150_), .ZN(new_n4214_));
  NOR2_X1    g01716(.A1(new_n4165_), .A2(new_n4131_), .ZN(new_n4215_));
  NAND2_X1   g01717(.A1(new_n3427_), .A2(new_n4215_), .ZN(new_n4216_));
  NOR2_X1    g01718(.A1(new_n4155_), .A2(new_n2587_), .ZN(new_n4217_));
  OAI21_X1   g01719(.A1(new_n4153_), .A2(new_n4216_), .B(new_n4217_), .ZN(new_n4218_));
  AOI21_X1   g01720(.A1(new_n4214_), .A2(new_n4148_), .B(new_n4218_), .ZN(new_n4219_));
  NOR2_X1    g01721(.A1(new_n4127_), .A2(new_n4114_), .ZN(new_n4220_));
  AOI21_X1   g01722(.A1(new_n3421_), .A2(new_n4220_), .B(new_n4124_), .ZN(new_n4221_));
  OAI21_X1   g01723(.A1(new_n4219_), .A2(pi0039), .B(new_n4221_), .ZN(new_n4222_));
  NOR4_X1    g01724(.A1(new_n4173_), .A2(new_n3472_), .A3(new_n4131_), .A4(new_n4165_), .ZN(new_n4223_));
  NAND2_X1   g01725(.A1(new_n4175_), .A2(new_n2525_), .ZN(new_n4224_));
  NOR2_X1    g01726(.A1(new_n3310_), .A2(new_n2524_), .ZN(new_n4225_));
  AOI21_X1   g01727(.A1(new_n3283_), .A2(pi0862), .B(pi0216), .ZN(new_n4226_));
  INV_X1     g01728(.I(new_n4226_), .ZN(new_n4227_));
  OAI21_X1   g01729(.A1(new_n4225_), .A2(new_n4227_), .B(new_n4144_), .ZN(new_n4228_));
  NAND2_X1   g01730(.A1(new_n4228_), .A2(new_n4150_), .ZN(new_n4229_));
  NAND4_X1   g01731(.A1(new_n4224_), .A2(new_n4145_), .A3(new_n4149_), .A4(new_n4229_), .ZN(new_n4230_));
  NAND2_X1   g01732(.A1(new_n4230_), .A2(new_n4160_), .ZN(new_n4231_));
  NOR4_X1    g01733(.A1(new_n4123_), .A2(new_n4114_), .A3(new_n2438_), .A4(new_n4127_), .ZN(new_n4232_));
  NOR2_X1    g01734(.A1(new_n4232_), .A2(new_n3671_), .ZN(new_n4233_));
  OAI21_X1   g01735(.A1(new_n4231_), .A2(new_n4223_), .B(new_n4233_), .ZN(new_n4234_));
  NOR2_X1    g01736(.A1(new_n4184_), .A2(new_n3288_), .ZN(new_n4235_));
  AOI21_X1   g01737(.A1(new_n4235_), .A2(pi0299), .B(new_n4232_), .ZN(new_n4236_));
  AOI21_X1   g01738(.A1(new_n4236_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4237_));
  INV_X1     g01739(.I(new_n4232_), .ZN(new_n4238_));
  AOI22_X1   g01740(.A1(new_n4167_), .A2(new_n4160_), .B1(new_n4229_), .B2(new_n4148_), .ZN(new_n4239_));
  OAI21_X1   g01741(.A1(new_n4239_), .A2(new_n2587_), .B(new_n4238_), .ZN(new_n4240_));
  NOR2_X1    g01742(.A1(pi0038), .A2(pi0100), .ZN(new_n4241_));
  OAI21_X1   g01743(.A1(new_n4240_), .A2(pi0039), .B(new_n4241_), .ZN(new_n4242_));
  AOI21_X1   g01744(.A1(new_n4234_), .A2(new_n4237_), .B(new_n4242_), .ZN(new_n4243_));
  AOI21_X1   g01745(.A1(new_n4222_), .A2(new_n4243_), .B(pi0087), .ZN(new_n4244_));
  NOR2_X1    g01746(.A1(new_n4236_), .A2(new_n3197_), .ZN(new_n4245_));
  AOI21_X1   g01747(.A1(new_n4240_), .A2(new_n3197_), .B(new_n4245_), .ZN(new_n4246_));
  NOR2_X1    g01748(.A1(new_n4246_), .A2(new_n3177_), .ZN(new_n4247_));
  OAI21_X1   g01749(.A1(new_n4244_), .A2(pi0075), .B(new_n4247_), .ZN(new_n4248_));
  NOR4_X1    g01750(.A1(new_n4246_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4236_), .ZN(new_n4249_));
  AOI21_X1   g01751(.A1(new_n4236_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4250_));
  AND2_X2    g01752(.A1(new_n4236_), .A2(pi0075), .Z(new_n4251_));
  NOR4_X1    g01753(.A1(new_n4249_), .A2(new_n3330_), .A3(new_n4250_), .A4(new_n4251_), .ZN(new_n4252_));
  INV_X1     g01754(.I(new_n4235_), .ZN(new_n4253_));
  NAND4_X1   g01755(.A1(new_n4239_), .A2(new_n3335_), .A3(new_n2548_), .A4(new_n4253_), .ZN(new_n4254_));
  NAND2_X1   g01756(.A1(new_n4254_), .A2(new_n2533_), .ZN(new_n4255_));
  AOI21_X1   g01757(.A1(new_n4248_), .A2(new_n4252_), .B(new_n4255_), .ZN(new_n4256_));
  NOR2_X1    g01758(.A1(new_n4256_), .A2(new_n3405_), .ZN(new_n4257_));
  INV_X1     g01759(.I(pi0247), .ZN(new_n4258_));
  OAI21_X1   g01760(.A1(new_n4235_), .A2(new_n2571_), .B(new_n4258_), .ZN(new_n4259_));
  OAI22_X1   g01761(.A1(new_n4209_), .A2(new_n4210_), .B1(new_n4257_), .B2(new_n4259_), .ZN(po0160));
  INV_X1     g01762(.I(pi1138), .ZN(new_n4261_));
  INV_X1     g01763(.I(pi0940), .ZN(new_n4262_));
  NOR3_X1    g01764(.A1(new_n2555_), .A2(new_n4262_), .A3(pi1138), .ZN(new_n4263_));
  AOI21_X1   g01765(.A1(new_n2554_), .A2(new_n4262_), .B(new_n4261_), .ZN(new_n4264_));
  OAI21_X1   g01766(.A1(new_n4263_), .A2(new_n4264_), .B(pi0221), .ZN(new_n4265_));
  INV_X1     g01767(.I(new_n4265_), .ZN(new_n4266_));
  AOI21_X1   g01768(.A1(pi0216), .A2(pi0269), .B(pi0221), .ZN(new_n4267_));
  MUX2_X1    g01769(.I0(new_n3428_), .I1(new_n3377_), .S(pi0877), .Z(new_n4268_));
  INV_X1     g01770(.I(pi0877), .ZN(new_n4269_));
  AOI21_X1   g01771(.A1(new_n3426_), .A2(new_n4269_), .B(pi0169), .ZN(new_n4270_));
  AOI21_X1   g01772(.A1(new_n4268_), .A2(pi0169), .B(new_n4270_), .ZN(new_n4271_));
  INV_X1     g01773(.I(pi0169), .ZN(new_n4272_));
  NOR2_X1    g01774(.A1(new_n2438_), .A2(new_n4269_), .ZN(new_n4273_));
  NAND4_X1   g01775(.A1(new_n4273_), .A2(pi0105), .A3(new_n4272_), .A4(new_n2523_), .ZN(new_n4274_));
  INV_X1     g01776(.I(new_n4274_), .ZN(new_n4275_));
  NOR2_X1    g01777(.A1(new_n4275_), .A2(pi0216), .ZN(new_n4276_));
  INV_X1     g01778(.I(new_n4276_), .ZN(new_n4277_));
  NOR2_X1    g01779(.A1(new_n3559_), .A2(new_n4277_), .ZN(new_n4278_));
  OAI21_X1   g01780(.A1(new_n4271_), .A2(pi0228), .B(new_n4278_), .ZN(new_n4279_));
  AOI21_X1   g01781(.A1(new_n4279_), .A2(new_n4267_), .B(new_n4266_), .ZN(new_n4280_));
  MUX2_X1    g01782(.I0(new_n4280_), .I1(new_n4261_), .S(pi0215), .Z(new_n4281_));
  NAND3_X1   g01783(.A1(new_n2589_), .A2(pi0940), .A3(new_n4261_), .ZN(new_n4282_));
  OAI21_X1   g01784(.A1(new_n2593_), .A2(pi0940), .B(pi1138), .ZN(new_n4283_));
  AOI21_X1   g01785(.A1(new_n4283_), .A2(new_n4282_), .B(new_n2588_), .ZN(new_n4284_));
  INV_X1     g01786(.I(new_n4284_), .ZN(new_n4285_));
  AOI21_X1   g01787(.A1(pi0224), .A2(pi0269), .B(pi0222), .ZN(new_n4286_));
  OAI21_X1   g01788(.A1(new_n4273_), .A2(pi0224), .B(new_n4286_), .ZN(new_n4287_));
  NAND2_X1   g01789(.A1(new_n4285_), .A2(new_n4287_), .ZN(new_n4288_));
  NAND3_X1   g01790(.A1(new_n4288_), .A2(new_n2604_), .A3(pi1138), .ZN(new_n4289_));
  OAI21_X1   g01791(.A1(new_n4288_), .A2(pi0223), .B(new_n4261_), .ZN(new_n4290_));
  NAND3_X1   g01792(.A1(new_n4290_), .A2(new_n4289_), .A3(new_n2587_), .ZN(new_n4291_));
  NOR2_X1    g01793(.A1(new_n4291_), .A2(new_n3297_), .ZN(new_n4292_));
  INV_X1     g01794(.I(new_n4292_), .ZN(new_n4293_));
  NOR2_X1    g01795(.A1(new_n2566_), .A2(new_n4261_), .ZN(new_n4294_));
  NOR3_X1    g01796(.A1(new_n2490_), .A2(new_n4272_), .A3(new_n4269_), .ZN(new_n4295_));
  AOI21_X1   g01797(.A1(new_n2491_), .A2(new_n4272_), .B(pi0877), .ZN(new_n4296_));
  NOR4_X1    g01798(.A1(new_n4296_), .A2(pi0228), .A3(new_n3282_), .A4(new_n4295_), .ZN(new_n4297_));
  NOR2_X1    g01799(.A1(new_n4276_), .A2(new_n4267_), .ZN(new_n4298_));
  INV_X1     g01800(.I(new_n4298_), .ZN(new_n4299_));
  OAI21_X1   g01801(.A1(new_n4297_), .A2(new_n4299_), .B(new_n4265_), .ZN(new_n4300_));
  AOI21_X1   g01802(.A1(new_n4300_), .A2(new_n2566_), .B(new_n4294_), .ZN(new_n4301_));
  AOI21_X1   g01803(.A1(new_n4301_), .A2(pi0299), .B(new_n4293_), .ZN(new_n4302_));
  OAI21_X1   g01804(.A1(new_n4302_), .A2(new_n3154_), .B(new_n3172_), .ZN(new_n4303_));
  OAI21_X1   g01805(.A1(new_n3422_), .A2(new_n4269_), .B(new_n2595_), .ZN(new_n4304_));
  AOI21_X1   g01806(.A1(new_n4304_), .A2(new_n4286_), .B(new_n4284_), .ZN(new_n4305_));
  NAND2_X1   g01807(.A1(new_n3422_), .A2(new_n4286_), .ZN(new_n4306_));
  NOR2_X1    g01808(.A1(pi0223), .A2(pi0299), .ZN(new_n4307_));
  OAI21_X1   g01809(.A1(new_n4305_), .A2(new_n4306_), .B(new_n4307_), .ZN(new_n4308_));
  INV_X1     g01810(.I(new_n4294_), .ZN(new_n4309_));
  AOI21_X1   g01811(.A1(new_n4272_), .A2(new_n2523_), .B(new_n4267_), .ZN(new_n4310_));
  NAND2_X1   g01812(.A1(new_n4276_), .A2(new_n4310_), .ZN(new_n4311_));
  NAND2_X1   g01813(.A1(new_n4311_), .A2(new_n4265_), .ZN(new_n4312_));
  NAND2_X1   g01814(.A1(new_n4312_), .A2(new_n2566_), .ZN(new_n4313_));
  NAND2_X1   g01815(.A1(new_n4313_), .A2(new_n4309_), .ZN(new_n4314_));
  INV_X1     g01816(.I(new_n4314_), .ZN(new_n4315_));
  AOI21_X1   g01817(.A1(pi0216), .A2(pi0269), .B(new_n3886_), .ZN(new_n4316_));
  NOR2_X1    g01818(.A1(new_n4315_), .A2(new_n4316_), .ZN(new_n4317_));
  INV_X1     g01819(.I(new_n4317_), .ZN(new_n4318_));
  AOI21_X1   g01820(.A1(new_n4318_), .A2(pi0299), .B(new_n4293_), .ZN(new_n4319_));
  INV_X1     g01821(.I(new_n4319_), .ZN(new_n4320_));
  OAI21_X1   g01822(.A1(new_n4320_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n4321_));
  NAND4_X1   g01823(.A1(new_n4308_), .A2(new_n3154_), .A3(new_n4303_), .A4(new_n4321_), .ZN(new_n4322_));
  AOI21_X1   g01824(.A1(new_n4281_), .A2(pi0299), .B(new_n4322_), .ZN(new_n4323_));
  NOR3_X1    g01825(.A1(new_n3257_), .A2(new_n4272_), .A3(new_n4269_), .ZN(new_n4324_));
  AOI21_X1   g01826(.A1(new_n3256_), .A2(new_n4272_), .B(pi0877), .ZN(new_n4325_));
  NOR3_X1    g01827(.A1(new_n4324_), .A2(pi0228), .A3(new_n4325_), .ZN(new_n4326_));
  NAND2_X1   g01828(.A1(new_n4326_), .A2(new_n3283_), .ZN(new_n4327_));
  AOI21_X1   g01829(.A1(new_n4327_), .A2(new_n4298_), .B(new_n4266_), .ZN(new_n4328_));
  OAI21_X1   g01830(.A1(new_n4328_), .A2(pi0215), .B(new_n4309_), .ZN(new_n4329_));
  NAND2_X1   g01831(.A1(new_n4329_), .A2(new_n2587_), .ZN(new_n4330_));
  NOR2_X1    g01832(.A1(new_n4293_), .A2(new_n2545_), .ZN(new_n4331_));
  OAI21_X1   g01833(.A1(new_n4320_), .A2(new_n2544_), .B(pi0100), .ZN(new_n4332_));
  AOI21_X1   g01834(.A1(new_n4330_), .A2(new_n4331_), .B(new_n4332_), .ZN(new_n4333_));
  OAI21_X1   g01835(.A1(new_n4323_), .A2(new_n4333_), .B(new_n3177_), .ZN(new_n4334_));
  NAND2_X1   g01836(.A1(new_n4320_), .A2(new_n3198_), .ZN(new_n4335_));
  OAI21_X1   g01837(.A1(new_n3198_), .A2(new_n4302_), .B(new_n4335_), .ZN(new_n4336_));
  NAND2_X1   g01838(.A1(new_n4336_), .A2(pi0087), .ZN(new_n4337_));
  AOI21_X1   g01839(.A1(new_n4334_), .A2(new_n2628_), .B(new_n4337_), .ZN(new_n4338_));
  NAND4_X1   g01840(.A1(new_n4336_), .A2(new_n3203_), .A3(new_n2534_), .A4(new_n4320_), .ZN(new_n4339_));
  OAI21_X1   g01841(.A1(new_n4320_), .A2(new_n2538_), .B(new_n3227_), .ZN(new_n4340_));
  NAND2_X1   g01842(.A1(new_n4319_), .A2(pi0075), .ZN(new_n4341_));
  NAND4_X1   g01843(.A1(new_n4339_), .A2(new_n3329_), .A3(new_n4340_), .A4(new_n4341_), .ZN(new_n4342_));
  INV_X1     g01844(.I(new_n4301_), .ZN(new_n4343_));
  MUX2_X1    g01845(.I0(new_n4343_), .I1(new_n4317_), .S(new_n3336_), .Z(new_n4344_));
  NOR2_X1    g01846(.A1(new_n4343_), .A2(new_n3234_), .ZN(new_n4345_));
  OAI21_X1   g01847(.A1(new_n4317_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n4346_));
  OAI21_X1   g01848(.A1(new_n4345_), .A2(new_n4346_), .B(new_n2533_), .ZN(new_n4347_));
  AOI21_X1   g01849(.A1(pi0056), .A2(new_n4344_), .B(new_n4347_), .ZN(new_n4348_));
  OAI21_X1   g01850(.A1(new_n4338_), .A2(new_n4342_), .B(new_n4348_), .ZN(new_n4349_));
  NAND2_X1   g01851(.A1(new_n4301_), .A2(new_n3343_), .ZN(new_n4350_));
  AOI21_X1   g01852(.A1(new_n4318_), .A2(new_n3400_), .B(pi0062), .ZN(new_n4351_));
  NAND2_X1   g01853(.A1(new_n2571_), .A2(pi0246), .ZN(new_n4352_));
  AOI21_X1   g01854(.A1(new_n4351_), .A2(new_n4350_), .B(new_n4352_), .ZN(new_n4353_));
  NAND4_X1   g01855(.A1(new_n4315_), .A2(pi0246), .A3(new_n3405_), .A4(new_n4316_), .ZN(new_n4354_));
  NAND2_X1   g01856(.A1(pi0223), .A2(pi1138), .ZN(new_n4355_));
  NAND2_X1   g01857(.A1(new_n4308_), .A2(new_n3154_), .ZN(new_n4356_));
  NAND4_X1   g01858(.A1(new_n4356_), .A2(new_n2587_), .A3(new_n4305_), .A4(new_n4355_), .ZN(new_n4365_));
  NOR2_X1    g01859(.A1(new_n4277_), .A2(new_n4267_), .ZN(new_n4366_));
  AOI21_X1   g01860(.A1(new_n4326_), .A2(new_n4366_), .B(new_n4266_), .ZN(new_n4367_));
  MUX2_X1    g01861(.I0(new_n4367_), .I1(new_n4261_), .S(new_n2566_), .Z(new_n4368_));
  NOR2_X1    g01862(.A1(new_n4291_), .A2(new_n2545_), .ZN(new_n4369_));
  OAI21_X1   g01863(.A1(new_n4368_), .A2(pi0299), .B(new_n4369_), .ZN(new_n4370_));
  AOI21_X1   g01864(.A1(new_n4315_), .A2(pi0299), .B(new_n4291_), .ZN(new_n4371_));
  AOI21_X1   g01865(.A1(new_n4371_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4372_));
  NOR3_X1    g01866(.A1(new_n4296_), .A2(pi0228), .A3(new_n4295_), .ZN(new_n4373_));
  NAND2_X1   g01867(.A1(new_n4373_), .A2(new_n4366_), .ZN(new_n4374_));
  AOI21_X1   g01868(.A1(new_n4374_), .A2(new_n4265_), .B(pi0215), .ZN(new_n4375_));
  AOI21_X1   g01869(.A1(pi0215), .A2(new_n4261_), .B(new_n4375_), .ZN(new_n4376_));
  NAND3_X1   g01870(.A1(new_n4290_), .A2(new_n4289_), .A3(new_n2587_), .ZN(new_n4377_));
  NOR2_X1    g01871(.A1(pi0038), .A2(pi0100), .ZN(new_n4378_));
  OAI21_X1   g01872(.A1(new_n4377_), .A2(pi0039), .B(new_n4378_), .ZN(new_n4379_));
  AOI21_X1   g01873(.A1(new_n4370_), .A2(new_n4372_), .B(new_n4379_), .ZN(new_n4380_));
  AOI21_X1   g01874(.A1(new_n4380_), .A2(new_n4365_), .B(pi0087), .ZN(new_n4381_));
  NOR2_X1    g01875(.A1(new_n4371_), .A2(new_n3197_), .ZN(new_n4382_));
  AOI21_X1   g01876(.A1(new_n3197_), .A2(new_n4377_), .B(new_n4382_), .ZN(new_n4383_));
  NOR2_X1    g01877(.A1(new_n4383_), .A2(new_n3177_), .ZN(new_n4384_));
  OAI21_X1   g01878(.A1(new_n4381_), .A2(pi0075), .B(new_n4384_), .ZN(new_n4385_));
  NOR4_X1    g01879(.A1(new_n4383_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4371_), .ZN(new_n4386_));
  AOI21_X1   g01880(.A1(new_n4371_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4387_));
  AND2_X2    g01881(.A1(new_n4371_), .A2(pi0075), .Z(new_n4388_));
  NOR4_X1    g01882(.A1(new_n4386_), .A2(new_n3330_), .A3(new_n4387_), .A4(new_n4388_), .ZN(new_n4389_));
  MUX2_X1    g01883(.I0(new_n4376_), .I1(new_n4315_), .S(new_n3336_), .Z(new_n4390_));
  NAND2_X1   g01884(.A1(new_n4376_), .A2(new_n3233_), .ZN(new_n4391_));
  AOI21_X1   g01885(.A1(new_n4315_), .A2(new_n3234_), .B(pi0055), .ZN(new_n4392_));
  AOI21_X1   g01886(.A1(new_n4391_), .A2(new_n4392_), .B(new_n3503_), .ZN(new_n4393_));
  OAI21_X1   g01887(.A1(new_n3335_), .A2(new_n4390_), .B(new_n4393_), .ZN(new_n4394_));
  AOI21_X1   g01888(.A1(new_n4385_), .A2(new_n4389_), .B(new_n4394_), .ZN(new_n4395_));
  AND2_X2    g01889(.A1(new_n4376_), .A2(new_n3343_), .Z(new_n4396_));
  OAI21_X1   g01890(.A1(new_n3343_), .A2(new_n4314_), .B(new_n3240_), .ZN(new_n4397_));
  NOR2_X1    g01891(.A1(new_n3405_), .A2(pi0246), .ZN(new_n4398_));
  OAI21_X1   g01892(.A1(new_n4396_), .A2(new_n4397_), .B(new_n4398_), .ZN(new_n4399_));
  OAI21_X1   g01893(.A1(new_n4395_), .A2(new_n4399_), .B(new_n4354_), .ZN(new_n4400_));
  AOI21_X1   g01894(.A1(new_n4349_), .A2(new_n4353_), .B(new_n4400_), .ZN(po0161));
  INV_X1     g01895(.I(pi1137), .ZN(new_n4402_));
  INV_X1     g01896(.I(pi0933), .ZN(new_n4403_));
  NOR3_X1    g01897(.A1(new_n2555_), .A2(new_n4403_), .A3(pi1137), .ZN(new_n4404_));
  AOI21_X1   g01898(.A1(new_n2554_), .A2(new_n4403_), .B(new_n4402_), .ZN(new_n4405_));
  OAI21_X1   g01899(.A1(new_n4404_), .A2(new_n4405_), .B(pi0221), .ZN(new_n4406_));
  INV_X1     g01900(.I(new_n4406_), .ZN(new_n4407_));
  AOI21_X1   g01901(.A1(pi0216), .A2(pi0280), .B(pi0221), .ZN(new_n4408_));
  MUX2_X1    g01902(.I0(new_n3428_), .I1(new_n3377_), .S(pi0878), .Z(new_n4409_));
  INV_X1     g01903(.I(pi0878), .ZN(new_n4410_));
  AOI21_X1   g01904(.A1(new_n3426_), .A2(new_n4410_), .B(pi0168), .ZN(new_n4411_));
  AOI21_X1   g01905(.A1(new_n4409_), .A2(pi0168), .B(new_n4411_), .ZN(new_n4412_));
  INV_X1     g01906(.I(pi0168), .ZN(new_n4413_));
  NOR2_X1    g01907(.A1(new_n2438_), .A2(new_n4410_), .ZN(new_n4414_));
  NAND4_X1   g01908(.A1(new_n4414_), .A2(pi0105), .A3(new_n4413_), .A4(new_n2523_), .ZN(new_n4415_));
  INV_X1     g01909(.I(new_n4415_), .ZN(new_n4416_));
  NOR2_X1    g01910(.A1(new_n4416_), .A2(pi0216), .ZN(new_n4417_));
  INV_X1     g01911(.I(new_n4417_), .ZN(new_n4418_));
  NOR2_X1    g01912(.A1(new_n3559_), .A2(new_n4418_), .ZN(new_n4419_));
  OAI21_X1   g01913(.A1(new_n4412_), .A2(pi0228), .B(new_n4419_), .ZN(new_n4420_));
  AOI21_X1   g01914(.A1(new_n4420_), .A2(new_n4408_), .B(new_n4407_), .ZN(new_n4421_));
  MUX2_X1    g01915(.I0(new_n4421_), .I1(new_n4402_), .S(pi0215), .Z(new_n4422_));
  NAND3_X1   g01916(.A1(new_n2589_), .A2(pi0933), .A3(new_n4402_), .ZN(new_n4423_));
  OAI21_X1   g01917(.A1(new_n2593_), .A2(pi0933), .B(pi1137), .ZN(new_n4424_));
  AOI21_X1   g01918(.A1(new_n4424_), .A2(new_n4423_), .B(new_n2588_), .ZN(new_n4425_));
  INV_X1     g01919(.I(new_n4425_), .ZN(new_n4426_));
  AOI21_X1   g01920(.A1(pi0224), .A2(pi0280), .B(pi0222), .ZN(new_n4427_));
  OAI21_X1   g01921(.A1(new_n4414_), .A2(pi0224), .B(new_n4427_), .ZN(new_n4428_));
  NAND2_X1   g01922(.A1(new_n4426_), .A2(new_n4428_), .ZN(new_n4429_));
  NAND3_X1   g01923(.A1(new_n4429_), .A2(new_n2604_), .A3(pi1137), .ZN(new_n4430_));
  OAI21_X1   g01924(.A1(new_n4429_), .A2(pi0223), .B(new_n4402_), .ZN(new_n4431_));
  NAND3_X1   g01925(.A1(new_n4431_), .A2(new_n4430_), .A3(new_n2587_), .ZN(new_n4432_));
  NOR2_X1    g01926(.A1(new_n4432_), .A2(new_n3297_), .ZN(new_n4433_));
  INV_X1     g01927(.I(new_n4433_), .ZN(new_n4434_));
  NOR2_X1    g01928(.A1(new_n2566_), .A2(new_n4402_), .ZN(new_n4435_));
  NOR3_X1    g01929(.A1(new_n2490_), .A2(new_n4413_), .A3(new_n4410_), .ZN(new_n4436_));
  AOI21_X1   g01930(.A1(new_n2491_), .A2(new_n4413_), .B(pi0878), .ZN(new_n4437_));
  NOR4_X1    g01931(.A1(new_n4437_), .A2(pi0228), .A3(new_n3282_), .A4(new_n4436_), .ZN(new_n4438_));
  NOR2_X1    g01932(.A1(new_n4417_), .A2(new_n4408_), .ZN(new_n4439_));
  INV_X1     g01933(.I(new_n4439_), .ZN(new_n4440_));
  OAI21_X1   g01934(.A1(new_n4438_), .A2(new_n4440_), .B(new_n4406_), .ZN(new_n4441_));
  AOI21_X1   g01935(.A1(new_n4441_), .A2(new_n2566_), .B(new_n4435_), .ZN(new_n4442_));
  AOI21_X1   g01936(.A1(new_n4442_), .A2(pi0299), .B(new_n4434_), .ZN(new_n4443_));
  OAI21_X1   g01937(.A1(new_n4443_), .A2(new_n3154_), .B(new_n3172_), .ZN(new_n4444_));
  OAI21_X1   g01938(.A1(new_n3422_), .A2(new_n4410_), .B(new_n2595_), .ZN(new_n4445_));
  AOI21_X1   g01939(.A1(new_n4445_), .A2(new_n4427_), .B(new_n4425_), .ZN(new_n4446_));
  NAND2_X1   g01940(.A1(new_n3422_), .A2(new_n4427_), .ZN(new_n4447_));
  NOR2_X1    g01941(.A1(pi0223), .A2(pi0299), .ZN(new_n4448_));
  OAI21_X1   g01942(.A1(new_n4446_), .A2(new_n4447_), .B(new_n4448_), .ZN(new_n4449_));
  INV_X1     g01943(.I(new_n4435_), .ZN(new_n4450_));
  AOI21_X1   g01944(.A1(new_n4413_), .A2(new_n2523_), .B(new_n4408_), .ZN(new_n4451_));
  NAND2_X1   g01945(.A1(new_n4417_), .A2(new_n4451_), .ZN(new_n4452_));
  NAND2_X1   g01946(.A1(new_n4452_), .A2(new_n4406_), .ZN(new_n4453_));
  NAND2_X1   g01947(.A1(new_n4453_), .A2(new_n2566_), .ZN(new_n4454_));
  NAND2_X1   g01948(.A1(new_n4454_), .A2(new_n4450_), .ZN(new_n4455_));
  INV_X1     g01949(.I(new_n4455_), .ZN(new_n4456_));
  AOI21_X1   g01950(.A1(pi0216), .A2(pi0280), .B(new_n3886_), .ZN(new_n4457_));
  NOR2_X1    g01951(.A1(new_n4456_), .A2(new_n4457_), .ZN(new_n4458_));
  INV_X1     g01952(.I(new_n4458_), .ZN(new_n4459_));
  AOI21_X1   g01953(.A1(new_n4459_), .A2(pi0299), .B(new_n4434_), .ZN(new_n4460_));
  INV_X1     g01954(.I(new_n4460_), .ZN(new_n4461_));
  OAI21_X1   g01955(.A1(new_n4461_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n4462_));
  NAND4_X1   g01956(.A1(new_n4449_), .A2(new_n3154_), .A3(new_n4444_), .A4(new_n4462_), .ZN(new_n4463_));
  AOI21_X1   g01957(.A1(new_n4422_), .A2(pi0299), .B(new_n4463_), .ZN(new_n4464_));
  NOR3_X1    g01958(.A1(new_n3257_), .A2(new_n4413_), .A3(new_n4410_), .ZN(new_n4465_));
  AOI21_X1   g01959(.A1(new_n3256_), .A2(new_n4413_), .B(pi0878), .ZN(new_n4466_));
  NOR3_X1    g01960(.A1(new_n4465_), .A2(pi0228), .A3(new_n4466_), .ZN(new_n4467_));
  NAND2_X1   g01961(.A1(new_n4467_), .A2(new_n3283_), .ZN(new_n4468_));
  AOI21_X1   g01962(.A1(new_n4468_), .A2(new_n4439_), .B(new_n4407_), .ZN(new_n4469_));
  OAI21_X1   g01963(.A1(new_n4469_), .A2(pi0215), .B(new_n4450_), .ZN(new_n4470_));
  NAND2_X1   g01964(.A1(new_n4470_), .A2(new_n2587_), .ZN(new_n4471_));
  NOR2_X1    g01965(.A1(new_n4434_), .A2(new_n2545_), .ZN(new_n4472_));
  OAI21_X1   g01966(.A1(new_n4461_), .A2(new_n2544_), .B(pi0100), .ZN(new_n4473_));
  AOI21_X1   g01967(.A1(new_n4471_), .A2(new_n4472_), .B(new_n4473_), .ZN(new_n4474_));
  OAI21_X1   g01968(.A1(new_n4464_), .A2(new_n4474_), .B(new_n3177_), .ZN(new_n4475_));
  NAND2_X1   g01969(.A1(new_n4461_), .A2(new_n3198_), .ZN(new_n4476_));
  OAI21_X1   g01970(.A1(new_n3198_), .A2(new_n4443_), .B(new_n4476_), .ZN(new_n4477_));
  NAND2_X1   g01971(.A1(new_n4477_), .A2(pi0087), .ZN(new_n4478_));
  AOI21_X1   g01972(.A1(new_n4475_), .A2(new_n2628_), .B(new_n4478_), .ZN(new_n4479_));
  NAND4_X1   g01973(.A1(new_n4477_), .A2(new_n3203_), .A3(new_n2534_), .A4(new_n4461_), .ZN(new_n4480_));
  OAI21_X1   g01974(.A1(new_n4461_), .A2(new_n2538_), .B(new_n3227_), .ZN(new_n4481_));
  NAND2_X1   g01975(.A1(new_n4460_), .A2(pi0075), .ZN(new_n4482_));
  NAND4_X1   g01976(.A1(new_n4480_), .A2(new_n3329_), .A3(new_n4481_), .A4(new_n4482_), .ZN(new_n4483_));
  INV_X1     g01977(.I(new_n4442_), .ZN(new_n4484_));
  MUX2_X1    g01978(.I0(new_n4484_), .I1(new_n4458_), .S(new_n3336_), .Z(new_n4485_));
  NOR2_X1    g01979(.A1(new_n4484_), .A2(new_n3234_), .ZN(new_n4486_));
  OAI21_X1   g01980(.A1(new_n4458_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n4487_));
  OAI21_X1   g01981(.A1(new_n4486_), .A2(new_n4487_), .B(new_n2533_), .ZN(new_n4488_));
  AOI21_X1   g01982(.A1(pi0056), .A2(new_n4485_), .B(new_n4488_), .ZN(new_n4489_));
  OAI21_X1   g01983(.A1(new_n4479_), .A2(new_n4483_), .B(new_n4489_), .ZN(new_n4490_));
  NAND2_X1   g01984(.A1(new_n4442_), .A2(new_n3343_), .ZN(new_n4491_));
  AOI21_X1   g01985(.A1(new_n4459_), .A2(new_n3400_), .B(pi0062), .ZN(new_n4492_));
  NAND2_X1   g01986(.A1(new_n2571_), .A2(pi0240), .ZN(new_n4493_));
  AOI21_X1   g01987(.A1(new_n4492_), .A2(new_n4491_), .B(new_n4493_), .ZN(new_n4494_));
  NAND4_X1   g01988(.A1(new_n4456_), .A2(pi0240), .A3(new_n3405_), .A4(new_n4457_), .ZN(new_n4495_));
  NAND2_X1   g01989(.A1(pi0223), .A2(pi1137), .ZN(new_n4496_));
  NAND2_X1   g01990(.A1(new_n4449_), .A2(new_n3154_), .ZN(new_n4497_));
  NAND4_X1   g01991(.A1(new_n4497_), .A2(new_n2587_), .A3(new_n4446_), .A4(new_n4496_), .ZN(new_n4506_));
  NOR2_X1    g01992(.A1(new_n4418_), .A2(new_n4408_), .ZN(new_n4507_));
  AOI21_X1   g01993(.A1(new_n4467_), .A2(new_n4507_), .B(new_n4407_), .ZN(new_n4508_));
  MUX2_X1    g01994(.I0(new_n4508_), .I1(new_n4402_), .S(new_n2566_), .Z(new_n4509_));
  NOR2_X1    g01995(.A1(new_n4432_), .A2(new_n2545_), .ZN(new_n4510_));
  OAI21_X1   g01996(.A1(new_n4509_), .A2(pi0299), .B(new_n4510_), .ZN(new_n4511_));
  AOI21_X1   g01997(.A1(new_n4456_), .A2(pi0299), .B(new_n4432_), .ZN(new_n4512_));
  AOI21_X1   g01998(.A1(new_n4512_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4513_));
  NOR3_X1    g01999(.A1(new_n4437_), .A2(pi0228), .A3(new_n4436_), .ZN(new_n4514_));
  NAND2_X1   g02000(.A1(new_n4514_), .A2(new_n4507_), .ZN(new_n4515_));
  AOI21_X1   g02001(.A1(new_n4515_), .A2(new_n4406_), .B(pi0215), .ZN(new_n4516_));
  AOI21_X1   g02002(.A1(pi0215), .A2(new_n4402_), .B(new_n4516_), .ZN(new_n4517_));
  NAND3_X1   g02003(.A1(new_n4431_), .A2(new_n4430_), .A3(new_n2587_), .ZN(new_n4518_));
  NOR2_X1    g02004(.A1(pi0038), .A2(pi0100), .ZN(new_n4519_));
  OAI21_X1   g02005(.A1(new_n4518_), .A2(pi0039), .B(new_n4519_), .ZN(new_n4520_));
  AOI21_X1   g02006(.A1(new_n4511_), .A2(new_n4513_), .B(new_n4520_), .ZN(new_n4521_));
  AOI21_X1   g02007(.A1(new_n4521_), .A2(new_n4506_), .B(pi0087), .ZN(new_n4522_));
  NOR2_X1    g02008(.A1(new_n4512_), .A2(new_n3197_), .ZN(new_n4523_));
  AOI21_X1   g02009(.A1(new_n3197_), .A2(new_n4518_), .B(new_n4523_), .ZN(new_n4524_));
  NOR2_X1    g02010(.A1(new_n4524_), .A2(new_n3177_), .ZN(new_n4525_));
  OAI21_X1   g02011(.A1(new_n4522_), .A2(pi0075), .B(new_n4525_), .ZN(new_n4526_));
  NOR4_X1    g02012(.A1(new_n4524_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4512_), .ZN(new_n4527_));
  AOI21_X1   g02013(.A1(new_n4512_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4528_));
  AND2_X2    g02014(.A1(new_n4512_), .A2(pi0075), .Z(new_n4529_));
  NOR4_X1    g02015(.A1(new_n4527_), .A2(new_n3330_), .A3(new_n4528_), .A4(new_n4529_), .ZN(new_n4530_));
  MUX2_X1    g02016(.I0(new_n4517_), .I1(new_n4456_), .S(new_n3336_), .Z(new_n4531_));
  NAND2_X1   g02017(.A1(new_n4517_), .A2(new_n3233_), .ZN(new_n4532_));
  AOI21_X1   g02018(.A1(new_n4456_), .A2(new_n3234_), .B(pi0055), .ZN(new_n4533_));
  AOI21_X1   g02019(.A1(new_n4532_), .A2(new_n4533_), .B(new_n3503_), .ZN(new_n4534_));
  OAI21_X1   g02020(.A1(new_n3335_), .A2(new_n4531_), .B(new_n4534_), .ZN(new_n4535_));
  AOI21_X1   g02021(.A1(new_n4526_), .A2(new_n4530_), .B(new_n4535_), .ZN(new_n4536_));
  AND2_X2    g02022(.A1(new_n4517_), .A2(new_n3343_), .Z(new_n4537_));
  OAI21_X1   g02023(.A1(new_n3343_), .A2(new_n4455_), .B(new_n3240_), .ZN(new_n4538_));
  NOR2_X1    g02024(.A1(new_n3405_), .A2(pi0240), .ZN(new_n4539_));
  OAI21_X1   g02025(.A1(new_n4537_), .A2(new_n4538_), .B(new_n4539_), .ZN(new_n4540_));
  OAI21_X1   g02026(.A1(new_n4536_), .A2(new_n4540_), .B(new_n4495_), .ZN(new_n4541_));
  AOI21_X1   g02027(.A1(new_n4490_), .A2(new_n4494_), .B(new_n4541_), .ZN(po0162));
  INV_X1     g02028(.I(pi1136), .ZN(new_n4543_));
  NAND3_X1   g02029(.A1(new_n2554_), .A2(pi0928), .A3(new_n4543_), .ZN(new_n4544_));
  OAI21_X1   g02030(.A1(new_n2555_), .A2(pi0928), .B(pi1136), .ZN(new_n4545_));
  AOI21_X1   g02031(.A1(new_n4545_), .A2(new_n4544_), .B(new_n2550_), .ZN(new_n4546_));
  INV_X1     g02032(.I(new_n4546_), .ZN(new_n4547_));
  OAI21_X1   g02033(.A1(new_n3377_), .A2(pi0166), .B(pi0875), .ZN(new_n4548_));
  INV_X1     g02034(.I(pi0166), .ZN(new_n4549_));
  INV_X1     g02035(.I(pi0875), .ZN(new_n4550_));
  NOR2_X1    g02036(.A1(new_n2438_), .A2(new_n4550_), .ZN(new_n4551_));
  INV_X1     g02037(.I(new_n4551_), .ZN(new_n4552_));
  MUX2_X1    g02038(.I0(new_n4552_), .I1(new_n4549_), .S(new_n2522_), .Z(new_n4553_));
  NAND2_X1   g02039(.A1(new_n3430_), .A2(new_n4553_), .ZN(new_n4554_));
  AOI21_X1   g02040(.A1(new_n4554_), .A2(new_n2523_), .B(pi0216), .ZN(new_n4555_));
  NAND2_X1   g02041(.A1(pi0166), .A2(pi0875), .ZN(new_n4556_));
  OAI21_X1   g02042(.A1(new_n3651_), .A2(new_n4556_), .B(new_n4555_), .ZN(new_n4557_));
  AOI21_X1   g02043(.A1(new_n4548_), .A2(new_n2523_), .B(new_n4557_), .ZN(new_n4558_));
  INV_X1     g02044(.I(pi0266), .ZN(new_n4559_));
  OAI21_X1   g02045(.A1(new_n2562_), .A2(new_n4559_), .B(new_n2550_), .ZN(new_n4560_));
  OAI21_X1   g02046(.A1(new_n4558_), .A2(new_n4560_), .B(new_n4547_), .ZN(new_n4561_));
  MUX2_X1    g02047(.I0(new_n4561_), .I1(pi1136), .S(pi0215), .Z(new_n4562_));
  NOR2_X1    g02048(.A1(new_n2438_), .A2(pi0224), .ZN(new_n4563_));
  INV_X1     g02049(.I(new_n4563_), .ZN(new_n4564_));
  AOI21_X1   g02050(.A1(new_n4559_), .A2(pi0224), .B(pi0222), .ZN(new_n4565_));
  OAI21_X1   g02051(.A1(new_n4564_), .A2(pi0875), .B(new_n4565_), .ZN(new_n4566_));
  INV_X1     g02052(.I(new_n4566_), .ZN(new_n4567_));
  INV_X1     g02053(.I(pi0928), .ZN(new_n4568_));
  NOR3_X1    g02054(.A1(new_n2593_), .A2(new_n4568_), .A3(pi1136), .ZN(new_n4569_));
  AOI21_X1   g02055(.A1(new_n2589_), .A2(new_n4568_), .B(new_n4543_), .ZN(new_n4570_));
  OAI21_X1   g02056(.A1(new_n4569_), .A2(new_n4570_), .B(pi0222), .ZN(new_n4571_));
  INV_X1     g02057(.I(new_n4571_), .ZN(new_n4572_));
  NOR2_X1    g02058(.A1(new_n4572_), .A2(new_n4567_), .ZN(new_n4573_));
  NAND3_X1   g02059(.A1(new_n4573_), .A2(new_n2604_), .A3(pi1136), .ZN(new_n4574_));
  OAI21_X1   g02060(.A1(new_n4573_), .A2(pi0223), .B(new_n4543_), .ZN(new_n4575_));
  NOR2_X1    g02061(.A1(new_n2566_), .A2(new_n4543_), .ZN(new_n4576_));
  NOR2_X1    g02062(.A1(new_n2490_), .A2(pi0166), .ZN(new_n4577_));
  OAI21_X1   g02063(.A1(new_n2491_), .A2(pi0875), .B(new_n2523_), .ZN(new_n4578_));
  OAI22_X1   g02064(.A1(new_n4578_), .A2(new_n4577_), .B1(new_n2523_), .B2(new_n4553_), .ZN(new_n4579_));
  NOR2_X1    g02065(.A1(new_n4579_), .A2(new_n3282_), .ZN(new_n4580_));
  NAND3_X1   g02066(.A1(new_n4580_), .A2(new_n2562_), .A3(pi0266), .ZN(new_n4581_));
  OAI21_X1   g02067(.A1(new_n4580_), .A2(pi0216), .B(new_n4559_), .ZN(new_n4582_));
  NOR2_X1    g02068(.A1(new_n4546_), .A2(pi0221), .ZN(new_n4583_));
  NAND3_X1   g02069(.A1(new_n4582_), .A2(new_n4581_), .A3(new_n4583_), .ZN(new_n4584_));
  AOI21_X1   g02070(.A1(new_n4584_), .A2(new_n2566_), .B(new_n4576_), .ZN(new_n4585_));
  NAND3_X1   g02071(.A1(new_n4575_), .A2(new_n4574_), .A3(new_n2587_), .ZN(new_n4586_));
  AOI21_X1   g02072(.A1(new_n4586_), .A2(pi0039), .B(pi0038), .ZN(new_n4587_));
  NAND3_X1   g02073(.A1(new_n4575_), .A2(new_n4574_), .A3(new_n2587_), .ZN(new_n4588_));
  NOR2_X1    g02074(.A1(pi0166), .A2(pi0228), .ZN(new_n4589_));
  AOI21_X1   g02075(.A1(new_n4553_), .A2(pi0228), .B(new_n4589_), .ZN(new_n4590_));
  NOR3_X1    g02076(.A1(new_n4590_), .A2(pi0216), .A3(new_n4559_), .ZN(new_n4591_));
  AOI21_X1   g02077(.A1(new_n4590_), .A2(new_n2562_), .B(pi0266), .ZN(new_n4592_));
  INV_X1     g02078(.I(new_n4592_), .ZN(new_n4593_));
  NAND2_X1   g02079(.A1(new_n4593_), .A2(new_n4583_), .ZN(new_n4594_));
  OAI21_X1   g02080(.A1(new_n4594_), .A2(new_n4591_), .B(new_n2566_), .ZN(new_n4595_));
  OAI21_X1   g02081(.A1(new_n2566_), .A2(new_n4543_), .B(new_n4595_), .ZN(new_n4596_));
  INV_X1     g02082(.I(new_n4596_), .ZN(new_n4597_));
  NOR2_X1    g02083(.A1(new_n4597_), .A2(new_n3288_), .ZN(new_n4598_));
  INV_X1     g02084(.I(new_n4598_), .ZN(new_n4599_));
  AOI21_X1   g02085(.A1(new_n4599_), .A2(pi0299), .B(new_n4588_), .ZN(new_n4600_));
  AOI21_X1   g02086(.A1(new_n4600_), .A2(pi0038), .B(pi0100), .ZN(new_n4601_));
  AOI21_X1   g02087(.A1(pi0223), .A2(pi1136), .B(pi0299), .ZN(new_n4602_));
  NOR2_X1    g02088(.A1(new_n3421_), .A2(new_n3155_), .ZN(new_n4603_));
  INV_X1     g02089(.I(new_n4603_), .ZN(new_n4604_));
  NAND2_X1   g02090(.A1(new_n4604_), .A2(new_n4573_), .ZN(new_n4605_));
  NAND2_X1   g02091(.A1(new_n4605_), .A2(new_n2604_), .ZN(new_n4606_));
  AOI21_X1   g02092(.A1(new_n4606_), .A2(new_n4602_), .B(pi0039), .ZN(new_n4607_));
  NOR3_X1    g02093(.A1(new_n4601_), .A2(new_n4587_), .A3(new_n4607_), .ZN(new_n4608_));
  OAI21_X1   g02094(.A1(new_n4562_), .A2(new_n2587_), .B(new_n4608_), .ZN(new_n4609_));
  NOR2_X1    g02095(.A1(new_n4553_), .A2(new_n2523_), .ZN(new_n4610_));
  INV_X1     g02096(.I(new_n3253_), .ZN(new_n4611_));
  MUX2_X1    g02097(.I0(new_n4611_), .I1(new_n3608_), .S(new_n2574_), .Z(new_n4612_));
  NOR2_X1    g02098(.A1(new_n4611_), .A2(pi0875), .ZN(new_n4613_));
  OAI22_X1   g02099(.A1(new_n4612_), .A2(new_n4550_), .B1(new_n4549_), .B2(new_n4613_), .ZN(new_n4614_));
  AOI21_X1   g02100(.A1(new_n4614_), .A2(new_n2523_), .B(new_n4610_), .ZN(new_n4615_));
  AND2_X2    g02101(.A1(new_n4615_), .A2(new_n3283_), .Z(new_n4616_));
  NAND3_X1   g02102(.A1(new_n4616_), .A2(new_n2562_), .A3(pi0266), .ZN(new_n4617_));
  OAI21_X1   g02103(.A1(new_n4616_), .A2(pi0216), .B(new_n4559_), .ZN(new_n4618_));
  NAND3_X1   g02104(.A1(new_n4618_), .A2(new_n4617_), .A3(new_n4583_), .ZN(new_n4619_));
  AOI21_X1   g02105(.A1(new_n4619_), .A2(new_n2566_), .B(new_n4576_), .ZN(new_n4620_));
  NAND4_X1   g02106(.A1(new_n4575_), .A2(new_n4574_), .A3(new_n2587_), .A4(new_n2545_), .ZN(new_n4621_));
  AOI21_X1   g02107(.A1(new_n4600_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4622_));
  OAI21_X1   g02108(.A1(new_n4620_), .A2(new_n4621_), .B(new_n4622_), .ZN(new_n4623_));
  AOI21_X1   g02109(.A1(new_n4609_), .A2(new_n4623_), .B(pi0087), .ZN(new_n4624_));
  NOR2_X1    g02110(.A1(new_n4600_), .A2(new_n3197_), .ZN(new_n4625_));
  AOI21_X1   g02111(.A1(new_n3197_), .A2(new_n4586_), .B(new_n4625_), .ZN(new_n4626_));
  NOR2_X1    g02112(.A1(new_n4626_), .A2(new_n3177_), .ZN(new_n4627_));
  OAI21_X1   g02113(.A1(new_n4624_), .A2(pi0075), .B(new_n4627_), .ZN(new_n4628_));
  NOR4_X1    g02114(.A1(new_n4626_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4600_), .ZN(new_n4629_));
  AOI21_X1   g02115(.A1(new_n4600_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4630_));
  AND2_X2    g02116(.A1(new_n4600_), .A2(pi0075), .Z(new_n4631_));
  NOR4_X1    g02117(.A1(new_n4629_), .A2(new_n3330_), .A3(new_n4630_), .A4(new_n4631_), .ZN(new_n4632_));
  MUX2_X1    g02118(.I0(new_n4585_), .I1(new_n4599_), .S(new_n3336_), .Z(new_n4633_));
  NAND2_X1   g02119(.A1(new_n4585_), .A2(new_n3233_), .ZN(new_n4634_));
  AOI21_X1   g02120(.A1(new_n4599_), .A2(new_n3234_), .B(pi0055), .ZN(new_n4635_));
  AOI21_X1   g02121(.A1(new_n4635_), .A2(new_n4634_), .B(new_n3503_), .ZN(new_n4636_));
  OAI21_X1   g02122(.A1(new_n3335_), .A2(new_n4633_), .B(new_n4636_), .ZN(new_n4637_));
  AOI21_X1   g02123(.A1(new_n4628_), .A2(new_n4632_), .B(new_n4637_), .ZN(new_n4638_));
  AND2_X2    g02124(.A1(new_n4585_), .A2(new_n3343_), .Z(new_n4639_));
  OAI21_X1   g02125(.A1(new_n4598_), .A2(new_n3343_), .B(new_n3240_), .ZN(new_n4640_));
  OAI21_X1   g02126(.A1(new_n4639_), .A2(new_n4640_), .B(new_n2571_), .ZN(new_n4641_));
  NOR2_X1    g02127(.A1(new_n4638_), .A2(new_n4641_), .ZN(new_n4642_));
  OAI21_X1   g02128(.A1(new_n4599_), .A2(new_n2571_), .B(pi0245), .ZN(new_n4643_));
  AOI21_X1   g02129(.A1(new_n3651_), .A2(new_n4549_), .B(new_n3428_), .ZN(new_n4644_));
  INV_X1     g02130(.I(new_n3428_), .ZN(new_n4645_));
  NOR3_X1    g02131(.A1(new_n3651_), .A2(pi0166), .A3(new_n4645_), .ZN(new_n4646_));
  OAI21_X1   g02132(.A1(new_n4646_), .A2(new_n4644_), .B(pi0875), .ZN(new_n4647_));
  NAND2_X1   g02133(.A1(new_n3376_), .A2(new_n4550_), .ZN(new_n4648_));
  NAND3_X1   g02134(.A1(new_n3430_), .A2(new_n2562_), .A3(pi0228), .ZN(new_n4649_));
  AOI21_X1   g02135(.A1(new_n4648_), .A2(new_n4549_), .B(new_n4649_), .ZN(new_n4650_));
  AOI22_X1   g02136(.A1(new_n4647_), .A2(new_n4650_), .B1(pi0216), .B2(pi0266), .ZN(new_n4651_));
  OAI21_X1   g02137(.A1(new_n4651_), .A2(pi0221), .B(new_n4547_), .ZN(new_n4652_));
  MUX2_X1    g02138(.I0(new_n4652_), .I1(new_n4543_), .S(pi0215), .Z(new_n4653_));
  NOR4_X1    g02139(.A1(new_n4604_), .A2(new_n4567_), .A3(new_n4572_), .A4(new_n4602_), .ZN(new_n4654_));
  AOI21_X1   g02140(.A1(new_n4653_), .A2(pi0299), .B(new_n4654_), .ZN(new_n4655_));
  NAND2_X1   g02141(.A1(new_n4606_), .A2(new_n4602_), .ZN(new_n4656_));
  NOR3_X1    g02142(.A1(new_n4588_), .A2(new_n3156_), .A3(new_n4552_), .ZN(new_n4657_));
  AOI21_X1   g02143(.A1(new_n4579_), .A2(new_n2562_), .B(new_n4560_), .ZN(new_n4658_));
  NAND2_X1   g02144(.A1(new_n4547_), .A2(new_n2566_), .ZN(new_n4659_));
  OAI22_X1   g02145(.A1(new_n4658_), .A2(new_n4659_), .B1(new_n2566_), .B2(pi1136), .ZN(new_n4660_));
  NOR2_X1    g02146(.A1(new_n4660_), .A2(new_n2587_), .ZN(new_n4661_));
  NOR2_X1    g02147(.A1(new_n4661_), .A2(new_n4657_), .ZN(new_n4662_));
  NAND3_X1   g02148(.A1(new_n4656_), .A2(pi0038), .A3(new_n3154_), .ZN(new_n4663_));
  NOR2_X1    g02149(.A1(new_n4615_), .A2(pi0216), .ZN(new_n4664_));
  OAI21_X1   g02150(.A1(new_n4664_), .A2(new_n4560_), .B(new_n4547_), .ZN(new_n4665_));
  MUX2_X1    g02151(.I0(new_n4665_), .I1(new_n4543_), .S(new_n2566_), .Z(new_n4666_));
  NOR2_X1    g02152(.A1(new_n4657_), .A2(new_n2545_), .ZN(new_n4667_));
  OAI21_X1   g02153(.A1(new_n4666_), .A2(pi0299), .B(new_n4667_), .ZN(new_n4668_));
  AOI21_X1   g02154(.A1(new_n4597_), .A2(pi0299), .B(new_n4657_), .ZN(new_n4669_));
  AOI21_X1   g02155(.A1(new_n4669_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4670_));
  INV_X1     g02156(.I(new_n4669_), .ZN(new_n4671_));
  OAI21_X1   g02157(.A1(new_n4671_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n4672_));
  AOI21_X1   g02158(.A1(new_n4668_), .A2(new_n4670_), .B(new_n4672_), .ZN(new_n4673_));
  OAI21_X1   g02159(.A1(new_n4655_), .A2(new_n4663_), .B(new_n4673_), .ZN(new_n4674_));
  AOI21_X1   g02160(.A1(new_n4674_), .A2(new_n3177_), .B(pi0075), .ZN(new_n4675_));
  NOR2_X1    g02161(.A1(new_n4662_), .A2(new_n3198_), .ZN(new_n4676_));
  AOI21_X1   g02162(.A1(new_n3198_), .A2(new_n4671_), .B(new_n4676_), .ZN(new_n4677_));
  OR2_X2     g02163(.A1(new_n4677_), .A2(new_n3177_), .Z(new_n4678_));
  NOR4_X1    g02164(.A1(new_n4677_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4669_), .ZN(new_n4679_));
  AOI21_X1   g02165(.A1(new_n4669_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4680_));
  NOR2_X1    g02166(.A1(new_n4671_), .A2(new_n2628_), .ZN(new_n4681_));
  NOR4_X1    g02167(.A1(new_n4679_), .A2(new_n3330_), .A3(new_n4680_), .A4(new_n4681_), .ZN(new_n4682_));
  OAI21_X1   g02168(.A1(new_n4675_), .A2(new_n4678_), .B(new_n4682_), .ZN(new_n4683_));
  MUX2_X1    g02169(.I0(new_n4660_), .I1(new_n4596_), .S(new_n3336_), .Z(new_n4684_));
  NOR2_X1    g02170(.A1(new_n4660_), .A2(new_n3234_), .ZN(new_n4685_));
  OAI21_X1   g02171(.A1(new_n4596_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n4686_));
  OAI21_X1   g02172(.A1(new_n4685_), .A2(new_n4686_), .B(new_n2533_), .ZN(new_n4687_));
  AOI21_X1   g02173(.A1(pi0056), .A2(new_n4684_), .B(new_n4687_), .ZN(new_n4688_));
  NOR2_X1    g02174(.A1(new_n4660_), .A2(new_n3400_), .ZN(new_n4689_));
  OAI21_X1   g02175(.A1(new_n4596_), .A2(new_n3343_), .B(new_n3240_), .ZN(new_n4690_));
  OAI21_X1   g02176(.A1(new_n4689_), .A2(new_n4690_), .B(new_n2571_), .ZN(new_n4691_));
  AOI21_X1   g02177(.A1(new_n4683_), .A2(new_n4688_), .B(new_n4691_), .ZN(new_n4692_));
  INV_X1     g02178(.I(pi0245), .ZN(new_n4693_));
  OAI21_X1   g02179(.A1(new_n4597_), .A2(new_n2571_), .B(new_n4693_), .ZN(new_n4694_));
  OAI22_X1   g02180(.A1(new_n4692_), .A2(new_n4694_), .B1(new_n4642_), .B2(new_n4643_), .ZN(po0163));
  INV_X1     g02181(.I(pi1135), .ZN(new_n4696_));
  NAND3_X1   g02182(.A1(new_n2554_), .A2(pi0938), .A3(new_n4696_), .ZN(new_n4697_));
  OAI21_X1   g02183(.A1(new_n2555_), .A2(pi0938), .B(pi1135), .ZN(new_n4698_));
  AOI21_X1   g02184(.A1(new_n4698_), .A2(new_n4697_), .B(new_n2550_), .ZN(new_n4699_));
  OAI21_X1   g02185(.A1(new_n3377_), .A2(pi0161), .B(pi0879), .ZN(new_n4700_));
  INV_X1     g02186(.I(pi0161), .ZN(new_n4701_));
  INV_X1     g02187(.I(pi0879), .ZN(new_n4702_));
  NOR2_X1    g02188(.A1(new_n2438_), .A2(new_n4702_), .ZN(new_n4703_));
  INV_X1     g02189(.I(new_n4703_), .ZN(new_n4704_));
  MUX2_X1    g02190(.I0(new_n4704_), .I1(new_n4701_), .S(new_n2522_), .Z(new_n4705_));
  NAND2_X1   g02191(.A1(new_n3430_), .A2(new_n4705_), .ZN(new_n4706_));
  AOI21_X1   g02192(.A1(new_n4706_), .A2(new_n2523_), .B(pi0216), .ZN(new_n4707_));
  NAND2_X1   g02193(.A1(pi0161), .A2(pi0879), .ZN(new_n4708_));
  OAI21_X1   g02194(.A1(new_n3651_), .A2(new_n4708_), .B(new_n4707_), .ZN(new_n4709_));
  AOI21_X1   g02195(.A1(new_n4700_), .A2(new_n2523_), .B(new_n4709_), .ZN(new_n4710_));
  INV_X1     g02196(.I(pi0279), .ZN(new_n4711_));
  OAI21_X1   g02197(.A1(new_n2562_), .A2(new_n4711_), .B(new_n2550_), .ZN(new_n4712_));
  NOR2_X1    g02198(.A1(new_n4710_), .A2(new_n4712_), .ZN(new_n4713_));
  NOR2_X1    g02199(.A1(new_n4713_), .A2(new_n4699_), .ZN(new_n4714_));
  MUX2_X1    g02200(.I0(new_n4714_), .I1(new_n4696_), .S(pi0215), .Z(new_n4715_));
  NAND2_X1   g02201(.A1(new_n4715_), .A2(pi0299), .ZN(new_n4716_));
  NOR2_X1    g02202(.A1(new_n2566_), .A2(new_n4696_), .ZN(new_n4717_));
  INV_X1     g02203(.I(new_n4717_), .ZN(new_n4718_));
  OR2_X2     g02204(.A1(new_n4705_), .A2(new_n2523_), .Z(new_n4719_));
  NAND3_X1   g02205(.A1(new_n3248_), .A2(new_n3250_), .A3(new_n4549_), .ZN(new_n4720_));
  XOR2_X1    g02206(.A1(new_n4720_), .A2(new_n3253_), .Z(new_n4721_));
  NOR2_X1    g02207(.A1(new_n4721_), .A2(new_n4702_), .ZN(new_n4722_));
  AOI21_X1   g02208(.A1(new_n3253_), .A2(new_n4702_), .B(new_n4701_), .ZN(new_n4723_));
  OAI21_X1   g02209(.A1(new_n4722_), .A2(new_n4723_), .B(new_n2523_), .ZN(new_n4724_));
  NAND3_X1   g02210(.A1(new_n4724_), .A2(new_n3283_), .A3(new_n4719_), .ZN(new_n4725_));
  NOR3_X1    g02211(.A1(new_n4725_), .A2(pi0216), .A3(new_n4711_), .ZN(new_n4726_));
  NOR2_X1    g02212(.A1(new_n4699_), .A2(pi0221), .ZN(new_n4727_));
  INV_X1     g02213(.I(new_n4727_), .ZN(new_n4728_));
  AOI21_X1   g02214(.A1(new_n4725_), .A2(new_n2562_), .B(pi0279), .ZN(new_n4729_));
  NOR3_X1    g02215(.A1(new_n4726_), .A2(new_n4729_), .A3(new_n4728_), .ZN(new_n4730_));
  OAI21_X1   g02216(.A1(new_n4730_), .A2(pi0215), .B(new_n4718_), .ZN(new_n4731_));
  INV_X1     g02217(.I(pi0938), .ZN(new_n4732_));
  NOR3_X1    g02218(.A1(new_n2593_), .A2(new_n4732_), .A3(pi1135), .ZN(new_n4733_));
  AOI21_X1   g02219(.A1(new_n2589_), .A2(new_n4732_), .B(new_n4696_), .ZN(new_n4734_));
  OAI21_X1   g02220(.A1(new_n4733_), .A2(new_n4734_), .B(pi0222), .ZN(new_n4735_));
  INV_X1     g02221(.I(new_n4735_), .ZN(new_n4736_));
  AOI21_X1   g02222(.A1(new_n4711_), .A2(pi0224), .B(pi0222), .ZN(new_n4737_));
  OAI21_X1   g02223(.A1(new_n4564_), .A2(pi0879), .B(new_n4737_), .ZN(new_n4738_));
  INV_X1     g02224(.I(new_n4738_), .ZN(new_n4739_));
  NOR2_X1    g02225(.A1(new_n4736_), .A2(new_n4739_), .ZN(new_n4740_));
  NAND3_X1   g02226(.A1(new_n4740_), .A2(new_n2604_), .A3(pi1135), .ZN(new_n4741_));
  OAI21_X1   g02227(.A1(new_n4740_), .A2(pi0223), .B(new_n4696_), .ZN(new_n4742_));
  NAND3_X1   g02228(.A1(new_n4742_), .A2(new_n4741_), .A3(new_n2587_), .ZN(new_n4743_));
  NOR2_X1    g02229(.A1(new_n4743_), .A2(new_n3671_), .ZN(new_n4744_));
  NAND2_X1   g02230(.A1(new_n4731_), .A2(new_n4744_), .ZN(new_n4745_));
  NOR2_X1    g02231(.A1(pi0161), .A2(pi0228), .ZN(new_n4746_));
  AOI21_X1   g02232(.A1(new_n4705_), .A2(pi0228), .B(new_n4746_), .ZN(new_n4747_));
  NOR3_X1    g02233(.A1(new_n4747_), .A2(pi0216), .A3(new_n4711_), .ZN(new_n4748_));
  AOI21_X1   g02234(.A1(new_n4747_), .A2(new_n2562_), .B(pi0279), .ZN(new_n4749_));
  OR2_X2     g02235(.A1(new_n4749_), .A2(new_n4728_), .Z(new_n4750_));
  OAI21_X1   g02236(.A1(new_n4750_), .A2(new_n4748_), .B(new_n2566_), .ZN(new_n4751_));
  NAND2_X1   g02237(.A1(new_n4751_), .A2(new_n4718_), .ZN(new_n4752_));
  INV_X1     g02238(.I(new_n4752_), .ZN(new_n4753_));
  NOR2_X1    g02239(.A1(new_n4753_), .A2(new_n3288_), .ZN(new_n4754_));
  INV_X1     g02240(.I(new_n4754_), .ZN(new_n4755_));
  AOI21_X1   g02241(.A1(new_n4755_), .A2(pi0299), .B(new_n4743_), .ZN(new_n4756_));
  AOI21_X1   g02242(.A1(new_n4756_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4757_));
  NOR2_X1    g02243(.A1(new_n2490_), .A2(pi0161), .ZN(new_n4758_));
  OAI21_X1   g02244(.A1(new_n2491_), .A2(pi0879), .B(new_n2523_), .ZN(new_n4759_));
  OAI21_X1   g02245(.A1(new_n4759_), .A2(new_n4758_), .B(new_n4719_), .ZN(new_n4760_));
  NOR2_X1    g02246(.A1(new_n4760_), .A2(new_n3282_), .ZN(new_n4761_));
  NAND3_X1   g02247(.A1(new_n4761_), .A2(new_n2562_), .A3(pi0279), .ZN(new_n4762_));
  OAI21_X1   g02248(.A1(new_n4761_), .A2(pi0216), .B(new_n4711_), .ZN(new_n4763_));
  NAND3_X1   g02249(.A1(new_n4763_), .A2(new_n4762_), .A3(new_n4727_), .ZN(new_n4764_));
  AOI21_X1   g02250(.A1(new_n4764_), .A2(new_n2566_), .B(new_n4717_), .ZN(new_n4765_));
  AOI21_X1   g02251(.A1(new_n4765_), .A2(pi0299), .B(new_n4743_), .ZN(new_n4766_));
  NAND2_X1   g02252(.A1(new_n4766_), .A2(new_n3154_), .ZN(new_n4767_));
  NAND2_X1   g02253(.A1(new_n4756_), .A2(pi0038), .ZN(new_n4768_));
  NAND2_X1   g02254(.A1(new_n4604_), .A2(new_n4740_), .ZN(new_n4769_));
  NOR2_X1    g02255(.A1(new_n2587_), .A2(pi0223), .ZN(new_n4770_));
  NAND2_X1   g02256(.A1(new_n4769_), .A2(new_n4770_), .ZN(new_n4771_));
  NAND4_X1   g02257(.A1(new_n4768_), .A2(new_n4767_), .A3(new_n2546_), .A4(new_n4771_), .ZN(new_n4772_));
  AOI21_X1   g02258(.A1(new_n4745_), .A2(new_n4757_), .B(new_n4772_), .ZN(new_n4773_));
  AOI21_X1   g02259(.A1(new_n4716_), .A2(new_n4773_), .B(pi0087), .ZN(new_n4774_));
  INV_X1     g02260(.I(new_n4756_), .ZN(new_n4775_));
  NOR2_X1    g02261(.A1(new_n4766_), .A2(new_n3198_), .ZN(new_n4776_));
  AOI21_X1   g02262(.A1(new_n3198_), .A2(new_n4775_), .B(new_n4776_), .ZN(new_n4777_));
  NOR2_X1    g02263(.A1(new_n4777_), .A2(new_n3177_), .ZN(new_n4778_));
  OAI21_X1   g02264(.A1(new_n4774_), .A2(pi0075), .B(new_n4778_), .ZN(new_n4779_));
  NOR4_X1    g02265(.A1(new_n4777_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4756_), .ZN(new_n4780_));
  AOI21_X1   g02266(.A1(new_n4756_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4781_));
  NOR2_X1    g02267(.A1(new_n4775_), .A2(new_n2628_), .ZN(new_n4782_));
  NOR4_X1    g02268(.A1(new_n4780_), .A2(new_n3330_), .A3(new_n4781_), .A4(new_n4782_), .ZN(new_n4783_));
  MUX2_X1    g02269(.I0(new_n4765_), .I1(new_n4755_), .S(new_n3336_), .Z(new_n4784_));
  NAND2_X1   g02270(.A1(new_n4765_), .A2(new_n3233_), .ZN(new_n4785_));
  AOI21_X1   g02271(.A1(new_n4755_), .A2(new_n3234_), .B(pi0055), .ZN(new_n4786_));
  AOI21_X1   g02272(.A1(new_n4786_), .A2(new_n4785_), .B(new_n3503_), .ZN(new_n4787_));
  OAI21_X1   g02273(.A1(new_n3335_), .A2(new_n4784_), .B(new_n4787_), .ZN(new_n4788_));
  AOI21_X1   g02274(.A1(new_n4779_), .A2(new_n4783_), .B(new_n4788_), .ZN(new_n4789_));
  AND2_X2    g02275(.A1(new_n4765_), .A2(new_n3343_), .Z(new_n4790_));
  OAI21_X1   g02276(.A1(new_n4754_), .A2(new_n3343_), .B(new_n3240_), .ZN(new_n4791_));
  OAI21_X1   g02277(.A1(new_n4790_), .A2(new_n4791_), .B(new_n2571_), .ZN(new_n4792_));
  NOR2_X1    g02278(.A1(new_n4789_), .A2(new_n4792_), .ZN(new_n4793_));
  OAI21_X1   g02279(.A1(new_n4755_), .A2(new_n2571_), .B(pi0244), .ZN(new_n4794_));
  OAI21_X1   g02280(.A1(new_n3426_), .A2(pi0161), .B(new_n4645_), .ZN(new_n4795_));
  NAND3_X1   g02281(.A1(new_n3426_), .A2(new_n4701_), .A3(new_n3428_), .ZN(new_n4796_));
  AOI21_X1   g02282(.A1(new_n4795_), .A2(new_n4796_), .B(new_n4702_), .ZN(new_n4797_));
  OAI21_X1   g02283(.A1(new_n3377_), .A2(pi0879), .B(new_n4701_), .ZN(new_n4798_));
  NAND4_X1   g02284(.A1(new_n4798_), .A2(pi0228), .A3(new_n3430_), .A4(new_n4707_), .ZN(new_n4799_));
  OAI22_X1   g02285(.A1(new_n4799_), .A2(new_n4797_), .B1(new_n2562_), .B2(new_n4711_), .ZN(new_n4800_));
  AOI21_X1   g02286(.A1(new_n4800_), .A2(new_n2550_), .B(new_n4699_), .ZN(new_n4801_));
  MUX2_X1    g02287(.I0(new_n4801_), .I1(pi1135), .S(pi0215), .Z(new_n4802_));
  INV_X1     g02288(.I(new_n4699_), .ZN(new_n4803_));
  AOI21_X1   g02289(.A1(new_n4724_), .A2(new_n4719_), .B(pi0216), .ZN(new_n4804_));
  OAI21_X1   g02290(.A1(new_n4804_), .A2(new_n4712_), .B(new_n4803_), .ZN(new_n4805_));
  MUX2_X1    g02291(.I0(new_n4805_), .I1(new_n4696_), .S(new_n2566_), .Z(new_n4806_));
  NOR3_X1    g02292(.A1(new_n4743_), .A2(new_n3156_), .A3(new_n4704_), .ZN(new_n4807_));
  NOR2_X1    g02293(.A1(new_n4807_), .A2(new_n2545_), .ZN(new_n4808_));
  OAI21_X1   g02294(.A1(new_n4806_), .A2(pi0299), .B(new_n4808_), .ZN(new_n4809_));
  AOI21_X1   g02295(.A1(new_n4753_), .A2(pi0299), .B(new_n4807_), .ZN(new_n4810_));
  AOI21_X1   g02296(.A1(new_n4810_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4811_));
  INV_X1     g02297(.I(new_n4807_), .ZN(new_n4812_));
  AOI21_X1   g02298(.A1(new_n4760_), .A2(new_n2562_), .B(new_n4712_), .ZN(new_n4813_));
  NAND2_X1   g02299(.A1(new_n4803_), .A2(new_n2566_), .ZN(new_n4814_));
  OAI22_X1   g02300(.A1(new_n4813_), .A2(new_n4814_), .B1(new_n2566_), .B2(pi1135), .ZN(new_n4815_));
  OAI21_X1   g02301(.A1(new_n4815_), .A2(new_n2587_), .B(new_n4812_), .ZN(new_n4816_));
  INV_X1     g02302(.I(new_n4770_), .ZN(new_n4817_));
  AOI21_X1   g02303(.A1(new_n4604_), .A2(new_n4739_), .B(new_n4736_), .ZN(new_n4818_));
  OAI21_X1   g02304(.A1(new_n4818_), .A2(new_n4817_), .B(new_n2546_), .ZN(new_n4819_));
  AOI21_X1   g02305(.A1(pi0038), .A2(new_n4810_), .B(new_n4819_), .ZN(new_n4820_));
  OAI21_X1   g02306(.A1(new_n4816_), .A2(pi0039), .B(new_n4820_), .ZN(new_n4821_));
  AOI21_X1   g02307(.A1(new_n4809_), .A2(new_n4811_), .B(new_n4821_), .ZN(new_n4822_));
  OAI21_X1   g02308(.A1(new_n4802_), .A2(new_n2587_), .B(new_n4822_), .ZN(new_n4823_));
  AOI21_X1   g02309(.A1(new_n4823_), .A2(new_n3177_), .B(pi0075), .ZN(new_n4824_));
  NOR2_X1    g02310(.A1(new_n4810_), .A2(new_n3197_), .ZN(new_n4825_));
  AOI21_X1   g02311(.A1(new_n4816_), .A2(new_n3197_), .B(new_n4825_), .ZN(new_n4826_));
  OR2_X2     g02312(.A1(new_n4826_), .A2(new_n3177_), .Z(new_n4827_));
  NOR4_X1    g02313(.A1(new_n4826_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4810_), .ZN(new_n4828_));
  AOI21_X1   g02314(.A1(new_n4810_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4829_));
  AND2_X2    g02315(.A1(new_n4810_), .A2(pi0075), .Z(new_n4830_));
  NOR4_X1    g02316(.A1(new_n4828_), .A2(new_n3330_), .A3(new_n4829_), .A4(new_n4830_), .ZN(new_n4831_));
  OAI21_X1   g02317(.A1(new_n4824_), .A2(new_n4827_), .B(new_n4831_), .ZN(new_n4832_));
  MUX2_X1    g02318(.I0(new_n4815_), .I1(new_n4752_), .S(new_n3336_), .Z(new_n4833_));
  NOR2_X1    g02319(.A1(new_n4815_), .A2(new_n3234_), .ZN(new_n4834_));
  OAI21_X1   g02320(.A1(new_n4752_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n4835_));
  OAI21_X1   g02321(.A1(new_n4834_), .A2(new_n4835_), .B(new_n2533_), .ZN(new_n4836_));
  AOI21_X1   g02322(.A1(pi0056), .A2(new_n4833_), .B(new_n4836_), .ZN(new_n4837_));
  NOR2_X1    g02323(.A1(new_n4815_), .A2(new_n3400_), .ZN(new_n4838_));
  OAI21_X1   g02324(.A1(new_n4752_), .A2(new_n3343_), .B(new_n3240_), .ZN(new_n4839_));
  OAI21_X1   g02325(.A1(new_n4838_), .A2(new_n4839_), .B(new_n2571_), .ZN(new_n4840_));
  AOI21_X1   g02326(.A1(new_n4832_), .A2(new_n4837_), .B(new_n4840_), .ZN(new_n4841_));
  INV_X1     g02327(.I(pi0244), .ZN(new_n4842_));
  OAI21_X1   g02328(.A1(new_n4753_), .A2(new_n2571_), .B(new_n4842_), .ZN(new_n4843_));
  OAI22_X1   g02329(.A1(new_n4793_), .A2(new_n4794_), .B1(new_n4841_), .B2(new_n4843_), .ZN(po0164));
  NOR3_X1    g02330(.A1(new_n2555_), .A2(new_n2550_), .A3(pi0930), .ZN(new_n4845_));
  INV_X1     g02331(.I(pi0846), .ZN(new_n4846_));
  NOR2_X1    g02332(.A1(new_n2438_), .A2(new_n4846_), .ZN(new_n4847_));
  INV_X1     g02333(.I(new_n4847_), .ZN(new_n4848_));
  MUX2_X1    g02334(.I0(new_n4848_), .I1(new_n3250_), .S(new_n2522_), .Z(new_n4849_));
  NOR2_X1    g02335(.A1(new_n4849_), .A2(new_n2523_), .ZN(new_n4850_));
  INV_X1     g02336(.I(new_n4850_), .ZN(new_n4851_));
  AOI21_X1   g02337(.A1(new_n2490_), .A2(new_n4846_), .B(pi0228), .ZN(new_n4852_));
  OAI21_X1   g02338(.A1(pi0152), .A2(new_n2490_), .B(new_n4852_), .ZN(new_n4853_));
  NAND2_X1   g02339(.A1(new_n2562_), .A2(pi0221), .ZN(new_n4854_));
  AOI21_X1   g02340(.A1(new_n4853_), .A2(new_n4851_), .B(new_n4854_), .ZN(new_n4855_));
  OAI21_X1   g02341(.A1(new_n4855_), .A2(new_n4845_), .B(new_n2566_), .ZN(new_n4856_));
  INV_X1     g02342(.I(new_n4845_), .ZN(new_n4857_));
  AOI21_X1   g02343(.A1(pi0216), .A2(pi0278), .B(pi0221), .ZN(new_n4858_));
  NOR2_X1    g02344(.A1(new_n3250_), .A2(pi0228), .ZN(new_n4859_));
  OAI21_X1   g02345(.A1(new_n4850_), .A2(new_n4859_), .B(new_n2562_), .ZN(new_n4860_));
  NAND2_X1   g02346(.A1(new_n4860_), .A2(new_n4858_), .ZN(new_n4861_));
  AOI21_X1   g02347(.A1(new_n4861_), .A2(new_n4857_), .B(pi0215), .ZN(new_n4862_));
  OAI21_X1   g02348(.A1(new_n3343_), .A2(new_n4862_), .B(new_n3240_), .ZN(new_n4863_));
  AOI21_X1   g02349(.A1(new_n4856_), .A2(new_n3343_), .B(new_n4863_), .ZN(new_n4864_));
  MUX2_X1    g02350(.I0(new_n4645_), .I1(new_n3426_), .S(new_n3250_), .Z(new_n4865_));
  OAI21_X1   g02351(.A1(new_n3377_), .A2(pi0846), .B(new_n3250_), .ZN(new_n4866_));
  NOR3_X1    g02352(.A1(new_n2522_), .A2(pi0152), .A3(pi0228), .ZN(new_n4867_));
  NOR2_X1    g02353(.A1(new_n3422_), .A2(pi0846), .ZN(new_n4868_));
  OAI21_X1   g02354(.A1(new_n4868_), .A2(new_n2522_), .B(new_n4867_), .ZN(new_n4869_));
  NAND2_X1   g02355(.A1(new_n4869_), .A2(new_n2562_), .ZN(new_n4870_));
  NAND2_X1   g02356(.A1(new_n2523_), .A2(pi0846), .ZN(new_n4871_));
  AOI21_X1   g02357(.A1(new_n3422_), .A2(new_n4867_), .B(new_n4871_), .ZN(new_n4872_));
  NAND4_X1   g02358(.A1(new_n4866_), .A2(new_n4865_), .A3(new_n4870_), .A4(new_n4872_), .ZN(new_n4873_));
  AOI21_X1   g02359(.A1(new_n4873_), .A2(new_n4858_), .B(new_n4845_), .ZN(new_n4874_));
  AOI21_X1   g02360(.A1(pi0224), .A2(pi0278), .B(pi0222), .ZN(new_n4875_));
  OAI21_X1   g02361(.A1(new_n4848_), .A2(pi0224), .B(new_n4875_), .ZN(new_n4876_));
  INV_X1     g02362(.I(new_n4876_), .ZN(new_n4877_));
  NOR2_X1    g02363(.A1(new_n2588_), .A2(pi0224), .ZN(new_n4878_));
  INV_X1     g02364(.I(new_n4878_), .ZN(new_n4879_));
  NOR3_X1    g02365(.A1(new_n4879_), .A2(new_n2553_), .A3(pi0930), .ZN(new_n4880_));
  NOR2_X1    g02366(.A1(new_n4877_), .A2(new_n4880_), .ZN(new_n4881_));
  NOR2_X1    g02367(.A1(new_n4881_), .A2(new_n2591_), .ZN(new_n4882_));
  NOR2_X1    g02368(.A1(new_n4882_), .A2(pi0299), .ZN(new_n4883_));
  NOR2_X1    g02369(.A1(new_n4883_), .A2(new_n3591_), .ZN(new_n4884_));
  AOI21_X1   g02370(.A1(new_n4884_), .A2(new_n2591_), .B(pi0299), .ZN(new_n4885_));
  INV_X1     g02371(.I(new_n4885_), .ZN(new_n4886_));
  AOI21_X1   g02372(.A1(new_n2604_), .A2(new_n4877_), .B(new_n4886_), .ZN(new_n4887_));
  INV_X1     g02373(.I(new_n4887_), .ZN(new_n4888_));
  NAND2_X1   g02374(.A1(new_n4856_), .A2(pi0299), .ZN(new_n4889_));
  NAND2_X1   g02375(.A1(new_n4888_), .A2(new_n4889_), .ZN(new_n4890_));
  AOI21_X1   g02376(.A1(new_n4890_), .A2(pi0039), .B(pi0038), .ZN(new_n4891_));
  INV_X1     g02377(.I(new_n4880_), .ZN(new_n4892_));
  OAI21_X1   g02378(.A1(new_n4868_), .A2(pi0224), .B(new_n4875_), .ZN(new_n4893_));
  NAND3_X1   g02379(.A1(new_n4893_), .A2(new_n3293_), .A3(new_n4892_), .ZN(new_n4894_));
  NAND2_X1   g02380(.A1(new_n4894_), .A2(new_n3154_), .ZN(new_n4895_));
  NOR2_X1    g02381(.A1(new_n4847_), .A2(new_n4875_), .ZN(new_n4896_));
  OAI21_X1   g02382(.A1(new_n3420_), .A2(pi0224), .B(new_n4896_), .ZN(new_n4897_));
  NOR2_X1    g02383(.A1(new_n4897_), .A2(new_n3294_), .ZN(new_n4898_));
  NOR2_X1    g02384(.A1(new_n2587_), .A2(pi0215), .ZN(new_n4899_));
  OAI21_X1   g02385(.A1(new_n4895_), .A2(new_n4898_), .B(new_n4899_), .ZN(new_n4900_));
  OR3_X2     g02386(.A1(new_n4874_), .A2(new_n4891_), .A3(new_n4900_), .Z(new_n4901_));
  NAND2_X1   g02387(.A1(new_n3252_), .A2(pi0846), .ZN(new_n4902_));
  NAND3_X1   g02388(.A1(new_n4902_), .A2(new_n2523_), .A3(new_n3255_), .ZN(new_n4903_));
  AOI21_X1   g02389(.A1(new_n4903_), .A2(new_n4851_), .B(new_n4854_), .ZN(new_n4904_));
  NOR2_X1    g02390(.A1(pi0215), .A2(pi0299), .ZN(new_n4905_));
  OAI21_X1   g02391(.A1(new_n4904_), .A2(new_n4845_), .B(new_n4905_), .ZN(new_n4906_));
  NAND3_X1   g02392(.A1(new_n4906_), .A2(new_n2544_), .A3(new_n4888_), .ZN(new_n4907_));
  INV_X1     g02393(.I(new_n4862_), .ZN(new_n4908_));
  AOI21_X1   g02394(.A1(pi0299), .A2(new_n4908_), .B(new_n4887_), .ZN(new_n4909_));
  AOI21_X1   g02395(.A1(new_n4909_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4910_));
  INV_X1     g02396(.I(new_n4909_), .ZN(new_n4911_));
  OAI21_X1   g02397(.A1(new_n4911_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n4912_));
  AOI21_X1   g02398(.A1(new_n4907_), .A2(new_n4910_), .B(new_n4912_), .ZN(new_n4913_));
  AOI21_X1   g02399(.A1(new_n4901_), .A2(new_n4913_), .B(pi0087), .ZN(new_n4914_));
  NOR2_X1    g02400(.A1(new_n4909_), .A2(new_n3197_), .ZN(new_n4915_));
  AOI21_X1   g02401(.A1(new_n3197_), .A2(new_n4890_), .B(new_n4915_), .ZN(new_n4916_));
  NOR2_X1    g02402(.A1(new_n4916_), .A2(new_n3177_), .ZN(new_n4917_));
  OAI21_X1   g02403(.A1(new_n4914_), .A2(pi0075), .B(new_n4917_), .ZN(new_n4918_));
  NOR4_X1    g02404(.A1(new_n4916_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4909_), .ZN(new_n4919_));
  AOI21_X1   g02405(.A1(new_n4909_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4920_));
  NOR2_X1    g02406(.A1(new_n4911_), .A2(new_n2628_), .ZN(new_n4921_));
  NOR4_X1    g02407(.A1(new_n4919_), .A2(new_n3330_), .A3(new_n4920_), .A4(new_n4921_), .ZN(new_n4922_));
  MUX2_X1    g02408(.I0(new_n4856_), .I1(new_n4908_), .S(new_n3336_), .Z(new_n4923_));
  NAND2_X1   g02409(.A1(new_n4856_), .A2(new_n3233_), .ZN(new_n4924_));
  AOI21_X1   g02410(.A1(new_n4908_), .A2(new_n3234_), .B(pi0055), .ZN(new_n4925_));
  AOI21_X1   g02411(.A1(new_n4924_), .A2(new_n4925_), .B(new_n3503_), .ZN(new_n4926_));
  OAI21_X1   g02412(.A1(new_n3335_), .A2(new_n4923_), .B(new_n4926_), .ZN(new_n4927_));
  AOI21_X1   g02413(.A1(new_n4918_), .A2(new_n4922_), .B(new_n4927_), .ZN(new_n4928_));
  INV_X1     g02414(.I(pi0242), .ZN(new_n4929_));
  AOI21_X1   g02415(.A1(new_n4908_), .A2(new_n4929_), .B(new_n2571_), .ZN(new_n4930_));
  OAI21_X1   g02416(.A1(new_n4928_), .A2(new_n4864_), .B(new_n4930_), .ZN(new_n4931_));
  OAI21_X1   g02417(.A1(pi0152), .A2(new_n3428_), .B(new_n3651_), .ZN(new_n4932_));
  NOR2_X1    g02418(.A1(pi0228), .A2(pi0846), .ZN(new_n4933_));
  NAND3_X1   g02419(.A1(new_n3426_), .A2(new_n3250_), .A3(new_n3428_), .ZN(new_n4934_));
  OAI21_X1   g02420(.A1(new_n3377_), .A2(pi0152), .B(new_n4846_), .ZN(new_n4935_));
  NAND4_X1   g02421(.A1(new_n4935_), .A2(new_n4932_), .A3(new_n4933_), .A4(new_n4934_), .ZN(new_n4936_));
  NOR2_X1    g02422(.A1(new_n4870_), .A2(new_n4858_), .ZN(new_n4937_));
  AOI21_X1   g02423(.A1(new_n4936_), .A2(new_n4937_), .B(new_n4845_), .ZN(new_n4938_));
  NOR2_X1    g02424(.A1(new_n4850_), .A2(new_n3282_), .ZN(new_n4939_));
  NAND2_X1   g02425(.A1(new_n4853_), .A2(new_n4939_), .ZN(new_n4940_));
  NAND2_X1   g02426(.A1(new_n4940_), .A2(new_n2562_), .ZN(new_n4941_));
  NAND2_X1   g02427(.A1(new_n4941_), .A2(new_n4858_), .ZN(new_n4942_));
  AOI21_X1   g02428(.A1(new_n4942_), .A2(new_n4857_), .B(pi0215), .ZN(new_n4943_));
  NOR2_X1    g02429(.A1(new_n4943_), .A2(new_n2587_), .ZN(new_n4944_));
  NOR2_X1    g02430(.A1(new_n4944_), .A2(new_n4885_), .ZN(new_n4945_));
  OAI21_X1   g02431(.A1(new_n4945_), .A2(new_n3154_), .B(new_n3172_), .ZN(new_n4946_));
  NAND3_X1   g02432(.A1(new_n4895_), .A2(new_n4946_), .A3(new_n4899_), .ZN(new_n4947_));
  INV_X1     g02433(.I(new_n4858_), .ZN(new_n4948_));
  NAND2_X1   g02434(.A1(new_n4903_), .A2(new_n4939_), .ZN(new_n4949_));
  AOI21_X1   g02435(.A1(new_n4949_), .A2(new_n2562_), .B(new_n4948_), .ZN(new_n4950_));
  OAI21_X1   g02436(.A1(new_n4950_), .A2(new_n4845_), .B(new_n4905_), .ZN(new_n4951_));
  NAND3_X1   g02437(.A1(new_n4951_), .A2(new_n2544_), .A3(new_n4886_), .ZN(new_n4952_));
  NOR2_X1    g02438(.A1(new_n4908_), .A2(new_n3288_), .ZN(new_n4953_));
  OAI21_X1   g02439(.A1(new_n4953_), .A2(new_n2587_), .B(new_n4886_), .ZN(new_n4954_));
  INV_X1     g02440(.I(new_n4954_), .ZN(new_n4955_));
  AOI21_X1   g02441(.A1(new_n4955_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4956_));
  OAI21_X1   g02442(.A1(new_n4954_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n4957_));
  AOI21_X1   g02443(.A1(new_n4952_), .A2(new_n4956_), .B(new_n4957_), .ZN(new_n4958_));
  OAI21_X1   g02444(.A1(new_n4938_), .A2(new_n4947_), .B(new_n4958_), .ZN(new_n4959_));
  AOI21_X1   g02445(.A1(new_n4959_), .A2(new_n3177_), .B(pi0075), .ZN(new_n4960_));
  NOR2_X1    g02446(.A1(new_n4945_), .A2(new_n3198_), .ZN(new_n4961_));
  AOI21_X1   g02447(.A1(new_n3198_), .A2(new_n4954_), .B(new_n4961_), .ZN(new_n4962_));
  OR2_X2     g02448(.A1(new_n4962_), .A2(new_n3177_), .Z(new_n4963_));
  NOR4_X1    g02449(.A1(new_n4962_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4955_), .ZN(new_n4964_));
  AOI21_X1   g02450(.A1(new_n4955_), .A2(new_n2539_), .B(pi0055), .ZN(new_n4965_));
  NOR2_X1    g02451(.A1(new_n4954_), .A2(new_n2628_), .ZN(new_n4966_));
  NOR4_X1    g02452(.A1(new_n4964_), .A2(new_n3330_), .A3(new_n4965_), .A4(new_n4966_), .ZN(new_n4967_));
  OAI21_X1   g02453(.A1(new_n4960_), .A2(new_n4963_), .B(new_n4967_), .ZN(new_n4968_));
  MUX2_X1    g02454(.I0(new_n4943_), .I1(new_n4953_), .S(new_n3336_), .Z(new_n4969_));
  NOR2_X1    g02455(.A1(new_n4943_), .A2(new_n3234_), .ZN(new_n4970_));
  OAI21_X1   g02456(.A1(new_n4953_), .A2(new_n3233_), .B(new_n3227_), .ZN(new_n4971_));
  OAI21_X1   g02457(.A1(new_n4970_), .A2(new_n4971_), .B(new_n2533_), .ZN(new_n4972_));
  AOI21_X1   g02458(.A1(pi0056), .A2(new_n4969_), .B(new_n4972_), .ZN(new_n4973_));
  NOR2_X1    g02459(.A1(new_n4943_), .A2(new_n3400_), .ZN(new_n4974_));
  OAI21_X1   g02460(.A1(new_n4953_), .A2(new_n3343_), .B(new_n3240_), .ZN(new_n4975_));
  NOR3_X1    g02461(.A1(new_n3405_), .A2(pi0242), .A3(pi1134), .ZN(new_n4976_));
  OAI21_X1   g02462(.A1(new_n4974_), .A2(new_n4975_), .B(new_n4976_), .ZN(new_n4977_));
  AOI21_X1   g02463(.A1(new_n4968_), .A2(new_n4973_), .B(new_n4977_), .ZN(new_n4978_));
  INV_X1     g02464(.I(new_n4884_), .ZN(new_n4979_));
  NAND2_X1   g02465(.A1(new_n2555_), .A2(pi0221), .ZN(new_n4980_));
  NAND2_X1   g02466(.A1(new_n4980_), .A2(new_n2566_), .ZN(new_n4981_));
  NOR2_X1    g02467(.A1(new_n4981_), .A2(new_n4845_), .ZN(new_n4982_));
  INV_X1     g02468(.I(new_n4982_), .ZN(new_n4983_));
  AOI21_X1   g02469(.A1(new_n4941_), .A2(new_n4858_), .B(new_n4983_), .ZN(new_n4984_));
  OAI21_X1   g02470(.A1(new_n4984_), .A2(new_n2587_), .B(new_n4979_), .ZN(new_n4985_));
  AOI21_X1   g02471(.A1(new_n4985_), .A2(pi0039), .B(pi0038), .ZN(new_n4986_));
  NAND2_X1   g02472(.A1(new_n4980_), .A2(new_n4899_), .ZN(new_n4987_));
  NAND2_X1   g02473(.A1(new_n4893_), .A2(new_n4892_), .ZN(new_n4988_));
  NOR2_X1    g02474(.A1(new_n2590_), .A2(new_n3294_), .ZN(new_n4989_));
  AOI21_X1   g02475(.A1(new_n4988_), .A2(new_n4989_), .B(pi0039), .ZN(new_n4990_));
  NOR3_X1    g02476(.A1(new_n4990_), .A2(new_n4986_), .A3(new_n4987_), .ZN(new_n4991_));
  NAND2_X1   g02477(.A1(new_n4938_), .A2(new_n4991_), .ZN(new_n4992_));
  OAI21_X1   g02478(.A1(new_n4950_), .A2(new_n4983_), .B(pi0299), .ZN(new_n4993_));
  NAND3_X1   g02479(.A1(new_n4993_), .A2(new_n2544_), .A3(new_n4979_), .ZN(new_n4994_));
  NAND2_X1   g02480(.A1(new_n4861_), .A2(new_n4982_), .ZN(new_n4995_));
  INV_X1     g02481(.I(new_n4995_), .ZN(new_n4996_));
  NOR2_X1    g02482(.A1(new_n4996_), .A2(new_n3288_), .ZN(new_n4997_));
  AOI21_X1   g02483(.A1(new_n4997_), .A2(pi0299), .B(new_n4884_), .ZN(new_n4998_));
  AOI21_X1   g02484(.A1(new_n4998_), .A2(new_n2545_), .B(new_n3173_), .ZN(new_n4999_));
  INV_X1     g02485(.I(new_n4998_), .ZN(new_n5000_));
  OAI21_X1   g02486(.A1(new_n5000_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n5001_));
  AOI21_X1   g02487(.A1(new_n4994_), .A2(new_n4999_), .B(new_n5001_), .ZN(new_n5002_));
  AOI21_X1   g02488(.A1(new_n4992_), .A2(new_n5002_), .B(pi0087), .ZN(new_n5003_));
  NOR2_X1    g02489(.A1(new_n4998_), .A2(new_n3197_), .ZN(new_n5004_));
  AOI21_X1   g02490(.A1(new_n3197_), .A2(new_n4985_), .B(new_n5004_), .ZN(new_n5005_));
  NOR2_X1    g02491(.A1(new_n5005_), .A2(new_n3177_), .ZN(new_n5006_));
  OAI21_X1   g02492(.A1(new_n5003_), .A2(pi0075), .B(new_n5006_), .ZN(new_n5007_));
  NOR4_X1    g02493(.A1(new_n5005_), .A2(pi0092), .A3(new_n2535_), .A4(new_n4998_), .ZN(new_n5008_));
  OAI21_X1   g02494(.A1(new_n5000_), .A2(new_n2628_), .B(new_n3203_), .ZN(new_n5009_));
  NOR2_X1    g02495(.A1(new_n5008_), .A2(new_n5009_), .ZN(new_n5010_));
  OAI21_X1   g02496(.A1(new_n5000_), .A2(new_n2538_), .B(new_n3227_), .ZN(new_n5011_));
  NAND3_X1   g02497(.A1(new_n5011_), .A2(pi0056), .A3(new_n2539_), .ZN(new_n5012_));
  AOI21_X1   g02498(.A1(new_n5007_), .A2(new_n5010_), .B(new_n5012_), .ZN(new_n5013_));
  INV_X1     g02499(.I(new_n4997_), .ZN(new_n5014_));
  NAND4_X1   g02500(.A1(new_n4984_), .A2(new_n5014_), .A3(new_n3335_), .A4(new_n2548_), .ZN(new_n5015_));
  NAND2_X1   g02501(.A1(new_n5015_), .A2(new_n3406_), .ZN(new_n5016_));
  AOI21_X1   g02502(.A1(new_n5014_), .A2(new_n3405_), .B(new_n4929_), .ZN(new_n5017_));
  OAI21_X1   g02503(.A1(new_n5013_), .A2(new_n5016_), .B(new_n5017_), .ZN(new_n5018_));
  NOR2_X1    g02504(.A1(new_n4855_), .A2(new_n4983_), .ZN(new_n5019_));
  OAI21_X1   g02505(.A1(new_n4881_), .A2(new_n2591_), .B(new_n2587_), .ZN(new_n5020_));
  AOI21_X1   g02506(.A1(new_n5020_), .A2(pi0039), .B(pi0038), .ZN(new_n5021_));
  AOI21_X1   g02507(.A1(new_n4897_), .A2(new_n4892_), .B(new_n4989_), .ZN(new_n5022_));
  NOR4_X1    g02508(.A1(new_n5022_), .A2(pi0039), .A3(new_n4987_), .A4(new_n5021_), .ZN(new_n5023_));
  NOR3_X1    g02509(.A1(new_n4882_), .A2(pi0299), .A3(new_n2545_), .ZN(new_n5024_));
  NOR2_X1    g02510(.A1(new_n4882_), .A2(pi0299), .ZN(new_n5025_));
  INV_X1     g02511(.I(new_n5025_), .ZN(new_n5026_));
  OAI21_X1   g02512(.A1(new_n5026_), .A2(new_n2544_), .B(pi0100), .ZN(new_n5027_));
  AOI21_X1   g02513(.A1(new_n5025_), .A2(pi0038), .B(pi0100), .ZN(new_n5028_));
  OAI21_X1   g02514(.A1(new_n5027_), .A2(new_n5024_), .B(new_n5028_), .ZN(new_n5029_));
  AOI21_X1   g02515(.A1(new_n4874_), .A2(new_n5023_), .B(new_n5029_), .ZN(new_n5030_));
  OAI21_X1   g02516(.A1(new_n5030_), .A2(pi0087), .B(new_n2628_), .ZN(new_n5031_));
  NAND2_X1   g02517(.A1(new_n5020_), .A2(new_n3197_), .ZN(new_n5032_));
  NAND2_X1   g02518(.A1(new_n5026_), .A2(new_n3198_), .ZN(new_n5033_));
  AOI21_X1   g02519(.A1(new_n5033_), .A2(new_n5032_), .B(new_n3177_), .ZN(new_n5034_));
  NAND2_X1   g02520(.A1(new_n5033_), .A2(new_n5032_), .ZN(new_n5035_));
  NAND4_X1   g02521(.A1(new_n5035_), .A2(new_n3203_), .A3(new_n2534_), .A4(new_n5026_), .ZN(new_n5036_));
  OAI21_X1   g02522(.A1(new_n5026_), .A2(new_n2538_), .B(new_n3227_), .ZN(new_n5037_));
  NAND2_X1   g02523(.A1(new_n5025_), .A2(pi0075), .ZN(new_n5038_));
  NAND4_X1   g02524(.A1(new_n5036_), .A2(new_n3329_), .A3(new_n5037_), .A4(new_n5038_), .ZN(new_n5039_));
  AOI21_X1   g02525(.A1(new_n5031_), .A2(new_n5034_), .B(new_n5039_), .ZN(new_n5040_));
  INV_X1     g02526(.I(new_n5019_), .ZN(new_n5041_));
  MUX2_X1    g02527(.I0(new_n5041_), .I1(new_n4995_), .S(new_n3336_), .Z(new_n5042_));
  NAND2_X1   g02528(.A1(new_n5041_), .A2(new_n3233_), .ZN(new_n5043_));
  AOI21_X1   g02529(.A1(new_n4995_), .A2(new_n3234_), .B(pi0055), .ZN(new_n5044_));
  AOI21_X1   g02530(.A1(new_n5043_), .A2(new_n5044_), .B(new_n3503_), .ZN(new_n5045_));
  OAI21_X1   g02531(.A1(new_n3335_), .A2(new_n5042_), .B(new_n5045_), .ZN(new_n5046_));
  NAND2_X1   g02532(.A1(new_n5041_), .A2(new_n3343_), .ZN(new_n5047_));
  AOI21_X1   g02533(.A1(new_n3400_), .A2(new_n4995_), .B(pi0062), .ZN(new_n5048_));
  AOI21_X1   g02534(.A1(new_n5047_), .A2(new_n5048_), .B(new_n3405_), .ZN(new_n5049_));
  OAI21_X1   g02535(.A1(new_n5040_), .A2(new_n5046_), .B(new_n5049_), .ZN(new_n5050_));
  AOI21_X1   g02536(.A1(new_n4996_), .A2(new_n3405_), .B(pi0242), .ZN(new_n5051_));
  AOI21_X1   g02537(.A1(new_n5050_), .A2(new_n5051_), .B(pi1134), .ZN(new_n5052_));
  AOI22_X1   g02538(.A1(new_n4931_), .A2(new_n4978_), .B1(new_n5018_), .B2(new_n5052_), .ZN(po0165));
  INV_X1     g02539(.I(pi0057), .ZN(new_n5055_));
  NOR2_X1    g02540(.A1(new_n3162_), .A2(new_n3198_), .ZN(new_n5056_));
  AOI21_X1   g02541(.A1(new_n5056_), .A2(new_n2542_), .B(new_n3335_), .ZN(new_n5057_));
  AOI21_X1   g02542(.A1(new_n2669_), .A2(new_n2902_), .B(new_n2841_), .ZN(new_n5058_));
  INV_X1     g02543(.I(new_n5058_), .ZN(new_n5059_));
  NAND3_X1   g02544(.A1(new_n2813_), .A2(new_n2682_), .A3(new_n2684_), .ZN(new_n5060_));
  AOI21_X1   g02545(.A1(new_n5060_), .A2(new_n2821_), .B(new_n2689_), .ZN(new_n5061_));
  INV_X1     g02546(.I(pi0108), .ZN(new_n5062_));
  NOR2_X1    g02547(.A1(new_n2828_), .A2(new_n5062_), .ZN(new_n5063_));
  NOR3_X1    g02548(.A1(new_n2833_), .A2(pi0108), .A3(pi0110), .ZN(new_n5064_));
  OAI21_X1   g02549(.A1(pi0046), .A2(new_n5063_), .B(new_n5064_), .ZN(new_n5065_));
  NOR2_X1    g02550(.A1(new_n2835_), .A2(new_n2679_), .ZN(new_n5066_));
  OAI21_X1   g02551(.A1(new_n5061_), .A2(new_n5065_), .B(new_n5066_), .ZN(new_n5067_));
  NOR2_X1    g02552(.A1(new_n2459_), .A2(new_n2476_), .ZN(new_n5068_));
  AOI21_X1   g02553(.A1(new_n5068_), .A2(pi0058), .B(pi0090), .ZN(new_n5069_));
  INV_X1     g02554(.I(new_n5069_), .ZN(new_n5070_));
  NOR2_X1    g02555(.A1(new_n2843_), .A2(new_n2638_), .ZN(new_n5071_));
  NAND2_X1   g02556(.A1(new_n5071_), .A2(new_n5070_), .ZN(new_n5072_));
  AOI21_X1   g02557(.A1(new_n5067_), .A2(new_n2661_), .B(new_n5072_), .ZN(new_n5073_));
  OAI21_X1   g02558(.A1(new_n5073_), .A2(new_n2840_), .B(new_n2841_), .ZN(new_n5074_));
  NAND2_X1   g02559(.A1(new_n5074_), .A2(new_n5059_), .ZN(new_n5075_));
  MUX2_X1    g02560(.I0(new_n5075_), .I1(new_n2851_), .S(pi0035), .Z(new_n5076_));
  AOI21_X1   g02561(.A1(new_n5076_), .A2(new_n2849_), .B(pi0051), .ZN(new_n5077_));
  NOR3_X1    g02562(.A1(new_n5077_), .A2(new_n2676_), .A3(new_n3105_), .ZN(new_n5078_));
  NOR2_X1    g02563(.A1(new_n2601_), .A2(pi0299), .ZN(new_n5079_));
  AOI21_X1   g02564(.A1(pi0210), .A2(pi0299), .B(new_n5079_), .ZN(new_n5080_));
  INV_X1     g02565(.I(new_n5080_), .ZN(new_n5081_));
  NOR2_X1    g02566(.A1(new_n2507_), .A2(pi0035), .ZN(new_n5082_));
  INV_X1     g02567(.I(new_n5082_), .ZN(new_n5083_));
  NOR3_X1    g02568(.A1(new_n2904_), .A2(pi0040), .A3(new_n5083_), .ZN(new_n5084_));
  AOI21_X1   g02569(.A1(new_n3363_), .A2(new_n5081_), .B(pi0032), .ZN(new_n5085_));
  OAI21_X1   g02570(.A1(new_n5081_), .A2(new_n5084_), .B(new_n5085_), .ZN(new_n5086_));
  AND2_X2    g02571(.A1(new_n5086_), .A2(new_n2437_), .Z(new_n5087_));
  OAI21_X1   g02572(.A1(new_n5078_), .A2(new_n3008_), .B(new_n5087_), .ZN(new_n5088_));
  NOR4_X1    g02573(.A1(pi0970), .A2(pi0972), .A3(pi0975), .A4(pi0978), .ZN(new_n5089_));
  NOR3_X1    g02574(.A1(new_n5089_), .A2(pi0960), .A3(pi0963), .ZN(new_n5090_));
  INV_X1     g02575(.I(new_n5090_), .ZN(new_n5091_));
  NOR2_X1    g02576(.A1(pi0907), .A2(pi0947), .ZN(new_n5092_));
  INV_X1     g02577(.I(new_n5092_), .ZN(new_n5093_));
  NOR2_X1    g02578(.A1(new_n5091_), .A2(new_n5093_), .ZN(new_n5094_));
  INV_X1     g02579(.I(pi0680), .ZN(new_n5095_));
  NOR2_X1    g02580(.A1(new_n5095_), .A2(pi0662), .ZN(new_n5096_));
  INV_X1     g02581(.I(new_n5096_), .ZN(new_n5097_));
  NOR2_X1    g02582(.A1(new_n5097_), .A2(pi0661), .ZN(new_n5098_));
  INV_X1     g02583(.I(new_n5098_), .ZN(new_n5099_));
  NOR2_X1    g02584(.A1(new_n5099_), .A2(pi0681), .ZN(new_n5100_));
  INV_X1     g02585(.I(pi0603), .ZN(new_n5101_));
  NOR2_X1    g02586(.A1(new_n5101_), .A2(pi0642), .ZN(new_n5102_));
  INV_X1     g02587(.I(new_n5102_), .ZN(new_n5103_));
  NOR2_X1    g02588(.A1(pi0614), .A2(pi0616), .ZN(new_n5104_));
  INV_X1     g02589(.I(new_n5104_), .ZN(new_n5105_));
  NOR2_X1    g02590(.A1(new_n5103_), .A2(new_n5105_), .ZN(new_n5106_));
  NOR2_X1    g02591(.A1(new_n5100_), .A2(new_n5106_), .ZN(new_n5107_));
  NOR2_X1    g02592(.A1(pi0332), .A2(pi0468), .ZN(new_n5108_));
  INV_X1     g02593(.I(new_n5108_), .ZN(new_n5109_));
  NOR2_X1    g02594(.A1(new_n3162_), .A2(new_n5109_), .ZN(new_n5110_));
  INV_X1     g02595(.I(new_n5110_), .ZN(new_n5111_));
  INV_X1     g02596(.I(new_n5107_), .ZN(po1101));
  NOR2_X1    g02597(.A1(new_n2921_), .A2(new_n2924_), .ZN(new_n5113_));
  NOR2_X1    g02598(.A1(pi0824), .A2(pi0829), .ZN(new_n5114_));
  NAND3_X1   g02599(.A1(new_n5114_), .A2(pi0824), .A3(new_n2918_), .ZN(new_n5115_));
  NOR2_X1    g02600(.A1(new_n5113_), .A2(new_n5115_), .ZN(new_n5116_));
  INV_X1     g02601(.I(new_n5116_), .ZN(new_n5117_));
  INV_X1     g02602(.I(pi0835), .ZN(new_n5118_));
  INV_X1     g02603(.I(pi0979), .ZN(new_n5119_));
  NAND2_X1   g02604(.A1(pi0835), .A2(pi0984), .ZN(new_n5120_));
  INV_X1     g02605(.I(pi1001), .ZN(new_n5121_));
  NAND2_X1   g02606(.A1(new_n3181_), .A2(new_n5121_), .ZN(new_n5122_));
  NAND3_X1   g02607(.A1(new_n5122_), .A2(new_n5119_), .A3(new_n5120_), .ZN(new_n5123_));
  NOR4_X1    g02608(.A1(new_n5123_), .A2(pi0287), .A3(new_n5118_), .A4(new_n2928_), .ZN(new_n5124_));
  INV_X1     g02609(.I(new_n5124_), .ZN(new_n5125_));
  NOR3_X1    g02610(.A1(new_n5117_), .A2(new_n2923_), .A3(new_n5125_), .ZN(new_n5126_));
  OAI21_X1   g02611(.A1(new_n5126_), .A2(new_n5108_), .B(po1101), .ZN(new_n5127_));
  OAI22_X1   g02612(.A1(new_n5111_), .A2(new_n5107_), .B1(new_n2490_), .B2(new_n5127_), .ZN(new_n5128_));
  INV_X1     g02613(.I(new_n5126_), .ZN(new_n5129_));
  NOR2_X1    g02614(.A1(po1101), .A2(new_n5108_), .ZN(new_n5130_));
  OAI21_X1   g02615(.A1(new_n5130_), .A2(new_n5129_), .B(new_n2490_), .ZN(new_n5131_));
  NAND4_X1   g02616(.A1(new_n5128_), .A2(new_n2566_), .A3(new_n5094_), .A4(new_n5131_), .ZN(new_n5132_));
  AOI21_X1   g02617(.A1(new_n5094_), .A2(new_n5108_), .B(new_n5130_), .ZN(new_n5133_));
  NOR2_X1    g02618(.A1(new_n3082_), .A2(new_n5125_), .ZN(new_n5134_));
  NAND4_X1   g02619(.A1(new_n5133_), .A2(pi0216), .A3(pi0221), .A4(new_n5134_), .ZN(new_n5135_));
  NAND2_X1   g02620(.A1(new_n5135_), .A2(new_n2490_), .ZN(new_n5136_));
  AOI21_X1   g02621(.A1(new_n5136_), .A2(new_n2566_), .B(new_n2587_), .ZN(new_n5137_));
  AOI21_X1   g02622(.A1(new_n5132_), .A2(new_n5137_), .B(new_n3154_), .ZN(new_n5138_));
  NOR4_X1    g02623(.A1(pi0969), .A2(pi0971), .A3(pi0974), .A4(pi0977), .ZN(new_n5139_));
  NOR4_X1    g02624(.A1(pi0587), .A2(pi0602), .A3(pi0961), .A4(pi0967), .ZN(new_n5140_));
  NOR2_X1    g02625(.A1(new_n5139_), .A2(new_n5140_), .ZN(new_n5141_));
  NAND4_X1   g02626(.A1(new_n5128_), .A2(new_n2604_), .A3(new_n5131_), .A4(new_n5141_), .ZN(new_n5142_));
  NOR2_X1    g02627(.A1(new_n5107_), .A2(new_n5108_), .ZN(new_n5143_));
  NOR2_X1    g02628(.A1(new_n5141_), .A2(new_n5109_), .ZN(new_n5144_));
  NOR2_X1    g02629(.A1(new_n5143_), .A2(new_n5144_), .ZN(new_n5145_));
  INV_X1     g02630(.I(new_n5145_), .ZN(new_n5146_));
  NAND4_X1   g02631(.A1(new_n5146_), .A2(pi0222), .A3(pi0224), .A4(new_n5134_), .ZN(new_n5147_));
  NAND2_X1   g02632(.A1(new_n5147_), .A2(new_n2490_), .ZN(new_n5148_));
  AOI21_X1   g02633(.A1(new_n5148_), .A2(new_n2604_), .B(pi0299), .ZN(new_n5149_));
  NAND2_X1   g02634(.A1(new_n5142_), .A2(new_n5149_), .ZN(new_n5150_));
  OAI21_X1   g02635(.A1(new_n5138_), .A2(new_n5150_), .B(new_n3154_), .ZN(new_n5151_));
  AOI21_X1   g02636(.A1(new_n5088_), .A2(new_n2872_), .B(new_n5151_), .ZN(new_n5152_));
  NOR2_X1    g02637(.A1(new_n3162_), .A2(pi0039), .ZN(new_n5153_));
  INV_X1     g02638(.I(new_n5153_), .ZN(new_n5154_));
  MUX2_X1    g02639(.I0(new_n5154_), .I1(new_n5152_), .S(new_n3172_), .Z(new_n5155_));
  NOR2_X1    g02640(.A1(new_n2491_), .A2(pi0039), .ZN(new_n5156_));
  INV_X1     g02641(.I(new_n5156_), .ZN(new_n5157_));
  NOR2_X1    g02642(.A1(new_n3173_), .A2(pi0038), .ZN(new_n5158_));
  INV_X1     g02643(.I(new_n5158_), .ZN(new_n5159_));
  NOR2_X1    g02644(.A1(new_n5157_), .A2(new_n5159_), .ZN(new_n5160_));
  NOR2_X1    g02645(.A1(new_n2605_), .A2(pi0142), .ZN(new_n5161_));
  NOR2_X1    g02646(.A1(new_n5161_), .A2(pi0299), .ZN(new_n5162_));
  AOI21_X1   g02647(.A1(new_n3025_), .A2(pi0299), .B(new_n5162_), .ZN(new_n5163_));
  NOR4_X1    g02648(.A1(pi0113), .A2(pi0114), .A3(pi0115), .A4(pi0116), .ZN(new_n5164_));
  NOR2_X1    g02649(.A1(pi0042), .A2(pi0043), .ZN(new_n5165_));
  INV_X1     g02650(.I(new_n5165_), .ZN(new_n5166_));
  NOR2_X1    g02651(.A1(new_n5166_), .A2(pi0052), .ZN(new_n5167_));
  INV_X1     g02652(.I(new_n5167_), .ZN(new_n5168_));
  NOR2_X1    g02653(.A1(new_n5168_), .A2(new_n5164_), .ZN(new_n5169_));
  INV_X1     g02654(.I(new_n5169_), .ZN(new_n5170_));
  NOR2_X1    g02655(.A1(pi0041), .A2(pi0099), .ZN(new_n5171_));
  INV_X1     g02656(.I(new_n5171_), .ZN(new_n5172_));
  NOR2_X1    g02657(.A1(new_n5172_), .A2(pi0101), .ZN(new_n5173_));
  INV_X1     g02658(.I(new_n5173_), .ZN(new_n5174_));
  NOR2_X1    g02659(.A1(new_n5170_), .A2(new_n5174_), .ZN(new_n5175_));
  INV_X1     g02660(.I(new_n5175_), .ZN(new_n5176_));
  NOR2_X1    g02661(.A1(new_n5176_), .A2(pi0044), .ZN(new_n5177_));
  INV_X1     g02662(.I(pi0683), .ZN(new_n5178_));
  INV_X1     g02663(.I(new_n5177_), .ZN(po1057));
  INV_X1     g02664(.I(pi0250), .ZN(new_n5180_));
  NOR2_X1    g02665(.A1(new_n5114_), .A2(new_n2955_), .ZN(new_n5181_));
  INV_X1     g02666(.I(new_n5181_), .ZN(new_n5182_));
  NOR2_X1    g02667(.A1(new_n5182_), .A2(pi1093), .ZN(po0740));
  NOR2_X1    g02668(.A1(new_n5180_), .A2(pi0129), .ZN(new_n5184_));
  AOI21_X1   g02669(.A1(po0740), .A2(new_n5180_), .B(new_n5184_), .ZN(new_n5185_));
  INV_X1     g02670(.I(new_n5185_), .ZN(new_n5186_));
  AOI21_X1   g02671(.A1(po1057), .A2(new_n5178_), .B(new_n5186_), .ZN(new_n5187_));
  OR3_X2     g02672(.A1(new_n5160_), .A2(new_n3245_), .A3(new_n5163_), .Z(new_n5188_));
  NAND2_X1   g02673(.A1(new_n5188_), .A2(new_n3177_), .ZN(new_n5189_));
  NOR3_X1    g02674(.A1(new_n5155_), .A2(pi0100), .A3(new_n5189_), .ZN(new_n5190_));
  NOR2_X1    g02675(.A1(new_n5056_), .A2(new_n3177_), .ZN(new_n5191_));
  NOR2_X1    g02676(.A1(new_n5191_), .A2(pi0075), .ZN(new_n5192_));
  NOR2_X1    g02677(.A1(pi0054), .A2(pi0092), .ZN(new_n5193_));
  NAND2_X1   g02678(.A1(new_n5192_), .A2(new_n5193_), .ZN(new_n5194_));
  INV_X1     g02679(.I(new_n5056_), .ZN(new_n5195_));
  NOR2_X1    g02680(.A1(new_n2537_), .A2(pi0054), .ZN(new_n5196_));
  INV_X1     g02681(.I(new_n5196_), .ZN(new_n5197_));
  NOR3_X1    g02682(.A1(new_n5195_), .A2(pi0074), .A3(new_n5197_), .ZN(new_n5198_));
  NOR2_X1    g02683(.A1(new_n5198_), .A2(pi0055), .ZN(new_n5199_));
  NOR2_X1    g02684(.A1(new_n5199_), .A2(pi0074), .ZN(new_n5200_));
  OAI21_X1   g02685(.A1(new_n5190_), .A2(new_n5194_), .B(new_n5200_), .ZN(new_n5201_));
  AOI21_X1   g02686(.A1(new_n5201_), .A2(new_n3335_), .B(new_n5057_), .ZN(new_n5202_));
  NOR2_X1    g02687(.A1(new_n3405_), .A2(pi0062), .ZN(new_n5203_));
  INV_X1     g02688(.I(new_n5203_), .ZN(new_n5204_));
  INV_X1     g02689(.I(pi0059), .ZN(new_n5205_));
  NOR2_X1    g02690(.A1(new_n5055_), .A2(new_n5205_), .ZN(new_n5206_));
  OR3_X2     g02691(.A1(new_n3336_), .A2(new_n3503_), .A3(new_n5206_), .Z(new_n5207_));
  OAI21_X1   g02692(.A1(new_n5207_), .A2(new_n2491_), .B(new_n3405_), .ZN(new_n5208_));
  INV_X1     g02693(.I(new_n5208_), .ZN(new_n5209_));
  OAI22_X1   g02694(.A1(new_n5202_), .A2(new_n5204_), .B1(new_n5055_), .B2(new_n5209_), .ZN(po0167));
  INV_X1     g02695(.I(pi1090), .ZN(po0170));
  NAND3_X1   g02696(.A1(new_n3233_), .A2(new_n2490_), .A3(new_n2523_), .ZN(new_n5212_));
  INV_X1     g02697(.I(pi0030), .ZN(new_n5213_));
  NOR2_X1    g02698(.A1(new_n5213_), .A2(new_n2523_), .ZN(new_n5214_));
  INV_X1     g02699(.I(new_n5214_), .ZN(new_n5215_));
  XOR2_X1    g02700(.A1(new_n5212_), .A2(new_n5215_), .Z(new_n5216_));
  INV_X1     g02701(.I(new_n5100_), .ZN(new_n5217_));
  NOR2_X1    g02702(.A1(new_n5217_), .A2(new_n5108_), .ZN(new_n5218_));
  AOI21_X1   g02703(.A1(pi0907), .A2(new_n5108_), .B(new_n5218_), .ZN(new_n5219_));
  INV_X1     g02704(.I(new_n5219_), .ZN(new_n5220_));
  NAND2_X1   g02705(.A1(new_n5216_), .A2(new_n5220_), .ZN(new_n5221_));
  NOR2_X1    g02706(.A1(new_n3503_), .A2(pi0055), .ZN(new_n5222_));
  NAND2_X1   g02707(.A1(new_n5222_), .A2(new_n5205_), .ZN(new_n5223_));
  INV_X1     g02708(.I(new_n5223_), .ZN(new_n5224_));
  OAI21_X1   g02709(.A1(new_n5224_), .A2(pi0228), .B(pi0057), .ZN(new_n5225_));
  NOR2_X1    g02710(.A1(new_n3228_), .A2(pi0054), .ZN(new_n5226_));
  AOI21_X1   g02711(.A1(pi0602), .A2(new_n5108_), .B(new_n5218_), .ZN(new_n5227_));
  MUX2_X1    g02712(.I0(new_n5227_), .I1(new_n5219_), .S(pi0299), .Z(new_n5228_));
  NOR2_X1    g02713(.A1(new_n5228_), .A2(new_n5215_), .ZN(new_n5229_));
  NOR2_X1    g02714(.A1(new_n5229_), .A2(new_n5226_), .ZN(new_n5230_));
  AOI21_X1   g02715(.A1(new_n3311_), .A2(new_n5215_), .B(pi0039), .ZN(new_n5231_));
  INV_X1     g02716(.I(new_n5231_), .ZN(new_n5232_));
  NOR2_X1    g02717(.A1(new_n5232_), .A2(new_n5228_), .ZN(new_n5233_));
  AOI22_X1   g02718(.A1(new_n5233_), .A2(new_n3207_), .B1(new_n2629_), .B2(new_n5229_), .ZN(new_n5234_));
  INV_X1     g02719(.I(new_n5234_), .ZN(new_n5235_));
  AOI21_X1   g02720(.A1(new_n5235_), .A2(new_n5226_), .B(new_n5230_), .ZN(new_n5236_));
  OAI21_X1   g02721(.A1(new_n5236_), .A2(pi0074), .B(new_n3227_), .ZN(new_n5237_));
  INV_X1     g02722(.I(new_n5227_), .ZN(new_n5238_));
  INV_X1     g02723(.I(new_n2665_), .ZN(new_n5239_));
  NAND4_X1   g02724(.A1(new_n5068_), .A2(new_n2841_), .A3(new_n2902_), .A4(new_n2479_), .ZN(new_n5240_));
  NOR3_X1    g02725(.A1(new_n5240_), .A2(new_n5239_), .A3(new_n2963_), .ZN(new_n5241_));
  INV_X1     g02726(.I(new_n5241_), .ZN(new_n5242_));
  NOR4_X1    g02727(.A1(new_n5242_), .A2(new_n2632_), .A3(pi0095), .A4(pi0198), .ZN(new_n5243_));
  INV_X1     g02728(.I(new_n5243_), .ZN(new_n5244_));
  NOR2_X1    g02729(.A1(new_n2862_), .A2(new_n2515_), .ZN(new_n5245_));
  NOR2_X1    g02730(.A1(new_n2679_), .A2(new_n2678_), .ZN(new_n5246_));
  NOR3_X1    g02731(.A1(new_n2823_), .A2(pi0046), .A3(new_n2831_), .ZN(new_n5247_));
  NAND2_X1   g02732(.A1(new_n2455_), .A2(new_n2454_), .ZN(po1049));
  NOR2_X1    g02733(.A1(new_n2794_), .A2(po1049), .ZN(new_n5249_));
  INV_X1     g02734(.I(pi0071), .ZN(new_n5250_));
  NOR2_X1    g02735(.A1(new_n2762_), .A2(new_n2766_), .ZN(new_n5251_));
  NAND2_X1   g02736(.A1(new_n2751_), .A2(pi0085), .ZN(new_n5252_));
  NAND2_X1   g02737(.A1(new_n5252_), .A2(pi0073), .ZN(new_n5253_));
  XOR2_X1    g02738(.A1(new_n5253_), .A2(new_n2759_), .Z(new_n5254_));
  NAND2_X1   g02739(.A1(new_n5254_), .A2(new_n2731_), .ZN(new_n5255_));
  OAI21_X1   g02740(.A1(new_n5255_), .A2(new_n2730_), .B(pi0084), .ZN(new_n5256_));
  AOI21_X1   g02741(.A1(new_n2730_), .A2(new_n5255_), .B(new_n5256_), .ZN(new_n5257_));
  XOR2_X1    g02742(.A1(new_n5257_), .A2(new_n2762_), .Z(new_n5258_));
  NAND2_X1   g02743(.A1(new_n5258_), .A2(new_n2757_), .ZN(new_n5259_));
  XNOR2_X1   g02744(.A1(new_n5259_), .A2(new_n5251_), .ZN(new_n5260_));
  NAND2_X1   g02745(.A1(new_n5260_), .A2(new_n2775_), .ZN(new_n5261_));
  AOI21_X1   g02746(.A1(new_n5261_), .A2(new_n2765_), .B(new_n2769_), .ZN(new_n5262_));
  NOR2_X1    g02747(.A1(new_n2780_), .A2(new_n2768_), .ZN(new_n5263_));
  NOR2_X1    g02748(.A1(new_n5262_), .A2(new_n5263_), .ZN(new_n5264_));
  OAI21_X1   g02749(.A1(new_n2789_), .A2(new_n2788_), .B(new_n2785_), .ZN(new_n5265_));
  OAI21_X1   g02750(.A1(new_n5264_), .A2(new_n5265_), .B(new_n5250_), .ZN(new_n5266_));
  AOI21_X1   g02751(.A1(new_n5266_), .A2(new_n5249_), .B(pi0081), .ZN(new_n5267_));
  NOR4_X1    g02752(.A1(new_n2721_), .A2(pi0081), .A3(new_n2452_), .A4(new_n2457_), .ZN(new_n5268_));
  NAND3_X1   g02753(.A1(new_n5268_), .A2(new_n2462_), .A3(new_n2698_), .ZN(new_n5269_));
  NOR3_X1    g02754(.A1(new_n2706_), .A2(new_n2708_), .A3(new_n5269_), .ZN(new_n5270_));
  AOI21_X1   g02755(.A1(new_n5267_), .A2(new_n5270_), .B(new_n2697_), .ZN(new_n5271_));
  OAI21_X1   g02756(.A1(new_n5271_), .A2(new_n2694_), .B(new_n2691_), .ZN(new_n5272_));
  NAND2_X1   g02757(.A1(new_n5272_), .A2(new_n5247_), .ZN(new_n5273_));
  NAND2_X1   g02758(.A1(new_n5273_), .A2(new_n2833_), .ZN(new_n5274_));
  AOI21_X1   g02759(.A1(new_n5274_), .A2(new_n5246_), .B(pi0091), .ZN(new_n5275_));
  INV_X1     g02760(.I(pi0314), .ZN(new_n5276_));
  NAND2_X1   g02761(.A1(new_n2660_), .A2(new_n5276_), .ZN(new_n5277_));
  INV_X1     g02762(.I(new_n5247_), .ZN(new_n5278_));
  INV_X1     g02763(.I(new_n2706_), .ZN(new_n5279_));
  NAND4_X1   g02764(.A1(new_n5267_), .A2(new_n2796_), .A3(new_n5249_), .A4(new_n5269_), .ZN(new_n5280_));
  NAND4_X1   g02765(.A1(new_n5280_), .A2(new_n2697_), .A3(new_n5279_), .A4(new_n2708_), .ZN(new_n5281_));
  OAI21_X1   g02766(.A1(new_n2692_), .A2(new_n2693_), .B(new_n5281_), .ZN(new_n5282_));
  NAND3_X1   g02767(.A1(new_n5282_), .A2(new_n2691_), .A3(new_n5278_), .ZN(new_n5283_));
  INV_X1     g02768(.I(new_n5246_), .ZN(new_n5284_));
  AOI21_X1   g02769(.A1(new_n5283_), .A2(new_n2833_), .B(new_n5284_), .ZN(new_n5285_));
  AOI21_X1   g02770(.A1(new_n2843_), .A2(pi0091), .B(pi0058), .ZN(new_n5286_));
  NOR2_X1    g02771(.A1(new_n5286_), .A2(pi0314), .ZN(new_n5287_));
  OAI21_X1   g02772(.A1(new_n5285_), .A2(new_n5277_), .B(new_n5287_), .ZN(new_n5288_));
  OAI21_X1   g02773(.A1(new_n5288_), .A2(new_n5275_), .B(pi0090), .ZN(new_n5289_));
  NOR2_X1    g02774(.A1(new_n2902_), .A2(pi0093), .ZN(new_n5290_));
  AOI21_X1   g02775(.A1(new_n2669_), .A2(new_n5290_), .B(pi0035), .ZN(new_n5291_));
  OAI21_X1   g02776(.A1(new_n2642_), .A2(new_n2839_), .B(new_n2841_), .ZN(new_n5292_));
  NOR2_X1    g02777(.A1(new_n5292_), .A2(new_n5291_), .ZN(new_n5293_));
  AOI21_X1   g02778(.A1(new_n5289_), .A2(new_n5293_), .B(pi0070), .ZN(new_n5294_));
  OAI21_X1   g02779(.A1(new_n5294_), .A2(new_n3066_), .B(new_n2861_), .ZN(new_n5295_));
  NAND2_X1   g02780(.A1(new_n5295_), .A2(new_n5245_), .ZN(new_n5296_));
  NAND2_X1   g02781(.A1(new_n5296_), .A2(new_n3100_), .ZN(new_n5297_));
  NAND2_X1   g02782(.A1(new_n5297_), .A2(new_n5244_), .ZN(new_n5298_));
  NOR2_X1    g02783(.A1(new_n5298_), .A2(pi0228), .ZN(new_n5299_));
  NOR2_X1    g02784(.A1(new_n2523_), .A2(pi0030), .ZN(new_n5300_));
  NOR2_X1    g02785(.A1(new_n5299_), .A2(new_n5300_), .ZN(new_n5301_));
  AOI21_X1   g02786(.A1(new_n5301_), .A2(new_n5238_), .B(pi0299), .ZN(new_n5302_));
  INV_X1     g02787(.I(new_n5286_), .ZN(new_n5303_));
  INV_X1     g02788(.I(new_n2639_), .ZN(new_n5304_));
  INV_X1     g02789(.I(new_n2832_), .ZN(new_n5305_));
  AOI21_X1   g02790(.A1(new_n5273_), .A2(new_n5305_), .B(new_n5304_), .ZN(new_n5306_));
  NOR3_X1    g02791(.A1(new_n5306_), .A2(pi0091), .A3(new_n5276_), .ZN(new_n5307_));
  NAND2_X1   g02792(.A1(new_n5283_), .A2(new_n5305_), .ZN(new_n5308_));
  AOI21_X1   g02793(.A1(new_n5308_), .A2(new_n2639_), .B(new_n5277_), .ZN(new_n5309_));
  OAI21_X1   g02794(.A1(new_n5309_), .A2(new_n5307_), .B(new_n5303_), .ZN(new_n5310_));
  NOR2_X1    g02795(.A1(new_n2840_), .A2(pi0090), .ZN(new_n5311_));
  NAND2_X1   g02796(.A1(new_n5310_), .A2(new_n5311_), .ZN(new_n5312_));
  NAND3_X1   g02797(.A1(new_n5312_), .A2(new_n2841_), .A3(new_n5291_), .ZN(new_n5313_));
  AOI21_X1   g02798(.A1(new_n5313_), .A2(new_n2849_), .B(new_n3066_), .ZN(new_n5314_));
  NOR2_X1    g02799(.A1(new_n2515_), .A2(pi0072), .ZN(new_n5315_));
  INV_X1     g02800(.I(new_n5315_), .ZN(new_n5316_));
  OAI21_X1   g02801(.A1(new_n5314_), .A2(new_n5316_), .B(new_n3100_), .ZN(new_n5317_));
  OAI21_X1   g02802(.A1(new_n5317_), .A2(new_n5243_), .B(new_n5108_), .ZN(new_n5318_));
  INV_X1     g02803(.I(new_n5298_), .ZN(new_n5319_));
  OAI21_X1   g02804(.A1(new_n5319_), .A2(new_n5108_), .B(new_n5318_), .ZN(new_n5320_));
  MUX2_X1    g02805(.I0(new_n5320_), .I1(new_n5213_), .S(new_n2523_), .Z(new_n5321_));
  OR2_X2     g02806(.A1(new_n5321_), .A2(new_n5238_), .Z(new_n5322_));
  INV_X1     g02807(.I(pi0145), .ZN(new_n5323_));
  INV_X1     g02808(.I(pi0180), .ZN(new_n5324_));
  INV_X1     g02809(.I(pi0181), .ZN(new_n5325_));
  INV_X1     g02810(.I(pi0182), .ZN(new_n5326_));
  NOR4_X1    g02811(.A1(new_n5323_), .A2(new_n5324_), .A3(new_n5325_), .A4(new_n5326_), .ZN(new_n5327_));
  AOI21_X1   g02812(.A1(new_n2587_), .A2(new_n5327_), .B(new_n5302_), .ZN(new_n5328_));
  AOI21_X1   g02813(.A1(new_n5322_), .A2(new_n5327_), .B(new_n5328_), .ZN(new_n5329_));
  NOR4_X1    g02814(.A1(new_n5242_), .A2(new_n2632_), .A3(pi0095), .A4(pi0210), .ZN(new_n5330_));
  INV_X1     g02815(.I(new_n5330_), .ZN(new_n5331_));
  NAND2_X1   g02816(.A1(new_n5297_), .A2(new_n5331_), .ZN(new_n5332_));
  INV_X1     g02817(.I(new_n5332_), .ZN(new_n5333_));
  NOR2_X1    g02818(.A1(new_n5333_), .A2(new_n5108_), .ZN(new_n5334_));
  OAI21_X1   g02819(.A1(new_n5317_), .A2(new_n5330_), .B(new_n5108_), .ZN(new_n5335_));
  INV_X1     g02820(.I(new_n5335_), .ZN(new_n5336_));
  NOR2_X1    g02821(.A1(new_n5334_), .A2(new_n5336_), .ZN(new_n5337_));
  INV_X1     g02822(.I(pi0160), .ZN(new_n5338_));
  INV_X1     g02823(.I(pi0197), .ZN(new_n5339_));
  INV_X1     g02824(.I(pi0158), .ZN(new_n5340_));
  INV_X1     g02825(.I(pi0159), .ZN(new_n5341_));
  NOR2_X1    g02826(.A1(new_n5340_), .A2(new_n5341_), .ZN(new_n5342_));
  INV_X1     g02827(.I(new_n5342_), .ZN(new_n5343_));
  NOR3_X1    g02828(.A1(new_n5343_), .A2(new_n5338_), .A3(new_n5339_), .ZN(new_n5344_));
  OAI21_X1   g02829(.A1(new_n5337_), .A2(new_n5219_), .B(new_n5344_), .ZN(new_n5345_));
  INV_X1     g02830(.I(new_n5344_), .ZN(new_n5346_));
  NAND2_X1   g02831(.A1(new_n5332_), .A2(new_n5220_), .ZN(new_n5347_));
  NAND2_X1   g02832(.A1(new_n5347_), .A2(new_n5346_), .ZN(new_n5348_));
  OAI21_X1   g02833(.A1(new_n5219_), .A2(new_n5215_), .B(pi0299), .ZN(new_n5349_));
  NOR2_X1    g02834(.A1(pi0228), .A2(pi0232), .ZN(new_n5350_));
  NAND4_X1   g02835(.A1(new_n5345_), .A2(new_n5348_), .A3(new_n5349_), .A4(new_n5350_), .ZN(new_n5351_));
  NAND2_X1   g02836(.A1(new_n5349_), .A2(new_n2523_), .ZN(new_n5352_));
  NOR2_X1    g02837(.A1(new_n5347_), .A2(new_n5352_), .ZN(new_n5353_));
  NOR2_X1    g02838(.A1(new_n5353_), .A2(pi0232), .ZN(new_n5354_));
  OAI22_X1   g02839(.A1(new_n5329_), .A2(new_n5351_), .B1(new_n5302_), .B2(new_n5354_), .ZN(new_n5355_));
  NOR2_X1    g02840(.A1(new_n2550_), .A2(pi0215), .ZN(new_n5356_));
  INV_X1     g02841(.I(new_n5356_), .ZN(new_n5357_));
  NOR2_X1    g02842(.A1(new_n2491_), .A2(pi0287), .ZN(new_n5358_));
  INV_X1     g02843(.I(new_n5358_), .ZN(new_n5359_));
  NOR2_X1    g02844(.A1(new_n5359_), .A2(new_n5123_), .ZN(new_n5360_));
  INV_X1     g02845(.I(new_n5360_), .ZN(new_n5361_));
  NOR2_X1    g02846(.A1(new_n5361_), .A2(new_n5118_), .ZN(new_n5362_));
  NOR2_X1    g02847(.A1(new_n2920_), .A2(pi0829), .ZN(new_n5363_));
  NOR2_X1    g02848(.A1(new_n5363_), .A2(new_n2918_), .ZN(new_n5364_));
  INV_X1     g02849(.I(new_n5364_), .ZN(new_n5365_));
  INV_X1     g02850(.I(pi0824), .ZN(new_n5366_));
  NOR2_X1    g02851(.A1(new_n5366_), .A2(new_n2924_), .ZN(new_n5367_));
  INV_X1     g02852(.I(new_n5367_), .ZN(new_n5368_));
  NOR2_X1    g02853(.A1(new_n5368_), .A2(new_n2955_), .ZN(new_n5369_));
  NAND3_X1   g02854(.A1(new_n5362_), .A2(new_n5365_), .A3(new_n5369_), .ZN(new_n5370_));
  INV_X1     g02855(.I(new_n5370_), .ZN(new_n5371_));
  NOR2_X1    g02856(.A1(new_n5371_), .A2(pi0216), .ZN(new_n5372_));
  MUX2_X1    g02857(.I0(new_n5372_), .I1(pi0030), .S(new_n2523_), .Z(new_n5373_));
  AND2_X2    g02858(.A1(new_n5373_), .A2(new_n5357_), .Z(new_n5374_));
  NAND2_X1   g02859(.A1(pi0030), .A2(pi0228), .ZN(new_n5375_));
  OAI21_X1   g02860(.A1(new_n5227_), .A2(new_n5375_), .B(new_n2587_), .ZN(new_n5376_));
  NAND2_X1   g02861(.A1(new_n5220_), .A2(new_n2587_), .ZN(new_n5377_));
  AOI21_X1   g02862(.A1(new_n5376_), .A2(pi0039), .B(new_n5377_), .ZN(new_n5378_));
  OAI21_X1   g02863(.A1(new_n5374_), .A2(new_n5214_), .B(new_n5378_), .ZN(new_n5379_));
  AOI21_X1   g02864(.A1(new_n5379_), .A2(new_n3172_), .B(pi0039), .ZN(new_n5380_));
  AOI21_X1   g02865(.A1(new_n5110_), .A2(new_n2491_), .B(new_n5217_), .ZN(new_n5381_));
  NAND2_X1   g02866(.A1(new_n5381_), .A2(pi0252), .ZN(new_n5382_));
  INV_X1     g02867(.I(new_n5161_), .ZN(new_n5383_));
  NOR4_X1    g02868(.A1(new_n5177_), .A2(new_n5178_), .A3(new_n2491_), .A4(new_n5186_), .ZN(new_n5384_));
  INV_X1     g02869(.I(new_n5384_), .ZN(new_n5385_));
  AOI21_X1   g02870(.A1(new_n5217_), .A2(new_n5109_), .B(new_n5385_), .ZN(new_n5386_));
  NAND3_X1   g02871(.A1(new_n5382_), .A2(pi0252), .A3(new_n5383_), .ZN(new_n5387_));
  NAND3_X1   g02872(.A1(new_n5382_), .A2(pi0252), .A3(new_n5383_), .ZN(new_n5388_));
  INV_X1     g02873(.I(new_n5386_), .ZN(new_n5389_));
  NOR2_X1    g02874(.A1(new_n5389_), .A2(new_n5383_), .ZN(new_n5390_));
  NAND2_X1   g02875(.A1(new_n5388_), .A2(new_n5390_), .ZN(new_n5391_));
  NAND2_X1   g02876(.A1(new_n5238_), .A2(new_n5214_), .ZN(new_n5392_));
  OAI21_X1   g02877(.A1(new_n5109_), .A2(pi0907), .B(new_n2523_), .ZN(new_n5393_));
  INV_X1     g02878(.I(pi0602), .ZN(new_n5394_));
  NAND2_X1   g02879(.A1(new_n5108_), .A2(new_n5394_), .ZN(new_n5395_));
  NAND4_X1   g02880(.A1(new_n5395_), .A2(new_n2545_), .A3(new_n2523_), .A4(new_n2587_), .ZN(new_n5396_));
  NOR2_X1    g02881(.A1(new_n3025_), .A2(new_n5396_), .ZN(new_n5397_));
  NAND4_X1   g02882(.A1(new_n5392_), .A2(new_n5349_), .A3(new_n5393_), .A4(new_n5397_), .ZN(new_n5398_));
  AOI21_X1   g02883(.A1(new_n5389_), .A2(new_n2577_), .B(new_n5398_), .ZN(new_n5399_));
  AND4_X2    g02884(.A1(new_n5382_), .A2(new_n5391_), .A3(new_n5387_), .A4(new_n5399_), .Z(new_n5400_));
  NOR2_X1    g02885(.A1(new_n2544_), .A2(pi0100), .ZN(new_n5401_));
  NAND2_X1   g02886(.A1(new_n5229_), .A2(new_n5401_), .ZN(new_n5402_));
  OAI21_X1   g02887(.A1(new_n5400_), .A2(new_n5402_), .B(new_n3177_), .ZN(new_n5403_));
  AOI21_X1   g02888(.A1(new_n5232_), .A2(new_n5215_), .B(new_n5228_), .ZN(new_n5404_));
  AOI21_X1   g02889(.A1(new_n5404_), .A2(new_n3172_), .B(pi0100), .ZN(new_n5405_));
  NAND2_X1   g02890(.A1(new_n5403_), .A2(new_n5405_), .ZN(new_n5406_));
  AOI21_X1   g02891(.A1(new_n5355_), .A2(new_n5380_), .B(new_n5406_), .ZN(new_n5407_));
  INV_X1     g02892(.I(new_n5229_), .ZN(new_n5408_));
  MUX2_X1    g02893(.I0(new_n5234_), .I1(new_n5408_), .S(new_n2628_), .Z(new_n5409_));
  INV_X1     g02894(.I(new_n5193_), .ZN(new_n5410_));
  NOR2_X1    g02895(.A1(new_n5410_), .A2(pi0075), .ZN(new_n5411_));
  OAI21_X1   g02896(.A1(new_n5408_), .A2(new_n3177_), .B(new_n5411_), .ZN(new_n5412_));
  AOI21_X1   g02897(.A1(new_n5235_), .A2(pi0075), .B(new_n5412_), .ZN(new_n5413_));
  OAI21_X1   g02898(.A1(pi0092), .A2(new_n5409_), .B(new_n5413_), .ZN(new_n5414_));
  NOR4_X1    g02899(.A1(new_n5234_), .A2(pi0054), .A3(new_n3228_), .A4(new_n5229_), .ZN(new_n5415_));
  NOR2_X1    g02900(.A1(new_n5415_), .A2(pi0074), .ZN(new_n5416_));
  OAI21_X1   g02901(.A1(new_n5407_), .A2(new_n5414_), .B(new_n5416_), .ZN(new_n5417_));
  NOR2_X1    g02902(.A1(new_n2533_), .A2(pi0055), .ZN(new_n5418_));
  NAND3_X1   g02903(.A1(new_n5216_), .A2(new_n5220_), .A3(new_n5418_), .ZN(new_n5419_));
  AOI21_X1   g02904(.A1(new_n5417_), .A2(new_n5237_), .B(new_n5419_), .ZN(new_n5420_));
  OAI21_X1   g02905(.A1(new_n5222_), .A2(pi0228), .B(new_n5205_), .ZN(new_n5421_));
  NOR2_X1    g02906(.A1(new_n5215_), .A2(new_n2533_), .ZN(new_n5422_));
  NAND2_X1   g02907(.A1(new_n5220_), .A2(new_n5422_), .ZN(new_n5423_));
  AOI21_X1   g02908(.A1(new_n5423_), .A2(new_n5205_), .B(pi0057), .ZN(new_n5424_));
  OAI21_X1   g02909(.A1(new_n5221_), .A2(new_n5421_), .B(new_n5424_), .ZN(new_n5425_));
  OAI22_X1   g02910(.A1(new_n5420_), .A2(new_n5425_), .B1(new_n5221_), .B2(new_n5225_), .ZN(po0171));
  INV_X1     g02911(.I(new_n5106_), .ZN(new_n5427_));
  NOR2_X1    g02912(.A1(new_n5427_), .A2(new_n5108_), .ZN(new_n5428_));
  AOI21_X1   g02913(.A1(pi0947), .A2(new_n5108_), .B(new_n5428_), .ZN(new_n5429_));
  INV_X1     g02914(.I(new_n5429_), .ZN(new_n5430_));
  NAND2_X1   g02915(.A1(new_n5216_), .A2(new_n5430_), .ZN(new_n5431_));
  AOI21_X1   g02916(.A1(pi0587), .A2(new_n5108_), .B(new_n5428_), .ZN(new_n5432_));
  MUX2_X1    g02917(.I0(new_n5432_), .I1(new_n5429_), .S(pi0299), .Z(new_n5433_));
  NOR2_X1    g02918(.A1(new_n5433_), .A2(new_n5215_), .ZN(new_n5434_));
  NOR2_X1    g02919(.A1(new_n5434_), .A2(new_n5226_), .ZN(new_n5435_));
  NOR2_X1    g02920(.A1(new_n5232_), .A2(new_n5433_), .ZN(new_n5436_));
  AOI22_X1   g02921(.A1(new_n5436_), .A2(new_n3207_), .B1(new_n2629_), .B2(new_n5434_), .ZN(new_n5437_));
  INV_X1     g02922(.I(new_n5437_), .ZN(new_n5438_));
  AOI21_X1   g02923(.A1(new_n5438_), .A2(new_n5226_), .B(new_n5435_), .ZN(new_n5439_));
  OAI21_X1   g02924(.A1(new_n5439_), .A2(pi0074), .B(new_n3227_), .ZN(new_n5440_));
  INV_X1     g02925(.I(new_n5321_), .ZN(new_n5441_));
  INV_X1     g02926(.I(new_n5327_), .ZN(new_n5442_));
  INV_X1     g02927(.I(new_n5301_), .ZN(new_n5443_));
  NOR2_X1    g02928(.A1(new_n5443_), .A2(new_n5432_), .ZN(new_n5444_));
  NAND4_X1   g02929(.A1(new_n5441_), .A2(new_n5442_), .A3(new_n5432_), .A4(new_n5444_), .ZN(new_n5445_));
  INV_X1     g02930(.I(new_n5432_), .ZN(new_n5446_));
  OAI22_X1   g02931(.A1(new_n5321_), .A2(new_n5446_), .B1(new_n5444_), .B2(new_n5327_), .ZN(new_n5447_));
  OAI21_X1   g02932(.A1(new_n5334_), .A2(new_n5336_), .B(new_n5430_), .ZN(new_n5448_));
  NOR2_X1    g02933(.A1(new_n5333_), .A2(new_n5429_), .ZN(new_n5449_));
  INV_X1     g02934(.I(new_n5449_), .ZN(new_n5450_));
  NAND2_X1   g02935(.A1(new_n5450_), .A2(new_n5346_), .ZN(new_n5451_));
  AOI21_X1   g02936(.A1(new_n5430_), .A2(new_n5214_), .B(new_n2587_), .ZN(new_n5452_));
  INV_X1     g02937(.I(new_n5452_), .ZN(new_n5453_));
  NAND4_X1   g02938(.A1(new_n5451_), .A2(new_n2587_), .A3(new_n5350_), .A4(new_n5453_), .ZN(new_n5454_));
  AOI21_X1   g02939(.A1(new_n5344_), .A2(new_n5448_), .B(new_n5454_), .ZN(new_n5455_));
  NAND3_X1   g02940(.A1(new_n5455_), .A2(new_n5445_), .A3(new_n5447_), .ZN(new_n5456_));
  NOR3_X1    g02941(.A1(new_n5450_), .A2(pi0228), .A3(new_n5452_), .ZN(new_n5457_));
  OAI22_X1   g02942(.A1(new_n5444_), .A2(pi0299), .B1(new_n5457_), .B2(pi0232), .ZN(new_n5458_));
  NAND2_X1   g02943(.A1(new_n5456_), .A2(new_n5458_), .ZN(new_n5459_));
  INV_X1     g02944(.I(pi0142), .ZN(new_n5460_));
  NOR2_X1    g02945(.A1(new_n5106_), .A2(new_n5108_), .ZN(new_n5461_));
  NOR2_X1    g02946(.A1(new_n5385_), .A2(new_n5461_), .ZN(new_n5462_));
  INV_X1     g02947(.I(new_n5462_), .ZN(new_n5463_));
  AOI21_X1   g02948(.A1(new_n5110_), .A2(new_n2491_), .B(new_n5427_), .ZN(new_n5464_));
  NAND2_X1   g02949(.A1(new_n5464_), .A2(pi0252), .ZN(new_n5465_));
  MUX2_X1    g02950(.I0(new_n5465_), .I1(new_n5463_), .S(new_n5460_), .Z(new_n5466_));
  OAI21_X1   g02951(.A1(new_n5428_), .A2(pi0587), .B(new_n2523_), .ZN(new_n5467_));
  INV_X1     g02952(.I(pi0587), .ZN(new_n5468_));
  AOI22_X1   g02953(.A1(new_n5446_), .A2(new_n5214_), .B1(new_n2523_), .B2(new_n2605_), .ZN(new_n5470_));
  OAI21_X1   g02954(.A1(new_n5466_), .A2(new_n5467_), .B(new_n5470_), .ZN(new_n5471_));
  OAI21_X1   g02955(.A1(new_n5428_), .A2(pi0947), .B(new_n3025_), .ZN(new_n5472_));
  INV_X1     g02956(.I(pi0947), .ZN(new_n5473_));
  AOI21_X1   g02957(.A1(new_n5473_), .A2(new_n5108_), .B(new_n3025_), .ZN(new_n5474_));
  AOI21_X1   g02958(.A1(new_n5462_), .A2(new_n5474_), .B(pi0228), .ZN(new_n5475_));
  OAI21_X1   g02959(.A1(new_n5465_), .A2(new_n5472_), .B(new_n5475_), .ZN(new_n5476_));
  NOR2_X1    g02960(.A1(new_n5453_), .A2(new_n2544_), .ZN(new_n5477_));
  AOI21_X1   g02961(.A1(new_n5476_), .A2(new_n5477_), .B(pi0299), .ZN(new_n5478_));
  NAND2_X1   g02962(.A1(new_n5434_), .A2(new_n5401_), .ZN(new_n5479_));
  AOI21_X1   g02963(.A1(new_n5471_), .A2(new_n5478_), .B(new_n5479_), .ZN(new_n5480_));
  NAND3_X1   g02964(.A1(new_n5446_), .A2(pi0030), .A3(pi0228), .ZN(new_n5481_));
  AOI21_X1   g02965(.A1(new_n5481_), .A2(new_n2587_), .B(new_n3154_), .ZN(new_n5482_));
  NOR2_X1    g02966(.A1(new_n5357_), .A2(new_n2587_), .ZN(new_n5483_));
  NOR4_X1    g02967(.A1(new_n5482_), .A2(new_n5429_), .A3(new_n5452_), .A4(new_n5483_), .ZN(new_n5484_));
  INV_X1     g02968(.I(new_n5434_), .ZN(new_n5485_));
  INV_X1     g02969(.I(new_n5436_), .ZN(new_n5486_));
  NAND4_X1   g02970(.A1(new_n5486_), .A2(new_n3172_), .A3(new_n3173_), .A4(new_n5485_), .ZN(new_n5487_));
  AOI21_X1   g02971(.A1(new_n5374_), .A2(new_n5484_), .B(new_n5487_), .ZN(new_n5488_));
  OAI21_X1   g02972(.A1(pi0087), .A2(new_n5480_), .B(new_n5488_), .ZN(new_n5489_));
  AOI21_X1   g02973(.A1(new_n5459_), .A2(new_n3154_), .B(new_n5489_), .ZN(new_n5490_));
  MUX2_X1    g02974(.I0(new_n5437_), .I1(new_n5485_), .S(new_n2628_), .Z(new_n5491_));
  OAI21_X1   g02975(.A1(new_n5485_), .A2(new_n3177_), .B(new_n5411_), .ZN(new_n5492_));
  AOI21_X1   g02976(.A1(new_n5438_), .A2(pi0075), .B(new_n5492_), .ZN(new_n5493_));
  OAI21_X1   g02977(.A1(new_n5491_), .A2(pi0092), .B(new_n5493_), .ZN(new_n5494_));
  NOR4_X1    g02978(.A1(new_n5437_), .A2(pi0054), .A3(new_n3228_), .A4(new_n5434_), .ZN(new_n5495_));
  NOR2_X1    g02979(.A1(new_n5495_), .A2(pi0074), .ZN(new_n5496_));
  OAI21_X1   g02980(.A1(new_n5490_), .A2(new_n5494_), .B(new_n5496_), .ZN(new_n5497_));
  NAND3_X1   g02981(.A1(new_n5216_), .A2(new_n5418_), .A3(new_n5430_), .ZN(new_n5498_));
  AOI21_X1   g02982(.A1(new_n5497_), .A2(new_n5440_), .B(new_n5498_), .ZN(new_n5499_));
  NAND2_X1   g02983(.A1(new_n5430_), .A2(new_n5422_), .ZN(new_n5500_));
  AOI21_X1   g02984(.A1(new_n5500_), .A2(new_n5205_), .B(pi0057), .ZN(new_n5501_));
  OAI21_X1   g02985(.A1(new_n5431_), .A2(new_n5421_), .B(new_n5501_), .ZN(new_n5502_));
  OAI22_X1   g02986(.A1(new_n5499_), .A2(new_n5502_), .B1(new_n5225_), .B2(new_n5431_), .ZN(po0172));
  INV_X1     g02987(.I(pi0970), .ZN(new_n5504_));
  NAND2_X1   g02988(.A1(new_n5110_), .A2(new_n2523_), .ZN(new_n5505_));
  NOR2_X1    g02989(.A1(new_n5505_), .A2(new_n5504_), .ZN(new_n5506_));
  NAND2_X1   g02990(.A1(new_n5506_), .A2(new_n3233_), .ZN(new_n5507_));
  NOR2_X1    g02991(.A1(new_n5507_), .A2(new_n5223_), .ZN(new_n5508_));
  NOR3_X1    g02992(.A1(new_n5109_), .A2(new_n5213_), .A3(new_n2523_), .ZN(new_n5509_));
  INV_X1     g02993(.I(new_n5509_), .ZN(new_n5510_));
  NOR2_X1    g02994(.A1(new_n5510_), .A2(new_n5504_), .ZN(new_n5511_));
  INV_X1     g02995(.I(new_n5511_), .ZN(new_n5512_));
  NAND2_X1   g02996(.A1(new_n5512_), .A2(pi0057), .ZN(new_n5513_));
  INV_X1     g02997(.I(pi0967), .ZN(new_n5514_));
  NAND2_X1   g02998(.A1(new_n3162_), .A2(pi0228), .ZN(new_n5515_));
  AOI21_X1   g02999(.A1(new_n5515_), .A2(new_n5215_), .B(new_n5109_), .ZN(new_n5516_));
  INV_X1     g03000(.I(new_n5516_), .ZN(new_n5517_));
  OAI21_X1   g03001(.A1(new_n5517_), .A2(new_n5514_), .B(new_n2587_), .ZN(new_n5518_));
  NOR2_X1    g03002(.A1(new_n5511_), .A2(new_n2587_), .ZN(new_n5519_));
  INV_X1     g03003(.I(new_n5519_), .ZN(new_n5520_));
  NAND2_X1   g03004(.A1(new_n5506_), .A2(new_n5520_), .ZN(new_n5521_));
  NAND3_X1   g03005(.A1(new_n5518_), .A2(new_n5521_), .A3(new_n3154_), .ZN(new_n5522_));
  MUX2_X1    g03006(.I0(new_n5514_), .I1(new_n5504_), .S(pi0299), .Z(new_n5523_));
  NOR2_X1    g03007(.A1(new_n5510_), .A2(new_n5523_), .ZN(new_n5524_));
  NOR2_X1    g03008(.A1(new_n3154_), .A2(pi0038), .ZN(new_n5525_));
  NAND2_X1   g03009(.A1(new_n5524_), .A2(new_n5525_), .ZN(new_n5526_));
  NOR4_X1    g03010(.A1(new_n5109_), .A2(new_n5213_), .A3(pi0039), .A4(pi0228), .ZN(new_n5527_));
  NAND2_X1   g03011(.A1(new_n2587_), .A2(pi0228), .ZN(new_n5528_));
  NOR2_X1    g03012(.A1(new_n5372_), .A2(new_n5357_), .ZN(new_n5529_));
  AOI21_X1   g03013(.A1(new_n5529_), .A2(new_n5108_), .B(pi0228), .ZN(new_n5530_));
  OR2_X2     g03014(.A1(new_n5530_), .A2(new_n2587_), .Z(new_n5531_));
  OAI22_X1   g03015(.A1(new_n5531_), .A2(new_n5504_), .B1(new_n5514_), .B2(new_n5528_), .ZN(new_n5532_));
  AOI21_X1   g03016(.A1(new_n5532_), .A2(new_n5527_), .B(pi0038), .ZN(new_n5533_));
  NOR2_X1    g03017(.A1(new_n5443_), .A2(new_n5109_), .ZN(new_n5534_));
  AOI21_X1   g03018(.A1(new_n5534_), .A2(pi0967), .B(pi0299), .ZN(new_n5535_));
  NOR2_X1    g03019(.A1(new_n5109_), .A2(pi0228), .ZN(new_n5536_));
  NAND2_X1   g03020(.A1(new_n5332_), .A2(new_n5536_), .ZN(new_n5537_));
  NOR3_X1    g03021(.A1(new_n5537_), .A2(new_n5504_), .A3(new_n5519_), .ZN(new_n5538_));
  OR3_X2     g03022(.A1(new_n5535_), .A2(pi0232), .A3(new_n5538_), .Z(new_n5539_));
  NAND2_X1   g03023(.A1(new_n5339_), .A2(pi0160), .ZN(new_n5540_));
  MUX2_X1    g03024(.I0(new_n5335_), .I1(new_n5332_), .S(new_n5540_), .Z(new_n5541_));
  INV_X1     g03025(.I(new_n5541_), .ZN(new_n5542_));
  AOI21_X1   g03026(.A1(new_n5542_), .A2(new_n5536_), .B(new_n5509_), .ZN(new_n5543_));
  NAND2_X1   g03027(.A1(new_n5342_), .A2(new_n2587_), .ZN(new_n5544_));
  NOR2_X1    g03028(.A1(new_n5538_), .A2(new_n5544_), .ZN(new_n5545_));
  OAI21_X1   g03029(.A1(new_n5543_), .A2(new_n5504_), .B(new_n5545_), .ZN(new_n5546_));
  NOR2_X1    g03030(.A1(new_n5318_), .A2(pi0228), .ZN(new_n5547_));
  OAI21_X1   g03031(.A1(new_n5319_), .A2(new_n5327_), .B(new_n5510_), .ZN(new_n5548_));
  OAI22_X1   g03032(.A1(new_n5534_), .A2(new_n5327_), .B1(new_n5547_), .B2(new_n5548_), .ZN(new_n5549_));
  OAI21_X1   g03033(.A1(new_n5549_), .A2(new_n5514_), .B(new_n2587_), .ZN(new_n5550_));
  NAND3_X1   g03034(.A1(new_n5550_), .A2(pi0232), .A3(new_n5546_), .ZN(new_n5551_));
  AOI21_X1   g03035(.A1(new_n5551_), .A2(new_n5539_), .B(pi0039), .ZN(new_n5552_));
  OAI22_X1   g03036(.A1(new_n5552_), .A2(new_n5533_), .B1(new_n5522_), .B2(new_n5526_), .ZN(new_n5553_));
  NOR2_X1    g03037(.A1(new_n5111_), .A2(new_n3181_), .ZN(new_n5554_));
  NOR2_X1    g03038(.A1(new_n5385_), .A2(new_n5109_), .ZN(new_n5555_));
  INV_X1     g03039(.I(new_n5555_), .ZN(new_n5556_));
  NOR3_X1    g03040(.A1(new_n5554_), .A2(new_n5556_), .A3(new_n3025_), .ZN(new_n5557_));
  INV_X1     g03041(.I(new_n5554_), .ZN(new_n5558_));
  AOI21_X1   g03042(.A1(new_n2577_), .A2(new_n5556_), .B(new_n5558_), .ZN(new_n5559_));
  OAI21_X1   g03043(.A1(new_n5559_), .A2(new_n5557_), .B(new_n2523_), .ZN(new_n5560_));
  NOR2_X1    g03044(.A1(new_n5109_), .A2(new_n5213_), .ZN(new_n5561_));
  NOR2_X1    g03045(.A1(new_n5556_), .A2(new_n5383_), .ZN(new_n5562_));
  NOR2_X1    g03046(.A1(new_n5554_), .A2(new_n5383_), .ZN(new_n5563_));
  NOR4_X1    g03047(.A1(new_n5563_), .A2(new_n5562_), .A3(pi0228), .A4(new_n5561_), .ZN(new_n5564_));
  OAI21_X1   g03048(.A1(new_n5564_), .A2(new_n5514_), .B(new_n2587_), .ZN(new_n5565_));
  NAND4_X1   g03049(.A1(new_n5565_), .A2(pi0970), .A3(new_n2545_), .A4(new_n5520_), .ZN(new_n5566_));
  INV_X1     g03050(.I(new_n5401_), .ZN(new_n5567_));
  INV_X1     g03051(.I(new_n5524_), .ZN(new_n5568_));
  NOR2_X1    g03052(.A1(new_n5568_), .A2(new_n5567_), .ZN(new_n5569_));
  OAI21_X1   g03053(.A1(new_n5566_), .A2(new_n5560_), .B(new_n5569_), .ZN(new_n5570_));
  AOI21_X1   g03054(.A1(new_n5570_), .A2(new_n3177_), .B(pi0100), .ZN(new_n5571_));
  AOI22_X1   g03055(.A1(new_n5522_), .A2(new_n3207_), .B1(new_n2629_), .B2(new_n5524_), .ZN(new_n5572_));
  MUX2_X1    g03056(.I0(new_n5572_), .I1(new_n5568_), .S(new_n2628_), .Z(new_n5573_));
  INV_X1     g03057(.I(new_n5572_), .ZN(new_n5574_));
  OAI21_X1   g03058(.A1(new_n5568_), .A2(new_n3177_), .B(new_n5411_), .ZN(new_n5575_));
  AOI21_X1   g03059(.A1(new_n5574_), .A2(pi0075), .B(new_n5575_), .ZN(new_n5576_));
  OAI21_X1   g03060(.A1(pi0092), .A2(new_n5573_), .B(new_n5576_), .ZN(new_n5577_));
  AOI21_X1   g03061(.A1(new_n5553_), .A2(new_n5571_), .B(new_n5577_), .ZN(new_n5578_));
  NOR2_X1    g03062(.A1(new_n5574_), .A2(new_n3228_), .ZN(new_n5579_));
  OAI21_X1   g03063(.A1(new_n5568_), .A2(new_n3209_), .B(pi0054), .ZN(new_n5580_));
  OAI21_X1   g03064(.A1(new_n5579_), .A2(new_n5580_), .B(new_n3202_), .ZN(new_n5581_));
  INV_X1     g03065(.I(new_n5226_), .ZN(new_n5582_));
  NOR2_X1    g03066(.A1(new_n5582_), .A2(pi0074), .ZN(new_n5583_));
  AOI21_X1   g03067(.A1(new_n5574_), .A2(new_n5583_), .B(pi0055), .ZN(new_n5584_));
  OAI21_X1   g03068(.A1(new_n5578_), .A2(new_n5581_), .B(new_n5584_), .ZN(new_n5585_));
  INV_X1     g03069(.I(new_n5418_), .ZN(new_n5586_));
  AOI21_X1   g03070(.A1(new_n5507_), .A2(new_n5512_), .B(new_n5586_), .ZN(new_n5587_));
  NAND2_X1   g03071(.A1(new_n5512_), .A2(new_n5224_), .ZN(new_n5588_));
  AOI21_X1   g03072(.A1(new_n5511_), .A2(new_n3503_), .B(pi0059), .ZN(new_n5589_));
  OAI21_X1   g03073(.A1(new_n5507_), .A2(new_n5588_), .B(new_n5589_), .ZN(new_n5590_));
  AOI21_X1   g03074(.A1(new_n5585_), .A2(new_n5587_), .B(new_n5590_), .ZN(new_n5591_));
  OAI22_X1   g03075(.A1(new_n5591_), .A2(pi0057), .B1(new_n5508_), .B2(new_n5513_), .ZN(po0173));
  INV_X1     g03076(.I(pi0972), .ZN(new_n5593_));
  NOR2_X1    g03077(.A1(new_n5505_), .A2(new_n5593_), .ZN(new_n5594_));
  NAND2_X1   g03078(.A1(new_n5594_), .A2(new_n3233_), .ZN(new_n5595_));
  NOR2_X1    g03079(.A1(new_n5595_), .A2(new_n5223_), .ZN(new_n5596_));
  NOR2_X1    g03080(.A1(new_n5510_), .A2(new_n5593_), .ZN(new_n5597_));
  INV_X1     g03081(.I(new_n5597_), .ZN(new_n5598_));
  NAND2_X1   g03082(.A1(new_n5598_), .A2(pi0057), .ZN(new_n5599_));
  INV_X1     g03083(.I(pi0961), .ZN(new_n5600_));
  OAI21_X1   g03084(.A1(new_n5517_), .A2(new_n5600_), .B(new_n2587_), .ZN(new_n5601_));
  NOR2_X1    g03085(.A1(new_n5597_), .A2(new_n2587_), .ZN(new_n5602_));
  INV_X1     g03086(.I(new_n5602_), .ZN(new_n5603_));
  NAND2_X1   g03087(.A1(new_n5594_), .A2(new_n5603_), .ZN(new_n5604_));
  NAND3_X1   g03088(.A1(new_n5601_), .A2(new_n5604_), .A3(new_n3154_), .ZN(new_n5605_));
  MUX2_X1    g03089(.I0(new_n5600_), .I1(new_n5593_), .S(pi0299), .Z(new_n5606_));
  NOR2_X1    g03090(.A1(new_n5510_), .A2(new_n5606_), .ZN(new_n5607_));
  NAND2_X1   g03091(.A1(new_n5607_), .A2(new_n5525_), .ZN(new_n5608_));
  OAI22_X1   g03092(.A1(new_n5531_), .A2(new_n5593_), .B1(new_n5600_), .B2(new_n5528_), .ZN(new_n5609_));
  AOI21_X1   g03093(.A1(new_n5609_), .A2(new_n5527_), .B(pi0038), .ZN(new_n5610_));
  AOI21_X1   g03094(.A1(new_n5534_), .A2(pi0961), .B(pi0299), .ZN(new_n5611_));
  NOR3_X1    g03095(.A1(new_n5537_), .A2(new_n5593_), .A3(new_n5602_), .ZN(new_n5612_));
  OR3_X2     g03096(.A1(new_n5611_), .A2(pi0232), .A3(new_n5612_), .Z(new_n5613_));
  NOR2_X1    g03097(.A1(new_n5612_), .A2(new_n5544_), .ZN(new_n5614_));
  OAI21_X1   g03098(.A1(new_n5543_), .A2(new_n5593_), .B(new_n5614_), .ZN(new_n5615_));
  OAI21_X1   g03099(.A1(new_n5549_), .A2(new_n5600_), .B(new_n2587_), .ZN(new_n5616_));
  NAND3_X1   g03100(.A1(new_n5616_), .A2(pi0232), .A3(new_n5615_), .ZN(new_n5617_));
  AOI21_X1   g03101(.A1(new_n5617_), .A2(new_n5613_), .B(pi0039), .ZN(new_n5618_));
  OAI22_X1   g03102(.A1(new_n5618_), .A2(new_n5610_), .B1(new_n5605_), .B2(new_n5608_), .ZN(new_n5619_));
  OAI21_X1   g03103(.A1(new_n5564_), .A2(new_n5600_), .B(new_n2587_), .ZN(new_n5620_));
  NAND4_X1   g03104(.A1(new_n5620_), .A2(pi0972), .A3(new_n2545_), .A4(new_n5603_), .ZN(new_n5621_));
  INV_X1     g03105(.I(new_n5607_), .ZN(new_n5622_));
  NOR2_X1    g03106(.A1(new_n5622_), .A2(new_n5567_), .ZN(new_n5623_));
  OAI21_X1   g03107(.A1(new_n5621_), .A2(new_n5560_), .B(new_n5623_), .ZN(new_n5624_));
  AOI21_X1   g03108(.A1(new_n5624_), .A2(new_n3177_), .B(pi0100), .ZN(new_n5625_));
  AOI22_X1   g03109(.A1(new_n5605_), .A2(new_n3207_), .B1(new_n2629_), .B2(new_n5607_), .ZN(new_n5626_));
  MUX2_X1    g03110(.I0(new_n5626_), .I1(new_n5622_), .S(new_n2628_), .Z(new_n5627_));
  INV_X1     g03111(.I(new_n5626_), .ZN(new_n5628_));
  OAI21_X1   g03112(.A1(new_n5622_), .A2(new_n3177_), .B(new_n5411_), .ZN(new_n5629_));
  AOI21_X1   g03113(.A1(new_n5628_), .A2(pi0075), .B(new_n5629_), .ZN(new_n5630_));
  OAI21_X1   g03114(.A1(pi0092), .A2(new_n5627_), .B(new_n5630_), .ZN(new_n5631_));
  AOI21_X1   g03115(.A1(new_n5619_), .A2(new_n5625_), .B(new_n5631_), .ZN(new_n5632_));
  NOR2_X1    g03116(.A1(new_n5628_), .A2(new_n3228_), .ZN(new_n5633_));
  OAI21_X1   g03117(.A1(new_n5622_), .A2(new_n3209_), .B(pi0054), .ZN(new_n5634_));
  OAI21_X1   g03118(.A1(new_n5633_), .A2(new_n5634_), .B(new_n3202_), .ZN(new_n5635_));
  NOR2_X1    g03119(.A1(new_n5582_), .A2(pi0074), .ZN(new_n5636_));
  AOI21_X1   g03120(.A1(new_n5628_), .A2(new_n5636_), .B(pi0055), .ZN(new_n5637_));
  OAI21_X1   g03121(.A1(new_n5632_), .A2(new_n5635_), .B(new_n5637_), .ZN(new_n5638_));
  AOI21_X1   g03122(.A1(new_n5595_), .A2(new_n5598_), .B(new_n5586_), .ZN(new_n5639_));
  NAND2_X1   g03123(.A1(new_n5598_), .A2(new_n5224_), .ZN(new_n5640_));
  AOI21_X1   g03124(.A1(new_n5597_), .A2(new_n3503_), .B(pi0059), .ZN(new_n5641_));
  OAI21_X1   g03125(.A1(new_n5595_), .A2(new_n5640_), .B(new_n5641_), .ZN(new_n5642_));
  AOI21_X1   g03126(.A1(new_n5638_), .A2(new_n5639_), .B(new_n5642_), .ZN(new_n5643_));
  OAI22_X1   g03127(.A1(new_n5643_), .A2(pi0057), .B1(new_n5596_), .B2(new_n5599_), .ZN(po0174));
  INV_X1     g03128(.I(pi0960), .ZN(new_n5645_));
  NOR2_X1    g03129(.A1(new_n5505_), .A2(new_n5645_), .ZN(new_n5646_));
  NAND2_X1   g03130(.A1(new_n5646_), .A2(new_n3233_), .ZN(new_n5647_));
  NOR2_X1    g03131(.A1(new_n5647_), .A2(new_n5223_), .ZN(new_n5648_));
  NOR2_X1    g03132(.A1(new_n5510_), .A2(new_n5645_), .ZN(new_n5649_));
  INV_X1     g03133(.I(new_n5649_), .ZN(new_n5650_));
  NAND2_X1   g03134(.A1(new_n5650_), .A2(pi0057), .ZN(new_n5651_));
  INV_X1     g03135(.I(pi0977), .ZN(new_n5652_));
  OAI21_X1   g03136(.A1(new_n5517_), .A2(new_n5652_), .B(new_n2587_), .ZN(new_n5653_));
  NOR2_X1    g03137(.A1(new_n5649_), .A2(new_n2587_), .ZN(new_n5654_));
  INV_X1     g03138(.I(new_n5654_), .ZN(new_n5655_));
  NAND2_X1   g03139(.A1(new_n5646_), .A2(new_n5655_), .ZN(new_n5656_));
  NAND3_X1   g03140(.A1(new_n5653_), .A2(new_n5656_), .A3(new_n3154_), .ZN(new_n5657_));
  MUX2_X1    g03141(.I0(new_n5652_), .I1(new_n5645_), .S(pi0299), .Z(new_n5658_));
  NOR2_X1    g03142(.A1(new_n5510_), .A2(new_n5658_), .ZN(new_n5659_));
  NAND2_X1   g03143(.A1(new_n5659_), .A2(new_n5525_), .ZN(new_n5660_));
  OAI22_X1   g03144(.A1(new_n5531_), .A2(new_n5645_), .B1(new_n5652_), .B2(new_n5528_), .ZN(new_n5661_));
  AOI21_X1   g03145(.A1(new_n5661_), .A2(new_n5527_), .B(pi0038), .ZN(new_n5662_));
  AOI21_X1   g03146(.A1(new_n5534_), .A2(pi0977), .B(pi0299), .ZN(new_n5663_));
  NOR3_X1    g03147(.A1(new_n5537_), .A2(new_n5645_), .A3(new_n5654_), .ZN(new_n5664_));
  OR3_X2     g03148(.A1(new_n5663_), .A2(pi0232), .A3(new_n5664_), .Z(new_n5665_));
  NOR2_X1    g03149(.A1(new_n5664_), .A2(new_n5544_), .ZN(new_n5666_));
  OAI21_X1   g03150(.A1(new_n5543_), .A2(new_n5645_), .B(new_n5666_), .ZN(new_n5667_));
  OAI21_X1   g03151(.A1(new_n5549_), .A2(new_n5652_), .B(new_n2587_), .ZN(new_n5668_));
  NAND3_X1   g03152(.A1(new_n5668_), .A2(pi0232), .A3(new_n5667_), .ZN(new_n5669_));
  AOI21_X1   g03153(.A1(new_n5669_), .A2(new_n5665_), .B(pi0039), .ZN(new_n5670_));
  OAI22_X1   g03154(.A1(new_n5670_), .A2(new_n5662_), .B1(new_n5657_), .B2(new_n5660_), .ZN(new_n5671_));
  OAI21_X1   g03155(.A1(new_n5564_), .A2(new_n5652_), .B(new_n2587_), .ZN(new_n5672_));
  NAND4_X1   g03156(.A1(new_n5672_), .A2(pi0960), .A3(new_n2545_), .A4(new_n5655_), .ZN(new_n5673_));
  INV_X1     g03157(.I(new_n5659_), .ZN(new_n5674_));
  NOR2_X1    g03158(.A1(new_n5674_), .A2(new_n5567_), .ZN(new_n5675_));
  OAI21_X1   g03159(.A1(new_n5673_), .A2(new_n5560_), .B(new_n5675_), .ZN(new_n5676_));
  AOI21_X1   g03160(.A1(new_n5676_), .A2(new_n3177_), .B(pi0100), .ZN(new_n5677_));
  AOI22_X1   g03161(.A1(new_n5657_), .A2(new_n3207_), .B1(new_n2629_), .B2(new_n5659_), .ZN(new_n5678_));
  MUX2_X1    g03162(.I0(new_n5678_), .I1(new_n5674_), .S(new_n2628_), .Z(new_n5679_));
  INV_X1     g03163(.I(new_n5678_), .ZN(new_n5680_));
  OAI21_X1   g03164(.A1(new_n5674_), .A2(new_n3177_), .B(new_n5411_), .ZN(new_n5681_));
  AOI21_X1   g03165(.A1(new_n5680_), .A2(pi0075), .B(new_n5681_), .ZN(new_n5682_));
  OAI21_X1   g03166(.A1(pi0092), .A2(new_n5679_), .B(new_n5682_), .ZN(new_n5683_));
  AOI21_X1   g03167(.A1(new_n5671_), .A2(new_n5677_), .B(new_n5683_), .ZN(new_n5684_));
  NOR2_X1    g03168(.A1(new_n5680_), .A2(new_n3228_), .ZN(new_n5685_));
  OAI21_X1   g03169(.A1(new_n5674_), .A2(new_n3209_), .B(pi0054), .ZN(new_n5686_));
  OAI21_X1   g03170(.A1(new_n5685_), .A2(new_n5686_), .B(new_n3202_), .ZN(new_n5687_));
  NOR2_X1    g03171(.A1(new_n5582_), .A2(pi0074), .ZN(new_n5688_));
  AOI21_X1   g03172(.A1(new_n5680_), .A2(new_n5688_), .B(pi0055), .ZN(new_n5689_));
  OAI21_X1   g03173(.A1(new_n5684_), .A2(new_n5687_), .B(new_n5689_), .ZN(new_n5690_));
  AOI21_X1   g03174(.A1(new_n5647_), .A2(new_n5650_), .B(new_n5586_), .ZN(new_n5691_));
  NAND2_X1   g03175(.A1(new_n5650_), .A2(new_n5224_), .ZN(new_n5692_));
  AOI21_X1   g03176(.A1(new_n5649_), .A2(new_n3503_), .B(pi0059), .ZN(new_n5693_));
  OAI21_X1   g03177(.A1(new_n5647_), .A2(new_n5692_), .B(new_n5693_), .ZN(new_n5694_));
  AOI21_X1   g03178(.A1(new_n5690_), .A2(new_n5691_), .B(new_n5694_), .ZN(new_n5695_));
  OAI22_X1   g03179(.A1(new_n5695_), .A2(pi0057), .B1(new_n5648_), .B2(new_n5651_), .ZN(po0175));
  INV_X1     g03180(.I(pi0963), .ZN(new_n5697_));
  NOR2_X1    g03181(.A1(new_n5505_), .A2(new_n5697_), .ZN(new_n5698_));
  NAND2_X1   g03182(.A1(new_n5698_), .A2(new_n3233_), .ZN(new_n5699_));
  NOR2_X1    g03183(.A1(new_n5699_), .A2(new_n5223_), .ZN(new_n5700_));
  NOR2_X1    g03184(.A1(new_n5510_), .A2(new_n5697_), .ZN(new_n5701_));
  INV_X1     g03185(.I(new_n5701_), .ZN(new_n5702_));
  NAND2_X1   g03186(.A1(new_n5702_), .A2(pi0057), .ZN(new_n5703_));
  INV_X1     g03187(.I(pi0969), .ZN(new_n5704_));
  OAI21_X1   g03188(.A1(new_n5517_), .A2(new_n5704_), .B(new_n2587_), .ZN(new_n5705_));
  NOR2_X1    g03189(.A1(new_n5701_), .A2(new_n2587_), .ZN(new_n5706_));
  INV_X1     g03190(.I(new_n5706_), .ZN(new_n5707_));
  NAND2_X1   g03191(.A1(new_n5698_), .A2(new_n5707_), .ZN(new_n5708_));
  NAND3_X1   g03192(.A1(new_n5705_), .A2(new_n5708_), .A3(new_n3154_), .ZN(new_n5709_));
  MUX2_X1    g03193(.I0(new_n5704_), .I1(new_n5697_), .S(pi0299), .Z(new_n5710_));
  NOR2_X1    g03194(.A1(new_n5510_), .A2(new_n5710_), .ZN(new_n5711_));
  NAND2_X1   g03195(.A1(new_n5711_), .A2(new_n5525_), .ZN(new_n5712_));
  OAI22_X1   g03196(.A1(new_n5531_), .A2(new_n5697_), .B1(new_n5704_), .B2(new_n5528_), .ZN(new_n5713_));
  AOI21_X1   g03197(.A1(new_n5713_), .A2(new_n5527_), .B(pi0038), .ZN(new_n5714_));
  AOI21_X1   g03198(.A1(new_n5534_), .A2(pi0969), .B(pi0299), .ZN(new_n5715_));
  NOR3_X1    g03199(.A1(new_n5537_), .A2(new_n5697_), .A3(new_n5706_), .ZN(new_n5716_));
  OR3_X2     g03200(.A1(new_n5715_), .A2(pi0232), .A3(new_n5716_), .Z(new_n5717_));
  NOR2_X1    g03201(.A1(new_n5716_), .A2(new_n5544_), .ZN(new_n5718_));
  OAI21_X1   g03202(.A1(new_n5543_), .A2(new_n5697_), .B(new_n5718_), .ZN(new_n5719_));
  OAI21_X1   g03203(.A1(new_n5549_), .A2(new_n5704_), .B(new_n2587_), .ZN(new_n5720_));
  NAND3_X1   g03204(.A1(new_n5720_), .A2(pi0232), .A3(new_n5719_), .ZN(new_n5721_));
  AOI21_X1   g03205(.A1(new_n5721_), .A2(new_n5717_), .B(pi0039), .ZN(new_n5722_));
  OAI22_X1   g03206(.A1(new_n5722_), .A2(new_n5714_), .B1(new_n5709_), .B2(new_n5712_), .ZN(new_n5723_));
  OAI21_X1   g03207(.A1(new_n5564_), .A2(new_n5704_), .B(new_n2587_), .ZN(new_n5724_));
  NAND4_X1   g03208(.A1(new_n5724_), .A2(pi0963), .A3(new_n2545_), .A4(new_n5707_), .ZN(new_n5725_));
  INV_X1     g03209(.I(new_n5711_), .ZN(new_n5726_));
  NOR2_X1    g03210(.A1(new_n5726_), .A2(new_n5567_), .ZN(new_n5727_));
  OAI21_X1   g03211(.A1(new_n5725_), .A2(new_n5560_), .B(new_n5727_), .ZN(new_n5728_));
  AOI21_X1   g03212(.A1(new_n5728_), .A2(new_n3177_), .B(pi0100), .ZN(new_n5729_));
  AOI22_X1   g03213(.A1(new_n5709_), .A2(new_n3207_), .B1(new_n2629_), .B2(new_n5711_), .ZN(new_n5730_));
  MUX2_X1    g03214(.I0(new_n5730_), .I1(new_n5726_), .S(new_n2628_), .Z(new_n5731_));
  INV_X1     g03215(.I(new_n5730_), .ZN(new_n5732_));
  OAI21_X1   g03216(.A1(new_n5726_), .A2(new_n3177_), .B(new_n5411_), .ZN(new_n5733_));
  AOI21_X1   g03217(.A1(new_n5732_), .A2(pi0075), .B(new_n5733_), .ZN(new_n5734_));
  OAI21_X1   g03218(.A1(pi0092), .A2(new_n5731_), .B(new_n5734_), .ZN(new_n5735_));
  AOI21_X1   g03219(.A1(new_n5723_), .A2(new_n5729_), .B(new_n5735_), .ZN(new_n5736_));
  NOR2_X1    g03220(.A1(new_n5732_), .A2(new_n3228_), .ZN(new_n5737_));
  OAI21_X1   g03221(.A1(new_n5726_), .A2(new_n3209_), .B(pi0054), .ZN(new_n5738_));
  OAI21_X1   g03222(.A1(new_n5737_), .A2(new_n5738_), .B(new_n3202_), .ZN(new_n5739_));
  NOR2_X1    g03223(.A1(new_n5582_), .A2(pi0074), .ZN(new_n5740_));
  AOI21_X1   g03224(.A1(new_n5732_), .A2(new_n5740_), .B(pi0055), .ZN(new_n5741_));
  OAI21_X1   g03225(.A1(new_n5736_), .A2(new_n5739_), .B(new_n5741_), .ZN(new_n5742_));
  AOI21_X1   g03226(.A1(new_n5699_), .A2(new_n5702_), .B(new_n5586_), .ZN(new_n5743_));
  NAND2_X1   g03227(.A1(new_n5702_), .A2(new_n5224_), .ZN(new_n5744_));
  AOI21_X1   g03228(.A1(new_n5701_), .A2(new_n3503_), .B(pi0059), .ZN(new_n5745_));
  OAI21_X1   g03229(.A1(new_n5699_), .A2(new_n5744_), .B(new_n5745_), .ZN(new_n5746_));
  AOI21_X1   g03230(.A1(new_n5742_), .A2(new_n5743_), .B(new_n5746_), .ZN(new_n5747_));
  OAI22_X1   g03231(.A1(new_n5747_), .A2(pi0057), .B1(new_n5700_), .B2(new_n5703_), .ZN(po0176));
  INV_X1     g03232(.I(pi0975), .ZN(new_n5749_));
  NOR2_X1    g03233(.A1(new_n5505_), .A2(new_n5749_), .ZN(new_n5750_));
  NAND2_X1   g03234(.A1(new_n5750_), .A2(new_n3233_), .ZN(new_n5751_));
  NOR2_X1    g03235(.A1(new_n5751_), .A2(new_n5223_), .ZN(new_n5752_));
  NOR2_X1    g03236(.A1(new_n5510_), .A2(new_n5749_), .ZN(new_n5753_));
  INV_X1     g03237(.I(new_n5753_), .ZN(new_n5754_));
  NAND2_X1   g03238(.A1(new_n5754_), .A2(pi0057), .ZN(new_n5755_));
  INV_X1     g03239(.I(pi0971), .ZN(new_n5756_));
  OAI21_X1   g03240(.A1(new_n5517_), .A2(new_n5756_), .B(new_n2587_), .ZN(new_n5757_));
  NOR2_X1    g03241(.A1(new_n5753_), .A2(new_n2587_), .ZN(new_n5758_));
  INV_X1     g03242(.I(new_n5758_), .ZN(new_n5759_));
  NAND2_X1   g03243(.A1(new_n5750_), .A2(new_n5759_), .ZN(new_n5760_));
  NAND3_X1   g03244(.A1(new_n5757_), .A2(new_n5760_), .A3(new_n3154_), .ZN(new_n5761_));
  MUX2_X1    g03245(.I0(new_n5756_), .I1(new_n5749_), .S(pi0299), .Z(new_n5762_));
  NOR2_X1    g03246(.A1(new_n5510_), .A2(new_n5762_), .ZN(new_n5763_));
  NAND2_X1   g03247(.A1(new_n5763_), .A2(new_n5525_), .ZN(new_n5764_));
  OAI22_X1   g03248(.A1(new_n5531_), .A2(new_n5749_), .B1(new_n5756_), .B2(new_n5528_), .ZN(new_n5765_));
  AOI21_X1   g03249(.A1(new_n5765_), .A2(new_n5527_), .B(pi0038), .ZN(new_n5766_));
  AOI21_X1   g03250(.A1(new_n5534_), .A2(pi0971), .B(pi0299), .ZN(new_n5767_));
  NOR3_X1    g03251(.A1(new_n5537_), .A2(new_n5749_), .A3(new_n5758_), .ZN(new_n5768_));
  OR3_X2     g03252(.A1(new_n5767_), .A2(pi0232), .A3(new_n5768_), .Z(new_n5769_));
  NOR2_X1    g03253(.A1(new_n5768_), .A2(new_n5544_), .ZN(new_n5770_));
  OAI21_X1   g03254(.A1(new_n5543_), .A2(new_n5749_), .B(new_n5770_), .ZN(new_n5771_));
  OAI21_X1   g03255(.A1(new_n5549_), .A2(new_n5756_), .B(new_n2587_), .ZN(new_n5772_));
  NAND3_X1   g03256(.A1(new_n5772_), .A2(pi0232), .A3(new_n5771_), .ZN(new_n5773_));
  AOI21_X1   g03257(.A1(new_n5773_), .A2(new_n5769_), .B(pi0039), .ZN(new_n5774_));
  OAI22_X1   g03258(.A1(new_n5774_), .A2(new_n5766_), .B1(new_n5761_), .B2(new_n5764_), .ZN(new_n5775_));
  OAI21_X1   g03259(.A1(new_n5564_), .A2(new_n5756_), .B(new_n2587_), .ZN(new_n5776_));
  NAND4_X1   g03260(.A1(new_n5776_), .A2(pi0975), .A3(new_n2545_), .A4(new_n5759_), .ZN(new_n5777_));
  INV_X1     g03261(.I(new_n5763_), .ZN(new_n5778_));
  NOR2_X1    g03262(.A1(new_n5778_), .A2(new_n5567_), .ZN(new_n5779_));
  OAI21_X1   g03263(.A1(new_n5777_), .A2(new_n5560_), .B(new_n5779_), .ZN(new_n5780_));
  AOI21_X1   g03264(.A1(new_n5780_), .A2(new_n3177_), .B(pi0100), .ZN(new_n5781_));
  AOI22_X1   g03265(.A1(new_n5761_), .A2(new_n3207_), .B1(new_n2629_), .B2(new_n5763_), .ZN(new_n5782_));
  MUX2_X1    g03266(.I0(new_n5782_), .I1(new_n5778_), .S(new_n2628_), .Z(new_n5783_));
  INV_X1     g03267(.I(new_n5782_), .ZN(new_n5784_));
  OAI21_X1   g03268(.A1(new_n5778_), .A2(new_n3177_), .B(new_n5411_), .ZN(new_n5785_));
  AOI21_X1   g03269(.A1(new_n5784_), .A2(pi0075), .B(new_n5785_), .ZN(new_n5786_));
  OAI21_X1   g03270(.A1(pi0092), .A2(new_n5783_), .B(new_n5786_), .ZN(new_n5787_));
  AOI21_X1   g03271(.A1(new_n5775_), .A2(new_n5781_), .B(new_n5787_), .ZN(new_n5788_));
  NOR2_X1    g03272(.A1(new_n5784_), .A2(new_n3228_), .ZN(new_n5789_));
  OAI21_X1   g03273(.A1(new_n5778_), .A2(new_n3209_), .B(pi0054), .ZN(new_n5790_));
  OAI21_X1   g03274(.A1(new_n5789_), .A2(new_n5790_), .B(new_n3202_), .ZN(new_n5791_));
  NOR2_X1    g03275(.A1(new_n5582_), .A2(pi0074), .ZN(new_n5792_));
  AOI21_X1   g03276(.A1(new_n5784_), .A2(new_n5792_), .B(pi0055), .ZN(new_n5793_));
  OAI21_X1   g03277(.A1(new_n5788_), .A2(new_n5791_), .B(new_n5793_), .ZN(new_n5794_));
  AOI21_X1   g03278(.A1(new_n5751_), .A2(new_n5754_), .B(new_n5586_), .ZN(new_n5795_));
  NAND2_X1   g03279(.A1(new_n5754_), .A2(new_n5224_), .ZN(new_n5796_));
  AOI21_X1   g03280(.A1(new_n5753_), .A2(new_n3503_), .B(pi0059), .ZN(new_n5797_));
  OAI21_X1   g03281(.A1(new_n5751_), .A2(new_n5796_), .B(new_n5797_), .ZN(new_n5798_));
  AOI21_X1   g03282(.A1(new_n5794_), .A2(new_n5795_), .B(new_n5798_), .ZN(new_n5799_));
  OAI22_X1   g03283(.A1(new_n5799_), .A2(pi0057), .B1(new_n5752_), .B2(new_n5755_), .ZN(po0177));
  NAND4_X1   g03284(.A1(new_n5110_), .A2(new_n2523_), .A3(pi0978), .A4(new_n3233_), .ZN(new_n5801_));
  NOR2_X1    g03285(.A1(new_n5801_), .A2(new_n5223_), .ZN(new_n5802_));
  INV_X1     g03286(.I(pi0978), .ZN(new_n5803_));
  NOR2_X1    g03287(.A1(new_n5510_), .A2(new_n5803_), .ZN(new_n5804_));
  INV_X1     g03288(.I(new_n5804_), .ZN(new_n5805_));
  NAND2_X1   g03289(.A1(new_n5805_), .A2(pi0057), .ZN(new_n5806_));
  INV_X1     g03290(.I(pi0974), .ZN(new_n5807_));
  MUX2_X1    g03291(.I0(new_n5807_), .I1(new_n5803_), .S(pi0299), .Z(new_n5808_));
  NOR2_X1    g03292(.A1(new_n5517_), .A2(new_n5808_), .ZN(new_n5809_));
  INV_X1     g03293(.I(new_n5809_), .ZN(new_n5810_));
  NOR2_X1    g03294(.A1(new_n5510_), .A2(new_n5808_), .ZN(new_n5811_));
  INV_X1     g03295(.I(new_n5811_), .ZN(new_n5812_));
  NAND4_X1   g03296(.A1(new_n5810_), .A2(new_n3172_), .A3(pi0039), .A4(new_n5812_), .ZN(new_n5813_));
  OAI22_X1   g03297(.A1(new_n5531_), .A2(new_n5803_), .B1(new_n5807_), .B2(new_n5528_), .ZN(new_n5814_));
  AOI21_X1   g03298(.A1(new_n5814_), .A2(new_n5527_), .B(pi0038), .ZN(new_n5815_));
  AOI21_X1   g03299(.A1(new_n5534_), .A2(pi0974), .B(pi0299), .ZN(new_n5816_));
  NOR2_X1    g03300(.A1(new_n5804_), .A2(new_n2587_), .ZN(new_n5817_));
  NOR3_X1    g03301(.A1(new_n5537_), .A2(new_n5803_), .A3(new_n5817_), .ZN(new_n5818_));
  OR3_X2     g03302(.A1(new_n5816_), .A2(pi0232), .A3(new_n5818_), .Z(new_n5819_));
  NOR2_X1    g03303(.A1(new_n5818_), .A2(new_n5544_), .ZN(new_n5820_));
  OAI21_X1   g03304(.A1(new_n5543_), .A2(new_n5803_), .B(new_n5820_), .ZN(new_n5821_));
  OAI21_X1   g03305(.A1(new_n5549_), .A2(new_n5807_), .B(new_n2587_), .ZN(new_n5822_));
  NAND3_X1   g03306(.A1(new_n5822_), .A2(pi0232), .A3(new_n5821_), .ZN(new_n5823_));
  AOI21_X1   g03307(.A1(new_n5823_), .A2(new_n5819_), .B(pi0039), .ZN(new_n5824_));
  OAI21_X1   g03308(.A1(new_n5824_), .A2(new_n5815_), .B(new_n5813_), .ZN(new_n5825_));
  OAI21_X1   g03309(.A1(new_n5564_), .A2(new_n5807_), .B(new_n2587_), .ZN(new_n5826_));
  NOR3_X1    g03310(.A1(new_n5817_), .A2(new_n5803_), .A3(new_n2544_), .ZN(new_n5827_));
  NAND2_X1   g03311(.A1(new_n5826_), .A2(new_n5827_), .ZN(new_n5828_));
  NOR2_X1    g03312(.A1(new_n5812_), .A2(new_n5567_), .ZN(new_n5829_));
  OAI21_X1   g03313(.A1(new_n5828_), .A2(new_n5560_), .B(new_n5829_), .ZN(new_n5830_));
  AOI21_X1   g03314(.A1(new_n5830_), .A2(new_n3177_), .B(pi0100), .ZN(new_n5831_));
  AOI21_X1   g03315(.A1(new_n2523_), .A2(new_n2629_), .B(new_n5810_), .ZN(new_n5832_));
  INV_X1     g03316(.I(new_n5832_), .ZN(new_n5833_));
  OAI21_X1   g03317(.A1(new_n5833_), .A2(new_n5811_), .B(pi0075), .ZN(new_n5834_));
  NOR2_X1    g03318(.A1(new_n5812_), .A2(new_n3177_), .ZN(new_n5835_));
  NOR4_X1    g03319(.A1(new_n5832_), .A2(pi0075), .A3(new_n5410_), .A4(new_n5835_), .ZN(new_n5836_));
  OAI21_X1   g03320(.A1(new_n5834_), .A2(new_n3203_), .B(new_n5836_), .ZN(new_n5837_));
  AOI21_X1   g03321(.A1(new_n5825_), .A2(new_n5831_), .B(new_n5837_), .ZN(new_n5838_));
  NOR2_X1    g03322(.A1(new_n5833_), .A2(new_n3228_), .ZN(new_n5839_));
  OAI21_X1   g03323(.A1(new_n5812_), .A2(new_n3209_), .B(pi0054), .ZN(new_n5840_));
  OAI21_X1   g03324(.A1(new_n5839_), .A2(new_n5840_), .B(new_n3202_), .ZN(new_n5841_));
  NAND2_X1   g03325(.A1(new_n5833_), .A2(new_n3214_), .ZN(new_n5842_));
  NAND2_X1   g03326(.A1(new_n5812_), .A2(new_n5582_), .ZN(new_n5843_));
  AOI21_X1   g03327(.A1(new_n5843_), .A2(pi0074), .B(new_n3209_), .ZN(new_n5844_));
  AOI21_X1   g03328(.A1(new_n5842_), .A2(new_n5844_), .B(pi0055), .ZN(new_n5845_));
  OAI21_X1   g03329(.A1(new_n5838_), .A2(new_n5841_), .B(new_n5845_), .ZN(new_n5846_));
  AOI21_X1   g03330(.A1(new_n5801_), .A2(new_n5805_), .B(new_n5586_), .ZN(new_n5847_));
  NAND2_X1   g03331(.A1(new_n5805_), .A2(new_n5224_), .ZN(new_n5848_));
  AOI21_X1   g03332(.A1(new_n5804_), .A2(new_n3503_), .B(pi0059), .ZN(new_n5849_));
  OAI21_X1   g03333(.A1(new_n5801_), .A2(new_n5848_), .B(new_n5849_), .ZN(new_n5850_));
  AOI21_X1   g03334(.A1(new_n5846_), .A2(new_n5847_), .B(new_n5850_), .ZN(new_n5851_));
  OAI22_X1   g03335(.A1(new_n5851_), .A2(pi0057), .B1(new_n5802_), .B2(new_n5806_), .ZN(po0178));
  NOR3_X1    g03336(.A1(new_n5332_), .A2(new_n2587_), .A3(new_n5342_), .ZN(new_n5853_));
  NOR2_X1    g03337(.A1(new_n2587_), .A2(pi0232), .ZN(new_n5854_));
  INV_X1     g03338(.I(new_n5854_), .ZN(new_n5855_));
  NOR4_X1    g03339(.A1(new_n5334_), .A2(new_n5343_), .A3(new_n5853_), .A4(new_n5855_), .ZN(new_n5856_));
  AOI21_X1   g03340(.A1(new_n5108_), .A2(new_n5327_), .B(new_n5319_), .ZN(new_n5857_));
  NOR2_X1    g03341(.A1(new_n5318_), .A2(new_n5442_), .ZN(new_n5858_));
  OAI21_X1   g03342(.A1(new_n5857_), .A2(pi0299), .B(new_n5858_), .ZN(new_n5859_));
  AOI21_X1   g03343(.A1(new_n5541_), .A2(new_n5856_), .B(new_n5859_), .ZN(new_n5860_));
  AOI21_X1   g03344(.A1(new_n2587_), .A2(new_n5298_), .B(new_n5332_), .ZN(new_n5861_));
  NOR3_X1    g03345(.A1(new_n5333_), .A2(pi0299), .A3(new_n5298_), .ZN(new_n5862_));
  NOR2_X1    g03346(.A1(pi0039), .A2(pi0232), .ZN(new_n5863_));
  INV_X1     g03347(.I(new_n5863_), .ZN(new_n5864_));
  NOR4_X1    g03348(.A1(new_n5860_), .A2(new_n5861_), .A3(new_n5862_), .A4(new_n5864_), .ZN(new_n5865_));
  INV_X1     g03349(.I(new_n5133_), .ZN(new_n5866_));
  NOR3_X1    g03350(.A1(new_n5866_), .A2(new_n3154_), .A3(new_n2587_), .ZN(new_n5867_));
  AOI21_X1   g03351(.A1(new_n5529_), .A2(new_n5867_), .B(pi0038), .ZN(new_n5868_));
  INV_X1     g03352(.I(new_n5868_), .ZN(new_n5869_));
  AOI21_X1   g03353(.A1(new_n5153_), .A2(pi0038), .B(new_n3173_), .ZN(new_n5870_));
  OAI21_X1   g03354(.A1(new_n5865_), .A2(new_n5869_), .B(new_n5870_), .ZN(new_n5871_));
  NOR2_X1    g03355(.A1(new_n5157_), .A2(pi0038), .ZN(new_n5872_));
  INV_X1     g03356(.I(new_n5872_), .ZN(new_n5873_));
  OAI21_X1   g03357(.A1(new_n3173_), .A2(new_n5873_), .B(new_n5871_), .ZN(new_n5874_));
  NOR2_X1    g03358(.A1(new_n5157_), .A2(new_n3208_), .ZN(new_n5875_));
  NOR2_X1    g03359(.A1(new_n5875_), .A2(new_n2628_), .ZN(new_n5876_));
  NOR2_X1    g03360(.A1(new_n2535_), .A2(new_n2622_), .ZN(new_n5877_));
  NAND2_X1   g03361(.A1(new_n5156_), .A2(new_n5877_), .ZN(new_n5878_));
  INV_X1     g03362(.I(new_n5878_), .ZN(new_n5879_));
  NOR2_X1    g03363(.A1(new_n5879_), .A2(new_n3203_), .ZN(new_n5880_));
  NOR2_X1    g03364(.A1(new_n5876_), .A2(new_n5880_), .ZN(new_n5881_));
  NOR2_X1    g03365(.A1(new_n5881_), .A2(new_n3228_), .ZN(new_n5882_));
  INV_X1     g03366(.I(new_n5882_), .ZN(new_n5883_));
  AOI21_X1   g03367(.A1(new_n5874_), .A2(new_n5189_), .B(new_n5883_), .ZN(new_n5884_));
  OAI21_X1   g03368(.A1(new_n5884_), .A2(pi0054), .B(new_n3202_), .ZN(new_n5886_));
  NOR2_X1    g03369(.A1(new_n5195_), .A2(new_n2541_), .ZN(new_n5887_));
  INV_X1     g03370(.I(new_n5887_), .ZN(new_n5888_));
  NOR2_X1    g03371(.A1(new_n5888_), .A2(pi0055), .ZN(new_n5889_));
  NOR2_X1    g03372(.A1(new_n5889_), .A2(pi0056), .ZN(new_n5890_));
  NOR2_X1    g03373(.A1(new_n5890_), .A2(pi0062), .ZN(new_n5891_));
  INV_X1     g03374(.I(new_n5891_), .ZN(new_n5892_));
  AOI21_X1   g03375(.A1(new_n5886_), .A2(new_n5199_), .B(new_n5892_), .ZN(new_n5893_));
  OAI21_X1   g03376(.A1(new_n5893_), .A2(new_n3405_), .B(new_n5208_), .ZN(new_n5894_));
  INV_X1     g03377(.I(pi0024), .ZN(new_n5895_));
  NAND2_X1   g03378(.A1(new_n5895_), .A2(pi0954), .ZN(new_n5896_));
  OAI21_X1   g03379(.A1(new_n5894_), .A2(pi0954), .B(new_n5896_), .ZN(po0182));
  OAI21_X1   g03380(.A1(new_n5161_), .A2(new_n3181_), .B(new_n2587_), .ZN(new_n5898_));
  OAI22_X1   g03381(.A1(new_n3256_), .A2(new_n2587_), .B1(new_n2491_), .B2(new_n5898_), .ZN(new_n5899_));
  INV_X1     g03382(.I(new_n5899_), .ZN(new_n5900_));
  NOR3_X1    g03383(.A1(new_n5900_), .A2(new_n3173_), .A3(new_n3311_), .ZN(new_n5901_));
  NOR2_X1    g03384(.A1(pi0100), .A2(pi0228), .ZN(new_n5902_));
  NOR4_X1    g03385(.A1(new_n3377_), .A2(pi0039), .A3(new_n5901_), .A4(new_n5902_), .ZN(new_n5903_));
  NOR2_X1    g03386(.A1(pi0039), .A2(pi0100), .ZN(new_n5904_));
  AOI21_X1   g03387(.A1(new_n3310_), .A2(new_n5904_), .B(pi0038), .ZN(new_n5905_));
  OAI21_X1   g03388(.A1(new_n5903_), .A2(new_n5905_), .B(new_n2525_), .ZN(new_n5906_));
  NOR2_X1    g03389(.A1(new_n3311_), .A2(new_n2547_), .ZN(new_n5907_));
  OAI21_X1   g03390(.A1(new_n5907_), .A2(new_n2524_), .B(pi0087), .ZN(new_n5908_));
  NAND2_X1   g03391(.A1(new_n5908_), .A2(new_n2628_), .ZN(new_n5909_));
  NOR2_X1    g03392(.A1(new_n3311_), .A2(new_n3323_), .ZN(new_n5910_));
  NOR2_X1    g03393(.A1(new_n2538_), .A2(new_n3203_), .ZN(new_n5911_));
  OAI21_X1   g03394(.A1(new_n5910_), .A2(new_n2524_), .B(new_n5911_), .ZN(new_n5912_));
  OAI21_X1   g03395(.A1(new_n2524_), .A2(new_n2628_), .B(new_n3203_), .ZN(new_n5913_));
  NAND3_X1   g03396(.A1(new_n5909_), .A2(new_n5912_), .A3(new_n5913_), .ZN(new_n5914_));
  AOI21_X1   g03397(.A1(new_n5906_), .A2(new_n3177_), .B(new_n5914_), .ZN(new_n5915_));
  NOR2_X1    g03398(.A1(new_n2524_), .A2(new_n2538_), .ZN(new_n5916_));
  OAI21_X1   g03399(.A1(new_n5915_), .A2(pi0055), .B(new_n5916_), .ZN(new_n5917_));
  NOR2_X1    g03400(.A1(new_n5197_), .A2(new_n2547_), .ZN(new_n5918_));
  NAND3_X1   g03401(.A1(new_n3310_), .A2(new_n3202_), .A3(new_n5918_), .ZN(new_n5919_));
  AOI21_X1   g03402(.A1(new_n5919_), .A2(new_n2525_), .B(pi0055), .ZN(new_n5920_));
  NAND2_X1   g03403(.A1(new_n3310_), .A2(new_n2548_), .ZN(new_n5921_));
  OAI21_X1   g03404(.A1(new_n5921_), .A2(new_n2524_), .B(new_n3335_), .ZN(new_n5922_));
  NOR2_X1    g03405(.A1(new_n5920_), .A2(new_n5922_), .ZN(new_n5923_));
  AOI21_X1   g03406(.A1(new_n5917_), .A2(new_n5923_), .B(pi0062), .ZN(new_n5924_));
  NAND2_X1   g03407(.A1(new_n5907_), .A2(new_n3341_), .ZN(new_n5925_));
  NAND3_X1   g03408(.A1(new_n5925_), .A2(pi0062), .A3(new_n2525_), .ZN(new_n5926_));
  NAND2_X1   g03409(.A1(new_n5926_), .A2(new_n2571_), .ZN(new_n5927_));
  OAI22_X1   g03410(.A1(new_n5924_), .A2(new_n5927_), .B1(new_n2525_), .B2(new_n2571_), .ZN(po0183));
  INV_X1     g03411(.I(pi0119), .ZN(new_n5929_));
  NAND2_X1   g03412(.A1(new_n2523_), .A2(pi0252), .ZN(new_n5930_));
  AOI21_X1   g03413(.A1(new_n5930_), .A2(new_n5929_), .B(pi0468), .ZN(new_n5931_));
  NAND2_X1   g03414(.A1(pi0119), .A2(pi1056), .ZN(new_n5932_));
  NAND2_X1   g03415(.A1(new_n5931_), .A2(new_n5932_), .ZN(po0184));
  NAND2_X1   g03416(.A1(pi0119), .A2(pi1077), .ZN(new_n5934_));
  NAND2_X1   g03417(.A1(new_n5931_), .A2(new_n5934_), .ZN(po0185));
  NAND2_X1   g03418(.A1(pi0119), .A2(pi1073), .ZN(new_n5936_));
  NAND2_X1   g03419(.A1(new_n5931_), .A2(new_n5936_), .ZN(po0186));
  NAND2_X1   g03420(.A1(pi0119), .A2(pi1041), .ZN(new_n5938_));
  NAND2_X1   g03421(.A1(new_n5931_), .A2(new_n5938_), .ZN(po0187));
  INV_X1     g03422(.I(pi0591), .ZN(new_n5940_));
  NOR2_X1    g03423(.A1(new_n5410_), .A2(pi0074), .ZN(new_n5941_));
  INV_X1     g03424(.I(new_n5941_), .ZN(new_n5942_));
  INV_X1     g03425(.I(po0740), .ZN(new_n5943_));
  NOR2_X1    g03426(.A1(new_n2491_), .A2(new_n5943_), .ZN(new_n5944_));
  NOR2_X1    g03427(.A1(new_n2927_), .A2(pi0122), .ZN(new_n5945_));
  INV_X1     g03428(.I(new_n5945_), .ZN(new_n5946_));
  NOR2_X1    g03429(.A1(new_n5946_), .A2(new_n2955_), .ZN(new_n5947_));
  INV_X1     g03430(.I(new_n5947_), .ZN(new_n5948_));
  NAND2_X1   g03431(.A1(new_n2641_), .A2(new_n2902_), .ZN(new_n5949_));
  OAI21_X1   g03432(.A1(new_n5949_), .A2(new_n2839_), .B(new_n2841_), .ZN(new_n5950_));
  NOR2_X1    g03433(.A1(pi0035), .A2(pi0070), .ZN(new_n5951_));
  NAND2_X1   g03434(.A1(new_n5059_), .A2(new_n5951_), .ZN(new_n5952_));
  OAI21_X1   g03435(.A1(new_n5950_), .A2(new_n5952_), .B(new_n2658_), .ZN(new_n5953_));
  INV_X1     g03436(.I(new_n5953_), .ZN(new_n5954_));
  NOR2_X1    g03437(.A1(pi0050), .A2(pi0077), .ZN(new_n5955_));
  INV_X1     g03438(.I(new_n5955_), .ZN(new_n5956_));
  NOR2_X1    g03439(.A1(new_n5956_), .A2(pi0094), .ZN(new_n5957_));
  INV_X1     g03440(.I(new_n5957_), .ZN(new_n5958_));
  NOR2_X1    g03441(.A1(new_n2703_), .A2(new_n5958_), .ZN(new_n5959_));
  NAND4_X1   g03442(.A1(new_n5959_), .A2(new_n2710_), .A3(pi0098), .A4(new_n2467_), .ZN(new_n5960_));
  INV_X1     g03443(.I(new_n5960_), .ZN(new_n5961_));
  NOR2_X1    g03444(.A1(new_n5961_), .A2(pi0097), .ZN(new_n5962_));
  NOR2_X1    g03445(.A1(new_n5962_), .A2(new_n2890_), .ZN(new_n5963_));
  NOR2_X1    g03446(.A1(new_n2650_), .A2(pi0035), .ZN(new_n5964_));
  INV_X1     g03447(.I(new_n5964_), .ZN(new_n5965_));
  NOR2_X1    g03448(.A1(new_n5965_), .A2(pi0070), .ZN(new_n5966_));
  NAND2_X1   g03449(.A1(new_n5963_), .A2(new_n5966_), .ZN(new_n5967_));
  OAI22_X1   g03450(.A1(new_n5954_), .A2(new_n5967_), .B1(new_n2658_), .B2(new_n2673_), .ZN(new_n5968_));
  NOR2_X1    g03451(.A1(new_n5968_), .A2(pi0096), .ZN(new_n5969_));
  NOR4_X1    g03452(.A1(new_n2501_), .A2(pi0093), .A3(pi0841), .A4(new_n2480_), .ZN(new_n5970_));
  AOI21_X1   g03453(.A1(new_n5970_), .A2(new_n2665_), .B(new_n2659_), .ZN(new_n5971_));
  NOR2_X1    g03454(.A1(new_n5971_), .A2(new_n2485_), .ZN(new_n5972_));
  INV_X1     g03455(.I(new_n5972_), .ZN(new_n5973_));
  NOR3_X1    g03456(.A1(new_n5969_), .A2(new_n5948_), .A3(new_n5973_), .ZN(new_n5974_));
  NOR2_X1    g03457(.A1(new_n2485_), .A2(pi0096), .ZN(new_n5975_));
  NAND2_X1   g03458(.A1(new_n5968_), .A2(new_n5975_), .ZN(new_n5976_));
  NOR3_X1    g03459(.A1(new_n5976_), .A2(new_n5182_), .A3(new_n5945_), .ZN(new_n5977_));
  NOR3_X1    g03460(.A1(new_n5974_), .A2(new_n5977_), .A3(pi1093), .ZN(new_n5978_));
  NOR2_X1    g03461(.A1(new_n2547_), .A2(pi0075), .ZN(new_n5979_));
  INV_X1     g03462(.I(new_n5979_), .ZN(new_n5980_));
  NAND4_X1   g03463(.A1(new_n5978_), .A2(new_n3177_), .A3(new_n5944_), .A4(new_n5980_), .ZN(new_n5981_));
  INV_X1     g03464(.I(new_n5981_), .ZN(new_n5982_));
  NOR2_X1    g03465(.A1(new_n2576_), .A2(new_n2587_), .ZN(new_n5983_));
  NOR2_X1    g03466(.A1(new_n2605_), .A2(pi0299), .ZN(new_n5984_));
  NOR2_X1    g03467(.A1(new_n5983_), .A2(new_n5984_), .ZN(new_n5985_));
  INV_X1     g03468(.I(new_n5985_), .ZN(new_n5986_));
  INV_X1     g03469(.I(pi0232), .ZN(new_n5987_));
  NOR2_X1    g03470(.A1(new_n5109_), .A2(new_n5987_), .ZN(new_n5988_));
  INV_X1     g03471(.I(new_n5988_), .ZN(new_n5989_));
  NOR2_X1    g03472(.A1(new_n5986_), .A2(new_n5989_), .ZN(new_n5990_));
  NOR2_X1    g03473(.A1(new_n5990_), .A2(new_n2629_), .ZN(new_n5991_));
  NOR2_X1    g03474(.A1(new_n3181_), .A2(pi0024), .ZN(new_n5992_));
  INV_X1     g03475(.I(new_n5992_), .ZN(new_n5993_));
  NOR2_X1    g03476(.A1(new_n2491_), .A2(new_n5993_), .ZN(new_n5994_));
  NOR2_X1    g03477(.A1(new_n5177_), .A2(new_n2920_), .ZN(new_n5995_));
  NOR2_X1    g03478(.A1(new_n5948_), .A2(new_n2918_), .ZN(new_n5996_));
  NAND3_X1   g03479(.A1(new_n5995_), .A2(new_n5994_), .A3(new_n5996_), .ZN(new_n5997_));
  NOR2_X1    g03480(.A1(new_n5997_), .A2(new_n2924_), .ZN(new_n5998_));
  AOI21_X1   g03481(.A1(new_n5998_), .A2(new_n5991_), .B(new_n2628_), .ZN(new_n5999_));
  NAND2_X1   g03482(.A1(new_n2920_), .A2(pi1093), .ZN(new_n6000_));
  NAND3_X1   g03483(.A1(new_n2490_), .A2(new_n5181_), .A3(new_n6000_), .ZN(new_n6001_));
  INV_X1     g03484(.I(new_n6001_), .ZN(new_n6002_));
  NOR2_X1    g03485(.A1(new_n2924_), .A2(pi1091), .ZN(new_n6003_));
  NOR2_X1    g03486(.A1(new_n2955_), .A2(new_n5366_), .ZN(new_n6004_));
  INV_X1     g03487(.I(new_n6004_), .ZN(new_n6005_));
  NOR2_X1    g03488(.A1(new_n2491_), .A2(new_n6005_), .ZN(new_n6006_));
  NOR2_X1    g03489(.A1(new_n6002_), .A2(new_n6003_), .ZN(new_n6007_));
  NOR3_X1    g03490(.A1(new_n6007_), .A2(pi0087), .A3(new_n3197_), .ZN(new_n6008_));
  INV_X1     g03491(.I(new_n6008_), .ZN(new_n6009_));
  NOR2_X1    g03492(.A1(new_n5948_), .A2(new_n2924_), .ZN(new_n6010_));
  INV_X1     g03493(.I(new_n5995_), .ZN(new_n6011_));
  NOR2_X1    g03494(.A1(new_n6011_), .A2(new_n2491_), .ZN(new_n6012_));
  NAND2_X1   g03495(.A1(new_n6012_), .A2(new_n6010_), .ZN(new_n6013_));
  NOR2_X1    g03496(.A1(new_n6013_), .A2(new_n2918_), .ZN(new_n6014_));
  NOR4_X1    g03497(.A1(new_n5990_), .A2(pi0100), .A3(new_n2523_), .A4(new_n2545_), .ZN(new_n6015_));
  NAND2_X1   g03498(.A1(new_n6014_), .A2(new_n6015_), .ZN(new_n6016_));
  INV_X1     g03499(.I(new_n5952_), .ZN(new_n6017_));
  INV_X1     g03500(.I(new_n2844_), .ZN(new_n6018_));
  NOR2_X1    g03501(.A1(new_n6018_), .A2(pi0024), .ZN(new_n6019_));
  INV_X1     g03502(.I(new_n6019_), .ZN(new_n6020_));
  NAND2_X1   g03503(.A1(new_n5062_), .A2(pi0097), .ZN(new_n6021_));
  NOR4_X1    g03504(.A1(new_n5304_), .A2(pi0046), .A3(pi0091), .A4(new_n6021_), .ZN(new_n6022_));
  NAND2_X1   g03505(.A1(new_n2688_), .A2(new_n6022_), .ZN(new_n6023_));
  NAND2_X1   g03506(.A1(new_n6020_), .A2(new_n6023_), .ZN(new_n6024_));
  NAND3_X1   g03507(.A1(new_n6024_), .A2(new_n2479_), .A3(new_n6017_), .ZN(new_n6025_));
  AOI21_X1   g03508(.A1(new_n6025_), .A2(new_n5954_), .B(new_n2674_), .ZN(new_n6026_));
  NOR2_X1    g03509(.A1(new_n5973_), .A2(new_n2957_), .ZN(new_n6027_));
  OAI21_X1   g03510(.A1(new_n6026_), .A2(pi0096), .B(new_n6027_), .ZN(new_n6028_));
  INV_X1     g03511(.I(pi0122), .ZN(new_n6029_));
  NOR2_X1    g03512(.A1(new_n2676_), .A2(new_n2485_), .ZN(new_n6030_));
  NAND2_X1   g03513(.A1(new_n5953_), .A2(new_n6030_), .ZN(new_n6031_));
  NOR2_X1    g03514(.A1(new_n6031_), .A2(new_n6005_), .ZN(new_n6032_));
  AOI21_X1   g03515(.A1(new_n6032_), .A2(new_n2927_), .B(new_n6029_), .ZN(new_n6033_));
  NAND2_X1   g03516(.A1(new_n6028_), .A2(new_n6033_), .ZN(new_n6034_));
  NOR3_X1    g03517(.A1(new_n6031_), .A2(pi0122), .A3(new_n5182_), .ZN(new_n6035_));
  NOR2_X1    g03518(.A1(new_n2920_), .A2(new_n2924_), .ZN(new_n6036_));
  INV_X1     g03519(.I(new_n6036_), .ZN(new_n6037_));
  AOI21_X1   g03520(.A1(new_n6034_), .A2(new_n6035_), .B(new_n6037_), .ZN(new_n6038_));
  OAI21_X1   g03521(.A1(new_n6034_), .A2(new_n6035_), .B(new_n6038_), .ZN(new_n6039_));
  NAND2_X1   g03522(.A1(new_n6039_), .A2(pi1091), .ZN(new_n6040_));
  NOR2_X1    g03523(.A1(new_n5978_), .A2(pi1091), .ZN(new_n6041_));
  INV_X1     g03524(.I(new_n6041_), .ZN(new_n6042_));
  OAI21_X1   g03525(.A1(new_n6040_), .A2(new_n5978_), .B(new_n6042_), .ZN(new_n6043_));
  NAND3_X1   g03526(.A1(new_n5362_), .A2(new_n2958_), .A3(new_n2929_), .ZN(new_n6044_));
  NOR2_X1    g03527(.A1(new_n6044_), .A2(new_n2926_), .ZN(new_n6045_));
  INV_X1     g03528(.I(new_n6045_), .ZN(new_n6046_));
  NOR2_X1    g03529(.A1(new_n6046_), .A2(new_n2918_), .ZN(new_n6047_));
  INV_X1     g03530(.I(new_n6047_), .ZN(new_n6048_));
  NOR2_X1    g03531(.A1(new_n6048_), .A2(new_n5145_), .ZN(new_n6049_));
  NOR2_X1    g03532(.A1(new_n2588_), .A2(pi0223), .ZN(new_n6050_));
  INV_X1     g03533(.I(new_n6050_), .ZN(new_n6051_));
  NOR4_X1    g03534(.A1(new_n6051_), .A2(pi0039), .A3(pi0224), .A4(pi0299), .ZN(new_n6052_));
  NAND2_X1   g03535(.A1(new_n6049_), .A2(new_n6052_), .ZN(new_n6053_));
  NOR2_X1    g03536(.A1(new_n6048_), .A2(new_n5866_), .ZN(new_n6054_));
  NOR3_X1    g03537(.A1(new_n5357_), .A2(pi0216), .A3(new_n2587_), .ZN(new_n6055_));
  NAND3_X1   g03538(.A1(new_n6053_), .A2(new_n6054_), .A3(new_n6055_), .ZN(new_n6056_));
  NAND2_X1   g03539(.A1(new_n6056_), .A2(new_n3172_), .ZN(new_n6057_));
  NOR2_X1    g03540(.A1(new_n6057_), .A2(pi0039), .ZN(new_n6058_));
  AOI21_X1   g03541(.A1(new_n6058_), .A2(new_n6043_), .B(pi0100), .ZN(new_n6059_));
  INV_X1     g03542(.I(new_n6059_), .ZN(new_n6060_));
  INV_X1     g03543(.I(new_n5369_), .ZN(new_n6061_));
  INV_X1     g03544(.I(new_n6040_), .ZN(new_n6062_));
  INV_X1     g03545(.I(new_n6057_), .ZN(new_n6063_));
  NOR4_X1    g03546(.A1(new_n6063_), .A2(new_n6061_), .A3(new_n6031_), .A4(new_n6062_), .ZN(new_n6064_));
  OAI21_X1   g03547(.A1(new_n6060_), .A2(new_n6064_), .B(new_n6016_), .ZN(new_n6065_));
  NAND2_X1   g03548(.A1(new_n6065_), .A2(new_n3177_), .ZN(new_n6066_));
  AOI21_X1   g03549(.A1(new_n6066_), .A2(new_n6009_), .B(pi0075), .ZN(new_n6067_));
  NOR2_X1    g03550(.A1(new_n6067_), .A2(new_n5999_), .ZN(new_n6068_));
  NOR3_X1    g03551(.A1(new_n5982_), .A2(pi0567), .A3(new_n5942_), .ZN(new_n6069_));
  INV_X1     g03552(.I(new_n6069_), .ZN(new_n6070_));
  INV_X1     g03553(.I(new_n5999_), .ZN(new_n6071_));
  NOR3_X1    g03554(.A1(new_n2545_), .A2(new_n3177_), .A3(pi0100), .ZN(new_n6072_));
  NAND2_X1   g03555(.A1(new_n6002_), .A2(new_n2918_), .ZN(new_n6073_));
  NOR2_X1    g03556(.A1(new_n5944_), .A2(pi1091), .ZN(new_n6074_));
  INV_X1     g03557(.I(new_n6074_), .ZN(new_n6075_));
  AOI21_X1   g03558(.A1(new_n6075_), .A2(new_n6073_), .B(new_n6072_), .ZN(new_n6076_));
  INV_X1     g03559(.I(new_n6016_), .ZN(new_n6077_));
  NOR2_X1    g03560(.A1(new_n6077_), .A2(pi0087), .ZN(new_n6078_));
  INV_X1     g03561(.I(new_n6078_), .ZN(new_n6079_));
  OAI22_X1   g03562(.A1(new_n6059_), .A2(new_n6079_), .B1(pi0075), .B2(new_n6076_), .ZN(new_n6080_));
  NAND2_X1   g03563(.A1(new_n6080_), .A2(new_n6071_), .ZN(new_n6081_));
  NAND2_X1   g03564(.A1(new_n6081_), .A2(pi0567), .ZN(new_n6082_));
  NOR2_X1    g03565(.A1(new_n6082_), .A2(pi0592), .ZN(new_n6083_));
  INV_X1     g03566(.I(pi0592), .ZN(new_n6084_));
  NOR2_X1    g03567(.A1(new_n6070_), .A2(new_n6084_), .ZN(new_n6085_));
  NOR2_X1    g03568(.A1(new_n6083_), .A2(new_n6085_), .ZN(new_n6086_));
  INV_X1     g03569(.I(new_n6086_), .ZN(new_n6087_));
  INV_X1     g03570(.I(pi1199), .ZN(new_n6088_));
  NOR2_X1    g03571(.A1(new_n6088_), .A2(pi0351), .ZN(new_n6089_));
  INV_X1     g03572(.I(pi1197), .ZN(new_n6090_));
  XNOR2_X1   g03573(.A1(pi0345), .A2(pi0346), .ZN(new_n6091_));
  NOR2_X1    g03574(.A1(pi0345), .A2(pi0346), .ZN(new_n6092_));
  INV_X1     g03575(.I(pi0345), .ZN(new_n6093_));
  INV_X1     g03576(.I(pi0346), .ZN(new_n6094_));
  NOR2_X1    g03577(.A1(new_n6093_), .A2(new_n6094_), .ZN(new_n6095_));
  OAI21_X1   g03578(.A1(new_n6095_), .A2(new_n6092_), .B(pi0323), .ZN(new_n6096_));
  OAI21_X1   g03579(.A1(pi0323), .A2(new_n6091_), .B(new_n6096_), .ZN(new_n6097_));
  XNOR2_X1   g03580(.A1(pi0358), .A2(pi0450), .ZN(new_n6098_));
  XNOR2_X1   g03581(.A1(pi0358), .A2(pi0450), .ZN(new_n6099_));
  NAND2_X1   g03582(.A1(new_n6097_), .A2(new_n6099_), .ZN(new_n6100_));
  OAI21_X1   g03583(.A1(new_n6097_), .A2(new_n6098_), .B(new_n6100_), .ZN(new_n6101_));
  INV_X1     g03584(.I(pi0362), .ZN(new_n6102_));
  XOR2_X1    g03585(.A1(pi0327), .A2(pi0343), .Z(new_n6103_));
  XOR2_X1    g03586(.A1(new_n6103_), .A2(new_n6102_), .Z(new_n6104_));
  XOR2_X1    g03587(.A1(new_n6104_), .A2(pi0344), .Z(new_n6105_));
  XOR2_X1    g03588(.A1(new_n6105_), .A2(new_n6101_), .Z(new_n6106_));
  NOR2_X1    g03589(.A1(new_n6106_), .A2(new_n6090_), .ZN(new_n6107_));
  INV_X1     g03590(.I(pi0350), .ZN(new_n6108_));
  NOR2_X1    g03591(.A1(new_n6108_), .A2(pi0592), .ZN(new_n6109_));
  INV_X1     g03592(.I(new_n6109_), .ZN(new_n6110_));
  INV_X1     g03593(.I(new_n6082_), .ZN(new_n6111_));
  XOR2_X1    g03594(.A1(pi0322), .A2(pi0359), .Z(new_n6112_));
  INV_X1     g03595(.I(pi0322), .ZN(new_n6113_));
  NOR2_X1    g03596(.A1(new_n6113_), .A2(pi0359), .ZN(new_n6114_));
  INV_X1     g03597(.I(pi0359), .ZN(new_n6115_));
  NOR2_X1    g03598(.A1(new_n6115_), .A2(pi0322), .ZN(new_n6116_));
  OAI21_X1   g03599(.A1(new_n6114_), .A2(new_n6116_), .B(pi0315), .ZN(new_n6117_));
  OAI21_X1   g03600(.A1(pi0315), .A2(new_n6112_), .B(new_n6117_), .ZN(new_n6118_));
  XNOR2_X1   g03601(.A1(new_n6118_), .A2(pi0316), .ZN(new_n6119_));
  XOR2_X1    g03602(.A1(new_n6119_), .A2(pi0349), .Z(new_n6120_));
  XOR2_X1    g03603(.A1(new_n6120_), .A2(pi0348), .Z(new_n6121_));
  XOR2_X1    g03604(.A1(pi0321), .A2(pi0347), .Z(new_n6122_));
  INV_X1     g03605(.I(new_n6122_), .ZN(new_n6123_));
  XNOR2_X1   g03606(.A1(pi0321), .A2(pi0347), .ZN(new_n6124_));
  NOR2_X1    g03607(.A1(new_n6121_), .A2(new_n6124_), .ZN(new_n6125_));
  AOI21_X1   g03608(.A1(new_n6121_), .A2(new_n6123_), .B(new_n6125_), .ZN(new_n6126_));
  OAI21_X1   g03609(.A1(new_n6111_), .A2(new_n6110_), .B(new_n6126_), .ZN(new_n6127_));
  INV_X1     g03610(.I(pi0355), .ZN(new_n6130_));
  INV_X1     g03611(.I(pi0458), .ZN(new_n6131_));
  INV_X1     g03612(.I(pi0320), .ZN(new_n6132_));
  INV_X1     g03613(.I(pi0342), .ZN(new_n6133_));
  NOR2_X1    g03614(.A1(new_n6133_), .A2(pi0460), .ZN(new_n6134_));
  INV_X1     g03615(.I(pi0460), .ZN(new_n6135_));
  NOR2_X1    g03616(.A1(new_n6135_), .A2(pi0342), .ZN(new_n6136_));
  OAI21_X1   g03617(.A1(new_n6134_), .A2(new_n6136_), .B(new_n6132_), .ZN(new_n6137_));
  NOR2_X1    g03618(.A1(pi0342), .A2(pi0460), .ZN(new_n6138_));
  NOR2_X1    g03619(.A1(new_n6133_), .A2(new_n6135_), .ZN(new_n6139_));
  OAI21_X1   g03620(.A1(new_n6139_), .A2(new_n6138_), .B(pi0320), .ZN(new_n6140_));
  NAND2_X1   g03621(.A1(new_n6140_), .A2(new_n6137_), .ZN(new_n6141_));
  XOR2_X1    g03622(.A1(pi0361), .A2(pi0441), .Z(new_n6142_));
  NOR2_X1    g03623(.A1(new_n6141_), .A2(new_n6142_), .ZN(new_n6143_));
  INV_X1     g03624(.I(new_n6141_), .ZN(new_n6144_));
  XNOR2_X1   g03625(.A1(pi0361), .A2(pi0441), .ZN(new_n6145_));
  NOR2_X1    g03626(.A1(new_n6144_), .A2(new_n6145_), .ZN(new_n6146_));
  NOR2_X1    g03627(.A1(new_n6146_), .A2(new_n6143_), .ZN(new_n6147_));
  XOR2_X1    g03628(.A1(new_n6147_), .A2(new_n6131_), .Z(new_n6148_));
  XOR2_X1    g03629(.A1(pi0452), .A2(pi0455), .Z(new_n6149_));
  XOR2_X1    g03630(.A1(new_n6148_), .A2(new_n6149_), .Z(new_n6150_));
  XOR2_X1    g03631(.A1(new_n6150_), .A2(new_n6130_), .Z(new_n6151_));
  NAND2_X1   g03632(.A1(new_n6151_), .A2(pi1196), .ZN(new_n6152_));
  NOR2_X1    g03633(.A1(pi0350), .A2(pi0592), .ZN(new_n6153_));
  AOI21_X1   g03634(.A1(new_n6082_), .A2(new_n6153_), .B(new_n6126_), .ZN(new_n6154_));
  INV_X1     g03635(.I(pi1198), .ZN(new_n6156_));
  XOR2_X1    g03636(.A1(pi0452), .A2(pi0455), .Z(new_n6160_));
  XNOR2_X1   g03637(.A1(pi0357), .A2(pi0461), .ZN(new_n6180_));
  INV_X1     g03638(.I(pi0351), .ZN(new_n6181_));
  NOR2_X1    g03639(.A1(new_n6181_), .A2(pi1199), .ZN(new_n6182_));
  INV_X1     g03640(.I(pi0354), .ZN(new_n6192_));
  INV_X1     g03641(.I(pi0462), .ZN(new_n6193_));
  XOR2_X1    g03642(.A1(pi0352), .A2(pi0353), .Z(new_n6194_));
  XOR2_X1    g03643(.A1(new_n6194_), .A2(new_n6193_), .Z(new_n6195_));
  XOR2_X1    g03644(.A1(new_n6195_), .A2(pi0360), .Z(new_n6196_));
  XOR2_X1    g03645(.A1(new_n6196_), .A2(new_n6192_), .Z(new_n6197_));
  INV_X1     g03646(.I(pi0356), .ZN(new_n6198_));
  NOR3_X1    g03647(.A1(new_n6070_), .A2(pi0590), .A3(new_n5940_), .ZN(new_n6202_));
  INV_X1     g03648(.I(pi0590), .ZN(new_n6203_));
  INV_X1     g03649(.I(pi0334), .ZN(new_n6204_));
  INV_X1     g03650(.I(pi0393), .ZN(new_n6205_));
  XNOR2_X1   g03651(.A1(pi0391), .A2(pi0392), .ZN(new_n6206_));
  INV_X1     g03652(.I(new_n6206_), .ZN(new_n6207_));
  NOR2_X1    g03653(.A1(new_n6090_), .A2(pi0333), .ZN(new_n6208_));
  INV_X1     g03654(.I(pi1196), .ZN(new_n6209_));
  INV_X1     g03655(.I(pi0411), .ZN(new_n6210_));
  INV_X1     g03656(.I(pi0397), .ZN(new_n6211_));
  INV_X1     g03657(.I(pi0319), .ZN(new_n6212_));
  INV_X1     g03658(.I(pi0324), .ZN(new_n6213_));
  NOR2_X1    g03659(.A1(new_n6213_), .A2(pi0456), .ZN(new_n6214_));
  INV_X1     g03660(.I(pi0456), .ZN(new_n6215_));
  NOR2_X1    g03661(.A1(new_n6215_), .A2(pi0324), .ZN(new_n6216_));
  OAI21_X1   g03662(.A1(new_n6214_), .A2(new_n6216_), .B(new_n6212_), .ZN(new_n6217_));
  NOR2_X1    g03663(.A1(pi0324), .A2(pi0456), .ZN(new_n6218_));
  NOR2_X1    g03664(.A1(new_n6213_), .A2(new_n6215_), .ZN(new_n6219_));
  OAI21_X1   g03665(.A1(new_n6219_), .A2(new_n6218_), .B(pi0319), .ZN(new_n6220_));
  NAND2_X1   g03666(.A1(new_n6220_), .A2(new_n6217_), .ZN(new_n6221_));
  XOR2_X1    g03667(.A1(new_n6221_), .A2(new_n6211_), .Z(new_n6222_));
  XOR2_X1    g03668(.A1(new_n6222_), .A2(pi0412), .Z(new_n6223_));
  XOR2_X1    g03669(.A1(new_n6223_), .A2(pi0404), .Z(new_n6224_));
  XOR2_X1    g03670(.A1(pi0390), .A2(pi0410), .Z(new_n6225_));
  INV_X1     g03671(.I(new_n6225_), .ZN(new_n6226_));
  AND2_X2    g03672(.A1(new_n6224_), .A2(new_n6226_), .Z(new_n6227_));
  XNOR2_X1   g03673(.A1(pi0390), .A2(pi0410), .ZN(new_n6228_));
  NOR2_X1    g03674(.A1(new_n6224_), .A2(new_n6228_), .ZN(new_n6229_));
  NOR3_X1    g03675(.A1(new_n6227_), .A2(new_n6210_), .A3(new_n6229_), .ZN(new_n6230_));
  NOR2_X1    g03676(.A1(new_n6227_), .A2(new_n6229_), .ZN(new_n6231_));
  NOR2_X1    g03677(.A1(new_n6231_), .A2(pi0411), .ZN(new_n6232_));
  NOR2_X1    g03678(.A1(new_n6232_), .A2(new_n6230_), .ZN(new_n6233_));
  INV_X1     g03679(.I(new_n6233_), .ZN(new_n6234_));
  NAND4_X1   g03680(.A1(new_n6060_), .A2(new_n6079_), .A3(new_n6064_), .A4(new_n6234_), .ZN(new_n6235_));
  INV_X1     g03681(.I(new_n6072_), .ZN(new_n6236_));
  NOR3_X1    g03682(.A1(new_n6002_), .A2(new_n6236_), .A3(new_n6003_), .ZN(new_n6237_));
  INV_X1     g03683(.I(new_n6006_), .ZN(new_n6238_));
  OAI21_X1   g03684(.A1(new_n6233_), .A2(new_n6238_), .B(new_n6003_), .ZN(new_n6239_));
  NAND2_X1   g03685(.A1(new_n6239_), .A2(new_n6237_), .ZN(new_n6240_));
  NOR2_X1    g03686(.A1(pi0075), .A2(pi0592), .ZN(new_n6241_));
  NAND4_X1   g03687(.A1(new_n6235_), .A2(pi1196), .A3(new_n6240_), .A4(new_n6241_), .ZN(new_n6242_));
  NAND2_X1   g03688(.A1(new_n6242_), .A2(new_n6088_), .ZN(new_n6243_));
  AOI21_X1   g03689(.A1(new_n6067_), .A2(new_n6209_), .B(new_n6243_), .ZN(new_n6244_));
  XNOR2_X1   g03690(.A1(pi0325), .A2(pi0326), .ZN(new_n6245_));
  XOR2_X1    g03691(.A1(new_n6245_), .A2(pi0405), .Z(new_n6246_));
  XOR2_X1    g03692(.A1(new_n6246_), .A2(pi0403), .Z(new_n6247_));
  XOR2_X1    g03693(.A1(new_n6247_), .A2(pi0401), .Z(new_n6248_));
  XOR2_X1    g03694(.A1(new_n6248_), .A2(pi0406), .Z(new_n6249_));
  XOR2_X1    g03695(.A1(new_n6249_), .A2(pi0402), .Z(new_n6250_));
  INV_X1     g03696(.I(new_n6250_), .ZN(new_n6251_));
  XOR2_X1    g03697(.A1(pi0318), .A2(pi0409), .Z(new_n6252_));
  NOR2_X1    g03698(.A1(new_n6251_), .A2(new_n6252_), .ZN(new_n6253_));
  XNOR2_X1   g03699(.A1(pi0318), .A2(pi0409), .ZN(new_n6254_));
  NOR2_X1    g03700(.A1(new_n6250_), .A2(new_n6254_), .ZN(new_n6255_));
  NOR2_X1    g03701(.A1(new_n6253_), .A2(new_n6255_), .ZN(new_n6256_));
  OAI21_X1   g03702(.A1(new_n6234_), .A2(pi0075), .B(new_n6209_), .ZN(new_n6257_));
  NAND2_X1   g03703(.A1(new_n6257_), .A2(new_n6256_), .ZN(new_n6258_));
  NAND4_X1   g03704(.A1(new_n6060_), .A2(new_n6079_), .A3(new_n6064_), .A4(new_n6258_), .ZN(new_n6259_));
  INV_X1     g03705(.I(new_n6256_), .ZN(new_n6260_));
  NOR4_X1    g03706(.A1(new_n6260_), .A2(new_n6003_), .A3(new_n6238_), .A4(new_n6237_), .ZN(new_n6261_));
  INV_X1     g03707(.I(new_n6241_), .ZN(new_n6262_));
  NOR2_X1    g03708(.A1(new_n6262_), .A2(new_n6088_), .ZN(new_n6263_));
  NOR4_X1    g03709(.A1(new_n6261_), .A2(new_n6209_), .A3(new_n6239_), .A4(new_n6263_), .ZN(new_n6264_));
  AOI21_X1   g03710(.A1(new_n6259_), .A2(new_n6264_), .B(pi0567), .ZN(new_n6265_));
  OAI21_X1   g03711(.A1(new_n6068_), .A2(new_n6241_), .B(new_n6265_), .ZN(new_n6266_));
  INV_X1     g03712(.I(pi0567), .ZN(new_n6267_));
  NAND3_X1   g03713(.A1(new_n5981_), .A2(new_n6267_), .A3(new_n5941_), .ZN(new_n6268_));
  XNOR2_X1   g03714(.A1(pi0328), .A2(pi0394), .ZN(new_n6269_));
  XOR2_X1    g03715(.A1(new_n6269_), .A2(pi0408), .Z(new_n6270_));
  XOR2_X1    g03716(.A1(new_n6270_), .A2(pi0396), .Z(new_n6271_));
  XNOR2_X1   g03717(.A1(pi0329), .A2(pi0395), .ZN(new_n6272_));
  XOR2_X1    g03718(.A1(new_n6272_), .A2(pi0399), .Z(new_n6273_));
  XOR2_X1    g03719(.A1(new_n6273_), .A2(pi0398), .Z(new_n6274_));
  XNOR2_X1   g03720(.A1(new_n6274_), .A2(pi0400), .ZN(new_n6275_));
  XOR2_X1    g03721(.A1(new_n6274_), .A2(pi0400), .Z(new_n6276_));
  MUX2_X1    g03722(.I0(new_n6276_), .I1(new_n6275_), .S(new_n6271_), .Z(new_n6277_));
  INV_X1     g03723(.I(new_n6277_), .ZN(new_n6278_));
  NOR2_X1    g03724(.A1(new_n6278_), .A2(new_n6156_), .ZN(new_n6279_));
  NOR2_X1    g03725(.A1(new_n6268_), .A2(new_n6279_), .ZN(new_n6280_));
  OAI21_X1   g03726(.A1(new_n6266_), .A2(new_n6244_), .B(new_n6280_), .ZN(new_n6281_));
  NAND2_X1   g03727(.A1(new_n6087_), .A2(new_n6279_), .ZN(new_n6282_));
  XOR2_X1    g03728(.A1(new_n6281_), .A2(new_n6282_), .Z(new_n6283_));
  MUX2_X1    g03729(.I0(new_n6283_), .I1(new_n6086_), .S(new_n6208_), .Z(new_n6284_));
  NOR2_X1    g03730(.A1(new_n6284_), .A2(new_n6207_), .ZN(new_n6285_));
  INV_X1     g03731(.I(pi0333), .ZN(new_n6286_));
  NOR2_X1    g03732(.A1(new_n6286_), .A2(pi1197), .ZN(new_n6287_));
  MUX2_X1    g03733(.I0(new_n6283_), .I1(new_n6087_), .S(new_n6287_), .Z(new_n6288_));
  NAND2_X1   g03734(.A1(new_n6288_), .A2(new_n6207_), .ZN(new_n6289_));
  XOR2_X1    g03735(.A1(new_n6285_), .A2(new_n6289_), .Z(new_n6290_));
  NAND2_X1   g03736(.A1(new_n6290_), .A2(new_n6205_), .ZN(new_n6291_));
  NOR2_X1    g03737(.A1(new_n6288_), .A2(new_n6207_), .ZN(new_n6292_));
  NAND2_X1   g03738(.A1(new_n6284_), .A2(new_n6207_), .ZN(new_n6293_));
  XNOR2_X1   g03739(.A1(new_n6292_), .A2(new_n6293_), .ZN(new_n6294_));
  OR2_X2     g03740(.A1(new_n6294_), .A2(new_n6205_), .Z(new_n6295_));
  NAND2_X1   g03741(.A1(new_n6295_), .A2(new_n6291_), .ZN(new_n6296_));
  INV_X1     g03742(.I(new_n6296_), .ZN(new_n6297_));
  NOR2_X1    g03743(.A1(new_n6294_), .A2(pi0393), .ZN(new_n6298_));
  AOI21_X1   g03744(.A1(pi0393), .A2(new_n6290_), .B(new_n6298_), .ZN(new_n6299_));
  AOI21_X1   g03745(.A1(new_n6204_), .A2(new_n6299_), .B(new_n6297_), .ZN(new_n6300_));
  NOR3_X1    g03746(.A1(new_n6296_), .A2(new_n6299_), .A3(pi0334), .ZN(new_n6301_));
  XNOR2_X1   g03747(.A1(pi0335), .A2(pi0407), .ZN(new_n6302_));
  XOR2_X1    g03748(.A1(new_n6302_), .A2(pi0463), .Z(new_n6303_));
  XOR2_X1    g03749(.A1(new_n6303_), .A2(pi0413), .Z(new_n6304_));
  NAND4_X1   g03750(.A1(new_n6297_), .A2(new_n6299_), .A3(pi0334), .A4(new_n6304_), .ZN(new_n6305_));
  NAND2_X1   g03751(.A1(new_n6305_), .A2(new_n6304_), .ZN(new_n6306_));
  NOR3_X1    g03752(.A1(new_n6306_), .A2(new_n6300_), .A3(new_n6301_), .ZN(new_n6307_));
  OAI21_X1   g03753(.A1(new_n6307_), .A2(pi0591), .B(new_n6203_), .ZN(new_n6308_));
  NOR2_X1    g03754(.A1(new_n6082_), .A2(new_n6084_), .ZN(new_n6309_));
  AOI21_X1   g03755(.A1(new_n6084_), .A2(new_n6069_), .B(new_n6309_), .ZN(new_n6310_));
  INV_X1     g03756(.I(new_n6310_), .ZN(new_n6311_));
  XOR2_X1    g03757(.A1(pi0365), .A2(pi0447), .Z(new_n6312_));
  INV_X1     g03758(.I(new_n6312_), .ZN(new_n6313_));
  INV_X1     g03759(.I(pi0383), .ZN(new_n6314_));
  XOR2_X1    g03760(.A1(pi0336), .A2(pi0364), .Z(new_n6315_));
  XOR2_X1    g03761(.A1(new_n6315_), .A2(new_n6314_), .Z(new_n6316_));
  XOR2_X1    g03762(.A1(new_n6316_), .A2(pi0366), .Z(new_n6317_));
  XOR2_X1    g03763(.A1(new_n6317_), .A2(new_n6313_), .Z(new_n6318_));
  INV_X1     g03764(.I(pi0389), .ZN(new_n6319_));
  NOR2_X1    g03765(.A1(new_n6319_), .A2(pi0368), .ZN(new_n6320_));
  INV_X1     g03766(.I(pi0368), .ZN(new_n6321_));
  NOR2_X1    g03767(.A1(new_n6321_), .A2(pi0389), .ZN(new_n6322_));
  NOR2_X1    g03768(.A1(new_n6320_), .A2(new_n6322_), .ZN(new_n6323_));
  XOR2_X1    g03769(.A1(new_n6318_), .A2(new_n6323_), .Z(new_n6324_));
  XOR2_X1    g03770(.A1(new_n6324_), .A2(pi0367), .Z(new_n6325_));
  NAND2_X1   g03771(.A1(new_n6325_), .A2(new_n6090_), .ZN(new_n6326_));
  INV_X1     g03772(.I(new_n6326_), .ZN(new_n6327_));
  NOR2_X1    g03773(.A1(new_n6327_), .A2(pi1196), .ZN(new_n6328_));
  OAI21_X1   g03774(.A1(new_n6070_), .A2(new_n6328_), .B(new_n6311_), .ZN(new_n6329_));
  XOR2_X1    g03775(.A1(pi0372), .A2(pi0386), .Z(new_n6330_));
  INV_X1     g03776(.I(pi0372), .ZN(new_n6331_));
  NOR2_X1    g03777(.A1(new_n6331_), .A2(pi0386), .ZN(new_n6332_));
  INV_X1     g03778(.I(pi0386), .ZN(new_n6333_));
  NOR2_X1    g03779(.A1(new_n6333_), .A2(pi0372), .ZN(new_n6334_));
  OAI21_X1   g03780(.A1(new_n6332_), .A2(new_n6334_), .B(pi0363), .ZN(new_n6335_));
  OAI21_X1   g03781(.A1(pi0363), .A2(new_n6330_), .B(new_n6335_), .ZN(new_n6336_));
  INV_X1     g03782(.I(pi0387), .ZN(new_n6337_));
  XOR2_X1    g03783(.A1(pi0337), .A2(pi0339), .Z(new_n6338_));
  XOR2_X1    g03784(.A1(new_n6338_), .A2(new_n6337_), .Z(new_n6339_));
  XOR2_X1    g03785(.A1(new_n6339_), .A2(pi0380), .Z(new_n6340_));
  XOR2_X1    g03786(.A1(new_n6340_), .A2(new_n6336_), .Z(new_n6341_));
  XOR2_X1    g03787(.A1(new_n6341_), .A2(pi0388), .Z(new_n6342_));
  XOR2_X1    g03788(.A1(new_n6342_), .A2(pi0338), .Z(new_n6343_));
  INV_X1     g03789(.I(new_n6343_), .ZN(new_n6344_));
  NOR3_X1    g03790(.A1(new_n6311_), .A2(new_n6069_), .A3(new_n6328_), .ZN(new_n6345_));
  NOR2_X1    g03791(.A1(new_n6345_), .A2(new_n6344_), .ZN(new_n6346_));
  AOI21_X1   g03792(.A1(new_n6070_), .A2(new_n6326_), .B(new_n6343_), .ZN(new_n6347_));
  OAI21_X1   g03793(.A1(new_n6311_), .A2(new_n6326_), .B(new_n6347_), .ZN(new_n6348_));
  NAND2_X1   g03794(.A1(new_n6348_), .A2(new_n6088_), .ZN(new_n6349_));
  AOI21_X1   g03795(.A1(new_n6329_), .A2(new_n6346_), .B(new_n6349_), .ZN(new_n6350_));
  NOR2_X1    g03796(.A1(new_n6344_), .A2(new_n6209_), .ZN(new_n6351_));
  NOR2_X1    g03797(.A1(new_n6351_), .A2(new_n6327_), .ZN(new_n6352_));
  INV_X1     g03798(.I(new_n6352_), .ZN(new_n6353_));
  INV_X1     g03799(.I(pi0377), .ZN(new_n6354_));
  INV_X1     g03800(.I(pi0376), .ZN(new_n6355_));
  INV_X1     g03801(.I(pi0317), .ZN(new_n6356_));
  NOR2_X1    g03802(.A1(pi0378), .A2(pi0385), .ZN(new_n6357_));
  INV_X1     g03803(.I(pi0378), .ZN(new_n6358_));
  INV_X1     g03804(.I(pi0385), .ZN(new_n6359_));
  NOR2_X1    g03805(.A1(new_n6358_), .A2(new_n6359_), .ZN(new_n6360_));
  OAI21_X1   g03806(.A1(new_n6360_), .A2(new_n6357_), .B(new_n6356_), .ZN(new_n6361_));
  NOR2_X1    g03807(.A1(new_n6358_), .A2(pi0385), .ZN(new_n6362_));
  NOR2_X1    g03808(.A1(new_n6359_), .A2(pi0378), .ZN(new_n6363_));
  OAI21_X1   g03809(.A1(new_n6362_), .A2(new_n6363_), .B(pi0317), .ZN(new_n6364_));
  NAND2_X1   g03810(.A1(new_n6361_), .A2(new_n6364_), .ZN(new_n6365_));
  XOR2_X1    g03811(.A1(new_n6365_), .A2(new_n6355_), .Z(new_n6366_));
  XOR2_X1    g03812(.A1(new_n6366_), .A2(pi0439), .Z(new_n6367_));
  XOR2_X1    g03813(.A1(new_n6367_), .A2(pi0381), .Z(new_n6368_));
  XOR2_X1    g03814(.A1(pi0379), .A2(pi0382), .Z(new_n6369_));
  INV_X1     g03815(.I(new_n6369_), .ZN(new_n6370_));
  XNOR2_X1   g03816(.A1(pi0379), .A2(pi0382), .ZN(new_n6371_));
  NOR2_X1    g03817(.A1(new_n6368_), .A2(new_n6371_), .ZN(new_n6372_));
  AOI21_X1   g03818(.A1(new_n6368_), .A2(new_n6370_), .B(new_n6372_), .ZN(new_n6373_));
  NAND2_X1   g03819(.A1(new_n6373_), .A2(new_n6084_), .ZN(new_n6374_));
  AOI21_X1   g03820(.A1(new_n6082_), .A2(new_n6354_), .B(new_n6374_), .ZN(new_n6375_));
  OAI21_X1   g03821(.A1(pi0377), .A2(new_n6084_), .B(new_n6070_), .ZN(new_n6376_));
  NOR2_X1    g03822(.A1(new_n6354_), .A2(new_n6084_), .ZN(new_n6377_));
  INV_X1     g03823(.I(new_n6377_), .ZN(new_n6378_));
  OAI21_X1   g03824(.A1(new_n6111_), .A2(new_n6378_), .B(new_n6373_), .ZN(new_n6379_));
  NAND2_X1   g03825(.A1(new_n6070_), .A2(new_n6378_), .ZN(new_n6380_));
  AOI22_X1   g03826(.A1(new_n6379_), .A2(new_n6380_), .B1(new_n6375_), .B2(new_n6376_), .ZN(new_n6381_));
  MUX2_X1    g03827(.I0(new_n6381_), .I1(new_n6310_), .S(new_n6353_), .Z(new_n6382_));
  NOR2_X1    g03828(.A1(new_n6382_), .A2(new_n6088_), .ZN(new_n6383_));
  OR2_X2     g03829(.A1(new_n6350_), .A2(new_n6383_), .Z(new_n6384_));
  NOR2_X1    g03830(.A1(new_n6383_), .A2(pi1198), .ZN(new_n6385_));
  NOR2_X1    g03831(.A1(new_n6310_), .A2(new_n6156_), .ZN(new_n6386_));
  XOR2_X1    g03832(.A1(new_n6385_), .A2(new_n6386_), .Z(new_n6387_));
  AOI21_X1   g03833(.A1(new_n6156_), .A2(new_n6350_), .B(new_n6387_), .ZN(new_n6388_));
  XNOR2_X1   g03834(.A1(pi0369), .A2(pi0374), .ZN(new_n6389_));
  MUX2_X1    g03835(.I0(new_n6388_), .I1(new_n6384_), .S(new_n6389_), .Z(new_n6390_));
  XNOR2_X1   g03836(.A1(pi0369), .A2(pi0374), .ZN(new_n6391_));
  XNOR2_X1   g03837(.A1(pi0370), .A2(pi0371), .ZN(new_n6392_));
  NOR2_X1    g03838(.A1(new_n6391_), .A2(new_n6392_), .ZN(new_n6393_));
  XOR2_X1    g03839(.A1(new_n6390_), .A2(new_n6393_), .Z(new_n6394_));
  NOR2_X1    g03840(.A1(new_n6394_), .A2(pi0373), .ZN(new_n6395_));
  INV_X1     g03841(.I(pi0373), .ZN(new_n6396_));
  INV_X1     g03842(.I(new_n6392_), .ZN(new_n6397_));
  NAND2_X1   g03843(.A1(new_n6397_), .A2(new_n6391_), .ZN(new_n6398_));
  XNOR2_X1   g03844(.A1(new_n6390_), .A2(new_n6398_), .ZN(new_n6399_));
  NOR2_X1    g03845(.A1(new_n6399_), .A2(new_n6396_), .ZN(new_n6400_));
  XNOR2_X1   g03846(.A1(pi0370), .A2(pi0371), .ZN(new_n6401_));
  OAI22_X1   g03847(.A1(new_n6400_), .A2(new_n6395_), .B1(pi0375), .B2(new_n6401_), .ZN(new_n6402_));
  NOR2_X1    g03848(.A1(new_n6400_), .A2(new_n6395_), .ZN(new_n6403_));
  NOR2_X1    g03849(.A1(new_n6401_), .A2(pi0375), .ZN(new_n6404_));
  NAND2_X1   g03850(.A1(new_n6403_), .A2(new_n6404_), .ZN(new_n6405_));
  NOR2_X1    g03851(.A1(new_n6399_), .A2(pi0373), .ZN(new_n6406_));
  NOR2_X1    g03852(.A1(new_n6394_), .A2(new_n6396_), .ZN(new_n6407_));
  NOR2_X1    g03853(.A1(new_n6406_), .A2(new_n6407_), .ZN(new_n6408_));
  INV_X1     g03854(.I(pi0384), .ZN(new_n6409_));
  INV_X1     g03855(.I(pi0440), .ZN(new_n6410_));
  NOR2_X1    g03856(.A1(new_n6410_), .A2(pi0442), .ZN(new_n6411_));
  INV_X1     g03857(.I(pi0442), .ZN(new_n6412_));
  NOR2_X1    g03858(.A1(new_n6412_), .A2(pi0440), .ZN(new_n6413_));
  OAI21_X1   g03859(.A1(new_n6411_), .A2(new_n6413_), .B(new_n6409_), .ZN(new_n6414_));
  NOR2_X1    g03860(.A1(pi0440), .A2(pi0442), .ZN(new_n6415_));
  NOR2_X1    g03861(.A1(new_n6410_), .A2(new_n6412_), .ZN(new_n6416_));
  OAI21_X1   g03862(.A1(new_n6416_), .A2(new_n6415_), .B(pi0384), .ZN(new_n6417_));
  NAND2_X1   g03863(.A1(new_n6417_), .A2(new_n6414_), .ZN(new_n6418_));
  INV_X1     g03864(.I(new_n6418_), .ZN(new_n6419_));
  NAND4_X1   g03865(.A1(new_n6403_), .A2(new_n6408_), .A3(pi0375), .A4(new_n6419_), .ZN(new_n6420_));
  NOR2_X1    g03866(.A1(new_n6418_), .A2(pi0591), .ZN(new_n6421_));
  NAND4_X1   g03867(.A1(new_n6420_), .A2(new_n6402_), .A3(new_n6405_), .A4(new_n6421_), .ZN(new_n6422_));
  AOI21_X1   g03868(.A1(new_n6422_), .A2(new_n6308_), .B(new_n6202_), .ZN(new_n6423_));
  NOR2_X1    g03869(.A1(new_n2924_), .A2(pi0122), .ZN(new_n6424_));
  INV_X1     g03870(.I(new_n6424_), .ZN(new_n6425_));
  NOR2_X1    g03871(.A1(new_n6005_), .A2(new_n6425_), .ZN(new_n6426_));
  INV_X1     g03872(.I(new_n6426_), .ZN(new_n6427_));
  NOR2_X1    g03873(.A1(new_n6427_), .A2(pi1091), .ZN(new_n6428_));
  INV_X1     g03874(.I(new_n6428_), .ZN(new_n6429_));
  NOR2_X1    g03875(.A1(new_n6429_), .A2(pi0098), .ZN(new_n6430_));
  INV_X1     g03876(.I(new_n6430_), .ZN(new_n6431_));
  NOR2_X1    g03877(.A1(new_n6431_), .A2(new_n6267_), .ZN(new_n6432_));
  NOR2_X1    g03878(.A1(new_n6432_), .A2(new_n5941_), .ZN(new_n6433_));
  INV_X1     g03879(.I(new_n5991_), .ZN(new_n6434_));
  INV_X1     g03880(.I(new_n5994_), .ZN(new_n6435_));
  INV_X1     g03881(.I(new_n6010_), .ZN(new_n6436_));
  NOR4_X1    g03882(.A1(new_n6011_), .A2(pi1091), .A3(new_n6435_), .A4(new_n6436_), .ZN(new_n6437_));
  OR2_X2     g03883(.A1(new_n6437_), .A2(new_n6434_), .Z(new_n6438_));
  NOR2_X1    g03884(.A1(new_n6005_), .A2(pi0098), .ZN(new_n6440_));
  INV_X1     g03885(.I(new_n6440_), .ZN(new_n6441_));
  NOR2_X1    g03886(.A1(new_n6441_), .A2(new_n6425_), .ZN(new_n6442_));
  INV_X1     g03887(.I(new_n5094_), .ZN(new_n6445_));
  INV_X1     g03888(.I(new_n5130_), .ZN(new_n6446_));
  INV_X1     g03889(.I(new_n6442_), .ZN(new_n6448_));
  NOR2_X1    g03890(.A1(new_n5357_), .A2(pi0216), .ZN(new_n6452_));
  INV_X1     g03891(.I(new_n6452_), .ZN(new_n6453_));
  INV_X1     g03892(.I(new_n5141_), .ZN(new_n6460_));
  NOR2_X1    g03893(.A1(new_n4879_), .A2(pi0223), .ZN(new_n6462_));
  NOR2_X1    g03894(.A1(new_n6040_), .A2(new_n5978_), .ZN(new_n6467_));
  NOR2_X1    g03895(.A1(new_n6467_), .A2(pi0039), .ZN(new_n6468_));
  INV_X1     g03896(.I(new_n6032_), .ZN(new_n6469_));
  NAND2_X1   g03897(.A1(new_n6469_), .A2(pi0122), .ZN(new_n6470_));
  NAND2_X1   g03898(.A1(new_n6441_), .A2(new_n6029_), .ZN(new_n6471_));
  NAND4_X1   g03899(.A1(new_n6042_), .A2(pi1093), .A3(new_n6470_), .A4(new_n6471_), .ZN(new_n6472_));
  NOR2_X1    g03900(.A1(new_n6468_), .A2(new_n6472_), .ZN(new_n6473_));
  MUX2_X1    g03901(.I0(new_n6441_), .I1(new_n6238_), .S(pi0122), .Z(new_n6475_));
  NAND4_X1   g03902(.A1(new_n6075_), .A2(pi1093), .A3(new_n3198_), .A4(new_n6073_), .ZN(new_n6476_));
  NOR2_X1    g03903(.A1(new_n6476_), .A2(new_n6475_), .ZN(new_n6477_));
  INV_X1     g03904(.I(new_n6477_), .ZN(new_n6478_));
  NOR2_X1    g03905(.A1(new_n5990_), .A2(new_n2523_), .ZN(new_n6481_));
  NOR2_X1    g03906(.A1(new_n6448_), .A2(pi1091), .ZN(new_n6482_));
  AOI21_X1   g03907(.A1(new_n5981_), .A2(new_n6267_), .B(new_n5942_), .ZN(new_n6488_));
  AND2_X2    g03908(.A1(new_n6488_), .A2(new_n6433_), .Z(new_n6489_));
  NOR2_X1    g03909(.A1(new_n6488_), .A2(new_n6433_), .ZN(new_n6490_));
  NOR2_X1    g03910(.A1(new_n6489_), .A2(new_n6490_), .ZN(new_n6491_));
  INV_X1     g03911(.I(new_n6491_), .ZN(new_n6492_));
  INV_X1     g03912(.I(new_n6089_), .ZN(new_n6493_));
  NOR2_X1    g03913(.A1(new_n6491_), .A2(new_n6084_), .ZN(new_n6494_));
  NOR2_X1    g03914(.A1(new_n6111_), .A2(pi0592), .ZN(new_n6495_));
  NOR2_X1    g03915(.A1(new_n6495_), .A2(new_n6494_), .ZN(new_n6496_));
  INV_X1     g03916(.I(new_n6496_), .ZN(new_n6497_));
  XOR2_X1    g03917(.A1(new_n6148_), .A2(pi0355), .Z(new_n6498_));
  INV_X1     g03918(.I(new_n6498_), .ZN(new_n6499_));
  INV_X1     g03919(.I(pi0452), .ZN(new_n6500_));
  NOR2_X1    g03920(.A1(new_n6492_), .A2(pi0455), .ZN(new_n6501_));
  AOI21_X1   g03921(.A1(new_n6496_), .A2(pi0455), .B(new_n6501_), .ZN(new_n6502_));
  INV_X1     g03922(.I(pi0455), .ZN(new_n6503_));
  NOR2_X1    g03923(.A1(new_n6492_), .A2(new_n6503_), .ZN(new_n6504_));
  AOI21_X1   g03924(.A1(new_n6496_), .A2(new_n6503_), .B(new_n6504_), .ZN(new_n6505_));
  MUX2_X1    g03925(.I0(new_n6505_), .I1(new_n6502_), .S(new_n6500_), .Z(new_n6506_));
  NAND2_X1   g03926(.A1(new_n6502_), .A2(pi0452), .ZN(new_n6507_));
  NAND3_X1   g03927(.A1(new_n6507_), .A2(new_n6209_), .A3(new_n6499_), .ZN(new_n6508_));
  AOI21_X1   g03928(.A1(new_n6500_), .A2(new_n6505_), .B(new_n6508_), .ZN(new_n6509_));
  OAI21_X1   g03929(.A1(new_n6506_), .A2(new_n6499_), .B(new_n6509_), .ZN(new_n6510_));
  OR2_X2     g03930(.A1(new_n6154_), .A2(new_n6153_), .Z(new_n6511_));
  INV_X1     g03931(.I(new_n6152_), .ZN(new_n6512_));
  NOR2_X1    g03932(.A1(new_n6512_), .A2(new_n6109_), .ZN(new_n6513_));
  NAND4_X1   g03933(.A1(new_n6511_), .A2(new_n6127_), .A3(new_n6492_), .A4(new_n6513_), .ZN(new_n6514_));
  NAND4_X1   g03934(.A1(new_n6514_), .A2(new_n6156_), .A3(new_n6152_), .A4(new_n6496_), .ZN(new_n6515_));
  NOR2_X1    g03935(.A1(new_n6491_), .A2(pi1196), .ZN(new_n6516_));
  INV_X1     g03936(.I(new_n6516_), .ZN(new_n6517_));
  NAND4_X1   g03937(.A1(new_n6510_), .A2(new_n6156_), .A3(new_n6515_), .A4(new_n6517_), .ZN(new_n6518_));
  MUX2_X1    g03938(.I0(new_n6518_), .I1(new_n6496_), .S(new_n6107_), .Z(new_n6519_));
  MUX2_X1    g03939(.I0(new_n6519_), .I1(new_n6497_), .S(new_n6493_), .Z(new_n6520_));
  NOR2_X1    g03940(.A1(new_n6181_), .A2(new_n6088_), .ZN(new_n6521_));
  INV_X1     g03941(.I(new_n6521_), .ZN(new_n6522_));
  MUX2_X1    g03942(.I0(new_n6519_), .I1(new_n6497_), .S(new_n6522_), .Z(new_n6523_));
  XOR2_X1    g03943(.A1(new_n6523_), .A2(new_n6520_), .Z(new_n6524_));
  INV_X1     g03944(.I(new_n6524_), .ZN(new_n6525_));
  NOR2_X1    g03945(.A1(new_n6525_), .A2(new_n6180_), .ZN(new_n6526_));
  XNOR2_X1   g03946(.A1(new_n6526_), .A2(new_n6520_), .ZN(new_n6527_));
  NOR2_X1    g03947(.A1(new_n6524_), .A2(new_n6180_), .ZN(new_n6528_));
  XOR2_X1    g03948(.A1(new_n6528_), .A2(new_n6520_), .Z(new_n6529_));
  NOR2_X1    g03949(.A1(new_n6529_), .A2(new_n6198_), .ZN(new_n6530_));
  AOI21_X1   g03950(.A1(new_n6198_), .A2(new_n6527_), .B(new_n6530_), .ZN(new_n6531_));
  NOR2_X1    g03951(.A1(new_n6529_), .A2(pi0356), .ZN(new_n6532_));
  AOI21_X1   g03952(.A1(pi0356), .A2(new_n6527_), .B(new_n6532_), .ZN(new_n6533_));
  MUX2_X1    g03953(.I0(new_n6533_), .I1(new_n6531_), .S(new_n6197_), .Z(new_n6534_));
  NAND4_X1   g03954(.A1(new_n6534_), .A2(new_n6203_), .A3(new_n5940_), .A4(new_n6492_), .ZN(new_n6535_));
  INV_X1     g03955(.I(pi0288), .ZN(new_n6536_));
  NOR3_X1    g03956(.A1(pi0285), .A2(pi0286), .A3(pi0289), .ZN(new_n6537_));
  NAND2_X1   g03957(.A1(new_n6537_), .A2(new_n6536_), .ZN(new_n6538_));
  INV_X1     g03958(.I(new_n6279_), .ZN(new_n6539_));
  NOR2_X1    g03959(.A1(new_n6234_), .A2(new_n6075_), .ZN(new_n6540_));
  INV_X1     g03960(.I(new_n6482_), .ZN(new_n6541_));
  NOR2_X1    g03961(.A1(new_n6233_), .A2(new_n6541_), .ZN(new_n6542_));
  AOI21_X1   g03962(.A1(new_n6542_), .A2(new_n3198_), .B(new_n3177_), .ZN(new_n6543_));
  OAI21_X1   g03963(.A1(new_n6478_), .A2(new_n6540_), .B(new_n6543_), .ZN(new_n6544_));
  INV_X1     g03964(.I(new_n6542_), .ZN(new_n6545_));
  INV_X1     g03965(.I(new_n6473_), .ZN(new_n6546_));
  AOI21_X1   g03966(.A1(new_n6041_), .A2(new_n6233_), .B(new_n6546_), .ZN(new_n6547_));
  INV_X1     g03967(.I(new_n5143_), .ZN(new_n6548_));
  NOR2_X1    g03968(.A1(new_n6048_), .A2(new_n6548_), .ZN(new_n6549_));
  NOR2_X1    g03969(.A1(new_n6048_), .A2(new_n5130_), .ZN(new_n6551_));
  AOI21_X1   g03970(.A1(new_n6542_), .A2(new_n6453_), .B(new_n2587_), .ZN(new_n6554_));
  INV_X1     g03971(.I(new_n6549_), .ZN(new_n6556_));
  INV_X1     g03972(.I(new_n6551_), .ZN(new_n6558_));
  INV_X1     g03973(.I(new_n6462_), .ZN(new_n6559_));
  NOR3_X1    g03974(.A1(new_n6545_), .A2(new_n3172_), .A3(new_n3173_), .ZN(new_n6565_));
  NOR2_X1    g03975(.A1(new_n6542_), .A2(new_n6016_), .ZN(new_n6566_));
  OAI21_X1   g03976(.A1(new_n6565_), .A2(new_n6566_), .B(new_n3177_), .ZN(new_n6567_));
  AOI21_X1   g03977(.A1(new_n6567_), .A2(new_n6544_), .B(pi0075), .ZN(new_n6568_));
  NAND2_X1   g03978(.A1(new_n6234_), .A2(new_n6442_), .ZN(new_n6569_));
  AOI21_X1   g03979(.A1(new_n6569_), .A2(new_n2918_), .B(new_n6438_), .ZN(new_n6570_));
  NOR4_X1    g03980(.A1(new_n6570_), .A2(pi0075), .A3(new_n6434_), .A4(new_n6542_), .ZN(new_n6571_));
  NOR2_X1    g03981(.A1(new_n6209_), .A2(pi0592), .ZN(new_n6572_));
  INV_X1     g03982(.I(new_n6572_), .ZN(new_n6573_));
  NOR3_X1    g03983(.A1(new_n6545_), .A2(new_n6267_), .A3(new_n5941_), .ZN(new_n6574_));
  OAI21_X1   g03984(.A1(new_n6574_), .A2(new_n6573_), .B(pi0567), .ZN(new_n6575_));
  NOR2_X1    g03985(.A1(new_n6571_), .A2(new_n6575_), .ZN(new_n6576_));
  NAND2_X1   g03986(.A1(new_n6576_), .A2(new_n6268_), .ZN(new_n6577_));
  OAI21_X1   g03987(.A1(new_n6577_), .A2(new_n6568_), .B(new_n6088_), .ZN(new_n6578_));
  OAI21_X1   g03988(.A1(new_n6516_), .A2(new_n6578_), .B(new_n6539_), .ZN(new_n6579_));
  NOR2_X1    g03989(.A1(new_n6260_), .A2(new_n6541_), .ZN(new_n6580_));
  NOR2_X1    g03990(.A1(new_n5941_), .A2(new_n6267_), .ZN(new_n6581_));
  NAND2_X1   g03991(.A1(new_n6084_), .A2(new_n6209_), .ZN(new_n6582_));
  AOI21_X1   g03992(.A1(new_n6580_), .A2(new_n6581_), .B(new_n6582_), .ZN(new_n6583_));
  OAI21_X1   g03993(.A1(new_n6256_), .A2(new_n6075_), .B(new_n6477_), .ZN(new_n6584_));
  NAND4_X1   g03994(.A1(new_n6580_), .A2(new_n3177_), .A3(new_n3198_), .A4(new_n6584_), .ZN(new_n6585_));
  INV_X1     g03995(.I(new_n6580_), .ZN(new_n6586_));
  OAI21_X1   g03996(.A1(new_n6586_), .A2(new_n6452_), .B(pi0299), .ZN(new_n6591_));
  NOR2_X1    g03997(.A1(new_n6586_), .A2(new_n6462_), .ZN(new_n6592_));
  NOR2_X1    g03998(.A1(pi0039), .A2(pi0299), .ZN(new_n6593_));
  INV_X1     g03999(.I(new_n6593_), .ZN(new_n6594_));
  OAI21_X1   g04000(.A1(new_n6260_), .A2(new_n6469_), .B(pi0122), .ZN(new_n6598_));
  OAI21_X1   g04001(.A1(new_n6260_), .A2(new_n6441_), .B(new_n6029_), .ZN(new_n6599_));
  NAND2_X1   g04002(.A1(new_n6598_), .A2(new_n6599_), .ZN(new_n6600_));
  NAND3_X1   g04003(.A1(new_n6600_), .A2(new_n2924_), .A3(new_n6042_), .ZN(new_n6601_));
  NOR3_X1    g04004(.A1(new_n6586_), .A2(new_n3172_), .A3(new_n3173_), .ZN(new_n6603_));
  NOR2_X1    g04005(.A1(new_n6580_), .A2(new_n6016_), .ZN(new_n6604_));
  OAI21_X1   g04006(.A1(new_n6603_), .A2(new_n6604_), .B(new_n3177_), .ZN(new_n6605_));
  AOI21_X1   g04007(.A1(new_n6605_), .A2(new_n6585_), .B(pi0075), .ZN(new_n6606_));
  NAND2_X1   g04008(.A1(new_n6256_), .A2(new_n6442_), .ZN(new_n6607_));
  AOI21_X1   g04009(.A1(new_n6607_), .A2(new_n2918_), .B(new_n6438_), .ZN(new_n6608_));
  NOR4_X1    g04010(.A1(new_n6608_), .A2(pi0075), .A3(new_n6580_), .A4(new_n6434_), .ZN(new_n6609_));
  OAI21_X1   g04011(.A1(new_n6606_), .A2(new_n6609_), .B(new_n6583_), .ZN(new_n6610_));
  NOR2_X1    g04012(.A1(new_n6260_), .A2(new_n6545_), .ZN(new_n6611_));
  NAND2_X1   g04013(.A1(new_n6611_), .A2(new_n5401_), .ZN(new_n6619_));
  INV_X1     g04014(.I(new_n6611_), .ZN(new_n6620_));
  NAND2_X1   g04015(.A1(new_n6620_), .A2(new_n6558_), .ZN(new_n6621_));
  NAND2_X1   g04016(.A1(new_n6621_), .A2(new_n6460_), .ZN(new_n6622_));
  NAND2_X1   g04017(.A1(new_n6620_), .A2(new_n6556_), .ZN(new_n6623_));
  AOI21_X1   g04018(.A1(new_n6623_), .A2(new_n5141_), .B(new_n6462_), .ZN(new_n6624_));
  NAND2_X1   g04019(.A1(new_n6592_), .A2(new_n6542_), .ZN(new_n6625_));
  NAND2_X1   g04020(.A1(new_n6625_), .A2(new_n2587_), .ZN(new_n6626_));
  AOI21_X1   g04021(.A1(new_n6622_), .A2(new_n6624_), .B(new_n6626_), .ZN(new_n6627_));
  INV_X1     g04022(.I(new_n6554_), .ZN(new_n6628_));
  NAND2_X1   g04023(.A1(new_n6621_), .A2(new_n6445_), .ZN(new_n6629_));
  AOI21_X1   g04024(.A1(new_n6623_), .A2(new_n5094_), .B(new_n6452_), .ZN(new_n6630_));
  AOI22_X1   g04025(.A1(new_n6630_), .A2(new_n6629_), .B1(new_n6628_), .B2(new_n6591_), .ZN(new_n6631_));
  OAI21_X1   g04026(.A1(new_n6627_), .A2(new_n3154_), .B(new_n6631_), .ZN(new_n6632_));
  NAND2_X1   g04027(.A1(new_n6547_), .A2(new_n6601_), .ZN(new_n6633_));
  AOI21_X1   g04028(.A1(new_n6633_), .A2(new_n6632_), .B(pi0038), .ZN(new_n6634_));
  NOR3_X1    g04029(.A1(new_n6586_), .A2(new_n3172_), .A3(new_n6545_), .ZN(new_n6635_));
  OR3_X2     g04030(.A1(new_n6634_), .A2(pi0100), .A3(new_n6635_), .Z(new_n6636_));
  NOR4_X1    g04031(.A1(new_n6586_), .A2(pi0087), .A3(new_n3197_), .A4(new_n6545_), .ZN(new_n6637_));
  NOR2_X1    g04032(.A1(new_n6584_), .A2(new_n6540_), .ZN(new_n6638_));
  OAI21_X1   g04033(.A1(new_n6637_), .A2(new_n6638_), .B(new_n3177_), .ZN(new_n6639_));
  AOI21_X1   g04034(.A1(new_n6636_), .A2(new_n6619_), .B(new_n6639_), .ZN(new_n6640_));
  AOI21_X1   g04035(.A1(new_n6620_), .A2(new_n2918_), .B(new_n6438_), .ZN(new_n6641_));
  NOR2_X1    g04036(.A1(new_n6545_), .A2(new_n6267_), .ZN(new_n6642_));
  NOR2_X1    g04037(.A1(new_n5941_), .A2(new_n6572_), .ZN(new_n6643_));
  NAND4_X1   g04038(.A1(new_n6642_), .A2(new_n6256_), .A3(new_n6440_), .A4(new_n6643_), .ZN(new_n6644_));
  NAND4_X1   g04039(.A1(new_n6580_), .A2(new_n2628_), .A3(new_n6434_), .A4(new_n6542_), .ZN(new_n6645_));
  NAND2_X1   g04040(.A1(new_n6645_), .A2(new_n6644_), .ZN(new_n6646_));
  NOR2_X1    g04041(.A1(new_n6646_), .A2(new_n6641_), .ZN(new_n6647_));
  OAI21_X1   g04042(.A1(new_n6640_), .A2(pi0075), .B(new_n6647_), .ZN(new_n6648_));
  INV_X1     g04043(.I(new_n6583_), .ZN(new_n6649_));
  AOI21_X1   g04044(.A1(new_n6649_), .A2(new_n6644_), .B(pi1199), .ZN(new_n6650_));
  AOI21_X1   g04045(.A1(new_n6650_), .A2(new_n6268_), .B(new_n6267_), .ZN(new_n6651_));
  NAND4_X1   g04046(.A1(new_n6648_), .A2(new_n6579_), .A3(new_n6610_), .A4(new_n6651_), .ZN(new_n6652_));
  AOI21_X1   g04047(.A1(new_n6495_), .A2(new_n6279_), .B(new_n6494_), .ZN(new_n6653_));
  NAND2_X1   g04048(.A1(new_n6652_), .A2(new_n6653_), .ZN(new_n6654_));
  XOR2_X1    g04049(.A1(new_n6654_), .A2(new_n6497_), .Z(new_n6655_));
  NAND2_X1   g04050(.A1(new_n6655_), .A2(new_n6208_), .ZN(new_n6656_));
  XOR2_X1    g04051(.A1(new_n6656_), .A2(new_n6496_), .Z(new_n6657_));
  NAND3_X1   g04052(.A1(new_n6655_), .A2(pi0333), .A3(pi1197), .ZN(new_n6658_));
  XOR2_X1    g04053(.A1(new_n6658_), .A2(new_n6496_), .Z(new_n6659_));
  AOI21_X1   g04054(.A1(new_n6659_), .A2(new_n6207_), .B(new_n6657_), .ZN(new_n6660_));
  XOR2_X1    g04055(.A1(new_n6304_), .A2(new_n6204_), .Z(new_n6661_));
  XOR2_X1    g04056(.A1(new_n6661_), .A2(new_n6205_), .Z(new_n6662_));
  INV_X1     g04057(.I(new_n6657_), .ZN(new_n6663_));
  NOR3_X1    g04058(.A1(new_n6663_), .A2(new_n6206_), .A3(new_n6659_), .ZN(new_n6664_));
  NOR3_X1    g04059(.A1(new_n6664_), .A2(new_n6660_), .A3(new_n6662_), .ZN(new_n6665_));
  XOR2_X1    g04060(.A1(new_n6658_), .A2(new_n6497_), .Z(new_n6666_));
  AOI21_X1   g04061(.A1(new_n6666_), .A2(new_n6207_), .B(new_n6657_), .ZN(new_n6667_));
  NAND3_X1   g04062(.A1(new_n6659_), .A2(new_n6657_), .A3(new_n6207_), .ZN(new_n6668_));
  NAND2_X1   g04063(.A1(new_n6668_), .A2(new_n6662_), .ZN(new_n6669_));
  OAI21_X1   g04064(.A1(new_n6669_), .A2(new_n6667_), .B(pi0591), .ZN(new_n6670_));
  OAI21_X1   g04065(.A1(new_n6670_), .A2(new_n6665_), .B(new_n6203_), .ZN(new_n6671_));
  INV_X1     g04066(.I(pi0371), .ZN(new_n6672_));
  INV_X1     g04067(.I(new_n6309_), .ZN(new_n6673_));
  OAI21_X1   g04068(.A1(pi0592), .A2(new_n6492_), .B(new_n6673_), .ZN(new_n6674_));
  NOR2_X1    g04069(.A1(new_n6379_), .A2(new_n6378_), .ZN(new_n6675_));
  NOR2_X1    g04070(.A1(new_n6084_), .A2(pi0377), .ZN(new_n6676_));
  OAI21_X1   g04071(.A1(new_n6675_), .A2(new_n6676_), .B(new_n6491_), .ZN(new_n6677_));
  NOR2_X1    g04072(.A1(new_n6677_), .A2(new_n6353_), .ZN(new_n6678_));
  NOR2_X1    g04073(.A1(new_n6492_), .A2(new_n6353_), .ZN(new_n6679_));
  OAI21_X1   g04074(.A1(pi1199), .A2(new_n6679_), .B(new_n6678_), .ZN(new_n6680_));
  NAND2_X1   g04075(.A1(new_n6674_), .A2(new_n6353_), .ZN(new_n6681_));
  NAND4_X1   g04076(.A1(new_n6677_), .A2(new_n6088_), .A3(new_n6352_), .A4(new_n6491_), .ZN(new_n6682_));
  NAND3_X1   g04077(.A1(new_n6680_), .A2(new_n6681_), .A3(new_n6682_), .ZN(new_n6683_));
  XOR2_X1    g04078(.A1(new_n6683_), .A2(new_n6674_), .Z(new_n6684_));
  NAND2_X1   g04079(.A1(pi0374), .A2(pi1198), .ZN(new_n6685_));
  NOR2_X1    g04080(.A1(new_n6684_), .A2(new_n6685_), .ZN(new_n6686_));
  XNOR2_X1   g04081(.A1(new_n6686_), .A2(new_n6674_), .ZN(new_n6687_));
  XNOR2_X1   g04082(.A1(pi0369), .A2(pi0370), .ZN(new_n6688_));
  INV_X1     g04083(.I(pi0374), .ZN(new_n6689_));
  NAND2_X1   g04084(.A1(new_n6689_), .A2(pi1198), .ZN(new_n6690_));
  NOR2_X1    g04085(.A1(new_n6684_), .A2(new_n6690_), .ZN(new_n6691_));
  XOR2_X1    g04086(.A1(new_n6691_), .A2(new_n6674_), .Z(new_n6692_));
  XOR2_X1    g04087(.A1(new_n6687_), .A2(new_n6692_), .Z(new_n6693_));
  NOR2_X1    g04088(.A1(new_n6693_), .A2(new_n6688_), .ZN(new_n6694_));
  XOR2_X1    g04089(.A1(new_n6694_), .A2(new_n6687_), .Z(new_n6695_));
  XOR2_X1    g04090(.A1(pi0373), .A2(pi0375), .Z(new_n6696_));
  NOR2_X1    g04091(.A1(new_n6418_), .A2(new_n6696_), .ZN(new_n6697_));
  XOR2_X1    g04092(.A1(pi0373), .A2(pi0375), .Z(new_n6698_));
  AOI21_X1   g04093(.A1(new_n6418_), .A2(new_n6698_), .B(new_n6697_), .ZN(new_n6699_));
  INV_X1     g04094(.I(new_n6693_), .ZN(new_n6700_));
  NOR2_X1    g04095(.A1(new_n6700_), .A2(new_n6688_), .ZN(new_n6701_));
  AOI21_X1   g04096(.A1(new_n6701_), .A2(new_n6687_), .B(new_n6672_), .ZN(new_n6702_));
  OAI21_X1   g04097(.A1(new_n6687_), .A2(new_n6701_), .B(new_n6702_), .ZN(new_n6703_));
  NAND2_X1   g04098(.A1(new_n6703_), .A2(new_n6699_), .ZN(new_n6704_));
  AOI21_X1   g04099(.A1(new_n6672_), .A2(new_n6695_), .B(new_n6704_), .ZN(new_n6705_));
  NOR2_X1    g04100(.A1(new_n6695_), .A2(new_n6672_), .ZN(new_n6706_));
  NAND3_X1   g04101(.A1(new_n6703_), .A2(new_n5940_), .A3(new_n6699_), .ZN(new_n6707_));
  OR3_X2     g04102(.A1(new_n6705_), .A2(new_n6706_), .A3(new_n6707_), .Z(new_n6708_));
  AOI21_X1   g04103(.A1(new_n6708_), .A2(new_n6671_), .B(new_n6538_), .ZN(new_n6709_));
  AOI21_X1   g04104(.A1(new_n6709_), .A2(new_n6535_), .B(pi0588), .ZN(new_n6710_));
  INV_X1     g04105(.I(pi0588), .ZN(new_n6711_));
  XNOR2_X1   g04106(.A1(pi0426), .A2(pi0430), .ZN(new_n6712_));
  INV_X1     g04107(.I(pi0454), .ZN(new_n6713_));
  INV_X1     g04108(.I(pi0459), .ZN(new_n6714_));
  XOR2_X1    g04109(.A1(pi0421), .A2(pi0432), .Z(new_n6715_));
  XOR2_X1    g04110(.A1(new_n6715_), .A2(new_n6714_), .Z(new_n6716_));
  XOR2_X1    g04111(.A1(new_n6716_), .A2(new_n6713_), .Z(new_n6717_));
  XOR2_X1    g04112(.A1(pi0419), .A2(pi0420), .Z(new_n6718_));
  XOR2_X1    g04113(.A1(new_n6718_), .A2(pi0424), .Z(new_n6719_));
  XOR2_X1    g04114(.A1(new_n6719_), .A2(pi0423), .Z(new_n6720_));
  XOR2_X1    g04115(.A1(new_n6717_), .A2(new_n6720_), .Z(new_n6721_));
  XOR2_X1    g04116(.A1(new_n6721_), .A2(pi0425), .Z(new_n6722_));
  NAND2_X1   g04117(.A1(new_n6722_), .A2(new_n6156_), .ZN(new_n6723_));
  INV_X1     g04118(.I(pi0417), .ZN(new_n6724_));
  INV_X1     g04119(.I(pi0418), .ZN(new_n6725_));
  NOR2_X1    g04120(.A1(new_n6725_), .A2(pi0437), .ZN(new_n6726_));
  INV_X1     g04121(.I(pi0437), .ZN(new_n6727_));
  NOR2_X1    g04122(.A1(new_n6727_), .A2(pi0418), .ZN(new_n6728_));
  OAI21_X1   g04123(.A1(new_n6726_), .A2(new_n6728_), .B(new_n6724_), .ZN(new_n6729_));
  NOR2_X1    g04124(.A1(pi0418), .A2(pi0437), .ZN(new_n6730_));
  NOR2_X1    g04125(.A1(new_n6725_), .A2(new_n6727_), .ZN(new_n6731_));
  OAI21_X1   g04126(.A1(new_n6731_), .A2(new_n6730_), .B(pi0417), .ZN(new_n6732_));
  NAND2_X1   g04127(.A1(new_n6732_), .A2(new_n6729_), .ZN(new_n6733_));
  XOR2_X1    g04128(.A1(pi0453), .A2(pi0464), .Z(new_n6734_));
  XOR2_X1    g04129(.A1(pi0453), .A2(pi0464), .Z(new_n6735_));
  NAND2_X1   g04130(.A1(new_n6733_), .A2(new_n6735_), .ZN(new_n6736_));
  OAI21_X1   g04131(.A1(new_n6733_), .A2(new_n6734_), .B(new_n6736_), .ZN(new_n6737_));
  XOR2_X1    g04132(.A1(pi0415), .A2(pi0416), .Z(new_n6738_));
  XOR2_X1    g04133(.A1(new_n6738_), .A2(pi0438), .Z(new_n6739_));
  XOR2_X1    g04134(.A1(new_n6739_), .A2(pi0431), .Z(new_n6740_));
  XOR2_X1    g04135(.A1(new_n6740_), .A2(new_n6737_), .Z(new_n6741_));
  NAND2_X1   g04136(.A1(new_n6741_), .A2(new_n6090_), .ZN(new_n6742_));
  NAND2_X1   g04137(.A1(new_n6723_), .A2(new_n6742_), .ZN(new_n6743_));
  NOR2_X1    g04138(.A1(new_n6496_), .A2(new_n6743_), .ZN(new_n6744_));
  INV_X1     g04139(.I(pi0443), .ZN(new_n6745_));
  NOR2_X1    g04140(.A1(new_n6745_), .A2(pi0592), .ZN(new_n6746_));
  XNOR2_X1   g04141(.A1(pi0414), .A2(pi0422), .ZN(new_n6747_));
  XOR2_X1    g04142(.A1(new_n6747_), .A2(pi0446), .Z(new_n6748_));
  NOR2_X1    g04143(.A1(new_n6748_), .A2(pi0434), .ZN(new_n6749_));
  AND2_X2    g04144(.A1(new_n6748_), .A2(pi0434), .Z(new_n6750_));
  NOR2_X1    g04145(.A1(new_n6750_), .A2(new_n6749_), .ZN(new_n6751_));
  XOR2_X1    g04146(.A1(pi0429), .A2(pi0435), .Z(new_n6752_));
  NAND2_X1   g04147(.A1(new_n6751_), .A2(new_n6752_), .ZN(new_n6753_));
  XOR2_X1    g04148(.A1(pi0429), .A2(pi0435), .Z(new_n6754_));
  OAI21_X1   g04149(.A1(new_n6751_), .A2(new_n6754_), .B(new_n6753_), .ZN(new_n6755_));
  XOR2_X1    g04150(.A1(pi0436), .A2(pi0444), .Z(new_n6756_));
  XOR2_X1    g04151(.A1(new_n6755_), .A2(new_n6756_), .Z(new_n6757_));
  AOI21_X1   g04152(.A1(new_n6082_), .A2(new_n6746_), .B(new_n6757_), .ZN(new_n6758_));
  NOR4_X1    g04153(.A1(new_n6758_), .A2(pi1196), .A3(new_n6491_), .A4(new_n6746_), .ZN(new_n6759_));
  NAND2_X1   g04154(.A1(new_n6745_), .A2(new_n6084_), .ZN(new_n6760_));
  OAI21_X1   g04155(.A1(new_n6111_), .A2(new_n6760_), .B(new_n6757_), .ZN(new_n6761_));
  NAND3_X1   g04156(.A1(new_n6761_), .A2(new_n6492_), .A3(new_n6760_), .ZN(new_n6762_));
  OAI21_X1   g04157(.A1(new_n6762_), .A2(new_n6759_), .B(new_n6517_), .ZN(new_n6763_));
  NAND2_X1   g04158(.A1(new_n6763_), .A2(new_n6743_), .ZN(new_n6764_));
  XNOR2_X1   g04159(.A1(new_n6764_), .A2(new_n6744_), .ZN(new_n6765_));
  XNOR2_X1   g04160(.A1(pi0427), .A2(pi0428), .ZN(new_n6766_));
  MUX2_X1    g04161(.I0(new_n6497_), .I1(new_n6765_), .S(new_n6766_), .Z(new_n6767_));
  INV_X1     g04162(.I(new_n6765_), .ZN(new_n6768_));
  MUX2_X1    g04163(.I0(new_n6497_), .I1(new_n6768_), .S(new_n6766_), .Z(new_n6769_));
  MUX2_X1    g04164(.I0(new_n6769_), .I1(new_n6767_), .S(new_n6712_), .Z(new_n6770_));
  NOR2_X1    g04165(.A1(new_n6770_), .A2(pi0445), .ZN(new_n6771_));
  INV_X1     g04166(.I(pi0445), .ZN(new_n6772_));
  INV_X1     g04167(.I(new_n6712_), .ZN(new_n6773_));
  NOR2_X1    g04168(.A1(new_n6769_), .A2(new_n6773_), .ZN(new_n6774_));
  NOR2_X1    g04169(.A1(new_n6767_), .A2(new_n6712_), .ZN(new_n6775_));
  XOR2_X1    g04170(.A1(new_n6774_), .A2(new_n6775_), .Z(new_n6776_));
  NOR2_X1    g04171(.A1(new_n6776_), .A2(new_n6772_), .ZN(new_n6777_));
  NOR2_X1    g04172(.A1(new_n6776_), .A2(pi0445), .ZN(new_n6778_));
  NOR2_X1    g04173(.A1(new_n6770_), .A2(new_n6772_), .ZN(new_n6779_));
  NOR2_X1    g04174(.A1(new_n6778_), .A2(new_n6779_), .ZN(new_n6780_));
  INV_X1     g04175(.I(pi0448), .ZN(new_n6781_));
  INV_X1     g04176(.I(pi0433), .ZN(new_n6782_));
  NOR2_X1    g04177(.A1(pi0449), .A2(pi0451), .ZN(new_n6783_));
  INV_X1     g04178(.I(pi0449), .ZN(new_n6784_));
  INV_X1     g04179(.I(pi0451), .ZN(new_n6785_));
  NOR2_X1    g04180(.A1(new_n6784_), .A2(new_n6785_), .ZN(new_n6786_));
  OAI21_X1   g04181(.A1(new_n6786_), .A2(new_n6783_), .B(new_n6782_), .ZN(new_n6787_));
  NOR2_X1    g04182(.A1(new_n6784_), .A2(pi0451), .ZN(new_n6788_));
  NOR2_X1    g04183(.A1(new_n6785_), .A2(pi0449), .ZN(new_n6789_));
  OAI21_X1   g04184(.A1(new_n6788_), .A2(new_n6789_), .B(pi0433), .ZN(new_n6790_));
  NAND2_X1   g04185(.A1(new_n6787_), .A2(new_n6790_), .ZN(new_n6791_));
  XOR2_X1    g04186(.A1(new_n6791_), .A2(new_n6781_), .Z(new_n6792_));
  OAI22_X1   g04187(.A1(new_n6780_), .A2(new_n6792_), .B1(new_n6771_), .B2(new_n6777_), .ZN(new_n6793_));
  NOR2_X1    g04188(.A1(new_n6777_), .A2(new_n6771_), .ZN(new_n6794_));
  INV_X1     g04189(.I(new_n6792_), .ZN(new_n6795_));
  NAND3_X1   g04190(.A1(new_n6780_), .A2(new_n6794_), .A3(new_n6795_), .ZN(new_n6796_));
  NOR2_X1    g04191(.A1(pi0590), .A2(pi0591), .ZN(new_n6797_));
  INV_X1     g04192(.I(new_n6797_), .ZN(new_n6798_));
  AOI21_X1   g04193(.A1(new_n6765_), .A2(new_n6088_), .B(new_n6798_), .ZN(new_n6799_));
  AOI21_X1   g04194(.A1(new_n6491_), .A2(new_n6798_), .B(new_n6538_), .ZN(new_n6800_));
  NOR3_X1    g04195(.A1(new_n6799_), .A2(new_n6088_), .A3(new_n6800_), .ZN(new_n6801_));
  NAND3_X1   g04196(.A1(new_n6793_), .A2(new_n6796_), .A3(new_n6801_), .ZN(new_n6802_));
  INV_X1     g04197(.I(new_n6743_), .ZN(new_n6803_));
  INV_X1     g04198(.I(pi0444), .ZN(new_n6804_));
  NAND2_X1   g04199(.A1(new_n6111_), .A2(new_n6746_), .ZN(new_n6805_));
  OAI21_X1   g04200(.A1(new_n6070_), .A2(new_n6746_), .B(new_n6805_), .ZN(new_n6806_));
  NAND2_X1   g04201(.A1(new_n6806_), .A2(new_n6804_), .ZN(new_n6807_));
  NAND2_X1   g04202(.A1(new_n6069_), .A2(new_n6760_), .ZN(new_n6808_));
  OAI21_X1   g04203(.A1(new_n6082_), .A2(new_n6760_), .B(new_n6808_), .ZN(new_n6809_));
  NAND2_X1   g04204(.A1(new_n6809_), .A2(pi0444), .ZN(new_n6810_));
  NAND2_X1   g04205(.A1(new_n6807_), .A2(new_n6810_), .ZN(new_n6811_));
  NAND2_X1   g04206(.A1(new_n6806_), .A2(pi0444), .ZN(new_n6812_));
  INV_X1     g04207(.I(pi0436), .ZN(new_n6813_));
  AOI21_X1   g04208(.A1(new_n6809_), .A2(new_n6804_), .B(new_n6813_), .ZN(new_n6814_));
  AOI21_X1   g04209(.A1(new_n6812_), .A2(new_n6814_), .B(new_n6755_), .ZN(new_n6815_));
  OAI21_X1   g04210(.A1(pi0436), .A2(new_n6811_), .B(new_n6815_), .ZN(new_n6816_));
  NAND2_X1   g04211(.A1(new_n6812_), .A2(new_n6814_), .ZN(new_n6817_));
  NAND2_X1   g04212(.A1(new_n6811_), .A2(pi0436), .ZN(new_n6818_));
  NAND2_X1   g04213(.A1(new_n6818_), .A2(new_n6817_), .ZN(new_n6819_));
  AOI21_X1   g04214(.A1(new_n6819_), .A2(new_n6755_), .B(new_n6209_), .ZN(new_n6820_));
  AOI22_X1   g04215(.A1(new_n6820_), .A2(new_n6816_), .B1(new_n6209_), .B2(new_n6070_), .ZN(new_n6821_));
  MUX2_X1    g04216(.I0(new_n6821_), .I1(new_n6087_), .S(new_n6803_), .Z(new_n6822_));
  MUX2_X1    g04217(.I0(new_n6822_), .I1(new_n6086_), .S(new_n6766_), .Z(new_n6823_));
  INV_X1     g04218(.I(new_n6766_), .ZN(new_n6824_));
  NOR2_X1    g04219(.A1(new_n6822_), .A2(new_n6824_), .ZN(new_n6825_));
  NOR2_X1    g04220(.A1(new_n6086_), .A2(new_n6766_), .ZN(new_n6826_));
  XOR2_X1    g04221(.A1(new_n6825_), .A2(new_n6826_), .Z(new_n6827_));
  XNOR2_X1   g04222(.A1(new_n6827_), .A2(new_n6823_), .ZN(new_n6828_));
  NOR2_X1    g04223(.A1(new_n6828_), .A2(new_n6712_), .ZN(new_n6829_));
  XOR2_X1    g04224(.A1(new_n6829_), .A2(new_n6823_), .Z(new_n6830_));
  NOR2_X1    g04225(.A1(new_n6712_), .A2(pi0445), .ZN(new_n6831_));
  NOR2_X1    g04226(.A1(new_n6830_), .A2(new_n6831_), .ZN(new_n6832_));
  AND2_X2    g04227(.A1(new_n6830_), .A2(new_n6831_), .Z(new_n6833_));
  XOR2_X1    g04228(.A1(new_n6791_), .A2(new_n6781_), .Z(new_n6834_));
  INV_X1     g04229(.I(new_n6830_), .ZN(new_n6835_));
  NAND2_X1   g04230(.A1(new_n6828_), .A2(new_n6773_), .ZN(new_n6836_));
  XOR2_X1    g04231(.A1(new_n6836_), .A2(new_n6823_), .Z(new_n6837_));
  NOR4_X1    g04232(.A1(new_n6835_), .A2(new_n6837_), .A3(new_n6772_), .A4(new_n6834_), .ZN(new_n6838_));
  NOR4_X1    g04233(.A1(new_n6838_), .A2(new_n6832_), .A3(new_n6833_), .A4(new_n6834_), .ZN(new_n6839_));
  OAI21_X1   g04234(.A1(new_n6822_), .A2(new_n6798_), .B(new_n6088_), .ZN(new_n6840_));
  NOR3_X1    g04235(.A1(new_n6070_), .A2(new_n6797_), .A3(new_n6538_), .ZN(new_n6841_));
  OAI21_X1   g04236(.A1(new_n6839_), .A2(new_n6840_), .B(new_n6841_), .ZN(new_n6842_));
  AOI21_X1   g04237(.A1(new_n6842_), .A2(new_n6802_), .B(new_n6711_), .ZN(new_n6843_));
  INV_X1     g04238(.I(new_n6538_), .ZN(new_n6844_));
  NOR2_X1    g04239(.A1(new_n5223_), .A2(pi0057), .ZN(new_n6845_));
  NAND2_X1   g04240(.A1(new_n6845_), .A2(new_n6844_), .ZN(new_n6846_));
  NOR4_X1    g04241(.A1(new_n6710_), .A2(new_n6423_), .A3(new_n6843_), .A4(new_n6846_), .ZN(new_n6847_));
  NAND3_X1   g04242(.A1(new_n6492_), .A2(new_n6069_), .A3(new_n6844_), .ZN(new_n6848_));
  OAI21_X1   g04243(.A1(new_n6492_), .A2(new_n6538_), .B(new_n6070_), .ZN(new_n6849_));
  NAND3_X1   g04244(.A1(new_n6849_), .A2(new_n6848_), .A3(new_n6845_), .ZN(new_n6850_));
  INV_X1     g04245(.I(new_n6432_), .ZN(new_n6851_));
  NOR2_X1    g04246(.A1(new_n6851_), .A2(new_n6084_), .ZN(new_n6852_));
  INV_X1     g04247(.I(new_n6852_), .ZN(new_n6853_));
  NAND2_X1   g04248(.A1(new_n6233_), .A2(pi1196), .ZN(new_n6854_));
  NAND4_X1   g04249(.A1(new_n6580_), .A2(pi0567), .A3(new_n6084_), .A4(new_n6854_), .ZN(new_n6855_));
  NAND2_X1   g04250(.A1(new_n6855_), .A2(new_n6853_), .ZN(new_n6856_));
  NAND2_X1   g04251(.A1(new_n6856_), .A2(new_n6088_), .ZN(new_n6857_));
  NAND2_X1   g04252(.A1(new_n6642_), .A2(new_n6572_), .ZN(new_n6858_));
  NAND2_X1   g04253(.A1(new_n6851_), .A2(new_n6572_), .ZN(new_n6859_));
  NAND4_X1   g04254(.A1(new_n6857_), .A2(new_n6088_), .A3(new_n6858_), .A4(new_n6859_), .ZN(new_n6860_));
  NOR2_X1    g04255(.A1(new_n6853_), .A2(new_n6090_), .ZN(new_n6861_));
  AOI21_X1   g04256(.A1(new_n6860_), .A2(new_n6090_), .B(new_n6861_), .ZN(new_n6862_));
  NOR3_X1    g04257(.A1(new_n6860_), .A2(new_n6156_), .A3(new_n6852_), .ZN(new_n6863_));
  NOR2_X1    g04258(.A1(new_n6863_), .A2(new_n6278_), .ZN(new_n6864_));
  OAI21_X1   g04259(.A1(pi0333), .A2(new_n6860_), .B(new_n6864_), .ZN(new_n6865_));
  AOI21_X1   g04260(.A1(pi0333), .A2(new_n6862_), .B(new_n6865_), .ZN(new_n6866_));
  NAND2_X1   g04261(.A1(new_n6864_), .A2(new_n6860_), .ZN(new_n6867_));
  AOI21_X1   g04262(.A1(new_n6286_), .A2(new_n6862_), .B(new_n6867_), .ZN(new_n6868_));
  XOR2_X1    g04263(.A1(new_n6866_), .A2(new_n6868_), .Z(new_n6869_));
  NAND2_X1   g04264(.A1(new_n6869_), .A2(new_n6207_), .ZN(new_n6870_));
  XOR2_X1    g04265(.A1(new_n6870_), .A2(new_n6866_), .Z(new_n6871_));
  NAND2_X1   g04266(.A1(new_n6662_), .A2(new_n6206_), .ZN(new_n6872_));
  XOR2_X1    g04267(.A1(new_n6871_), .A2(new_n6872_), .Z(new_n6873_));
  OAI21_X1   g04268(.A1(new_n6873_), .A2(pi0590), .B(new_n6851_), .ZN(new_n6874_));
  NAND3_X1   g04269(.A1(new_n6873_), .A2(new_n6203_), .A3(new_n6432_), .ZN(new_n6875_));
  AOI21_X1   g04270(.A1(new_n6874_), .A2(new_n6875_), .B(new_n5940_), .ZN(new_n6876_));
  XOR2_X1    g04271(.A1(new_n6126_), .A2(new_n6108_), .Z(new_n6877_));
  NOR2_X1    g04272(.A1(new_n6877_), .A2(new_n6512_), .ZN(new_n6878_));
  NOR2_X1    g04273(.A1(new_n6851_), .A2(pi0592), .ZN(new_n6879_));
  NAND3_X1   g04274(.A1(new_n6878_), .A2(pi1198), .A3(new_n6879_), .ZN(new_n6880_));
  XOR2_X1    g04275(.A1(new_n6149_), .A2(pi0355), .Z(new_n6881_));
  XOR2_X1    g04276(.A1(new_n6881_), .A2(pi0458), .Z(new_n6882_));
  XOR2_X1    g04277(.A1(new_n6882_), .A2(pi0361), .Z(new_n6883_));
  XOR2_X1    g04278(.A1(new_n6883_), .A2(pi0441), .Z(new_n6884_));
  NAND2_X1   g04279(.A1(new_n6432_), .A2(new_n6141_), .ZN(new_n6885_));
  AOI21_X1   g04280(.A1(new_n6884_), .A2(new_n6084_), .B(new_n6885_), .ZN(new_n6886_));
  XNOR2_X1   g04281(.A1(new_n6148_), .A2(new_n6881_), .ZN(new_n6887_));
  NAND2_X1   g04282(.A1(new_n6887_), .A2(new_n6084_), .ZN(new_n6888_));
  NAND4_X1   g04283(.A1(new_n6888_), .A2(new_n6209_), .A3(new_n6144_), .A4(new_n6432_), .ZN(new_n6889_));
  OAI21_X1   g04284(.A1(new_n6889_), .A2(new_n6886_), .B(new_n6156_), .ZN(new_n6890_));
  AOI21_X1   g04285(.A1(new_n6880_), .A2(new_n6890_), .B(new_n6107_), .ZN(new_n6891_));
  OR3_X2     g04286(.A1(new_n6891_), .A2(pi0592), .A3(new_n6851_), .Z(new_n6892_));
  NAND2_X1   g04287(.A1(new_n6892_), .A2(new_n6521_), .ZN(new_n6893_));
  XOR2_X1    g04288(.A1(new_n6893_), .A2(new_n6853_), .Z(new_n6894_));
  NAND2_X1   g04289(.A1(new_n6892_), .A2(new_n6089_), .ZN(new_n6895_));
  XOR2_X1    g04290(.A1(new_n6895_), .A2(new_n6852_), .Z(new_n6896_));
  XOR2_X1    g04291(.A1(new_n6896_), .A2(new_n6894_), .Z(new_n6897_));
  NOR2_X1    g04292(.A1(new_n6897_), .A2(new_n6180_), .ZN(new_n6898_));
  XOR2_X1    g04293(.A1(new_n6898_), .A2(new_n6894_), .Z(new_n6899_));
  INV_X1     g04294(.I(new_n6897_), .ZN(new_n6900_));
  NOR2_X1    g04295(.A1(new_n6900_), .A2(new_n6180_), .ZN(new_n6901_));
  XNOR2_X1   g04296(.A1(new_n6901_), .A2(new_n6894_), .ZN(new_n6902_));
  XOR2_X1    g04297(.A1(new_n6197_), .A2(pi0356), .Z(new_n6903_));
  OAI21_X1   g04298(.A1(new_n6902_), .A2(new_n6903_), .B(new_n6899_), .ZN(new_n6904_));
  INV_X1     g04299(.I(new_n6902_), .ZN(new_n6905_));
  NOR3_X1    g04300(.A1(new_n6905_), .A2(new_n6899_), .A3(new_n6903_), .ZN(new_n6906_));
  NOR2_X1    g04301(.A1(new_n6906_), .A2(new_n6203_), .ZN(new_n6907_));
  XOR2_X1    g04302(.A1(new_n6373_), .A2(new_n6354_), .Z(new_n6908_));
  NOR2_X1    g04303(.A1(new_n6353_), .A2(new_n6908_), .ZN(new_n6909_));
  INV_X1     g04304(.I(new_n6909_), .ZN(new_n6910_));
  NOR3_X1    g04305(.A1(new_n6432_), .A2(new_n6084_), .A3(pi1199), .ZN(new_n6911_));
  AOI22_X1   g04306(.A1(new_n6910_), .A2(new_n6911_), .B1(pi0592), .B2(new_n6353_), .ZN(new_n6912_));
  NAND2_X1   g04307(.A1(new_n6912_), .A2(new_n6852_), .ZN(new_n6913_));
  XOR2_X1    g04308(.A1(new_n6688_), .A2(pi0374), .Z(new_n6914_));
  XOR2_X1    g04309(.A1(new_n6914_), .A2(pi0371), .Z(new_n6915_));
  XOR2_X1    g04310(.A1(new_n6915_), .A2(new_n6418_), .Z(new_n6916_));
  XOR2_X1    g04311(.A1(new_n6916_), .A2(pi0375), .Z(new_n6917_));
  OAI21_X1   g04312(.A1(new_n6917_), .A2(pi0373), .B(pi1198), .ZN(new_n6918_));
  AOI21_X1   g04313(.A1(pi0373), .A2(new_n6917_), .B(new_n6918_), .ZN(new_n6919_));
  AOI21_X1   g04314(.A1(new_n6913_), .A2(new_n6919_), .B(new_n6879_), .ZN(new_n6920_));
  NAND2_X1   g04315(.A1(new_n6920_), .A2(new_n6203_), .ZN(new_n6921_));
  NAND2_X1   g04316(.A1(new_n6921_), .A2(new_n5940_), .ZN(new_n6922_));
  AOI21_X1   g04317(.A1(new_n6907_), .A2(new_n6904_), .B(new_n6922_), .ZN(new_n6923_));
  INV_X1     g04318(.I(new_n6791_), .ZN(new_n6924_));
  INV_X1     g04319(.I(new_n6879_), .ZN(new_n6925_));
  NAND2_X1   g04320(.A1(new_n6804_), .A2(pi0443), .ZN(new_n6926_));
  NAND2_X1   g04321(.A1(new_n6745_), .A2(pi0444), .ZN(new_n6927_));
  AOI21_X1   g04322(.A1(new_n6926_), .A2(new_n6927_), .B(pi0436), .ZN(new_n6928_));
  XNOR2_X1   g04323(.A1(pi0443), .A2(pi0444), .ZN(new_n6929_));
  AOI21_X1   g04324(.A1(pi0436), .A2(new_n6929_), .B(new_n6928_), .ZN(new_n6930_));
  XNOR2_X1   g04325(.A1(new_n6755_), .A2(new_n6930_), .ZN(new_n6931_));
  NAND3_X1   g04326(.A1(new_n6803_), .A2(new_n6572_), .A3(new_n6931_), .ZN(new_n6932_));
  NOR2_X1    g04327(.A1(new_n6932_), .A2(new_n6925_), .ZN(new_n6933_));
  XNOR2_X1   g04328(.A1(pi0426), .A2(pi0427), .ZN(new_n6934_));
  XOR2_X1    g04329(.A1(new_n6934_), .A2(pi0430), .Z(new_n6935_));
  XOR2_X1    g04330(.A1(new_n6935_), .A2(pi0428), .Z(new_n6936_));
  XOR2_X1    g04331(.A1(new_n6936_), .A2(pi0445), .Z(new_n6937_));
  XOR2_X1    g04332(.A1(new_n6937_), .A2(new_n6781_), .Z(new_n6938_));
  AOI21_X1   g04333(.A1(new_n6933_), .A2(new_n6938_), .B(new_n6852_), .ZN(new_n6939_));
  INV_X1     g04334(.I(new_n6933_), .ZN(new_n6940_));
  AOI21_X1   g04335(.A1(new_n6940_), .A2(new_n6938_), .B(new_n6852_), .ZN(new_n6941_));
  MUX2_X1    g04336(.I0(new_n6941_), .I1(new_n6939_), .S(new_n6924_), .Z(new_n6942_));
  OR2_X2     g04337(.A1(new_n6942_), .A2(new_n6088_), .Z(new_n6943_));
  NOR2_X1    g04338(.A1(new_n6852_), .A2(pi1199), .ZN(new_n6944_));
  OAI21_X1   g04339(.A1(new_n6851_), .A2(new_n6797_), .B(pi0588), .ZN(new_n6945_));
  NAND4_X1   g04340(.A1(new_n6945_), .A2(new_n6797_), .A3(new_n6844_), .A4(new_n6845_), .ZN(new_n6946_));
  AOI21_X1   g04341(.A1(new_n6940_), .A2(new_n6944_), .B(new_n6946_), .ZN(new_n6947_));
  AOI21_X1   g04342(.A1(new_n6943_), .A2(new_n6947_), .B(pi0588), .ZN(new_n6948_));
  OAI21_X1   g04343(.A1(new_n6876_), .A2(new_n6923_), .B(new_n6948_), .ZN(new_n6949_));
  INV_X1     g04344(.I(new_n6845_), .ZN(po1038));
  NAND2_X1   g04345(.A1(po1038), .A2(new_n6844_), .ZN(new_n6951_));
  NOR3_X1    g04346(.A1(new_n6851_), .A2(pi0217), .A3(new_n6951_), .ZN(new_n6952_));
  NOR3_X1    g04347(.A1(pi1161), .A2(pi1162), .A3(pi1163), .ZN(new_n6953_));
  NOR3_X1    g04348(.A1(new_n6952_), .A2(pi0217), .A3(new_n6953_), .ZN(new_n6954_));
  NAND3_X1   g04349(.A1(new_n6949_), .A2(new_n6850_), .A3(new_n6954_), .ZN(new_n6955_));
  INV_X1     g04350(.I(pi1163), .ZN(new_n6956_));
  NAND3_X1   g04351(.A1(new_n2925_), .A2(pi1161), .A3(new_n6956_), .ZN(new_n6957_));
  INV_X1     g04352(.I(pi0031), .ZN(new_n6958_));
  NAND2_X1   g04353(.A1(new_n6958_), .A2(pi1162), .ZN(new_n6959_));
  OAI22_X1   g04354(.A1(new_n6847_), .A2(new_n6955_), .B1(new_n6957_), .B2(new_n6959_), .ZN(po0189));
  NAND2_X1   g04355(.A1(new_n2533_), .A2(new_n2571_), .ZN(new_n6961_));
  NOR2_X1    g04356(.A1(pi0055), .A2(pi0074), .ZN(new_n6962_));
  INV_X1     g04357(.I(new_n6962_), .ZN(new_n6963_));
  NOR2_X1    g04358(.A1(new_n6961_), .A2(new_n6963_), .ZN(new_n6964_));
  INV_X1     g04359(.I(new_n6964_), .ZN(new_n6965_));
  NOR2_X1    g04360(.A1(new_n6965_), .A2(new_n5410_), .ZN(new_n6966_));
  INV_X1     g04361(.I(new_n6966_), .ZN(new_n6967_));
  INV_X1     g04362(.I(new_n2671_), .ZN(new_n6968_));
  NOR2_X1    g04363(.A1(new_n6968_), .A2(pi0024), .ZN(new_n6969_));
  INV_X1     g04364(.I(new_n6969_), .ZN(new_n6970_));
  NOR4_X1    g04365(.A1(new_n6970_), .A2(pi0051), .A3(new_n2485_), .A4(new_n2644_), .ZN(new_n6971_));
  NOR2_X1    g04366(.A1(new_n5177_), .A2(new_n5990_), .ZN(new_n6972_));
  INV_X1     g04367(.I(new_n6972_), .ZN(new_n6973_));
  NAND2_X1   g04368(.A1(new_n6973_), .A2(pi0252), .ZN(new_n6974_));
  INV_X1     g04369(.I(new_n5163_), .ZN(new_n6975_));
  NOR2_X1    g04370(.A1(new_n5177_), .A2(new_n6975_), .ZN(new_n6976_));
  NAND2_X1   g04371(.A1(new_n2924_), .A2(pi0829), .ZN(new_n6977_));
  NOR2_X1    g04372(.A1(new_n6977_), .A2(new_n2955_), .ZN(new_n6978_));
  NOR2_X1    g04373(.A1(new_n2964_), .A2(new_n6978_), .ZN(new_n6979_));
  INV_X1     g04374(.I(new_n6979_), .ZN(po0840));
  NOR2_X1    g04375(.A1(new_n2545_), .A2(pi0087), .ZN(new_n6981_));
  NAND3_X1   g04376(.A1(new_n6981_), .A2(pi0075), .A3(new_n3173_), .ZN(new_n6982_));
  NOR4_X1    g04377(.A1(new_n6976_), .A2(pi0137), .A3(po0840), .A4(new_n6982_), .ZN(new_n6983_));
  NAND3_X1   g04378(.A1(new_n6971_), .A2(new_n6974_), .A3(new_n6983_), .ZN(new_n6984_));
  NOR2_X1    g04379(.A1(new_n2705_), .A2(new_n2460_), .ZN(new_n6985_));
  INV_X1     g04380(.I(new_n2638_), .ZN(new_n6986_));
  NAND3_X1   g04381(.A1(new_n2887_), .A2(new_n2466_), .A3(new_n2468_), .ZN(new_n6987_));
  NOR3_X1    g04382(.A1(new_n6987_), .A2(pi0047), .A3(new_n6986_), .ZN(new_n6988_));
  INV_X1     g04383(.I(new_n2467_), .ZN(new_n6989_));
  NOR2_X1    g04384(.A1(new_n6989_), .A2(pi0093), .ZN(new_n6990_));
  NOR4_X1    g04385(.A1(new_n5083_), .A2(pi0024), .A3(pi0040), .A4(pi0090), .ZN(new_n6991_));
  NAND4_X1   g04386(.A1(new_n6985_), .A2(new_n6988_), .A3(new_n6990_), .A4(new_n6991_), .ZN(new_n6992_));
  OAI21_X1   g04387(.A1(new_n5084_), .A2(new_n6992_), .B(pi0032), .ZN(new_n6993_));
  NOR2_X1    g04388(.A1(new_n6993_), .A2(new_n5080_), .ZN(new_n6994_));
  NOR2_X1    g04389(.A1(pi0024), .A2(pi0841), .ZN(new_n6995_));
  NAND2_X1   g04390(.A1(new_n2655_), .A2(pi0032), .ZN(new_n6996_));
  INV_X1     g04391(.I(new_n6985_), .ZN(new_n6997_));
  NOR2_X1    g04392(.A1(new_n2469_), .A2(new_n2640_), .ZN(new_n6998_));
  INV_X1     g04393(.I(new_n6998_), .ZN(new_n6999_));
  NAND2_X1   g04394(.A1(new_n2799_), .A2(new_n2800_), .ZN(new_n7000_));
  NOR2_X1    g04395(.A1(pi0089), .A2(pi0102), .ZN(new_n7001_));
  NAND2_X1   g04396(.A1(new_n5955_), .A2(new_n7001_), .ZN(new_n7002_));
  NOR4_X1    g04397(.A1(pi0049), .A2(pi0066), .A3(pi0068), .A4(pi0073), .ZN(new_n7003_));
  NOR4_X1    g04398(.A1(new_n7002_), .A2(pi0081), .A3(new_n7000_), .A4(new_n7003_), .ZN(new_n7004_));
  NOR2_X1    g04399(.A1(new_n2724_), .A2(new_n2785_), .ZN(new_n7005_));
  NOR2_X1    g04400(.A1(pi0045), .A2(pi0048), .ZN(new_n7006_));
  NAND4_X1   g04401(.A1(new_n7005_), .A2(new_n2492_), .A3(new_n2747_), .A4(new_n7006_), .ZN(new_n7007_));
  INV_X1     g04402(.I(new_n2463_), .ZN(new_n7008_));
  NOR4_X1    g04403(.A1(new_n2497_), .A2(new_n7008_), .A3(new_n2769_), .A4(pi0103), .ZN(new_n7009_));
  NAND4_X1   g04404(.A1(new_n7009_), .A2(new_n2454_), .A3(pi0076), .A4(new_n2444_), .ZN(new_n7010_));
  NOR2_X1    g04405(.A1(new_n7010_), .A2(new_n7007_), .ZN(new_n7011_));
  NAND2_X1   g04406(.A1(new_n7011_), .A2(new_n7004_), .ZN(new_n7012_));
  AOI21_X1   g04407(.A1(new_n6997_), .A2(new_n7012_), .B(new_n6999_), .ZN(new_n7013_));
  INV_X1     g04408(.I(new_n6988_), .ZN(new_n7014_));
  NOR2_X1    g04409(.A1(new_n7012_), .A2(new_n6989_), .ZN(new_n7015_));
  INV_X1     g04410(.I(new_n7015_), .ZN(new_n7016_));
  NOR2_X1    g04411(.A1(new_n7016_), .A2(new_n7014_), .ZN(new_n7017_));
  INV_X1     g04412(.I(new_n7017_), .ZN(new_n7018_));
  AOI21_X1   g04413(.A1(new_n7013_), .A2(new_n7018_), .B(new_n5895_), .ZN(new_n7019_));
  NOR2_X1    g04414(.A1(po0840), .A2(new_n6538_), .ZN(new_n7020_));
  NOR2_X1    g04415(.A1(new_n2963_), .A2(new_n2505_), .ZN(new_n7021_));
  INV_X1     g04416(.I(new_n7021_), .ZN(new_n7022_));
  NOR4_X1    g04417(.A1(new_n7020_), .A2(pi0137), .A3(new_n5965_), .A4(new_n7022_), .ZN(new_n7023_));
  NOR2_X1    g04418(.A1(new_n7020_), .A2(pi0137), .ZN(new_n7024_));
  NOR2_X1    g04419(.A1(new_n6992_), .A2(new_n7024_), .ZN(new_n7025_));
  AOI21_X1   g04420(.A1(new_n7019_), .A2(new_n7023_), .B(new_n7025_), .ZN(new_n7026_));
  OAI22_X1   g04421(.A1(new_n7026_), .A2(pi0032), .B1(new_n6995_), .B2(new_n6996_), .ZN(new_n7027_));
  AOI21_X1   g04422(.A1(new_n7027_), .A2(new_n5080_), .B(new_n6994_), .ZN(new_n7028_));
  NAND2_X1   g04423(.A1(new_n2546_), .A2(new_n2437_), .ZN(new_n7029_));
  NOR4_X1    g04424(.A1(po1057), .A2(new_n2491_), .A3(new_n6975_), .A4(new_n5186_), .ZN(new_n7030_));
  NAND2_X1   g04425(.A1(new_n7030_), .A2(new_n2436_), .ZN(new_n7031_));
  INV_X1     g04426(.I(new_n3191_), .ZN(new_n7032_));
  NAND2_X1   g04427(.A1(new_n2490_), .A2(pi0129), .ZN(new_n7033_));
  INV_X1     g04428(.I(new_n7033_), .ZN(new_n7034_));
  NOR4_X1    g04429(.A1(new_n6972_), .A2(pi0137), .A3(new_n3181_), .A4(new_n5163_), .ZN(new_n7035_));
  AOI21_X1   g04430(.A1(new_n7035_), .A2(new_n7034_), .B(new_n7032_), .ZN(new_n7036_));
  AOI21_X1   g04431(.A1(new_n7036_), .A2(new_n7031_), .B(new_n2535_), .ZN(new_n7037_));
  OAI21_X1   g04432(.A1(new_n7028_), .A2(new_n7029_), .B(new_n7037_), .ZN(new_n7038_));
  AOI21_X1   g04433(.A1(new_n7038_), .A2(new_n6984_), .B(new_n6967_), .ZN(po0190));
  INV_X1     g04434(.I(pi0954), .ZN(po1110));
  NOR2_X1    g04435(.A1(pi0075), .A2(pi0100), .ZN(new_n7041_));
  XNOR2_X1   g04436(.A1(pi0149), .A2(pi0157), .ZN(new_n7042_));
  NOR2_X1    g04437(.A1(new_n7042_), .A2(new_n5109_), .ZN(new_n7043_));
  INV_X1     g04438(.I(new_n7043_), .ZN(new_n7044_));
  NOR2_X1    g04439(.A1(new_n7044_), .A2(new_n5987_), .ZN(new_n7045_));
  NOR2_X1    g04440(.A1(new_n7045_), .A2(new_n7041_), .ZN(new_n7046_));
  INV_X1     g04441(.I(new_n7046_), .ZN(new_n7047_));
  INV_X1     g04442(.I(new_n7041_), .ZN(new_n7048_));
  NOR2_X1    g04443(.A1(new_n5989_), .A2(new_n7048_), .ZN(new_n7049_));
  INV_X1     g04444(.I(new_n7049_), .ZN(new_n7050_));
  NOR4_X1    g04445(.A1(new_n7047_), .A2(pi0074), .A3(new_n4272_), .A4(new_n7050_), .ZN(new_n7051_));
  AOI21_X1   g04446(.A1(pi0164), .A2(new_n7049_), .B(new_n7046_), .ZN(new_n7052_));
  NOR2_X1    g04447(.A1(new_n7052_), .A2(pi0074), .ZN(new_n7053_));
  OAI21_X1   g04448(.A1(new_n2571_), .A2(new_n7051_), .B(new_n7053_), .ZN(new_n7054_));
  INV_X1     g04449(.I(new_n7051_), .ZN(new_n7055_));
  NOR2_X1    g04450(.A1(new_n7052_), .A2(new_n3214_), .ZN(new_n7056_));
  INV_X1     g04451(.I(new_n7056_), .ZN(new_n7057_));
  INV_X1     g04452(.I(pi0164), .ZN(new_n7058_));
  NOR3_X1    g04453(.A1(new_n5989_), .A2(new_n3172_), .A3(new_n7058_), .ZN(new_n7059_));
  AOI21_X1   g04454(.A1(new_n7041_), .A2(new_n7059_), .B(new_n7046_), .ZN(new_n7060_));
  NAND2_X1   g04455(.A1(new_n7057_), .A2(new_n7060_), .ZN(new_n7061_));
  NAND2_X1   g04456(.A1(new_n7061_), .A2(new_n3202_), .ZN(new_n7062_));
  AOI21_X1   g04457(.A1(new_n7062_), .A2(new_n7055_), .B(new_n2533_), .ZN(new_n7063_));
  NOR2_X1    g04458(.A1(new_n7063_), .A2(new_n3405_), .ZN(new_n7064_));
  AOI21_X1   g04459(.A1(new_n5988_), .A2(pi0164), .B(new_n3172_), .ZN(new_n7065_));
  NOR2_X1    g04460(.A1(new_n7065_), .A2(new_n3206_), .ZN(new_n7066_));
  INV_X1     g04461(.I(pi0149), .ZN(new_n7067_));
  NOR2_X1    g04462(.A1(pi0053), .A2(pi0060), .ZN(new_n7068_));
  NOR2_X1    g04463(.A1(new_n2698_), .A2(pi0050), .ZN(new_n7069_));
  INV_X1     g04464(.I(new_n7069_), .ZN(new_n7070_));
  NOR2_X1    g04465(.A1(pi0064), .A2(pi0081), .ZN(new_n7071_));
  INV_X1     g04466(.I(new_n7071_), .ZN(new_n7072_));
  NOR2_X1    g04467(.A1(new_n7072_), .A2(pi0102), .ZN(new_n7073_));
  INV_X1     g04468(.I(new_n7073_), .ZN(new_n7074_));
  NOR2_X1    g04469(.A1(new_n7074_), .A2(new_n2724_), .ZN(new_n7075_));
  INV_X1     g04470(.I(new_n7075_), .ZN(new_n7076_));
  NOR3_X1    g04471(.A1(new_n2723_), .A2(new_n7070_), .A3(new_n7076_), .ZN(new_n7077_));
  NOR2_X1    g04472(.A1(new_n2888_), .A2(new_n2683_), .ZN(new_n7078_));
  NAND3_X1   g04473(.A1(new_n7077_), .A2(new_n7068_), .A3(new_n7078_), .ZN(new_n7079_));
  NOR2_X1    g04474(.A1(new_n7079_), .A2(pi0058), .ZN(new_n7080_));
  INV_X1     g04475(.I(new_n7080_), .ZN(new_n7081_));
  NOR2_X1    g04476(.A1(new_n7081_), .A2(new_n5965_), .ZN(new_n7082_));
  NAND3_X1   g04477(.A1(new_n7082_), .A2(new_n2632_), .A3(new_n2506_), .ZN(new_n7083_));
  NOR2_X1    g04478(.A1(new_n7083_), .A2(pi0095), .ZN(new_n7084_));
  NOR4_X1    g04479(.A1(new_n7084_), .A2(pi0039), .A3(new_n7067_), .A4(new_n5989_), .ZN(new_n7085_));
  NOR2_X1    g04480(.A1(new_n7000_), .A2(pi0040), .ZN(new_n7086_));
  INV_X1     g04481(.I(new_n7086_), .ZN(new_n7087_));
  OAI21_X1   g04482(.A1(new_n7085_), .A2(new_n7087_), .B(new_n3172_), .ZN(new_n7088_));
  INV_X1     g04483(.I(new_n7045_), .ZN(new_n7089_));
  OAI21_X1   g04484(.A1(new_n7086_), .A2(pi0038), .B(new_n3173_), .ZN(new_n7090_));
  NOR2_X1    g04485(.A1(new_n7065_), .A2(new_n7090_), .ZN(new_n7091_));
  AOI22_X1   g04486(.A1(new_n7089_), .A2(pi0100), .B1(pi0087), .B2(new_n7091_), .ZN(new_n7092_));
  AOI21_X1   g04487(.A1(new_n7088_), .A2(new_n7066_), .B(new_n7092_), .ZN(new_n7093_));
  MUX2_X1    g04488(.I0(new_n7093_), .I1(new_n7045_), .S(pi0075), .Z(new_n7094_));
  NAND2_X1   g04489(.A1(new_n7091_), .A2(new_n2628_), .ZN(new_n7095_));
  NOR2_X1    g04490(.A1(new_n7046_), .A2(new_n3203_), .ZN(new_n7096_));
  AOI22_X1   g04491(.A1(new_n7094_), .A2(new_n3203_), .B1(new_n7095_), .B2(new_n7096_), .ZN(new_n7097_));
  AOI21_X1   g04492(.A1(new_n7052_), .A2(pi0054), .B(pi0074), .ZN(new_n7098_));
  OAI21_X1   g04493(.A1(new_n7097_), .A2(pi0054), .B(new_n7098_), .ZN(new_n7099_));
  NOR2_X1    g04494(.A1(new_n7051_), .A2(new_n3227_), .ZN(new_n7100_));
  XNOR2_X1   g04495(.A1(pi0178), .A2(pi0183), .ZN(new_n7101_));
  NOR2_X1    g04496(.A1(new_n7101_), .A2(new_n5109_), .ZN(new_n7102_));
  MUX2_X1    g04497(.I0(new_n7102_), .I1(new_n7043_), .S(pi0299), .Z(new_n7103_));
  NAND2_X1   g04498(.A1(new_n7103_), .A2(pi0232), .ZN(new_n7104_));
  INV_X1     g04499(.I(new_n7104_), .ZN(new_n7105_));
  NOR2_X1    g04500(.A1(new_n7105_), .A2(new_n3173_), .ZN(new_n7106_));
  NOR2_X1    g04501(.A1(new_n7105_), .A2(new_n2628_), .ZN(new_n7107_));
  NOR2_X1    g04502(.A1(new_n7106_), .A2(new_n7107_), .ZN(new_n7108_));
  INV_X1     g04503(.I(pi0186), .ZN(new_n7109_));
  MUX2_X1    g04504(.I0(new_n7109_), .I1(new_n7058_), .S(pi0299), .Z(new_n7110_));
  NOR2_X1    g04505(.A1(new_n5989_), .A2(new_n7110_), .ZN(new_n7111_));
  INV_X1     g04506(.I(new_n7111_), .ZN(new_n7112_));
  NOR4_X1    g04507(.A1(new_n7108_), .A2(pi0054), .A3(new_n7048_), .A4(new_n7112_), .ZN(new_n7113_));
  AOI21_X1   g04508(.A1(new_n3271_), .A2(pi0299), .B(new_n5987_), .ZN(new_n7114_));
  INV_X1     g04509(.I(new_n7114_), .ZN(new_n7115_));
  NOR2_X1    g04510(.A1(pi0176), .A2(pi0299), .ZN(new_n7116_));
  NOR3_X1    g04511(.A1(new_n7115_), .A2(new_n5109_), .A3(new_n7116_), .ZN(new_n7117_));
  INV_X1     g04512(.I(new_n7084_), .ZN(new_n7118_));
  NOR2_X1    g04513(.A1(new_n7118_), .A2(new_n2624_), .ZN(new_n7119_));
  INV_X1     g04514(.I(new_n7119_), .ZN(new_n7120_));
  NOR2_X1    g04515(.A1(new_n7087_), .A2(new_n2622_), .ZN(new_n7121_));
  OAI21_X1   g04516(.A1(new_n7120_), .A2(new_n7117_), .B(new_n7121_), .ZN(new_n7122_));
  NOR2_X1    g04517(.A1(new_n3203_), .A2(pi0075), .ZN(new_n7123_));
  INV_X1     g04518(.I(new_n7123_), .ZN(new_n7124_));
  NAND2_X1   g04519(.A1(new_n7111_), .A2(pi0038), .ZN(new_n7125_));
  NAND2_X1   g04520(.A1(new_n7125_), .A2(new_n3173_), .ZN(new_n7126_));
  NOR2_X1    g04521(.A1(new_n7104_), .A2(new_n3173_), .ZN(new_n7127_));
  XNOR2_X1   g04522(.A1(new_n7127_), .A2(new_n7126_), .ZN(new_n7128_));
  INV_X1     g04523(.I(new_n7128_), .ZN(new_n7129_));
  NAND3_X1   g04524(.A1(new_n7122_), .A2(new_n7124_), .A3(new_n7129_), .ZN(new_n7130_));
  NAND2_X1   g04525(.A1(new_n7127_), .A2(new_n3177_), .ZN(new_n7131_));
  OR3_X2     g04526(.A1(new_n7128_), .A2(new_n3177_), .A3(new_n7121_), .Z(new_n7132_));
  OAI21_X1   g04527(.A1(new_n7105_), .A2(new_n2628_), .B(new_n3228_), .ZN(new_n7133_));
  AOI21_X1   g04528(.A1(new_n7132_), .A2(new_n7131_), .B(new_n7133_), .ZN(new_n7134_));
  AOI21_X1   g04529(.A1(new_n7130_), .A2(new_n7134_), .B(pi0054), .ZN(new_n7135_));
  OAI21_X1   g04530(.A1(new_n7135_), .A2(new_n7113_), .B(new_n3202_), .ZN(new_n7136_));
  NOR2_X1    g04531(.A1(pi0191), .A2(pi0299), .ZN(new_n7137_));
  AOI21_X1   g04532(.A1(new_n4272_), .A2(pi0299), .B(new_n7137_), .ZN(new_n7138_));
  AOI21_X1   g04533(.A1(new_n7049_), .A2(new_n7138_), .B(pi0074), .ZN(new_n7139_));
  NAND2_X1   g04534(.A1(new_n7108_), .A2(new_n7139_), .ZN(new_n7140_));
  NAND4_X1   g04535(.A1(new_n7136_), .A2(new_n3227_), .A3(new_n3503_), .A4(new_n7140_), .ZN(new_n7141_));
  AOI21_X1   g04536(.A1(new_n7099_), .A2(new_n7100_), .B(new_n7141_), .ZN(new_n7142_));
  NOR2_X1    g04537(.A1(new_n7087_), .A2(pi0038), .ZN(new_n7143_));
  INV_X1     g04538(.I(new_n7143_), .ZN(new_n7144_));
  NOR2_X1    g04539(.A1(new_n7144_), .A2(new_n7048_), .ZN(new_n7145_));
  INV_X1     g04540(.I(new_n7145_), .ZN(new_n7146_));
  NOR2_X1    g04541(.A1(new_n7146_), .A2(new_n2539_), .ZN(new_n7147_));
  AOI21_X1   g04542(.A1(new_n3503_), .A2(new_n7147_), .B(new_n7142_), .ZN(new_n7148_));
  OAI21_X1   g04543(.A1(new_n7148_), .A2(new_n7064_), .B(new_n7054_), .ZN(new_n7149_));
  INV_X1     g04544(.I(pi0176), .ZN(new_n7150_));
  INV_X1     g04545(.I(pi0174), .ZN(new_n7151_));
  INV_X1     g04546(.I(new_n5144_), .ZN(new_n7152_));
  NOR2_X1    g04547(.A1(new_n6051_), .A2(new_n2595_), .ZN(new_n7153_));
  INV_X1     g04548(.I(new_n7153_), .ZN(new_n7154_));
  NOR2_X1    g04549(.A1(new_n7152_), .A2(new_n7154_), .ZN(new_n7155_));
  INV_X1     g04550(.I(new_n7155_), .ZN(new_n7156_));
  NAND2_X1   g04551(.A1(new_n6047_), .A2(new_n7155_), .ZN(new_n7157_));
  AOI21_X1   g04552(.A1(new_n7151_), .A2(new_n7156_), .B(new_n7157_), .ZN(new_n7158_));
  NOR3_X1    g04553(.A1(new_n6047_), .A2(pi0174), .A3(new_n7156_), .ZN(new_n7159_));
  NOR4_X1    g04554(.A1(new_n7158_), .A2(new_n7150_), .A3(pi0299), .A4(new_n7159_), .ZN(new_n7160_));
  NOR2_X1    g04555(.A1(new_n5370_), .A2(new_n7152_), .ZN(new_n7161_));
  INV_X1     g04556(.I(new_n7161_), .ZN(new_n7162_));
  NOR2_X1    g04557(.A1(new_n7162_), .A2(new_n7154_), .ZN(new_n7163_));
  AOI21_X1   g04558(.A1(new_n7163_), .A2(new_n7151_), .B(pi0299), .ZN(new_n7164_));
  OAI21_X1   g04559(.A1(new_n7164_), .A2(pi0176), .B(new_n5987_), .ZN(new_n7165_));
  NOR2_X1    g04560(.A1(new_n5094_), .A2(new_n5109_), .ZN(new_n7166_));
  INV_X1     g04561(.I(new_n7166_), .ZN(new_n7167_));
  NOR2_X1    g04562(.A1(new_n6048_), .A2(new_n7167_), .ZN(new_n7168_));
  NAND3_X1   g04563(.A1(new_n7168_), .A2(pi0152), .A3(pi0154), .ZN(new_n7169_));
  NOR2_X1    g04564(.A1(new_n5357_), .A2(new_n2562_), .ZN(new_n7170_));
  NOR2_X1    g04565(.A1(new_n5370_), .A2(new_n7167_), .ZN(new_n7171_));
  AOI21_X1   g04566(.A1(new_n7167_), .A2(pi0154), .B(pi0152), .ZN(new_n7172_));
  OAI21_X1   g04567(.A1(new_n7171_), .A2(pi0154), .B(new_n7172_), .ZN(new_n7173_));
  NAND3_X1   g04568(.A1(new_n7169_), .A2(new_n7170_), .A3(new_n7173_), .ZN(new_n7174_));
  AOI21_X1   g04569(.A1(new_n7174_), .A2(pi0299), .B(new_n3154_), .ZN(new_n7175_));
  OAI21_X1   g04570(.A1(new_n7160_), .A2(new_n7165_), .B(new_n7175_), .ZN(new_n7176_));
  NOR2_X1    g04571(.A1(new_n5987_), .A2(pi0039), .ZN(new_n7177_));
  INV_X1     g04572(.I(new_n7177_), .ZN(new_n7178_));
  INV_X1     g04573(.I(pi0193), .ZN(new_n7179_));
  INV_X1     g04574(.I(pi0183), .ZN(new_n7180_));
  NOR2_X1    g04575(.A1(new_n3066_), .A2(new_n2485_), .ZN(new_n7181_));
  NOR2_X1    g04576(.A1(new_n5949_), .A2(pi0090), .ZN(new_n7182_));
  NAND3_X1   g04577(.A1(new_n7182_), .A2(new_n2478_), .A3(new_n5070_), .ZN(new_n7183_));
  INV_X1     g04578(.I(pi0060), .ZN(new_n7184_));
  AOI21_X1   g04579(.A1(new_n6985_), .A2(new_n7184_), .B(new_n2697_), .ZN(new_n7185_));
  INV_X1     g04580(.I(new_n7185_), .ZN(new_n7186_));
  NOR4_X1    g04581(.A1(new_n2884_), .A2(pi0090), .A3(new_n2478_), .A4(new_n2890_), .ZN(new_n7187_));
  AOI21_X1   g04582(.A1(new_n7186_), .A2(new_n7187_), .B(pi0070), .ZN(new_n7188_));
  NAND2_X1   g04583(.A1(new_n7188_), .A2(new_n7183_), .ZN(new_n7189_));
  NAND2_X1   g04584(.A1(new_n7189_), .A2(new_n7181_), .ZN(new_n7190_));
  INV_X1     g04585(.I(new_n7190_), .ZN(new_n7191_));
  NOR2_X1    g04586(.A1(new_n7191_), .A2(new_n5243_), .ZN(new_n7192_));
  NOR2_X1    g04587(.A1(new_n7192_), .A2(new_n5109_), .ZN(new_n7193_));
  INV_X1     g04588(.I(new_n2484_), .ZN(new_n7194_));
  NOR2_X1    g04589(.A1(new_n5109_), .A2(new_n7194_), .ZN(new_n7195_));
  INV_X1     g04590(.I(new_n7195_), .ZN(new_n7196_));
  NOR2_X1    g04591(.A1(new_n7196_), .A2(pi0040), .ZN(new_n7197_));
  INV_X1     g04592(.I(new_n7197_), .ZN(new_n7198_));
  NOR2_X1    g04593(.A1(pi0072), .A2(pi0093), .ZN(new_n7199_));
  INV_X1     g04594(.I(new_n7199_), .ZN(new_n7200_));
  NOR3_X1    g04595(.A1(new_n7182_), .A2(new_n2648_), .A3(new_n7200_), .ZN(new_n7201_));
  INV_X1     g04596(.I(new_n7201_), .ZN(new_n7202_));
  NOR2_X1    g04597(.A1(new_n7202_), .A2(new_n5069_), .ZN(new_n7203_));
  INV_X1     g04598(.I(new_n7203_), .ZN(new_n7204_));
  NOR2_X1    g04599(.A1(new_n7204_), .A2(new_n7198_), .ZN(new_n7205_));
  INV_X1     g04600(.I(new_n7205_), .ZN(new_n7206_));
  AOI21_X1   g04601(.A1(new_n7206_), .A2(new_n7180_), .B(pi0174), .ZN(new_n7207_));
  OAI21_X1   g04602(.A1(new_n7193_), .A2(new_n7180_), .B(new_n7207_), .ZN(new_n7208_));
  AOI21_X1   g04603(.A1(new_n7068_), .A2(new_n7077_), .B(new_n7185_), .ZN(new_n7209_));
  INV_X1     g04604(.I(new_n7068_), .ZN(new_n7210_));
  NOR2_X1    g04605(.A1(new_n7076_), .A2(new_n7070_), .ZN(new_n7211_));
  INV_X1     g04606(.I(pi0111), .ZN(new_n7212_));
  NAND4_X1   g04607(.A1(new_n2445_), .A2(new_n2449_), .A3(new_n2451_), .A4(new_n7212_), .ZN(new_n7213_));
  NOR2_X1    g04608(.A1(pi0082), .A2(pi0084), .ZN(new_n7214_));
  INV_X1     g04609(.I(new_n7214_), .ZN(new_n7215_));
  NOR4_X1    g04610(.A1(new_n7213_), .A2(pi0066), .A3(new_n2728_), .A4(new_n7215_), .ZN(new_n7216_));
  NAND3_X1   g04611(.A1(new_n7211_), .A2(new_n2729_), .A3(new_n7216_), .ZN(new_n7217_));
  AND3_X2    g04612(.A1(new_n7217_), .A2(new_n7000_), .A3(new_n7210_), .Z(new_n7218_));
  AOI21_X1   g04613(.A1(new_n7209_), .A2(new_n7218_), .B(new_n2683_), .ZN(new_n7219_));
  AND2_X2    g04614(.A1(new_n7187_), .A2(new_n2455_), .Z(new_n7220_));
  AOI21_X1   g04615(.A1(new_n7219_), .A2(new_n7220_), .B(pi0070), .ZN(new_n7221_));
  INV_X1     g04616(.I(new_n7221_), .ZN(new_n7222_));
  NAND2_X1   g04617(.A1(new_n7222_), .A2(new_n7183_), .ZN(new_n7223_));
  NAND2_X1   g04618(.A1(new_n7223_), .A2(new_n7181_), .ZN(new_n7224_));
  INV_X1     g04619(.I(new_n7224_), .ZN(new_n7225_));
  INV_X1     g04620(.I(new_n7181_), .ZN(new_n7226_));
  NAND2_X1   g04621(.A1(new_n2437_), .A2(pi0032), .ZN(new_n7227_));
  OAI22_X1   g04622(.A1(new_n7222_), .A2(new_n7226_), .B1(new_n5242_), .B2(new_n7227_), .ZN(new_n7228_));
  NOR2_X1    g04623(.A1(new_n7228_), .A2(pi0198), .ZN(new_n7229_));
  NOR2_X1    g04624(.A1(new_n7225_), .A2(new_n7229_), .ZN(new_n7230_));
  INV_X1     g04625(.I(new_n7230_), .ZN(new_n7231_));
  NOR2_X1    g04626(.A1(new_n7217_), .A2(new_n6999_), .ZN(new_n7232_));
  NAND2_X1   g04627(.A1(new_n7232_), .A2(new_n2455_), .ZN(new_n7233_));
  AOI21_X1   g04628(.A1(new_n5069_), .A2(new_n7233_), .B(new_n7202_), .ZN(new_n7234_));
  INV_X1     g04629(.I(new_n7234_), .ZN(new_n7235_));
  NOR2_X1    g04630(.A1(new_n7235_), .A2(new_n7198_), .ZN(new_n7236_));
  NAND4_X1   g04631(.A1(new_n7231_), .A2(pi0174), .A3(pi0183), .A4(new_n5108_), .ZN(new_n7237_));
  AOI21_X1   g04632(.A1(new_n7237_), .A2(new_n7208_), .B(new_n7179_), .ZN(new_n7238_));
  NOR2_X1    g04633(.A1(new_n7222_), .A2(new_n7226_), .ZN(new_n7239_));
  NOR2_X1    g04634(.A1(new_n7239_), .A2(new_n5330_), .ZN(new_n7240_));
  NOR4_X1    g04635(.A1(new_n7240_), .A2(new_n7224_), .A3(pi0152), .A4(new_n3707_), .ZN(new_n7241_));
  NOR2_X1    g04636(.A1(new_n7190_), .A2(new_n3707_), .ZN(new_n7242_));
  NOR2_X1    g04637(.A1(new_n7226_), .A2(new_n7188_), .ZN(new_n7243_));
  NOR2_X1    g04638(.A1(new_n7243_), .A2(new_n5330_), .ZN(new_n7244_));
  NAND2_X1   g04639(.A1(new_n7244_), .A2(pi0152), .ZN(new_n7245_));
  NOR2_X1    g04640(.A1(new_n5109_), .A2(new_n7067_), .ZN(new_n7246_));
  OAI21_X1   g04641(.A1(new_n7245_), .A2(new_n7242_), .B(new_n7246_), .ZN(new_n7247_));
  NOR2_X1    g04642(.A1(new_n5109_), .A2(pi0040), .ZN(new_n7248_));
  NOR3_X1    g04643(.A1(new_n2648_), .A2(pi0090), .A3(new_n7200_), .ZN(new_n7249_));
  INV_X1     g04644(.I(new_n7249_), .ZN(new_n7250_));
  NOR2_X1    g04645(.A1(new_n7233_), .A2(new_n7250_), .ZN(new_n7251_));
  INV_X1     g04646(.I(new_n7251_), .ZN(new_n7252_));
  NOR2_X1    g04647(.A1(new_n7252_), .A2(new_n7194_), .ZN(new_n7253_));
  NAND2_X1   g04648(.A1(new_n7253_), .A2(new_n7248_), .ZN(new_n7254_));
  INV_X1     g04649(.I(new_n7254_), .ZN(new_n7255_));
  AOI21_X1   g04650(.A1(new_n7236_), .A2(new_n3250_), .B(new_n7205_), .ZN(new_n7256_));
  NAND3_X1   g04651(.A1(new_n7255_), .A2(new_n3250_), .A3(new_n3707_), .ZN(new_n7257_));
  NAND3_X1   g04652(.A1(new_n7255_), .A2(new_n3250_), .A3(new_n3707_), .ZN(new_n7258_));
  NOR2_X1    g04653(.A1(new_n7256_), .A2(new_n3707_), .ZN(new_n7259_));
  AOI21_X1   g04654(.A1(new_n7259_), .A2(new_n7258_), .B(pi0149), .ZN(new_n7260_));
  NOR2_X1    g04655(.A1(new_n3100_), .A2(new_n5109_), .ZN(new_n7261_));
  INV_X1     g04656(.I(new_n7261_), .ZN(new_n7262_));
  OAI21_X1   g04657(.A1(new_n7262_), .A2(new_n5340_), .B(pi0299), .ZN(new_n7263_));
  AOI21_X1   g04658(.A1(new_n7260_), .A2(new_n7257_), .B(new_n7263_), .ZN(new_n7264_));
  OAI21_X1   g04659(.A1(new_n7241_), .A2(new_n7247_), .B(new_n7264_), .ZN(new_n7265_));
  NOR2_X1    g04660(.A1(new_n7239_), .A2(new_n5243_), .ZN(new_n7266_));
  NAND2_X1   g04661(.A1(new_n5108_), .A2(pi0183), .ZN(new_n7267_));
  NOR2_X1    g04662(.A1(new_n7243_), .A2(new_n5243_), .ZN(new_n7268_));
  INV_X1     g04663(.I(new_n7268_), .ZN(new_n7269_));
  NAND3_X1   g04664(.A1(new_n7269_), .A2(pi0174), .A3(new_n7267_), .ZN(new_n7270_));
  NAND2_X1   g04665(.A1(new_n7151_), .A2(new_n7180_), .ZN(new_n7271_));
  OAI22_X1   g04666(.A1(new_n7266_), .A2(new_n7270_), .B1(new_n7254_), .B2(new_n7271_), .ZN(new_n7272_));
  NAND2_X1   g04667(.A1(new_n7272_), .A2(new_n7179_), .ZN(new_n7273_));
  NAND2_X1   g04668(.A1(new_n7261_), .A2(pi0180), .ZN(new_n7274_));
  NAND4_X1   g04669(.A1(new_n7265_), .A2(new_n2587_), .A3(new_n7273_), .A4(new_n7274_), .ZN(new_n7275_));
  OAI21_X1   g04670(.A1(new_n7275_), .A2(new_n7238_), .B(new_n7178_), .ZN(new_n7276_));
  NAND2_X1   g04671(.A1(new_n7276_), .A2(new_n7176_), .ZN(new_n7277_));
  NAND2_X1   g04672(.A1(new_n7058_), .A2(pi0186), .ZN(new_n7278_));
  NOR3_X1    g04673(.A1(new_n5153_), .A2(new_n2587_), .A3(new_n5989_), .ZN(new_n7279_));
  INV_X1     g04674(.I(new_n7279_), .ZN(new_n7280_));
  NOR2_X1    g04675(.A1(new_n5156_), .A2(new_n5989_), .ZN(new_n7281_));
  OAI21_X1   g04676(.A1(new_n7280_), .A2(new_n7281_), .B(pi0186), .ZN(new_n7282_));
  NOR3_X1    g04677(.A1(new_n5153_), .A2(pi0299), .A3(new_n5989_), .ZN(new_n7283_));
  INV_X1     g04678(.I(new_n7283_), .ZN(new_n7284_));
  OAI22_X1   g04679(.A1(new_n7282_), .A2(new_n7058_), .B1(new_n7278_), .B2(new_n7284_), .ZN(new_n7285_));
  MUX2_X1    g04680(.I0(new_n7285_), .I1(new_n7277_), .S(new_n3172_), .Z(new_n7286_));
  NAND2_X1   g04681(.A1(new_n7286_), .A2(new_n3177_), .ZN(new_n7287_));
  OAI21_X1   g04682(.A1(new_n7125_), .A2(pi0087), .B(new_n3173_), .ZN(new_n7288_));
  AOI21_X1   g04683(.A1(new_n7287_), .A2(new_n7288_), .B(new_n7106_), .ZN(new_n7289_));
  NOR2_X1    g04684(.A1(pi0038), .A2(pi0087), .ZN(new_n7290_));
  NAND4_X1   g04685(.A1(new_n7117_), .A2(new_n3173_), .A3(new_n7124_), .A4(new_n7290_), .ZN(new_n7291_));
  NOR2_X1    g04686(.A1(new_n5154_), .A2(new_n7291_), .ZN(new_n7292_));
  AOI21_X1   g04687(.A1(new_n7292_), .A2(new_n7128_), .B(new_n7107_), .ZN(new_n7293_));
  OAI21_X1   g04688(.A1(new_n7289_), .A2(new_n3228_), .B(new_n7293_), .ZN(new_n7294_));
  AOI21_X1   g04689(.A1(new_n7294_), .A2(new_n3214_), .B(new_n7113_), .ZN(new_n7295_));
  NAND3_X1   g04690(.A1(new_n7140_), .A2(new_n3227_), .A3(new_n3202_), .ZN(new_n7296_));
  NOR3_X1    g04691(.A1(new_n5154_), .A2(new_n7067_), .A3(new_n5989_), .ZN(new_n7297_));
  NAND2_X1   g04692(.A1(new_n7059_), .A2(pi0087), .ZN(new_n7298_));
  NAND2_X1   g04693(.A1(new_n7298_), .A2(new_n3173_), .ZN(new_n7299_));
  NAND2_X1   g04694(.A1(new_n7045_), .A2(pi0100), .ZN(new_n7300_));
  OAI21_X1   g04695(.A1(new_n7299_), .A2(new_n7300_), .B(new_n7066_), .ZN(new_n7301_));
  AOI21_X1   g04696(.A1(new_n7299_), .A2(new_n7300_), .B(new_n7301_), .ZN(new_n7302_));
  OAI21_X1   g04697(.A1(new_n7297_), .A2(pi0038), .B(new_n7302_), .ZN(new_n7303_));
  MUX2_X1    g04698(.I0(new_n7303_), .I1(new_n7089_), .S(pi0075), .Z(new_n7304_));
  NOR2_X1    g04699(.A1(new_n7304_), .A2(pi0092), .ZN(new_n7305_));
  NAND2_X1   g04700(.A1(new_n7060_), .A2(pi0092), .ZN(new_n7306_));
  NAND3_X1   g04701(.A1(new_n7057_), .A2(new_n7306_), .A3(new_n3214_), .ZN(new_n7307_));
  OAI21_X1   g04702(.A1(new_n7305_), .A2(new_n7307_), .B(new_n3202_), .ZN(new_n7308_));
  OAI21_X1   g04703(.A1(new_n7063_), .A2(new_n3405_), .B(new_n5418_), .ZN(new_n7309_));
  AOI21_X1   g04704(.A1(new_n7308_), .A2(new_n7055_), .B(new_n7309_), .ZN(new_n7310_));
  OAI21_X1   g04705(.A1(new_n7295_), .A2(new_n7296_), .B(new_n7310_), .ZN(new_n7311_));
  NAND2_X1   g04706(.A1(new_n7311_), .A2(new_n7054_), .ZN(new_n7312_));
  INV_X1     g04707(.I(pi0033), .ZN(new_n7313_));
  INV_X1     g04708(.I(pi0034), .ZN(new_n7314_));
  INV_X1     g04709(.I(pi0079), .ZN(new_n7315_));
  NOR4_X1    g04710(.A1(pi0138), .A2(pi0139), .A3(pi0195), .A4(pi0196), .ZN(new_n7316_));
  NOR2_X1    g04711(.A1(new_n7316_), .A2(pi0118), .ZN(new_n7317_));
  NAND3_X1   g04712(.A1(new_n7317_), .A2(new_n7314_), .A3(new_n7315_), .ZN(new_n7318_));
  NAND2_X1   g04713(.A1(new_n7318_), .A2(new_n7313_), .ZN(new_n7319_));
  MUX2_X1    g04714(.I0(new_n7312_), .I1(new_n7149_), .S(new_n7319_), .Z(new_n7320_));
  OR2_X2     g04715(.A1(new_n7149_), .A2(new_n7313_), .Z(new_n7321_));
  NAND2_X1   g04716(.A1(new_n7312_), .A2(pi0033), .ZN(new_n7322_));
  AOI21_X1   g04717(.A1(new_n7322_), .A2(new_n7321_), .B(po1110), .ZN(new_n7323_));
  AOI21_X1   g04718(.A1(po1110), .A2(new_n7320_), .B(new_n7323_), .ZN(po0191));
  INV_X1     g04719(.I(pi0162), .ZN(new_n7325_));
  NOR2_X1    g04720(.A1(pi0149), .A2(pi0157), .ZN(new_n7326_));
  XOR2_X1    g04721(.A1(new_n7326_), .A2(new_n7325_), .Z(new_n7327_));
  XOR2_X1    g04722(.A1(new_n7327_), .A2(new_n5339_), .Z(new_n7328_));
  NAND2_X1   g04723(.A1(new_n7328_), .A2(new_n5109_), .ZN(new_n7329_));
  NOR2_X1    g04724(.A1(new_n7329_), .A2(new_n5987_), .ZN(new_n7330_));
  NOR4_X1    g04725(.A1(new_n5989_), .A2(new_n7048_), .A3(pi0074), .A4(new_n4130_), .ZN(new_n7331_));
  INV_X1     g04726(.I(new_n7330_), .ZN(new_n7332_));
  NOR2_X1    g04727(.A1(new_n7332_), .A2(new_n7041_), .ZN(new_n7333_));
  INV_X1     g04728(.I(pi0167), .ZN(new_n7334_));
  NOR2_X1    g04729(.A1(new_n7050_), .A2(new_n7334_), .ZN(new_n7335_));
  NOR2_X1    g04730(.A1(new_n7333_), .A2(new_n7335_), .ZN(new_n7336_));
  AOI21_X1   g04731(.A1(new_n7336_), .A2(new_n3202_), .B(new_n7331_), .ZN(new_n7337_));
  NAND2_X1   g04732(.A1(new_n7337_), .A2(new_n3405_), .ZN(new_n7338_));
  INV_X1     g04733(.I(pi0140), .ZN(new_n7339_));
  NOR2_X1    g04734(.A1(new_n7339_), .A2(new_n5323_), .ZN(new_n7340_));
  NOR3_X1    g04735(.A1(new_n7340_), .A2(pi0178), .A3(pi0183), .ZN(new_n7341_));
  INV_X1     g04736(.I(new_n7341_), .ZN(new_n7342_));
  NOR2_X1    g04737(.A1(pi0140), .A2(pi0145), .ZN(new_n7343_));
  NOR2_X1    g04738(.A1(new_n5109_), .A2(new_n7343_), .ZN(new_n7344_));
  INV_X1     g04739(.I(pi0178), .ZN(new_n7345_));
  AOI21_X1   g04740(.A1(new_n7345_), .A2(new_n7180_), .B(new_n5109_), .ZN(new_n7346_));
  OAI21_X1   g04741(.A1(new_n7340_), .A2(new_n7343_), .B(new_n7346_), .ZN(new_n7347_));
  NOR2_X1    g04742(.A1(pi0232), .A2(pi0299), .ZN(new_n7348_));
  NAND2_X1   g04743(.A1(new_n7347_), .A2(new_n7348_), .ZN(new_n7349_));
  AOI21_X1   g04744(.A1(new_n7342_), .A2(new_n7344_), .B(new_n7349_), .ZN(new_n7350_));
  NAND3_X1   g04745(.A1(new_n7350_), .A2(new_n5109_), .A3(new_n7328_), .ZN(new_n7351_));
  INV_X1     g04746(.I(new_n7351_), .ZN(new_n7352_));
  NOR2_X1    g04747(.A1(new_n7352_), .A2(new_n3173_), .ZN(new_n7353_));
  NOR2_X1    g04748(.A1(new_n7352_), .A2(new_n2628_), .ZN(new_n7354_));
  NOR2_X1    g04749(.A1(new_n7353_), .A2(new_n7354_), .ZN(new_n7355_));
  INV_X1     g04750(.I(pi0188), .ZN(new_n7356_));
  MUX2_X1    g04751(.I0(new_n7356_), .I1(new_n7334_), .S(pi0299), .Z(new_n7357_));
  NOR2_X1    g04752(.A1(new_n5989_), .A2(new_n7357_), .ZN(new_n7358_));
  NOR2_X1    g04753(.A1(new_n7358_), .A2(pi0100), .ZN(new_n7359_));
  INV_X1     g04754(.I(new_n7359_), .ZN(new_n7360_));
  NOR2_X1    g04755(.A1(pi0054), .A2(pi0075), .ZN(new_n7361_));
  INV_X1     g04756(.I(new_n7361_), .ZN(new_n7362_));
  NOR3_X1    g04757(.A1(new_n7355_), .A2(new_n7360_), .A3(new_n7362_), .ZN(new_n7363_));
  INV_X1     g04758(.I(new_n7363_), .ZN(new_n7364_));
  OAI21_X1   g04759(.A1(new_n7082_), .A2(new_n7000_), .B(pi0070), .ZN(new_n7365_));
  AOI21_X1   g04760(.A1(new_n2478_), .A2(new_n2455_), .B(pi0070), .ZN(new_n7366_));
  INV_X1     g04761(.I(new_n7366_), .ZN(new_n7367_));
  INV_X1     g04762(.I(pi0058), .ZN(new_n7368_));
  AOI21_X1   g04763(.A1(new_n7079_), .A2(new_n2455_), .B(new_n7368_), .ZN(new_n7369_));
  INV_X1     g04764(.I(new_n7369_), .ZN(new_n7370_));
  INV_X1     g04765(.I(new_n7219_), .ZN(new_n7371_));
  AOI21_X1   g04766(.A1(new_n7000_), .A2(new_n2683_), .B(new_n2888_), .ZN(new_n7372_));
  OAI21_X1   g04767(.A1(new_n2888_), .A2(new_n2455_), .B(new_n7368_), .ZN(new_n7373_));
  AOI21_X1   g04768(.A1(new_n7371_), .A2(new_n7372_), .B(new_n7373_), .ZN(new_n7374_));
  NOR2_X1    g04769(.A1(new_n7081_), .A2(pi0841), .ZN(new_n7375_));
  INV_X1     g04770(.I(new_n7375_), .ZN(new_n7376_));
  NOR3_X1    g04771(.A1(new_n7000_), .A2(pi0090), .A3(new_n2477_), .ZN(new_n7377_));
  AOI21_X1   g04772(.A1(new_n7376_), .A2(new_n7377_), .B(pi0090), .ZN(new_n7378_));
  INV_X1     g04773(.I(new_n7378_), .ZN(new_n7379_));
  AOI21_X1   g04774(.A1(new_n7374_), .A2(new_n7370_), .B(new_n7379_), .ZN(new_n7380_));
  OAI21_X1   g04775(.A1(new_n7380_), .A2(new_n7367_), .B(new_n7365_), .ZN(new_n7381_));
  NOR2_X1    g04776(.A1(new_n2503_), .A2(pi0051), .ZN(new_n7382_));
  AOI21_X1   g04777(.A1(new_n2455_), .A2(new_n7382_), .B(new_n7381_), .ZN(new_n7383_));
  NAND3_X1   g04778(.A1(new_n7381_), .A2(new_n7000_), .A3(new_n7382_), .ZN(new_n7384_));
  NAND2_X1   g04779(.A1(new_n7384_), .A2(new_n3364_), .ZN(new_n7385_));
  OAI21_X1   g04780(.A1(new_n7385_), .A2(new_n7383_), .B(new_n2632_), .ZN(new_n7386_));
  OAI21_X1   g04781(.A1(new_n2632_), .A2(new_n7086_), .B(new_n7386_), .ZN(new_n7387_));
  NAND2_X1   g04782(.A1(new_n7387_), .A2(new_n2437_), .ZN(new_n7388_));
  NAND2_X1   g04783(.A1(new_n7083_), .A2(new_n2455_), .ZN(new_n7389_));
  INV_X1     g04784(.I(new_n7389_), .ZN(new_n7390_));
  NOR3_X1    g04785(.A1(pi0040), .A2(pi0095), .A3(pi0479), .ZN(new_n7391_));
  NAND2_X1   g04786(.A1(new_n7390_), .A2(new_n7391_), .ZN(new_n7392_));
  NAND2_X1   g04787(.A1(new_n7388_), .A2(new_n7392_), .ZN(new_n7393_));
  INV_X1     g04788(.I(new_n7393_), .ZN(new_n7394_));
  AOI21_X1   g04789(.A1(new_n7375_), .A2(new_n7249_), .B(new_n7087_), .ZN(new_n7395_));
  NOR2_X1    g04790(.A1(new_n7395_), .A2(new_n2632_), .ZN(new_n7396_));
  INV_X1     g04791(.I(new_n7396_), .ZN(new_n7397_));
  NAND2_X1   g04792(.A1(new_n7386_), .A2(new_n7397_), .ZN(new_n7398_));
  NAND2_X1   g04793(.A1(new_n7398_), .A2(new_n2437_), .ZN(new_n7399_));
  NOR3_X1    g04794(.A1(new_n7394_), .A2(new_n5081_), .A3(new_n7399_), .ZN(new_n7400_));
  NOR2_X1    g04795(.A1(new_n2587_), .A2(pi0159), .ZN(new_n7401_));
  INV_X1     g04796(.I(new_n7392_), .ZN(new_n7402_));
  AOI21_X1   g04797(.A1(new_n2437_), .A2(new_n7087_), .B(new_n7402_), .ZN(new_n7403_));
  NOR2_X1    g04798(.A1(new_n7399_), .A2(pi0210), .ZN(new_n7405_));
  NOR2_X1    g04799(.A1(new_n7393_), .A2(new_n7405_), .ZN(new_n7406_));
  AOI21_X1   g04800(.A1(new_n7000_), .A2(pi0032), .B(pi0040), .ZN(new_n7409_));
  INV_X1     g04801(.I(new_n7409_), .ZN(new_n7410_));
  AOI21_X1   g04802(.A1(new_n7376_), .A2(pi0090), .B(new_n2455_), .ZN(new_n7411_));
  OAI21_X1   g04803(.A1(pi0090), .A2(new_n7369_), .B(new_n7411_), .ZN(new_n7412_));
  NAND2_X1   g04804(.A1(new_n7412_), .A2(new_n2841_), .ZN(new_n7413_));
  AOI21_X1   g04805(.A1(new_n5083_), .A2(new_n2455_), .B(pi0032), .ZN(new_n7414_));
  OAI21_X1   g04806(.A1(new_n2841_), .A2(new_n2455_), .B(new_n5082_), .ZN(new_n7415_));
  NOR2_X1    g04807(.A1(new_n7414_), .A2(new_n7415_), .ZN(new_n7416_));
  AOI21_X1   g04808(.A1(new_n7413_), .A2(new_n7416_), .B(new_n7410_), .ZN(new_n7417_));
  NOR2_X1    g04809(.A1(new_n7417_), .A2(pi0095), .ZN(new_n7418_));
  INV_X1     g04810(.I(new_n7418_), .ZN(new_n7419_));
  AOI21_X1   g04811(.A1(new_n7419_), .A2(new_n7392_), .B(new_n5109_), .ZN(new_n7420_));
  NAND3_X1   g04812(.A1(new_n7412_), .A2(new_n2839_), .A3(new_n7232_), .ZN(new_n7423_));
  NOR4_X1    g04813(.A1(new_n7414_), .A2(pi0093), .A3(new_n7409_), .A4(new_n7415_), .ZN(new_n7424_));
  NAND2_X1   g04814(.A1(new_n7423_), .A2(new_n7424_), .ZN(new_n7425_));
  NAND2_X1   g04815(.A1(new_n7392_), .A2(new_n5109_), .ZN(new_n7426_));
  AOI21_X1   g04816(.A1(new_n7425_), .A2(new_n2437_), .B(new_n7426_), .ZN(new_n7427_));
  NAND3_X1   g04817(.A1(new_n5082_), .A2(new_n2649_), .A3(new_n6998_), .ZN(new_n7430_));
  NOR4_X1    g04818(.A1(new_n7217_), .A2(pi0032), .A3(new_n7086_), .A4(new_n7430_), .ZN(new_n7431_));
  INV_X1     g04819(.I(new_n7078_), .ZN(new_n7440_));
  NOR3_X1    g04820(.A1(new_n7209_), .A2(new_n2455_), .A3(new_n7440_), .ZN(new_n7441_));
  NOR2_X1    g04821(.A1(new_n7441_), .A2(pi0058), .ZN(new_n7442_));
  AOI21_X1   g04822(.A1(new_n7442_), .A2(new_n7370_), .B(new_n7379_), .ZN(new_n7443_));
  OAI21_X1   g04823(.A1(new_n7443_), .A2(new_n7367_), .B(new_n7365_), .ZN(new_n7444_));
  MUX2_X1    g04824(.I0(new_n7444_), .I1(new_n2455_), .S(new_n7382_), .Z(new_n7445_));
  AOI21_X1   g04825(.A1(new_n7445_), .A2(new_n3364_), .B(pi0032), .ZN(new_n7446_));
  OAI21_X1   g04826(.A1(new_n7446_), .A2(new_n7396_), .B(new_n2437_), .ZN(new_n7447_));
  NOR2_X1    g04827(.A1(new_n7447_), .A2(pi0210), .ZN(new_n7448_));
  NOR2_X1    g04828(.A1(new_n7086_), .A2(new_n2632_), .ZN(new_n7449_));
  OAI21_X1   g04829(.A1(new_n7446_), .A2(new_n7449_), .B(new_n2437_), .ZN(new_n7450_));
  NAND2_X1   g04830(.A1(new_n7450_), .A2(new_n7392_), .ZN(new_n7451_));
  NOR2_X1    g04831(.A1(new_n7448_), .A2(new_n7451_), .ZN(new_n7452_));
  INV_X1     g04832(.I(new_n7452_), .ZN(new_n7453_));
  NOR2_X1    g04833(.A1(new_n7453_), .A2(new_n5109_), .ZN(new_n7454_));
  INV_X1     g04834(.I(new_n7365_), .ZN(new_n7459_));
  NAND2_X1   g04835(.A1(new_n2509_), .A2(new_n7000_), .ZN(new_n7460_));
  OR2_X2     g04836(.A1(new_n7374_), .A2(new_n5965_), .Z(new_n7461_));
  AOI21_X1   g04837(.A1(new_n7461_), .A2(new_n7460_), .B(pi0070), .ZN(new_n7462_));
  AOI21_X1   g04838(.A1(new_n2861_), .A2(new_n2659_), .B(pi0051), .ZN(new_n7463_));
  OAI21_X1   g04839(.A1(new_n7462_), .A2(new_n7459_), .B(new_n7463_), .ZN(new_n7464_));
  AOI21_X1   g04840(.A1(new_n2503_), .A2(new_n2455_), .B(pi0040), .ZN(new_n7465_));
  NAND2_X1   g04841(.A1(new_n7464_), .A2(new_n7465_), .ZN(new_n7466_));
  NOR2_X1    g04842(.A1(new_n2455_), .A2(pi0040), .ZN(new_n7467_));
  INV_X1     g04843(.I(new_n7467_), .ZN(new_n7468_));
  NOR2_X1    g04844(.A1(new_n7468_), .A2(new_n2632_), .ZN(new_n7469_));
  AOI21_X1   g04845(.A1(new_n7466_), .A2(new_n2632_), .B(new_n7469_), .ZN(new_n7470_));
  OAI21_X1   g04846(.A1(new_n2962_), .A2(new_n7086_), .B(new_n7470_), .ZN(new_n7471_));
  NAND2_X1   g04847(.A1(new_n7471_), .A2(new_n2437_), .ZN(new_n7472_));
  NOR2_X1    g04848(.A1(new_n7472_), .A2(new_n7402_), .ZN(new_n7473_));
  NOR2_X1    g04849(.A1(new_n7086_), .A2(new_n2437_), .ZN(new_n7474_));
  NOR2_X1    g04850(.A1(new_n7472_), .A2(new_n7474_), .ZN(new_n7475_));
  OAI21_X1   g04851(.A1(new_n7395_), .A2(pi0040), .B(pi0032), .ZN(new_n7476_));
  OAI21_X1   g04852(.A1(new_n7466_), .A2(pi0032), .B(new_n7476_), .ZN(new_n7477_));
  NAND2_X1   g04853(.A1(new_n7477_), .A2(new_n2437_), .ZN(new_n7478_));
  NOR2_X1    g04854(.A1(new_n7467_), .A2(new_n2437_), .ZN(new_n7479_));
  NOR2_X1    g04855(.A1(new_n7478_), .A2(new_n7479_), .ZN(new_n7480_));
  INV_X1     g04856(.I(new_n7480_), .ZN(new_n7481_));
  NAND2_X1   g04857(.A1(new_n7475_), .A2(new_n7481_), .ZN(new_n7482_));
  AOI21_X1   g04858(.A1(new_n7482_), .A2(new_n2631_), .B(new_n5109_), .ZN(new_n7483_));
  NOR2_X1    g04859(.A1(new_n7086_), .A2(new_n5109_), .ZN(new_n7484_));
  OAI21_X1   g04860(.A1(new_n7483_), .A2(new_n7484_), .B(new_n7473_), .ZN(new_n7485_));
  OAI21_X1   g04861(.A1(new_n7442_), .A2(new_n5965_), .B(new_n7460_), .ZN(new_n7486_));
  AOI21_X1   g04862(.A1(new_n7486_), .A2(new_n2849_), .B(new_n7459_), .ZN(new_n7487_));
  MUX2_X1    g04863(.I0(new_n7487_), .I1(new_n2455_), .S(new_n7382_), .Z(new_n7488_));
  NAND2_X1   g04864(.A1(new_n7488_), .A2(new_n3364_), .ZN(new_n7489_));
  NAND2_X1   g04865(.A1(new_n7489_), .A2(new_n2632_), .ZN(new_n7490_));
  INV_X1     g04866(.I(new_n7490_), .ZN(new_n7491_));
  OAI21_X1   g04867(.A1(new_n7491_), .A2(new_n7449_), .B(new_n2437_), .ZN(new_n7492_));
  INV_X1     g04868(.I(new_n7492_), .ZN(new_n7493_));
  NOR2_X1    g04869(.A1(new_n7493_), .A2(new_n7402_), .ZN(new_n7494_));
  AOI21_X1   g04870(.A1(new_n7490_), .A2(new_n7397_), .B(pi0095), .ZN(new_n7495_));
  NOR2_X1    g04871(.A1(new_n5108_), .A2(pi0210), .ZN(new_n7496_));
  OAI21_X1   g04872(.A1(new_n7495_), .A2(new_n7474_), .B(new_n7496_), .ZN(new_n7497_));
  OAI21_X1   g04873(.A1(new_n5109_), .A2(new_n7086_), .B(new_n7497_), .ZN(new_n7498_));
  AND2_X2    g04874(.A1(new_n7498_), .A2(new_n7494_), .Z(new_n7499_));
  INV_X1     g04875(.I(pi0144), .ZN(new_n7504_));
  NOR2_X1    g04876(.A1(new_n7399_), .A2(pi0198), .ZN(new_n7505_));
  NOR2_X1    g04877(.A1(new_n7393_), .A2(new_n7505_), .ZN(new_n7506_));
  INV_X1     g04878(.I(new_n7506_), .ZN(new_n7511_));
  NAND2_X1   g04879(.A1(new_n7495_), .A2(new_n2601_), .ZN(new_n7513_));
  NAND2_X1   g04880(.A1(new_n7494_), .A2(new_n7513_), .ZN(new_n7514_));
  NOR2_X1    g04881(.A1(new_n7447_), .A2(pi0198), .ZN(new_n7517_));
  NOR2_X1    g04882(.A1(new_n7517_), .A2(new_n7451_), .ZN(new_n7518_));
  INV_X1     g04883(.I(new_n7518_), .ZN(new_n7519_));
  OAI21_X1   g04884(.A1(new_n7488_), .A2(pi0040), .B(new_n2632_), .ZN(new_n7531_));
  AOI21_X1   g04885(.A1(new_n7531_), .A2(new_n7476_), .B(pi0095), .ZN(new_n7532_));
  NOR2_X1    g04886(.A1(new_n7532_), .A2(new_n7479_), .ZN(new_n7533_));
  NOR2_X1    g04887(.A1(new_n7467_), .A2(new_n2632_), .ZN(new_n7534_));
  INV_X1     g04888(.I(new_n7534_), .ZN(new_n7535_));
  AOI21_X1   g04889(.A1(new_n7531_), .A2(new_n7535_), .B(pi0095), .ZN(new_n7536_));
  NOR3_X1    g04890(.A1(new_n7536_), .A2(new_n2601_), .A3(new_n7479_), .ZN(new_n7537_));
  AOI21_X1   g04891(.A1(new_n2601_), .A2(new_n7533_), .B(new_n7537_), .ZN(new_n7538_));
  AOI21_X1   g04892(.A1(new_n7482_), .A2(new_n2601_), .B(new_n5109_), .ZN(new_n7556_));
  OAI21_X1   g04893(.A1(new_n2437_), .A2(new_n7086_), .B(new_n7388_), .ZN(new_n7559_));
  NOR2_X1    g04894(.A1(new_n7559_), .A2(new_n7505_), .ZN(new_n7560_));
  NOR2_X1    g04895(.A1(new_n7556_), .A2(new_n7484_), .ZN(new_n7564_));
  NOR3_X1    g04896(.A1(new_n7564_), .A2(new_n7402_), .A3(new_n7472_), .ZN(new_n7565_));
  NOR2_X1    g04897(.A1(new_n7559_), .A2(new_n7405_), .ZN(new_n7573_));
  NOR2_X1    g04898(.A1(new_n5341_), .A2(new_n2587_), .ZN(new_n7593_));
  NOR2_X1    g04899(.A1(new_n7400_), .A2(pi0232), .ZN(new_n7595_));
  NOR2_X1    g04900(.A1(new_n7087_), .A2(new_n7170_), .ZN(new_n7596_));
  NOR2_X1    g04901(.A1(new_n7596_), .A2(new_n2587_), .ZN(new_n7597_));
  INV_X1     g04902(.I(new_n5134_), .ZN(new_n7598_));
  NOR3_X1    g04903(.A1(new_n5364_), .A2(new_n2923_), .A3(new_n5368_), .ZN(new_n7599_));
  NAND2_X1   g04904(.A1(new_n7599_), .A2(new_n5124_), .ZN(new_n7600_));
  AOI21_X1   g04905(.A1(new_n7598_), .A2(new_n7600_), .B(new_n7118_), .ZN(new_n7601_));
  AOI21_X1   g04906(.A1(new_n7601_), .A2(new_n5143_), .B(new_n7087_), .ZN(new_n7602_));
  NAND2_X1   g04907(.A1(new_n7601_), .A2(new_n7484_), .ZN(new_n7603_));
  NAND3_X1   g04908(.A1(new_n7602_), .A2(new_n7603_), .A3(new_n6445_), .ZN(new_n7604_));
  NOR2_X1    g04909(.A1(new_n7087_), .A2(new_n7153_), .ZN(new_n7605_));
  INV_X1     g04910(.I(new_n7603_), .ZN(new_n7606_));
  NOR2_X1    g04911(.A1(new_n7606_), .A2(new_n5141_), .ZN(new_n7607_));
  AOI21_X1   g04912(.A1(new_n7607_), .A2(new_n7602_), .B(new_n7605_), .ZN(new_n7608_));
  AOI22_X1   g04913(.A1(new_n7608_), .A2(new_n2587_), .B1(new_n7604_), .B2(new_n7597_), .ZN(new_n7609_));
  NOR3_X1    g04914(.A1(new_n7118_), .A2(new_n7598_), .A3(new_n7152_), .ZN(new_n7610_));
  AOI21_X1   g04915(.A1(new_n7610_), .A2(new_n7153_), .B(new_n7087_), .ZN(new_n7611_));
  INV_X1     g04916(.I(new_n7602_), .ZN(new_n7612_));
  NOR2_X1    g04917(.A1(pi0177), .A2(pi0299), .ZN(new_n7615_));
  INV_X1     g04918(.I(new_n7615_), .ZN(new_n7616_));
  INV_X1     g04919(.I(pi0177), .ZN(new_n7620_));
  NOR2_X1    g04920(.A1(new_n7620_), .A2(pi0299), .ZN(new_n7621_));
  INV_X1     g04921(.I(new_n7621_), .ZN(new_n7622_));
  NOR2_X1    g04922(.A1(new_n7118_), .A2(new_n7600_), .ZN(new_n7623_));
  AOI21_X1   g04923(.A1(new_n7623_), .A2(new_n7484_), .B(new_n5141_), .ZN(new_n7624_));
  NOR2_X1    g04924(.A1(new_n7609_), .A2(pi0232), .ZN(new_n7627_));
  INV_X1     g04925(.I(new_n7597_), .ZN(new_n7628_));
  NOR2_X1    g04926(.A1(new_n7118_), .A2(new_n7598_), .ZN(new_n7629_));
  AOI21_X1   g04927(.A1(new_n7629_), .A2(new_n6446_), .B(new_n7087_), .ZN(new_n7630_));
  NAND3_X1   g04928(.A1(new_n7630_), .A2(new_n4701_), .A3(new_n5108_), .ZN(new_n7631_));
  AOI21_X1   g04929(.A1(new_n7604_), .A2(new_n7631_), .B(new_n7170_), .ZN(new_n7632_));
  NOR4_X1    g04930(.A1(new_n7632_), .A2(pi0038), .A3(pi0155), .A4(new_n7628_), .ZN(new_n7633_));
  INV_X1     g04931(.I(new_n7170_), .ZN(new_n7634_));
  INV_X1     g04932(.I(new_n7623_), .ZN(new_n7635_));
  NAND2_X1   g04933(.A1(new_n7087_), .A2(new_n5109_), .ZN(new_n7636_));
  NOR4_X1    g04934(.A1(new_n7635_), .A2(new_n4701_), .A3(new_n5094_), .A4(new_n7636_), .ZN(new_n7637_));
  NOR3_X1    g04935(.A1(new_n7612_), .A2(new_n7637_), .A3(new_n7634_), .ZN(new_n7638_));
  INV_X1     g04936(.I(pi0155), .ZN(new_n7639_));
  NOR2_X1    g04937(.A1(new_n7639_), .A2(pi0038), .ZN(new_n7640_));
  NAND2_X1   g04938(.A1(new_n7597_), .A2(new_n7640_), .ZN(new_n7641_));
  OAI21_X1   g04939(.A1(new_n7638_), .A2(new_n7641_), .B(pi0232), .ZN(new_n7642_));
  OAI22_X1   g04940(.A1(new_n7627_), .A2(pi0038), .B1(new_n7633_), .B2(new_n7642_), .ZN(new_n7643_));
  AOI21_X1   g04941(.A1(new_n7358_), .A2(pi0038), .B(new_n7143_), .ZN(new_n7644_));
  NAND2_X1   g04942(.A1(new_n3177_), .A2(new_n3173_), .ZN(new_n7645_));
  AOI21_X1   g04943(.A1(new_n7643_), .A2(pi0039), .B(new_n7645_), .ZN(new_n7646_));
  OAI21_X1   g04944(.A1(new_n7595_), .A2(new_n2545_), .B(new_n7646_), .ZN(new_n7647_));
  INV_X1     g04945(.I(new_n7644_), .ZN(new_n7648_));
  OAI21_X1   g04946(.A1(pi0177), .A2(pi0299), .B(pi0155), .ZN(new_n7649_));
  NAND3_X1   g04947(.A1(new_n7639_), .A2(new_n2587_), .A3(pi0177), .ZN(new_n7650_));
  NAND4_X1   g04948(.A1(new_n5988_), .A2(new_n3172_), .A3(new_n7649_), .A4(new_n7650_), .ZN(new_n7651_));
  NOR3_X1    g04949(.A1(new_n7119_), .A2(new_n7648_), .A3(new_n7651_), .ZN(new_n7652_));
  NAND3_X1   g04950(.A1(new_n7351_), .A2(pi0100), .A3(new_n7124_), .ZN(new_n7653_));
  OAI22_X1   g04951(.A1(new_n7652_), .A2(new_n7653_), .B1(new_n2628_), .B2(new_n7352_), .ZN(new_n7654_));
  AOI21_X1   g04952(.A1(new_n7647_), .A2(new_n3209_), .B(new_n7654_), .ZN(new_n7655_));
  OAI21_X1   g04953(.A1(new_n7655_), .A2(pi0054), .B(new_n7364_), .ZN(new_n7656_));
  NOR2_X1    g04954(.A1(pi0141), .A2(pi0299), .ZN(new_n7657_));
  AOI21_X1   g04955(.A1(new_n4130_), .A2(pi0299), .B(new_n7657_), .ZN(new_n7658_));
  NAND2_X1   g04956(.A1(new_n5988_), .A2(new_n7658_), .ZN(new_n7659_));
  INV_X1     g04957(.I(new_n7659_), .ZN(new_n7660_));
  NOR2_X1    g04958(.A1(new_n3227_), .A2(pi0074), .ZN(new_n7661_));
  NAND2_X1   g04959(.A1(new_n5108_), .A2(pi0162), .ZN(new_n7662_));
  AOI21_X1   g04960(.A1(new_n7119_), .A2(new_n7662_), .B(new_n7144_), .ZN(new_n7663_));
  OAI22_X1   g04961(.A1(new_n7663_), .A2(pi0100), .B1(pi0232), .B2(new_n7120_), .ZN(new_n7664_));
  NAND3_X1   g04962(.A1(new_n5988_), .A2(pi0038), .A3(pi0167), .ZN(new_n7665_));
  AOI22_X1   g04963(.A1(new_n7664_), .A2(new_n7665_), .B1(pi0100), .B2(new_n7332_), .ZN(new_n7666_));
  MUX2_X1    g04964(.I0(new_n7666_), .I1(new_n7330_), .S(pi0075), .Z(new_n7667_));
  AOI21_X1   g04965(.A1(new_n7335_), .A2(pi0038), .B(pi0054), .ZN(new_n7668_));
  OAI21_X1   g04966(.A1(new_n7332_), .A2(new_n7041_), .B(new_n7668_), .ZN(new_n7669_));
  NAND2_X1   g04967(.A1(new_n7669_), .A2(new_n7146_), .ZN(new_n7670_));
  AOI22_X1   g04968(.A1(new_n7667_), .A2(new_n3203_), .B1(new_n5410_), .B2(new_n7670_), .ZN(new_n7671_));
  NOR3_X1    g04969(.A1(new_n7333_), .A2(new_n3214_), .A3(new_n7335_), .ZN(new_n7672_));
  NOR2_X1    g04970(.A1(new_n7331_), .A2(new_n3227_), .ZN(new_n7673_));
  NOR3_X1    g04971(.A1(new_n7673_), .A2(pi0074), .A3(new_n2533_), .ZN(new_n7674_));
  OAI21_X1   g04972(.A1(new_n7671_), .A2(new_n7672_), .B(new_n7674_), .ZN(new_n7675_));
  AOI21_X1   g04973(.A1(new_n7656_), .A2(new_n7661_), .B(new_n7675_), .ZN(new_n7676_));
  NAND2_X1   g04974(.A1(new_n7669_), .A2(new_n3202_), .ZN(new_n7677_));
  NOR2_X1    g04975(.A1(new_n3405_), .A2(new_n2533_), .ZN(new_n7678_));
  OAI21_X1   g04976(.A1(new_n7337_), .A2(new_n7677_), .B(new_n7678_), .ZN(new_n7679_));
  INV_X1     g04977(.I(new_n7147_), .ZN(new_n7680_));
  AOI21_X1   g04978(.A1(new_n7680_), .A2(new_n3503_), .B(new_n3405_), .ZN(new_n7681_));
  INV_X1     g04979(.I(new_n7681_), .ZN(new_n7682_));
  AND2_X2    g04980(.A1(new_n7679_), .A2(new_n7682_), .Z(new_n7683_));
  OAI21_X1   g04981(.A1(new_n7676_), .A2(new_n7683_), .B(new_n7338_), .ZN(new_n7684_));
  INV_X1     g04982(.I(new_n7661_), .ZN(new_n7685_));
  NAND2_X1   g04983(.A1(new_n7225_), .A2(new_n5460_), .ZN(new_n7686_));
  NAND3_X1   g04984(.A1(new_n7686_), .A2(pi0140), .A3(new_n7266_), .ZN(new_n7687_));
  NOR2_X1    g04985(.A1(new_n7236_), .A2(new_n5460_), .ZN(new_n7688_));
  OAI21_X1   g04986(.A1(new_n7254_), .A2(new_n5460_), .B(new_n7339_), .ZN(new_n7689_));
  NOR2_X1    g04987(.A1(new_n7688_), .A2(new_n7689_), .ZN(new_n7690_));
  OAI21_X1   g04988(.A1(new_n5108_), .A2(new_n7339_), .B(new_n7504_), .ZN(new_n7694_));
  AOI21_X1   g04989(.A1(new_n7687_), .A2(new_n7690_), .B(new_n7694_), .ZN(new_n7695_));
  INV_X1     g04990(.I(new_n7240_), .ZN(new_n7696_));
  NAND3_X1   g04991(.A1(new_n7696_), .A2(new_n7225_), .A3(new_n3560_), .ZN(new_n7697_));
  NOR4_X1    g04992(.A1(new_n7244_), .A2(new_n7190_), .A3(pi0146), .A4(pi0161), .ZN(new_n7698_));
  NOR4_X1    g04993(.A1(new_n7262_), .A2(new_n5341_), .A3(pi0162), .A4(pi0299), .ZN(new_n7699_));
  NAND4_X1   g04994(.A1(new_n7662_), .A2(pi0159), .A3(new_n4701_), .A4(new_n2587_), .ZN(new_n7700_));
  NOR4_X1    g04995(.A1(new_n7698_), .A2(new_n3100_), .A3(new_n7699_), .A4(new_n7700_), .ZN(new_n7701_));
  MUX2_X1    g04996(.I0(new_n7255_), .I1(new_n7236_), .S(new_n3560_), .Z(new_n7702_));
  NAND2_X1   g04997(.A1(new_n3560_), .A2(pi0161), .ZN(new_n7703_));
  OAI21_X1   g04998(.A1(new_n7206_), .A2(new_n7703_), .B(new_n7325_), .ZN(new_n7704_));
  AOI21_X1   g04999(.A1(new_n7702_), .A2(new_n4701_), .B(new_n7704_), .ZN(new_n7705_));
  AOI21_X1   g05000(.A1(new_n7697_), .A2(new_n7701_), .B(new_n7705_), .ZN(new_n7706_));
  NOR2_X1    g05001(.A1(new_n7262_), .A2(new_n5325_), .ZN(new_n7707_));
  NOR4_X1    g05002(.A1(new_n7695_), .A2(pi0299), .A3(new_n7706_), .A4(new_n7707_), .ZN(new_n7708_));
  NAND2_X1   g05003(.A1(new_n2545_), .A2(new_n5987_), .ZN(new_n7709_));
  OAI21_X1   g05004(.A1(new_n6047_), .A2(new_n4701_), .B(new_n7166_), .ZN(new_n7710_));
  NOR2_X1    g05005(.A1(new_n7710_), .A2(new_n7634_), .ZN(new_n7711_));
  INV_X1     g05006(.I(new_n7711_), .ZN(new_n7712_));
  NAND3_X1   g05007(.A1(new_n7171_), .A2(new_n4701_), .A3(new_n7170_), .ZN(new_n7713_));
  AOI21_X1   g05008(.A1(new_n7639_), .A2(new_n7713_), .B(new_n7712_), .ZN(new_n7714_));
  NOR3_X1    g05009(.A1(new_n7711_), .A2(pi0155), .A3(new_n7713_), .ZN(new_n7715_));
  NOR4_X1    g05010(.A1(new_n7714_), .A2(pi0038), .A3(new_n2587_), .A4(new_n7715_), .ZN(new_n7716_));
  OAI21_X1   g05011(.A1(new_n7155_), .A2(pi0144), .B(new_n7622_), .ZN(new_n7717_));
  AOI21_X1   g05012(.A1(new_n7157_), .A2(pi0144), .B(new_n7717_), .ZN(new_n7718_));
  NAND2_X1   g05013(.A1(new_n7163_), .A2(new_n7504_), .ZN(new_n7719_));
  NAND2_X1   g05014(.A1(new_n7719_), .A2(new_n7615_), .ZN(new_n7720_));
  OAI21_X1   g05015(.A1(new_n7718_), .A2(new_n7720_), .B(new_n5987_), .ZN(new_n7721_));
  NAND2_X1   g05016(.A1(new_n7721_), .A2(new_n3172_), .ZN(new_n7722_));
  NOR2_X1    g05017(.A1(new_n7716_), .A2(new_n7722_), .ZN(new_n7723_));
  OAI22_X1   g05018(.A1(new_n7708_), .A2(new_n7709_), .B1(new_n7723_), .B2(new_n3154_), .ZN(new_n7724_));
  AOI21_X1   g05019(.A1(new_n7724_), .A2(new_n3173_), .B(new_n7353_), .ZN(new_n7725_));
  INV_X1     g05020(.I(new_n7353_), .ZN(new_n7726_));
  NOR2_X1    g05021(.A1(new_n7359_), .A2(new_n2621_), .ZN(new_n7727_));
  AOI21_X1   g05022(.A1(new_n7726_), .A2(new_n7727_), .B(new_n3177_), .ZN(new_n7728_));
  NOR4_X1    g05023(.A1(new_n7728_), .A2(pi0075), .A3(pi0092), .A4(new_n7354_), .ZN(new_n7735_));
  OAI21_X1   g05024(.A1(new_n7725_), .A2(pi0087), .B(new_n7735_), .ZN(new_n7736_));
  NOR2_X1    g05025(.A1(new_n7363_), .A2(pi0054), .ZN(new_n7737_));
  AOI21_X1   g05026(.A1(new_n7736_), .A2(new_n7737_), .B(new_n7685_), .ZN(new_n7738_));
  INV_X1     g05027(.I(new_n7290_), .ZN(new_n7739_));
  NOR4_X1    g05028(.A1(new_n7178_), .A2(pi0092), .A3(new_n7325_), .A4(new_n7739_), .ZN(new_n7740_));
  NAND2_X1   g05029(.A1(new_n5110_), .A2(new_n7740_), .ZN(new_n7741_));
  AOI21_X1   g05030(.A1(new_n7741_), .A2(new_n7665_), .B(new_n7048_), .ZN(new_n7742_));
  NOR3_X1    g05031(.A1(new_n7050_), .A2(new_n3214_), .A3(new_n7334_), .ZN(new_n7743_));
  NOR3_X1    g05032(.A1(new_n7333_), .A2(pi0074), .A3(new_n7743_), .ZN(new_n7744_));
  OAI21_X1   g05033(.A1(new_n7742_), .A2(new_n3214_), .B(new_n7744_), .ZN(new_n7745_));
  NAND4_X1   g05034(.A1(new_n7745_), .A2(new_n3503_), .A3(new_n7673_), .A4(new_n7679_), .ZN(new_n7746_));
  OAI21_X1   g05035(.A1(new_n7738_), .A2(new_n7746_), .B(new_n7338_), .ZN(new_n7747_));
  INV_X1     g05036(.I(pi0118), .ZN(new_n7748_));
  NAND2_X1   g05037(.A1(new_n7315_), .A2(new_n7748_), .ZN(new_n7749_));
  AOI21_X1   g05038(.A1(new_n7749_), .A2(new_n7316_), .B(pi0034), .ZN(new_n7750_));
  NOR2_X1    g05039(.A1(pi0033), .A2(pi0954), .ZN(new_n7751_));
  NOR4_X1    g05040(.A1(new_n7684_), .A2(new_n7747_), .A3(new_n7750_), .A4(new_n7751_), .ZN(new_n7752_));
  AOI21_X1   g05041(.A1(new_n7747_), .A2(pi0034), .B(new_n7751_), .ZN(new_n7753_));
  OAI21_X1   g05042(.A1(new_n7684_), .A2(new_n7314_), .B(new_n7753_), .ZN(new_n7754_));
  NOR2_X1    g05043(.A1(new_n7752_), .A2(new_n7754_), .ZN(po0192));
  INV_X1     g05044(.I(new_n2959_), .ZN(new_n7756_));
  NOR2_X1    g05045(.A1(new_n7756_), .A2(new_n2958_), .ZN(new_n7757_));
  NOR2_X1    g05046(.A1(new_n7757_), .A2(new_n6005_), .ZN(new_n7758_));
  NAND2_X1   g05047(.A1(new_n7758_), .A2(pi0683), .ZN(new_n7759_));
  NAND3_X1   g05048(.A1(po1057), .A2(pi0252), .A3(new_n7759_), .ZN(new_n7760_));
  NOR2_X1    g05049(.A1(new_n6973_), .A2(new_n5163_), .ZN(new_n7761_));
  AOI22_X1   g05050(.A1(new_n5983_), .A2(pi0146), .B1(pi0142), .B2(new_n5984_), .ZN(new_n7762_));
  NAND2_X1   g05051(.A1(new_n7760_), .A2(new_n7762_), .ZN(new_n7763_));
  NAND2_X1   g05052(.A1(new_n7763_), .A2(new_n5986_), .ZN(new_n7764_));
  NOR2_X1    g05053(.A1(new_n7760_), .A2(new_n5988_), .ZN(new_n7765_));
  AOI21_X1   g05054(.A1(new_n2436_), .A2(pi0252), .B(new_n7765_), .ZN(new_n7766_));
  AOI22_X1   g05055(.A1(new_n7766_), .A2(new_n7764_), .B1(new_n7760_), .B2(new_n7761_), .ZN(new_n7767_));
  AOI21_X1   g05056(.A1(new_n7030_), .A2(pi0137), .B(new_n7032_), .ZN(new_n7768_));
  OAI21_X1   g05057(.A1(new_n7767_), .A2(new_n7033_), .B(new_n7768_), .ZN(new_n7769_));
  NAND3_X1   g05058(.A1(new_n5068_), .A2(pi0058), .A3(new_n2839_), .ZN(new_n7770_));
  NAND3_X1   g05059(.A1(new_n5059_), .A2(new_n2841_), .A3(new_n7770_), .ZN(new_n7771_));
  NAND2_X1   g05060(.A1(new_n7771_), .A2(new_n2876_), .ZN(new_n7772_));
  AOI21_X1   g05061(.A1(new_n2649_), .A2(new_n7017_), .B(new_n7772_), .ZN(new_n7773_));
  NOR2_X1    g05062(.A1(new_n7772_), .A2(new_n5081_), .ZN(new_n7774_));
  AOI21_X1   g05063(.A1(new_n2904_), .A2(pi0035), .B(new_n7022_), .ZN(new_n7775_));
  INV_X1     g05064(.I(new_n7775_), .ZN(new_n7776_));
  NAND2_X1   g05065(.A1(new_n5080_), .A2(new_n2436_), .ZN(new_n7777_));
  NAND4_X1   g05066(.A1(new_n6010_), .A2(new_n2921_), .A3(new_n6844_), .A4(new_n7777_), .ZN(new_n7778_));
  NOR2_X1    g05067(.A1(po0740), .A2(pi0122), .ZN(new_n7779_));
  NAND3_X1   g05068(.A1(new_n7779_), .A2(new_n6538_), .A3(new_n7777_), .ZN(new_n7780_));
  NAND3_X1   g05069(.A1(new_n7778_), .A2(new_n7780_), .A3(new_n2484_), .ZN(new_n7781_));
  NOR4_X1    g05070(.A1(new_n7776_), .A2(new_n7773_), .A3(new_n7774_), .A4(new_n7781_), .ZN(new_n7782_));
  AOI21_X1   g05071(.A1(new_n2876_), .A2(new_n7771_), .B(new_n7776_), .ZN(new_n7783_));
  NOR2_X1    g05072(.A1(new_n7783_), .A2(new_n2859_), .ZN(new_n7784_));
  NAND2_X1   g05073(.A1(new_n2484_), .A2(pi1082), .ZN(new_n7785_));
  OAI21_X1   g05074(.A1(new_n7784_), .A2(new_n7785_), .B(new_n3172_), .ZN(new_n7786_));
  NOR2_X1    g05075(.A1(new_n7786_), .A2(new_n7782_), .ZN(new_n7787_));
  INV_X1     g05076(.I(new_n5949_), .ZN(new_n7788_));
  NAND4_X1   g05077(.A1(new_n7788_), .A2(pi0032), .A3(new_n2841_), .A4(new_n6991_), .ZN(new_n7789_));
  NAND2_X1   g05078(.A1(new_n7783_), .A2(new_n2632_), .ZN(new_n7790_));
  NAND2_X1   g05079(.A1(new_n5080_), .A2(new_n2437_), .ZN(new_n7791_));
  AOI21_X1   g05080(.A1(new_n7790_), .A2(new_n7789_), .B(new_n7791_), .ZN(new_n7792_));
  INV_X1     g05081(.I(new_n6971_), .ZN(new_n7793_));
  OAI21_X1   g05082(.A1(new_n7793_), .A2(pi0038), .B(new_n5904_), .ZN(new_n7794_));
  OAI21_X1   g05083(.A1(new_n7787_), .A2(new_n7792_), .B(new_n7794_), .ZN(new_n7795_));
  AOI21_X1   g05084(.A1(new_n7795_), .A2(new_n7769_), .B(new_n2535_), .ZN(new_n7796_));
  INV_X1     g05085(.I(new_n6982_), .ZN(new_n7797_));
  OAI21_X1   g05086(.A1(new_n6976_), .A2(po0840), .B(new_n2436_), .ZN(new_n7798_));
  NAND4_X1   g05087(.A1(new_n6971_), .A2(new_n6974_), .A3(new_n7797_), .A4(new_n7798_), .ZN(new_n7799_));
  NAND2_X1   g05088(.A1(new_n7799_), .A2(new_n3203_), .ZN(new_n7800_));
  AOI21_X1   g05089(.A1(new_n5895_), .A2(new_n3203_), .B(pi0054), .ZN(new_n7801_));
  NAND2_X1   g05090(.A1(new_n5878_), .A2(new_n7801_), .ZN(new_n7802_));
  NOR2_X1    g05091(.A1(new_n3503_), .A2(new_n6963_), .ZN(new_n7803_));
  AOI21_X1   g05092(.A1(new_n7802_), .A2(new_n7803_), .B(pi0054), .ZN(new_n7804_));
  OAI21_X1   g05093(.A1(new_n7796_), .A2(new_n7800_), .B(new_n7804_), .ZN(new_n7805_));
  NOR3_X1    g05094(.A1(new_n7793_), .A2(new_n3503_), .A3(new_n3234_), .ZN(new_n7806_));
  INV_X1     g05095(.I(new_n7806_), .ZN(new_n7807_));
  NOR2_X1    g05096(.A1(new_n7807_), .A2(pi0055), .ZN(new_n7808_));
  INV_X1     g05097(.I(new_n7808_), .ZN(new_n7809_));
  MUX2_X1    g05098(.I0(new_n7809_), .I1(new_n7805_), .S(new_n5205_), .Z(new_n7810_));
  NOR2_X1    g05099(.A1(new_n7810_), .A2(pi0057), .ZN(po0193));
  NAND3_X1   g05100(.A1(new_n2777_), .A2(new_n2784_), .A3(new_n2775_), .ZN(new_n7812_));
  NOR4_X1    g05101(.A1(new_n7074_), .A2(new_n7000_), .A3(new_n7008_), .A4(pi0065), .ZN(new_n7813_));
  NOR3_X1    g05102(.A1(pi0069), .A2(pi0071), .A3(pi0103), .ZN(new_n7814_));
  NAND4_X1   g05103(.A1(new_n7813_), .A2(pi0036), .A3(new_n2768_), .A4(new_n7814_), .ZN(new_n7815_));
  NOR2_X1    g05104(.A1(new_n7812_), .A2(new_n7815_), .ZN(new_n7816_));
  INV_X1     g05105(.I(new_n7816_), .ZN(new_n7817_));
  NOR2_X1    g05106(.A1(new_n2890_), .A2(new_n2687_), .ZN(new_n7818_));
  INV_X1     g05107(.I(new_n7818_), .ZN(new_n7819_));
  NOR2_X1    g05108(.A1(new_n7817_), .A2(new_n7819_), .ZN(new_n7820_));
  AOI21_X1   g05109(.A1(new_n7368_), .A2(new_n6019_), .B(new_n7820_), .ZN(new_n7821_));
  NOR2_X1    g05110(.A1(po1038), .A2(new_n2539_), .ZN(new_n7822_));
  INV_X1     g05111(.I(new_n7822_), .ZN(new_n7823_));
  NOR2_X1    g05112(.A1(new_n7823_), .A2(new_n3325_), .ZN(new_n7824_));
  INV_X1     g05113(.I(new_n7824_), .ZN(new_n7825_));
  NOR2_X1    g05114(.A1(new_n2515_), .A2(new_n2650_), .ZN(new_n7826_));
  NAND2_X1   g05115(.A1(new_n5082_), .A2(new_n7826_), .ZN(new_n7827_));
  NOR2_X1    g05116(.A1(new_n7825_), .A2(new_n7827_), .ZN(new_n7828_));
  INV_X1     g05117(.I(new_n7828_), .ZN(new_n7829_));
  NOR3_X1    g05118(.A1(new_n7821_), .A2(new_n5943_), .A3(new_n7829_), .ZN(po0194));
  INV_X1     g05119(.I(new_n5894_), .ZN(po0195));
  NOR2_X1    g05120(.A1(po1038), .A2(new_n3232_), .ZN(new_n7832_));
  INV_X1     g05121(.I(new_n7832_), .ZN(new_n7833_));
  INV_X1     g05122(.I(new_n7213_), .ZN(new_n7834_));
  INV_X1     g05123(.I(pi0049), .ZN(new_n7835_));
  NAND2_X1   g05124(.A1(new_n2732_), .A2(new_n7835_), .ZN(new_n7836_));
  NOR2_X1    g05125(.A1(new_n2758_), .A2(new_n7836_), .ZN(new_n7837_));
  NAND4_X1   g05126(.A1(new_n7214_), .A2(new_n2734_), .A3(new_n2806_), .A4(pi0089), .ZN(new_n7838_));
  NOR2_X1    g05127(.A1(new_n7837_), .A2(new_n7838_), .ZN(new_n7839_));
  NOR4_X1    g05128(.A1(new_n7000_), .A2(new_n2442_), .A3(pi0071), .A4(pi0104), .ZN(new_n7840_));
  NAND3_X1   g05129(.A1(new_n7839_), .A2(new_n7834_), .A3(new_n7840_), .ZN(new_n7841_));
  OAI21_X1   g05130(.A1(new_n7841_), .A2(new_n2563_), .B(new_n2454_), .ZN(new_n7842_));
  INV_X1     g05131(.I(new_n2662_), .ZN(new_n7843_));
  NOR2_X1    g05132(.A1(new_n7843_), .A2(new_n2474_), .ZN(new_n7844_));
  INV_X1     g05133(.I(new_n7844_), .ZN(new_n7845_));
  NOR3_X1    g05134(.A1(new_n7845_), .A2(new_n2509_), .A3(new_n2515_), .ZN(new_n7846_));
  INV_X1     g05135(.I(new_n7846_), .ZN(new_n7847_));
  NOR2_X1    g05136(.A1(new_n7847_), .A2(new_n2507_), .ZN(new_n7848_));
  NOR4_X1    g05137(.A1(new_n2464_), .A2(pi0039), .A3(pi0081), .A4(pi0841), .ZN(new_n7849_));
  NAND4_X1   g05138(.A1(new_n7848_), .A2(new_n2727_), .A3(new_n7842_), .A4(new_n7849_), .ZN(new_n7850_));
  NOR4_X1    g05139(.A1(new_n2654_), .A2(new_n5895_), .A3(pi0039), .A4(new_n2485_), .ZN(new_n7851_));
  INV_X1     g05140(.I(new_n7851_), .ZN(new_n7852_));
  MUX2_X1    g05141(.I0(new_n7852_), .I1(new_n7850_), .S(new_n3172_), .Z(new_n7853_));
  NOR2_X1    g05142(.A1(new_n7853_), .A2(new_n7833_), .ZN(po0196));
  NOR2_X1    g05143(.A1(new_n7833_), .A2(pi0038), .ZN(new_n7855_));
  INV_X1     g05144(.I(new_n7855_), .ZN(new_n7856_));
  OAI21_X1   g05145(.A1(pi0252), .A2(pi1001), .B(new_n5119_), .ZN(new_n7857_));
  INV_X1     g05146(.I(pi0984), .ZN(new_n7858_));
  NAND2_X1   g05147(.A1(new_n2955_), .A2(new_n7858_), .ZN(new_n7859_));
  NAND3_X1   g05148(.A1(new_n7857_), .A2(new_n7859_), .A3(pi0835), .ZN(new_n7860_));
  INV_X1     g05149(.I(new_n7860_), .ZN(new_n7861_));
  NOR2_X1    g05150(.A1(new_n5117_), .A2(new_n7861_), .ZN(new_n7862_));
  AOI21_X1   g05151(.A1(new_n5143_), .A2(new_n7862_), .B(new_n5361_), .ZN(new_n7863_));
  INV_X1     g05152(.I(new_n7863_), .ZN(new_n7864_));
  AOI21_X1   g05153(.A1(new_n6446_), .A2(new_n7862_), .B(new_n5361_), .ZN(new_n7865_));
  INV_X1     g05154(.I(new_n7865_), .ZN(new_n7866_));
  AOI21_X1   g05155(.A1(new_n6460_), .A2(new_n7866_), .B(new_n7864_), .ZN(new_n7867_));
  NOR3_X1    g05156(.A1(new_n7866_), .A2(new_n5141_), .A3(new_n7863_), .ZN(new_n7868_));
  NOR3_X1    g05157(.A1(new_n7867_), .A2(new_n7868_), .A3(pi0299), .ZN(new_n7869_));
  AOI21_X1   g05158(.A1(pi1093), .A2(new_n7862_), .B(new_n5361_), .ZN(new_n7870_));
  AOI21_X1   g05159(.A1(new_n2604_), .A2(new_n7870_), .B(new_n7869_), .ZN(new_n7871_));
  OAI21_X1   g05160(.A1(new_n7863_), .A2(new_n6445_), .B(new_n2587_), .ZN(new_n7872_));
  AOI21_X1   g05161(.A1(new_n6445_), .A2(new_n7866_), .B(new_n7872_), .ZN(new_n7873_));
  NAND2_X1   g05162(.A1(new_n7870_), .A2(new_n2566_), .ZN(new_n7874_));
  NAND2_X1   g05163(.A1(new_n7873_), .A2(new_n7874_), .ZN(new_n7875_));
  INV_X1     g05164(.I(pi0786), .ZN(new_n7876_));
  NOR2_X1    g05165(.A1(new_n7876_), .A2(pi1082), .ZN(new_n7877_));
  INV_X1     g05166(.I(new_n7877_), .ZN(new_n7878_));
  NOR2_X1    g05167(.A1(new_n5145_), .A2(new_n3294_), .ZN(new_n7879_));
  INV_X1     g05168(.I(new_n4899_), .ZN(new_n7880_));
  NOR2_X1    g05169(.A1(new_n5866_), .A2(new_n7880_), .ZN(new_n7881_));
  NOR4_X1    g05170(.A1(new_n7881_), .A2(new_n5943_), .A3(new_n7878_), .A4(new_n7879_), .ZN(new_n7882_));
  AOI21_X1   g05171(.A1(new_n7882_), .A2(new_n5362_), .B(new_n7877_), .ZN(new_n7883_));
  NAND2_X1   g05172(.A1(new_n7875_), .A2(new_n7883_), .ZN(new_n7884_));
  OAI21_X1   g05173(.A1(new_n7871_), .A2(new_n7884_), .B(pi0039), .ZN(new_n7885_));
  INV_X1     g05174(.I(new_n2887_), .ZN(new_n7886_));
  NOR2_X1    g05175(.A1(new_n5063_), .A2(new_n7886_), .ZN(new_n7887_));
  INV_X1     g05176(.I(new_n2449_), .ZN(new_n7888_));
  INV_X1     g05177(.I(pi0082), .ZN(new_n7889_));
  NAND4_X1   g05178(.A1(new_n2757_), .A2(new_n2728_), .A3(new_n7889_), .A4(pi0048), .ZN(new_n7890_));
  NOR4_X1    g05179(.A1(new_n7890_), .A2(new_n7002_), .A3(pi0111), .A4(new_n7888_), .ZN(new_n7891_));
  NOR4_X1    g05180(.A1(pi0064), .A2(pi0066), .A3(pi0081), .A4(pi0084), .ZN(new_n7892_));
  NOR3_X1    g05181(.A1(new_n7892_), .A2(pi0065), .A3(pi0069), .ZN(new_n7893_));
  INV_X1     g05182(.I(new_n7840_), .ZN(new_n7894_));
  NOR4_X1    g05183(.A1(new_n7894_), .A2(new_n7008_), .A3(new_n2769_), .A4(new_n7836_), .ZN(new_n7895_));
  NAND3_X1   g05184(.A1(new_n7895_), .A2(new_n7891_), .A3(new_n7893_), .ZN(new_n7896_));
  INV_X1     g05185(.I(new_n7896_), .ZN(new_n7897_));
  NOR3_X1    g05186(.A1(new_n7210_), .A2(new_n2683_), .A3(pi0841), .ZN(new_n7898_));
  NAND4_X1   g05187(.A1(new_n7887_), .A2(new_n2680_), .A3(new_n7897_), .A4(new_n7898_), .ZN(new_n7899_));
  OAI21_X1   g05188(.A1(po0740), .A2(pi0986), .B(pi0252), .ZN(new_n7900_));
  AND2_X2    g05189(.A1(new_n7900_), .A2(pi0314), .Z(new_n7901_));
  NAND2_X1   g05190(.A1(new_n5071_), .A2(new_n7901_), .ZN(new_n7902_));
  NAND4_X1   g05191(.A1(new_n2686_), .A2(new_n2680_), .A3(pi0108), .A4(new_n2887_), .ZN(new_n7903_));
  OR4_X2     g05192(.A1(pi0102), .A2(new_n2459_), .A3(new_n7008_), .A4(new_n7903_), .Z(new_n7904_));
  NAND4_X1   g05193(.A1(new_n7899_), .A2(new_n2661_), .A3(new_n7902_), .A4(new_n7904_), .ZN(new_n7905_));
  NOR3_X1    g05194(.A1(new_n7896_), .A2(pi0047), .A3(pi0841), .ZN(new_n7906_));
  OAI21_X1   g05195(.A1(new_n2661_), .A2(new_n2635_), .B(new_n7906_), .ZN(new_n7907_));
  NOR3_X1    g05196(.A1(new_n7906_), .A2(new_n2661_), .A3(new_n2635_), .ZN(new_n7908_));
  NOR4_X1    g05197(.A1(new_n7908_), .A2(new_n7843_), .A3(new_n6986_), .A4(new_n7901_), .ZN(new_n7909_));
  AOI21_X1   g05198(.A1(new_n7909_), .A2(new_n7907_), .B(new_n2650_), .ZN(new_n7910_));
  AOI21_X1   g05199(.A1(new_n7905_), .A2(new_n7910_), .B(pi0035), .ZN(new_n7911_));
  NAND2_X1   g05200(.A1(new_n5970_), .A2(new_n2876_), .ZN(new_n7912_));
  NAND3_X1   g05201(.A1(new_n7912_), .A2(new_n2506_), .A3(new_n2512_), .ZN(new_n7913_));
  NOR3_X1    g05202(.A1(new_n5242_), .A2(new_n2632_), .A3(new_n5080_), .ZN(new_n7914_));
  NOR3_X1    g05203(.A1(new_n7914_), .A2(pi0039), .A3(pi0095), .ZN(new_n7915_));
  OAI21_X1   g05204(.A1(new_n7911_), .A2(new_n7913_), .B(new_n7915_), .ZN(new_n7916_));
  AOI21_X1   g05205(.A1(new_n7885_), .A2(new_n7916_), .B(new_n7856_), .ZN(po0197));
  NOR2_X1    g05206(.A1(new_n3365_), .A2(new_n7194_), .ZN(new_n7918_));
  NOR4_X1    g05207(.A1(new_n2480_), .A2(pi0081), .A3(pi0093), .A4(new_n2462_), .ZN(new_n7919_));
  NAND2_X1   g05208(.A1(new_n7919_), .A2(new_n7069_), .ZN(new_n7920_));
  NOR4_X1    g05209(.A1(new_n7845_), .A2(new_n2699_), .A3(new_n5083_), .A4(new_n7920_), .ZN(new_n7921_));
  OAI21_X1   g05210(.A1(pi0040), .A2(new_n7921_), .B(new_n7918_), .ZN(new_n7922_));
  NAND2_X1   g05211(.A1(new_n7922_), .A2(pi1082), .ZN(new_n7923_));
  NAND3_X1   g05212(.A1(new_n7921_), .A2(pi1082), .A3(new_n2514_), .ZN(new_n7924_));
  AOI21_X1   g05213(.A1(new_n7923_), .A2(new_n7924_), .B(new_n7825_), .ZN(po0198));
  NOR2_X1    g05214(.A1(new_n3154_), .A2(new_n5987_), .ZN(new_n7926_));
  INV_X1     g05215(.I(new_n7926_), .ZN(new_n7927_));
  NOR2_X1    g05216(.A1(new_n5109_), .A2(pi0166), .ZN(new_n7928_));
  NAND3_X1   g05217(.A1(new_n7928_), .A2(new_n3250_), .A3(pi0161), .ZN(new_n7929_));
  NOR2_X1    g05218(.A1(new_n7929_), .A2(new_n7927_), .ZN(new_n7930_));
  INV_X1     g05219(.I(pi0041), .ZN(new_n7931_));
  NAND4_X1   g05220(.A1(new_n6845_), .A2(pi0039), .A3(new_n7931_), .A4(new_n2861_), .ZN(new_n7932_));
  INV_X1     g05221(.I(pi0044), .ZN(new_n7933_));
  NOR2_X1    g05222(.A1(new_n7933_), .A2(pi0072), .ZN(new_n7934_));
  INV_X1     g05223(.I(new_n5976_), .ZN(new_n7935_));
  NOR2_X1    g05224(.A1(new_n5971_), .A2(new_n2515_), .ZN(new_n7936_));
  OAI21_X1   g05225(.A1(pi0072), .A2(new_n5948_), .B(new_n7936_), .ZN(new_n7937_));
  NOR2_X1    g05226(.A1(new_n5969_), .A2(new_n7937_), .ZN(new_n7938_));
  NAND2_X1   g05227(.A1(new_n5948_), .A2(new_n2861_), .ZN(new_n7939_));
  OAI22_X1   g05228(.A1(new_n7938_), .A2(pi1093), .B1(new_n7935_), .B2(new_n7939_), .ZN(new_n7940_));
  NOR2_X1    g05229(.A1(new_n5962_), .A2(new_n2935_), .ZN(new_n7941_));
  AOI21_X1   g05230(.A1(new_n7941_), .A2(new_n2934_), .B(new_n6019_), .ZN(new_n7942_));
  OAI21_X1   g05231(.A1(new_n7942_), .A2(new_n2480_), .B(new_n5950_), .ZN(new_n7943_));
  AOI21_X1   g05232(.A1(new_n7943_), .A2(new_n6017_), .B(new_n2658_), .ZN(new_n7944_));
  NAND4_X1   g05233(.A1(new_n2500_), .A2(new_n2441_), .A3(new_n2475_), .A4(new_n2481_), .ZN(new_n7945_));
  NOR2_X1    g05234(.A1(new_n7945_), .A2(new_n2658_), .ZN(new_n7946_));
  NOR3_X1    g05235(.A1(new_n7944_), .A2(pi0096), .A3(new_n7946_), .ZN(new_n7947_));
  NAND4_X1   g05236(.A1(new_n7947_), .A2(new_n2861_), .A3(new_n5947_), .A4(new_n7936_), .ZN(new_n7948_));
  OAI21_X1   g05237(.A1(new_n5947_), .A2(new_n5976_), .B(new_n7948_), .ZN(new_n7949_));
  NAND3_X1   g05238(.A1(new_n7949_), .A2(new_n2861_), .A3(new_n2924_), .ZN(new_n7950_));
  NAND2_X1   g05239(.A1(new_n7950_), .A2(new_n7940_), .ZN(new_n7951_));
  AOI21_X1   g05240(.A1(new_n7951_), .A2(new_n7933_), .B(new_n7934_), .ZN(new_n7952_));
  NOR3_X1    g05241(.A1(new_n7952_), .A2(new_n2861_), .A3(pi0101), .ZN(new_n7953_));
  INV_X1     g05242(.I(pi0101), .ZN(new_n7954_));
  AOI21_X1   g05243(.A1(new_n7952_), .A2(new_n7954_), .B(pi0072), .ZN(new_n7955_));
  NOR3_X1    g05244(.A1(new_n7953_), .A2(new_n7955_), .A3(pi0041), .ZN(new_n7956_));
  INV_X1     g05245(.I(new_n7956_), .ZN(new_n7957_));
  NOR2_X1    g05246(.A1(new_n5976_), .A2(new_n5947_), .ZN(new_n7958_));
  NOR3_X1    g05247(.A1(new_n5974_), .A2(new_n7958_), .A3(pi1093), .ZN(new_n7959_));
  NOR2_X1    g05248(.A1(new_n7959_), .A2(pi0044), .ZN(new_n7960_));
  NAND2_X1   g05249(.A1(new_n7949_), .A2(pi1093), .ZN(new_n7961_));
  NAND2_X1   g05250(.A1(new_n7961_), .A2(new_n7960_), .ZN(new_n7962_));
  NOR2_X1    g05251(.A1(new_n7962_), .A2(pi0101), .ZN(new_n7963_));
  INV_X1     g05252(.I(new_n7963_), .ZN(new_n7964_));
  NOR4_X1    g05253(.A1(new_n7957_), .A2(pi0041), .A3(new_n2921_), .A4(new_n7964_), .ZN(new_n7965_));
  NAND3_X1   g05254(.A1(new_n7940_), .A2(new_n2861_), .A3(new_n5976_), .ZN(new_n7966_));
  INV_X1     g05255(.I(new_n7966_), .ZN(new_n7967_));
  AOI21_X1   g05256(.A1(new_n7967_), .A2(new_n7933_), .B(new_n7934_), .ZN(new_n7968_));
  INV_X1     g05257(.I(new_n7968_), .ZN(new_n7969_));
  NAND3_X1   g05258(.A1(new_n7969_), .A2(pi0072), .A3(new_n7954_), .ZN(new_n7970_));
  OAI21_X1   g05259(.A1(new_n7969_), .A2(pi0101), .B(new_n2861_), .ZN(new_n7971_));
  NAND3_X1   g05260(.A1(new_n7971_), .A2(new_n7970_), .A3(new_n7931_), .ZN(new_n7972_));
  INV_X1     g05261(.I(new_n7972_), .ZN(new_n7973_));
  OAI21_X1   g05262(.A1(new_n2924_), .A2(new_n7935_), .B(new_n7960_), .ZN(new_n7974_));
  NOR2_X1    g05263(.A1(new_n7974_), .A2(pi0101), .ZN(new_n7975_));
  NAND2_X1   g05264(.A1(new_n7975_), .A2(new_n7931_), .ZN(new_n7976_));
  NAND4_X1   g05265(.A1(new_n7973_), .A2(pi0228), .A3(new_n2922_), .A4(new_n7976_), .ZN(new_n7977_));
  NOR2_X1    g05266(.A1(new_n2831_), .A2(new_n2886_), .ZN(new_n7978_));
  AOI21_X1   g05267(.A1(new_n2820_), .A2(new_n7978_), .B(pi0110), .ZN(new_n7979_));
  INV_X1     g05268(.I(pi0480), .ZN(new_n7980_));
  NAND4_X1   g05269(.A1(new_n2651_), .A2(new_n2661_), .A3(new_n7980_), .A4(pi0949), .ZN(new_n7981_));
  NOR4_X1    g05270(.A1(new_n7979_), .A2(new_n6986_), .A3(new_n2835_), .A4(new_n7981_), .ZN(new_n7982_));
  INV_X1     g05271(.I(pi0959), .ZN(new_n7983_));
  NAND2_X1   g05272(.A1(new_n2820_), .A2(new_n2889_), .ZN(new_n7984_));
  NOR2_X1    g05273(.A1(new_n7984_), .A2(new_n2652_), .ZN(new_n7985_));
  OAI21_X1   g05274(.A1(new_n7980_), .A2(pi0949), .B(new_n7985_), .ZN(new_n7986_));
  NAND3_X1   g05275(.A1(new_n7986_), .A2(pi0901), .A3(new_n7983_), .ZN(new_n7987_));
  INV_X1     g05276(.I(pi0949), .ZN(new_n7988_));
  NOR4_X1    g05277(.A1(new_n2637_), .A2(pi0047), .A3(pi0109), .A4(new_n6986_), .ZN(new_n7989_));
  NAND2_X1   g05278(.A1(new_n7989_), .A2(pi0110), .ZN(new_n7990_));
  NOR4_X1    g05279(.A1(new_n7990_), .A2(pi0480), .A3(new_n7988_), .A4(new_n2652_), .ZN(new_n7991_));
  AOI21_X1   g05280(.A1(pi0901), .A2(new_n7983_), .B(new_n7991_), .ZN(new_n7992_));
  NOR4_X1    g05281(.A1(new_n7992_), .A2(pi0250), .A3(new_n3181_), .A4(new_n2515_), .ZN(new_n7993_));
  OAI21_X1   g05282(.A1(new_n7987_), .A2(new_n7982_), .B(new_n7993_), .ZN(new_n7994_));
  AOI21_X1   g05283(.A1(pi0250), .A2(new_n3181_), .B(new_n2515_), .ZN(new_n7995_));
  NAND2_X1   g05284(.A1(new_n7991_), .A2(new_n7995_), .ZN(new_n7996_));
  AND3_X2    g05285(.A1(new_n7994_), .A2(new_n2861_), .A3(new_n7996_), .Z(new_n7997_));
  AOI21_X1   g05286(.A1(new_n7997_), .A2(new_n7933_), .B(new_n7934_), .ZN(new_n7998_));
  NOR3_X1    g05287(.A1(new_n7998_), .A2(new_n2861_), .A3(pi0101), .ZN(new_n7999_));
  AOI21_X1   g05288(.A1(new_n7998_), .A2(new_n7954_), .B(pi0072), .ZN(new_n8000_));
  NOR3_X1    g05289(.A1(new_n7999_), .A2(new_n8000_), .A3(pi0041), .ZN(new_n8001_));
  NOR2_X1    g05290(.A1(new_n7990_), .A2(new_n7827_), .ZN(new_n8002_));
  NOR4_X1    g05291(.A1(new_n5180_), .A2(pi0252), .A3(pi0480), .A4(pi0949), .ZN(new_n8003_));
  NOR2_X1    g05292(.A1(new_n7994_), .A2(pi0072), .ZN(new_n8004_));
  AOI21_X1   g05293(.A1(new_n8002_), .A2(new_n8003_), .B(new_n8004_), .ZN(new_n8005_));
  NAND3_X1   g05294(.A1(new_n8005_), .A2(new_n7933_), .A3(new_n7954_), .ZN(new_n8006_));
  NAND2_X1   g05295(.A1(new_n8006_), .A2(pi0041), .ZN(new_n8007_));
  NAND2_X1   g05296(.A1(new_n8001_), .A2(new_n8007_), .ZN(new_n8008_));
  AOI21_X1   g05297(.A1(new_n8008_), .A2(new_n2523_), .B(pi0039), .ZN(new_n8009_));
  OAI21_X1   g05298(.A1(new_n7965_), .A2(new_n7977_), .B(new_n8009_), .ZN(new_n8010_));
  NOR2_X1    g05299(.A1(new_n5109_), .A2(pi0189), .ZN(new_n8011_));
  INV_X1     g05300(.I(new_n8011_), .ZN(new_n8012_));
  NOR2_X1    g05301(.A1(new_n8012_), .A2(new_n7504_), .ZN(new_n8013_));
  NAND2_X1   g05302(.A1(new_n8013_), .A2(new_n7151_), .ZN(new_n8014_));
  NAND2_X1   g05303(.A1(new_n8014_), .A2(new_n2587_), .ZN(new_n8015_));
  OAI21_X1   g05304(.A1(pi0299), .A2(new_n2605_), .B(new_n7929_), .ZN(new_n8016_));
  NAND3_X1   g05305(.A1(new_n8015_), .A2(pi0232), .A3(new_n8016_), .ZN(new_n8017_));
  INV_X1     g05306(.I(pi0287), .ZN(new_n8018_));
  NOR2_X1    g05307(.A1(new_n2491_), .A2(new_n8018_), .ZN(new_n8019_));
  OR2_X2     g05308(.A1(new_n8019_), .A2(new_n8017_), .Z(new_n8020_));
  AOI21_X1   g05309(.A1(new_n8017_), .A2(pi0072), .B(new_n3154_), .ZN(new_n8021_));
  AOI21_X1   g05310(.A1(new_n8020_), .A2(new_n8021_), .B(new_n2622_), .ZN(new_n8022_));
  NOR2_X1    g05311(.A1(pi0041), .A2(pi0072), .ZN(new_n8023_));
  INV_X1     g05312(.I(new_n8023_), .ZN(new_n8024_));
  INV_X1     g05313(.I(new_n6481_), .ZN(new_n8025_));
  NOR2_X1    g05314(.A1(new_n8025_), .A2(new_n2922_), .ZN(new_n8026_));
  AOI21_X1   g05315(.A1(new_n8026_), .A2(new_n8024_), .B(pi0039), .ZN(new_n8027_));
  NOR2_X1    g05316(.A1(new_n7954_), .A2(pi0072), .ZN(new_n8028_));
  NOR2_X1    g05317(.A1(new_n8028_), .A2(pi0041), .ZN(new_n8029_));
  NOR2_X1    g05318(.A1(new_n2654_), .A2(new_n2515_), .ZN(new_n8030_));
  INV_X1     g05319(.I(new_n8030_), .ZN(new_n8031_));
  NOR2_X1    g05320(.A1(new_n8031_), .A2(pi0044), .ZN(new_n8032_));
  AOI22_X1   g05321(.A1(new_n8032_), .A2(new_n8029_), .B1(new_n7931_), .B2(pi0072), .ZN(new_n8033_));
  AOI21_X1   g05322(.A1(new_n2861_), .A2(new_n6436_), .B(new_n8033_), .ZN(new_n8034_));
  NOR3_X1    g05323(.A1(new_n2491_), .A2(pi0044), .A3(pi0101), .ZN(new_n8035_));
  INV_X1     g05324(.I(new_n8035_), .ZN(new_n8036_));
  NOR2_X1    g05325(.A1(new_n8036_), .A2(new_n6436_), .ZN(new_n8037_));
  NOR2_X1    g05326(.A1(new_n8037_), .A2(new_n7931_), .ZN(new_n8038_));
  NAND2_X1   g05327(.A1(new_n7931_), .A2(pi0072), .ZN(new_n8039_));
  NOR2_X1    g05328(.A1(new_n5170_), .A2(pi0099), .ZN(new_n8040_));
  NAND4_X1   g05329(.A1(new_n6481_), .A2(new_n2922_), .A3(new_n8039_), .A4(new_n8040_), .ZN(new_n8041_));
  OR3_X2     g05330(.A1(new_n8034_), .A2(new_n8038_), .A3(new_n8041_), .Z(new_n8042_));
  AOI21_X1   g05331(.A1(new_n8017_), .A2(new_n2861_), .B(new_n3154_), .ZN(new_n8043_));
  INV_X1     g05332(.I(new_n8043_), .ZN(new_n8044_));
  NAND2_X1   g05333(.A1(new_n8044_), .A2(new_n5159_), .ZN(new_n8045_));
  AOI21_X1   g05334(.A1(new_n8042_), .A2(new_n8027_), .B(new_n8045_), .ZN(new_n8046_));
  NOR2_X1    g05335(.A1(new_n8023_), .A2(pi0039), .ZN(new_n8047_));
  NOR2_X1    g05336(.A1(new_n8043_), .A2(new_n8047_), .ZN(new_n8048_));
  NAND2_X1   g05337(.A1(new_n8048_), .A2(new_n3172_), .ZN(new_n8049_));
  NAND2_X1   g05338(.A1(new_n8049_), .A2(new_n3177_), .ZN(new_n8050_));
  INV_X1     g05339(.I(new_n8047_), .ZN(new_n8051_));
  OAI21_X1   g05340(.A1(new_n8051_), .A2(new_n2621_), .B(pi0087), .ZN(new_n8052_));
  INV_X1     g05341(.I(new_n8033_), .ZN(new_n8053_));
  NOR2_X1    g05342(.A1(new_n3197_), .A2(new_n2523_), .ZN(new_n8054_));
  OAI21_X1   g05343(.A1(new_n8035_), .A2(new_n7931_), .B(new_n8054_), .ZN(new_n8055_));
  OAI21_X1   g05344(.A1(new_n8053_), .A2(new_n8055_), .B(new_n8044_), .ZN(new_n8056_));
  AOI21_X1   g05345(.A1(new_n8056_), .A2(new_n8052_), .B(pi0075), .ZN(new_n8057_));
  OAI21_X1   g05346(.A1(new_n8046_), .A2(new_n8050_), .B(new_n8057_), .ZN(new_n8058_));
  AOI21_X1   g05347(.A1(new_n8010_), .A2(new_n8022_), .B(new_n8058_), .ZN(new_n8059_));
  NOR2_X1    g05348(.A1(new_n2654_), .A2(pi0024), .ZN(new_n8061_));
  NAND4_X1   g05349(.A1(new_n8061_), .A2(pi0252), .A3(new_n2514_), .A4(new_n6010_), .ZN(new_n8062_));
  NOR2_X1    g05350(.A1(new_n8062_), .A2(pi0044), .ZN(new_n8063_));
  NAND2_X1   g05351(.A1(new_n8063_), .A2(new_n8029_), .ZN(new_n8064_));
  INV_X1     g05352(.I(new_n8037_), .ZN(new_n8067_));
  NAND4_X1   g05353(.A1(new_n8044_), .A2(new_n2628_), .A3(new_n3208_), .A4(new_n8051_), .ZN(new_n8070_));
  NOR2_X1    g05354(.A1(new_n6845_), .A2(new_n5942_), .ZN(new_n8071_));
  NAND2_X1   g05355(.A1(new_n8070_), .A2(new_n8071_), .ZN(new_n8072_));
  OAI22_X1   g05356(.A1(new_n8059_), .A2(new_n8072_), .B1(new_n7930_), .B2(new_n7932_), .ZN(po0199));
  INV_X1     g05357(.I(pi0042), .ZN(new_n8074_));
  NOR2_X1    g05358(.A1(new_n8074_), .A2(pi0072), .ZN(new_n8075_));
  INV_X1     g05359(.I(pi0212), .ZN(new_n8076_));
  INV_X1     g05360(.I(pi0211), .ZN(new_n8077_));
  INV_X1     g05361(.I(pi0214), .ZN(new_n8078_));
  NOR2_X1    g05362(.A1(new_n8077_), .A2(new_n8078_), .ZN(new_n8079_));
  INV_X1     g05363(.I(new_n8079_), .ZN(new_n8080_));
  NOR2_X1    g05364(.A1(new_n8080_), .A2(new_n8076_), .ZN(new_n8081_));
  NOR2_X1    g05365(.A1(new_n8081_), .A2(pi0219), .ZN(new_n8082_));
  AOI21_X1   g05366(.A1(new_n5988_), .A2(new_n4549_), .B(pi0072), .ZN(new_n8083_));
  INV_X1     g05367(.I(new_n8083_), .ZN(new_n8084_));
  NOR2_X1    g05368(.A1(new_n8084_), .A2(new_n8082_), .ZN(new_n8085_));
  MUX2_X1    g05369(.I0(new_n8085_), .I1(new_n8075_), .S(new_n3154_), .Z(new_n8086_));
  INV_X1     g05370(.I(pi0207), .ZN(new_n8087_));
  INV_X1     g05371(.I(pi0208), .ZN(new_n8088_));
  NOR2_X1    g05372(.A1(new_n8087_), .A2(new_n8088_), .ZN(new_n8089_));
  INV_X1     g05373(.I(new_n8089_), .ZN(new_n8090_));
  NOR2_X1    g05374(.A1(new_n8011_), .A2(pi0072), .ZN(new_n8091_));
  INV_X1     g05375(.I(new_n8091_), .ZN(new_n8092_));
  AOI21_X1   g05376(.A1(new_n2861_), .A2(pi0199), .B(pi0232), .ZN(new_n8093_));
  INV_X1     g05377(.I(pi0199), .ZN(new_n8094_));
  NOR2_X1    g05378(.A1(new_n8094_), .A2(pi0232), .ZN(new_n8095_));
  OAI21_X1   g05379(.A1(new_n8093_), .A2(pi0299), .B(new_n8095_), .ZN(new_n8096_));
  NOR2_X1    g05380(.A1(new_n8092_), .A2(new_n8096_), .ZN(new_n8097_));
  INV_X1     g05381(.I(pi0200), .ZN(new_n8098_));
  NOR2_X1    g05382(.A1(new_n8098_), .A2(pi0072), .ZN(new_n8099_));
  OAI21_X1   g05383(.A1(new_n8099_), .A2(pi0232), .B(new_n2587_), .ZN(new_n8100_));
  NAND4_X1   g05384(.A1(new_n8091_), .A2(pi0200), .A3(new_n5987_), .A4(new_n8100_), .ZN(new_n8101_));
  NAND2_X1   g05385(.A1(new_n8101_), .A2(pi0039), .ZN(new_n8102_));
  NOR2_X1    g05386(.A1(new_n8102_), .A2(new_n8097_), .ZN(new_n8103_));
  NOR2_X1    g05387(.A1(new_n8075_), .A2(pi0039), .ZN(new_n8104_));
  INV_X1     g05388(.I(new_n8104_), .ZN(new_n8105_));
  NAND2_X1   g05389(.A1(new_n5942_), .A2(new_n8105_), .ZN(new_n8106_));
  OAI21_X1   g05390(.A1(new_n8103_), .A2(new_n8106_), .B(new_n8089_), .ZN(new_n8107_));
  INV_X1     g05391(.I(new_n8075_), .ZN(new_n8108_));
  INV_X1     g05392(.I(pi0116), .ZN(new_n8109_));
  NOR2_X1    g05393(.A1(new_n8109_), .A2(pi0072), .ZN(new_n8110_));
  INV_X1     g05394(.I(pi0113), .ZN(new_n8111_));
  NOR2_X1    g05395(.A1(new_n8111_), .A2(pi0072), .ZN(new_n8112_));
  INV_X1     g05396(.I(new_n8112_), .ZN(new_n8113_));
  NOR2_X1    g05397(.A1(new_n8113_), .A2(new_n5171_), .ZN(new_n8114_));
  INV_X1     g05398(.I(pi0099), .ZN(new_n8115_));
  NAND2_X1   g05399(.A1(new_n7972_), .A2(new_n8115_), .ZN(new_n8116_));
  AOI21_X1   g05400(.A1(new_n8116_), .A2(pi0113), .B(new_n8114_), .ZN(new_n8117_));
  INV_X1     g05401(.I(new_n8117_), .ZN(new_n8118_));
  AOI21_X1   g05402(.A1(new_n8118_), .A2(new_n8109_), .B(new_n8110_), .ZN(new_n8119_));
  NOR3_X1    g05403(.A1(new_n5172_), .A2(pi0113), .A3(pi0116), .ZN(new_n8120_));
  NAND2_X1   g05404(.A1(new_n7975_), .A2(new_n8120_), .ZN(new_n8121_));
  AOI21_X1   g05405(.A1(new_n8074_), .A2(new_n8121_), .B(new_n8119_), .ZN(new_n8122_));
  INV_X1     g05406(.I(new_n8119_), .ZN(new_n8123_));
  NOR3_X1    g05407(.A1(new_n8123_), .A2(pi0042), .A3(new_n8121_), .ZN(new_n8124_));
  INV_X1     g05408(.I(pi0115), .ZN(new_n8125_));
  AOI21_X1   g05409(.A1(new_n2922_), .A2(new_n8125_), .B(pi0114), .ZN(new_n8126_));
  INV_X1     g05410(.I(new_n8126_), .ZN(new_n8127_));
  NOR3_X1    g05411(.A1(new_n8124_), .A2(new_n8122_), .A3(new_n8127_), .ZN(new_n8128_));
  NOR2_X1    g05412(.A1(new_n2922_), .A2(pi0115), .ZN(new_n8129_));
  INV_X1     g05413(.I(new_n8129_), .ZN(new_n8130_));
  NAND2_X1   g05414(.A1(new_n7957_), .A2(new_n8115_), .ZN(new_n8131_));
  AOI21_X1   g05415(.A1(new_n8131_), .A2(pi0113), .B(new_n8114_), .ZN(new_n8132_));
  INV_X1     g05416(.I(new_n8132_), .ZN(new_n8133_));
  AOI21_X1   g05417(.A1(new_n8133_), .A2(new_n8109_), .B(new_n8110_), .ZN(new_n8134_));
  INV_X1     g05418(.I(new_n8134_), .ZN(new_n8135_));
  NOR2_X1    g05419(.A1(new_n8135_), .A2(pi0114), .ZN(new_n8136_));
  INV_X1     g05420(.I(new_n8136_), .ZN(new_n8137_));
  INV_X1     g05421(.I(pi0114), .ZN(new_n8138_));
  NOR2_X1    g05422(.A1(new_n8075_), .A2(new_n8138_), .ZN(new_n8139_));
  INV_X1     g05423(.I(new_n8139_), .ZN(new_n8140_));
  NOR2_X1    g05424(.A1(pi0113), .A2(pi0116), .ZN(new_n8141_));
  INV_X1     g05425(.I(new_n8141_), .ZN(new_n8142_));
  NOR3_X1    g05426(.A1(new_n7964_), .A2(new_n5172_), .A3(new_n8142_), .ZN(new_n8143_));
  AOI21_X1   g05427(.A1(new_n8143_), .A2(new_n8140_), .B(pi0042), .ZN(new_n8144_));
  AOI21_X1   g05428(.A1(new_n8137_), .A2(new_n8144_), .B(new_n8130_), .ZN(new_n8145_));
  NAND2_X1   g05429(.A1(new_n8125_), .A2(new_n2523_), .ZN(new_n8146_));
  NOR4_X1    g05430(.A1(new_n8145_), .A2(new_n8108_), .A3(new_n8128_), .A4(new_n8146_), .ZN(new_n8147_));
  AOI22_X1   g05431(.A1(new_n8001_), .A2(pi0099), .B1(pi0072), .B2(new_n5172_), .ZN(new_n8148_));
  OAI21_X1   g05432(.A1(new_n8148_), .A2(pi0113), .B(new_n8113_), .ZN(new_n8149_));
  AOI21_X1   g05433(.A1(new_n8149_), .A2(new_n8109_), .B(new_n8110_), .ZN(new_n8150_));
  NAND2_X1   g05434(.A1(new_n8150_), .A2(new_n8138_), .ZN(new_n8151_));
  NOR2_X1    g05435(.A1(new_n8006_), .A2(new_n5172_), .ZN(new_n8152_));
  NAND2_X1   g05436(.A1(new_n8152_), .A2(new_n8141_), .ZN(new_n8153_));
  INV_X1     g05437(.I(new_n8153_), .ZN(new_n8154_));
  AOI21_X1   g05438(.A1(new_n8154_), .A2(new_n8140_), .B(pi0042), .ZN(new_n8155_));
  NAND2_X1   g05439(.A1(new_n8151_), .A2(new_n8155_), .ZN(new_n8156_));
  MUX2_X1    g05440(.I0(new_n8156_), .I1(new_n8108_), .S(pi0115), .Z(new_n8157_));
  OAI21_X1   g05441(.A1(new_n8157_), .A2(pi0228), .B(new_n3154_), .ZN(new_n8158_));
  MUX2_X1    g05442(.I0(new_n8019_), .I1(new_n2861_), .S(new_n8012_), .Z(new_n8159_));
  NOR2_X1    g05443(.A1(pi0199), .A2(pi0200), .ZN(new_n8160_));
  INV_X1     g05444(.I(new_n8160_), .ZN(new_n8161_));
  NAND3_X1   g05445(.A1(new_n8159_), .A2(new_n5987_), .A3(new_n8161_), .ZN(new_n8162_));
  INV_X1     g05446(.I(new_n7928_), .ZN(new_n8163_));
  INV_X1     g05447(.I(new_n8019_), .ZN(new_n8164_));
  NOR2_X1    g05448(.A1(new_n8164_), .A2(new_n8163_), .ZN(new_n8165_));
  NOR2_X1    g05449(.A1(new_n5987_), .A2(new_n2587_), .ZN(new_n8166_));
  INV_X1     g05450(.I(new_n8166_), .ZN(new_n8167_));
  NOR3_X1    g05451(.A1(new_n8165_), .A2(new_n8083_), .A3(new_n8167_), .ZN(new_n8168_));
  NOR2_X1    g05452(.A1(pi0199), .A2(pi0299), .ZN(new_n8169_));
  INV_X1     g05453(.I(new_n8169_), .ZN(new_n8170_));
  NOR4_X1    g05454(.A1(new_n8170_), .A2(pi0072), .A3(new_n8098_), .A4(pi0232), .ZN(new_n8171_));
  NOR4_X1    g05455(.A1(new_n8162_), .A2(new_n8168_), .A3(new_n6594_), .A4(new_n8171_), .ZN(new_n8172_));
  NOR3_X1    g05456(.A1(new_n8147_), .A2(new_n8158_), .A3(new_n8172_), .ZN(new_n8173_));
  AOI21_X1   g05457(.A1(new_n6481_), .A2(new_n8108_), .B(new_n8129_), .ZN(new_n8174_));
  INV_X1     g05458(.I(new_n8032_), .ZN(new_n8175_));
  NOR2_X1    g05459(.A1(new_n8175_), .A2(new_n5174_), .ZN(new_n8176_));
  INV_X1     g05460(.I(new_n8176_), .ZN(new_n8177_));
  NOR2_X1    g05461(.A1(new_n8177_), .A2(new_n8142_), .ZN(new_n8178_));
  AOI21_X1   g05462(.A1(new_n8178_), .A2(new_n6010_), .B(pi0072), .ZN(new_n8179_));
  INV_X1     g05463(.I(new_n8179_), .ZN(new_n8180_));
  NAND2_X1   g05464(.A1(new_n8035_), .A2(new_n8120_), .ZN(new_n8181_));
  NOR2_X1    g05465(.A1(new_n8181_), .A2(new_n6436_), .ZN(new_n8182_));
  INV_X1     g05466(.I(new_n8182_), .ZN(new_n8183_));
  NOR3_X1    g05467(.A1(new_n8183_), .A2(pi0114), .A3(new_n5167_), .ZN(new_n8184_));
  NAND3_X1   g05468(.A1(new_n8180_), .A2(new_n8074_), .A3(new_n8184_), .ZN(new_n8185_));
  OAI21_X1   g05469(.A1(pi0042), .A2(new_n8184_), .B(new_n8179_), .ZN(new_n8186_));
  NAND4_X1   g05470(.A1(new_n8185_), .A2(new_n8138_), .A3(new_n8140_), .A4(new_n8186_), .ZN(new_n8187_));
  AOI22_X1   g05471(.A1(new_n8187_), .A2(new_n8174_), .B1(new_n8025_), .B2(new_n8108_), .ZN(new_n8188_));
  NOR2_X1    g05472(.A1(new_n8188_), .A2(pi0039), .ZN(new_n8189_));
  NOR2_X1    g05473(.A1(new_n8084_), .A2(new_n2587_), .ZN(new_n8190_));
  NOR2_X1    g05474(.A1(new_n8190_), .A2(new_n3154_), .ZN(new_n8191_));
  INV_X1     g05475(.I(new_n8191_), .ZN(new_n8192_));
  NOR3_X1    g05476(.A1(new_n8192_), .A2(new_n8097_), .A3(new_n8102_), .ZN(new_n8193_));
  INV_X1     g05477(.I(new_n8193_), .ZN(new_n8194_));
  AOI21_X1   g05478(.A1(new_n8189_), .A2(new_n8194_), .B(new_n5159_), .ZN(new_n8195_));
  OAI21_X1   g05479(.A1(new_n8102_), .A2(new_n8097_), .B(new_n8105_), .ZN(new_n8196_));
  NOR2_X1    g05480(.A1(new_n8192_), .A2(new_n8097_), .ZN(new_n8197_));
  NOR2_X1    g05481(.A1(new_n8197_), .A2(new_n8104_), .ZN(new_n8198_));
  NOR4_X1    g05482(.A1(new_n8198_), .A2(new_n3172_), .A3(pi0087), .A4(new_n8196_), .ZN(new_n8199_));
  OAI21_X1   g05483(.A1(new_n8195_), .A2(new_n8199_), .B(new_n2621_), .ZN(new_n8200_));
  NAND2_X1   g05484(.A1(new_n8176_), .A2(pi0228), .ZN(new_n8201_));
  OAI21_X1   g05485(.A1(new_n8201_), .A2(new_n5164_), .B(new_n8075_), .ZN(new_n8202_));
  NOR2_X1    g05486(.A1(new_n8181_), .A2(new_n2523_), .ZN(new_n8203_));
  NAND3_X1   g05487(.A1(new_n8203_), .A2(new_n8138_), .A3(new_n8125_), .ZN(new_n8204_));
  NOR3_X1    g05488(.A1(new_n8204_), .A2(pi0042), .A3(new_n3197_), .ZN(new_n8205_));
  NAND2_X1   g05489(.A1(new_n8202_), .A2(new_n8205_), .ZN(new_n8206_));
  AOI21_X1   g05490(.A1(new_n8104_), .A2(new_n2622_), .B(new_n3177_), .ZN(new_n8207_));
  INV_X1     g05491(.I(new_n8207_), .ZN(new_n8208_));
  NOR2_X1    g05492(.A1(new_n8193_), .A2(new_n8208_), .ZN(new_n8209_));
  AOI21_X1   g05493(.A1(new_n8206_), .A2(new_n8209_), .B(pi0075), .ZN(new_n8210_));
  OAI21_X1   g05494(.A1(new_n8173_), .A2(new_n8200_), .B(new_n8210_), .ZN(new_n8211_));
  NOR2_X1    g05495(.A1(new_n5941_), .A2(new_n2628_), .ZN(new_n8212_));
  INV_X1     g05496(.I(new_n8212_), .ZN(new_n8213_));
  NAND2_X1   g05497(.A1(new_n8184_), .A2(new_n5994_), .ZN(new_n8214_));
  NOR2_X1    g05498(.A1(new_n8214_), .A2(pi0042), .ZN(new_n8215_));
  INV_X1     g05499(.I(new_n8063_), .ZN(new_n8216_));
  NOR2_X1    g05500(.A1(new_n8216_), .A2(new_n5174_), .ZN(new_n8217_));
  INV_X1     g05501(.I(new_n8217_), .ZN(new_n8218_));
  NOR2_X1    g05502(.A1(new_n8218_), .A2(new_n8142_), .ZN(new_n8219_));
  OAI21_X1   g05503(.A1(new_n8219_), .A2(new_n8108_), .B(new_n8138_), .ZN(new_n8220_));
  OAI21_X1   g05504(.A1(new_n8220_), .A2(new_n8215_), .B(new_n8140_), .ZN(new_n8221_));
  NAND2_X1   g05505(.A1(new_n8221_), .A2(new_n8174_), .ZN(new_n8222_));
  AOI21_X1   g05506(.A1(new_n8025_), .A2(new_n8108_), .B(new_n3208_), .ZN(new_n8223_));
  OAI21_X1   g05507(.A1(new_n3208_), .A2(new_n8075_), .B(new_n3154_), .ZN(new_n8224_));
  AOI21_X1   g05508(.A1(new_n8222_), .A2(new_n8223_), .B(new_n8224_), .ZN(new_n8225_));
  AOI21_X1   g05509(.A1(new_n8225_), .A2(new_n8194_), .B(new_n8213_), .ZN(new_n8226_));
  AOI21_X1   g05510(.A1(new_n8211_), .A2(new_n8226_), .B(new_n8107_), .ZN(new_n8227_));
  AOI21_X1   g05511(.A1(new_n8198_), .A2(new_n5942_), .B(new_n8082_), .ZN(new_n8228_));
  OAI21_X1   g05512(.A1(new_n8227_), .A2(new_n8090_), .B(new_n8228_), .ZN(new_n8229_));
  NOR2_X1    g05513(.A1(new_n8147_), .A2(new_n8158_), .ZN(new_n8230_));
  INV_X1     g05514(.I(new_n8159_), .ZN(new_n8231_));
  OAI21_X1   g05515(.A1(new_n8231_), .A2(new_n8096_), .B(pi0039), .ZN(new_n8232_));
  AOI21_X1   g05516(.A1(new_n8230_), .A2(new_n8232_), .B(new_n2622_), .ZN(new_n8233_));
  NOR2_X1    g05517(.A1(new_n8097_), .A2(new_n3154_), .ZN(new_n8234_));
  NOR3_X1    g05518(.A1(new_n8188_), .A2(pi0039), .A3(new_n8234_), .ZN(new_n8235_));
  INV_X1     g05519(.I(new_n8234_), .ZN(new_n8236_));
  AOI21_X1   g05520(.A1(new_n8225_), .A2(new_n8236_), .B(new_n8213_), .ZN(new_n8237_));
  NAND3_X1   g05521(.A1(new_n8206_), .A2(new_n8207_), .A3(new_n8236_), .ZN(new_n8238_));
  NAND2_X1   g05522(.A1(new_n8238_), .A2(new_n2628_), .ZN(new_n8239_));
  NOR3_X1    g05523(.A1(new_n3173_), .A2(pi0038), .A3(pi0087), .ZN(new_n8240_));
  NAND2_X1   g05524(.A1(new_n8239_), .A2(new_n8240_), .ZN(new_n8241_));
  NOR4_X1    g05525(.A1(new_n8233_), .A2(new_n8235_), .A3(new_n8237_), .A4(new_n8241_), .ZN(new_n8242_));
  OAI21_X1   g05526(.A1(new_n8234_), .A2(new_n8106_), .B(new_n8090_), .ZN(new_n8243_));
  OAI21_X1   g05527(.A1(new_n8242_), .A2(new_n8243_), .B(new_n8107_), .ZN(new_n8244_));
  AOI21_X1   g05528(.A1(new_n8244_), .A2(new_n8082_), .B(po1038), .ZN(new_n8245_));
  AOI22_X1   g05529(.A1(new_n8245_), .A2(new_n8229_), .B1(po1038), .B2(new_n8086_), .ZN(po0200));
  INV_X1     g05530(.I(pi0219), .ZN(new_n8247_));
  NOR2_X1    g05531(.A1(new_n8076_), .A2(new_n8078_), .ZN(new_n8248_));
  NOR2_X1    g05532(.A1(new_n8248_), .A2(new_n8077_), .ZN(new_n8249_));
  INV_X1     g05533(.I(new_n8248_), .ZN(new_n8250_));
  NOR2_X1    g05534(.A1(new_n8250_), .A2(pi0211), .ZN(new_n8251_));
  AOI21_X1   g05535(.A1(new_n8251_), .A2(new_n8247_), .B(new_n8249_), .ZN(new_n8252_));
  INV_X1     g05536(.I(new_n8252_), .ZN(new_n8253_));
  NOR2_X1    g05537(.A1(new_n8119_), .A2(new_n2921_), .ZN(new_n8254_));
  NOR2_X1    g05538(.A1(new_n8134_), .A2(new_n2922_), .ZN(new_n8255_));
  OAI21_X1   g05539(.A1(new_n8255_), .A2(new_n8254_), .B(pi0228), .ZN(new_n8256_));
  OAI21_X1   g05540(.A1(pi0228), .A2(new_n8150_), .B(new_n8256_), .ZN(new_n8257_));
  NOR3_X1    g05541(.A1(pi0042), .A2(pi0114), .A3(pi0115), .ZN(new_n8258_));
  INV_X1     g05542(.I(pi0043), .ZN(new_n8259_));
  NOR2_X1    g05543(.A1(new_n8259_), .A2(pi0072), .ZN(new_n8260_));
  NOR2_X1    g05544(.A1(new_n8260_), .A2(new_n8258_), .ZN(new_n8261_));
  NOR2_X1    g05545(.A1(new_n7964_), .A2(new_n5172_), .ZN(new_n8262_));
  NOR2_X1    g05546(.A1(new_n8262_), .A2(new_n2922_), .ZN(new_n8263_));
  AOI21_X1   g05547(.A1(new_n7975_), .A2(new_n5171_), .B(new_n2921_), .ZN(new_n8264_));
  NOR4_X1    g05548(.A1(new_n8263_), .A2(new_n2523_), .A3(new_n8142_), .A4(new_n8264_), .ZN(new_n8265_));
  AOI21_X1   g05549(.A1(new_n2523_), .A2(new_n8154_), .B(new_n8265_), .ZN(new_n8266_));
  NAND3_X1   g05550(.A1(new_n8261_), .A2(pi0043), .A3(new_n8258_), .ZN(new_n8267_));
  NOR2_X1    g05551(.A1(new_n8160_), .A2(pi0299), .ZN(new_n8268_));
  INV_X1     g05552(.I(new_n8268_), .ZN(new_n8269_));
  AOI21_X1   g05553(.A1(new_n8269_), .A2(new_n2861_), .B(pi0232), .ZN(new_n8270_));
  NOR2_X1    g05554(.A1(new_n8270_), .A2(pi0299), .ZN(new_n8271_));
  INV_X1     g05555(.I(new_n8271_), .ZN(new_n8272_));
  NAND2_X1   g05556(.A1(new_n8159_), .A2(new_n8160_), .ZN(new_n8273_));
  AOI21_X1   g05557(.A1(new_n8273_), .A2(pi0232), .B(new_n8272_), .ZN(new_n8274_));
  OAI21_X1   g05558(.A1(new_n8257_), .A2(new_n8267_), .B(new_n3154_), .ZN(new_n8275_));
  AOI21_X1   g05559(.A1(new_n8091_), .A2(new_n8160_), .B(new_n7178_), .ZN(new_n8276_));
  NAND2_X1   g05560(.A1(new_n8272_), .A2(new_n8276_), .ZN(new_n8277_));
  INV_X1     g05561(.I(new_n8277_), .ZN(new_n8278_));
  INV_X1     g05562(.I(new_n8260_), .ZN(new_n8279_));
  AOI21_X1   g05563(.A1(new_n2921_), .A2(new_n8258_), .B(new_n8025_), .ZN(new_n8280_));
  INV_X1     g05564(.I(new_n8280_), .ZN(new_n8284_));
  NOR2_X1    g05565(.A1(new_n8260_), .A2(pi0039), .ZN(new_n8287_));
  NOR2_X1    g05566(.A1(new_n8278_), .A2(new_n8287_), .ZN(new_n8288_));
  INV_X1     g05567(.I(new_n8288_), .ZN(new_n8289_));
  NOR2_X1    g05568(.A1(pi0038), .A2(pi0100), .ZN(new_n8291_));
  NAND2_X1   g05569(.A1(new_n8275_), .A2(new_n8291_), .ZN(new_n8292_));
  NAND4_X1   g05570(.A1(new_n8182_), .A2(new_n8259_), .A3(pi0052), .A4(new_n5994_), .ZN(new_n8293_));
  NOR2_X1    g05571(.A1(new_n8219_), .A2(pi0072), .ZN(new_n8294_));
  NAND2_X1   g05572(.A1(new_n8294_), .A2(pi0043), .ZN(new_n8295_));
  XOR2_X1    g05573(.A1(new_n8295_), .A2(new_n8293_), .Z(new_n8296_));
  MUX2_X1    g05574(.I0(new_n8296_), .I1(new_n8260_), .S(new_n8284_), .Z(new_n8297_));
  OAI21_X1   g05575(.A1(new_n3207_), .A2(new_n8260_), .B(new_n8297_), .ZN(new_n8298_));
  OR3_X2     g05576(.A1(new_n8297_), .A2(new_n3207_), .A3(new_n8279_), .Z(new_n8299_));
  NAND4_X1   g05577(.A1(new_n8299_), .A2(new_n3154_), .A3(new_n8277_), .A4(new_n8298_), .ZN(new_n8300_));
  NOR2_X1    g05578(.A1(new_n8289_), .A2(new_n5941_), .ZN(new_n8301_));
  INV_X1     g05579(.I(new_n8287_), .ZN(new_n8302_));
  NAND2_X1   g05580(.A1(new_n8258_), .A2(pi0228), .ZN(new_n8303_));
  INV_X1     g05581(.I(new_n8181_), .ZN(new_n8304_));
  NOR2_X1    g05582(.A1(new_n8178_), .A2(pi0072), .ZN(new_n8305_));
  MUX2_X1    g05583(.I0(new_n8305_), .I1(new_n8304_), .S(new_n8259_), .Z(new_n8306_));
  NOR4_X1    g05584(.A1(new_n8306_), .A2(new_n3197_), .A3(new_n8260_), .A4(new_n8303_), .ZN(new_n8307_));
  NOR2_X1    g05585(.A1(new_n2621_), .A2(pi0087), .ZN(new_n8308_));
  INV_X1     g05586(.I(new_n8308_), .ZN(new_n8309_));
  NOR2_X1    g05587(.A1(new_n8288_), .A2(new_n2546_), .ZN(new_n8310_));
  NOR4_X1    g05588(.A1(new_n8307_), .A2(new_n8302_), .A3(new_n8309_), .A4(new_n8310_), .ZN(new_n8311_));
  OAI22_X1   g05589(.A1(new_n8311_), .A2(pi0075), .B1(new_n8090_), .B2(new_n8301_), .ZN(new_n8312_));
  AOI21_X1   g05590(.A1(new_n8300_), .A2(new_n8212_), .B(new_n8312_), .ZN(new_n8313_));
  AOI21_X1   g05591(.A1(new_n8292_), .A2(new_n8313_), .B(new_n8253_), .ZN(new_n8314_));
  NAND2_X1   g05592(.A1(new_n8191_), .A2(new_n8101_), .ZN(new_n8315_));
  NOR2_X1    g05593(.A1(new_n5941_), .A2(new_n8287_), .ZN(new_n8316_));
  AOI21_X1   g05594(.A1(new_n8315_), .A2(new_n8316_), .B(new_n8089_), .ZN(new_n8317_));
  OAI21_X1   g05595(.A1(new_n8317_), .A2(new_n8252_), .B(new_n6845_), .ZN(new_n8318_));
  NOR2_X1    g05596(.A1(new_n8252_), .A2(new_n8084_), .ZN(new_n8319_));
  NAND2_X1   g05597(.A1(new_n6845_), .A2(pi0039), .ZN(new_n8320_));
  OAI22_X1   g05598(.A1(new_n8314_), .A2(new_n8318_), .B1(new_n8319_), .B2(new_n8320_), .ZN(po0201));
  INV_X1     g05599(.I(new_n7934_), .ZN(new_n8322_));
  NAND3_X1   g05600(.A1(new_n2576_), .A2(new_n5988_), .A3(new_n2861_), .ZN(new_n8323_));
  MUX2_X1    g05601(.I0(new_n8323_), .I1(new_n8322_), .S(new_n3154_), .Z(new_n8324_));
  AOI21_X1   g05602(.A1(pi0044), .A2(pi0072), .B(new_n2918_), .ZN(new_n8325_));
  NAND2_X1   g05603(.A1(new_n5995_), .A2(new_n8325_), .ZN(new_n8326_));
  NOR4_X1    g05604(.A1(new_n2491_), .A2(pi0044), .A3(new_n5993_), .A4(new_n6436_), .ZN(new_n8327_));
  AOI21_X1   g05605(.A1(new_n8062_), .A2(pi0044), .B(new_n8327_), .ZN(new_n8328_));
  AOI21_X1   g05606(.A1(new_n8025_), .A2(new_n8322_), .B(pi0039), .ZN(new_n8329_));
  AOI21_X1   g05607(.A1(new_n2922_), .A2(new_n7934_), .B(new_n8025_), .ZN(new_n8330_));
  INV_X1     g05608(.I(new_n8330_), .ZN(new_n8331_));
  NOR2_X1    g05609(.A1(new_n8331_), .A2(new_n8329_), .ZN(new_n8332_));
  OAI21_X1   g05610(.A1(new_n8328_), .A2(new_n8326_), .B(new_n8332_), .ZN(new_n8333_));
  INV_X1     g05611(.I(new_n5990_), .ZN(new_n8334_));
  NOR3_X1    g05612(.A1(new_n8334_), .A2(new_n3154_), .A3(pi0072), .ZN(new_n8335_));
  NOR2_X1    g05613(.A1(new_n8335_), .A2(new_n3208_), .ZN(new_n8336_));
  NAND2_X1   g05614(.A1(new_n8333_), .A2(new_n8336_), .ZN(new_n8337_));
  AOI21_X1   g05615(.A1(new_n3154_), .A2(new_n7933_), .B(pi0072), .ZN(new_n8338_));
  OAI21_X1   g05616(.A1(new_n5990_), .A2(new_n3154_), .B(new_n8338_), .ZN(new_n8339_));
  INV_X1     g05617(.I(new_n8339_), .ZN(new_n8340_));
  NOR2_X1    g05618(.A1(new_n3208_), .A2(pi0075), .ZN(new_n8341_));
  INV_X1     g05619(.I(new_n8341_), .ZN(new_n8342_));
  NOR2_X1    g05620(.A1(new_n8340_), .A2(new_n8342_), .ZN(new_n8343_));
  NAND4_X1   g05621(.A1(new_n7951_), .A2(new_n7962_), .A3(pi0044), .A4(new_n2922_), .ZN(new_n8344_));
  NAND2_X1   g05622(.A1(new_n7967_), .A2(pi0044), .ZN(new_n8345_));
  NAND4_X1   g05623(.A1(new_n8344_), .A2(new_n2922_), .A3(new_n7974_), .A4(new_n8345_), .ZN(new_n8346_));
  NAND3_X1   g05624(.A1(new_n7997_), .A2(pi0044), .A3(pi0228), .ZN(new_n8347_));
  NAND2_X1   g05625(.A1(new_n8347_), .A2(new_n3154_), .ZN(new_n8348_));
  AOI21_X1   g05626(.A1(new_n8346_), .A2(pi0228), .B(new_n8348_), .ZN(new_n8349_));
  NAND2_X1   g05627(.A1(new_n8030_), .A2(pi0287), .ZN(new_n8350_));
  NAND2_X1   g05628(.A1(new_n8350_), .A2(new_n2861_), .ZN(new_n8351_));
  INV_X1     g05629(.I(new_n8351_), .ZN(new_n8352_));
  NAND3_X1   g05630(.A1(new_n8352_), .A2(new_n3319_), .A3(new_n5990_), .ZN(new_n8353_));
  NAND2_X1   g05631(.A1(new_n2491_), .A2(new_n7933_), .ZN(new_n8354_));
  XOR2_X1    g05632(.A1(new_n6010_), .A2(new_n7933_), .Z(new_n8355_));
  OAI21_X1   g05633(.A1(new_n8030_), .A2(new_n6436_), .B(new_n8355_), .ZN(new_n8356_));
  OAI21_X1   g05634(.A1(new_n8340_), .A2(new_n3172_), .B(new_n3177_), .ZN(new_n8357_));
  NOR2_X1    g05635(.A1(new_n8335_), .A2(new_n5159_), .ZN(new_n8358_));
  NOR4_X1    g05636(.A1(new_n8326_), .A2(new_n8329_), .A3(new_n8330_), .A4(new_n8358_), .ZN(new_n8359_));
  NAND2_X1   g05637(.A1(new_n8359_), .A2(new_n8357_), .ZN(new_n8360_));
  AOI21_X1   g05638(.A1(new_n8356_), .A2(new_n8354_), .B(new_n8360_), .ZN(new_n8361_));
  OAI21_X1   g05639(.A1(new_n8349_), .A2(new_n8353_), .B(new_n8361_), .ZN(new_n8362_));
  NOR4_X1    g05640(.A1(new_n8031_), .A2(new_n2523_), .A3(new_n2622_), .A4(new_n7934_), .ZN(new_n8363_));
  NOR4_X1    g05641(.A1(new_n2491_), .A2(pi0044), .A3(new_n2523_), .A4(new_n2622_), .ZN(new_n8364_));
  OR3_X2     g05642(.A1(new_n8363_), .A2(pi0039), .A3(new_n8364_), .Z(new_n8365_));
  NOR3_X1    g05643(.A1(new_n8334_), .A2(pi0072), .A3(new_n2624_), .ZN(new_n8366_));
  AOI21_X1   g05644(.A1(new_n8365_), .A2(new_n8366_), .B(pi0075), .ZN(new_n8367_));
  AOI22_X1   g05645(.A1(new_n8362_), .A2(new_n8367_), .B1(new_n8337_), .B2(new_n8343_), .ZN(new_n8368_));
  NAND2_X1   g05646(.A1(po1038), .A2(new_n5941_), .ZN(new_n8369_));
  OAI22_X1   g05647(.A1(new_n8368_), .A2(new_n8369_), .B1(new_n6845_), .B2(new_n8324_), .ZN(po0202));
  NAND2_X1   g05648(.A1(new_n7832_), .A2(new_n5525_), .ZN(new_n8371_));
  NOR3_X1    g05649(.A1(new_n5359_), .A2(new_n5119_), .A3(new_n8371_), .ZN(po0203));
  NOR2_X1    g05650(.A1(new_n5305_), .A2(new_n2640_), .ZN(new_n8373_));
  NOR3_X1    g05651(.A1(new_n7000_), .A2(new_n2492_), .A3(pi0071), .ZN(new_n8374_));
  AND4_X2    g05652(.A1(new_n5955_), .A2(new_n7009_), .A3(new_n7006_), .A4(new_n8374_), .Z(new_n8375_));
  NOR4_X1    g05653(.A1(pi0049), .A2(pi0068), .A3(pi0073), .A4(pi0076), .ZN(new_n8376_));
  NOR3_X1    g05654(.A1(pi0102), .A2(pi0104), .A3(pi0111), .ZN(new_n8377_));
  INV_X1     g05655(.I(new_n8377_), .ZN(new_n8378_));
  NAND2_X1   g05656(.A1(new_n7889_), .A2(new_n2784_), .ZN(new_n8379_));
  NOR4_X1    g05657(.A1(new_n8378_), .A2(pi0089), .A3(new_n8379_), .A4(new_n8376_), .ZN(new_n8380_));
  NAND4_X1   g05658(.A1(new_n8375_), .A2(new_n6998_), .A3(new_n8380_), .A4(new_n7893_), .ZN(new_n8381_));
  OAI21_X1   g05659(.A1(pi0841), .A2(new_n8381_), .B(new_n7828_), .ZN(new_n8382_));
  AOI21_X1   g05660(.A1(new_n8373_), .A2(pi0024), .B(new_n8382_), .ZN(po0204));
  NOR2_X1    g05661(.A1(new_n2745_), .A2(pi0089), .ZN(new_n8384_));
  INV_X1     g05662(.I(new_n2764_), .ZN(new_n8385_));
  NOR4_X1    g05663(.A1(new_n7837_), .A2(new_n2747_), .A3(new_n8385_), .A4(new_n7215_), .ZN(new_n8386_));
  NAND2_X1   g05664(.A1(new_n8384_), .A2(new_n8386_), .ZN(new_n8387_));
  NAND2_X1   g05665(.A1(new_n7005_), .A2(new_n7073_), .ZN(new_n8388_));
  NOR3_X1    g05666(.A1(new_n7000_), .A2(pi0067), .A3(pi0103), .ZN(new_n8389_));
  INV_X1     g05667(.I(new_n8389_), .ZN(new_n8390_));
  NOR4_X1    g05668(.A1(new_n8388_), .A2(new_n8390_), .A3(pi0036), .A4(pi0098), .ZN(new_n8391_));
  NAND2_X1   g05669(.A1(new_n8387_), .A2(new_n8391_), .ZN(new_n8392_));
  OAI21_X1   g05670(.A1(new_n2778_), .A2(new_n8392_), .B(new_n2710_), .ZN(new_n8393_));
  INV_X1     g05671(.I(pi0098), .ZN(new_n8394_));
  NAND4_X1   g05672(.A1(new_n2702_), .A2(new_n2710_), .A3(new_n8394_), .A4(new_n5956_), .ZN(new_n8395_));
  NOR2_X1    g05673(.A1(new_n8395_), .A2(new_n2663_), .ZN(new_n8396_));
  NAND2_X1   g05674(.A1(new_n8393_), .A2(new_n8396_), .ZN(new_n8397_));
  INV_X1     g05675(.I(new_n8397_), .ZN(new_n8398_));
  NAND2_X1   g05676(.A1(new_n8398_), .A2(new_n2660_), .ZN(new_n8399_));
  NAND2_X1   g05677(.A1(new_n8399_), .A2(new_n6020_), .ZN(new_n8400_));
  AOI21_X1   g05678(.A1(new_n8400_), .A2(new_n7368_), .B(new_n7827_), .ZN(new_n8401_));
  INV_X1     g05679(.I(new_n8401_), .ZN(new_n8402_));
  NAND2_X1   g05680(.A1(new_n8402_), .A2(pi1093), .ZN(new_n8403_));
  INV_X1     g05681(.I(new_n2955_), .ZN(new_n8404_));
  INV_X1     g05682(.I(new_n5114_), .ZN(new_n8405_));
  NAND3_X1   g05683(.A1(new_n8387_), .A2(new_n8391_), .A3(new_n2767_), .ZN(new_n8406_));
  AOI21_X1   g05684(.A1(new_n8406_), .A2(new_n2710_), .B(new_n8395_), .ZN(new_n8407_));
  NAND2_X1   g05685(.A1(new_n7848_), .A2(new_n8407_), .ZN(new_n8408_));
  NOR3_X1    g05686(.A1(new_n8408_), .A2(new_n2955_), .A3(new_n8405_), .ZN(new_n8409_));
  OAI21_X1   g05687(.A1(new_n8402_), .A2(new_n8404_), .B(new_n8409_), .ZN(new_n8410_));
  MUX2_X1    g05688(.I0(new_n8403_), .I1(new_n8410_), .S(new_n2958_), .Z(new_n8411_));
  NOR2_X1    g05689(.A1(new_n8402_), .A2(new_n6004_), .ZN(new_n8412_));
  NOR2_X1    g05690(.A1(new_n5363_), .A2(new_n6003_), .ZN(new_n8413_));
  NOR3_X1    g05691(.A1(new_n7821_), .A2(new_n6005_), .A3(new_n7827_), .ZN(new_n8414_));
  NOR2_X1    g05692(.A1(new_n8414_), .A2(new_n8413_), .ZN(new_n8415_));
  OAI21_X1   g05693(.A1(new_n8412_), .A2(new_n8415_), .B(new_n7824_), .ZN(new_n8416_));
  OAI21_X1   g05694(.A1(pi0829), .A2(new_n8412_), .B(new_n8410_), .ZN(new_n8417_));
  NAND4_X1   g05695(.A1(new_n8417_), .A2(new_n2918_), .A3(new_n2924_), .A4(new_n8416_), .ZN(new_n8418_));
  NOR2_X1    g05696(.A1(new_n8418_), .A2(new_n8411_), .ZN(po0205));
  NOR3_X1    g05697(.A1(new_n2644_), .A2(pi0072), .A3(new_n2902_), .ZN(new_n8420_));
  NAND2_X1   g05698(.A1(new_n8420_), .A2(new_n2658_), .ZN(new_n8421_));
  NOR4_X1    g05699(.A1(new_n7825_), .A2(new_n7847_), .A3(new_n7896_), .A4(new_n8421_), .ZN(po0206));
  INV_X1     g05700(.I(new_n5918_), .ZN(new_n8423_));
  NOR4_X1    g05701(.A1(new_n8378_), .A2(pi0045), .A3(new_n7835_), .A4(pi0082), .ZN(new_n8424_));
  OR3_X2     g05702(.A1(new_n2769_), .A2(pi0103), .A3(new_n7892_), .Z(new_n8425_));
  NAND3_X1   g05703(.A1(new_n7005_), .A2(new_n2757_), .A3(new_n2728_), .ZN(new_n8426_));
  NOR2_X1    g05704(.A1(new_n8426_), .A2(new_n8425_), .ZN(new_n8427_));
  NOR2_X1    g05705(.A1(new_n7070_), .A2(new_n7000_), .ZN(new_n8428_));
  NAND4_X1   g05706(.A1(new_n8427_), .A2(new_n8384_), .A3(new_n8428_), .A4(new_n8424_), .ZN(new_n8429_));
  NOR3_X1    g05707(.A1(new_n8429_), .A2(new_n2646_), .A3(new_n6999_), .ZN(new_n8430_));
  NAND3_X1   g05708(.A1(new_n8430_), .A2(new_n7826_), .A3(new_n8420_), .ZN(new_n8431_));
  MUX2_X1    g05709(.I0(new_n8431_), .I1(new_n7793_), .S(pi0074), .Z(new_n8432_));
  NOR3_X1    g05710(.A1(new_n8432_), .A2(new_n8423_), .A3(po1038), .ZN(po0207));
  NAND4_X1   g05711(.A1(new_n6971_), .A2(new_n6976_), .A3(new_n6979_), .A4(new_n7797_), .ZN(new_n8434_));
  NAND2_X1   g05712(.A1(new_n2534_), .A2(new_n2544_), .ZN(new_n8435_));
  AOI21_X1   g05713(.A1(new_n8434_), .A2(new_n8435_), .B(new_n6967_), .ZN(po0208));
  INV_X1     g05714(.I(new_n2663_), .ZN(new_n8437_));
  NAND3_X1   g05715(.A1(new_n7828_), .A2(new_n2638_), .A3(new_n8437_), .ZN(new_n8438_));
  NAND2_X1   g05716(.A1(new_n8428_), .A2(new_n7075_), .ZN(new_n8439_));
  INV_X1     g05717(.I(new_n8439_), .ZN(new_n8440_));
  NOR2_X1    g05718(.A1(new_n7888_), .A2(pi0069), .ZN(new_n8441_));
  NAND2_X1   g05719(.A1(new_n8440_), .A2(new_n8441_), .ZN(new_n8442_));
  NOR2_X1    g05720(.A1(new_n8442_), .A2(new_n2769_), .ZN(new_n8443_));
  INV_X1     g05721(.I(new_n8443_), .ZN(new_n8444_));
  NOR3_X1    g05722(.A1(new_n8438_), .A2(new_n2765_), .A3(new_n8444_), .ZN(po0209));
  NOR2_X1    g05723(.A1(new_n8248_), .A2(pi0211), .ZN(new_n8446_));
  INV_X1     g05724(.I(new_n8446_), .ZN(new_n8447_));
  NOR2_X1    g05725(.A1(new_n8447_), .A2(pi0219), .ZN(new_n8448_));
  INV_X1     g05726(.I(pi0052), .ZN(new_n8449_));
  NOR2_X1    g05727(.A1(new_n8449_), .A2(pi0072), .ZN(new_n8450_));
  NAND4_X1   g05728(.A1(new_n6845_), .A2(new_n8448_), .A3(pi0039), .A4(new_n8083_), .ZN(new_n8451_));
  INV_X1     g05729(.I(new_n8448_), .ZN(new_n8452_));
  OAI21_X1   g05730(.A1(new_n8143_), .A2(pi0052), .B(new_n8130_), .ZN(new_n8453_));
  AOI21_X1   g05731(.A1(new_n8134_), .A2(pi0052), .B(new_n8453_), .ZN(new_n8454_));
  INV_X1     g05732(.I(new_n8121_), .ZN(new_n8455_));
  NAND4_X1   g05733(.A1(new_n8123_), .A2(pi0052), .A3(new_n8125_), .A4(new_n2922_), .ZN(new_n8456_));
  NOR3_X1    g05734(.A1(new_n5166_), .A2(pi0114), .A3(pi0115), .ZN(new_n8457_));
  OAI21_X1   g05735(.A1(new_n8154_), .A2(pi0052), .B(new_n8457_), .ZN(new_n8458_));
  AOI21_X1   g05736(.A1(new_n8150_), .A2(pi0052), .B(new_n8458_), .ZN(new_n8459_));
  INV_X1     g05737(.I(new_n8450_), .ZN(new_n8460_));
  NAND2_X1   g05738(.A1(new_n8457_), .A2(new_n8460_), .ZN(new_n8461_));
  NAND2_X1   g05739(.A1(new_n8461_), .A2(new_n2523_), .ZN(new_n8462_));
  OAI21_X1   g05740(.A1(new_n8459_), .A2(new_n8462_), .B(new_n3154_), .ZN(new_n8463_));
  NOR2_X1    g05741(.A1(new_n5166_), .A2(pi0114), .ZN(new_n8464_));
  NAND2_X1   g05742(.A1(new_n8461_), .A2(pi0228), .ZN(new_n8465_));
  NAND4_X1   g05743(.A1(new_n8456_), .A2(new_n8463_), .A3(new_n8464_), .A4(new_n8465_), .ZN(new_n8466_));
  NOR2_X1    g05744(.A1(new_n8466_), .A2(new_n8454_), .ZN(new_n8467_));
  INV_X1     g05745(.I(new_n8467_), .ZN(new_n8468_));
  NAND3_X1   g05746(.A1(new_n5987_), .A2(new_n2587_), .A3(pi0072), .ZN(new_n8469_));
  NAND2_X1   g05747(.A1(new_n8469_), .A2(pi0039), .ZN(new_n8470_));
  AOI21_X1   g05748(.A1(new_n8468_), .A2(new_n8470_), .B(new_n2622_), .ZN(new_n8471_));
  INV_X1     g05749(.I(new_n8464_), .ZN(new_n8472_));
  NOR2_X1    g05750(.A1(new_n8025_), .A2(new_n8130_), .ZN(new_n8473_));
  INV_X1     g05751(.I(new_n8473_), .ZN(new_n8474_));
  NOR2_X1    g05752(.A1(new_n8474_), .A2(new_n8472_), .ZN(new_n8475_));
  NAND4_X1   g05753(.A1(new_n8178_), .A2(new_n6010_), .A3(new_n8460_), .A4(new_n8475_), .ZN(new_n8476_));
  INV_X1     g05754(.I(new_n8476_), .ZN(new_n8477_));
  NOR2_X1    g05755(.A1(new_n8477_), .A2(pi0039), .ZN(new_n8478_));
  OAI21_X1   g05756(.A1(new_n8478_), .A2(new_n8191_), .B(new_n5158_), .ZN(new_n8479_));
  NOR2_X1    g05757(.A1(new_n8450_), .A2(pi0039), .ZN(new_n8480_));
  NOR2_X1    g05758(.A1(new_n8191_), .A2(new_n8480_), .ZN(new_n8481_));
  AOI21_X1   g05759(.A1(new_n8481_), .A2(new_n3172_), .B(pi0087), .ZN(new_n8482_));
  NAND2_X1   g05760(.A1(new_n8479_), .A2(new_n8482_), .ZN(new_n8483_));
  AOI21_X1   g05761(.A1(new_n8481_), .A2(new_n2622_), .B(new_n3177_), .ZN(new_n8484_));
  NOR2_X1    g05762(.A1(new_n8305_), .A2(new_n8449_), .ZN(new_n8485_));
  AOI21_X1   g05763(.A1(new_n8449_), .A2(new_n8181_), .B(new_n8485_), .ZN(new_n8486_));
  NOR2_X1    g05764(.A1(new_n8457_), .A2(pi0228), .ZN(new_n8487_));
  MUX2_X1    g05765(.I0(new_n8460_), .I1(new_n8486_), .S(new_n8487_), .Z(new_n8488_));
  NOR2_X1    g05766(.A1(new_n8488_), .A2(pi0039), .ZN(new_n8489_));
  OR3_X2     g05767(.A1(new_n8489_), .A2(new_n2622_), .A3(new_n8191_), .Z(new_n8490_));
  AOI21_X1   g05768(.A1(new_n8490_), .A2(new_n8484_), .B(new_n8090_), .ZN(new_n8491_));
  OAI21_X1   g05769(.A1(new_n8471_), .A2(new_n8483_), .B(new_n8491_), .ZN(new_n8492_));
  NAND3_X1   g05770(.A1(new_n8231_), .A2(new_n7348_), .A3(new_n8161_), .ZN(new_n8493_));
  NOR2_X1    g05771(.A1(new_n8168_), .A2(new_n8270_), .ZN(new_n8494_));
  AOI21_X1   g05772(.A1(new_n8494_), .A2(new_n8493_), .B(new_n3154_), .ZN(new_n8495_));
  NOR2_X1    g05773(.A1(new_n8277_), .A2(new_n8190_), .ZN(new_n8496_));
  NOR2_X1    g05774(.A1(new_n8278_), .A2(new_n8480_), .ZN(new_n8498_));
  NOR2_X1    g05775(.A1(pi0038), .A2(pi0100), .ZN(new_n8499_));
  OAI21_X1   g05776(.A1(new_n8467_), .A2(new_n8495_), .B(new_n8499_), .ZN(new_n8500_));
  INV_X1     g05777(.I(new_n8498_), .ZN(new_n8501_));
  AOI21_X1   g05778(.A1(new_n8501_), .A2(new_n8484_), .B(new_n2621_), .ZN(new_n8502_));
  OAI21_X1   g05779(.A1(new_n8489_), .A2(new_n8496_), .B(new_n8502_), .ZN(new_n8503_));
  AOI21_X1   g05780(.A1(new_n8503_), .A2(new_n8090_), .B(pi0087), .ZN(new_n8504_));
  AOI21_X1   g05781(.A1(new_n8500_), .A2(new_n8504_), .B(pi0075), .ZN(new_n8505_));
  NOR2_X1    g05782(.A1(new_n8460_), .A2(pi0039), .ZN(new_n8506_));
  NAND2_X1   g05783(.A1(new_n8219_), .A2(new_n8475_), .ZN(new_n8507_));
  OAI21_X1   g05784(.A1(new_n8507_), .A2(new_n3208_), .B(new_n8506_), .ZN(new_n8508_));
  NAND2_X1   g05785(.A1(new_n8508_), .A2(new_n3154_), .ZN(new_n8509_));
  OAI21_X1   g05786(.A1(new_n8481_), .A2(new_n5941_), .B(new_n8448_), .ZN(new_n8510_));
  NAND4_X1   g05787(.A1(new_n8192_), .A2(new_n2628_), .A3(new_n5942_), .A4(new_n8089_), .ZN(new_n8511_));
  NOR2_X1    g05788(.A1(new_n8511_), .A2(new_n8496_), .ZN(new_n8512_));
  NAND3_X1   g05789(.A1(new_n8509_), .A2(new_n8510_), .A3(new_n8512_), .ZN(new_n8513_));
  AOI21_X1   g05790(.A1(new_n8492_), .A2(new_n8505_), .B(new_n8513_), .ZN(new_n8514_));
  NOR2_X1    g05791(.A1(new_n8274_), .A2(new_n3154_), .ZN(new_n8515_));
  NOR2_X1    g05792(.A1(new_n8467_), .A2(new_n8515_), .ZN(new_n8516_));
  NAND2_X1   g05793(.A1(new_n3172_), .A2(new_n3173_), .ZN(new_n8518_));
  NOR2_X1    g05794(.A1(new_n8489_), .A2(new_n8278_), .ZN(new_n8519_));
  MUX2_X1    g05795(.I0(new_n8519_), .I1(new_n8498_), .S(new_n2622_), .Z(new_n8520_));
  NAND2_X1   g05796(.A1(new_n8507_), .A2(new_n8450_), .ZN(new_n8521_));
  AOI21_X1   g05797(.A1(new_n8521_), .A2(new_n3154_), .B(new_n8278_), .ZN(new_n8522_));
  OAI21_X1   g05798(.A1(new_n8498_), .A2(new_n2628_), .B(new_n3208_), .ZN(new_n8523_));
  NOR3_X1    g05799(.A1(new_n5942_), .A2(new_n8089_), .A3(pi0075), .ZN(new_n8524_));
  OAI21_X1   g05800(.A1(new_n8522_), .A2(new_n8523_), .B(new_n8524_), .ZN(new_n8525_));
  AOI21_X1   g05801(.A1(new_n8520_), .A2(new_n3177_), .B(new_n8525_), .ZN(new_n8526_));
  OAI21_X1   g05802(.A1(new_n8516_), .A2(new_n8518_), .B(new_n8526_), .ZN(new_n8527_));
  INV_X1     g05803(.I(new_n8506_), .ZN(new_n8528_));
  NOR3_X1    g05804(.A1(new_n8468_), .A2(pi0100), .A3(new_n8476_), .ZN(new_n8529_));
  AOI21_X1   g05805(.A1(new_n8468_), .A2(new_n3173_), .B(new_n8477_), .ZN(new_n8530_));
  NOR3_X1    g05806(.A1(new_n8529_), .A2(new_n8530_), .A3(pi0039), .ZN(new_n8531_));
  MUX2_X1    g05807(.I0(new_n8531_), .I1(new_n8528_), .S(pi0038), .Z(new_n8532_));
  INV_X1     g05808(.I(new_n5525_), .ZN(new_n8533_));
  NOR2_X1    g05809(.A1(new_n8533_), .A2(pi0100), .ZN(new_n8534_));
  NOR2_X1    g05810(.A1(new_n8534_), .A2(new_n3177_), .ZN(new_n8535_));
  OAI21_X1   g05811(.A1(new_n8528_), .A2(pi0038), .B(pi0100), .ZN(new_n8536_));
  OAI22_X1   g05812(.A1(new_n8532_), .A2(pi0087), .B1(new_n8535_), .B2(new_n8536_), .ZN(new_n8537_));
  MUX2_X1    g05813(.I0(new_n8537_), .I1(new_n8508_), .S(pi0075), .Z(new_n8538_));
  AND2_X2    g05814(.A1(new_n8538_), .A2(new_n5941_), .Z(new_n8539_));
  OAI21_X1   g05815(.A1(new_n8506_), .A2(new_n5941_), .B(new_n8089_), .ZN(new_n8540_));
  OAI21_X1   g05816(.A1(new_n8539_), .A2(new_n8540_), .B(new_n8527_), .ZN(new_n8541_));
  AOI21_X1   g05817(.A1(new_n8541_), .A2(new_n8452_), .B(new_n8514_), .ZN(new_n8542_));
  NOR2_X1    g05818(.A1(new_n5941_), .A2(new_n8089_), .ZN(new_n8543_));
  OAI21_X1   g05819(.A1(new_n8498_), .A2(new_n8543_), .B(new_n6845_), .ZN(new_n8544_));
  OAI21_X1   g05820(.A1(new_n8542_), .A2(new_n8544_), .B(new_n8451_), .ZN(po0210));
  INV_X1     g05821(.I(new_n3378_), .ZN(new_n8546_));
  NAND4_X1   g05822(.A1(new_n2693_), .A2(pi0053), .A3(new_n2682_), .A4(new_n2889_), .ZN(new_n8547_));
  INV_X1     g05823(.I(new_n7827_), .ZN(new_n8548_));
  NAND2_X1   g05824(.A1(new_n8548_), .A2(pi0024), .ZN(new_n8549_));
  OAI21_X1   g05825(.A1(new_n8547_), .A2(new_n8549_), .B(pi0039), .ZN(new_n8550_));
  INV_X1     g05826(.I(new_n5120_), .ZN(new_n8551_));
  NOR2_X1    g05827(.A1(pi0287), .A2(pi0979), .ZN(new_n8552_));
  NOR3_X1    g05828(.A1(new_n8551_), .A2(pi0039), .A3(new_n8552_), .ZN(new_n8553_));
  INV_X1     g05829(.I(new_n8553_), .ZN(new_n8554_));
  NAND2_X1   g05830(.A1(new_n7855_), .A2(new_n8554_), .ZN(new_n8555_));
  AOI21_X1   g05831(.A1(new_n8550_), .A2(new_n8546_), .B(new_n8555_), .ZN(po0211));
  NOR2_X1    g05832(.A1(pi0060), .A2(pi0085), .ZN(new_n8557_));
  NAND4_X1   g05833(.A1(new_n2775_), .A2(new_n7001_), .A3(new_n8557_), .A4(pi0106), .ZN(new_n8558_));
  NOR4_X1    g05834(.A1(new_n7007_), .A2(new_n8376_), .A3(new_n8425_), .A4(new_n8558_), .ZN(new_n8559_));
  NAND2_X1   g05835(.A1(new_n8559_), .A2(new_n8428_), .ZN(new_n8560_));
  NOR4_X1    g05836(.A1(new_n8560_), .A2(pi0053), .A3(new_n7014_), .A4(new_n7440_), .ZN(new_n8561_));
  NOR4_X1    g05837(.A1(new_n2485_), .A2(new_n2644_), .A3(new_n2650_), .A4(pi0841), .ZN(new_n8562_));
  NOR2_X1    g05838(.A1(new_n2629_), .A2(new_n3228_), .ZN(new_n8563_));
  NAND4_X1   g05839(.A1(new_n8561_), .A2(new_n2645_), .A3(new_n8562_), .A4(new_n8563_), .ZN(new_n8564_));
  NOR2_X1    g05840(.A1(new_n7852_), .A2(new_n3208_), .ZN(new_n8565_));
  INV_X1     g05841(.I(new_n8565_), .ZN(new_n8566_));
  NOR2_X1    g05842(.A1(new_n8566_), .A2(new_n3228_), .ZN(new_n8567_));
  INV_X1     g05843(.I(new_n8567_), .ZN(new_n8568_));
  MUX2_X1    g05844(.I0(new_n8568_), .I1(new_n8564_), .S(new_n3214_), .Z(new_n8569_));
  NOR2_X1    g05845(.A1(new_n8569_), .A2(new_n6965_), .ZN(po0212));
  NAND4_X1   g05846(.A1(new_n2775_), .A2(new_n2455_), .A3(pi0045), .A4(new_n2747_), .ZN(new_n8571_));
  NOR4_X1    g05847(.A1(new_n8426_), .A2(new_n8571_), .A3(new_n2499_), .A4(new_n8425_), .ZN(new_n8572_));
  NOR4_X1    g05848(.A1(new_n3234_), .A2(new_n2464_), .A3(new_n2515_), .A4(new_n7430_), .ZN(new_n8573_));
  NAND2_X1   g05849(.A1(new_n8573_), .A2(new_n8572_), .ZN(new_n8574_));
  AOI21_X1   g05850(.A1(new_n8574_), .A2(new_n3227_), .B(new_n6961_), .ZN(new_n8575_));
  NOR4_X1    g05851(.A1(new_n8568_), .A2(pi0054), .A3(new_n6963_), .A4(new_n8575_), .ZN(po0213));
  INV_X1     g05852(.I(new_n5084_), .ZN(new_n8577_));
  NOR4_X1    g05853(.A1(new_n8577_), .A2(pi0056), .A3(new_n7194_), .A4(new_n3336_), .ZN(new_n8578_));
  AOI21_X1   g05854(.A1(pi0056), .A2(new_n3240_), .B(new_n2571_), .ZN(new_n8579_));
  NAND2_X1   g05855(.A1(new_n8578_), .A2(new_n8579_), .ZN(new_n8580_));
  AOI21_X1   g05856(.A1(pi0055), .A2(new_n7806_), .B(new_n8580_), .ZN(po0214));
  NOR2_X1    g05857(.A1(new_n8568_), .A2(pi0054), .ZN(new_n8582_));
  NAND3_X1   g05858(.A1(new_n8582_), .A2(new_n3202_), .A3(new_n5222_), .ZN(new_n8583_));
  NOR3_X1    g05859(.A1(new_n5242_), .A2(new_n7194_), .A3(new_n3336_), .ZN(new_n8584_));
  NOR4_X1    g05860(.A1(new_n8584_), .A2(new_n3335_), .A3(pi0062), .A4(pi0924), .ZN(new_n8585_));
  OAI21_X1   g05861(.A1(new_n8585_), .A2(pi0057), .B(new_n5205_), .ZN(new_n8586_));
  AOI21_X1   g05862(.A1(new_n8583_), .A2(pi0057), .B(new_n8586_), .ZN(po0215));
  INV_X1     g05863(.I(new_n5975_), .ZN(new_n8588_));
  NOR2_X1    g05864(.A1(new_n8588_), .A2(new_n5239_), .ZN(new_n8589_));
  NAND3_X1   g05865(.A1(new_n7824_), .A2(new_n2841_), .A3(new_n8589_), .ZN(new_n8590_));
  NOR3_X1    g05866(.A1(new_n8590_), .A2(new_n5949_), .A3(new_n2839_), .ZN(po0216));
  AND4_X2    g05867(.A1(new_n3335_), .A2(new_n8584_), .A3(pi0062), .A4(pi0924), .Z(new_n8592_));
  OAI21_X1   g05868(.A1(new_n8592_), .A2(pi0059), .B(new_n5055_), .ZN(new_n8593_));
  AOI21_X1   g05869(.A1(new_n8583_), .A2(pi0059), .B(new_n8593_), .ZN(po0217));
  NAND2_X1   g05870(.A1(new_n3181_), .A2(pi0039), .ZN(new_n8595_));
  NOR4_X1    g05871(.A1(new_n8551_), .A2(new_n8595_), .A3(pi0979), .A4(pi1001), .ZN(new_n8596_));
  AND2_X2    g05872(.A1(new_n5358_), .A2(new_n8596_), .Z(new_n8597_));
  NOR2_X1    g05873(.A1(new_n5895_), .A2(pi0039), .ZN(new_n8598_));
  NOR3_X1    g05874(.A1(new_n7014_), .A2(new_n7440_), .A3(pi0053), .ZN(new_n8599_));
  NAND4_X1   g05875(.A1(new_n8599_), .A2(pi0060), .A3(new_n8548_), .A4(new_n8598_), .ZN(new_n8600_));
  OAI21_X1   g05876(.A1(new_n8600_), .A2(new_n2635_), .B(new_n7855_), .ZN(new_n8601_));
  NOR2_X1    g05877(.A1(new_n8601_), .A2(new_n8597_), .ZN(po0218));
  NAND4_X1   g05878(.A1(new_n8599_), .A2(new_n5895_), .A3(pi0060), .A4(new_n2695_), .ZN(new_n8603_));
  OR2_X2     g05879(.A1(new_n8381_), .A2(new_n2902_), .Z(new_n8604_));
  AOI21_X1   g05880(.A1(new_n8603_), .A2(new_n8604_), .B(new_n7829_), .ZN(po0219));
  AOI21_X1   g05881(.A1(new_n8578_), .A2(pi0062), .B(pi0057), .ZN(new_n8606_));
  OAI21_X1   g05882(.A1(new_n7808_), .A2(new_n5055_), .B(new_n5205_), .ZN(new_n8607_));
  NOR2_X1    g05883(.A1(new_n8607_), .A2(new_n8606_), .ZN(po0220));
  INV_X1     g05884(.I(pi0999), .ZN(new_n8609_));
  NAND4_X1   g05885(.A1(new_n7077_), .A2(pi0063), .A3(new_n2800_), .A4(new_n6998_), .ZN(new_n8610_));
  OAI21_X1   g05886(.A1(new_n8609_), .A2(new_n8610_), .B(new_n7828_), .ZN(new_n8611_));
  AOI21_X1   g05887(.A1(new_n8373_), .A2(new_n5895_), .B(new_n8611_), .ZN(po0221));
  NAND3_X1   g05888(.A1(new_n7077_), .A2(new_n2799_), .A3(pi0107), .ZN(new_n8613_));
  NAND3_X1   g05889(.A1(new_n2725_), .A2(new_n2799_), .A3(pi0107), .ZN(new_n8614_));
  NAND4_X1   g05890(.A1(new_n2727_), .A2(new_n2454_), .A3(new_n2634_), .A4(new_n8614_), .ZN(new_n8615_));
  MUX2_X1    g05891(.I0(new_n8615_), .I1(new_n8613_), .S(new_n2902_), .Z(new_n8616_));
  NOR2_X1    g05892(.A1(new_n8616_), .A2(new_n8438_), .ZN(po0222));
  INV_X1     g05893(.I(new_n7869_), .ZN(new_n8618_));
  NOR2_X1    g05894(.A1(new_n7878_), .A2(new_n3154_), .ZN(new_n8619_));
  INV_X1     g05895(.I(new_n8619_), .ZN(new_n8620_));
  NOR4_X1    g05896(.A1(new_n8618_), .A2(new_n7873_), .A3(new_n7856_), .A4(new_n8620_), .ZN(po0223));
  NOR4_X1    g05897(.A1(new_n7430_), .A2(new_n5276_), .A3(new_n7070_), .A4(new_n2515_), .ZN(new_n8622_));
  INV_X1     g05898(.I(new_n8622_), .ZN(new_n8623_));
  NOR4_X1    g05899(.A1(new_n8623_), .A2(new_n2441_), .A3(pi0102), .A4(new_n2699_), .ZN(new_n8624_));
  NOR2_X1    g05900(.A1(new_n3230_), .A2(new_n2622_), .ZN(new_n8625_));
  NOR2_X1    g05901(.A1(new_n8094_), .A2(pi0299), .ZN(new_n8626_));
  NAND4_X1   g05902(.A1(new_n8624_), .A2(new_n2623_), .A3(new_n8625_), .A4(new_n8626_), .ZN(new_n8627_));
  AOI21_X1   g05903(.A1(new_n8627_), .A2(new_n8247_), .B(po1038), .ZN(new_n8628_));
  NAND2_X1   g05904(.A1(new_n8624_), .A2(new_n3233_), .ZN(new_n8629_));
  NOR4_X1    g05905(.A1(new_n8628_), .A2(pi0219), .A3(new_n8169_), .A4(new_n8629_), .ZN(po0224));
  NAND3_X1   g05906(.A1(new_n8440_), .A2(pi0083), .A3(new_n2795_), .ZN(new_n8631_));
  NOR4_X1    g05907(.A1(new_n7825_), .A2(new_n2788_), .A3(new_n8623_), .A4(new_n8631_), .ZN(po0225));
  NOR2_X1    g05908(.A1(new_n5370_), .A2(new_n5145_), .ZN(new_n8633_));
  NOR2_X1    g05909(.A1(new_n3300_), .A2(new_n3294_), .ZN(new_n8634_));
  NOR2_X1    g05910(.A1(new_n5370_), .A2(new_n5866_), .ZN(new_n8635_));
  NOR3_X1    g05911(.A1(new_n7880_), .A2(new_n2562_), .A3(pi0221), .ZN(new_n8636_));
  AOI22_X1   g05912(.A1(new_n8633_), .A2(new_n8634_), .B1(new_n8635_), .B2(new_n8636_), .ZN(new_n8637_));
  NOR2_X1    g05913(.A1(new_n8637_), .A2(new_n8371_), .ZN(po0226));
  NAND3_X1   g05914(.A1(new_n2770_), .A2(pi0069), .A3(new_n2795_), .ZN(new_n8639_));
  OAI21_X1   g05915(.A1(new_n7812_), .A2(new_n8639_), .B(new_n5250_), .ZN(new_n8640_));
  NOR3_X1    g05916(.A1(new_n2464_), .A2(pi0081), .A3(pi0314), .ZN(new_n8641_));
  NAND3_X1   g05917(.A1(new_n8640_), .A2(new_n5249_), .A3(new_n8641_), .ZN(new_n8642_));
  NOR2_X1    g05918(.A1(new_n5250_), .A2(new_n5276_), .ZN(new_n8643_));
  NAND4_X1   g05919(.A1(new_n2722_), .A2(new_n7813_), .A3(new_n5955_), .A4(new_n8643_), .ZN(new_n8644_));
  AOI21_X1   g05920(.A1(new_n8642_), .A2(new_n8644_), .B(new_n8438_), .ZN(po0227));
  NOR4_X1    g05921(.A1(new_n6968_), .A2(pi0051), .A3(new_n2849_), .A4(pi0096), .ZN(new_n8646_));
  NAND3_X1   g05922(.A1(new_n8646_), .A2(new_n3418_), .A3(new_n8598_), .ZN(new_n8647_));
  INV_X1     g05923(.I(new_n5123_), .ZN(new_n8648_));
  INV_X1     g05924(.I(pi0589), .ZN(new_n8649_));
  NOR4_X1    g05925(.A1(new_n5145_), .A2(new_n2601_), .A3(new_n8649_), .A4(new_n3296_), .ZN(new_n8650_));
  NOR3_X1    g05926(.A1(new_n5866_), .A2(new_n3285_), .A3(new_n7880_), .ZN(new_n8651_));
  NOR2_X1    g05927(.A1(new_n2631_), .A2(new_n8649_), .ZN(new_n8652_));
  AOI21_X1   g05928(.A1(new_n8651_), .A2(new_n8652_), .B(new_n8650_), .ZN(new_n8653_));
  OAI21_X1   g05929(.A1(new_n2918_), .A2(new_n2958_), .B(new_n5369_), .ZN(new_n8654_));
  NAND2_X1   g05930(.A1(new_n3082_), .A2(new_n8654_), .ZN(new_n8655_));
  NOR2_X1    g05931(.A1(new_n5118_), .A2(pi0593), .ZN(new_n8656_));
  NAND4_X1   g05932(.A1(new_n8653_), .A2(new_n8648_), .A3(new_n8655_), .A4(new_n8656_), .ZN(new_n8657_));
  NAND2_X1   g05933(.A1(new_n8657_), .A2(new_n8018_), .ZN(new_n8658_));
  NAND2_X1   g05934(.A1(new_n8658_), .A2(new_n3378_), .ZN(new_n8659_));
  AOI21_X1   g05935(.A1(new_n8659_), .A2(new_n8647_), .B(new_n7856_), .ZN(po0228));
  NOR4_X1    g05936(.A1(new_n5252_), .A2(new_n2717_), .A3(new_n2718_), .A4(new_n2758_), .ZN(new_n8661_));
  NOR2_X1    g05937(.A1(new_n8170_), .A2(new_n8098_), .ZN(new_n8662_));
  NOR2_X1    g05938(.A1(new_n8077_), .A2(pi0219), .ZN(new_n8663_));
  INV_X1     g05939(.I(new_n8663_), .ZN(new_n8664_));
  NOR2_X1    g05940(.A1(new_n8664_), .A2(new_n2587_), .ZN(new_n8665_));
  NOR2_X1    g05941(.A1(new_n8665_), .A2(new_n8662_), .ZN(new_n8666_));
  INV_X1     g05942(.I(new_n8666_), .ZN(new_n8667_));
  NOR2_X1    g05943(.A1(new_n8667_), .A2(new_n8388_), .ZN(new_n8668_));
  NAND4_X1   g05944(.A1(new_n8661_), .A2(new_n8389_), .A3(new_n8622_), .A4(new_n8668_), .ZN(new_n8669_));
  NAND4_X1   g05945(.A1(new_n8661_), .A2(new_n2454_), .A3(new_n7005_), .A4(new_n8389_), .ZN(new_n8670_));
  NOR3_X1    g05946(.A1(new_n5269_), .A2(pi0050), .A3(new_n6999_), .ZN(new_n8671_));
  NOR4_X1    g05947(.A1(new_n7827_), .A2(pi0081), .A3(new_n8666_), .A4(new_n5276_), .ZN(new_n8672_));
  NAND3_X1   g05948(.A1(new_n8670_), .A2(new_n8671_), .A3(new_n8672_), .ZN(new_n8673_));
  AOI21_X1   g05949(.A1(new_n8673_), .A2(new_n8669_), .B(new_n7825_), .ZN(po0229));
  NAND2_X1   g05950(.A1(new_n8633_), .A2(new_n6052_), .ZN(new_n8675_));
  NAND4_X1   g05951(.A1(new_n8675_), .A2(new_n6055_), .A3(new_n7856_), .A4(new_n8635_), .ZN(new_n8676_));
  NAND2_X1   g05952(.A1(pi0024), .A2(pi0072), .ZN(new_n8677_));
  NOR2_X1    g05953(.A1(new_n2703_), .A2(pi0098), .ZN(new_n8678_));
  NOR4_X1    g05954(.A1(new_n7819_), .A2(new_n2710_), .A3(new_n7250_), .A4(new_n8654_), .ZN(new_n8679_));
  NAND2_X1   g05955(.A1(new_n8679_), .A2(new_n8678_), .ZN(new_n8680_));
  OAI21_X1   g05956(.A1(new_n2654_), .A2(new_n8677_), .B(new_n8680_), .ZN(new_n8681_));
  AOI21_X1   g05957(.A1(new_n8681_), .A2(new_n2514_), .B(pi0039), .ZN(new_n8682_));
  NOR2_X1    g05958(.A1(new_n8676_), .A2(new_n8682_), .ZN(po0230));
  INV_X1     g05959(.I(pi1050), .ZN(new_n8684_));
  NOR2_X1    g05960(.A1(new_n7233_), .A2(new_n7827_), .ZN(new_n8685_));
  INV_X1     g05961(.I(new_n8685_), .ZN(new_n8686_));
  NOR3_X1    g05962(.A1(new_n8686_), .A2(pi0314), .A3(new_n8684_), .ZN(new_n8687_));
  AOI21_X1   g05963(.A1(new_n8635_), .A2(new_n7170_), .B(new_n2587_), .ZN(new_n8688_));
  NAND2_X1   g05964(.A1(new_n8633_), .A2(new_n7153_), .ZN(new_n8689_));
  AOI21_X1   g05965(.A1(new_n2587_), .A2(new_n8689_), .B(new_n8688_), .ZN(new_n8690_));
  INV_X1     g05966(.I(new_n8690_), .ZN(new_n8691_));
  OR3_X2     g05967(.A1(new_n8691_), .A2(new_n3154_), .A3(new_n8687_), .Z(new_n8692_));
  OAI21_X1   g05968(.A1(new_n8690_), .A2(new_n3154_), .B(new_n8687_), .ZN(new_n8693_));
  AOI21_X1   g05969(.A1(new_n8692_), .A2(new_n8693_), .B(new_n7856_), .ZN(po0231));
  INV_X1     g05970(.I(new_n2666_), .ZN(new_n8695_));
  NOR3_X1    g05971(.A1(new_n6023_), .A2(new_n5239_), .A3(new_n8695_), .ZN(new_n8696_));
  NOR2_X1    g05972(.A1(new_n8696_), .A2(pi0096), .ZN(new_n8697_));
  OAI21_X1   g05973(.A1(new_n5081_), .A2(pi0096), .B(pi0479), .ZN(new_n8698_));
  NAND2_X1   g05974(.A1(new_n6979_), .A2(new_n8698_), .ZN(new_n8699_));
  NAND3_X1   g05975(.A1(new_n6004_), .A2(new_n2659_), .A3(new_n2924_), .ZN(new_n8700_));
  NAND4_X1   g05976(.A1(new_n8699_), .A2(new_n3322_), .A3(new_n5941_), .A4(new_n8700_), .ZN(new_n8701_));
  OR3_X2     g05977(.A1(new_n5973_), .A2(new_n8697_), .A3(new_n8701_), .Z(new_n8702_));
  NAND2_X1   g05978(.A1(new_n8582_), .A2(pi0074), .ZN(new_n8703_));
  AOI21_X1   g05979(.A1(new_n8703_), .A2(new_n8702_), .B(po1038), .ZN(po0232));
  OAI22_X1   g05980(.A1(new_n8697_), .A2(new_n2960_), .B1(new_n2659_), .B2(pi1093), .ZN(new_n8705_));
  NAND3_X1   g05981(.A1(new_n8705_), .A2(new_n2625_), .A3(new_n6027_), .ZN(new_n8706_));
  NOR4_X1    g05982(.A1(new_n8566_), .A2(pi0075), .A3(new_n6966_), .A4(new_n8706_), .ZN(po0233));
  NOR3_X1    g05983(.A1(new_n7847_), .A2(new_n2507_), .A3(new_n7012_), .ZN(new_n8708_));
  INV_X1     g05984(.I(new_n8708_), .ZN(new_n8709_));
  NOR3_X1    g05985(.A1(new_n8709_), .A2(po1057), .A3(new_n7779_), .ZN(new_n8710_));
  NAND2_X1   g05986(.A1(new_n7985_), .A2(new_n3418_), .ZN(new_n8711_));
  AOI21_X1   g05987(.A1(pi0252), .A2(new_n2956_), .B(new_n8711_), .ZN(new_n8712_));
  NAND2_X1   g05988(.A1(new_n7984_), .A2(new_n7014_), .ZN(new_n8713_));
  AOI21_X1   g05989(.A1(new_n7016_), .A2(new_n2466_), .B(new_n7827_), .ZN(new_n8714_));
  NAND2_X1   g05990(.A1(new_n8713_), .A2(new_n8714_), .ZN(new_n8715_));
  INV_X1     g05991(.I(new_n8715_), .ZN(new_n8716_));
  NOR4_X1    g05992(.A1(new_n8716_), .A2(new_n3181_), .A3(new_n2956_), .A4(new_n8708_), .ZN(new_n8717_));
  NOR2_X1    g05993(.A1(new_n8716_), .A2(new_n2956_), .ZN(new_n8718_));
  NOR2_X1    g05994(.A1(new_n8717_), .A2(new_n8718_), .ZN(new_n8719_));
  NOR2_X1    g05995(.A1(new_n8719_), .A2(new_n6029_), .ZN(new_n8720_));
  OAI21_X1   g05996(.A1(new_n8712_), .A2(pi0122), .B(new_n2924_), .ZN(new_n8721_));
  INV_X1     g05997(.I(new_n8719_), .ZN(new_n8722_));
  INV_X1     g05998(.I(new_n8711_), .ZN(new_n8723_));
  AOI21_X1   g05999(.A1(new_n6004_), .A2(new_n8718_), .B(new_n8717_), .ZN(new_n8724_));
  OR3_X2     g06000(.A1(new_n8724_), .A2(new_n5181_), .A3(new_n8723_), .Z(new_n8725_));
  AOI21_X1   g06001(.A1(new_n8725_), .A2(new_n6029_), .B(new_n8722_), .ZN(new_n8726_));
  NOR3_X1    g06002(.A1(new_n8725_), .A2(pi0122), .A3(new_n8719_), .ZN(new_n8727_));
  NOR3_X1    g06003(.A1(new_n8727_), .A2(new_n8726_), .A3(pi1093), .ZN(new_n8728_));
  OAI21_X1   g06004(.A1(new_n8720_), .A2(new_n8721_), .B(new_n8728_), .ZN(new_n8729_));
  NOR4_X1    g06005(.A1(new_n8729_), .A2(new_n2436_), .A3(new_n2922_), .A4(new_n8712_), .ZN(new_n8730_));
  NAND4_X1   g06006(.A1(new_n8711_), .A2(new_n8715_), .A3(pi0122), .A4(new_n2924_), .ZN(new_n8731_));
  NAND2_X1   g06007(.A1(new_n8728_), .A2(new_n8731_), .ZN(new_n8732_));
  NAND2_X1   g06008(.A1(new_n8732_), .A2(new_n2922_), .ZN(new_n8733_));
  NOR2_X1    g06009(.A1(new_n2921_), .A2(pi0137), .ZN(new_n8734_));
  INV_X1     g06010(.I(new_n8734_), .ZN(new_n8735_));
  NOR3_X1    g06011(.A1(new_n3181_), .A2(new_n2923_), .A3(pi1093), .ZN(new_n8736_));
  NAND2_X1   g06012(.A1(new_n8736_), .A2(new_n2929_), .ZN(new_n8737_));
  NAND2_X1   g06013(.A1(new_n8737_), .A2(new_n2436_), .ZN(new_n8738_));
  AOI22_X1   g06014(.A1(new_n8733_), .A2(new_n8735_), .B1(new_n8723_), .B2(new_n8738_), .ZN(new_n8739_));
  NOR2_X1    g06015(.A1(new_n8739_), .A2(new_n8730_), .ZN(new_n8740_));
  INV_X1     g06016(.I(new_n8740_), .ZN(new_n8741_));
  MUX2_X1    g06017(.I0(new_n8741_), .I1(new_n2436_), .S(po1057), .Z(new_n8742_));
  NOR2_X1    g06018(.A1(new_n8742_), .A2(new_n8710_), .ZN(new_n8743_));
  NAND2_X1   g06019(.A1(new_n8743_), .A2(new_n2601_), .ZN(new_n8744_));
  NAND2_X1   g06020(.A1(new_n8729_), .A2(new_n2921_), .ZN(new_n8745_));
  NAND2_X1   g06021(.A1(new_n8745_), .A2(new_n8733_), .ZN(new_n8746_));
  INV_X1     g06022(.I(new_n8746_), .ZN(new_n8747_));
  NOR2_X1    g06023(.A1(new_n8747_), .A2(po1057), .ZN(new_n8748_));
  OR3_X2     g06024(.A1(new_n8748_), .A2(new_n2601_), .A3(new_n8710_), .Z(new_n8749_));
  NAND2_X1   g06025(.A1(new_n8744_), .A2(new_n8749_), .ZN(new_n8750_));
  INV_X1     g06026(.I(new_n8750_), .ZN(new_n8751_));
  NAND2_X1   g06027(.A1(new_n8747_), .A2(pi0198), .ZN(new_n8752_));
  OAI21_X1   g06028(.A1(new_n8741_), .A2(pi0198), .B(new_n8752_), .ZN(new_n8753_));
  NAND4_X1   g06029(.A1(new_n8751_), .A2(new_n2605_), .A3(new_n5108_), .A4(new_n8753_), .ZN(new_n8754_));
  NAND2_X1   g06030(.A1(new_n2605_), .A2(new_n5108_), .ZN(new_n8755_));
  OAI21_X1   g06031(.A1(new_n8755_), .A2(new_n8753_), .B(new_n8750_), .ZN(new_n8756_));
  AOI21_X1   g06032(.A1(new_n8754_), .A2(new_n8756_), .B(pi0299), .ZN(new_n8757_));
  NOR2_X1    g06033(.A1(new_n8163_), .A2(new_n2575_), .ZN(new_n8758_));
  NOR3_X1    g06034(.A1(new_n8748_), .A2(new_n2631_), .A3(new_n8710_), .ZN(new_n8759_));
  AOI21_X1   g06035(.A1(new_n8743_), .A2(new_n2631_), .B(new_n8759_), .ZN(new_n8760_));
  NAND2_X1   g06036(.A1(new_n8760_), .A2(new_n8758_), .ZN(new_n8761_));
  NOR2_X1    g06037(.A1(new_n8741_), .A2(pi0210), .ZN(new_n8762_));
  NOR2_X1    g06038(.A1(new_n8746_), .A2(new_n2631_), .ZN(new_n8763_));
  OAI21_X1   g06039(.A1(new_n8762_), .A2(new_n8763_), .B(new_n8758_), .ZN(new_n8764_));
  AOI21_X1   g06040(.A1(new_n8761_), .A2(new_n8764_), .B(new_n2587_), .ZN(new_n8765_));
  OAI21_X1   g06041(.A1(new_n8757_), .A2(new_n8765_), .B(pi0232), .ZN(new_n8766_));
  NAND2_X1   g06042(.A1(new_n8751_), .A2(new_n2587_), .ZN(new_n8767_));
  AOI21_X1   g06043(.A1(new_n8760_), .A2(pi0299), .B(pi0232), .ZN(new_n8768_));
  AOI21_X1   g06044(.A1(new_n8767_), .A2(new_n8768_), .B(new_n6844_), .ZN(new_n8769_));
  NAND2_X1   g06045(.A1(new_n8766_), .A2(new_n8769_), .ZN(new_n8770_));
  INV_X1     g06046(.I(new_n6978_), .ZN(new_n8771_));
  NOR2_X1    g06047(.A1(new_n8771_), .A2(pi0137), .ZN(new_n8772_));
  AOI21_X1   g06048(.A1(po1057), .A2(new_n8772_), .B(new_n2921_), .ZN(new_n8773_));
  NOR2_X1    g06049(.A1(new_n8715_), .A2(new_n2924_), .ZN(new_n8774_));
  NOR2_X1    g06050(.A1(new_n8711_), .A2(pi0252), .ZN(new_n8775_));
  MUX2_X1    g06051(.I0(new_n8775_), .I1(new_n8716_), .S(new_n2957_), .Z(new_n8776_));
  INV_X1     g06052(.I(new_n8776_), .ZN(new_n8777_));
  AOI21_X1   g06053(.A1(new_n8777_), .A2(new_n2436_), .B(pi1093), .ZN(new_n8778_));
  NOR2_X1    g06054(.A1(new_n8719_), .A2(pi1093), .ZN(new_n8779_));
  INV_X1     g06055(.I(new_n8779_), .ZN(new_n8780_));
  OAI22_X1   g06056(.A1(new_n8774_), .A2(new_n8778_), .B1(new_n8780_), .B2(new_n2436_), .ZN(new_n8781_));
  OAI21_X1   g06057(.A1(new_n8781_), .A2(new_n8708_), .B(po1057), .ZN(new_n8782_));
  NOR2_X1    g06058(.A1(new_n8782_), .A2(new_n8773_), .ZN(new_n8783_));
  NAND2_X1   g06059(.A1(new_n8777_), .A2(new_n6424_), .ZN(new_n8784_));
  XOR2_X1    g06060(.A1(new_n8784_), .A2(new_n8720_), .Z(new_n8785_));
  NOR2_X1    g06061(.A1(new_n8785_), .A2(new_n8779_), .ZN(new_n8786_));
  MUX2_X1    g06062(.I0(new_n8786_), .I1(new_n8776_), .S(new_n2436_), .Z(new_n8787_));
  INV_X1     g06063(.I(new_n8787_), .ZN(new_n8788_));
  OAI21_X1   g06064(.A1(new_n2436_), .A2(new_n6424_), .B(new_n2956_), .ZN(new_n8789_));
  NAND2_X1   g06065(.A1(new_n8789_), .A2(new_n2922_), .ZN(new_n8790_));
  NOR4_X1    g06066(.A1(new_n8788_), .A2(po1057), .A3(new_n8709_), .A4(new_n8790_), .ZN(new_n8791_));
  NOR2_X1    g06067(.A1(new_n8791_), .A2(new_n8783_), .ZN(new_n8792_));
  NOR2_X1    g06068(.A1(new_n8792_), .A2(pi0198), .ZN(new_n8793_));
  OAI21_X1   g06069(.A1(new_n2922_), .A2(new_n6436_), .B(new_n8708_), .ZN(new_n8794_));
  NAND2_X1   g06070(.A1(new_n8715_), .A2(pi1093), .ZN(new_n8795_));
  NOR3_X1    g06071(.A1(new_n8785_), .A2(new_n2921_), .A3(new_n8795_), .ZN(new_n8796_));
  INV_X1     g06072(.I(new_n8785_), .ZN(new_n8797_));
  AOI21_X1   g06073(.A1(new_n2922_), .A2(new_n8795_), .B(new_n8797_), .ZN(new_n8798_));
  NOR3_X1    g06074(.A1(new_n8798_), .A2(new_n8796_), .A3(new_n8779_), .ZN(new_n8799_));
  MUX2_X1    g06075(.I0(new_n8799_), .I1(new_n8794_), .S(po1057), .Z(new_n8800_));
  NOR2_X1    g06076(.A1(new_n8800_), .A2(new_n2601_), .ZN(new_n8801_));
  NOR2_X1    g06077(.A1(new_n8793_), .A2(new_n8801_), .ZN(new_n8802_));
  NOR2_X1    g06078(.A1(new_n8787_), .A2(new_n2922_), .ZN(new_n8803_));
  AOI21_X1   g06079(.A1(new_n2922_), .A2(new_n8781_), .B(new_n8803_), .ZN(new_n8804_));
  NOR2_X1    g06080(.A1(new_n8804_), .A2(pi0198), .ZN(new_n8805_));
  AOI21_X1   g06081(.A1(pi0198), .A2(new_n8799_), .B(new_n8805_), .ZN(new_n8806_));
  MUX2_X1    g06082(.I0(new_n8806_), .I1(new_n8802_), .S(new_n8755_), .Z(new_n8807_));
  OAI21_X1   g06083(.A1(new_n8791_), .A2(new_n8783_), .B(new_n2631_), .ZN(new_n8808_));
  OAI21_X1   g06084(.A1(new_n2631_), .A2(new_n8800_), .B(new_n8808_), .ZN(new_n8809_));
  MUX2_X1    g06085(.I0(new_n8804_), .I1(new_n8799_), .S(new_n2631_), .Z(new_n8810_));
  AOI21_X1   g06086(.A1(new_n8809_), .A2(new_n8810_), .B(new_n8758_), .ZN(new_n8811_));
  NAND2_X1   g06087(.A1(new_n8811_), .A2(new_n2587_), .ZN(new_n8812_));
  OAI21_X1   g06088(.A1(new_n8807_), .A2(pi0299), .B(new_n8812_), .ZN(new_n8813_));
  NOR3_X1    g06089(.A1(new_n8793_), .A2(pi0299), .A3(new_n8801_), .ZN(new_n8814_));
  OAI21_X1   g06090(.A1(new_n8809_), .A2(new_n2587_), .B(new_n5987_), .ZN(new_n8815_));
  OAI21_X1   g06091(.A1(new_n8815_), .A2(new_n8814_), .B(new_n6844_), .ZN(new_n8816_));
  AOI21_X1   g06092(.A1(new_n8813_), .A2(new_n5987_), .B(new_n8816_), .ZN(new_n8817_));
  AOI21_X1   g06093(.A1(new_n8770_), .A2(new_n8817_), .B(new_n7825_), .ZN(po0234));
  AOI21_X1   g06094(.A1(new_n2707_), .A2(new_n2684_), .B(pi0086), .ZN(new_n8819_));
  NOR3_X1    g06095(.A1(new_n5278_), .A2(new_n2640_), .A3(new_n8819_), .ZN(new_n8820_));
  INV_X1     g06096(.I(new_n8820_), .ZN(new_n8821_));
  NOR3_X1    g06097(.A1(new_n2819_), .A2(new_n2691_), .A3(new_n7014_), .ZN(new_n8822_));
  OAI21_X1   g06098(.A1(new_n8821_), .A2(new_n8822_), .B(pi0314), .ZN(new_n8823_));
  NOR2_X1    g06099(.A1(new_n8823_), .A2(new_n7829_), .ZN(po0235));
  NOR3_X1    g06100(.A1(new_n5929_), .A2(new_n5987_), .A3(pi0468), .ZN(po0236));
  INV_X1     g06101(.I(pi0163), .ZN(new_n8826_));
  NAND4_X1   g06102(.A1(new_n5108_), .A2(new_n7326_), .A3(pi0162), .A4(pi0197), .ZN(new_n8827_));
  NOR2_X1    g06103(.A1(pi0162), .A2(pi0197), .ZN(new_n8828_));
  NOR3_X1    g06104(.A1(new_n5109_), .A2(new_n7326_), .A3(new_n8828_), .ZN(new_n8829_));
  INV_X1     g06105(.I(new_n8829_), .ZN(new_n8830_));
  NAND2_X1   g06106(.A1(new_n5109_), .A2(pi0163), .ZN(new_n8831_));
  NAND3_X1   g06107(.A1(new_n8830_), .A2(new_n8827_), .A3(new_n8831_), .ZN(new_n8832_));
  XOR2_X1    g06108(.A1(new_n8832_), .A2(new_n8826_), .Z(new_n8833_));
  NOR2_X1    g06109(.A1(new_n8833_), .A2(new_n5987_), .ZN(new_n8834_));
  AOI21_X1   g06110(.A1(new_n8834_), .A2(new_n7048_), .B(new_n3202_), .ZN(new_n8835_));
  INV_X1     g06111(.I(pi0147), .ZN(new_n8836_));
  NOR4_X1    g06112(.A1(new_n8834_), .A2(new_n8836_), .A3(new_n7041_), .A4(new_n7050_), .ZN(new_n8837_));
  INV_X1     g06113(.I(new_n8837_), .ZN(new_n8838_));
  NOR3_X1    g06114(.A1(new_n8838_), .A2(new_n8835_), .A3(new_n2571_), .ZN(new_n8839_));
  NOR2_X1    g06115(.A1(new_n8837_), .A2(new_n3214_), .ZN(new_n8840_));
  NOR2_X1    g06116(.A1(new_n8834_), .A2(new_n3173_), .ZN(new_n8841_));
  NOR2_X1    g06117(.A1(pi0038), .A2(pi0040), .ZN(new_n8842_));
  NOR3_X1    g06118(.A1(new_n5989_), .A2(pi0038), .A3(new_n8836_), .ZN(new_n8843_));
  NOR2_X1    g06119(.A1(new_n8843_), .A2(pi0100), .ZN(new_n8844_));
  NOR2_X1    g06120(.A1(new_n8844_), .A2(new_n8842_), .ZN(new_n8845_));
  NOR2_X1    g06121(.A1(new_n8841_), .A2(new_n8845_), .ZN(new_n8846_));
  AOI21_X1   g06122(.A1(new_n8834_), .A2(pi0075), .B(pi0054), .ZN(new_n8847_));
  OAI21_X1   g06123(.A1(new_n8846_), .A2(new_n2628_), .B(new_n8847_), .ZN(new_n8848_));
  OAI21_X1   g06124(.A1(new_n8848_), .A2(new_n8840_), .B(new_n3202_), .ZN(new_n8849_));
  NOR2_X1    g06125(.A1(new_n8835_), .A2(new_n2533_), .ZN(new_n8850_));
  AOI21_X1   g06126(.A1(new_n8849_), .A2(new_n8850_), .B(new_n3405_), .ZN(new_n8851_));
  INV_X1     g06127(.I(new_n8851_), .ZN(new_n8852_));
  INV_X1     g06128(.I(new_n8833_), .ZN(new_n8853_));
  NOR4_X1    g06129(.A1(new_n7342_), .A2(pi0184), .A3(new_n5109_), .A4(new_n7343_), .ZN(new_n8854_));
  NAND2_X1   g06130(.A1(new_n7341_), .A2(new_n7344_), .ZN(new_n8855_));
  NAND3_X1   g06131(.A1(new_n8855_), .A2(pi0184), .A3(new_n5108_), .ZN(new_n8856_));
  NAND2_X1   g06132(.A1(new_n8856_), .A2(new_n7348_), .ZN(new_n8857_));
  NOR2_X1    g06133(.A1(new_n8857_), .A2(new_n8854_), .ZN(new_n8858_));
  NAND2_X1   g06134(.A1(new_n8853_), .A2(new_n8858_), .ZN(new_n8859_));
  INV_X1     g06135(.I(new_n8859_), .ZN(new_n8860_));
  INV_X1     g06136(.I(pi0187), .ZN(new_n8861_));
  MUX2_X1    g06137(.I0(new_n8861_), .I1(new_n8836_), .S(pi0299), .Z(new_n8862_));
  NOR2_X1    g06138(.A1(new_n5989_), .A2(new_n8862_), .ZN(new_n8863_));
  MUX2_X1    g06139(.I0(new_n8863_), .I1(new_n8860_), .S(new_n7041_), .Z(new_n8864_));
  NAND2_X1   g06140(.A1(new_n8864_), .A2(new_n3214_), .ZN(new_n8865_));
  NOR4_X1    g06141(.A1(new_n7390_), .A2(pi0040), .A3(pi0095), .A4(pi0479), .ZN(new_n8866_));
  INV_X1     g06142(.I(new_n8866_), .ZN(new_n8867_));
  NOR2_X1    g06143(.A1(new_n7560_), .A2(pi0040), .ZN(new_n8868_));
  OAI21_X1   g06144(.A1(new_n8868_), .A2(pi0095), .B(new_n8867_), .ZN(new_n8869_));
  INV_X1     g06145(.I(new_n8869_), .ZN(new_n8870_));
  NOR2_X1    g06146(.A1(pi0175), .A2(pi0299), .ZN(new_n8871_));
  INV_X1     g06147(.I(pi0189), .ZN(new_n8872_));
  NOR2_X1    g06148(.A1(new_n5109_), .A2(new_n8872_), .ZN(new_n8873_));
  OAI21_X1   g06149(.A1(new_n7445_), .A2(pi0040), .B(new_n2632_), .ZN(new_n8874_));
  AOI21_X1   g06150(.A1(new_n8874_), .A2(new_n7476_), .B(pi0095), .ZN(new_n8875_));
  OR2_X2     g06151(.A1(new_n8875_), .A2(new_n7479_), .Z(new_n8876_));
  AOI21_X1   g06152(.A1(new_n8874_), .A2(new_n7535_), .B(pi0095), .ZN(new_n8877_));
  NOR2_X1    g06153(.A1(new_n8877_), .A2(new_n7479_), .ZN(new_n8878_));
  OAI21_X1   g06154(.A1(new_n8876_), .A2(new_n8878_), .B(pi0198), .ZN(new_n8879_));
  NOR2_X1    g06155(.A1(new_n5326_), .A2(pi0184), .ZN(new_n8880_));
  OAI21_X1   g06156(.A1(new_n8879_), .A2(new_n8012_), .B(new_n8880_), .ZN(new_n8881_));
  AOI21_X1   g06157(.A1(new_n8868_), .A2(new_n8873_), .B(new_n8881_), .ZN(new_n8882_));
  INV_X1     g06158(.I(pi0184), .ZN(new_n8883_));
  OAI21_X1   g06159(.A1(new_n7417_), .A2(pi0040), .B(new_n2437_), .ZN(new_n8884_));
  NAND2_X1   g06160(.A1(new_n7425_), .A2(new_n3364_), .ZN(new_n8885_));
  NOR4_X1    g06161(.A1(new_n8866_), .A2(new_n5326_), .A3(new_n5108_), .A4(new_n7479_), .ZN(new_n8886_));
  NOR3_X1    g06162(.A1(new_n8885_), .A2(new_n8872_), .A3(new_n8886_), .ZN(new_n8887_));
  AOI21_X1   g06163(.A1(new_n8887_), .A2(new_n8884_), .B(new_n8883_), .ZN(new_n8888_));
  OAI21_X1   g06164(.A1(new_n8882_), .A2(new_n8888_), .B(new_n8871_), .ZN(new_n8889_));
  NAND3_X1   g06165(.A1(new_n7477_), .A2(new_n2437_), .A3(new_n8867_), .ZN(new_n8890_));
  AOI21_X1   g06166(.A1(new_n7470_), .A2(new_n2437_), .B(new_n8866_), .ZN(new_n8891_));
  XNOR2_X1   g06167(.A1(new_n8891_), .A2(new_n8890_), .ZN(new_n8892_));
  NAND2_X1   g06168(.A1(new_n8892_), .A2(pi0198), .ZN(new_n8893_));
  XOR2_X1    g06169(.A1(new_n8893_), .A2(new_n8890_), .Z(new_n8894_));
  NAND2_X1   g06170(.A1(new_n8894_), .A2(new_n8873_), .ZN(new_n8895_));
  INV_X1     g06171(.I(new_n8873_), .ZN(new_n8896_));
  NAND2_X1   g06172(.A1(new_n7467_), .A2(pi0095), .ZN(new_n8897_));
  OAI21_X1   g06173(.A1(new_n7470_), .A2(pi0095), .B(new_n8897_), .ZN(new_n8898_));
  OAI21_X1   g06174(.A1(new_n7481_), .A2(new_n8898_), .B(pi0198), .ZN(new_n8899_));
  OAI22_X1   g06175(.A1(new_n8899_), .A2(new_n8896_), .B1(new_n7538_), .B2(new_n8012_), .ZN(new_n8900_));
  INV_X1     g06176(.I(new_n8900_), .ZN(new_n8901_));
  AOI21_X1   g06177(.A1(pi0182), .A2(new_n8901_), .B(new_n8895_), .ZN(new_n8902_));
  NAND3_X1   g06178(.A1(new_n8895_), .A2(pi0182), .A3(new_n8900_), .ZN(new_n8903_));
  NAND2_X1   g06179(.A1(new_n5326_), .A2(pi0095), .ZN(new_n8904_));
  AND2_X2    g06180(.A1(new_n7538_), .A2(new_n8904_), .Z(new_n8905_));
  OAI21_X1   g06181(.A1(new_n8905_), .A2(new_n8866_), .B(new_n8012_), .ZN(new_n8906_));
  NAND3_X1   g06182(.A1(new_n8903_), .A2(new_n8883_), .A3(new_n8906_), .ZN(new_n8907_));
  NAND2_X1   g06183(.A1(new_n8866_), .A2(new_n5326_), .ZN(new_n8908_));
  OAI21_X1   g06184(.A1(pi0095), .A2(new_n8872_), .B(new_n2455_), .ZN(new_n8909_));
  NOR2_X1    g06185(.A1(new_n7431_), .A2(pi0040), .ZN(new_n8910_));
  NAND3_X1   g06186(.A1(new_n8904_), .A2(pi0184), .A3(new_n5108_), .ZN(new_n8911_));
  AOI21_X1   g06187(.A1(new_n8910_), .A2(new_n8909_), .B(new_n8911_), .ZN(new_n8912_));
  INV_X1     g06188(.I(pi0175), .ZN(new_n8913_));
  NOR2_X1    g06189(.A1(new_n8913_), .A2(pi0299), .ZN(new_n8914_));
  INV_X1     g06190(.I(new_n8914_), .ZN(new_n8915_));
  AOI21_X1   g06191(.A1(new_n8908_), .A2(new_n8912_), .B(new_n8915_), .ZN(new_n8916_));
  OAI21_X1   g06192(.A1(new_n8907_), .A2(new_n8902_), .B(new_n8916_), .ZN(new_n8917_));
  AOI22_X1   g06193(.A1(new_n8917_), .A2(new_n8889_), .B1(new_n5109_), .B2(new_n8870_), .ZN(new_n8918_));
  NOR2_X1    g06194(.A1(new_n7573_), .A2(pi0040), .ZN(new_n8919_));
  OAI21_X1   g06195(.A1(new_n8919_), .A2(pi0095), .B(new_n8867_), .ZN(new_n8920_));
  INV_X1     g06196(.I(new_n8920_), .ZN(new_n8921_));
  NAND2_X1   g06197(.A1(new_n8921_), .A2(pi0166), .ZN(new_n8922_));
  NOR2_X1    g06198(.A1(new_n8875_), .A2(new_n8866_), .ZN(new_n8923_));
  NOR2_X1    g06199(.A1(new_n8877_), .A2(new_n8866_), .ZN(new_n8924_));
  MUX2_X1    g06200(.I0(new_n8924_), .I1(new_n8923_), .S(new_n2631_), .Z(new_n8925_));
  AOI21_X1   g06201(.A1(new_n8925_), .A2(new_n7928_), .B(pi0153), .ZN(new_n8926_));
  NOR2_X1    g06202(.A1(new_n7928_), .A2(new_n2631_), .ZN(new_n8927_));
  OAI21_X1   g06203(.A1(new_n7536_), .A2(new_n8866_), .B(new_n8927_), .ZN(new_n8928_));
  NOR2_X1    g06204(.A1(new_n7532_), .A2(new_n8866_), .ZN(new_n8929_));
  NOR2_X1    g06205(.A1(new_n8929_), .A2(pi0210), .ZN(new_n8930_));
  NOR2_X1    g06206(.A1(new_n5109_), .A2(new_n4549_), .ZN(new_n8931_));
  NAND2_X1   g06207(.A1(new_n8892_), .A2(pi0210), .ZN(new_n8932_));
  XOR2_X1    g06208(.A1(new_n8932_), .A2(new_n8890_), .Z(new_n8933_));
  AOI22_X1   g06209(.A1(new_n8933_), .A2(new_n8931_), .B1(new_n8928_), .B2(new_n8930_), .ZN(new_n8934_));
  OAI21_X1   g06210(.A1(new_n8934_), .A2(pi0153), .B(new_n5338_), .ZN(new_n8935_));
  AOI21_X1   g06211(.A1(new_n8922_), .A2(new_n8926_), .B(new_n8935_), .ZN(new_n8936_));
  NOR2_X1    g06212(.A1(new_n7536_), .A2(new_n7479_), .ZN(new_n8937_));
  MUX2_X1    g06213(.I0(new_n8937_), .I1(new_n7533_), .S(new_n2631_), .Z(new_n8938_));
  NAND2_X1   g06214(.A1(new_n8938_), .A2(new_n7928_), .ZN(new_n8939_));
  NOR2_X1    g06215(.A1(new_n7480_), .A2(new_n2631_), .ZN(new_n8940_));
  AND2_X2    g06216(.A1(new_n8898_), .A2(pi0210), .Z(new_n8941_));
  OAI21_X1   g06217(.A1(new_n8940_), .A2(new_n8941_), .B(new_n8931_), .ZN(new_n8942_));
  NAND2_X1   g06218(.A1(new_n2526_), .A2(new_n5338_), .ZN(new_n8943_));
  AOI21_X1   g06219(.A1(new_n8942_), .A2(new_n8939_), .B(new_n8943_), .ZN(new_n8944_));
  NAND4_X1   g06220(.A1(new_n8919_), .A2(pi0153), .A3(pi0166), .A4(new_n5108_), .ZN(new_n8946_));
  NOR2_X1    g06221(.A1(new_n8885_), .A2(new_n4549_), .ZN(new_n8947_));
  NOR2_X1    g06222(.A1(new_n8947_), .A2(new_n8884_), .ZN(new_n8948_));
  OAI21_X1   g06223(.A1(new_n8948_), .A2(new_n7479_), .B(new_n5109_), .ZN(new_n8949_));
  INV_X1     g06224(.I(new_n8931_), .ZN(new_n8950_));
  NOR2_X1    g06225(.A1(new_n8950_), .A2(new_n7479_), .ZN(new_n8951_));
  OAI21_X1   g06226(.A1(new_n8910_), .A2(pi0095), .B(new_n8951_), .ZN(new_n8952_));
  NOR3_X1    g06227(.A1(new_n8163_), .A2(pi0153), .A3(new_n7468_), .ZN(new_n8953_));
  AOI21_X1   g06228(.A1(new_n8952_), .A2(new_n8953_), .B(pi0153), .ZN(new_n8954_));
  NAND2_X1   g06229(.A1(new_n8949_), .A2(new_n8954_), .ZN(new_n8955_));
  OAI22_X1   g06230(.A1(new_n8686_), .A2(pi0166), .B1(pi0095), .B2(new_n8910_), .ZN(new_n8956_));
  NAND2_X1   g06231(.A1(new_n5108_), .A2(new_n5338_), .ZN(new_n8957_));
  AOI21_X1   g06232(.A1(new_n8956_), .A2(pi0153), .B(new_n8957_), .ZN(new_n8958_));
  NAND2_X1   g06233(.A1(new_n2526_), .A2(new_n8826_), .ZN(new_n8959_));
  AOI21_X1   g06234(.A1(new_n8867_), .A2(new_n8958_), .B(new_n8959_), .ZN(new_n8960_));
  AOI21_X1   g06235(.A1(new_n8948_), .A2(new_n8960_), .B(pi0160), .ZN(new_n8961_));
  AOI21_X1   g06236(.A1(new_n8955_), .A2(new_n8961_), .B(pi0163), .ZN(new_n8962_));
  OAI21_X1   g06237(.A1(new_n8946_), .A2(new_n8944_), .B(new_n8962_), .ZN(new_n8963_));
  MUX2_X1    g06238(.I0(new_n8924_), .I1(new_n8923_), .S(new_n2601_), .Z(new_n8964_));
  NAND2_X1   g06239(.A1(new_n8964_), .A2(new_n8011_), .ZN(new_n8965_));
  NOR2_X1    g06240(.A1(pi0182), .A2(pi0184), .ZN(new_n8966_));
  NAND3_X1   g06241(.A1(new_n8965_), .A2(new_n8871_), .A3(new_n8966_), .ZN(new_n8967_));
  NOR2_X1    g06242(.A1(new_n8869_), .A2(new_n8011_), .ZN(new_n8968_));
  OAI21_X1   g06243(.A1(new_n8920_), .A2(new_n5108_), .B(new_n5854_), .ZN(new_n8969_));
  AOI21_X1   g06244(.A1(new_n8967_), .A2(new_n8968_), .B(new_n8969_), .ZN(new_n8970_));
  OAI21_X1   g06245(.A1(new_n8936_), .A2(new_n8963_), .B(new_n8970_), .ZN(new_n8971_));
  AOI21_X1   g06246(.A1(new_n2587_), .A2(new_n8869_), .B(new_n8920_), .ZN(new_n8972_));
  NOR3_X1    g06247(.A1(new_n8921_), .A2(pi0299), .A3(new_n8869_), .ZN(new_n8973_));
  INV_X1     g06248(.I(pi0156), .ZN(new_n8974_));
  NOR3_X1    g06249(.A1(new_n7634_), .A2(pi0299), .A3(new_n7467_), .ZN(new_n8975_));
  NOR2_X1    g06250(.A1(new_n5143_), .A2(new_n7468_), .ZN(new_n8976_));
  AOI22_X1   g06251(.A1(new_n7601_), .A2(new_n8976_), .B1(new_n5130_), .B2(new_n7467_), .ZN(new_n8977_));
  NOR4_X1    g06252(.A1(new_n8977_), .A2(new_n7000_), .A3(new_n7248_), .A4(new_n7629_), .ZN(new_n8978_));
  NOR2_X1    g06253(.A1(new_n5130_), .A2(new_n2455_), .ZN(new_n8979_));
  AOI21_X1   g06254(.A1(new_n7601_), .A2(new_n8979_), .B(pi0040), .ZN(new_n8980_));
  AOI21_X1   g06255(.A1(new_n8978_), .A2(new_n8980_), .B(new_n8872_), .ZN(new_n8981_));
  NOR2_X1    g06256(.A1(new_n5141_), .A2(pi0179), .ZN(new_n8982_));
  INV_X1     g06257(.I(pi0179), .ZN(new_n8983_));
  NOR2_X1    g06258(.A1(new_n7602_), .A2(pi0040), .ZN(new_n8984_));
  OAI21_X1   g06259(.A1(new_n8984_), .A2(new_n6460_), .B(new_n8983_), .ZN(new_n8985_));
  AOI21_X1   g06260(.A1(new_n8981_), .A2(new_n8982_), .B(new_n8985_), .ZN(new_n8986_));
  INV_X1     g06261(.I(new_n8986_), .ZN(new_n8987_));
  AOI21_X1   g06262(.A1(new_n7154_), .A2(new_n7468_), .B(new_n8987_), .ZN(new_n8988_));
  NOR3_X1    g06263(.A1(new_n8986_), .A2(new_n7153_), .A3(new_n7468_), .ZN(new_n8989_));
  NOR4_X1    g06264(.A1(new_n8988_), .A2(pi0299), .A3(new_n8975_), .A4(new_n8989_), .ZN(new_n8990_));
  NOR3_X1    g06265(.A1(new_n8990_), .A2(new_n8974_), .A3(new_n5987_), .ZN(new_n8991_));
  NAND2_X1   g06266(.A1(new_n8974_), .A2(pi0232), .ZN(new_n8992_));
  NAND2_X1   g06267(.A1(new_n8984_), .A2(new_n5094_), .ZN(new_n8993_));
  NAND2_X1   g06268(.A1(new_n8980_), .A2(new_n6445_), .ZN(new_n8994_));
  AOI21_X1   g06269(.A1(new_n8993_), .A2(new_n8994_), .B(new_n7628_), .ZN(new_n8995_));
  NAND2_X1   g06270(.A1(new_n8984_), .A2(new_n5141_), .ZN(new_n8996_));
  AOI21_X1   g06271(.A1(new_n8980_), .A2(new_n6460_), .B(new_n7154_), .ZN(new_n8997_));
  OAI21_X1   g06272(.A1(new_n7153_), .A2(new_n7467_), .B(new_n2587_), .ZN(new_n8998_));
  AOI21_X1   g06273(.A1(new_n8996_), .A2(new_n8997_), .B(new_n8998_), .ZN(new_n8999_));
  NOR4_X1    g06274(.A1(new_n8995_), .A2(new_n8999_), .A3(new_n3154_), .A4(pi0232), .ZN(new_n9000_));
  OAI21_X1   g06275(.A1(new_n8990_), .A2(new_n8992_), .B(new_n9000_), .ZN(new_n9001_));
  NOR2_X1    g06276(.A1(new_n8991_), .A2(new_n9001_), .ZN(new_n9002_));
  NOR4_X1    g06277(.A1(new_n8973_), .A2(new_n5864_), .A3(new_n8972_), .A4(new_n9002_), .ZN(new_n9003_));
  OAI21_X1   g06278(.A1(new_n8918_), .A2(new_n8971_), .B(new_n9003_), .ZN(new_n9004_));
  NOR2_X1    g06279(.A1(new_n8861_), .A2(pi0147), .ZN(new_n9005_));
  OAI21_X1   g06280(.A1(new_n7280_), .A2(new_n7281_), .B(pi0187), .ZN(new_n9006_));
  INV_X1     g06281(.I(new_n9006_), .ZN(new_n9007_));
  AOI22_X1   g06282(.A1(new_n9007_), .A2(pi0147), .B1(new_n7283_), .B2(new_n9005_), .ZN(new_n9008_));
  NOR2_X1    g06283(.A1(new_n8860_), .A2(new_n3173_), .ZN(new_n9009_));
  INV_X1     g06284(.I(new_n9009_), .ZN(new_n9010_));
  INV_X1     g06285(.I(new_n8842_), .ZN(new_n9011_));
  NOR3_X1    g06286(.A1(new_n9011_), .A2(new_n3177_), .A3(new_n2455_), .ZN(new_n9012_));
  OAI21_X1   g06287(.A1(new_n8863_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n9013_));
  NOR4_X1    g06288(.A1(new_n9010_), .A2(pi0087), .A3(pi0100), .A4(new_n3209_), .ZN(new_n9015_));
  OAI21_X1   g06289(.A1(new_n9008_), .A2(new_n3172_), .B(new_n9015_), .ZN(new_n9016_));
  AOI21_X1   g06290(.A1(new_n9004_), .A2(new_n3172_), .B(new_n9016_), .ZN(new_n9017_));
  AOI21_X1   g06291(.A1(new_n7118_), .A2(new_n2455_), .B(pi0040), .ZN(new_n9018_));
  MUX2_X1    g06292(.I0(pi0179), .I1(pi0156), .S(pi0299), .Z(new_n9019_));
  NAND3_X1   g06293(.A1(new_n5988_), .A2(new_n2455_), .A3(new_n9019_), .ZN(new_n9020_));
  AOI21_X1   g06294(.A1(new_n9018_), .A2(new_n9020_), .B(pi0039), .ZN(new_n9021_));
  AOI21_X1   g06295(.A1(new_n7468_), .A2(pi0039), .B(new_n7739_), .ZN(new_n9022_));
  OAI21_X1   g06296(.A1(new_n9013_), .A2(new_n9012_), .B(new_n9022_), .ZN(new_n9023_));
  OAI21_X1   g06297(.A1(new_n9021_), .A2(new_n9023_), .B(new_n9010_), .ZN(new_n9024_));
  AOI22_X1   g06298(.A1(new_n9024_), .A2(new_n7123_), .B1(pi0075), .B2(new_n8859_), .ZN(new_n9025_));
  OAI21_X1   g06299(.A1(new_n9017_), .A2(new_n9025_), .B(new_n3214_), .ZN(new_n9026_));
  AOI21_X1   g06300(.A1(new_n9026_), .A2(new_n8865_), .B(pi0074), .ZN(new_n9027_));
  AOI21_X1   g06301(.A1(new_n7084_), .A2(new_n5109_), .B(new_n7087_), .ZN(new_n9028_));
  INV_X1     g06302(.I(new_n9028_), .ZN(new_n9029_));
  OR3_X2     g06303(.A1(new_n9018_), .A2(new_n8826_), .A3(new_n5987_), .Z(new_n9030_));
  OAI21_X1   g06304(.A1(new_n9030_), .A2(new_n9029_), .B(new_n3154_), .ZN(new_n9031_));
  OR2_X2     g06305(.A1(new_n8844_), .A2(new_n9012_), .Z(new_n9032_));
  AOI21_X1   g06306(.A1(new_n9031_), .A2(new_n9022_), .B(new_n9032_), .ZN(new_n9033_));
  NOR2_X1    g06307(.A1(pi0075), .A2(pi0092), .ZN(new_n9034_));
  OAI21_X1   g06308(.A1(new_n9033_), .A2(new_n8841_), .B(new_n9034_), .ZN(new_n9035_));
  NOR2_X1    g06309(.A1(new_n8835_), .A2(pi0074), .ZN(new_n9036_));
  OAI21_X1   g06310(.A1(new_n3214_), .A2(new_n8838_), .B(new_n9036_), .ZN(new_n9037_));
  AOI21_X1   g06311(.A1(new_n9035_), .A2(pi0054), .B(new_n9037_), .ZN(new_n9038_));
  NAND2_X1   g06312(.A1(new_n7048_), .A2(new_n3202_), .ZN(new_n9039_));
  OAI21_X1   g06313(.A1(new_n8859_), .A2(new_n9039_), .B(new_n3227_), .ZN(new_n9040_));
  OAI21_X1   g06314(.A1(new_n9038_), .A2(new_n5586_), .B(new_n9040_), .ZN(new_n9041_));
  OAI22_X1   g06315(.A1(new_n9027_), .A2(new_n9041_), .B1(new_n2533_), .B2(new_n7680_), .ZN(new_n9042_));
  AOI21_X1   g06316(.A1(new_n9042_), .A2(new_n8852_), .B(new_n8839_), .ZN(new_n9043_));
  NAND2_X1   g06317(.A1(new_n9008_), .A2(pi0038), .ZN(new_n9044_));
  NOR2_X1    g06318(.A1(new_n7228_), .A2(pi0210), .ZN(new_n9051_));
  INV_X1     g06319(.I(new_n7244_), .ZN(new_n9065_));
  NAND3_X1   g06320(.A1(new_n3364_), .A2(new_n5987_), .A3(pi0038), .ZN(new_n9106_));
  NAND2_X1   g06321(.A1(new_n9044_), .A2(new_n9106_), .ZN(new_n9107_));
  NOR2_X1    g06322(.A1(pi0087), .A2(pi0100), .ZN(new_n9109_));
  NAND2_X1   g06323(.A1(new_n2628_), .A2(new_n3203_), .ZN(new_n9113_));
  AOI21_X1   g06324(.A1(new_n9107_), .A2(new_n9109_), .B(new_n9113_), .ZN(new_n9114_));
  NAND2_X1   g06325(.A1(new_n8865_), .A2(new_n3214_), .ZN(new_n9115_));
  NOR2_X1    g06326(.A1(new_n9040_), .A2(pi0074), .ZN(new_n9116_));
  OAI21_X1   g06327(.A1(new_n9114_), .A2(new_n9115_), .B(new_n9116_), .ZN(new_n9117_));
  OR4_X2     g06328(.A1(new_n2628_), .A2(new_n8834_), .A3(pi0100), .A4(new_n8843_), .Z(new_n9120_));
  AOI21_X1   g06329(.A1(pi0054), .A2(new_n9120_), .B(new_n9037_), .ZN(new_n9121_));
  NOR3_X1    g06330(.A1(new_n8851_), .A2(new_n9121_), .A3(new_n5586_), .ZN(new_n9122_));
  AOI21_X1   g06331(.A1(new_n9117_), .A2(new_n9122_), .B(new_n8839_), .ZN(new_n9123_));
  NOR2_X1    g06332(.A1(new_n7317_), .A2(pi0079), .ZN(new_n9124_));
  NAND2_X1   g06333(.A1(new_n7751_), .A2(new_n7314_), .ZN(new_n9125_));
  NAND4_X1   g06334(.A1(new_n9043_), .A2(new_n9123_), .A3(new_n9124_), .A4(new_n9125_), .ZN(new_n9126_));
  OAI21_X1   g06335(.A1(new_n9123_), .A2(new_n7315_), .B(new_n9125_), .ZN(new_n9127_));
  AOI21_X1   g06336(.A1(new_n9043_), .A2(pi0079), .B(new_n9127_), .ZN(new_n9128_));
  NAND2_X1   g06337(.A1(new_n9126_), .A2(new_n9128_), .ZN(po0237));
  NOR2_X1    g06338(.A1(new_n8394_), .A2(new_n2923_), .ZN(new_n9130_));
  INV_X1     g06339(.I(new_n9130_), .ZN(new_n9131_));
  NOR2_X1    g06340(.A1(new_n9131_), .A2(new_n2924_), .ZN(new_n9132_));
  NOR2_X1    g06341(.A1(new_n2926_), .A2(pi0567), .ZN(new_n9133_));
  NOR2_X1    g06342(.A1(new_n9132_), .A2(new_n9133_), .ZN(new_n9134_));
  INV_X1     g06343(.I(new_n9134_), .ZN(new_n9135_));
  AOI21_X1   g06344(.A1(new_n9135_), .A2(pi0591), .B(new_n6203_), .ZN(new_n9136_));
  INV_X1     g06345(.I(new_n9136_), .ZN(new_n9137_));
  NOR2_X1    g06346(.A1(new_n9135_), .A2(new_n6084_), .ZN(new_n9138_));
  INV_X1     g06347(.I(new_n9138_), .ZN(new_n9139_));
  NOR2_X1    g06348(.A1(new_n9135_), .A2(new_n5941_), .ZN(new_n9140_));
  INV_X1     g06349(.I(new_n6003_), .ZN(new_n9141_));
  INV_X1     g06350(.I(new_n9132_), .ZN(new_n9142_));
  NOR2_X1    g06351(.A1(new_n9142_), .A2(new_n2918_), .ZN(new_n9143_));
  INV_X1     g06352(.I(new_n9143_), .ZN(new_n9144_));
  NAND3_X1   g06353(.A1(new_n7978_), .A2(new_n2710_), .A3(new_n2467_), .ZN(new_n9145_));
  NOR3_X1    g06354(.A1(new_n9145_), .A2(new_n6986_), .A3(new_n2678_), .ZN(new_n9146_));
  NAND2_X1   g06355(.A1(new_n5959_), .A2(new_n9146_), .ZN(new_n9147_));
  XOR2_X1    g06356(.A1(pi0090), .A2(pi0093), .Z(new_n9148_));
  NOR2_X1    g06357(.A1(new_n5239_), .A2(pi0841), .ZN(new_n9149_));
  AOI22_X1   g06358(.A1(pi0051), .A2(new_n5966_), .B1(new_n9149_), .B2(new_n9148_), .ZN(new_n9150_));
  NOR2_X1    g06359(.A1(new_n9147_), .A2(new_n9150_), .ZN(new_n9151_));
  NAND4_X1   g06360(.A1(new_n3418_), .A2(new_n2659_), .A3(pi0824), .A4(pi0950), .ZN(new_n9152_));
  OAI21_X1   g06361(.A1(new_n9151_), .A2(new_n9152_), .B(new_n8394_), .ZN(new_n9153_));
  NAND2_X1   g06362(.A1(new_n9153_), .A2(pi1092), .ZN(new_n9154_));
  OAI21_X1   g06363(.A1(new_n9154_), .A2(new_n9141_), .B(new_n9144_), .ZN(new_n9155_));
  NAND2_X1   g06364(.A1(new_n9155_), .A2(new_n2625_), .ZN(new_n9156_));
  NOR2_X1    g06365(.A1(new_n5366_), .A2(new_n2928_), .ZN(new_n9157_));
  NAND3_X1   g06366(.A1(new_n5966_), .A2(new_n2488_), .A3(new_n9157_), .ZN(new_n9158_));
  OAI21_X1   g06367(.A1(new_n9147_), .A2(new_n9158_), .B(new_n8394_), .ZN(new_n9159_));
  NAND3_X1   g06368(.A1(new_n9159_), .A2(pi1092), .A3(new_n6003_), .ZN(new_n9160_));
  AOI21_X1   g06369(.A1(new_n9160_), .A2(new_n9144_), .B(new_n6236_), .ZN(new_n9161_));
  INV_X1     g06370(.I(new_n9161_), .ZN(new_n9162_));
  NOR2_X1    g06371(.A1(new_n9132_), .A2(new_n3198_), .ZN(new_n9163_));
  INV_X1     g06372(.I(new_n9163_), .ZN(new_n9164_));
  NAND3_X1   g06373(.A1(new_n9156_), .A2(new_n9162_), .A3(new_n9164_), .ZN(new_n9165_));
  MUX2_X1    g06374(.I0(new_n9165_), .I1(new_n9132_), .S(new_n2628_), .Z(new_n9166_));
  NAND2_X1   g06375(.A1(new_n9166_), .A2(new_n6267_), .ZN(new_n9167_));
  NOR2_X1    g06376(.A1(new_n9133_), .A2(new_n5942_), .ZN(new_n9168_));
  AOI21_X1   g06377(.A1(new_n9167_), .A2(new_n9168_), .B(new_n9140_), .ZN(new_n9169_));
  NAND2_X1   g06378(.A1(new_n9169_), .A2(new_n6084_), .ZN(new_n9170_));
  NAND2_X1   g06379(.A1(new_n9170_), .A2(new_n9139_), .ZN(new_n9171_));
  NAND2_X1   g06380(.A1(new_n9171_), .A2(new_n6107_), .ZN(new_n9172_));
  INV_X1     g06381(.I(new_n6878_), .ZN(new_n9173_));
  AOI21_X1   g06382(.A1(new_n9171_), .A2(new_n9135_), .B(new_n9173_), .ZN(new_n9174_));
  INV_X1     g06383(.I(new_n9171_), .ZN(new_n9175_));
  NOR2_X1    g06384(.A1(new_n9134_), .A2(new_n6149_), .ZN(new_n9176_));
  AOI21_X1   g06385(.A1(new_n9175_), .A2(new_n6149_), .B(new_n9176_), .ZN(new_n9177_));
  NOR2_X1    g06386(.A1(new_n9177_), .A2(pi0355), .ZN(new_n9178_));
  MUX2_X1    g06387(.I0(new_n9171_), .I1(new_n9134_), .S(new_n6160_), .Z(new_n9179_));
  NOR2_X1    g06388(.A1(new_n9179_), .A2(new_n6130_), .ZN(new_n9180_));
  NOR2_X1    g06389(.A1(new_n9180_), .A2(new_n9178_), .ZN(new_n9181_));
  NAND3_X1   g06390(.A1(new_n9181_), .A2(new_n6131_), .A3(new_n6147_), .ZN(new_n9184_));
  AOI21_X1   g06391(.A1(new_n9134_), .A2(new_n6156_), .B(pi1196), .ZN(new_n9185_));
  AOI22_X1   g06392(.A1(new_n9184_), .A2(new_n9185_), .B1(pi1198), .B2(new_n9174_), .ZN(new_n9186_));
  OAI21_X1   g06393(.A1(new_n9186_), .A2(new_n6107_), .B(new_n9172_), .ZN(new_n9187_));
  MUX2_X1    g06394(.I0(new_n9187_), .I1(new_n9171_), .S(new_n6182_), .Z(new_n9188_));
  XOR2_X1    g06395(.A1(new_n9187_), .A2(new_n9171_), .Z(new_n9189_));
  NOR2_X1    g06396(.A1(new_n9189_), .A2(new_n6089_), .ZN(new_n9190_));
  XOR2_X1    g06397(.A1(new_n9190_), .A2(new_n9171_), .Z(new_n9191_));
  XOR2_X1    g06398(.A1(new_n9191_), .A2(new_n9188_), .Z(new_n9192_));
  NOR2_X1    g06399(.A1(new_n9192_), .A2(new_n6180_), .ZN(new_n9193_));
  XNOR2_X1   g06400(.A1(new_n9193_), .A2(new_n9188_), .ZN(new_n9194_));
  OR2_X2     g06401(.A1(new_n9194_), .A2(pi0356), .Z(new_n9195_));
  INV_X1     g06402(.I(new_n9192_), .ZN(new_n9196_));
  NOR2_X1    g06403(.A1(new_n9196_), .A2(new_n6180_), .ZN(new_n9197_));
  XNOR2_X1   g06404(.A1(new_n9197_), .A2(new_n9188_), .ZN(new_n9198_));
  OAI21_X1   g06405(.A1(new_n6198_), .A2(new_n9198_), .B(new_n9195_), .ZN(new_n9199_));
  OR2_X2     g06406(.A1(new_n9194_), .A2(new_n6198_), .Z(new_n9200_));
  OAI21_X1   g06407(.A1(pi0356), .A2(new_n9198_), .B(new_n9200_), .ZN(new_n9201_));
  XOR2_X1    g06408(.A1(new_n9199_), .A2(new_n9201_), .Z(new_n9202_));
  NAND2_X1   g06409(.A1(new_n9202_), .A2(pi0354), .ZN(new_n9203_));
  XNOR2_X1   g06410(.A1(new_n9203_), .A2(new_n9199_), .ZN(new_n9204_));
  XOR2_X1    g06411(.A1(new_n9203_), .A2(new_n9201_), .Z(new_n9205_));
  OAI21_X1   g06412(.A1(new_n9205_), .A2(new_n6196_), .B(new_n5940_), .ZN(new_n9206_));
  AOI21_X1   g06413(.A1(new_n6196_), .A2(new_n9204_), .B(new_n9206_), .ZN(new_n9207_));
  XOR2_X1    g06414(.A1(pi0370), .A2(pi0371), .Z(new_n9208_));
  INV_X1     g06415(.I(new_n9208_), .ZN(new_n9209_));
  NOR2_X1    g06416(.A1(new_n6699_), .A2(new_n6392_), .ZN(new_n9210_));
  AOI21_X1   g06417(.A1(new_n6699_), .A2(new_n9209_), .B(new_n9210_), .ZN(new_n9211_));
  INV_X1     g06418(.I(new_n9211_), .ZN(new_n9212_));
  NOR2_X1    g06419(.A1(new_n9135_), .A2(pi0592), .ZN(new_n9213_));
  AOI21_X1   g06420(.A1(new_n9169_), .A2(pi0592), .B(new_n9213_), .ZN(new_n9214_));
  NAND4_X1   g06421(.A1(new_n9214_), .A2(new_n6088_), .A3(new_n6909_), .A4(new_n9135_), .ZN(new_n9215_));
  XOR2_X1    g06422(.A1(new_n6323_), .A2(pi0367), .Z(new_n9216_));
  NAND2_X1   g06423(.A1(new_n6318_), .A2(new_n9216_), .ZN(new_n9217_));
  XOR2_X1    g06424(.A1(new_n6323_), .A2(pi0367), .Z(new_n9218_));
  OAI21_X1   g06425(.A1(new_n6318_), .A2(new_n9218_), .B(new_n9217_), .ZN(new_n9219_));
  OAI21_X1   g06426(.A1(new_n9219_), .A2(new_n9134_), .B(new_n6090_), .ZN(new_n9220_));
  AOI21_X1   g06427(.A1(new_n9214_), .A2(new_n9219_), .B(new_n9220_), .ZN(new_n9221_));
  INV_X1     g06428(.I(new_n6351_), .ZN(new_n9222_));
  OAI21_X1   g06429(.A1(new_n9214_), .A2(new_n9222_), .B(new_n6088_), .ZN(new_n9223_));
  AOI21_X1   g06430(.A1(new_n6090_), .A2(new_n9135_), .B(new_n6351_), .ZN(new_n9224_));
  NAND2_X1   g06431(.A1(new_n9223_), .A2(new_n9224_), .ZN(new_n9225_));
  OAI21_X1   g06432(.A1(new_n9225_), .A2(new_n9221_), .B(new_n9215_), .ZN(new_n9226_));
  MUX2_X1    g06433(.I0(new_n9226_), .I1(new_n9214_), .S(new_n6685_), .Z(new_n9227_));
  INV_X1     g06434(.I(pi0369), .ZN(new_n9228_));
  INV_X1     g06435(.I(new_n9214_), .ZN(new_n9229_));
  XOR2_X1    g06436(.A1(new_n9226_), .A2(new_n9229_), .Z(new_n9230_));
  NOR2_X1    g06437(.A1(new_n9230_), .A2(new_n6690_), .ZN(new_n9231_));
  XOR2_X1    g06438(.A1(new_n9231_), .A2(new_n9229_), .Z(new_n9232_));
  XOR2_X1    g06439(.A1(new_n9232_), .A2(new_n9227_), .Z(new_n9233_));
  NOR2_X1    g06440(.A1(new_n9233_), .A2(new_n9228_), .ZN(new_n9234_));
  XOR2_X1    g06441(.A1(new_n9234_), .A2(new_n9227_), .Z(new_n9235_));
  NOR2_X1    g06442(.A1(new_n9235_), .A2(new_n9212_), .ZN(new_n9236_));
  XNOR2_X1   g06443(.A1(new_n9234_), .A2(new_n9232_), .ZN(new_n9237_));
  OAI21_X1   g06444(.A1(new_n9237_), .A2(new_n9211_), .B(new_n5940_), .ZN(new_n9238_));
  OAI21_X1   g06445(.A1(new_n9238_), .A2(new_n9236_), .B(new_n6203_), .ZN(new_n9239_));
  INV_X1     g06446(.I(new_n6661_), .ZN(new_n9240_));
  INV_X1     g06447(.I(pi0392), .ZN(new_n9241_));
  NAND2_X1   g06448(.A1(new_n6260_), .A2(new_n9154_), .ZN(new_n9242_));
  OAI21_X1   g06449(.A1(new_n6260_), .A2(new_n9130_), .B(new_n9242_), .ZN(new_n9243_));
  NOR2_X1    g06450(.A1(new_n9243_), .A2(new_n9156_), .ZN(new_n9244_));
  NAND2_X1   g06451(.A1(new_n9159_), .A2(pi1092), .ZN(new_n9245_));
  NOR2_X1    g06452(.A1(new_n6260_), .A2(new_n9130_), .ZN(new_n9246_));
  AOI21_X1   g06453(.A1(new_n6260_), .A2(new_n9245_), .B(new_n9246_), .ZN(new_n9247_));
  AOI22_X1   g06454(.A1(new_n9247_), .A2(new_n9161_), .B1(new_n3198_), .B2(new_n9132_), .ZN(new_n9248_));
  OAI22_X1   g06455(.A1(new_n9248_), .A2(new_n9244_), .B1(new_n6582_), .B2(new_n9140_), .ZN(new_n9249_));
  OAI21_X1   g06456(.A1(new_n9135_), .A2(new_n5941_), .B(new_n6572_), .ZN(new_n9250_));
  MUX2_X1    g06457(.I0(new_n9131_), .I1(new_n9154_), .S(new_n6233_), .Z(new_n9251_));
  OAI21_X1   g06458(.A1(new_n9251_), .A2(new_n9141_), .B(new_n9144_), .ZN(new_n9252_));
  NAND2_X1   g06459(.A1(new_n9252_), .A2(new_n2625_), .ZN(new_n9253_));
  NOR4_X1    g06460(.A1(new_n9147_), .A2(pi0098), .A3(new_n2923_), .A4(new_n9158_), .ZN(new_n9254_));
  NAND2_X1   g06461(.A1(new_n6234_), .A2(new_n9254_), .ZN(new_n9255_));
  XOR2_X1    g06462(.A1(new_n9255_), .A2(new_n9245_), .Z(new_n9256_));
  NAND2_X1   g06463(.A1(new_n9256_), .A2(new_n6003_), .ZN(new_n9257_));
  NAND2_X1   g06464(.A1(new_n9257_), .A2(new_n9144_), .ZN(new_n9258_));
  NAND2_X1   g06465(.A1(new_n9258_), .A2(new_n6072_), .ZN(new_n9259_));
  NAND3_X1   g06466(.A1(new_n9259_), .A2(new_n9164_), .A3(new_n9253_), .ZN(new_n9260_));
  NOR4_X1    g06467(.A1(new_n9260_), .A2(new_n6256_), .A3(new_n9162_), .A4(new_n9244_), .ZN(new_n9261_));
  OAI21_X1   g06468(.A1(new_n9261_), .A2(new_n9250_), .B(new_n9249_), .ZN(new_n9262_));
  NAND2_X1   g06469(.A1(new_n9262_), .A2(new_n2628_), .ZN(new_n9263_));
  INV_X1     g06470(.I(new_n9168_), .ZN(new_n9264_));
  OAI21_X1   g06471(.A1(new_n6262_), .A2(new_n9264_), .B(new_n9135_), .ZN(new_n9265_));
  AOI21_X1   g06472(.A1(new_n9265_), .A2(pi1199), .B(pi0567), .ZN(new_n9266_));
  AND2_X2    g06473(.A1(new_n9260_), .A2(new_n2628_), .Z(new_n9267_));
  OAI21_X1   g06474(.A1(new_n9134_), .A2(new_n6572_), .B(new_n6088_), .ZN(new_n9268_));
  NAND2_X1   g06475(.A1(new_n9142_), .A2(pi0075), .ZN(new_n9269_));
  NOR2_X1    g06476(.A1(new_n9168_), .A2(new_n6267_), .ZN(new_n9270_));
  NAND4_X1   g06477(.A1(new_n9250_), .A2(new_n9268_), .A3(new_n9269_), .A4(new_n9270_), .ZN(new_n9271_));
  OAI21_X1   g06478(.A1(new_n9267_), .A2(new_n9271_), .B(new_n6539_), .ZN(new_n9272_));
  AOI21_X1   g06479(.A1(new_n9263_), .A2(new_n9266_), .B(new_n9272_), .ZN(new_n9273_));
  NOR2_X1    g06480(.A1(new_n6279_), .A2(pi1197), .ZN(new_n9274_));
  NOR2_X1    g06481(.A1(new_n9171_), .A2(new_n9274_), .ZN(new_n9275_));
  AOI21_X1   g06482(.A1(new_n9273_), .A2(pi1197), .B(new_n9275_), .ZN(new_n9276_));
  NAND2_X1   g06483(.A1(new_n9175_), .A2(new_n6279_), .ZN(new_n9277_));
  AND2_X2    g06484(.A1(new_n9273_), .A2(new_n9277_), .Z(new_n9278_));
  XOR2_X1    g06485(.A1(new_n9278_), .A2(new_n9276_), .Z(new_n9279_));
  XNOR2_X1   g06486(.A1(pi0333), .A2(pi0391), .ZN(new_n9280_));
  INV_X1     g06487(.I(new_n9280_), .ZN(new_n9281_));
  NAND2_X1   g06488(.A1(new_n9279_), .A2(new_n9281_), .ZN(new_n9282_));
  XOR2_X1    g06489(.A1(new_n9282_), .A2(new_n9276_), .Z(new_n9283_));
  NAND2_X1   g06490(.A1(new_n9283_), .A2(new_n9241_), .ZN(new_n9284_));
  NOR2_X1    g06491(.A1(new_n9279_), .A2(new_n9280_), .ZN(new_n9285_));
  XOR2_X1    g06492(.A1(new_n9285_), .A2(new_n9276_), .Z(new_n9286_));
  OAI21_X1   g06493(.A1(new_n9241_), .A2(new_n9286_), .B(new_n9284_), .ZN(new_n9287_));
  XNOR2_X1   g06494(.A1(pi0333), .A2(pi0391), .ZN(new_n9288_));
  NOR2_X1    g06495(.A1(new_n9288_), .A2(new_n6205_), .ZN(new_n9289_));
  XOR2_X1    g06496(.A1(new_n9287_), .A2(new_n9289_), .Z(new_n9290_));
  NAND2_X1   g06497(.A1(new_n9290_), .A2(new_n9240_), .ZN(new_n9291_));
  NAND2_X1   g06498(.A1(new_n9283_), .A2(pi0392), .ZN(new_n9292_));
  OAI21_X1   g06499(.A1(pi0392), .A2(new_n9286_), .B(new_n9292_), .ZN(new_n9293_));
  XOR2_X1    g06500(.A1(new_n9293_), .A2(new_n9289_), .Z(new_n9294_));
  NAND2_X1   g06501(.A1(new_n9294_), .A2(new_n6661_), .ZN(new_n9295_));
  AOI21_X1   g06502(.A1(new_n9291_), .A2(new_n9295_), .B(pi0591), .ZN(new_n9296_));
  AOI21_X1   g06503(.A1(new_n9296_), .A2(new_n9239_), .B(pi0588), .ZN(new_n9297_));
  OAI21_X1   g06504(.A1(new_n9207_), .A2(new_n9137_), .B(new_n9297_), .ZN(new_n9298_));
  AOI21_X1   g06505(.A1(new_n9134_), .A2(new_n6798_), .B(new_n6711_), .ZN(new_n9299_));
  NOR2_X1    g06506(.A1(new_n9134_), .A2(pi1196), .ZN(new_n9300_));
  INV_X1     g06507(.I(pi0429), .ZN(new_n9301_));
  INV_X1     g06508(.I(pi0435), .ZN(new_n9302_));
  INV_X1     g06509(.I(new_n6756_), .ZN(new_n9303_));
  NOR2_X1    g06510(.A1(new_n9135_), .A2(pi0443), .ZN(new_n9304_));
  AOI21_X1   g06511(.A1(new_n9171_), .A2(pi0443), .B(new_n9304_), .ZN(new_n9305_));
  NOR2_X1    g06512(.A1(new_n9135_), .A2(new_n6745_), .ZN(new_n9306_));
  AOI21_X1   g06513(.A1(new_n9171_), .A2(new_n6745_), .B(new_n9306_), .ZN(new_n9307_));
  INV_X1     g06514(.I(new_n9307_), .ZN(new_n9308_));
  NOR2_X1    g06515(.A1(new_n9308_), .A2(new_n9303_), .ZN(new_n9309_));
  AOI21_X1   g06516(.A1(new_n9303_), .A2(new_n9305_), .B(new_n9309_), .ZN(new_n9310_));
  NOR2_X1    g06517(.A1(new_n9310_), .A2(new_n9302_), .ZN(new_n9311_));
  XNOR2_X1   g06518(.A1(pi0436), .A2(pi0444), .ZN(new_n9312_));
  MUX2_X1    g06519(.I0(new_n9308_), .I1(new_n9305_), .S(new_n9312_), .Z(new_n9313_));
  AOI21_X1   g06520(.A1(new_n9302_), .A2(new_n9313_), .B(new_n9311_), .ZN(new_n9314_));
  NAND2_X1   g06521(.A1(new_n9313_), .A2(pi0435), .ZN(new_n9315_));
  OAI21_X1   g06522(.A1(pi0435), .A2(new_n9310_), .B(new_n9315_), .ZN(new_n9316_));
  INV_X1     g06523(.I(new_n9316_), .ZN(new_n9317_));
  AOI21_X1   g06524(.A1(new_n9317_), .A2(new_n9301_), .B(new_n9314_), .ZN(new_n9318_));
  NAND3_X1   g06525(.A1(new_n9314_), .A2(new_n9301_), .A3(new_n9316_), .ZN(new_n9319_));
  NAND4_X1   g06526(.A1(new_n9317_), .A2(new_n9314_), .A3(pi0429), .A4(new_n6751_), .ZN(new_n9320_));
  NOR3_X1    g06527(.A1(new_n6750_), .A2(new_n6209_), .A3(new_n6749_), .ZN(new_n9321_));
  NAND3_X1   g06528(.A1(new_n9320_), .A2(new_n9319_), .A3(new_n9321_), .ZN(new_n9322_));
  NOR2_X1    g06529(.A1(new_n9322_), .A2(new_n9318_), .ZN(new_n9323_));
  NOR2_X1    g06530(.A1(new_n9323_), .A2(new_n9300_), .ZN(new_n9324_));
  MUX2_X1    g06531(.I0(new_n9171_), .I1(new_n9324_), .S(new_n6743_), .Z(new_n9325_));
  MUX2_X1    g06532(.I0(new_n9325_), .I1(new_n9175_), .S(new_n6824_), .Z(new_n9326_));
  MUX2_X1    g06533(.I0(new_n9325_), .I1(new_n9175_), .S(new_n6766_), .Z(new_n9327_));
  XOR2_X1    g06534(.A1(new_n9327_), .A2(new_n9326_), .Z(new_n9328_));
  NOR2_X1    g06535(.A1(new_n9328_), .A2(new_n6712_), .ZN(new_n9329_));
  XNOR2_X1   g06536(.A1(new_n9329_), .A2(new_n9326_), .ZN(new_n9330_));
  NAND2_X1   g06537(.A1(new_n9328_), .A2(new_n6773_), .ZN(new_n9331_));
  XOR2_X1    g06538(.A1(new_n9331_), .A2(new_n9326_), .Z(new_n9332_));
  OR2_X2     g06539(.A1(new_n9332_), .A2(new_n6772_), .Z(new_n9333_));
  OAI21_X1   g06540(.A1(pi0445), .A2(new_n9330_), .B(new_n9333_), .ZN(new_n9334_));
  NOR3_X1    g06541(.A1(new_n9334_), .A2(pi0448), .A3(new_n6791_), .ZN(new_n9337_));
  OAI21_X1   g06542(.A1(new_n9325_), .A2(new_n6798_), .B(new_n6088_), .ZN(new_n9338_));
  OAI21_X1   g06543(.A1(new_n9337_), .A2(new_n9338_), .B(new_n9299_), .ZN(new_n9339_));
  NAND3_X1   g06544(.A1(new_n9298_), .A2(new_n6538_), .A3(new_n9339_), .ZN(new_n9340_));
  NOR2_X1    g06545(.A1(new_n9143_), .A2(new_n3198_), .ZN(new_n9341_));
  INV_X1     g06546(.I(new_n9341_), .ZN(new_n9342_));
  NAND4_X1   g06547(.A1(new_n9154_), .A2(pi0087), .A3(new_n9245_), .A4(new_n9342_), .ZN(new_n9343_));
  NOR2_X1    g06548(.A1(new_n6428_), .A2(new_n9132_), .ZN(new_n9344_));
  AOI21_X1   g06549(.A1(new_n9344_), .A2(new_n6029_), .B(new_n9141_), .ZN(new_n9345_));
  OAI21_X1   g06550(.A1(new_n9345_), .A2(new_n9342_), .B(new_n2628_), .ZN(new_n9346_));
  AOI21_X1   g06551(.A1(new_n9343_), .A2(pi0122), .B(new_n9346_), .ZN(new_n9347_));
  OAI22_X1   g06552(.A1(new_n9344_), .A2(new_n5941_), .B1(pi0567), .B2(new_n2926_), .ZN(new_n9348_));
  NOR2_X1    g06553(.A1(new_n5942_), .A2(new_n6267_), .ZN(new_n9349_));
  NAND2_X1   g06554(.A1(new_n9344_), .A2(new_n5980_), .ZN(new_n9350_));
  NAND3_X1   g06555(.A1(new_n9348_), .A2(new_n9350_), .A3(new_n9349_), .ZN(new_n9351_));
  NOR2_X1    g06556(.A1(new_n9347_), .A2(new_n9351_), .ZN(new_n9352_));
  AOI21_X1   g06557(.A1(new_n9352_), .A2(new_n6084_), .B(new_n9138_), .ZN(new_n9353_));
  INV_X1     g06558(.I(new_n9353_), .ZN(new_n9354_));
  AOI21_X1   g06559(.A1(new_n9135_), .A2(new_n9354_), .B(new_n9173_), .ZN(new_n9355_));
  AOI21_X1   g06560(.A1(new_n9353_), .A2(new_n6149_), .B(new_n9176_), .ZN(new_n9356_));
  NOR2_X1    g06561(.A1(new_n9356_), .A2(pi0355), .ZN(new_n9357_));
  MUX2_X1    g06562(.I0(new_n9353_), .I1(new_n9135_), .S(new_n6160_), .Z(new_n9358_));
  INV_X1     g06563(.I(new_n9358_), .ZN(new_n9359_));
  NOR2_X1    g06564(.A1(new_n9359_), .A2(new_n6130_), .ZN(new_n9360_));
  NOR2_X1    g06565(.A1(new_n9356_), .A2(new_n6130_), .ZN(new_n9361_));
  NOR2_X1    g06566(.A1(new_n9359_), .A2(pi0355), .ZN(new_n9362_));
  NOR2_X1    g06567(.A1(new_n9362_), .A2(new_n9361_), .ZN(new_n9363_));
  INV_X1     g06568(.I(new_n9363_), .ZN(new_n9364_));
  OAI22_X1   g06569(.A1(new_n9364_), .A2(pi0458), .B1(new_n9357_), .B2(new_n9360_), .ZN(new_n9365_));
  NOR2_X1    g06570(.A1(new_n9360_), .A2(new_n9357_), .ZN(new_n9366_));
  NAND3_X1   g06571(.A1(new_n9364_), .A2(new_n6131_), .A3(new_n9366_), .ZN(new_n9367_));
  NAND4_X1   g06572(.A1(new_n9366_), .A2(new_n9363_), .A3(pi0458), .A4(new_n6147_), .ZN(new_n9368_));
  NAND4_X1   g06573(.A1(new_n9365_), .A2(new_n6147_), .A3(new_n9367_), .A4(new_n9368_), .ZN(new_n9369_));
  AOI22_X1   g06574(.A1(new_n9369_), .A2(new_n9185_), .B1(pi1198), .B2(new_n9355_), .ZN(new_n9370_));
  NOR2_X1    g06575(.A1(new_n9370_), .A2(new_n6107_), .ZN(new_n9371_));
  AOI21_X1   g06576(.A1(new_n6107_), .A2(new_n9354_), .B(new_n9371_), .ZN(new_n9372_));
  XOR2_X1    g06577(.A1(new_n9372_), .A2(new_n9353_), .Z(new_n9373_));
  NAND2_X1   g06578(.A1(new_n9373_), .A2(new_n6182_), .ZN(new_n9374_));
  XOR2_X1    g06579(.A1(new_n9374_), .A2(new_n9372_), .Z(new_n9375_));
  MUX2_X1    g06580(.I0(new_n9372_), .I1(new_n9354_), .S(new_n6089_), .Z(new_n9376_));
  XOR2_X1    g06581(.A1(new_n9375_), .A2(new_n9376_), .Z(new_n9377_));
  NOR2_X1    g06582(.A1(new_n9377_), .A2(new_n6180_), .ZN(new_n9378_));
  XNOR2_X1   g06583(.A1(new_n9378_), .A2(new_n9375_), .ZN(new_n9379_));
  OR2_X2     g06584(.A1(new_n9379_), .A2(pi0356), .Z(new_n9380_));
  INV_X1     g06585(.I(new_n9377_), .ZN(new_n9381_));
  NOR2_X1    g06586(.A1(new_n9381_), .A2(new_n6180_), .ZN(new_n9382_));
  XNOR2_X1   g06587(.A1(new_n9382_), .A2(new_n9375_), .ZN(new_n9383_));
  OAI21_X1   g06588(.A1(new_n6198_), .A2(new_n9383_), .B(new_n9380_), .ZN(new_n9384_));
  OR2_X2     g06589(.A1(new_n9379_), .A2(new_n6198_), .Z(new_n9385_));
  OAI21_X1   g06590(.A1(pi0356), .A2(new_n9383_), .B(new_n9385_), .ZN(new_n9386_));
  XOR2_X1    g06591(.A1(new_n9384_), .A2(new_n9386_), .Z(new_n9387_));
  NAND2_X1   g06592(.A1(new_n9387_), .A2(pi0354), .ZN(new_n9388_));
  XNOR2_X1   g06593(.A1(new_n9388_), .A2(new_n9384_), .ZN(new_n9389_));
  XOR2_X1    g06594(.A1(new_n9388_), .A2(new_n9386_), .Z(new_n9390_));
  OAI21_X1   g06595(.A1(new_n9390_), .A2(new_n6196_), .B(new_n5940_), .ZN(new_n9391_));
  AOI21_X1   g06596(.A1(new_n6196_), .A2(new_n9389_), .B(new_n9391_), .ZN(new_n9392_));
  INV_X1     g06597(.I(pi0404), .ZN(new_n9393_));
  NOR2_X1    g06598(.A1(new_n9393_), .A2(pi0411), .ZN(new_n9394_));
  NOR2_X1    g06599(.A1(new_n6210_), .A2(pi0404), .ZN(new_n9395_));
  OAI21_X1   g06600(.A1(new_n9394_), .A2(new_n9395_), .B(new_n6211_), .ZN(new_n9396_));
  NOR2_X1    g06601(.A1(pi0404), .A2(pi0411), .ZN(new_n9397_));
  NOR2_X1    g06602(.A1(new_n9393_), .A2(new_n6210_), .ZN(new_n9398_));
  OAI21_X1   g06603(.A1(new_n9398_), .A2(new_n9397_), .B(pi0397), .ZN(new_n9399_));
  NAND2_X1   g06604(.A1(new_n9399_), .A2(new_n9396_), .ZN(new_n9400_));
  NAND2_X1   g06605(.A1(new_n9400_), .A2(new_n6226_), .ZN(new_n9401_));
  OAI21_X1   g06606(.A1(new_n6228_), .A2(new_n9400_), .B(new_n9401_), .ZN(new_n9402_));
  AOI21_X1   g06607(.A1(new_n9402_), .A2(new_n6004_), .B(new_n9130_), .ZN(new_n9403_));
  NOR2_X1    g06608(.A1(new_n9403_), .A2(pi0412), .ZN(new_n9404_));
  INV_X1     g06609(.I(pi0412), .ZN(new_n9405_));
  OR2_X2     g06610(.A1(new_n9402_), .A2(new_n6005_), .Z(new_n9406_));
  AOI21_X1   g06611(.A1(new_n9406_), .A2(new_n9131_), .B(new_n9405_), .ZN(new_n9407_));
  NOR3_X1    g06612(.A1(new_n9407_), .A2(new_n6221_), .A3(new_n9404_), .ZN(new_n9408_));
  AOI21_X1   g06613(.A1(pi0412), .A2(new_n9403_), .B(new_n9407_), .ZN(new_n9409_));
  AOI21_X1   g06614(.A1(new_n6217_), .A2(new_n6220_), .B(new_n9409_), .ZN(new_n9410_));
  NOR3_X1    g06615(.A1(new_n9410_), .A2(new_n9408_), .A3(pi0122), .ZN(new_n9411_));
  INV_X1     g06616(.I(new_n9411_), .ZN(new_n9412_));
  AOI21_X1   g06617(.A1(new_n9412_), .A2(new_n9131_), .B(new_n9141_), .ZN(new_n9413_));
  NOR2_X1    g06618(.A1(new_n9413_), .A2(new_n9143_), .ZN(new_n9414_));
  INV_X1     g06619(.I(new_n9414_), .ZN(new_n9415_));
  OAI21_X1   g06620(.A1(new_n9251_), .A2(new_n6029_), .B(new_n9412_), .ZN(new_n9416_));
  AOI21_X1   g06621(.A1(new_n9416_), .A2(new_n6003_), .B(pi0087), .ZN(new_n9417_));
  NOR2_X1    g06622(.A1(new_n9342_), .A2(new_n3177_), .ZN(new_n9418_));
  INV_X1     g06623(.I(new_n9418_), .ZN(new_n9419_));
  NAND2_X1   g06624(.A1(new_n9256_), .A2(pi0122), .ZN(new_n9420_));
  NAND2_X1   g06625(.A1(new_n9420_), .A2(new_n9412_), .ZN(new_n9421_));
  AOI21_X1   g06626(.A1(new_n9421_), .A2(new_n6003_), .B(new_n9419_), .ZN(new_n9422_));
  NOR2_X1    g06627(.A1(new_n9415_), .A2(new_n3197_), .ZN(new_n9423_));
  NOR4_X1    g06628(.A1(new_n9422_), .A2(new_n9341_), .A3(new_n9417_), .A4(new_n9423_), .ZN(new_n9424_));
  MUX2_X1    g06629(.I0(new_n9424_), .I1(new_n9415_), .S(pi0075), .Z(new_n9425_));
  NOR2_X1    g06630(.A1(new_n2925_), .A2(pi0567), .ZN(new_n9426_));
  AOI21_X1   g06631(.A1(new_n9414_), .A2(pi0567), .B(new_n9426_), .ZN(new_n9427_));
  INV_X1     g06632(.I(new_n9427_), .ZN(new_n9428_));
  OAI21_X1   g06633(.A1(new_n9428_), .A2(new_n9168_), .B(new_n6573_), .ZN(new_n9429_));
  AOI21_X1   g06634(.A1(new_n9425_), .A2(new_n9349_), .B(new_n9429_), .ZN(new_n9430_));
  NOR2_X1    g06635(.A1(new_n6005_), .A2(pi0122), .ZN(new_n9431_));
  INV_X1     g06636(.I(new_n9431_), .ZN(new_n9432_));
  NAND4_X1   g06637(.A1(new_n9131_), .A2(new_n6029_), .A3(new_n2918_), .A4(pi1093), .ZN(new_n9442_));
  AOI21_X1   g06638(.A1(new_n6260_), .A2(new_n6004_), .B(new_n9442_), .ZN(new_n9443_));
  OAI21_X1   g06639(.A1(new_n9130_), .A2(new_n9431_), .B(new_n9443_), .ZN(new_n9447_));
  AOI21_X1   g06640(.A1(new_n9447_), .A2(pi0567), .B(new_n9426_), .ZN(new_n9448_));
  INV_X1     g06641(.I(new_n9448_), .ZN(new_n9449_));
  OAI21_X1   g06642(.A1(new_n6267_), .A2(new_n9414_), .B(new_n9449_), .ZN(new_n9450_));
  AOI21_X1   g06643(.A1(new_n9135_), .A2(pi0592), .B(pi1199), .ZN(new_n9462_));
  OAI21_X1   g06644(.A1(new_n9430_), .A2(new_n9300_), .B(new_n9462_), .ZN(new_n9463_));
  MUX2_X1    g06645(.I0(new_n9463_), .I1(new_n9354_), .S(new_n9274_), .Z(new_n9464_));
  NOR2_X1    g06646(.A1(new_n9464_), .A2(new_n9281_), .ZN(new_n9465_));
  NOR2_X1    g06647(.A1(new_n9463_), .A2(new_n6279_), .ZN(new_n9466_));
  AOI21_X1   g06648(.A1(new_n6279_), .A2(new_n9354_), .B(new_n9466_), .ZN(new_n9467_));
  NOR2_X1    g06649(.A1(new_n9467_), .A2(new_n9280_), .ZN(new_n9468_));
  XOR2_X1    g06650(.A1(new_n9468_), .A2(new_n9465_), .Z(new_n9469_));
  XNOR2_X1   g06651(.A1(pi0392), .A2(pi0393), .ZN(new_n9470_));
  NAND2_X1   g06652(.A1(new_n9469_), .A2(new_n9470_), .ZN(new_n9471_));
  MUX2_X1    g06653(.I0(new_n9467_), .I1(new_n9464_), .S(new_n9281_), .Z(new_n9472_));
  OR2_X2     g06654(.A1(new_n9472_), .A2(new_n9470_), .Z(new_n9473_));
  OAI21_X1   g06655(.A1(new_n9471_), .A2(new_n9473_), .B(new_n9240_), .ZN(new_n9474_));
  AOI21_X1   g06656(.A1(new_n9471_), .A2(new_n9473_), .B(new_n9474_), .ZN(new_n9475_));
  NAND2_X1   g06657(.A1(new_n9472_), .A2(new_n9470_), .ZN(new_n9476_));
  NOR2_X1    g06658(.A1(new_n9469_), .A2(new_n9470_), .ZN(new_n9477_));
  XNOR2_X1   g06659(.A1(new_n9477_), .A2(new_n9476_), .ZN(new_n9478_));
  NOR2_X1    g06660(.A1(new_n9478_), .A2(new_n6661_), .ZN(new_n9479_));
  OAI21_X1   g06661(.A1(new_n9479_), .A2(new_n9475_), .B(pi0591), .ZN(new_n9480_));
  NOR2_X1    g06662(.A1(new_n6910_), .A2(new_n9134_), .ZN(new_n9481_));
  AOI21_X1   g06663(.A1(new_n9352_), .A2(pi0592), .B(new_n9213_), .ZN(new_n9482_));
  INV_X1     g06664(.I(new_n9482_), .ZN(new_n9483_));
  NOR2_X1    g06665(.A1(new_n6909_), .A2(new_n9483_), .ZN(new_n9484_));
  OAI21_X1   g06666(.A1(new_n9481_), .A2(new_n9484_), .B(pi1199), .ZN(new_n9485_));
  INV_X1     g06667(.I(new_n9218_), .ZN(new_n9486_));
  MUX2_X1    g06668(.I0(new_n9482_), .I1(new_n9135_), .S(new_n9486_), .Z(new_n9487_));
  NOR2_X1    g06669(.A1(new_n9486_), .A2(new_n6313_), .ZN(new_n9489_));
  INV_X1     g06670(.I(new_n9489_), .ZN(new_n9490_));
  XOR2_X1    g06671(.A1(new_n9487_), .A2(new_n9490_), .Z(new_n9491_));
  NOR2_X1    g06672(.A1(new_n9491_), .A2(new_n6317_), .ZN(new_n9492_));
  NAND3_X1   g06673(.A1(new_n9483_), .A2(new_n6312_), .A3(new_n9218_), .ZN(new_n9493_));
  MUX2_X1    g06674(.I0(new_n9482_), .I1(new_n9134_), .S(new_n9486_), .Z(new_n9494_));
  NAND2_X1   g06675(.A1(new_n9494_), .A2(new_n9490_), .ZN(new_n9495_));
  NAND3_X1   g06676(.A1(new_n9495_), .A2(new_n6317_), .A3(new_n9493_), .ZN(new_n9496_));
  NOR2_X1    g06677(.A1(new_n9224_), .A2(pi1197), .ZN(new_n9497_));
  OAI21_X1   g06678(.A1(new_n9492_), .A2(new_n9496_), .B(new_n9497_), .ZN(new_n9498_));
  AOI21_X1   g06679(.A1(new_n9483_), .A2(new_n6351_), .B(pi1199), .ZN(new_n9499_));
  NAND3_X1   g06680(.A1(new_n9498_), .A2(new_n9485_), .A3(new_n9499_), .ZN(new_n9500_));
  MUX2_X1    g06681(.I0(new_n9485_), .I1(new_n9483_), .S(pi1198), .Z(new_n9501_));
  AOI21_X1   g06682(.A1(new_n9498_), .A2(new_n9499_), .B(pi1198), .ZN(new_n9502_));
  NOR2_X1    g06683(.A1(new_n9501_), .A2(new_n9502_), .ZN(new_n9503_));
  NAND2_X1   g06684(.A1(new_n9503_), .A2(pi0374), .ZN(new_n9504_));
  OAI21_X1   g06685(.A1(pi0374), .A2(new_n9500_), .B(new_n9504_), .ZN(new_n9505_));
  NOR2_X1    g06686(.A1(new_n9500_), .A2(new_n6689_), .ZN(new_n9506_));
  AOI21_X1   g06687(.A1(new_n9503_), .A2(new_n6689_), .B(new_n9506_), .ZN(new_n9507_));
  XOR2_X1    g06688(.A1(new_n9505_), .A2(new_n9507_), .Z(new_n9508_));
  NOR2_X1    g06689(.A1(new_n9508_), .A2(new_n9228_), .ZN(new_n9509_));
  XOR2_X1    g06690(.A1(new_n9509_), .A2(new_n9505_), .Z(new_n9510_));
  NAND2_X1   g06691(.A1(new_n9510_), .A2(new_n9211_), .ZN(new_n9511_));
  XNOR2_X1   g06692(.A1(new_n9509_), .A2(new_n9507_), .ZN(new_n9512_));
  AOI21_X1   g06693(.A1(new_n9512_), .A2(new_n9212_), .B(pi0591), .ZN(new_n9513_));
  AOI21_X1   g06694(.A1(new_n9513_), .A2(new_n9511_), .B(pi0590), .ZN(new_n9514_));
  AOI21_X1   g06695(.A1(new_n9480_), .A2(new_n9514_), .B(pi0588), .ZN(new_n9515_));
  OAI21_X1   g06696(.A1(new_n9392_), .A2(new_n9137_), .B(new_n9515_), .ZN(new_n9516_));
  NOR2_X1    g06697(.A1(new_n9354_), .A2(new_n6824_), .ZN(new_n9517_));
  AOI21_X1   g06698(.A1(new_n9354_), .A2(pi0443), .B(new_n9304_), .ZN(new_n9518_));
  NAND2_X1   g06699(.A1(new_n9518_), .A2(new_n9303_), .ZN(new_n9519_));
  INV_X1     g06700(.I(new_n9306_), .ZN(new_n9520_));
  OAI21_X1   g06701(.A1(new_n9353_), .A2(pi0443), .B(new_n9520_), .ZN(new_n9521_));
  OAI21_X1   g06702(.A1(new_n9303_), .A2(new_n9521_), .B(new_n9519_), .ZN(new_n9522_));
  MUX2_X1    g06703(.I0(new_n9521_), .I1(new_n9518_), .S(new_n9312_), .Z(new_n9523_));
  AND2_X2    g06704(.A1(new_n9523_), .A2(new_n9302_), .Z(new_n9524_));
  AOI21_X1   g06705(.A1(pi0435), .A2(new_n9522_), .B(new_n9524_), .ZN(new_n9525_));
  NAND2_X1   g06706(.A1(new_n9522_), .A2(new_n9302_), .ZN(new_n9526_));
  NAND2_X1   g06707(.A1(new_n9523_), .A2(pi0435), .ZN(new_n9527_));
  NAND2_X1   g06708(.A1(new_n9526_), .A2(new_n9527_), .ZN(new_n9528_));
  INV_X1     g06709(.I(new_n9528_), .ZN(new_n9529_));
  AOI21_X1   g06710(.A1(new_n9301_), .A2(new_n9529_), .B(new_n9525_), .ZN(new_n9530_));
  NAND3_X1   g06711(.A1(new_n9525_), .A2(new_n9301_), .A3(new_n9528_), .ZN(new_n9531_));
  NAND4_X1   g06712(.A1(new_n9525_), .A2(new_n9529_), .A3(pi0429), .A4(new_n6751_), .ZN(new_n9532_));
  NAND3_X1   g06713(.A1(new_n9532_), .A2(new_n9531_), .A3(new_n9321_), .ZN(new_n9533_));
  OAI22_X1   g06714(.A1(new_n9533_), .A2(new_n9530_), .B1(pi1196), .B2(new_n9134_), .ZN(new_n9534_));
  MUX2_X1    g06715(.I0(new_n9353_), .I1(new_n9534_), .S(new_n6743_), .Z(new_n9535_));
  NOR2_X1    g06716(.A1(new_n9535_), .A2(new_n6766_), .ZN(new_n9536_));
  XOR2_X1    g06717(.A1(new_n9536_), .A2(new_n9517_), .Z(new_n9537_));
  MUX2_X1    g06718(.I0(new_n9535_), .I1(new_n9354_), .S(new_n6824_), .Z(new_n9538_));
  XNOR2_X1   g06719(.A1(new_n9537_), .A2(new_n9538_), .ZN(new_n9539_));
  NAND2_X1   g06720(.A1(new_n9539_), .A2(new_n6773_), .ZN(new_n9540_));
  XNOR2_X1   g06721(.A1(new_n9540_), .A2(new_n9537_), .ZN(new_n9541_));
  NOR2_X1    g06722(.A1(new_n9541_), .A2(pi0445), .ZN(new_n9542_));
  MUX2_X1    g06723(.I0(new_n9538_), .I1(new_n9537_), .S(new_n6712_), .Z(new_n9543_));
  NOR2_X1    g06724(.A1(new_n9543_), .A2(new_n6772_), .ZN(new_n9544_));
  NOR2_X1    g06725(.A1(new_n9542_), .A2(new_n9544_), .ZN(new_n9545_));
  XNOR2_X1   g06726(.A1(pi0426), .A2(pi0430), .ZN(new_n9546_));
  NOR2_X1    g06727(.A1(new_n9546_), .A2(pi0448), .ZN(new_n9547_));
  NOR2_X1    g06728(.A1(new_n9545_), .A2(new_n9547_), .ZN(new_n9548_));
  NAND2_X1   g06729(.A1(new_n9545_), .A2(new_n9547_), .ZN(new_n9549_));
  NOR2_X1    g06730(.A1(new_n9543_), .A2(pi0445), .ZN(new_n9550_));
  NOR2_X1    g06731(.A1(new_n9541_), .A2(new_n6772_), .ZN(new_n9551_));
  NOR2_X1    g06732(.A1(new_n9551_), .A2(new_n9550_), .ZN(new_n9552_));
  NAND4_X1   g06733(.A1(new_n9545_), .A2(new_n9552_), .A3(pi0448), .A4(new_n6924_), .ZN(new_n9553_));
  NAND3_X1   g06734(.A1(new_n9553_), .A2(new_n6924_), .A3(new_n9549_), .ZN(new_n9554_));
  AOI21_X1   g06735(.A1(new_n9535_), .A2(new_n6797_), .B(pi1199), .ZN(new_n9555_));
  OAI21_X1   g06736(.A1(new_n9554_), .A2(new_n9548_), .B(new_n9555_), .ZN(new_n9556_));
  AOI21_X1   g06737(.A1(new_n9556_), .A2(new_n9299_), .B(new_n6538_), .ZN(new_n9557_));
  XOR2_X1    g06738(.A1(new_n6662_), .A2(new_n9241_), .Z(new_n9558_));
  NOR2_X1    g06739(.A1(new_n6879_), .A2(new_n9135_), .ZN(new_n9559_));
  INV_X1     g06740(.I(new_n9559_), .ZN(new_n9560_));
  NOR3_X1    g06741(.A1(new_n9428_), .A2(new_n6573_), .A3(new_n9134_), .ZN(new_n9561_));
  AOI21_X1   g06742(.A1(new_n6572_), .A2(new_n9134_), .B(new_n9427_), .ZN(new_n9562_));
  OAI21_X1   g06743(.A1(new_n9561_), .A2(new_n9562_), .B(new_n6088_), .ZN(new_n9563_));
  AOI21_X1   g06744(.A1(new_n9448_), .A2(new_n6209_), .B(pi0592), .ZN(new_n9564_));
  AOI21_X1   g06745(.A1(new_n9450_), .A2(new_n6572_), .B(new_n6088_), .ZN(new_n9565_));
  OAI21_X1   g06746(.A1(new_n9138_), .A2(new_n9564_), .B(new_n9565_), .ZN(new_n9566_));
  NAND2_X1   g06747(.A1(new_n9566_), .A2(new_n9563_), .ZN(new_n9567_));
  MUX2_X1    g06748(.I0(new_n9567_), .I1(new_n9560_), .S(new_n9274_), .Z(new_n9568_));
  INV_X1     g06749(.I(pi0391), .ZN(new_n9569_));
  NOR2_X1    g06750(.A1(new_n6539_), .A2(new_n9560_), .ZN(new_n9570_));
  AOI21_X1   g06751(.A1(new_n9567_), .A2(new_n6539_), .B(new_n9570_), .ZN(new_n9571_));
  NOR2_X1    g06752(.A1(new_n9571_), .A2(pi0333), .ZN(new_n9572_));
  NOR2_X1    g06753(.A1(new_n9572_), .A2(new_n9569_), .ZN(new_n9573_));
  OAI21_X1   g06754(.A1(new_n6286_), .A2(new_n9568_), .B(new_n9573_), .ZN(new_n9574_));
  NOR2_X1    g06755(.A1(new_n9568_), .A2(pi0333), .ZN(new_n9575_));
  NOR2_X1    g06756(.A1(new_n9571_), .A2(new_n6286_), .ZN(new_n9576_));
  OAI21_X1   g06757(.A1(new_n9575_), .A2(new_n9576_), .B(pi0391), .ZN(new_n9577_));
  AOI21_X1   g06758(.A1(new_n9574_), .A2(new_n9577_), .B(new_n9558_), .ZN(new_n9578_));
  NOR3_X1    g06759(.A1(new_n9575_), .A2(pi0391), .A3(new_n9576_), .ZN(new_n9579_));
  NAND2_X1   g06760(.A1(new_n9574_), .A2(new_n9558_), .ZN(new_n9580_));
  NOR2_X1    g06761(.A1(new_n9580_), .A2(new_n9579_), .ZN(new_n9581_));
  MUX2_X1    g06762(.I0(new_n6912_), .I1(pi0592), .S(new_n6156_), .Z(new_n9582_));
  AOI21_X1   g06763(.A1(new_n6920_), .A2(new_n6925_), .B(new_n6432_), .ZN(new_n9583_));
  AOI21_X1   g06764(.A1(new_n9583_), .A2(new_n9582_), .B(new_n9135_), .ZN(new_n9584_));
  AOI21_X1   g06765(.A1(new_n9584_), .A2(new_n6203_), .B(pi0591), .ZN(new_n9585_));
  OAI21_X1   g06766(.A1(new_n9581_), .A2(new_n9578_), .B(new_n9585_), .ZN(new_n9586_));
  NOR3_X1    g06767(.A1(new_n6891_), .A2(new_n6852_), .A3(new_n9135_), .ZN(new_n9587_));
  NOR2_X1    g06768(.A1(new_n9587_), .A2(new_n6522_), .ZN(new_n9588_));
  NOR2_X1    g06769(.A1(new_n9588_), .A2(new_n9559_), .ZN(new_n9589_));
  OAI21_X1   g06770(.A1(new_n9587_), .A2(new_n6493_), .B(new_n9560_), .ZN(new_n9590_));
  MUX2_X1    g06771(.I0(new_n9590_), .I1(new_n9589_), .S(new_n6180_), .Z(new_n9591_));
  NOR2_X1    g06772(.A1(new_n9591_), .A2(pi0356), .ZN(new_n9592_));
  NOR2_X1    g06773(.A1(new_n9587_), .A2(new_n6493_), .ZN(new_n9593_));
  NOR2_X1    g06774(.A1(new_n9593_), .A2(new_n9559_), .ZN(new_n9594_));
  MUX2_X1    g06775(.I0(new_n9594_), .I1(new_n9589_), .S(new_n6180_), .Z(new_n9595_));
  NOR2_X1    g06776(.A1(new_n9595_), .A2(new_n6198_), .ZN(new_n9596_));
  OR2_X2     g06777(.A1(new_n9595_), .A2(pi0356), .Z(new_n9597_));
  OAI21_X1   g06778(.A1(new_n9591_), .A2(new_n6198_), .B(new_n9597_), .ZN(new_n9598_));
  OAI22_X1   g06779(.A1(new_n9598_), .A2(pi0354), .B1(new_n9592_), .B2(new_n9596_), .ZN(new_n9599_));
  NOR2_X1    g06780(.A1(new_n9592_), .A2(new_n9596_), .ZN(new_n9600_));
  NAND3_X1   g06781(.A1(new_n9598_), .A2(new_n6192_), .A3(new_n9600_), .ZN(new_n9601_));
  NAND2_X1   g06782(.A1(new_n9598_), .A2(pi0354), .ZN(new_n9602_));
  AND3_X2    g06783(.A1(new_n9600_), .A2(pi0354), .A3(new_n6196_), .Z(new_n9603_));
  NAND2_X1   g06784(.A1(new_n6196_), .A2(new_n5940_), .ZN(new_n9604_));
  AOI21_X1   g06785(.A1(new_n9602_), .A2(new_n9603_), .B(new_n9604_), .ZN(new_n9605_));
  NAND3_X1   g06786(.A1(new_n9605_), .A2(new_n9599_), .A3(new_n9601_), .ZN(new_n9606_));
  AOI21_X1   g06787(.A1(new_n9606_), .A2(new_n9136_), .B(pi0588), .ZN(new_n9607_));
  INV_X1     g06788(.I(new_n9299_), .ZN(new_n9608_));
  OAI21_X1   g06789(.A1(new_n6084_), .A2(new_n6743_), .B(new_n6932_), .ZN(new_n9609_));
  AND3_X2    g06790(.A1(new_n9609_), .A2(new_n6851_), .A3(new_n9135_), .Z(new_n9610_));
  INV_X1     g06791(.I(new_n9610_), .ZN(new_n9611_));
  MUX2_X1    g06792(.I0(new_n9611_), .I1(new_n9560_), .S(new_n6766_), .Z(new_n9612_));
  XNOR2_X1   g06793(.A1(pi0427), .A2(pi0428), .ZN(new_n9613_));
  NOR2_X1    g06794(.A1(new_n6712_), .A2(new_n9613_), .ZN(new_n9614_));
  XOR2_X1    g06795(.A1(new_n9612_), .A2(new_n9614_), .Z(new_n9615_));
  NAND2_X1   g06796(.A1(new_n6773_), .A2(new_n9613_), .ZN(new_n9616_));
  XOR2_X1    g06797(.A1(new_n9612_), .A2(new_n9616_), .Z(new_n9617_));
  NAND2_X1   g06798(.A1(new_n9617_), .A2(pi0445), .ZN(new_n9618_));
  OAI21_X1   g06799(.A1(pi0445), .A2(new_n9615_), .B(new_n9618_), .ZN(new_n9619_));
  XNOR2_X1   g06800(.A1(pi0426), .A2(pi0430), .ZN(new_n9620_));
  NOR2_X1    g06801(.A1(new_n9620_), .A2(new_n6781_), .ZN(new_n9621_));
  XOR2_X1    g06802(.A1(new_n9619_), .A2(new_n9621_), .Z(new_n9622_));
  NAND2_X1   g06803(.A1(new_n9622_), .A2(new_n6924_), .ZN(new_n9623_));
  NAND2_X1   g06804(.A1(new_n9617_), .A2(new_n6772_), .ZN(new_n9624_));
  OAI21_X1   g06805(.A1(new_n6772_), .A2(new_n9615_), .B(new_n9624_), .ZN(new_n9625_));
  XOR2_X1    g06806(.A1(new_n9625_), .A2(new_n9621_), .Z(new_n9626_));
  NAND2_X1   g06807(.A1(new_n9626_), .A2(new_n6791_), .ZN(new_n9627_));
  OAI21_X1   g06808(.A1(new_n9611_), .A2(new_n6798_), .B(new_n6088_), .ZN(new_n9628_));
  AOI21_X1   g06809(.A1(new_n9623_), .A2(new_n9627_), .B(new_n9628_), .ZN(new_n9629_));
  OAI21_X1   g06810(.A1(new_n9629_), .A2(new_n9608_), .B(new_n6844_), .ZN(new_n9630_));
  AOI21_X1   g06811(.A1(new_n9586_), .A2(new_n9607_), .B(new_n9630_), .ZN(new_n9631_));
  INV_X1     g06812(.I(pi0080), .ZN(new_n9632_));
  NAND4_X1   g06813(.A1(new_n6845_), .A2(new_n9134_), .A3(new_n9632_), .A4(new_n6538_), .ZN(new_n9633_));
  NOR3_X1    g06814(.A1(po1038), .A2(pi0080), .A3(pi0217), .ZN(new_n9634_));
  OAI21_X1   g06815(.A1(new_n9631_), .A2(new_n9633_), .B(new_n9634_), .ZN(new_n9635_));
  AOI21_X1   g06816(.A1(new_n9516_), .A2(new_n9557_), .B(new_n9635_), .ZN(new_n9636_));
  INV_X1     g06817(.I(pi0217), .ZN(new_n9637_));
  NOR2_X1    g06818(.A1(new_n6953_), .A2(new_n9637_), .ZN(new_n9638_));
  OAI21_X1   g06819(.A1(new_n9134_), .A2(pi0080), .B(new_n9638_), .ZN(new_n9639_));
  AOI21_X1   g06820(.A1(new_n9340_), .A2(new_n9636_), .B(new_n9639_), .ZN(po0238));
  INV_X1     g06821(.I(new_n8573_), .ZN(new_n9641_));
  NOR3_X1    g06822(.A1(new_n2699_), .A2(new_n2441_), .A3(pi0314), .ZN(new_n9642_));
  NOR4_X1    g06823(.A1(new_n2757_), .A2(pi0036), .A3(pi0064), .A4(pi0081), .ZN(new_n9643_));
  NAND4_X1   g06824(.A1(new_n8389_), .A2(new_n7005_), .A3(new_n2775_), .A4(new_n9643_), .ZN(new_n9644_));
  NOR2_X1    g06825(.A1(new_n2776_), .A2(new_n9644_), .ZN(new_n9645_));
  NOR4_X1    g06826(.A1(new_n9641_), .A2(po1038), .A3(new_n9642_), .A4(new_n9645_), .ZN(po0239));
  NOR3_X1    g06827(.A1(new_n2783_), .A2(new_n5276_), .A3(pi0067), .ZN(new_n9647_));
  NOR3_X1    g06828(.A1(new_n2786_), .A2(new_n2731_), .A3(pi0073), .ZN(new_n9648_));
  AOI22_X1   g06829(.A1(new_n2779_), .A2(new_n9647_), .B1(new_n2448_), .B2(new_n9648_), .ZN(new_n9649_));
  NOR4_X1    g06830(.A1(new_n8438_), .A2(new_n7888_), .A3(new_n8439_), .A4(new_n9649_), .ZN(po0240));
  NAND3_X1   g06831(.A1(new_n2762_), .A2(new_n2767_), .A3(new_n2775_), .ZN(new_n9651_));
  NOR4_X1    g06832(.A1(new_n9651_), .A2(pi0068), .A3(new_n2766_), .A4(new_n2786_), .ZN(new_n9652_));
  NOR2_X1    g06833(.A1(new_n8439_), .A2(new_n6999_), .ZN(new_n9653_));
  OAI21_X1   g06834(.A1(new_n9652_), .A2(pi0083), .B(new_n9653_), .ZN(new_n9654_));
  OAI21_X1   g06835(.A1(new_n9654_), .A2(new_n2790_), .B(pi0314), .ZN(new_n9655_));
  NAND4_X1   g06836(.A1(new_n9652_), .A2(pi0314), .A3(new_n2449_), .A4(new_n9653_), .ZN(new_n9656_));
  AOI21_X1   g06837(.A1(new_n9655_), .A2(new_n9656_), .B(new_n7829_), .ZN(po0241));
  NOR2_X1    g06838(.A1(pi0211), .A2(pi0219), .ZN(new_n9658_));
  INV_X1     g06839(.I(new_n9658_), .ZN(new_n9659_));
  MUX2_X1    g06840(.I0(new_n9659_), .I1(new_n8161_), .S(new_n2587_), .Z(new_n9660_));
  NOR3_X1    g06841(.A1(new_n8629_), .A2(po1038), .A3(new_n9660_), .ZN(po0242));
  NAND3_X1   g06842(.A1(new_n8661_), .A2(new_n5276_), .A3(new_n8443_), .ZN(new_n9662_));
  NAND3_X1   g06843(.A1(new_n5263_), .A2(new_n8440_), .A3(new_n8441_), .ZN(new_n9663_));
  AOI21_X1   g06844(.A1(new_n9662_), .A2(new_n9663_), .B(new_n8438_), .ZN(po0243));
  AOI22_X1   g06845(.A1(new_n6049_), .A2(new_n8634_), .B1(new_n6054_), .B2(new_n8636_), .ZN(new_n9665_));
  NOR2_X1    g06846(.A1(new_n9665_), .A2(new_n8371_), .ZN(po0244));
  NOR2_X1    g06847(.A1(new_n8439_), .A2(new_n2469_), .ZN(new_n9667_));
  NAND2_X1   g06848(.A1(new_n2796_), .A2(new_n9667_), .ZN(new_n9668_));
  NOR4_X1    g06849(.A1(new_n7829_), .A2(new_n5276_), .A3(new_n2640_), .A4(new_n9668_), .ZN(po0245));
  OAI21_X1   g06850(.A1(new_n8408_), .A2(new_n6005_), .B(new_n2924_), .ZN(new_n9670_));
  NOR2_X1    g06851(.A1(new_n6986_), .A2(new_n2678_), .ZN(new_n9671_));
  NOR3_X1    g06852(.A1(new_n8406_), .A2(new_n5958_), .A3(new_n9145_), .ZN(new_n9672_));
  NAND4_X1   g06853(.A1(new_n9672_), .A2(new_n6004_), .A3(new_n8548_), .A4(new_n9671_), .ZN(new_n9673_));
  NOR4_X1    g06854(.A1(new_n9673_), .A2(pi1093), .A3(new_n3233_), .A4(new_n7757_), .ZN(new_n9674_));
  NAND2_X1   g06855(.A1(new_n9670_), .A2(new_n9674_), .ZN(new_n9675_));
  INV_X1     g06856(.I(new_n8678_), .ZN(new_n9676_));
  NOR2_X1    g06857(.A1(new_n2652_), .A2(new_n6005_), .ZN(new_n9677_));
  NOR3_X1    g06858(.A1(new_n2485_), .A2(new_n2710_), .A3(pi1093), .ZN(new_n9678_));
  NAND4_X1   g06859(.A1(new_n7818_), .A2(new_n3233_), .A3(new_n9677_), .A4(new_n9678_), .ZN(new_n9679_));
  OAI21_X1   g06860(.A1(new_n9676_), .A2(new_n9679_), .B(new_n6844_), .ZN(new_n9680_));
  NAND2_X1   g06861(.A1(new_n9680_), .A2(new_n6845_), .ZN(new_n9681_));
  AOI21_X1   g06862(.A1(new_n9675_), .A2(new_n6538_), .B(new_n9681_), .ZN(po0246));
  NOR4_X1    g06863(.A1(new_n7841_), .A2(new_n2464_), .A3(new_n6999_), .A4(new_n7072_), .ZN(new_n9683_));
  INV_X1     g06864(.I(new_n9683_), .ZN(new_n9684_));
  NOR3_X1    g06865(.A1(new_n9684_), .A2(new_n2902_), .A3(new_n5965_), .ZN(new_n9685_));
  NAND3_X1   g06866(.A1(new_n7824_), .A2(new_n2849_), .A3(new_n2488_), .ZN(new_n9686_));
  OAI21_X1   g06867(.A1(new_n9686_), .A2(new_n9685_), .B(new_n2849_), .ZN(new_n9687_));
  NOR2_X1    g06868(.A1(new_n6970_), .A2(new_n9687_), .ZN(po0247));
  NAND3_X1   g06869(.A1(new_n7232_), .A2(new_n8684_), .A3(new_n2455_), .ZN(new_n9689_));
  AOI21_X1   g06870(.A1(new_n9689_), .A2(new_n2839_), .B(new_n8590_), .ZN(new_n9690_));
  NOR4_X1    g06871(.A1(new_n9690_), .A2(pi0090), .A3(new_n2902_), .A4(new_n2642_), .ZN(po0248));
  AOI21_X1   g06872(.A1(new_n7368_), .A2(new_n2844_), .B(new_n7820_), .ZN(new_n9692_));
  NAND4_X1   g06873(.A1(new_n3082_), .A2(pi0024), .A3(new_n2666_), .A4(new_n8589_), .ZN(new_n9693_));
  NOR3_X1    g06874(.A1(new_n3082_), .A2(pi0039), .A3(new_n7827_), .ZN(new_n9694_));
  OAI21_X1   g06875(.A1(new_n6018_), .A2(new_n9693_), .B(new_n9694_), .ZN(new_n9695_));
  OAI21_X1   g06876(.A1(new_n9692_), .A2(new_n9695_), .B(new_n7832_), .ZN(new_n9696_));
  NOR2_X1    g06877(.A1(new_n6063_), .A2(new_n9696_), .ZN(po0249));
  NOR2_X1    g06878(.A1(new_n3203_), .A2(pi0314), .ZN(new_n9698_));
  NAND4_X1   g06879(.A1(new_n2490_), .A2(pi1050), .A3(new_n3322_), .A4(new_n9698_), .ZN(new_n9699_));
  NOR3_X1    g06880(.A1(new_n7880_), .A2(new_n2562_), .A3(new_n2550_), .ZN(new_n9700_));
  NAND2_X1   g06881(.A1(new_n6054_), .A2(new_n9700_), .ZN(new_n9701_));
  NOR3_X1    g06882(.A1(new_n3294_), .A2(new_n2588_), .A3(new_n2595_), .ZN(new_n9702_));
  NAND2_X1   g06883(.A1(new_n6049_), .A2(new_n9702_), .ZN(new_n9703_));
  NAND4_X1   g06884(.A1(new_n9701_), .A2(new_n9703_), .A3(new_n2536_), .A4(new_n8534_), .ZN(new_n9704_));
  AOI21_X1   g06885(.A1(new_n9704_), .A2(new_n9699_), .B(new_n7823_), .ZN(po0250));
  NAND4_X1   g06886(.A1(new_n2669_), .A2(pi0093), .A3(pi0841), .A4(new_n8589_), .ZN(new_n9706_));
  NAND2_X1   g06887(.A1(new_n9706_), .A2(new_n3203_), .ZN(new_n9707_));
  NOR2_X1    g06888(.A1(new_n7823_), .A2(new_n3323_), .ZN(new_n9708_));
  NAND3_X1   g06889(.A1(new_n2490_), .A2(new_n3203_), .A3(new_n8684_), .ZN(new_n9709_));
  AOI21_X1   g06890(.A1(new_n9707_), .A2(new_n9708_), .B(new_n9709_), .ZN(po0251));
  NAND2_X1   g06891(.A1(new_n8430_), .A2(new_n8562_), .ZN(new_n9711_));
  NAND3_X1   g06892(.A1(new_n2957_), .A2(new_n2921_), .A3(new_n2924_), .ZN(new_n9712_));
  INV_X1     g06893(.I(new_n8429_), .ZN(new_n9713_));
  AOI21_X1   g06894(.A1(new_n7898_), .A2(new_n9713_), .B(new_n2820_), .ZN(new_n9714_));
  NAND3_X1   g06895(.A1(new_n8548_), .A2(pi0252), .A3(new_n2889_), .ZN(new_n9715_));
  OAI22_X1   g06896(.A1(new_n9714_), .A2(new_n9715_), .B1(new_n9711_), .B2(new_n9712_), .ZN(new_n9716_));
  OAI21_X1   g06897(.A1(new_n9716_), .A2(po0840), .B(new_n9711_), .ZN(new_n9717_));
  NAND2_X1   g06898(.A1(new_n9716_), .A2(pi0252), .ZN(new_n9718_));
  NAND2_X1   g06899(.A1(new_n9717_), .A2(new_n9718_), .ZN(new_n9719_));
  NAND3_X1   g06900(.A1(new_n9719_), .A2(new_n6972_), .A3(new_n9711_), .ZN(new_n9720_));
  INV_X1     g06901(.I(new_n9711_), .ZN(new_n9721_));
  OAI21_X1   g06902(.A1(new_n9719_), .A2(new_n6973_), .B(new_n9721_), .ZN(new_n9722_));
  AOI21_X1   g06903(.A1(new_n9722_), .A2(new_n9720_), .B(new_n7825_), .ZN(po0252));
  NAND4_X1   g06904(.A1(new_n2483_), .A2(pi0024), .A3(new_n2632_), .A4(pi0095), .ZN(new_n9724_));
  NOR4_X1    g06905(.A1(new_n7827_), .A2(pi0332), .A3(pi0841), .A4(new_n2650_), .ZN(new_n9725_));
  AOI21_X1   g06906(.A1(new_n9725_), .A2(new_n9683_), .B(pi0039), .ZN(new_n9726_));
  OAI21_X1   g06907(.A1(new_n2654_), .A2(new_n9724_), .B(new_n9726_), .ZN(new_n9727_));
  NOR3_X1    g06908(.A1(new_n8651_), .A2(new_n2631_), .A3(new_n8649_), .ZN(new_n9728_));
  OAI21_X1   g06909(.A1(new_n2601_), .A2(new_n8649_), .B(new_n3295_), .ZN(new_n9729_));
  NOR2_X1    g06910(.A1(new_n5145_), .A2(new_n9729_), .ZN(new_n9730_));
  OAI21_X1   g06911(.A1(new_n9728_), .A2(new_n9730_), .B(new_n3154_), .ZN(new_n9731_));
  AOI21_X1   g06912(.A1(new_n7855_), .A2(new_n9727_), .B(new_n9731_), .ZN(po0253));
  NAND2_X1   g06913(.A1(new_n6979_), .A2(pi0479), .ZN(new_n9733_));
  NAND4_X1   g06914(.A1(new_n9733_), .A2(pi0096), .A3(new_n2512_), .A4(new_n5951_), .ZN(new_n9734_));
  NOR4_X1    g06915(.A1(new_n2904_), .A2(pi0051), .A3(pi0072), .A4(new_n9734_), .ZN(new_n9735_));
  NOR2_X1    g06916(.A1(new_n3101_), .A2(new_n9733_), .ZN(new_n9736_));
  OAI21_X1   g06917(.A1(new_n9735_), .A2(new_n9736_), .B(new_n2437_), .ZN(new_n9737_));
  NAND4_X1   g06918(.A1(new_n8061_), .A2(new_n2632_), .A3(pi0095), .A4(new_n2483_), .ZN(new_n9738_));
  AOI21_X1   g06919(.A1(new_n9737_), .A2(new_n9738_), .B(new_n7825_), .ZN(po0254));
  NAND3_X1   g06920(.A1(new_n8653_), .A2(pi0039), .A3(pi0593), .ZN(new_n9740_));
  OAI21_X1   g06921(.A1(new_n9733_), .A2(new_n5080_), .B(new_n5943_), .ZN(new_n9741_));
  NOR2_X1    g06922(.A1(pi0039), .A2(pi0096), .ZN(new_n9742_));
  NAND4_X1   g06923(.A1(new_n8696_), .A2(new_n3418_), .A3(new_n9741_), .A4(new_n9742_), .ZN(new_n9743_));
  AOI21_X1   g06924(.A1(new_n9740_), .A2(new_n9743_), .B(new_n7856_), .ZN(po0255));
  NAND3_X1   g06925(.A1(new_n8686_), .A2(pi0092), .A3(new_n2490_), .ZN(new_n9745_));
  OAI21_X1   g06926(.A1(new_n3203_), .A2(new_n2490_), .B(new_n8685_), .ZN(new_n9746_));
  NAND3_X1   g06927(.A1(new_n9708_), .A2(pi0314), .A3(pi1050), .ZN(new_n9747_));
  AOI21_X1   g06928(.A1(new_n9745_), .A2(new_n9746_), .B(new_n9747_), .ZN(po0256));
  NOR2_X1    g06929(.A1(new_n8115_), .A2(pi0072), .ZN(new_n9749_));
  INV_X1     g06930(.I(new_n9749_), .ZN(new_n9750_));
  NOR4_X1    g06931(.A1(new_n8163_), .A2(pi0072), .A3(new_n3250_), .A4(new_n4701_), .ZN(new_n9751_));
  NAND2_X1   g06932(.A1(new_n9751_), .A2(pi0232), .ZN(new_n9752_));
  MUX2_X1    g06933(.I0(new_n9752_), .I1(new_n9750_), .S(new_n3154_), .Z(new_n9753_));
  AOI22_X1   g06934(.A1(new_n8064_), .A2(new_n9749_), .B1(new_n5173_), .B2(new_n8327_), .ZN(new_n9754_));
  NOR3_X1    g06935(.A1(new_n8025_), .A2(new_n2922_), .A3(new_n8040_), .ZN(new_n9755_));
  INV_X1     g06936(.I(new_n9755_), .ZN(new_n9756_));
  AOI21_X1   g06937(.A1(new_n8026_), .A2(new_n9750_), .B(pi0039), .ZN(new_n9757_));
  OAI21_X1   g06938(.A1(new_n9754_), .A2(new_n9756_), .B(new_n9757_), .ZN(new_n9758_));
  NAND4_X1   g06939(.A1(new_n8013_), .A2(new_n2861_), .A3(pi0174), .A4(new_n2587_), .ZN(new_n9759_));
  NAND2_X1   g06940(.A1(new_n9751_), .A2(pi0299), .ZN(new_n9760_));
  XNOR2_X1   g06941(.A1(new_n9760_), .A2(new_n9759_), .ZN(new_n9761_));
  NAND2_X1   g06942(.A1(new_n9761_), .A2(pi0232), .ZN(new_n9762_));
  NAND2_X1   g06943(.A1(new_n9762_), .A2(pi0039), .ZN(new_n9763_));
  NAND3_X1   g06944(.A1(new_n9758_), .A2(new_n3207_), .A3(new_n9763_), .ZN(new_n9764_));
  INV_X1     g06945(.I(new_n9763_), .ZN(new_n9765_));
  AOI21_X1   g06946(.A1(new_n3154_), .A2(new_n9750_), .B(new_n9765_), .ZN(new_n9766_));
  INV_X1     g06947(.I(new_n9766_), .ZN(new_n9767_));
  NOR3_X1    g06948(.A1(new_n9767_), .A2(pi0075), .A3(new_n3207_), .ZN(new_n9768_));
  AOI21_X1   g06949(.A1(pi0041), .A2(pi0072), .B(new_n8115_), .ZN(new_n9769_));
  NAND2_X1   g06950(.A1(new_n7973_), .A2(new_n9769_), .ZN(new_n9770_));
  NAND2_X1   g06951(.A1(new_n9770_), .A2(new_n8264_), .ZN(new_n9771_));
  INV_X1     g06952(.I(new_n8263_), .ZN(new_n9772_));
  NAND3_X1   g06953(.A1(new_n9772_), .A2(new_n7956_), .A3(new_n9769_), .ZN(new_n9773_));
  AOI21_X1   g06954(.A1(new_n9773_), .A2(new_n9771_), .B(pi0228), .ZN(new_n9774_));
  NAND2_X1   g06955(.A1(new_n9761_), .A2(new_n7927_), .ZN(new_n9775_));
  NOR2_X1    g06956(.A1(pi0039), .A2(pi0228), .ZN(new_n9776_));
  OAI21_X1   g06957(.A1(new_n8350_), .A2(new_n9775_), .B(new_n9776_), .ZN(new_n9777_));
  NOR2_X1    g06958(.A1(new_n8152_), .A2(new_n9777_), .ZN(new_n9778_));
  OAI21_X1   g06959(.A1(new_n8001_), .A2(new_n9769_), .B(new_n9778_), .ZN(new_n9779_));
  NOR2_X1    g06960(.A1(new_n8034_), .A2(new_n9750_), .ZN(new_n9780_));
  OAI21_X1   g06961(.A1(new_n8067_), .A2(new_n5172_), .B(new_n9755_), .ZN(new_n9781_));
  OAI21_X1   g06962(.A1(new_n9780_), .A2(new_n9781_), .B(new_n9757_), .ZN(new_n9782_));
  NOR2_X1    g06963(.A1(new_n9765_), .A2(new_n5158_), .ZN(new_n9783_));
  OAI21_X1   g06964(.A1(new_n9767_), .A2(pi0038), .B(new_n8308_), .ZN(new_n9784_));
  AOI21_X1   g06965(.A1(new_n9782_), .A2(new_n9783_), .B(new_n9784_), .ZN(new_n9785_));
  OAI21_X1   g06966(.A1(new_n9774_), .A2(new_n9779_), .B(new_n9785_), .ZN(new_n9786_));
  NOR3_X1    g06967(.A1(new_n8036_), .A2(new_n2523_), .A3(new_n5172_), .ZN(new_n9787_));
  NOR4_X1    g06968(.A1(new_n9787_), .A2(new_n2523_), .A3(new_n2546_), .A4(new_n9749_), .ZN(new_n9788_));
  NAND3_X1   g06969(.A1(new_n8032_), .A2(new_n8029_), .A3(new_n9788_), .ZN(new_n9789_));
  AOI21_X1   g06970(.A1(new_n9767_), .A2(new_n2547_), .B(new_n3177_), .ZN(new_n9790_));
  AOI21_X1   g06971(.A1(new_n9790_), .A2(new_n9789_), .B(pi0075), .ZN(new_n9791_));
  AOI22_X1   g06972(.A1(new_n9786_), .A2(new_n9791_), .B1(new_n9764_), .B2(new_n9768_), .ZN(new_n9792_));
  NAND2_X1   g06973(.A1(po1038), .A2(new_n5941_), .ZN(new_n9793_));
  OAI22_X1   g06974(.A1(new_n9792_), .A2(new_n9793_), .B1(new_n6845_), .B2(new_n9753_), .ZN(po0257));
  NAND4_X1   g06975(.A1(new_n6974_), .A2(new_n5895_), .A3(po0840), .A4(new_n7797_), .ZN(new_n9795_));
  NOR2_X1    g06976(.A1(new_n5985_), .A2(pi0129), .ZN(new_n9796_));
  NAND2_X1   g06977(.A1(new_n7760_), .A2(pi0129), .ZN(new_n9797_));
  AOI22_X1   g06978(.A1(new_n7765_), .A2(new_n9796_), .B1(new_n9797_), .B2(new_n7762_), .ZN(new_n9798_));
  OR2_X2     g06979(.A1(new_n5187_), .A2(new_n6975_), .Z(new_n9799_));
  NOR3_X1    g06980(.A1(new_n5159_), .A2(pi0075), .A3(new_n2624_), .ZN(new_n9800_));
  OAI21_X1   g06981(.A1(new_n9798_), .A2(new_n9799_), .B(new_n9800_), .ZN(new_n9801_));
  NAND2_X1   g06982(.A1(new_n2490_), .A2(new_n6966_), .ZN(new_n9802_));
  AOI21_X1   g06983(.A1(new_n9801_), .A2(new_n9795_), .B(new_n9802_), .ZN(po0258));
  INV_X1     g06984(.I(new_n8028_), .ZN(new_n9804_));
  NOR3_X1    g06985(.A1(new_n3247_), .A2(new_n5109_), .A3(new_n3250_), .ZN(new_n9805_));
  INV_X1     g06986(.I(new_n9805_), .ZN(new_n9806_));
  NOR2_X1    g06987(.A1(new_n9806_), .A2(pi0072), .ZN(new_n9807_));
  NAND2_X1   g06988(.A1(new_n9807_), .A2(pi0232), .ZN(new_n9808_));
  MUX2_X1    g06989(.I0(new_n9808_), .I1(new_n9804_), .S(new_n3154_), .Z(new_n9809_));
  AOI21_X1   g06990(.A1(new_n7954_), .A2(new_n7974_), .B(new_n7968_), .ZN(new_n9810_));
  NOR3_X1    g06991(.A1(new_n7969_), .A2(pi0101), .A3(new_n7974_), .ZN(new_n9811_));
  AND2_X2    g06992(.A1(new_n7952_), .A2(pi0101), .Z(new_n9812_));
  AOI21_X1   g06993(.A1(new_n7961_), .A2(new_n7960_), .B(pi0101), .ZN(new_n9813_));
  OAI21_X1   g06994(.A1(new_n9812_), .A2(new_n9813_), .B(new_n2922_), .ZN(new_n9814_));
  NOR3_X1    g06995(.A1(new_n9814_), .A2(new_n9810_), .A3(new_n9811_), .ZN(new_n9815_));
  NOR2_X1    g06996(.A1(new_n7998_), .A2(new_n7954_), .ZN(new_n9816_));
  AOI21_X1   g06997(.A1(new_n8005_), .A2(new_n7933_), .B(new_n7954_), .ZN(new_n9817_));
  NOR4_X1    g06998(.A1(new_n9816_), .A2(pi0039), .A3(pi0228), .A4(new_n9817_), .ZN(new_n9818_));
  OAI21_X1   g06999(.A1(new_n9815_), .A2(new_n2523_), .B(new_n9818_), .ZN(new_n9819_));
  NAND4_X1   g07000(.A1(new_n8352_), .A2(new_n7504_), .A3(pi0174), .A4(new_n8011_), .ZN(new_n9820_));
  AOI21_X1   g07001(.A1(new_n9820_), .A2(new_n2587_), .B(new_n7927_), .ZN(new_n9821_));
  NOR2_X1    g07002(.A1(new_n8351_), .A2(new_n9806_), .ZN(new_n9822_));
  NOR4_X1    g07003(.A1(new_n9821_), .A2(new_n2587_), .A3(new_n2621_), .A4(new_n9822_), .ZN(new_n9823_));
  AOI21_X1   g07004(.A1(new_n8026_), .A2(new_n9804_), .B(pi0039), .ZN(new_n9824_));
  NOR3_X1    g07005(.A1(new_n8025_), .A2(new_n2922_), .A3(new_n5175_), .ZN(new_n9825_));
  NOR3_X1    g07006(.A1(new_n8175_), .A2(new_n6436_), .A3(new_n8028_), .ZN(new_n9826_));
  OAI21_X1   g07007(.A1(new_n9826_), .A2(new_n8037_), .B(new_n9825_), .ZN(new_n9827_));
  NOR4_X1    g07008(.A1(new_n9807_), .A2(pi0039), .A3(pi0232), .A4(new_n2587_), .ZN(new_n9829_));
  INV_X1     g07009(.I(new_n9829_), .ZN(new_n9830_));
  NAND2_X1   g07010(.A1(new_n9830_), .A2(new_n5159_), .ZN(new_n9831_));
  AOI21_X1   g07011(.A1(new_n9827_), .A2(new_n9824_), .B(new_n9831_), .ZN(new_n9832_));
  NAND2_X1   g07012(.A1(new_n9804_), .A2(new_n3154_), .ZN(new_n9833_));
  NAND2_X1   g07013(.A1(new_n9830_), .A2(new_n9833_), .ZN(new_n9834_));
  OAI21_X1   g07014(.A1(new_n9834_), .A2(pi0038), .B(new_n3177_), .ZN(new_n9835_));
  NAND4_X1   g07015(.A1(new_n8032_), .A2(pi0228), .A3(new_n2621_), .A4(new_n9804_), .ZN(new_n9836_));
  NAND2_X1   g07016(.A1(new_n8364_), .A2(new_n7954_), .ZN(new_n9837_));
  NAND4_X1   g07017(.A1(new_n9836_), .A2(new_n3154_), .A3(new_n9830_), .A4(new_n9837_), .ZN(new_n9838_));
  AOI21_X1   g07018(.A1(new_n9838_), .A2(new_n3177_), .B(pi0075), .ZN(new_n9839_));
  OAI21_X1   g07019(.A1(new_n9832_), .A2(new_n9835_), .B(new_n9839_), .ZN(new_n9840_));
  AOI21_X1   g07020(.A1(new_n9819_), .A2(new_n9823_), .B(new_n9840_), .ZN(new_n9841_));
  NAND4_X1   g07021(.A1(new_n9830_), .A2(new_n2628_), .A3(new_n3208_), .A4(new_n9833_), .ZN(new_n9847_));
  NOR2_X1    g07022(.A1(new_n6845_), .A2(new_n5942_), .ZN(new_n9849_));
  NAND2_X1   g07023(.A1(new_n9847_), .A2(new_n9849_), .ZN(new_n9850_));
  OAI22_X1   g07024(.A1(new_n9841_), .A2(new_n9850_), .B1(new_n6845_), .B2(new_n9809_), .ZN(po0259));
  NAND4_X1   g07025(.A1(new_n2807_), .A2(new_n2454_), .A3(new_n2441_), .A4(new_n2455_), .ZN(new_n9852_));
  NOR3_X1    g07026(.A1(new_n9641_), .A2(po1038), .A3(new_n9852_), .ZN(po0260));
  AOI21_X1   g07027(.A1(new_n2470_), .A2(new_n9668_), .B(new_n5284_), .ZN(new_n9854_));
  NOR4_X1    g07028(.A1(new_n2637_), .A2(new_n2470_), .A3(pi0314), .A4(new_n2678_), .ZN(new_n9855_));
  NAND2_X1   g07029(.A1(new_n2638_), .A2(new_n5276_), .ZN(new_n9856_));
  NOR4_X1    g07030(.A1(new_n7829_), .A2(new_n9854_), .A3(new_n9855_), .A4(new_n9856_), .ZN(po0261));
  NOR2_X1    g07031(.A1(new_n9673_), .A2(po1057), .ZN(new_n9858_));
  INV_X1     g07032(.I(new_n7757_), .ZN(new_n9859_));
  NAND2_X1   g07033(.A1(new_n8334_), .A2(new_n9859_), .ZN(new_n9860_));
  NOR2_X1    g07034(.A1(new_n9672_), .A2(pi0110), .ZN(new_n9861_));
  NAND3_X1   g07035(.A1(new_n8548_), .A2(new_n2661_), .A3(new_n6004_), .ZN(new_n9862_));
  NOR4_X1    g07036(.A1(new_n9861_), .A2(new_n6986_), .A3(new_n2835_), .A4(new_n9862_), .ZN(new_n9863_));
  OAI22_X1   g07037(.A1(po1057), .A2(new_n9863_), .B1(new_n9858_), .B2(new_n9860_), .ZN(new_n9864_));
  NOR2_X1    g07038(.A1(new_n8334_), .A2(new_n7757_), .ZN(new_n9865_));
  AOI21_X1   g07039(.A1(new_n9863_), .A2(new_n9865_), .B(new_n6538_), .ZN(new_n9866_));
  INV_X1     g07040(.I(new_n7758_), .ZN(new_n9867_));
  NAND3_X1   g07041(.A1(new_n6973_), .A2(new_n6538_), .A3(new_n9867_), .ZN(new_n9868_));
  OAI21_X1   g07042(.A1(new_n9868_), .A2(new_n8002_), .B(new_n7825_), .ZN(new_n9869_));
  AOI21_X1   g07043(.A1(new_n9864_), .A2(new_n9866_), .B(new_n9869_), .ZN(po0262));
  INV_X1     g07044(.I(new_n8547_), .ZN(new_n9871_));
  NAND2_X1   g07045(.A1(new_n9871_), .A2(new_n6995_), .ZN(new_n9872_));
  AOI21_X1   g07046(.A1(new_n2692_), .A2(new_n8560_), .B(new_n2884_), .ZN(new_n9873_));
  AND3_X2    g07047(.A1(new_n9873_), .A2(new_n5895_), .A3(new_n2889_), .Z(new_n9874_));
  NAND2_X1   g07048(.A1(new_n8561_), .A2(pi0024), .ZN(new_n9875_));
  OAI21_X1   g07049(.A1(new_n9874_), .A2(new_n9875_), .B(pi0841), .ZN(new_n9876_));
  AOI21_X1   g07050(.A1(new_n9874_), .A2(new_n9875_), .B(new_n9876_), .ZN(new_n9877_));
  NOR2_X1    g07051(.A1(new_n9877_), .A2(new_n9872_), .ZN(new_n9878_));
  AND2_X2    g07052(.A1(new_n9877_), .A2(new_n9872_), .Z(new_n9879_));
  NOR3_X1    g07053(.A1(new_n9879_), .A2(new_n7829_), .A3(new_n9878_), .ZN(po0264));
  NOR3_X1    g07054(.A1(new_n7829_), .A2(pi0999), .A3(new_n8610_), .ZN(po0265));
  INV_X1     g07055(.I(new_n7887_), .ZN(new_n9882_));
  AOI21_X1   g07056(.A1(new_n5961_), .A2(new_n2680_), .B(pi0108), .ZN(new_n9883_));
  NOR4_X1    g07057(.A1(new_n9882_), .A2(pi0047), .A3(new_n6986_), .A4(new_n9883_), .ZN(new_n9884_));
  INV_X1     g07058(.I(new_n9884_), .ZN(new_n9885_));
  OAI21_X1   g07059(.A1(new_n9885_), .A2(new_n5963_), .B(pi0314), .ZN(new_n9886_));
  NAND3_X1   g07060(.A1(new_n7900_), .A2(new_n2658_), .A3(new_n5966_), .ZN(new_n9887_));
  INV_X1     g07061(.I(new_n6030_), .ZN(new_n9888_));
  NOR2_X1    g07062(.A1(new_n9888_), .A2(new_n3198_), .ZN(new_n9889_));
  OAI21_X1   g07063(.A1(new_n9886_), .A2(new_n9887_), .B(new_n9889_), .ZN(new_n9890_));
  NAND2_X1   g07064(.A1(new_n5192_), .A2(new_n6966_), .ZN(new_n9891_));
  AOI21_X1   g07065(.A1(new_n9890_), .A2(new_n3177_), .B(new_n9891_), .ZN(po0266));
  NOR2_X1    g07066(.A1(new_n6999_), .A2(pi0050), .ZN(new_n9893_));
  NAND2_X1   g07067(.A1(new_n2707_), .A2(new_n9893_), .ZN(new_n9894_));
  NOR3_X1    g07068(.A1(new_n7829_), .A2(new_n5276_), .A3(new_n9894_), .ZN(po0267));
  NOR2_X1    g07069(.A1(new_n6973_), .A2(new_n9867_), .ZN(new_n9896_));
  INV_X1     g07070(.I(new_n9896_), .ZN(new_n9897_));
  NOR2_X1    g07071(.A1(new_n9897_), .A2(new_n7990_), .ZN(new_n9898_));
  INV_X1     g07072(.I(new_n2777_), .ZN(new_n9899_));
  NAND4_X1   g07073(.A1(new_n9671_), .A2(new_n7889_), .A3(new_n2470_), .A4(pi0111), .ZN(new_n9900_));
  NOR4_X1    g07074(.A1(new_n8444_), .A2(new_n2469_), .A3(new_n9899_), .A4(new_n9900_), .ZN(new_n9901_));
  INV_X1     g07075(.I(new_n9901_), .ZN(new_n9902_));
  OAI21_X1   g07076(.A1(new_n9902_), .A2(new_n5276_), .B(new_n7828_), .ZN(new_n9903_));
  NOR2_X1    g07077(.A1(new_n9898_), .A2(new_n9903_), .ZN(po0268));
  NAND2_X1   g07078(.A1(new_n9901_), .A2(new_n5276_), .ZN(new_n9905_));
  NOR2_X1    g07079(.A1(new_n7825_), .A2(new_n2515_), .ZN(new_n9906_));
  OAI21_X1   g07080(.A1(new_n9905_), .A2(new_n7250_), .B(new_n9906_), .ZN(new_n9907_));
  AOI21_X1   g07081(.A1(pi0072), .A2(new_n8061_), .B(new_n9907_), .ZN(po0269));
  INV_X1     g07082(.I(pi0468), .ZN(new_n9909_));
  NAND2_X1   g07083(.A1(new_n9909_), .A2(pi0124), .ZN(po0270));
  NOR2_X1    g07084(.A1(new_n8113_), .A2(pi0039), .ZN(new_n9911_));
  AOI22_X1   g07085(.A1(new_n8201_), .A2(new_n8112_), .B1(new_n8111_), .B2(new_n9787_), .ZN(new_n9912_));
  INV_X1     g07086(.I(new_n9911_), .ZN(new_n9913_));
  NOR2_X1    g07087(.A1(new_n9913_), .A2(new_n8309_), .ZN(new_n9914_));
  OAI21_X1   g07088(.A1(new_n9912_), .A2(new_n2547_), .B(new_n9914_), .ZN(new_n9915_));
  NOR2_X1    g07089(.A1(new_n7957_), .A2(new_n2922_), .ZN(new_n9916_));
  OAI21_X1   g07090(.A1(new_n7972_), .A2(new_n2921_), .B(new_n8115_), .ZN(new_n9917_));
  NOR3_X1    g07091(.A1(new_n5172_), .A2(pi0072), .A3(pi0113), .ZN(new_n9918_));
  OAI21_X1   g07092(.A1(new_n9916_), .A2(new_n9917_), .B(new_n9918_), .ZN(new_n9919_));
  NOR4_X1    g07093(.A1(new_n8263_), .A2(pi0113), .A3(pi0228), .A4(new_n8264_), .ZN(new_n9920_));
  INV_X1     g07094(.I(new_n8148_), .ZN(new_n9921_));
  OAI21_X1   g07095(.A1(pi0113), .A2(new_n8152_), .B(new_n9921_), .ZN(new_n9922_));
  NAND3_X1   g07096(.A1(new_n8148_), .A2(new_n8111_), .A3(new_n8152_), .ZN(new_n9923_));
  NAND3_X1   g07097(.A1(new_n9922_), .A2(new_n9776_), .A3(new_n9923_), .ZN(new_n9924_));
  AOI21_X1   g07098(.A1(new_n9919_), .A2(new_n9920_), .B(new_n9924_), .ZN(new_n9925_));
  INV_X1     g07099(.I(new_n8026_), .ZN(new_n9926_));
  NOR2_X1    g07100(.A1(new_n9926_), .A2(new_n5169_), .ZN(new_n9927_));
  NAND4_X1   g07101(.A1(new_n9927_), .A2(new_n8111_), .A3(new_n5171_), .A4(new_n8037_), .ZN(new_n9928_));
  NOR2_X1    g07102(.A1(new_n9926_), .A2(new_n8112_), .ZN(new_n9929_));
  NOR2_X1    g07103(.A1(new_n8177_), .A2(new_n6436_), .ZN(new_n9930_));
  OAI21_X1   g07104(.A1(new_n9930_), .A2(new_n5169_), .B(new_n9929_), .ZN(new_n9931_));
  NAND2_X1   g07105(.A1(new_n9931_), .A2(new_n9928_), .ZN(new_n9932_));
  NOR2_X1    g07106(.A1(new_n5158_), .A2(pi0039), .ZN(new_n9933_));
  OAI21_X1   g07107(.A1(new_n9913_), .A2(pi0038), .B(new_n3177_), .ZN(new_n9934_));
  AOI21_X1   g07108(.A1(new_n9932_), .A2(new_n9933_), .B(new_n9934_), .ZN(new_n9935_));
  OAI21_X1   g07109(.A1(new_n9925_), .A2(new_n2622_), .B(new_n9935_), .ZN(new_n9936_));
  OAI21_X1   g07110(.A1(new_n8217_), .A2(new_n5169_), .B(new_n9929_), .ZN(new_n9937_));
  OR2_X2     g07111(.A1(new_n9928_), .A2(new_n6435_), .Z(new_n9938_));
  AOI21_X1   g07112(.A1(new_n9937_), .A2(new_n9938_), .B(new_n2629_), .ZN(new_n9939_));
  NAND2_X1   g07113(.A1(new_n8341_), .A2(new_n9913_), .ZN(new_n9940_));
  OAI21_X1   g07114(.A1(new_n9939_), .A2(new_n9940_), .B(new_n2628_), .ZN(new_n9941_));
  AOI21_X1   g07115(.A1(new_n9936_), .A2(new_n9915_), .B(new_n9941_), .ZN(new_n9942_));
  MUX2_X1    g07116(.I0(new_n9942_), .I1(new_n9911_), .S(new_n6967_), .Z(po0271));
  NOR2_X1    g07117(.A1(new_n8138_), .A2(pi0072), .ZN(new_n9944_));
  INV_X1     g07118(.I(new_n9944_), .ZN(new_n9945_));
  NOR2_X1    g07119(.A1(new_n9945_), .A2(pi0039), .ZN(new_n9946_));
  NAND4_X1   g07120(.A1(new_n8294_), .A2(pi0114), .A3(new_n8214_), .A4(new_n8474_), .ZN(new_n9947_));
  AOI21_X1   g07121(.A1(new_n8474_), .A2(new_n9945_), .B(new_n2629_), .ZN(new_n9948_));
  NAND2_X1   g07122(.A1(new_n9947_), .A2(new_n9948_), .ZN(new_n9949_));
  NOR2_X1    g07123(.A1(new_n8342_), .A2(new_n9946_), .ZN(new_n9950_));
  NAND2_X1   g07124(.A1(new_n8257_), .A2(pi0114), .ZN(new_n9951_));
  OAI21_X1   g07125(.A1(pi0114), .A2(new_n8266_), .B(new_n9951_), .ZN(new_n9952_));
  MUX2_X1    g07126(.I0(new_n9952_), .I1(new_n9944_), .S(pi0115), .Z(new_n9953_));
  NAND2_X1   g07127(.A1(new_n9953_), .A2(new_n3154_), .ZN(new_n9954_));
  INV_X1     g07128(.I(new_n8184_), .ZN(new_n9955_));
  NAND4_X1   g07129(.A1(new_n8180_), .A2(new_n8138_), .A3(new_n9955_), .A4(new_n8474_), .ZN(new_n9956_));
  OAI21_X1   g07130(.A1(new_n9946_), .A2(new_n3172_), .B(new_n3177_), .ZN(new_n9957_));
  NAND2_X1   g07131(.A1(new_n9957_), .A2(new_n9933_), .ZN(new_n9958_));
  AOI21_X1   g07132(.A1(new_n8474_), .A2(new_n9945_), .B(new_n9958_), .ZN(new_n9959_));
  NAND2_X1   g07133(.A1(new_n8178_), .A2(pi0228), .ZN(new_n9960_));
  OAI21_X1   g07134(.A1(new_n2621_), .A2(new_n9946_), .B(new_n8535_), .ZN(new_n9961_));
  NOR2_X1    g07135(.A1(new_n2621_), .A2(pi0115), .ZN(new_n9962_));
  NAND4_X1   g07136(.A1(new_n8204_), .A2(new_n9945_), .A3(new_n9961_), .A4(new_n9962_), .ZN(new_n9963_));
  NOR2_X1    g07137(.A1(new_n2622_), .A2(pi0075), .ZN(new_n9964_));
  OAI21_X1   g07138(.A1(new_n9960_), .A2(new_n9963_), .B(new_n9964_), .ZN(new_n9965_));
  AOI21_X1   g07139(.A1(new_n9956_), .A2(new_n9959_), .B(new_n9965_), .ZN(new_n9966_));
  AOI22_X1   g07140(.A1(new_n9954_), .A2(new_n9966_), .B1(new_n9949_), .B2(new_n9950_), .ZN(new_n9967_));
  MUX2_X1    g07141(.I0(new_n9967_), .I1(new_n9946_), .S(new_n6967_), .Z(po0272));
  NAND2_X1   g07142(.A1(new_n3154_), .A2(new_n2861_), .ZN(new_n9969_));
  NOR2_X1    g07143(.A1(new_n9969_), .A2(new_n8125_), .ZN(new_n9970_));
  AOI21_X1   g07144(.A1(new_n2861_), .A2(pi0115), .B(new_n8026_), .ZN(new_n9971_));
  NAND2_X1   g07145(.A1(new_n8294_), .A2(pi0115), .ZN(new_n9972_));
  NOR4_X1    g07146(.A1(new_n8182_), .A2(pi0052), .A3(pi0115), .A4(new_n8472_), .ZN(new_n9973_));
  AOI21_X1   g07147(.A1(new_n9973_), .A2(new_n5994_), .B(new_n9926_), .ZN(new_n9974_));
  AOI21_X1   g07148(.A1(new_n9972_), .A2(new_n9974_), .B(new_n9971_), .ZN(new_n9975_));
  NOR3_X1    g07149(.A1(new_n3207_), .A2(new_n8125_), .A3(new_n9969_), .ZN(new_n9976_));
  OAI21_X1   g07150(.A1(new_n9976_), .A2(new_n2628_), .B(new_n2629_), .ZN(new_n9977_));
  NOR2_X1    g07151(.A1(new_n9975_), .A2(new_n9977_), .ZN(new_n9978_));
  AOI21_X1   g07152(.A1(new_n8266_), .A2(new_n8125_), .B(pi0039), .ZN(new_n9979_));
  OAI21_X1   g07153(.A1(new_n8257_), .A2(new_n8125_), .B(new_n9979_), .ZN(new_n9980_));
  OR3_X2     g07154(.A1(new_n9973_), .A2(pi0115), .A3(new_n8026_), .Z(new_n9981_));
  NOR2_X1    g07155(.A1(new_n9971_), .A2(pi0039), .ZN(new_n9982_));
  OAI21_X1   g07156(.A1(new_n8179_), .A2(new_n9981_), .B(new_n9982_), .ZN(new_n9983_));
  INV_X1     g07157(.I(new_n8203_), .ZN(new_n9985_));
  OAI21_X1   g07158(.A1(new_n8125_), .A2(new_n9969_), .B(new_n2622_), .ZN(new_n9987_));
  NOR4_X1    g07159(.A1(new_n9970_), .A2(new_n2535_), .A3(pi0038), .A4(pi0100), .ZN(new_n9988_));
  OAI21_X1   g07160(.A1(new_n8535_), .A2(new_n9987_), .B(new_n9988_), .ZN(new_n9989_));
  AOI21_X1   g07161(.A1(new_n9983_), .A2(new_n5158_), .B(new_n9989_), .ZN(new_n9990_));
  AOI21_X1   g07162(.A1(new_n9980_), .A2(new_n9990_), .B(new_n9978_), .ZN(new_n9991_));
  MUX2_X1    g07163(.I0(new_n9991_), .I1(new_n9970_), .S(new_n6967_), .Z(po0273));
  INV_X1     g07164(.I(new_n8110_), .ZN(new_n9993_));
  NOR2_X1    g07165(.A1(new_n9993_), .A2(pi0039), .ZN(new_n9994_));
  AOI21_X1   g07166(.A1(new_n8118_), .A2(pi0116), .B(new_n2921_), .ZN(new_n9995_));
  NOR3_X1    g07167(.A1(new_n8133_), .A2(pi0116), .A3(new_n2922_), .ZN(new_n9996_));
  NOR3_X1    g07168(.A1(new_n9996_), .A2(new_n8143_), .A3(new_n9995_), .ZN(new_n9997_));
  NAND3_X1   g07169(.A1(new_n8455_), .A2(new_n2523_), .A3(new_n2922_), .ZN(new_n9998_));
  NAND2_X1   g07170(.A1(new_n8153_), .A2(new_n9776_), .ZN(new_n9999_));
  AOI21_X1   g07171(.A1(new_n8149_), .A2(pi0116), .B(new_n9999_), .ZN(new_n10000_));
  OAI21_X1   g07172(.A1(new_n9997_), .A2(new_n9998_), .B(new_n10000_), .ZN(new_n10001_));
  INV_X1     g07173(.I(new_n9994_), .ZN(new_n10008_));
  NOR2_X1    g07174(.A1(pi0038), .A2(pi0100), .ZN(new_n10010_));
  OAI21_X1   g07175(.A1(new_n8201_), .A2(pi0113), .B(new_n8110_), .ZN(new_n10011_));
  NAND2_X1   g07176(.A1(new_n10011_), .A2(new_n9985_), .ZN(new_n10012_));
  OAI21_X1   g07177(.A1(new_n10008_), .A2(new_n3172_), .B(pi0100), .ZN(new_n10013_));
  AOI21_X1   g07178(.A1(new_n10012_), .A2(new_n3172_), .B(new_n10013_), .ZN(new_n10014_));
  NOR2_X1    g07179(.A1(new_n10008_), .A2(new_n3173_), .ZN(new_n10015_));
  OAI21_X1   g07180(.A1(new_n10014_), .A2(new_n10015_), .B(new_n8535_), .ZN(new_n10016_));
  NOR2_X1    g07181(.A1(new_n8218_), .A2(pi0113), .ZN(new_n10017_));
  OAI22_X1   g07182(.A1(new_n10017_), .A2(new_n9993_), .B1(new_n6435_), .B2(new_n8183_), .ZN(new_n10018_));
  AOI22_X1   g07183(.A1(new_n10018_), .A2(new_n9927_), .B1(new_n9926_), .B2(new_n8110_), .ZN(new_n10019_));
  NOR2_X1    g07184(.A1(new_n8342_), .A2(new_n9994_), .ZN(new_n10020_));
  OAI21_X1   g07185(.A1(new_n10019_), .A2(new_n2629_), .B(new_n10020_), .ZN(new_n10021_));
  NAND3_X1   g07186(.A1(new_n10021_), .A2(new_n2628_), .A3(new_n10016_), .ZN(new_n10022_));
  AOI21_X1   g07187(.A1(new_n10001_), .A2(new_n10010_), .B(new_n10022_), .ZN(new_n10023_));
  MUX2_X1    g07188(.I0(new_n10023_), .I1(new_n9994_), .S(new_n6967_), .Z(po0274));
  NOR2_X1    g07189(.A1(new_n5900_), .A2(pi0039), .ZN(new_n10025_));
  OAI21_X1   g07190(.A1(new_n3524_), .A2(pi0100), .B(new_n10025_), .ZN(new_n10026_));
  NOR3_X1    g07191(.A1(new_n3379_), .A2(pi0100), .A3(new_n10025_), .ZN(new_n10027_));
  NOR2_X1    g07192(.A1(new_n10027_), .A2(pi0038), .ZN(new_n10028_));
  NAND2_X1   g07193(.A1(new_n3177_), .A2(pi0075), .ZN(new_n10029_));
  AOI21_X1   g07194(.A1(new_n10028_), .A2(new_n10026_), .B(new_n10029_), .ZN(new_n10030_));
  NOR3_X1    g07195(.A1(new_n5880_), .A2(pi0054), .A3(pi0074), .ZN(new_n10031_));
  OAI21_X1   g07196(.A1(new_n10030_), .A2(pi0092), .B(new_n10031_), .ZN(new_n10032_));
  AOI21_X1   g07197(.A1(new_n10032_), .A2(new_n3227_), .B(new_n5888_), .ZN(new_n10033_));
  NOR3_X1    g07198(.A1(new_n10032_), .A2(pi0055), .A3(new_n5887_), .ZN(new_n10034_));
  NOR3_X1    g07199(.A1(new_n10034_), .A2(new_n10033_), .A3(pi0056), .ZN(new_n10035_));
  OAI21_X1   g07200(.A1(new_n10035_), .A2(new_n5057_), .B(new_n5203_), .ZN(po0275));
  NAND2_X1   g07201(.A1(new_n7049_), .A2(pi0165), .ZN(new_n10037_));
  INV_X1     g07202(.I(pi0150), .ZN(new_n10038_));
  NOR2_X1    g07203(.A1(new_n10038_), .A2(pi0163), .ZN(new_n10039_));
  NAND4_X1   g07204(.A1(new_n8830_), .A2(new_n5108_), .A3(new_n8827_), .A4(new_n10039_), .ZN(new_n10040_));
  NOR2_X1    g07205(.A1(new_n5109_), .A2(new_n8826_), .ZN(new_n10041_));
  OAI21_X1   g07206(.A1(new_n8853_), .A2(new_n10041_), .B(new_n10038_), .ZN(new_n10042_));
  NAND3_X1   g07207(.A1(new_n10042_), .A2(pi0232), .A3(new_n10040_), .ZN(new_n10043_));
  INV_X1     g07208(.I(new_n10043_), .ZN(new_n10044_));
  OAI21_X1   g07209(.A1(new_n10044_), .A2(new_n7041_), .B(new_n3202_), .ZN(new_n10045_));
  NAND3_X1   g07210(.A1(new_n10044_), .A2(pi0074), .A3(new_n7048_), .ZN(new_n10046_));
  AOI22_X1   g07211(.A1(new_n10045_), .A2(new_n10046_), .B1(new_n3405_), .B2(new_n10037_), .ZN(new_n10047_));
  INV_X1     g07212(.I(pi0143), .ZN(new_n10048_));
  OAI21_X1   g07213(.A1(new_n10048_), .A2(pi0165), .B(pi0299), .ZN(new_n10049_));
  NOR2_X1    g07214(.A1(new_n5989_), .A2(new_n10049_), .ZN(new_n10050_));
  INV_X1     g07215(.I(new_n10050_), .ZN(new_n10051_));
  NOR3_X1    g07216(.A1(new_n10051_), .A2(pi0054), .A3(new_n7041_), .ZN(new_n10052_));
  NOR4_X1    g07217(.A1(new_n7284_), .A2(pi0038), .A3(new_n10048_), .A4(pi0165), .ZN(new_n10054_));
  NOR2_X1    g07218(.A1(new_n10054_), .A2(new_n3206_), .ZN(new_n10055_));
  INV_X1     g07219(.I(pi0173), .ZN(new_n10056_));
  INV_X1     g07220(.I(new_n7403_), .ZN(new_n10057_));
  NAND3_X1   g07221(.A1(new_n7506_), .A2(new_n5108_), .A3(new_n10057_), .ZN(new_n10058_));
  OAI21_X1   g07222(.A1(new_n7506_), .A2(new_n5109_), .B(new_n7403_), .ZN(new_n10059_));
  AOI21_X1   g07223(.A1(new_n10059_), .A2(new_n10058_), .B(new_n10056_), .ZN(new_n10060_));
  NOR2_X1    g07224(.A1(new_n10057_), .A2(new_n5108_), .ZN(new_n10061_));
  OAI21_X1   g07225(.A1(new_n7565_), .A2(new_n10061_), .B(new_n10056_), .ZN(new_n10062_));
  NAND2_X1   g07226(.A1(new_n10062_), .A2(pi0185), .ZN(new_n10063_));
  NOR2_X1    g07227(.A1(new_n7403_), .A2(new_n5108_), .ZN(new_n10064_));
  NOR2_X1    g07228(.A1(new_n10064_), .A2(new_n7427_), .ZN(new_n10065_));
  INV_X1     g07229(.I(pi0185), .ZN(new_n10066_));
  NOR2_X1    g07230(.A1(new_n10056_), .A2(new_n10066_), .ZN(new_n10067_));
  NAND2_X1   g07231(.A1(new_n10065_), .A2(new_n10067_), .ZN(new_n10068_));
  OAI21_X1   g07232(.A1(new_n10063_), .A2(new_n10060_), .B(new_n10068_), .ZN(new_n10069_));
  OAI21_X1   g07233(.A1(new_n7514_), .A2(new_n7518_), .B(pi0173), .ZN(new_n10070_));
  NOR2_X1    g07234(.A1(new_n10070_), .A2(new_n5109_), .ZN(new_n10071_));
  OAI21_X1   g07235(.A1(new_n10057_), .A2(new_n5108_), .B(pi0185), .ZN(new_n10072_));
  NOR2_X1    g07236(.A1(new_n7420_), .A2(new_n10064_), .ZN(new_n10073_));
  INV_X1     g07237(.I(new_n10073_), .ZN(new_n10074_));
  AOI21_X1   g07238(.A1(new_n10056_), .A2(new_n10057_), .B(new_n10074_), .ZN(new_n10075_));
  NOR3_X1    g07239(.A1(new_n10073_), .A2(pi0173), .A3(new_n10057_), .ZN(new_n10076_));
  NOR4_X1    g07240(.A1(new_n10075_), .A2(pi0185), .A3(pi0190), .A4(new_n10076_), .ZN(new_n10077_));
  OAI21_X1   g07241(.A1(new_n10071_), .A2(new_n10072_), .B(new_n10077_), .ZN(new_n10078_));
  AOI21_X1   g07242(.A1(new_n10078_), .A2(new_n2587_), .B(pi0190), .ZN(new_n10079_));
  INV_X1     g07243(.I(new_n7499_), .ZN(new_n10080_));
  AOI21_X1   g07244(.A1(new_n4413_), .A2(new_n10080_), .B(new_n7485_), .ZN(new_n10081_));
  NAND3_X1   g07245(.A1(new_n7485_), .A2(new_n4413_), .A3(new_n7499_), .ZN(new_n10082_));
  NOR4_X1    g07246(.A1(new_n7454_), .A2(pi0151), .A3(pi0168), .A4(new_n10061_), .ZN(new_n10083_));
  NAND2_X1   g07247(.A1(new_n10082_), .A2(new_n10083_), .ZN(new_n10084_));
  NAND2_X1   g07248(.A1(new_n7406_), .A2(new_n5108_), .ZN(new_n10085_));
  NOR3_X1    g07249(.A1(new_n10061_), .A2(new_n3417_), .A3(new_n4413_), .ZN(new_n10086_));
  NOR2_X1    g07250(.A1(new_n5109_), .A2(new_n4413_), .ZN(new_n10088_));
  INV_X1     g07251(.I(new_n10088_), .ZN(new_n10089_));
  NAND3_X1   g07252(.A1(new_n5987_), .A2(new_n2587_), .A3(pi0150), .ZN(new_n10092_));
  AOI21_X1   g07253(.A1(new_n10085_), .A2(new_n10086_), .B(new_n10092_), .ZN(new_n10093_));
  OAI21_X1   g07254(.A1(new_n10084_), .A2(new_n10081_), .B(new_n10093_), .ZN(new_n10094_));
  AOI21_X1   g07255(.A1(new_n10069_), .A2(new_n10079_), .B(new_n10094_), .ZN(new_n10095_));
  INV_X1     g07256(.I(pi0190), .ZN(new_n10096_));
  NAND2_X1   g07257(.A1(new_n7611_), .A2(pi0178), .ZN(new_n10097_));
  NAND2_X1   g07258(.A1(new_n10097_), .A2(new_n10096_), .ZN(new_n10098_));
  NOR2_X1    g07259(.A1(new_n7635_), .A2(new_n4413_), .ZN(new_n10099_));
  NAND2_X1   g07260(.A1(new_n7629_), .A2(pi0157), .ZN(new_n10100_));
  NAND4_X1   g07261(.A1(new_n10100_), .A2(new_n6445_), .A3(new_n5108_), .A4(new_n7170_), .ZN(new_n10101_));
  OAI21_X1   g07262(.A1(new_n10101_), .A2(new_n10099_), .B(pi0299), .ZN(new_n10102_));
  AOI21_X1   g07263(.A1(new_n7345_), .A2(new_n2587_), .B(new_n7086_), .ZN(new_n10103_));
  AOI22_X1   g07264(.A1(new_n10102_), .A2(new_n10103_), .B1(new_n10098_), .B2(new_n2587_), .ZN(new_n10104_));
  OAI21_X1   g07265(.A1(new_n6460_), .A2(new_n7086_), .B(new_n7153_), .ZN(new_n10105_));
  NOR2_X1    g07266(.A1(new_n10096_), .A2(pi0299), .ZN(new_n10106_));
  INV_X1     g07267(.I(new_n10106_), .ZN(new_n10107_));
  OAI21_X1   g07268(.A1(new_n7605_), .A2(new_n10107_), .B(pi0178), .ZN(new_n10108_));
  NOR2_X1    g07269(.A1(new_n10108_), .A2(new_n10105_), .ZN(new_n10109_));
  NAND2_X1   g07270(.A1(new_n7607_), .A2(new_n10109_), .ZN(new_n10110_));
  AOI21_X1   g07271(.A1(new_n7086_), .A2(new_n5987_), .B(new_n3154_), .ZN(new_n10111_));
  NOR4_X1    g07272(.A1(new_n10105_), .A2(pi0178), .A3(pi0232), .A4(new_n10111_), .ZN(new_n10112_));
  NAND3_X1   g07273(.A1(new_n10110_), .A2(new_n7624_), .A3(new_n10112_), .ZN(new_n10113_));
  AOI21_X1   g07274(.A1(new_n7403_), .A2(new_n5987_), .B(new_n2545_), .ZN(new_n10114_));
  OAI21_X1   g07275(.A1(new_n10113_), .A2(new_n10104_), .B(new_n10114_), .ZN(new_n10115_));
  OAI21_X1   g07276(.A1(new_n10095_), .A2(new_n10115_), .B(new_n10055_), .ZN(new_n10116_));
  INV_X1     g07277(.I(pi0157), .ZN(new_n10117_));
  MUX2_X1    g07278(.I0(new_n7345_), .I1(new_n10117_), .S(pi0299), .Z(new_n10118_));
  NOR2_X1    g07279(.A1(new_n5989_), .A2(new_n10118_), .ZN(new_n10119_));
  AOI21_X1   g07280(.A1(new_n10051_), .A2(pi0038), .B(pi0100), .ZN(new_n10120_));
  INV_X1     g07281(.I(new_n10120_), .ZN(new_n10121_));
  NAND4_X1   g07282(.A1(new_n7119_), .A2(new_n7144_), .A3(new_n10119_), .A4(new_n10121_), .ZN(new_n10122_));
  AOI21_X1   g07283(.A1(new_n10122_), .A2(new_n3173_), .B(new_n7124_), .ZN(new_n10123_));
  NAND3_X1   g07284(.A1(new_n10050_), .A2(new_n3173_), .A3(new_n7290_), .ZN(new_n10124_));
  NOR2_X1    g07285(.A1(new_n10124_), .A2(new_n7143_), .ZN(new_n10125_));
  NOR4_X1    g07286(.A1(new_n10123_), .A2(new_n3209_), .A3(new_n7048_), .A4(new_n10125_), .ZN(new_n10126_));
  AOI21_X1   g07287(.A1(new_n10116_), .A2(new_n10126_), .B(pi0054), .ZN(new_n10127_));
  OAI21_X1   g07288(.A1(new_n10127_), .A2(new_n10052_), .B(new_n3202_), .ZN(new_n10128_));
  NOR2_X1    g07289(.A1(new_n10043_), .A2(new_n7041_), .ZN(new_n10129_));
  NOR2_X1    g07290(.A1(pi0038), .A2(pi0054), .ZN(new_n10130_));
  NAND3_X1   g07291(.A1(new_n5988_), .A2(pi0165), .A3(new_n10130_), .ZN(new_n10131_));
  NOR2_X1    g07292(.A1(new_n5989_), .A2(new_n10038_), .ZN(new_n10133_));
  NOR2_X1    g07293(.A1(new_n2533_), .A2(pi0055), .ZN(new_n10137_));
  NAND2_X1   g07294(.A1(new_n10043_), .A2(new_n7041_), .ZN(new_n10138_));
  NOR2_X1    g07295(.A1(new_n10131_), .A2(new_n7048_), .ZN(new_n10139_));
  NOR2_X1    g07296(.A1(new_n10139_), .A2(pi0074), .ZN(new_n10140_));
  NAND2_X1   g07297(.A1(new_n10138_), .A2(new_n10140_), .ZN(new_n10141_));
  NOR2_X1    g07298(.A1(new_n10129_), .A2(new_n3202_), .ZN(new_n10142_));
  NOR2_X1    g07299(.A1(new_n2533_), .A2(new_n2571_), .ZN(new_n10143_));
  OAI21_X1   g07300(.A1(new_n10142_), .A2(new_n10141_), .B(new_n10143_), .ZN(new_n10144_));
  AOI22_X1   g07301(.A1(new_n10128_), .A2(new_n10137_), .B1(new_n7682_), .B2(new_n10144_), .ZN(new_n10145_));
  NOR2_X1    g07302(.A1(new_n10145_), .A2(new_n10047_), .ZN(new_n10146_));
  INV_X1     g07303(.I(new_n10146_), .ZN(new_n10147_));
  INV_X1     g07304(.I(new_n10144_), .ZN(new_n10148_));
  OAI21_X1   g07305(.A1(new_n7235_), .A2(new_n7251_), .B(pi0173), .ZN(new_n10149_));
  OAI21_X1   g07306(.A1(new_n10149_), .A2(new_n2515_), .B(new_n10096_), .ZN(new_n10150_));
  NOR3_X1    g07307(.A1(new_n10096_), .A2(pi0173), .A3(pi0185), .ZN(new_n10151_));
  AOI21_X1   g07308(.A1(new_n7205_), .A2(new_n10151_), .B(new_n5108_), .ZN(new_n10152_));
  NOR3_X1    g07309(.A1(new_n7266_), .A2(new_n7224_), .A3(pi0173), .ZN(new_n10153_));
  INV_X1     g07310(.I(new_n10153_), .ZN(new_n10154_));
  NOR2_X1    g07311(.A1(pi0185), .A2(pi0190), .ZN(new_n10156_));
  AOI22_X1   g07312(.A1(new_n10154_), .A2(new_n10156_), .B1(new_n10150_), .B2(new_n10152_), .ZN(new_n10157_));
  NOR2_X1    g07313(.A1(new_n7230_), .A2(new_n5108_), .ZN(new_n10158_));
  OAI21_X1   g07314(.A1(new_n10157_), .A2(pi0299), .B(new_n10158_), .ZN(new_n10159_));
  NOR3_X1    g07315(.A1(new_n7240_), .A2(new_n7224_), .A3(pi0151), .ZN(new_n10160_));
  INV_X1     g07316(.I(new_n10160_), .ZN(new_n10161_));
  NOR3_X1    g07317(.A1(new_n7190_), .A2(pi0151), .A3(new_n10088_), .ZN(new_n10162_));
  AOI21_X1   g07318(.A1(new_n9065_), .A2(new_n10162_), .B(pi0168), .ZN(new_n10163_));
  AOI21_X1   g07319(.A1(new_n10161_), .A2(new_n10163_), .B(pi0150), .ZN(new_n10164_));
  NOR3_X1    g07320(.A1(new_n7204_), .A2(new_n7234_), .A3(new_n4413_), .ZN(new_n10165_));
  AOI21_X1   g07321(.A1(pi0168), .A2(new_n7204_), .B(new_n7235_), .ZN(new_n10166_));
  OAI21_X1   g07322(.A1(new_n10166_), .A2(new_n10165_), .B(new_n3417_), .ZN(new_n10167_));
  NOR3_X1    g07323(.A1(new_n7252_), .A2(new_n3417_), .A3(pi0168), .ZN(new_n10168_));
  NOR4_X1    g07324(.A1(new_n10168_), .A2(pi0040), .A3(new_n10038_), .A4(new_n7196_), .ZN(new_n10169_));
  AOI21_X1   g07325(.A1(new_n10167_), .A2(new_n10169_), .B(new_n5108_), .ZN(new_n10170_));
  OAI21_X1   g07326(.A1(new_n7225_), .A2(new_n9051_), .B(new_n10170_), .ZN(new_n10171_));
  OAI21_X1   g07327(.A1(new_n10164_), .A2(new_n10171_), .B(new_n2587_), .ZN(new_n10172_));
  AOI21_X1   g07328(.A1(new_n10159_), .A2(new_n10172_), .B(pi0232), .ZN(new_n10173_));
  NAND2_X1   g07329(.A1(new_n5145_), .A2(new_n7345_), .ZN(new_n10174_));
  NOR2_X1    g07330(.A1(new_n5143_), .A2(new_n7345_), .ZN(new_n10175_));
  AOI22_X1   g07331(.A1(new_n7162_), .A2(new_n10175_), .B1(new_n10096_), .B2(new_n10174_), .ZN(new_n10176_));
  NAND2_X1   g07332(.A1(new_n5144_), .A2(new_n7345_), .ZN(new_n10177_));
  OAI21_X1   g07333(.A1(new_n6048_), .A2(new_n10177_), .B(new_n6548_), .ZN(new_n10178_));
  AOI21_X1   g07334(.A1(new_n10178_), .A2(pi0190), .B(new_n10176_), .ZN(new_n10179_));
  INV_X1     g07335(.I(new_n9700_), .ZN(new_n10180_));
  NOR3_X1    g07336(.A1(new_n7166_), .A2(pi0157), .A3(pi0168), .ZN(new_n10181_));
  AOI21_X1   g07337(.A1(new_n7168_), .A2(new_n10181_), .B(new_n5143_), .ZN(new_n10182_));
  NOR2_X1    g07338(.A1(new_n9702_), .A2(pi0232), .ZN(new_n10183_));
  OAI21_X1   g07339(.A1(new_n10182_), .A2(new_n10180_), .B(new_n10183_), .ZN(new_n10184_));
  OAI21_X1   g07340(.A1(new_n5133_), .A2(new_n9700_), .B(new_n5987_), .ZN(new_n10185_));
  NAND3_X1   g07341(.A1(new_n5146_), .A2(new_n2587_), .A3(new_n7153_), .ZN(new_n10186_));
  AOI21_X1   g07342(.A1(new_n10185_), .A2(new_n10186_), .B(new_n3154_), .ZN(new_n10187_));
  OAI21_X1   g07343(.A1(new_n10184_), .A2(new_n10179_), .B(new_n10187_), .ZN(new_n10188_));
  NOR2_X1    g07344(.A1(new_n7228_), .A2(new_n5081_), .ZN(new_n10189_));
  OAI21_X1   g07345(.A1(new_n7225_), .A2(pi0232), .B(new_n10189_), .ZN(new_n10190_));
  NAND3_X1   g07346(.A1(new_n10188_), .A2(new_n3154_), .A3(new_n10190_), .ZN(new_n10191_));
  NOR2_X1    g07347(.A1(new_n10055_), .A2(pi0038), .ZN(new_n10192_));
  OAI21_X1   g07348(.A1(new_n10173_), .A2(new_n10191_), .B(new_n10192_), .ZN(new_n10193_));
  NAND2_X1   g07349(.A1(new_n10124_), .A2(new_n3173_), .ZN(new_n10194_));
  INV_X1     g07350(.I(new_n10194_), .ZN(new_n10195_));
  AOI21_X1   g07351(.A1(new_n10193_), .A2(new_n10195_), .B(new_n3209_), .ZN(new_n10196_));
  INV_X1     g07352(.I(new_n10196_), .ZN(new_n10197_));
  NOR4_X1    g07353(.A1(new_n2491_), .A2(pi0087), .A3(new_n2545_), .A4(new_n10119_), .ZN(new_n10198_));
  OAI21_X1   g07354(.A1(new_n10198_), .A2(new_n10121_), .B(new_n3173_), .ZN(new_n10199_));
  AOI21_X1   g07355(.A1(new_n10199_), .A2(new_n7123_), .B(new_n7362_), .ZN(new_n10200_));
  AOI21_X1   g07356(.A1(new_n10197_), .A2(new_n10200_), .B(new_n10052_), .ZN(new_n10201_));
  NOR2_X1    g07357(.A1(new_n2533_), .A2(pi0055), .ZN(new_n10207_));
  OAI21_X1   g07358(.A1(new_n10201_), .A2(pi0074), .B(new_n10207_), .ZN(new_n10208_));
  AOI21_X1   g07359(.A1(new_n10208_), .A2(new_n10148_), .B(new_n10047_), .ZN(new_n10209_));
  OAI21_X1   g07360(.A1(pi0118), .A2(new_n10209_), .B(new_n10147_), .ZN(new_n10210_));
  NAND3_X1   g07361(.A1(new_n10146_), .A2(new_n7748_), .A3(new_n10209_), .ZN(new_n10211_));
  NOR2_X1    g07362(.A1(new_n9125_), .A2(pi0079), .ZN(new_n10212_));
  INV_X1     g07363(.I(new_n10212_), .ZN(new_n10213_));
  NAND2_X1   g07364(.A1(new_n7316_), .A2(new_n7748_), .ZN(new_n10214_));
  INV_X1     g07365(.I(new_n10209_), .ZN(new_n10215_));
  AOI21_X1   g07366(.A1(new_n10215_), .A2(new_n10214_), .B(new_n10212_), .ZN(new_n10216_));
  OAI21_X1   g07367(.A1(new_n10147_), .A2(new_n10214_), .B(new_n10216_), .ZN(new_n10217_));
  NAND4_X1   g07368(.A1(new_n10210_), .A2(new_n10211_), .A3(new_n10217_), .A4(new_n10213_), .ZN(po0276));
  NAND2_X1   g07369(.A1(pi0128), .A2(pi0228), .ZN(new_n10219_));
  INV_X1     g07370(.I(new_n10219_), .ZN(new_n10220_));
  NOR3_X1    g07371(.A1(new_n5910_), .A2(new_n3203_), .A3(new_n10220_), .ZN(new_n10221_));
  NOR4_X1    g07372(.A1(new_n3311_), .A2(pi0087), .A3(pi0100), .A4(new_n2545_), .ZN(new_n10222_));
  OAI21_X1   g07373(.A1(new_n10222_), .A2(new_n10220_), .B(pi0075), .ZN(new_n10223_));
  NAND2_X1   g07374(.A1(new_n10223_), .A2(new_n3203_), .ZN(new_n10224_));
  NOR2_X1    g07375(.A1(new_n2523_), .A2(pi0128), .ZN(new_n10225_));
  NAND2_X1   g07376(.A1(new_n2669_), .A2(pi0093), .ZN(new_n10226_));
  OR3_X2     g07377(.A1(new_n5278_), .A2(new_n2964_), .A3(new_n8819_), .Z(new_n10227_));
  INV_X1     g07378(.I(new_n2685_), .ZN(new_n10228_));
  AOI21_X1   g07379(.A1(new_n10228_), .A2(new_n7816_), .B(new_n2822_), .ZN(new_n10229_));
  MUX2_X1    g07380(.I0(new_n5346_), .I1(new_n5442_), .S(new_n2587_), .Z(new_n10230_));
  NOR2_X1    g07381(.A1(new_n10230_), .A2(new_n5989_), .ZN(new_n10231_));
  NOR2_X1    g07382(.A1(new_n10231_), .A2(new_n2470_), .ZN(new_n10232_));
  NOR3_X1    g07383(.A1(new_n10230_), .A2(new_n5304_), .A3(new_n5989_), .ZN(new_n10233_));
  NAND4_X1   g07384(.A1(new_n2964_), .A2(new_n2465_), .A3(new_n2680_), .A4(new_n5062_), .ZN(new_n10234_));
  NOR4_X1    g07385(.A1(new_n10232_), .A2(new_n2689_), .A3(new_n10233_), .A4(new_n10234_), .ZN(new_n10235_));
  OAI21_X1   g07386(.A1(new_n5284_), .A2(new_n10231_), .B(new_n10235_), .ZN(new_n10236_));
  AOI21_X1   g07387(.A1(new_n10229_), .A2(new_n8819_), .B(new_n10236_), .ZN(new_n10237_));
  AOI21_X1   g07388(.A1(new_n10227_), .A2(new_n10237_), .B(new_n2660_), .ZN(new_n10238_));
  OAI21_X1   g07389(.A1(new_n10238_), .A2(new_n2844_), .B(new_n2666_), .ZN(new_n10239_));
  NAND2_X1   g07390(.A1(new_n8589_), .A2(new_n3154_), .ZN(new_n10240_));
  AOI21_X1   g07391(.A1(new_n10239_), .A2(new_n10226_), .B(new_n10240_), .ZN(new_n10241_));
  NAND3_X1   g07392(.A1(new_n6054_), .A2(new_n3285_), .A3(new_n4899_), .ZN(new_n10242_));
  NOR2_X1    g07393(.A1(new_n3294_), .A2(new_n2614_), .ZN(new_n10243_));
  NAND2_X1   g07394(.A1(new_n6049_), .A2(new_n10243_), .ZN(new_n10244_));
  AND3_X2    g07395(.A1(new_n10242_), .A2(pi0039), .A3(new_n10244_), .Z(new_n10245_));
  OAI21_X1   g07396(.A1(new_n10245_), .A2(new_n10241_), .B(new_n3172_), .ZN(new_n10246_));
  AOI21_X1   g07397(.A1(new_n10246_), .A2(new_n2523_), .B(new_n10225_), .ZN(new_n10247_));
  NAND2_X1   g07398(.A1(new_n3310_), .A2(new_n2544_), .ZN(new_n10248_));
  NAND2_X1   g07399(.A1(new_n10248_), .A2(new_n10219_), .ZN(new_n10249_));
  MUX2_X1    g07400(.I0(new_n10249_), .I1(new_n10247_), .S(new_n3173_), .Z(new_n10250_));
  AOI21_X1   g07401(.A1(new_n10219_), .A2(pi0087), .B(pi0075), .ZN(new_n10251_));
  OAI21_X1   g07402(.A1(new_n10250_), .A2(pi0087), .B(new_n10251_), .ZN(new_n10252_));
  AOI21_X1   g07403(.A1(new_n10252_), .A2(new_n10224_), .B(new_n10221_), .ZN(new_n10253_));
  MUX2_X1    g07404(.I0(new_n10253_), .I1(new_n10220_), .S(new_n7823_), .Z(po0277));
  NAND3_X1   g07405(.A1(new_n6958_), .A2(new_n9632_), .A3(pi0818), .ZN(new_n10255_));
  INV_X1     g07406(.I(new_n10255_), .ZN(new_n10256_));
  NOR4_X1    g07407(.A1(new_n9432_), .A2(pi0120), .A3(pi1091), .A4(pi1093), .ZN(new_n10257_));
  AOI21_X1   g07408(.A1(new_n6429_), .A2(pi0120), .B(new_n10257_), .ZN(new_n10258_));
  AOI21_X1   g07409(.A1(new_n2918_), .A2(new_n6427_), .B(new_n6437_), .ZN(new_n10259_));
  INV_X1     g07410(.I(new_n10259_), .ZN(new_n10260_));
  AOI21_X1   g07411(.A1(new_n10260_), .A2(pi0120), .B(new_n5990_), .ZN(new_n10261_));
  INV_X1     g07412(.I(new_n10261_), .ZN(new_n10262_));
  AND2_X2    g07413(.A1(new_n5997_), .A2(new_n10257_), .Z(new_n10263_));
  INV_X1     g07414(.I(new_n10258_), .ZN(new_n10264_));
  OAI22_X1   g07415(.A1(new_n10262_), .A2(new_n10263_), .B1(new_n8334_), .B2(new_n10264_), .ZN(new_n10265_));
  NOR4_X1    g07416(.A1(new_n10265_), .A2(pi0075), .A3(new_n2629_), .A4(new_n10258_), .ZN(new_n10266_));
  INV_X1     g07417(.I(pi0120), .ZN(new_n10267_));
  INV_X1     g07418(.I(new_n6014_), .ZN(new_n10268_));
  NAND2_X1   g07419(.A1(new_n10268_), .A2(new_n6429_), .ZN(new_n10269_));
  NAND2_X1   g07420(.A1(new_n6012_), .A2(new_n5996_), .ZN(new_n10270_));
  NAND3_X1   g07421(.A1(new_n10269_), .A2(new_n10267_), .A3(new_n10270_), .ZN(new_n10271_));
  NAND3_X1   g07422(.A1(new_n10268_), .A2(new_n10267_), .A3(pi1093), .ZN(new_n10272_));
  NAND2_X1   g07423(.A1(new_n6481_), .A2(new_n2544_), .ZN(new_n10273_));
  NAND3_X1   g07424(.A1(new_n10273_), .A2(new_n10264_), .A3(new_n3173_), .ZN(new_n10274_));
  AOI21_X1   g07425(.A1(new_n10271_), .A2(new_n10272_), .B(new_n10274_), .ZN(new_n10275_));
  NAND2_X1   g07426(.A1(new_n10258_), .A2(new_n6559_), .ZN(new_n10276_));
  NAND3_X1   g07427(.A1(new_n10258_), .A2(new_n2587_), .A3(new_n6453_), .ZN(new_n10277_));
  NAND4_X1   g07428(.A1(new_n10277_), .A2(new_n10276_), .A3(pi0039), .A4(new_n2587_), .ZN(new_n10278_));
  NOR2_X1    g07429(.A1(new_n5974_), .A2(new_n5977_), .ZN(new_n10279_));
  NOR2_X1    g07430(.A1(new_n10279_), .A2(pi1093), .ZN(new_n10280_));
  AOI21_X1   g07431(.A1(new_n10280_), .A2(pi0120), .B(pi0039), .ZN(new_n10281_));
  INV_X1     g07432(.I(new_n10281_), .ZN(new_n10282_));
  AND4_X2    g07433(.A1(new_n6029_), .A2(new_n7947_), .A3(new_n2958_), .A4(new_n6027_), .Z(new_n10283_));
  NOR2_X1    g07434(.A1(new_n5182_), .A2(pi0122), .ZN(new_n10284_));
  NOR2_X1    g07435(.A1(new_n6005_), .A2(pi0829), .ZN(new_n10285_));
  OAI21_X1   g07436(.A1(new_n10284_), .A2(new_n10285_), .B(new_n7935_), .ZN(new_n10286_));
  AOI21_X1   g07437(.A1(new_n10283_), .A2(new_n10286_), .B(new_n7756_), .ZN(new_n10287_));
  INV_X1     g07438(.I(new_n10287_), .ZN(new_n10288_));
  AOI21_X1   g07439(.A1(new_n7935_), .A2(new_n6004_), .B(new_n9141_), .ZN(new_n10289_));
  NAND2_X1   g07440(.A1(new_n10289_), .A2(new_n9432_), .ZN(new_n10290_));
  NAND2_X1   g07441(.A1(new_n10288_), .A2(new_n10290_), .ZN(new_n10291_));
  OAI21_X1   g07442(.A1(new_n10291_), .A2(new_n10282_), .B(new_n10278_), .ZN(new_n10292_));
  NOR2_X1    g07443(.A1(pi0120), .A2(pi1093), .ZN(new_n10293_));
  OAI21_X1   g07444(.A1(new_n6428_), .A2(new_n10293_), .B(pi0038), .ZN(new_n10294_));
  AOI22_X1   g07445(.A1(new_n10292_), .A2(new_n3172_), .B1(new_n3173_), .B2(new_n10294_), .ZN(new_n10295_));
  OAI21_X1   g07446(.A1(new_n10295_), .A2(new_n10275_), .B(new_n3177_), .ZN(new_n10296_));
  NAND4_X1   g07447(.A1(new_n2491_), .A2(pi0122), .A3(new_n6005_), .A4(new_n9141_), .ZN(new_n10297_));
  NAND4_X1   g07448(.A1(new_n10297_), .A2(new_n3197_), .A3(new_n6001_), .A4(new_n9141_), .ZN(new_n10298_));
  NAND4_X1   g07449(.A1(new_n10298_), .A2(new_n3177_), .A3(new_n3198_), .A4(new_n6428_), .ZN(new_n10299_));
  OR3_X2     g07450(.A1(new_n6009_), .A2(new_n10293_), .A3(new_n10299_), .Z(new_n10300_));
  AOI21_X1   g07451(.A1(new_n10296_), .A2(new_n10300_), .B(pi0075), .ZN(new_n10301_));
  AOI21_X1   g07452(.A1(new_n6428_), .A2(new_n5942_), .B(new_n6538_), .ZN(new_n10302_));
  INV_X1     g07453(.I(new_n10302_), .ZN(new_n10303_));
  NOR2_X1    g07454(.A1(new_n5941_), .A2(pi0120), .ZN(new_n10304_));
  AOI21_X1   g07455(.A1(new_n2924_), .A2(new_n10304_), .B(new_n10303_), .ZN(new_n10305_));
  NOR2_X1    g07456(.A1(new_n10305_), .A2(new_n5941_), .ZN(new_n10306_));
  OAI21_X1   g07457(.A1(new_n10301_), .A2(new_n10266_), .B(new_n10306_), .ZN(new_n10307_));
  INV_X1     g07458(.I(new_n10293_), .ZN(new_n10308_));
  NAND2_X1   g07459(.A1(new_n2587_), .A2(pi0039), .ZN(new_n10309_));
  NAND3_X1   g07460(.A1(new_n10293_), .A2(pi0038), .A3(pi0100), .ZN(new_n10320_));
  MUX2_X1    g07461(.I0(new_n10270_), .I1(new_n10268_), .S(pi0120), .Z(new_n10321_));
  OAI21_X1   g07462(.A1(new_n10321_), .A2(new_n10273_), .B(new_n10308_), .ZN(new_n10322_));
  AOI21_X1   g07463(.A1(new_n10322_), .A2(new_n3173_), .B(pi0087), .ZN(new_n10323_));
  AOI22_X1   g07464(.A1(new_n10323_), .A2(new_n10320_), .B1(new_n6008_), .B2(new_n10308_), .ZN(new_n10324_));
  NAND4_X1   g07465(.A1(new_n5999_), .A2(new_n2628_), .A3(new_n5942_), .A4(new_n10308_), .ZN(new_n10325_));
  AOI21_X1   g07466(.A1(new_n10304_), .A2(new_n2924_), .B(new_n6844_), .ZN(new_n10326_));
  OAI21_X1   g07467(.A1(new_n10324_), .A2(new_n10325_), .B(new_n10326_), .ZN(new_n10327_));
  AOI21_X1   g07468(.A1(new_n10307_), .A2(new_n10327_), .B(new_n10255_), .ZN(new_n10328_));
  NOR2_X1    g07469(.A1(new_n10264_), .A2(new_n6538_), .ZN(new_n10329_));
  NOR2_X1    g07470(.A1(po1038), .A2(new_n10256_), .ZN(new_n10330_));
  OAI21_X1   g07471(.A1(new_n10329_), .A2(new_n10293_), .B(new_n10330_), .ZN(new_n10331_));
  INV_X1     g07472(.I(new_n6953_), .ZN(new_n10332_));
  NAND3_X1   g07473(.A1(pi0951), .A2(pi0982), .A3(pi1092), .ZN(new_n10333_));
  NOR2_X1    g07474(.A1(new_n10333_), .A2(new_n2924_), .ZN(new_n10334_));
  NOR2_X1    g07475(.A1(new_n10334_), .A2(pi0120), .ZN(new_n10335_));
  OAI21_X1   g07476(.A1(new_n10329_), .A2(new_n10335_), .B(new_n10332_), .ZN(new_n10336_));
  NOR2_X1    g07477(.A1(new_n10331_), .A2(new_n10336_), .ZN(new_n10337_));
  INV_X1     g07478(.I(new_n10329_), .ZN(new_n10338_));
  NAND3_X1   g07479(.A1(new_n10331_), .A2(pi0120), .A3(new_n10338_), .ZN(new_n10339_));
  NAND2_X1   g07480(.A1(new_n10339_), .A2(new_n10332_), .ZN(new_n10340_));
  OAI22_X1   g07481(.A1(new_n10328_), .A2(po1038), .B1(new_n10337_), .B2(new_n10340_), .ZN(new_n10341_));
  INV_X1     g07482(.I(new_n10305_), .ZN(new_n10342_));
  NOR2_X1    g07483(.A1(new_n8334_), .A2(new_n10335_), .ZN(new_n10343_));
  OAI21_X1   g07484(.A1(new_n10335_), .A2(new_n2625_), .B(pi0075), .ZN(new_n10344_));
  AOI21_X1   g07485(.A1(new_n10343_), .A2(new_n2625_), .B(new_n10344_), .ZN(new_n10345_));
  NOR3_X1    g07486(.A1(new_n10287_), .A2(new_n10280_), .A3(new_n10289_), .ZN(new_n10346_));
  NAND2_X1   g07487(.A1(new_n10346_), .A2(pi0120), .ZN(new_n10347_));
  INV_X1     g07488(.I(new_n10333_), .ZN(new_n10348_));
  NOR4_X1    g07489(.A1(new_n2703_), .A2(pi0088), .A3(new_n8394_), .A4(new_n2687_), .ZN(new_n10349_));
  INV_X1     g07490(.I(new_n10349_), .ZN(new_n10350_));
  NOR4_X1    g07491(.A1(new_n5952_), .A2(pi0090), .A3(new_n2890_), .A4(new_n10350_), .ZN(new_n10351_));
  NOR2_X1    g07492(.A1(new_n9888_), .A2(new_n2928_), .ZN(new_n10352_));
  OAI21_X1   g07493(.A1(new_n5953_), .A2(new_n10351_), .B(new_n10352_), .ZN(new_n10353_));
  NAND4_X1   g07494(.A1(new_n10353_), .A2(pi0122), .A3(pi0829), .A4(new_n10348_), .ZN(new_n10354_));
  OAI21_X1   g07495(.A1(new_n10353_), .A2(new_n5366_), .B(new_n10348_), .ZN(new_n10355_));
  OAI21_X1   g07496(.A1(new_n10355_), .A2(pi0829), .B(new_n10354_), .ZN(new_n10356_));
  INV_X1     g07497(.I(new_n7946_), .ZN(new_n10357_));
  INV_X1     g07498(.I(new_n2934_), .ZN(new_n10358_));
  OAI21_X1   g07499(.A1(new_n10349_), .A2(pi0097), .B(new_n2936_), .ZN(new_n10359_));
  OAI21_X1   g07500(.A1(new_n10358_), .A2(new_n10359_), .B(new_n6020_), .ZN(new_n10360_));
  NOR2_X1    g07501(.A1(new_n5950_), .A2(new_n2480_), .ZN(new_n10361_));
  NAND2_X1   g07502(.A1(new_n6017_), .A2(new_n2658_), .ZN(new_n10362_));
  AOI21_X1   g07503(.A1(new_n10360_), .A2(new_n10361_), .B(new_n10362_), .ZN(new_n10363_));
  OAI21_X1   g07504(.A1(new_n10363_), .A2(new_n10357_), .B(new_n2659_), .ZN(new_n10364_));
  AOI21_X1   g07505(.A1(new_n10357_), .A2(new_n10363_), .B(new_n10364_), .ZN(new_n10365_));
  NAND3_X1   g07506(.A1(new_n7936_), .A2(new_n2861_), .A3(pi0950), .ZN(new_n10366_));
  NOR2_X1    g07507(.A1(new_n5946_), .A2(new_n10333_), .ZN(new_n10367_));
  OAI21_X1   g07508(.A1(new_n10365_), .A2(new_n10366_), .B(new_n10367_), .ZN(new_n10368_));
  AOI21_X1   g07509(.A1(new_n10368_), .A2(new_n10356_), .B(new_n6037_), .ZN(new_n10369_));
  INV_X1     g07510(.I(new_n10334_), .ZN(new_n10370_));
  NOR2_X1    g07511(.A1(new_n10370_), .A2(new_n2958_), .ZN(new_n10371_));
  OAI21_X1   g07512(.A1(new_n10369_), .A2(new_n10371_), .B(pi1091), .ZN(new_n10372_));
  INV_X1     g07513(.I(new_n10335_), .ZN(new_n10373_));
  NAND2_X1   g07514(.A1(new_n6556_), .A2(new_n10373_), .ZN(new_n10374_));
  NAND2_X1   g07515(.A1(new_n6558_), .A2(new_n10373_), .ZN(new_n10375_));
  NAND4_X1   g07516(.A1(new_n10374_), .A2(new_n10375_), .A3(new_n5094_), .A4(new_n6453_), .ZN(new_n10376_));
  AOI21_X1   g07517(.A1(new_n6453_), .A2(new_n10335_), .B(new_n2587_), .ZN(new_n10377_));
  NAND2_X1   g07518(.A1(new_n10376_), .A2(new_n10377_), .ZN(new_n10378_));
  NAND4_X1   g07519(.A1(new_n10374_), .A2(new_n10375_), .A3(new_n5141_), .A4(new_n6559_), .ZN(new_n10379_));
  NAND2_X1   g07520(.A1(new_n6559_), .A2(new_n10335_), .ZN(new_n10380_));
  NAND4_X1   g07521(.A1(new_n10378_), .A2(new_n2587_), .A3(new_n10379_), .A4(new_n10380_), .ZN(new_n10381_));
  NOR2_X1    g07522(.A1(new_n10370_), .A2(pi1091), .ZN(new_n10382_));
  OR3_X2     g07523(.A1(new_n10353_), .A2(new_n5366_), .A3(new_n10382_), .Z(new_n10383_));
  NAND3_X1   g07524(.A1(new_n10383_), .A2(new_n3154_), .A3(new_n10267_), .ZN(new_n10384_));
  AOI21_X1   g07525(.A1(new_n10381_), .A2(pi0039), .B(new_n10384_), .ZN(new_n10385_));
  NAND3_X1   g07526(.A1(new_n10385_), .A2(new_n10347_), .A3(new_n10372_), .ZN(new_n10386_));
  AOI21_X1   g07527(.A1(new_n3198_), .A2(new_n10335_), .B(new_n3177_), .ZN(new_n10387_));
  INV_X1     g07528(.I(new_n10382_), .ZN(new_n10388_));
  NAND3_X1   g07529(.A1(new_n2490_), .A2(new_n9157_), .A3(new_n10388_), .ZN(new_n10389_));
  NOR2_X1    g07530(.A1(new_n7756_), .A2(new_n10333_), .ZN(new_n10390_));
  NOR4_X1    g07531(.A1(new_n10390_), .A2(new_n2928_), .A3(new_n2920_), .A4(new_n5114_), .ZN(new_n10391_));
  NAND2_X1   g07532(.A1(new_n2490_), .A2(new_n10391_), .ZN(new_n10392_));
  AOI21_X1   g07533(.A1(new_n10389_), .A2(new_n10392_), .B(pi0120), .ZN(new_n10393_));
  OR3_X2     g07534(.A1(new_n6007_), .A2(new_n10267_), .A3(new_n3197_), .Z(new_n10394_));
  OAI21_X1   g07535(.A1(new_n10394_), .A2(new_n10393_), .B(new_n10387_), .ZN(new_n10395_));
  NAND2_X1   g07536(.A1(new_n10395_), .A2(new_n2628_), .ZN(new_n10396_));
  NAND2_X1   g07537(.A1(new_n10273_), .A2(new_n10335_), .ZN(new_n10397_));
  NAND2_X1   g07538(.A1(new_n3173_), .A2(pi0039), .ZN(new_n10398_));
  OAI21_X1   g07539(.A1(new_n6481_), .A2(new_n10398_), .B(new_n3172_), .ZN(new_n10399_));
  AOI21_X1   g07540(.A1(new_n10397_), .A2(new_n10399_), .B(pi0087), .ZN(new_n10400_));
  NAND2_X1   g07541(.A1(new_n10396_), .A2(new_n10400_), .ZN(new_n10401_));
  AOI21_X1   g07542(.A1(new_n10386_), .A2(new_n2621_), .B(new_n10401_), .ZN(new_n10402_));
  NOR2_X1    g07543(.A1(new_n10402_), .A2(new_n10345_), .ZN(new_n10403_));
  NOR2_X1    g07544(.A1(new_n5942_), .A2(new_n6538_), .ZN(new_n10404_));
  INV_X1     g07545(.I(new_n10404_), .ZN(new_n10405_));
  NOR2_X1    g07546(.A1(new_n10388_), .A2(new_n9431_), .ZN(new_n10406_));
  NOR4_X1    g07547(.A1(new_n6011_), .A2(new_n2928_), .A3(new_n5946_), .A4(new_n10390_), .ZN(new_n10407_));
  AOI21_X1   g07548(.A1(new_n10407_), .A2(new_n2490_), .B(new_n10406_), .ZN(new_n10408_));
  OAI21_X1   g07549(.A1(new_n10269_), .A2(new_n10267_), .B(new_n10408_), .ZN(new_n10409_));
  INV_X1     g07550(.I(new_n10408_), .ZN(new_n10410_));
  NAND3_X1   g07551(.A1(new_n10269_), .A2(pi0120), .A3(new_n10410_), .ZN(new_n10411_));
  NAND3_X1   g07552(.A1(new_n10409_), .A2(new_n10411_), .A3(new_n6481_), .ZN(new_n10412_));
  NOR2_X1    g07553(.A1(new_n10258_), .A2(new_n10335_), .ZN(new_n10413_));
  NOR3_X1    g07554(.A1(new_n10413_), .A2(new_n8025_), .A3(new_n2544_), .ZN(new_n10414_));
  OAI21_X1   g07555(.A1(new_n10413_), .A2(new_n2544_), .B(pi0100), .ZN(new_n10415_));
  AOI21_X1   g07556(.A1(new_n10412_), .A2(new_n10414_), .B(new_n10415_), .ZN(new_n10416_));
  INV_X1     g07557(.I(new_n10413_), .ZN(new_n10417_));
  AOI21_X1   g07558(.A1(new_n6044_), .A2(new_n10390_), .B(new_n10406_), .ZN(new_n10418_));
  NAND2_X1   g07559(.A1(new_n6048_), .A2(new_n6429_), .ZN(new_n10419_));
  MUX2_X1    g07560(.I0(new_n10419_), .I1(new_n10418_), .S(new_n10267_), .Z(new_n10420_));
  NOR2_X1    g07561(.A1(new_n6446_), .A2(new_n10413_), .ZN(new_n10421_));
  AOI21_X1   g07562(.A1(new_n10420_), .A2(new_n6446_), .B(new_n10421_), .ZN(new_n10422_));
  NOR2_X1    g07563(.A1(new_n10413_), .A2(new_n5143_), .ZN(new_n10423_));
  AOI21_X1   g07564(.A1(new_n10420_), .A2(new_n5143_), .B(new_n10423_), .ZN(new_n10424_));
  XOR2_X1    g07565(.A1(new_n10422_), .A2(new_n10424_), .Z(new_n10425_));
  NAND2_X1   g07566(.A1(new_n10425_), .A2(new_n5141_), .ZN(new_n10426_));
  XOR2_X1    g07567(.A1(new_n10426_), .A2(new_n10422_), .Z(new_n10427_));
  NAND2_X1   g07568(.A1(new_n10417_), .A2(new_n6559_), .ZN(new_n10428_));
  AOI22_X1   g07569(.A1(new_n10427_), .A2(new_n6462_), .B1(new_n2587_), .B2(new_n10428_), .ZN(new_n10429_));
  NAND2_X1   g07570(.A1(new_n10425_), .A2(new_n5094_), .ZN(new_n10430_));
  XOR2_X1    g07571(.A1(new_n10430_), .A2(new_n10422_), .Z(new_n10431_));
  OAI21_X1   g07572(.A1(new_n6429_), .A2(new_n6452_), .B(new_n10377_), .ZN(new_n10432_));
  AOI21_X1   g07573(.A1(new_n10431_), .A2(new_n6452_), .B(new_n10432_), .ZN(new_n10433_));
  OAI21_X1   g07574(.A1(new_n10429_), .A2(new_n10433_), .B(pi0039), .ZN(new_n10434_));
  MUX2_X1    g07575(.I0(new_n10434_), .I1(new_n10417_), .S(pi0038), .Z(new_n10435_));
  NOR2_X1    g07576(.A1(new_n10435_), .A2(pi0100), .ZN(new_n10436_));
  OAI21_X1   g07577(.A1(new_n10436_), .A2(new_n10416_), .B(new_n3177_), .ZN(new_n10437_));
  NAND2_X1   g07578(.A1(new_n10394_), .A2(new_n10298_), .ZN(new_n10438_));
  NAND2_X1   g07579(.A1(new_n6428_), .A2(new_n3198_), .ZN(new_n10439_));
  OAI21_X1   g07580(.A1(new_n9431_), .A2(new_n10388_), .B(new_n10392_), .ZN(new_n10440_));
  AOI22_X1   g07581(.A1(new_n10440_), .A2(new_n10393_), .B1(new_n10439_), .B2(new_n10387_), .ZN(new_n10441_));
  AOI21_X1   g07582(.A1(new_n10438_), .A2(new_n10441_), .B(pi0075), .ZN(new_n10442_));
  NAND4_X1   g07583(.A1(new_n2514_), .A2(new_n2665_), .A3(pi0950), .A4(new_n5945_), .ZN(new_n10443_));
  INV_X1     g07584(.I(new_n10390_), .ZN(new_n10444_));
  NAND4_X1   g07585(.A1(new_n10444_), .A2(new_n2502_), .A3(new_n2649_), .A4(new_n5992_), .ZN(new_n10445_));
  NOR4_X1    g07586(.A1(new_n6011_), .A2(new_n2642_), .A3(new_n10443_), .A4(new_n10445_), .ZN(new_n10446_));
  OAI21_X1   g07587(.A1(new_n10446_), .A2(new_n10406_), .B(new_n10267_), .ZN(new_n10447_));
  OAI22_X1   g07588(.A1(new_n10261_), .A2(new_n10447_), .B1(new_n8334_), .B2(new_n10413_), .ZN(new_n10448_));
  MUX2_X1    g07589(.I0(new_n10448_), .I1(new_n10417_), .S(new_n2629_), .Z(new_n10449_));
  OAI21_X1   g07590(.A1(new_n10449_), .A2(new_n2628_), .B(new_n5941_), .ZN(new_n10450_));
  AOI21_X1   g07591(.A1(new_n10437_), .A2(new_n10442_), .B(new_n10450_), .ZN(new_n10451_));
  OAI22_X1   g07592(.A1(new_n10451_), .A2(new_n10342_), .B1(new_n10403_), .B2(new_n10405_), .ZN(new_n10452_));
  INV_X1     g07593(.I(new_n10337_), .ZN(new_n10453_));
  AOI21_X1   g07594(.A1(new_n10304_), .A2(new_n10370_), .B(new_n10453_), .ZN(new_n10454_));
  NAND2_X1   g07595(.A1(new_n10260_), .A2(new_n5991_), .ZN(new_n10455_));
  AOI21_X1   g07596(.A1(new_n6434_), .A2(new_n6429_), .B(pi0075), .ZN(new_n10456_));
  NOR2_X1    g07597(.A1(new_n10291_), .A2(new_n10280_), .ZN(new_n10457_));
  NOR2_X1    g07598(.A1(new_n6429_), .A2(new_n6452_), .ZN(new_n10458_));
  MUX2_X1    g07599(.I0(new_n6427_), .I1(new_n6046_), .S(pi1091), .Z(new_n10459_));
  NAND2_X1   g07600(.A1(new_n5130_), .A2(new_n6428_), .ZN(new_n10460_));
  OAI21_X1   g07601(.A1(new_n10459_), .A2(new_n5130_), .B(new_n10460_), .ZN(new_n10461_));
  NAND4_X1   g07602(.A1(new_n6045_), .A2(pi1091), .A3(new_n5130_), .A4(new_n5143_), .ZN(new_n10462_));
  NAND4_X1   g07603(.A1(new_n6045_), .A2(pi1091), .A3(new_n6446_), .A4(new_n6548_), .ZN(new_n10463_));
  NAND2_X1   g07604(.A1(new_n10462_), .A2(new_n10463_), .ZN(new_n10464_));
  NAND2_X1   g07605(.A1(new_n10464_), .A2(new_n5094_), .ZN(new_n10465_));
  XNOR2_X1   g07606(.A1(new_n10461_), .A2(new_n10465_), .ZN(new_n10466_));
  AOI21_X1   g07607(.A1(new_n10466_), .A2(new_n6452_), .B(new_n10458_), .ZN(new_n10467_));
  NAND2_X1   g07608(.A1(new_n10464_), .A2(new_n5141_), .ZN(new_n10468_));
  XNOR2_X1   g07609(.A1(new_n10461_), .A2(new_n10468_), .ZN(new_n10469_));
  NAND2_X1   g07610(.A1(new_n10469_), .A2(new_n6462_), .ZN(new_n10470_));
  NAND2_X1   g07611(.A1(new_n6428_), .A2(new_n6559_), .ZN(new_n10471_));
  NAND4_X1   g07612(.A1(new_n10467_), .A2(new_n10470_), .A3(new_n2587_), .A4(new_n10471_), .ZN(new_n10472_));
  MUX2_X1    g07613(.I0(new_n10472_), .I1(new_n10457_), .S(new_n3154_), .Z(new_n10473_));
  AOI21_X1   g07614(.A1(new_n6428_), .A2(pi0038), .B(pi0100), .ZN(new_n10474_));
  OAI21_X1   g07615(.A1(new_n6016_), .A2(new_n6428_), .B(new_n10474_), .ZN(new_n10475_));
  AOI21_X1   g07616(.A1(new_n10473_), .A2(new_n3172_), .B(new_n10475_), .ZN(new_n10476_));
  OAI21_X1   g07617(.A1(new_n10476_), .A2(pi0087), .B(new_n10299_), .ZN(new_n10477_));
  AOI22_X1   g07618(.A1(new_n10477_), .A2(new_n2628_), .B1(new_n10455_), .B2(new_n10456_), .ZN(new_n10478_));
  OAI21_X1   g07619(.A1(new_n10346_), .A2(pi0039), .B(new_n6057_), .ZN(new_n10479_));
  NOR2_X1    g07620(.A1(new_n6077_), .A2(pi0100), .ZN(new_n10480_));
  AOI21_X1   g07621(.A1(new_n10479_), .A2(new_n10480_), .B(pi0087), .ZN(new_n10481_));
  NAND2_X1   g07622(.A1(new_n6009_), .A2(new_n2628_), .ZN(new_n10482_));
  OAI21_X1   g07623(.A1(new_n10481_), .A2(new_n10482_), .B(new_n6071_), .ZN(new_n10483_));
  NOR2_X1    g07624(.A1(new_n10304_), .A2(new_n6844_), .ZN(new_n10484_));
  AOI22_X1   g07625(.A1(new_n10483_), .A2(new_n10484_), .B1(new_n5942_), .B2(new_n10338_), .ZN(new_n10485_));
  NOR2_X1    g07626(.A1(new_n10485_), .A2(new_n10303_), .ZN(new_n10486_));
  NAND2_X1   g07627(.A1(new_n10340_), .A2(pi0120), .ZN(new_n10487_));
  AOI21_X1   g07628(.A1(new_n10478_), .A2(new_n10486_), .B(new_n10487_), .ZN(new_n10488_));
  AOI21_X1   g07629(.A1(new_n10452_), .A2(new_n10454_), .B(new_n10488_), .ZN(new_n10489_));
  OAI21_X1   g07630(.A1(new_n10489_), .A2(new_n10256_), .B(new_n10341_), .ZN(po0278));
  INV_X1     g07631(.I(new_n10041_), .ZN(new_n10491_));
  NOR4_X1    g07632(.A1(pi0067), .A2(pi0068), .A3(pi0071), .A4(pi0084), .ZN(new_n10492_));
  NOR4_X1    g07633(.A1(new_n5108_), .A2(new_n2658_), .A3(new_n3560_), .A4(pi0161), .ZN(new_n10493_));
  AOI21_X1   g07634(.A1(new_n10491_), .A2(new_n10493_), .B(new_n3177_), .ZN(new_n10494_));
  NAND2_X1   g07635(.A1(new_n10494_), .A2(pi0232), .ZN(new_n10495_));
  NOR2_X1    g07636(.A1(pi0135), .A2(pi0136), .ZN(new_n10496_));
  INV_X1     g07637(.I(new_n10496_), .ZN(new_n10497_));
  NOR3_X1    g07638(.A1(new_n10497_), .A2(pi0130), .A3(pi0134), .ZN(new_n10498_));
  NOR4_X1    g07639(.A1(new_n10498_), .A2(pi0121), .A3(pi0126), .A4(pi0132), .ZN(new_n10499_));
  INV_X1     g07640(.I(new_n10499_), .ZN(new_n10500_));
  NOR2_X1    g07641(.A1(pi0125), .A2(pi0133), .ZN(new_n10501_));
  XOR2_X1    g07642(.A1(new_n10501_), .A2(pi0121), .Z(new_n10502_));
  NAND2_X1   g07643(.A1(new_n10500_), .A2(new_n10502_), .ZN(new_n10503_));
  NOR2_X1    g07644(.A1(new_n10492_), .A2(pi0051), .ZN(new_n10504_));
  INV_X1     g07645(.I(new_n10504_), .ZN(new_n10505_));
  NOR2_X1    g07646(.A1(new_n10505_), .A2(pi0087), .ZN(new_n10506_));
  INV_X1     g07647(.I(new_n10506_), .ZN(new_n10507_));
  NAND4_X1   g07648(.A1(new_n10503_), .A2(new_n6845_), .A3(new_n10495_), .A4(new_n10507_), .ZN(new_n10508_));
  INV_X1     g07649(.I(new_n7813_), .ZN(new_n10509_));
  NOR4_X1    g07650(.A1(new_n9651_), .A2(pi0069), .A3(new_n7888_), .A4(new_n10509_), .ZN(new_n10510_));
  NAND4_X1   g07651(.A1(new_n10510_), .A2(new_n2460_), .A3(pi0077), .A4(new_n2467_), .ZN(new_n10511_));
  NOR2_X1    g07652(.A1(new_n5965_), .A2(new_n2644_), .ZN(new_n10512_));
  INV_X1     g07653(.I(new_n10512_), .ZN(new_n10513_));
  NOR3_X1    g07654(.A1(new_n10513_), .A2(pi0024), .A3(new_n5276_), .ZN(new_n10514_));
  NAND2_X1   g07655(.A1(new_n10514_), .A2(new_n6988_), .ZN(new_n10515_));
  NOR2_X1    g07656(.A1(new_n10511_), .A2(new_n10515_), .ZN(new_n10516_));
  NAND2_X1   g07657(.A1(new_n10516_), .A2(new_n3418_), .ZN(new_n10517_));
  INV_X1     g07658(.I(new_n10517_), .ZN(new_n10518_));
  NAND2_X1   g07659(.A1(new_n10510_), .A2(new_n10228_), .ZN(new_n10519_));
  OAI21_X1   g07660(.A1(new_n2691_), .A2(new_n10519_), .B(new_n10511_), .ZN(new_n10520_));
  AND3_X2    g07661(.A1(new_n10520_), .A2(pi0024), .A3(new_n6988_), .Z(new_n10521_));
  INV_X1     g07662(.I(new_n10519_), .ZN(new_n10522_));
  NOR3_X1    g07663(.A1(new_n7014_), .A2(pi0024), .A3(new_n2691_), .ZN(new_n10523_));
  AOI21_X1   g07664(.A1(new_n10522_), .A2(new_n10523_), .B(new_n10492_), .ZN(new_n10524_));
  INV_X1     g07665(.I(new_n10524_), .ZN(new_n10525_));
  INV_X1     g07666(.I(new_n10492_), .ZN(new_n10526_));
  AOI21_X1   g07667(.A1(new_n10513_), .A2(new_n10526_), .B(pi0051), .ZN(new_n10527_));
  OAI21_X1   g07668(.A1(new_n10521_), .A2(new_n10525_), .B(new_n10527_), .ZN(new_n10528_));
  NOR2_X1    g07669(.A1(new_n10528_), .A2(new_n2485_), .ZN(new_n10529_));
  INV_X1     g07670(.I(new_n10529_), .ZN(new_n10530_));
  NAND4_X1   g07671(.A1(new_n10522_), .A2(new_n7368_), .A3(new_n7078_), .A4(new_n10512_), .ZN(new_n10531_));
  NOR3_X1    g07672(.A1(new_n10531_), .A2(new_n2861_), .A3(new_n2515_), .ZN(new_n10532_));
  INV_X1     g07673(.I(new_n10532_), .ZN(new_n10533_));
  NAND3_X1   g07674(.A1(new_n10530_), .A2(new_n10504_), .A3(new_n10533_), .ZN(new_n10534_));
  NOR2_X1    g07675(.A1(new_n10534_), .A2(new_n10518_), .ZN(new_n10535_));
  NOR2_X1    g07676(.A1(new_n10535_), .A2(new_n5108_), .ZN(new_n10536_));
  NOR2_X1    g07677(.A1(new_n8031_), .A2(new_n2861_), .ZN(new_n10537_));
  INV_X1     g07678(.I(new_n10537_), .ZN(new_n10538_));
  AOI21_X1   g07679(.A1(new_n10538_), .A2(new_n2658_), .B(new_n5109_), .ZN(new_n10539_));
  XOR2_X1    g07680(.A1(new_n10536_), .A2(new_n10539_), .Z(new_n10540_));
  INV_X1     g07681(.I(new_n10540_), .ZN(new_n10541_));
  NAND2_X1   g07682(.A1(new_n10541_), .A2(new_n7504_), .ZN(new_n10542_));
  NOR2_X1    g07683(.A1(new_n5109_), .A2(new_n2658_), .ZN(new_n10543_));
  INV_X1     g07684(.I(new_n10543_), .ZN(new_n10544_));
  NOR2_X1    g07685(.A1(new_n10544_), .A2(pi0142), .ZN(new_n10545_));
  NOR2_X1    g07686(.A1(new_n10504_), .A2(new_n5109_), .ZN(new_n10546_));
  NOR2_X1    g07687(.A1(new_n10518_), .A2(new_n10505_), .ZN(new_n10547_));
  INV_X1     g07688(.I(new_n10547_), .ZN(new_n10548_));
  NOR2_X1    g07689(.A1(new_n10529_), .A2(new_n10548_), .ZN(new_n10549_));
  NOR2_X1    g07690(.A1(new_n10549_), .A2(new_n5108_), .ZN(new_n10550_));
  NOR2_X1    g07691(.A1(new_n10550_), .A2(new_n10546_), .ZN(new_n10551_));
  INV_X1     g07692(.I(new_n10551_), .ZN(new_n10552_));
  NOR2_X1    g07693(.A1(new_n10552_), .A2(new_n10532_), .ZN(new_n10553_));
  AOI21_X1   g07694(.A1(new_n10553_), .A2(pi0144), .B(new_n10545_), .ZN(new_n10554_));
  AOI21_X1   g07695(.A1(new_n10542_), .A2(new_n10554_), .B(new_n5324_), .ZN(new_n10555_));
  NAND4_X1   g07696(.A1(new_n2707_), .A2(new_n2658_), .A3(new_n10514_), .A4(new_n9893_), .ZN(new_n10556_));
  NOR2_X1    g07697(.A1(new_n2485_), .A2(new_n5109_), .ZN(new_n10557_));
  INV_X1     g07698(.I(new_n10557_), .ZN(new_n10558_));
  NOR2_X1    g07699(.A1(new_n10556_), .A2(new_n10558_), .ZN(new_n10559_));
  INV_X1     g07700(.I(new_n10559_), .ZN(new_n10560_));
  INV_X1     g07701(.I(new_n5245_), .ZN(new_n10561_));
  AOI21_X1   g07702(.A1(new_n2861_), .A2(new_n10556_), .B(new_n10561_), .ZN(new_n10562_));
  INV_X1     g07703(.I(new_n10562_), .ZN(new_n10563_));
  NOR2_X1    g07704(.A1(new_n10563_), .A2(new_n5109_), .ZN(new_n10564_));
  NOR2_X1    g07705(.A1(new_n10536_), .A2(new_n10564_), .ZN(new_n10565_));
  NAND2_X1   g07706(.A1(new_n10565_), .A2(new_n5460_), .ZN(new_n10566_));
  NAND2_X1   g07707(.A1(new_n10566_), .A2(new_n7504_), .ZN(new_n10567_));
  INV_X1     g07708(.I(new_n10553_), .ZN(new_n10568_));
  NOR2_X1    g07709(.A1(new_n10545_), .A2(new_n7504_), .ZN(new_n10569_));
  NOR3_X1    g07710(.A1(new_n10568_), .A2(new_n10518_), .A3(new_n10569_), .ZN(new_n10570_));
  NOR4_X1    g07711(.A1(new_n10570_), .A2(new_n5460_), .A3(pi0179), .A4(pi0180), .ZN(new_n10571_));
  NAND4_X1   g07712(.A1(new_n10571_), .A2(new_n10541_), .A3(new_n10560_), .A4(new_n10567_), .ZN(new_n10572_));
  NOR2_X1    g07713(.A1(new_n10572_), .A2(new_n10555_), .ZN(new_n10573_));
  AOI21_X1   g07714(.A1(new_n10530_), .A2(new_n10504_), .B(new_n5109_), .ZN(new_n10574_));
  NOR2_X1    g07715(.A1(new_n10526_), .A2(pi0051), .ZN(new_n10575_));
  NOR3_X1    g07716(.A1(new_n10528_), .A2(new_n2485_), .A3(new_n10575_), .ZN(new_n10576_));
  INV_X1     g07717(.I(new_n10575_), .ZN(new_n10577_));
  AOI21_X1   g07718(.A1(new_n10528_), .A2(new_n3418_), .B(new_n10577_), .ZN(new_n10578_));
  OAI21_X1   g07719(.A1(new_n10576_), .A2(new_n10578_), .B(new_n5108_), .ZN(new_n10579_));
  NOR2_X1    g07720(.A1(new_n10579_), .A2(new_n5460_), .ZN(new_n10580_));
  AOI21_X1   g07721(.A1(new_n5460_), .A2(new_n10574_), .B(new_n10580_), .ZN(new_n10581_));
  NAND2_X1   g07722(.A1(new_n10581_), .A2(new_n10552_), .ZN(new_n10582_));
  NOR2_X1    g07723(.A1(new_n5109_), .A2(pi0051), .ZN(new_n10583_));
  NAND2_X1   g07724(.A1(new_n10534_), .A2(new_n10583_), .ZN(new_n10584_));
  INV_X1     g07725(.I(new_n10584_), .ZN(new_n10585_));
  NOR3_X1    g07726(.A1(new_n10536_), .A2(new_n10585_), .A3(pi0144), .ZN(new_n10586_));
  INV_X1     g07727(.I(new_n8822_), .ZN(new_n10587_));
  MUX2_X1    g07728(.I0(new_n10587_), .I1(new_n8821_), .S(pi0024), .Z(new_n10588_));
  NOR2_X1    g07729(.A1(new_n10588_), .A2(new_n2652_), .ZN(new_n10589_));
  INV_X1     g07730(.I(new_n10589_), .ZN(new_n10590_));
  AOI21_X1   g07731(.A1(new_n10590_), .A2(new_n2861_), .B(new_n10561_), .ZN(new_n10591_));
  INV_X1     g07732(.I(new_n10591_), .ZN(new_n10592_));
  NOR2_X1    g07733(.A1(new_n10592_), .A2(new_n5109_), .ZN(new_n10593_));
  OR3_X2     g07734(.A1(new_n10593_), .A2(pi0142), .A3(new_n10536_), .Z(new_n10594_));
  NAND2_X1   g07735(.A1(new_n10594_), .A2(new_n7504_), .ZN(new_n10595_));
  INV_X1     g07736(.I(new_n10536_), .ZN(new_n10596_));
  NOR2_X1    g07737(.A1(new_n10590_), .A2(new_n10558_), .ZN(new_n10597_));
  OAI21_X1   g07738(.A1(new_n10597_), .A2(new_n10539_), .B(new_n10596_), .ZN(new_n10598_));
  NOR2_X1    g07739(.A1(new_n10598_), .A2(new_n5460_), .ZN(new_n10599_));
  AOI22_X1   g07740(.A1(new_n10595_), .A2(new_n10599_), .B1(new_n10582_), .B2(new_n10586_), .ZN(new_n10600_));
  OAI21_X1   g07741(.A1(new_n10600_), .A2(pi0180), .B(new_n8983_), .ZN(new_n10601_));
  NOR2_X1    g07742(.A1(pi0024), .A2(pi0314), .ZN(new_n10602_));
  MUX2_X1    g07743(.I0(new_n8822_), .I1(new_n8821_), .S(new_n10602_), .Z(new_n10603_));
  NOR2_X1    g07744(.A1(new_n10603_), .A2(new_n2652_), .ZN(new_n10604_));
  OAI21_X1   g07745(.A1(new_n10604_), .A2(pi0072), .B(new_n5245_), .ZN(new_n10605_));
  NOR2_X1    g07746(.A1(new_n10605_), .A2(new_n5109_), .ZN(new_n10606_));
  OR3_X2     g07747(.A1(new_n10606_), .A2(pi0142), .A3(new_n10536_), .Z(new_n10607_));
  NAND2_X1   g07748(.A1(new_n10607_), .A2(new_n7504_), .ZN(new_n10608_));
  INV_X1     g07749(.I(new_n10603_), .ZN(new_n10609_));
  NAND4_X1   g07750(.A1(new_n10609_), .A2(new_n3418_), .A3(new_n2643_), .A4(new_n5964_), .ZN(new_n10610_));
  NAND2_X1   g07751(.A1(new_n10610_), .A2(new_n2658_), .ZN(new_n10611_));
  INV_X1     g07752(.I(new_n10611_), .ZN(new_n10612_));
  NOR2_X1    g07753(.A1(new_n10612_), .A2(new_n10537_), .ZN(new_n10613_));
  INV_X1     g07754(.I(new_n10613_), .ZN(new_n10614_));
  NOR2_X1    g07755(.A1(new_n10614_), .A2(new_n5109_), .ZN(new_n10615_));
  AOI21_X1   g07756(.A1(new_n5109_), .A2(new_n10535_), .B(new_n10615_), .ZN(new_n10616_));
  NOR2_X1    g07757(.A1(new_n10616_), .A2(new_n5460_), .ZN(new_n10617_));
  INV_X1     g07758(.I(new_n10535_), .ZN(new_n10618_));
  OAI21_X1   g07759(.A1(new_n10618_), .A2(new_n10569_), .B(new_n5324_), .ZN(new_n10619_));
  AOI21_X1   g07760(.A1(new_n10617_), .A2(new_n10608_), .B(new_n10619_), .ZN(new_n10620_));
  AOI21_X1   g07761(.A1(new_n10620_), .A2(new_n10601_), .B(new_n10573_), .ZN(new_n10621_));
  NOR2_X1    g07762(.A1(new_n10544_), .A2(pi0146), .ZN(new_n10622_));
  NOR2_X1    g07763(.A1(new_n2587_), .A2(pi0158), .ZN(new_n10623_));
  INV_X1     g07764(.I(new_n10623_), .ZN(new_n10624_));
  NAND2_X1   g07765(.A1(new_n10574_), .A2(new_n3560_), .ZN(new_n10626_));
  OAI21_X1   g07766(.A1(new_n3560_), .A2(new_n10579_), .B(new_n10626_), .ZN(new_n10627_));
  NOR2_X1    g07767(.A1(new_n5340_), .A2(new_n2587_), .ZN(new_n10629_));
  NOR2_X1    g07768(.A1(new_n8974_), .A2(new_n4701_), .ZN(new_n10631_));
  NOR2_X1    g07769(.A1(new_n10531_), .A2(new_n2485_), .ZN(new_n10632_));
  NOR2_X1    g07770(.A1(new_n10632_), .A2(new_n10505_), .ZN(new_n10633_));
  OAI21_X1   g07771(.A1(new_n10633_), .A2(new_n10622_), .B(pi0161), .ZN(new_n10634_));
  INV_X1     g07772(.I(new_n10633_), .ZN(new_n10635_));
  NOR2_X1    g07773(.A1(new_n10635_), .A2(new_n5108_), .ZN(new_n10636_));
  AOI21_X1   g07774(.A1(new_n3162_), .A2(new_n5108_), .B(new_n10636_), .ZN(new_n10637_));
  INV_X1     g07775(.I(new_n10637_), .ZN(new_n10638_));
  NOR2_X1    g07776(.A1(new_n7945_), .A2(new_n8588_), .ZN(new_n10639_));
  NOR2_X1    g07777(.A1(new_n10639_), .A2(pi0051), .ZN(new_n10640_));
  INV_X1     g07778(.I(new_n10640_), .ZN(new_n10641_));
  NOR2_X1    g07779(.A1(new_n10641_), .A2(new_n5109_), .ZN(new_n10642_));
  NOR2_X1    g07780(.A1(new_n10636_), .A2(new_n10642_), .ZN(new_n10643_));
  INV_X1     g07781(.I(new_n10643_), .ZN(new_n10644_));
  MUX2_X1    g07782(.I0(new_n10644_), .I1(new_n10638_), .S(new_n3560_), .Z(new_n10645_));
  NAND2_X1   g07783(.A1(new_n10645_), .A2(new_n4701_), .ZN(new_n10646_));
  AOI21_X1   g07784(.A1(new_n10646_), .A2(new_n10634_), .B(new_n5357_), .ZN(new_n10647_));
  NOR2_X1    g07785(.A1(new_n5109_), .A2(pi0287), .ZN(new_n10648_));
  INV_X1     g07786(.I(new_n10648_), .ZN(new_n10649_));
  NOR2_X1    g07787(.A1(new_n10649_), .A2(pi0051), .ZN(new_n10650_));
  NOR2_X1    g07788(.A1(new_n10644_), .A2(new_n10650_), .ZN(new_n10651_));
  NOR2_X1    g07789(.A1(new_n10651_), .A2(pi0161), .ZN(new_n10652_));
  NOR2_X1    g07790(.A1(new_n10652_), .A2(new_n10622_), .ZN(new_n10653_));
  AOI21_X1   g07791(.A1(new_n10632_), .A2(new_n10649_), .B(new_n10505_), .ZN(new_n10654_));
  NAND2_X1   g07792(.A1(new_n10654_), .A2(pi0161), .ZN(new_n10655_));
  NOR2_X1    g07793(.A1(new_n5356_), .A2(new_n2562_), .ZN(new_n10656_));
  OAI21_X1   g07794(.A1(new_n10653_), .A2(new_n10655_), .B(new_n10656_), .ZN(new_n10657_));
  INV_X1     g07795(.I(new_n7593_), .ZN(new_n10658_));
  INV_X1     g07796(.I(new_n10493_), .ZN(new_n10659_));
  AOI21_X1   g07797(.A1(new_n10505_), .A2(new_n10659_), .B(new_n5356_), .ZN(new_n10660_));
  NOR2_X1    g07798(.A1(new_n10660_), .A2(new_n10658_), .ZN(new_n10661_));
  OAI21_X1   g07799(.A1(new_n10647_), .A2(new_n10657_), .B(new_n10661_), .ZN(new_n10662_));
  AOI21_X1   g07800(.A1(new_n10633_), .A2(new_n2658_), .B(new_n10543_), .ZN(new_n10663_));
  INV_X1     g07801(.I(new_n10663_), .ZN(new_n10664_));
  OAI21_X1   g07802(.A1(new_n10545_), .A2(new_n10504_), .B(new_n6051_), .ZN(new_n10665_));
  NOR2_X1    g07803(.A1(new_n2658_), .A2(new_n5460_), .ZN(new_n10666_));
  INV_X1     g07804(.I(new_n10666_), .ZN(new_n10667_));
  NOR2_X1    g07805(.A1(new_n6051_), .A2(pi0144), .ZN(new_n10668_));
  NAND4_X1   g07806(.A1(new_n10664_), .A2(new_n10665_), .A3(new_n10667_), .A4(new_n10668_), .ZN(new_n10669_));
  INV_X1     g07807(.I(new_n10546_), .ZN(new_n10670_));
  NOR2_X1    g07808(.A1(new_n10670_), .A2(new_n10666_), .ZN(new_n10671_));
  INV_X1     g07809(.I(new_n10671_), .ZN(new_n10672_));
  NOR2_X1    g07810(.A1(new_n10633_), .A2(pi0051), .ZN(new_n10673_));
  INV_X1     g07811(.I(new_n10673_), .ZN(new_n10674_));
  OAI21_X1   g07812(.A1(new_n10674_), .A2(new_n10575_), .B(pi0287), .ZN(new_n10675_));
  NOR2_X1    g07813(.A1(new_n10675_), .A2(new_n5109_), .ZN(new_n10676_));
  INV_X1     g07814(.I(new_n10676_), .ZN(new_n10677_));
  NAND2_X1   g07815(.A1(new_n7153_), .A2(new_n10526_), .ZN(new_n10678_));
  AOI21_X1   g07816(.A1(new_n10677_), .A2(new_n10672_), .B(new_n10678_), .ZN(new_n10679_));
  OAI21_X1   g07817(.A1(new_n10679_), .A2(new_n10669_), .B(pi0181), .ZN(new_n10680_));
  AOI21_X1   g07818(.A1(new_n10638_), .A2(new_n10643_), .B(new_n5460_), .ZN(new_n10681_));
  OAI21_X1   g07819(.A1(new_n10681_), .A2(pi0224), .B(new_n6050_), .ZN(new_n10682_));
  NOR2_X1    g07820(.A1(new_n10577_), .A2(new_n5109_), .ZN(new_n10683_));
  OR3_X2     g07821(.A1(new_n10683_), .A2(new_n10504_), .A3(new_n10545_), .Z(new_n10684_));
  AOI21_X1   g07822(.A1(new_n10684_), .A2(new_n6051_), .B(pi0144), .ZN(new_n10685_));
  NOR4_X1    g07823(.A1(new_n10644_), .A2(new_n2595_), .A3(new_n10545_), .A4(new_n10650_), .ZN(new_n10686_));
  NOR3_X1    g07824(.A1(new_n10682_), .A2(new_n10685_), .A3(new_n10686_), .ZN(new_n10687_));
  NAND2_X1   g07825(.A1(new_n10681_), .A2(new_n6050_), .ZN(new_n10688_));
  AND3_X2    g07826(.A1(new_n10669_), .A2(new_n5325_), .A3(new_n2587_), .Z(new_n10689_));
  OAI21_X1   g07827(.A1(new_n10688_), .A2(new_n10685_), .B(new_n10689_), .ZN(new_n10690_));
  AOI21_X1   g07828(.A1(new_n10687_), .A2(new_n10680_), .B(new_n10690_), .ZN(new_n10691_));
  NAND2_X1   g07829(.A1(new_n10662_), .A2(new_n10691_), .ZN(new_n10692_));
  INV_X1     g07830(.I(new_n10632_), .ZN(new_n10693_));
  NOR2_X1    g07831(.A1(new_n6051_), .A2(pi0299), .ZN(new_n10694_));
  NOR2_X1    g07832(.A1(new_n5483_), .A2(new_n10694_), .ZN(new_n10695_));
  OAI21_X1   g07833(.A1(new_n10693_), .A2(new_n10695_), .B(new_n5987_), .ZN(new_n10696_));
  NOR2_X1    g07834(.A1(new_n10504_), .A2(pi0039), .ZN(new_n10697_));
  OR2_X2     g07835(.A1(new_n10647_), .A2(new_n10660_), .Z(new_n10698_));
  NOR2_X1    g07836(.A1(new_n7401_), .A2(pi0232), .ZN(new_n10699_));
  AOI22_X1   g07837(.A1(new_n10698_), .A2(new_n10699_), .B1(new_n10696_), .B2(new_n10697_), .ZN(new_n10700_));
  AOI22_X1   g07838(.A1(new_n10700_), .A2(new_n10692_), .B1(new_n5863_), .B2(new_n10618_), .ZN(new_n10701_));
  NAND3_X1   g07839(.A1(new_n10533_), .A2(new_n10526_), .A3(new_n10583_), .ZN(new_n10702_));
  NOR2_X1    g07840(.A1(new_n10702_), .A2(new_n10518_), .ZN(new_n10703_));
  INV_X1     g07841(.I(new_n10703_), .ZN(new_n10704_));
  AOI22_X1   g07842(.A1(new_n10704_), .A2(new_n10544_), .B1(pi0146), .B2(new_n10505_), .ZN(new_n10705_));
  NOR4_X1    g07843(.A1(new_n10618_), .A2(pi0161), .A3(new_n5108_), .A4(new_n10705_), .ZN(new_n10706_));
  NOR4_X1    g07844(.A1(new_n10540_), .A2(new_n3560_), .A3(new_n4701_), .A4(new_n10559_), .ZN(new_n10707_));
  OAI21_X1   g07845(.A1(new_n10707_), .A2(new_n10706_), .B(new_n10623_), .ZN(new_n10708_));
  NOR4_X1    g07846(.A1(new_n10533_), .A2(pi0051), .A3(new_n5108_), .A4(new_n10526_), .ZN(new_n10709_));
  NOR4_X1    g07847(.A1(new_n10568_), .A2(new_n3560_), .A3(pi0161), .A4(new_n10536_), .ZN(new_n10710_));
  NOR3_X1    g07848(.A1(new_n10541_), .A2(pi0161), .A3(new_n10622_), .ZN(new_n10711_));
  OAI21_X1   g07849(.A1(new_n10711_), .A2(new_n10710_), .B(new_n10629_), .ZN(new_n10712_));
  AOI21_X1   g07850(.A1(new_n10712_), .A2(new_n10708_), .B(pi0156), .ZN(new_n10713_));
  NOR4_X1    g07851(.A1(new_n10701_), .A2(new_n10713_), .A3(new_n7178_), .A4(new_n10631_), .ZN(new_n10714_));
  OAI21_X1   g07852(.A1(new_n10621_), .A2(pi0299), .B(new_n10714_), .ZN(new_n10715_));
  NOR2_X1    g07853(.A1(new_n10672_), .A2(new_n10569_), .ZN(new_n10716_));
  INV_X1     g07854(.I(new_n10716_), .ZN(new_n10717_));
  NAND3_X1   g07855(.A1(new_n10717_), .A2(pi0299), .A3(new_n10493_), .ZN(new_n10718_));
  OAI21_X1   g07856(.A1(new_n2587_), .A2(new_n10493_), .B(new_n10716_), .ZN(new_n10719_));
  AOI21_X1   g07857(.A1(new_n10718_), .A2(new_n10719_), .B(new_n5987_), .ZN(new_n10720_));
  NOR4_X1    g07858(.A1(new_n10720_), .A2(pi0038), .A3(pi0100), .A4(new_n10504_), .ZN(new_n10721_));
  INV_X1     g07859(.I(new_n10720_), .ZN(new_n10722_));
  AOI21_X1   g07860(.A1(new_n10504_), .A2(pi0100), .B(new_n2541_), .ZN(new_n10723_));
  OAI21_X1   g07861(.A1(new_n10722_), .A2(new_n3173_), .B(new_n10723_), .ZN(new_n10724_));
  AOI21_X1   g07862(.A1(new_n10715_), .A2(new_n10721_), .B(new_n10724_), .ZN(new_n10725_));
  INV_X1     g07863(.I(new_n10622_), .ZN(new_n10726_));
  INV_X1     g07864(.I(new_n10597_), .ZN(new_n10727_));
  NAND2_X1   g07865(.A1(new_n10727_), .A2(new_n10726_), .ZN(new_n10728_));
  MUX2_X1    g07866(.I0(new_n10728_), .I1(new_n10627_), .S(new_n4701_), .Z(new_n10729_));
  NOR2_X1    g07867(.A1(new_n10611_), .A2(new_n5109_), .ZN(new_n10730_));
  INV_X1     g07868(.I(new_n10730_), .ZN(new_n10731_));
  AOI21_X1   g07869(.A1(pi0051), .A2(pi0146), .B(new_n10731_), .ZN(new_n10732_));
  NOR2_X1    g07870(.A1(new_n10521_), .A2(new_n10525_), .ZN(new_n10733_));
  NOR4_X1    g07871(.A1(new_n10516_), .A2(new_n2658_), .A3(new_n10492_), .A4(new_n10513_), .ZN(new_n10734_));
  NAND2_X1   g07872(.A1(new_n10733_), .A2(new_n10734_), .ZN(new_n10735_));
  MUX2_X1    g07873(.I0(new_n10577_), .I1(new_n10735_), .S(new_n3418_), .Z(new_n10736_));
  NOR2_X1    g07874(.A1(new_n10736_), .A2(new_n5109_), .ZN(new_n10737_));
  NOR2_X1    g07875(.A1(new_n10549_), .A2(new_n5109_), .ZN(new_n10738_));
  OAI21_X1   g07876(.A1(new_n10738_), .A2(new_n3560_), .B(new_n4701_), .ZN(new_n10739_));
  AOI21_X1   g07877(.A1(pi0146), .A2(new_n10737_), .B(new_n10739_), .ZN(new_n10740_));
  OAI21_X1   g07878(.A1(new_n10732_), .A2(new_n4701_), .B(new_n10740_), .ZN(new_n10741_));
  NAND2_X1   g07879(.A1(new_n10741_), .A2(new_n10629_), .ZN(new_n10742_));
  NAND4_X1   g07880(.A1(new_n10742_), .A2(new_n5987_), .A3(new_n10624_), .A4(new_n10729_), .ZN(new_n10743_));
  NOR3_X1    g07881(.A1(new_n10730_), .A2(pi0144), .A3(new_n10667_), .ZN(new_n10744_));
  NOR3_X1    g07882(.A1(new_n10736_), .A2(new_n5460_), .A3(new_n5109_), .ZN(new_n10745_));
  NOR2_X1    g07883(.A1(new_n10738_), .A2(new_n5460_), .ZN(new_n10746_));
  NOR4_X1    g07884(.A1(new_n10744_), .A2(pi0144), .A3(new_n10745_), .A4(new_n10746_), .ZN(new_n10747_));
  NAND2_X1   g07885(.A1(new_n10581_), .A2(new_n7504_), .ZN(new_n10748_));
  NAND3_X1   g07886(.A1(new_n10727_), .A2(new_n8983_), .A3(new_n10569_), .ZN(new_n10749_));
  OAI21_X1   g07887(.A1(new_n10749_), .A2(new_n10748_), .B(new_n5324_), .ZN(new_n10750_));
  NAND4_X1   g07888(.A1(new_n10516_), .A2(new_n2658_), .A3(new_n3418_), .A4(new_n10526_), .ZN(new_n10751_));
  XOR2_X1    g07889(.A1(new_n10751_), .A2(new_n10577_), .Z(new_n10752_));
  NAND2_X1   g07890(.A1(new_n10752_), .A2(new_n5108_), .ZN(new_n10753_));
  INV_X1     g07891(.I(new_n10753_), .ZN(new_n10754_));
  NOR2_X1    g07892(.A1(new_n10547_), .A2(new_n5109_), .ZN(new_n10755_));
  OAI21_X1   g07893(.A1(pi0142), .A2(new_n10755_), .B(new_n10754_), .ZN(new_n10756_));
  INV_X1     g07894(.I(new_n10755_), .ZN(new_n10757_));
  NOR3_X1    g07895(.A1(new_n10754_), .A2(pi0142), .A3(new_n10757_), .ZN(new_n10758_));
  NAND2_X1   g07896(.A1(new_n7504_), .A2(new_n5324_), .ZN(new_n10759_));
  NOR3_X1    g07897(.A1(new_n10758_), .A2(new_n10560_), .A3(new_n10759_), .ZN(new_n10760_));
  OAI21_X1   g07898(.A1(new_n10717_), .A2(pi0180), .B(new_n8983_), .ZN(new_n10761_));
  AOI21_X1   g07899(.A1(new_n10760_), .A2(new_n10756_), .B(new_n10761_), .ZN(new_n10762_));
  OAI21_X1   g07900(.A1(new_n10747_), .A2(new_n10750_), .B(new_n10762_), .ZN(new_n10763_));
  NAND2_X1   g07901(.A1(new_n10726_), .A2(pi0161), .ZN(new_n10766_));
  NAND4_X1   g07902(.A1(new_n10659_), .A2(new_n5340_), .A3(new_n5987_), .A4(pi0299), .ZN(new_n10769_));
  NAND2_X1   g07903(.A1(new_n10769_), .A2(new_n8974_), .ZN(new_n10770_));
  OAI21_X1   g07904(.A1(new_n10720_), .A2(new_n3172_), .B(new_n3173_), .ZN(new_n10771_));
  NAND3_X1   g07905(.A1(new_n10771_), .A2(new_n2545_), .A3(new_n10770_), .ZN(new_n10772_));
  NOR3_X1    g07906(.A1(new_n10493_), .A2(pi0159), .A3(new_n2587_), .ZN(new_n10773_));
  INV_X1     g07907(.I(new_n10639_), .ZN(new_n10774_));
  MUX2_X1    g07908(.I0(new_n10774_), .I1(new_n2491_), .S(pi0142), .Z(new_n10775_));
  NOR2_X1    g07909(.A1(new_n10677_), .A2(new_n7154_), .ZN(new_n10776_));
  NAND2_X1   g07910(.A1(new_n7153_), .A2(new_n10648_), .ZN(new_n10777_));
  NOR4_X1    g07911(.A1(new_n10569_), .A2(new_n10777_), .A3(pi0144), .A4(pi0181), .ZN(new_n10778_));
  NAND2_X1   g07912(.A1(new_n10778_), .A2(new_n10672_), .ZN(new_n10779_));
  NOR3_X1    g07913(.A1(new_n10776_), .A2(new_n10775_), .A3(new_n10779_), .ZN(new_n10780_));
  NOR2_X1    g07914(.A1(new_n10622_), .A2(pi0161), .ZN(new_n10781_));
  NOR2_X1    g07915(.A1(new_n5359_), .A2(new_n5109_), .ZN(new_n10782_));
  NAND3_X1   g07916(.A1(new_n10782_), .A2(new_n7634_), .A3(new_n10766_), .ZN(new_n10783_));
  AOI21_X1   g07917(.A1(new_n10677_), .A2(new_n10781_), .B(new_n10783_), .ZN(new_n10784_));
  NAND3_X1   g07918(.A1(new_n7634_), .A2(new_n10658_), .A3(new_n10493_), .ZN(new_n10785_));
  AOI21_X1   g07919(.A1(new_n10716_), .A2(new_n5325_), .B(pi0299), .ZN(new_n10786_));
  OAI21_X1   g07920(.A1(new_n10784_), .A2(new_n10785_), .B(new_n10786_), .ZN(new_n10787_));
  OAI22_X1   g07921(.A1(new_n10787_), .A2(new_n10780_), .B1(new_n7927_), .B2(new_n10773_), .ZN(new_n10788_));
  NOR2_X1    g07922(.A1(new_n10722_), .A2(new_n3173_), .ZN(new_n10789_));
  NOR4_X1    g07923(.A1(new_n10789_), .A2(new_n8974_), .A3(new_n2540_), .A4(new_n2545_), .ZN(new_n10790_));
  NAND3_X1   g07924(.A1(new_n10788_), .A2(new_n10772_), .A3(new_n10790_), .ZN(new_n10791_));
  AOI21_X1   g07925(.A1(new_n10763_), .A2(new_n2587_), .B(new_n10791_), .ZN(new_n10792_));
  NAND2_X1   g07926(.A1(pi0163), .A2(pi0299), .ZN(new_n10793_));
  OAI21_X1   g07927(.A1(new_n8883_), .A2(pi0299), .B(new_n10793_), .ZN(new_n10794_));
  AOI21_X1   g07928(.A1(new_n5988_), .A2(new_n10794_), .B(new_n3177_), .ZN(new_n10795_));
  NOR2_X1    g07929(.A1(new_n3229_), .A2(pi0087), .ZN(new_n10796_));
  NOR3_X1    g07930(.A1(new_n10503_), .A2(new_n10795_), .A3(new_n10796_), .ZN(new_n10797_));
  NAND2_X1   g07931(.A1(new_n10720_), .A2(new_n10797_), .ZN(new_n10798_));
  AOI21_X1   g07932(.A1(new_n10743_), .A2(new_n10792_), .B(new_n10798_), .ZN(new_n10799_));
  INV_X1     g07933(.I(new_n10796_), .ZN(new_n10800_));
  NOR2_X1    g07934(.A1(new_n10800_), .A2(new_n10504_), .ZN(new_n10801_));
  NOR2_X1    g07935(.A1(new_n10503_), .A2(new_n10795_), .ZN(new_n10802_));
  OAI21_X1   g07936(.A1(new_n10722_), .A2(new_n10801_), .B(new_n10802_), .ZN(new_n10803_));
  OAI21_X1   g07937(.A1(new_n10799_), .A2(po1038), .B(new_n10803_), .ZN(new_n10804_));
  OAI21_X1   g07938(.A1(new_n10725_), .A2(new_n10804_), .B(new_n10508_), .ZN(po0279));
  NOR3_X1    g07939(.A1(new_n10302_), .A2(new_n5942_), .A3(po1038), .ZN(new_n10806_));
  OAI21_X1   g07940(.A1(new_n10483_), .A2(new_n10405_), .B(new_n10806_), .ZN(new_n10807_));
  OAI22_X1   g07941(.A1(new_n10478_), .A2(new_n10807_), .B1(new_n6429_), .B2(new_n6951_), .ZN(po0280));
  NOR2_X1    g07942(.A1(new_n7600_), .A2(pi0110), .ZN(new_n10809_));
  NAND3_X1   g07943(.A1(new_n5133_), .A2(new_n5356_), .A3(new_n10809_), .ZN(new_n10810_));
  NOR2_X1    g07944(.A1(new_n2587_), .A2(pi0039), .ZN(new_n10811_));
  INV_X1     g07945(.I(new_n10811_), .ZN(new_n10812_));
  NOR2_X1    g07946(.A1(new_n10810_), .A2(new_n10812_), .ZN(new_n10813_));
  INV_X1     g07947(.I(new_n10813_), .ZN(new_n10814_));
  NOR2_X1    g07948(.A1(new_n2779_), .A2(new_n2783_), .ZN(new_n10815_));
  INV_X1     g07949(.I(new_n10815_), .ZN(new_n10816_));
  NAND2_X1   g07950(.A1(new_n2767_), .A2(new_n7889_), .ZN(new_n10817_));
  AOI21_X1   g07951(.A1(new_n9899_), .A2(pi0111), .B(new_n10817_), .ZN(new_n10818_));
  OAI21_X1   g07952(.A1(new_n5260_), .A2(pi0111), .B(new_n10818_), .ZN(new_n10819_));
  NAND2_X1   g07953(.A1(new_n10819_), .A2(pi0069), .ZN(new_n10820_));
  XOR2_X1    g07954(.A1(new_n10820_), .A2(new_n2780_), .Z(new_n10821_));
  NAND2_X1   g07955(.A1(new_n10821_), .A2(new_n2768_), .ZN(new_n10822_));
  INV_X1     g07956(.I(new_n10822_), .ZN(new_n10823_));
  NOR2_X1    g07957(.A1(new_n10823_), .A2(new_n10816_), .ZN(new_n10824_));
  INV_X1     g07958(.I(new_n10824_), .ZN(new_n10825_));
  AOI21_X1   g07959(.A1(new_n10823_), .A2(new_n10816_), .B(pi0083), .ZN(new_n10826_));
  AOI21_X1   g07960(.A1(new_n10825_), .A2(new_n10826_), .B(new_n2790_), .ZN(new_n10827_));
  OAI21_X1   g07961(.A1(new_n10827_), .A2(pi0071), .B(new_n5249_), .ZN(new_n10828_));
  NAND2_X1   g07962(.A1(new_n8671_), .A2(new_n2441_), .ZN(new_n10829_));
  INV_X1     g07963(.I(new_n10829_), .ZN(new_n10830_));
  AOI21_X1   g07964(.A1(new_n10828_), .A2(new_n10830_), .B(pi0090), .ZN(new_n10831_));
  OAI22_X1   g07965(.A1(new_n10831_), .A2(new_n2648_), .B1(pi0093), .B2(new_n2840_), .ZN(new_n10832_));
  NOR2_X1    g07966(.A1(new_n9896_), .A2(pi0072), .ZN(new_n10833_));
  AOI21_X1   g07967(.A1(new_n10832_), .A2(new_n10833_), .B(new_n5245_), .ZN(new_n10834_));
  INV_X1     g07968(.I(new_n10831_), .ZN(new_n10835_));
  NAND2_X1   g07969(.A1(new_n7989_), .A2(new_n2839_), .ZN(new_n10836_));
  NAND4_X1   g07970(.A1(new_n10835_), .A2(new_n2647_), .A3(new_n7199_), .A4(new_n10836_), .ZN(new_n10837_));
  NOR2_X1    g07971(.A1(new_n2652_), .A2(new_n2861_), .ZN(new_n10838_));
  AOI21_X1   g07972(.A1(new_n7989_), .A2(new_n10838_), .B(new_n2515_), .ZN(new_n10839_));
  AOI21_X1   g07973(.A1(new_n10837_), .A2(new_n10839_), .B(pi0110), .ZN(new_n10840_));
  OAI22_X1   g07974(.A1(new_n10840_), .A2(new_n9897_), .B1(pi0039), .B2(new_n10834_), .ZN(new_n10841_));
  NOR2_X1    g07975(.A1(new_n3232_), .A2(pi0038), .ZN(new_n10842_));
  INV_X1     g07976(.I(new_n10842_), .ZN(new_n10843_));
  AOI21_X1   g07977(.A1(new_n10841_), .A2(new_n10814_), .B(new_n10843_), .ZN(new_n10844_));
  AOI21_X1   g07978(.A1(new_n9896_), .A2(pi0110), .B(pi0039), .ZN(new_n10845_));
  OAI21_X1   g07979(.A1(new_n10845_), .A2(new_n10813_), .B(new_n10843_), .ZN(new_n10846_));
  NAND2_X1   g07980(.A1(new_n10846_), .A2(new_n6845_), .ZN(new_n10847_));
  NAND3_X1   g07981(.A1(new_n10810_), .A2(pi0039), .A3(new_n6845_), .ZN(new_n10850_));
  OAI21_X1   g07982(.A1(new_n10844_), .A2(new_n10847_), .B(new_n10850_), .ZN(po0281));
  NOR2_X1    g07983(.A1(new_n2490_), .A2(new_n5108_), .ZN(new_n10852_));
  AOI21_X1   g07984(.A1(new_n10674_), .A2(new_n5108_), .B(new_n10852_), .ZN(new_n10853_));
  INV_X1     g07985(.I(new_n10853_), .ZN(new_n10854_));
  NOR4_X1    g07986(.A1(new_n10677_), .A2(new_n2595_), .A3(new_n6050_), .A4(new_n10854_), .ZN(new_n10855_));
  AOI21_X1   g07987(.A1(new_n6051_), .A2(new_n10683_), .B(new_n10855_), .ZN(new_n10856_));
  INV_X1     g07988(.I(new_n10856_), .ZN(new_n10857_));
  NAND2_X1   g07989(.A1(new_n10857_), .A2(new_n7151_), .ZN(new_n10858_));
  AOI21_X1   g07990(.A1(new_n6559_), .A2(new_n10777_), .B(new_n2491_), .ZN(new_n10859_));
  NAND2_X1   g07991(.A1(new_n10859_), .A2(pi0174), .ZN(new_n10860_));
  AOI21_X1   g07992(.A1(new_n10858_), .A2(new_n7179_), .B(new_n10860_), .ZN(new_n10861_));
  NOR2_X1    g07993(.A1(new_n10635_), .A2(new_n5109_), .ZN(new_n10862_));
  NOR2_X1    g07994(.A1(new_n10862_), .A2(new_n10852_), .ZN(new_n10863_));
  INV_X1     g07995(.I(new_n10863_), .ZN(new_n10864_));
  NOR2_X1    g07996(.A1(new_n10693_), .A2(new_n10649_), .ZN(new_n10865_));
  NAND3_X1   g07997(.A1(new_n10865_), .A2(new_n2595_), .A3(new_n6051_), .ZN(new_n10866_));
  AOI22_X1   g07998(.A1(new_n10864_), .A2(new_n6462_), .B1(new_n10670_), .B2(new_n10866_), .ZN(new_n10867_));
  NOR2_X1    g07999(.A1(new_n10774_), .A2(new_n10649_), .ZN(new_n10868_));
  NOR2_X1    g08000(.A1(new_n10868_), .A2(new_n10543_), .ZN(new_n10869_));
  AOI21_X1   g08001(.A1(new_n10869_), .A2(pi0224), .B(new_n6051_), .ZN(new_n10870_));
  INV_X1     g08002(.I(new_n10870_), .ZN(new_n10871_));
  NOR2_X1    g08003(.A1(new_n10642_), .A2(new_n10852_), .ZN(new_n10872_));
  NOR2_X1    g08004(.A1(new_n10872_), .A2(new_n6559_), .ZN(new_n10873_));
  AOI21_X1   g08005(.A1(new_n10873_), .A2(new_n10871_), .B(new_n10543_), .ZN(new_n10874_));
  INV_X1     g08006(.I(new_n10874_), .ZN(new_n10875_));
  MUX2_X1    g08007(.I0(new_n10875_), .I1(new_n10867_), .S(pi0174), .Z(new_n10876_));
  AND2_X2    g08008(.A1(new_n10876_), .A2(new_n7179_), .Z(new_n10877_));
  NOR2_X1    g08009(.A1(new_n10546_), .A2(new_n6462_), .ZN(new_n10878_));
  OAI21_X1   g08010(.A1(new_n10854_), .A2(new_n10878_), .B(pi0174), .ZN(new_n10879_));
  NOR2_X1    g08011(.A1(new_n2491_), .A2(new_n6559_), .ZN(new_n10880_));
  OAI21_X1   g08012(.A1(new_n10544_), .A2(new_n7179_), .B(new_n5324_), .ZN(new_n10881_));
  AOI21_X1   g08013(.A1(new_n10880_), .A2(pi0174), .B(new_n10881_), .ZN(new_n10882_));
  NAND2_X1   g08014(.A1(new_n10879_), .A2(new_n10882_), .ZN(new_n10883_));
  AOI21_X1   g08015(.A1(new_n10883_), .A2(new_n2587_), .B(pi0180), .ZN(new_n10884_));
  OAI21_X1   g08016(.A1(new_n10861_), .A2(new_n10877_), .B(new_n10884_), .ZN(new_n10885_));
  NOR2_X1    g08017(.A1(new_n10865_), .A2(new_n10546_), .ZN(new_n10886_));
  NOR4_X1    g08018(.A1(new_n10886_), .A2(new_n3250_), .A3(pi0172), .A4(new_n10869_), .ZN(new_n10887_));
  NAND3_X1   g08019(.A1(new_n10677_), .A2(pi0152), .A3(new_n10782_), .ZN(new_n10888_));
  OAI21_X1   g08020(.A1(new_n3250_), .A2(new_n10782_), .B(new_n10676_), .ZN(new_n10889_));
  AOI21_X1   g08021(.A1(new_n10888_), .A2(new_n10889_), .B(pi0172), .ZN(new_n10890_));
  INV_X1     g08022(.I(new_n10872_), .ZN(new_n10891_));
  NAND2_X1   g08023(.A1(new_n10891_), .A2(pi0152), .ZN(new_n10892_));
  AOI22_X1   g08024(.A1(new_n10864_), .A2(new_n3250_), .B1(pi0051), .B2(new_n3707_), .ZN(new_n10893_));
  AOI21_X1   g08025(.A1(new_n10893_), .A2(new_n10892_), .B(pi0216), .ZN(new_n10894_));
  INV_X1     g08026(.I(new_n10629_), .ZN(new_n10895_));
  NOR2_X1    g08027(.A1(new_n10544_), .A2(new_n3707_), .ZN(new_n10896_));
  INV_X1     g08028(.I(new_n10683_), .ZN(new_n10897_));
  NOR2_X1    g08029(.A1(new_n10897_), .A2(pi0152), .ZN(new_n10898_));
  NOR2_X1    g08030(.A1(new_n10898_), .A2(new_n10896_), .ZN(new_n10899_));
  INV_X1     g08031(.I(new_n10899_), .ZN(new_n10900_));
  AOI21_X1   g08032(.A1(new_n10900_), .A2(new_n5357_), .B(new_n10895_), .ZN(new_n10901_));
  NOR4_X1    g08033(.A1(new_n10894_), .A2(pi0216), .A3(new_n5356_), .A4(new_n10901_), .ZN(new_n10902_));
  OAI21_X1   g08034(.A1(new_n10887_), .A2(new_n10890_), .B(new_n10902_), .ZN(new_n10903_));
  NAND2_X1   g08035(.A1(new_n10894_), .A2(new_n5356_), .ZN(new_n10904_));
  AOI21_X1   g08036(.A1(new_n10900_), .A2(new_n6452_), .B(new_n10624_), .ZN(new_n10905_));
  AOI22_X1   g08037(.A1(new_n10885_), .A2(new_n10903_), .B1(new_n10904_), .B2(new_n10905_), .ZN(new_n10906_));
  AOI21_X1   g08038(.A1(new_n10538_), .A2(new_n5987_), .B(pi0039), .ZN(new_n10907_));
  NOR2_X1    g08039(.A1(new_n6453_), .A2(new_n2587_), .ZN(new_n10908_));
  AOI21_X1   g08040(.A1(new_n2587_), .A2(new_n6462_), .B(new_n10908_), .ZN(new_n10909_));
  NAND3_X1   g08041(.A1(new_n3172_), .A2(new_n3154_), .A3(pi0232), .ZN(new_n10910_));
  NOR3_X1    g08042(.A1(new_n10906_), .A2(new_n10907_), .A3(new_n10910_), .ZN(new_n10911_));
  NOR2_X1    g08043(.A1(new_n10538_), .A2(new_n5108_), .ZN(new_n10912_));
  NOR2_X1    g08044(.A1(new_n10593_), .A2(new_n10912_), .ZN(new_n10913_));
  NOR2_X1    g08045(.A1(new_n10585_), .A2(new_n10912_), .ZN(new_n10914_));
  NOR3_X1    g08046(.A1(new_n10913_), .A2(new_n3250_), .A3(new_n3707_), .ZN(new_n10915_));
  NOR3_X1    g08047(.A1(new_n10597_), .A2(new_n10543_), .A3(new_n10537_), .ZN(new_n10916_));
  NOR2_X1    g08048(.A1(new_n10537_), .A2(new_n5108_), .ZN(new_n10917_));
  NOR2_X1    g08049(.A1(new_n10534_), .A2(new_n10702_), .ZN(new_n10918_));
  NOR2_X1    g08050(.A1(new_n10918_), .A2(new_n10917_), .ZN(new_n10919_));
  INV_X1     g08051(.I(new_n10919_), .ZN(new_n10920_));
  NAND4_X1   g08052(.A1(new_n10916_), .A2(new_n10920_), .A3(pi0152), .A4(new_n3707_), .ZN(new_n10921_));
  NAND2_X1   g08053(.A1(new_n10921_), .A2(new_n5339_), .ZN(new_n10922_));
  OAI21_X1   g08054(.A1(new_n10915_), .A2(new_n10922_), .B(new_n7640_), .ZN(new_n10923_));
  NOR2_X1    g08055(.A1(new_n10606_), .A2(new_n10912_), .ZN(new_n10924_));
  INV_X1     g08056(.I(new_n10924_), .ZN(new_n10925_));
  NAND2_X1   g08057(.A1(new_n10731_), .A2(new_n10538_), .ZN(new_n10926_));
  NOR4_X1    g08058(.A1(new_n10926_), .A2(pi0152), .A3(new_n3707_), .A4(new_n10925_), .ZN(new_n10927_));
  AOI21_X1   g08059(.A1(new_n10618_), .A2(new_n2658_), .B(new_n5109_), .ZN(new_n10928_));
  XOR2_X1    g08060(.A1(new_n10928_), .A2(new_n10917_), .Z(new_n10929_));
  INV_X1     g08061(.I(new_n10929_), .ZN(new_n10930_));
  INV_X1     g08062(.I(new_n10896_), .ZN(new_n10931_));
  NAND2_X1   g08063(.A1(new_n10931_), .A2(new_n3250_), .ZN(new_n10932_));
  OAI21_X1   g08064(.A1(new_n10930_), .A2(new_n10932_), .B(pi0197), .ZN(new_n10933_));
  NOR2_X1    g08065(.A1(new_n10927_), .A2(new_n10933_), .ZN(new_n10934_));
  NOR2_X1    g08066(.A1(new_n10564_), .A2(new_n10912_), .ZN(new_n10935_));
  NOR3_X1    g08067(.A1(new_n10537_), .A2(new_n10543_), .A3(new_n10559_), .ZN(new_n10936_));
  NAND3_X1   g08068(.A1(new_n10935_), .A2(new_n3707_), .A3(new_n10936_), .ZN(new_n10937_));
  OAI22_X1   g08069(.A1(new_n10564_), .A2(new_n10912_), .B1(pi0172), .B2(new_n10936_), .ZN(new_n10938_));
  AOI22_X1   g08070(.A1(new_n10937_), .A2(new_n10938_), .B1(pi0152), .B2(pi0197), .ZN(new_n10939_));
  OAI21_X1   g08071(.A1(new_n10703_), .A2(new_n10917_), .B(new_n10543_), .ZN(new_n10940_));
  AOI21_X1   g08072(.A1(new_n10940_), .A2(new_n3250_), .B(pi0197), .ZN(new_n10941_));
  AOI21_X1   g08073(.A1(new_n10709_), .A2(new_n3250_), .B(pi0197), .ZN(new_n10942_));
  NOR2_X1    g08074(.A1(new_n5109_), .A2(pi0152), .ZN(new_n10943_));
  NAND2_X1   g08075(.A1(new_n10538_), .A2(new_n10943_), .ZN(new_n10944_));
  OAI21_X1   g08076(.A1(new_n10942_), .A2(new_n10944_), .B(new_n10931_), .ZN(new_n10945_));
  OAI22_X1   g08077(.A1(new_n10941_), .A2(new_n10945_), .B1(pi0038), .B2(pi0155), .ZN(new_n10946_));
  OAI21_X1   g08078(.A1(new_n10939_), .A2(new_n10946_), .B(pi0299), .ZN(new_n10947_));
  AOI21_X1   g08079(.A1(new_n10934_), .A2(new_n10923_), .B(new_n10947_), .ZN(new_n10948_));
  AOI21_X1   g08080(.A1(new_n10913_), .A2(new_n5323_), .B(new_n10924_), .ZN(new_n10949_));
  NOR3_X1    g08081(.A1(new_n10913_), .A2(pi0145), .A3(new_n10925_), .ZN(new_n10950_));
  NOR3_X1    g08082(.A1(new_n10950_), .A2(new_n10949_), .A3(pi0193), .ZN(new_n10951_));
  OAI21_X1   g08083(.A1(new_n10544_), .A2(new_n7179_), .B(pi0145), .ZN(new_n10952_));
  NOR2_X1    g08084(.A1(new_n10930_), .A2(new_n10952_), .ZN(new_n10953_));
  NOR2_X1    g08085(.A1(new_n10914_), .A2(pi0193), .ZN(new_n10954_));
  NOR2_X1    g08086(.A1(new_n10954_), .A2(pi0145), .ZN(new_n10955_));
  NAND2_X1   g08087(.A1(new_n10919_), .A2(pi0193), .ZN(new_n10956_));
  OAI21_X1   g08088(.A1(new_n10955_), .A2(new_n10956_), .B(new_n7151_), .ZN(new_n10957_));
  OAI21_X1   g08089(.A1(new_n10953_), .A2(new_n10957_), .B(new_n7621_), .ZN(new_n10958_));
  NAND2_X1   g08090(.A1(new_n10958_), .A2(new_n7151_), .ZN(new_n10959_));
  NOR2_X1    g08091(.A1(new_n10912_), .A2(new_n10709_), .ZN(new_n10960_));
  NOR3_X1    g08092(.A1(new_n10940_), .A2(new_n5323_), .A3(new_n7151_), .ZN(new_n10961_));
  NAND2_X1   g08093(.A1(new_n10935_), .A2(pi0145), .ZN(new_n10962_));
  AOI21_X1   g08094(.A1(new_n10538_), .A2(new_n5323_), .B(pi0174), .ZN(new_n10963_));
  AOI21_X1   g08095(.A1(new_n10962_), .A2(new_n10963_), .B(new_n10961_), .ZN(new_n10964_));
  OAI21_X1   g08096(.A1(new_n10559_), .A2(new_n10543_), .B(pi0145), .ZN(new_n10965_));
  NAND3_X1   g08097(.A1(new_n10560_), .A2(new_n5323_), .A3(new_n10543_), .ZN(new_n10966_));
  NAND3_X1   g08098(.A1(new_n10538_), .A2(new_n10965_), .A3(new_n10966_), .ZN(new_n10967_));
  NOR2_X1    g08099(.A1(new_n10518_), .A2(new_n10543_), .ZN(new_n10968_));
  NAND2_X1   g08100(.A1(new_n10702_), .A2(pi0145), .ZN(new_n10969_));
  OAI21_X1   g08101(.A1(new_n10969_), .A2(new_n10968_), .B(new_n7151_), .ZN(new_n10970_));
  NAND2_X1   g08102(.A1(new_n7151_), .A2(new_n7179_), .ZN(new_n10971_));
  AOI21_X1   g08103(.A1(new_n10970_), .A2(new_n10917_), .B(new_n10971_), .ZN(new_n10972_));
  AOI21_X1   g08104(.A1(new_n10972_), .A2(new_n10967_), .B(new_n7616_), .ZN(new_n10973_));
  OAI21_X1   g08105(.A1(new_n10964_), .A2(pi0193), .B(new_n10973_), .ZN(new_n10974_));
  OAI21_X1   g08106(.A1(new_n10959_), .A2(new_n10951_), .B(new_n10974_), .ZN(new_n10975_));
  AOI21_X1   g08107(.A1(new_n10975_), .A2(new_n3172_), .B(new_n10948_), .ZN(new_n10976_));
  OAI22_X1   g08108(.A1(new_n10976_), .A2(new_n7178_), .B1(pi0100), .B2(new_n10911_), .ZN(new_n10977_));
  INV_X1     g08109(.I(new_n10549_), .ZN(new_n10978_));
  AOI21_X1   g08110(.A1(new_n10978_), .A2(new_n5987_), .B(pi0039), .ZN(new_n10979_));
  NOR2_X1    g08111(.A1(new_n10979_), .A2(pi0038), .ZN(new_n10980_));
  MUX2_X1    g08112(.I0(new_n10635_), .I1(new_n8019_), .S(new_n5108_), .Z(new_n10981_));
  AOI21_X1   g08113(.A1(new_n10505_), .A2(new_n5109_), .B(new_n7153_), .ZN(new_n10982_));
  INV_X1     g08114(.I(new_n10982_), .ZN(new_n10983_));
  OAI21_X1   g08115(.A1(new_n10981_), .A2(new_n7154_), .B(new_n10983_), .ZN(new_n10984_));
  AOI21_X1   g08116(.A1(new_n10632_), .A2(new_n7153_), .B(new_n10505_), .ZN(new_n10985_));
  INV_X1     g08117(.I(new_n10985_), .ZN(new_n10986_));
  NOR2_X1    g08118(.A1(new_n10654_), .A2(pi0051), .ZN(new_n10987_));
  NOR2_X1    g08119(.A1(new_n10987_), .A2(new_n5109_), .ZN(new_n10988_));
  INV_X1     g08120(.I(new_n10988_), .ZN(new_n10989_));
  NAND2_X1   g08121(.A1(new_n10989_), .A2(new_n10986_), .ZN(new_n10990_));
  MUX2_X1    g08122(.I0(new_n10990_), .I1(new_n10984_), .S(new_n7151_), .Z(new_n10991_));
  NOR2_X1    g08123(.A1(new_n10991_), .A2(new_n5324_), .ZN(new_n10992_));
  AOI21_X1   g08124(.A1(new_n10638_), .A2(new_n7153_), .B(new_n10982_), .ZN(new_n10993_));
  INV_X1     g08125(.I(new_n10993_), .ZN(new_n10994_));
  NOR2_X1    g08126(.A1(new_n10985_), .A2(new_n10543_), .ZN(new_n10995_));
  NAND3_X1   g08127(.A1(new_n10994_), .A2(pi0174), .A3(new_n10995_), .ZN(new_n10996_));
  OAI21_X1   g08128(.A1(new_n7151_), .A2(new_n10995_), .B(new_n10993_), .ZN(new_n10997_));
  AOI21_X1   g08129(.A1(new_n10996_), .A2(new_n10997_), .B(pi0180), .ZN(new_n10998_));
  NOR2_X1    g08130(.A1(new_n5324_), .A2(pi0174), .ZN(new_n10999_));
  NAND2_X1   g08131(.A1(new_n10654_), .A2(new_n10999_), .ZN(new_n11000_));
  AOI21_X1   g08132(.A1(new_n10650_), .A2(new_n10999_), .B(pi0193), .ZN(new_n11001_));
  OAI21_X1   g08133(.A1(new_n11000_), .A2(new_n10985_), .B(new_n11001_), .ZN(new_n11002_));
  AOI21_X1   g08134(.A1(new_n11002_), .A2(new_n2587_), .B(pi0193), .ZN(new_n11003_));
  OAI21_X1   g08135(.A1(new_n10998_), .A2(new_n10992_), .B(new_n11003_), .ZN(new_n11004_));
  AOI21_X1   g08136(.A1(new_n10633_), .A2(new_n10943_), .B(new_n10641_), .ZN(new_n11005_));
  INV_X1     g08137(.I(new_n10943_), .ZN(new_n11006_));
  NOR3_X1    g08138(.A1(new_n10633_), .A2(new_n10640_), .A3(new_n11006_), .ZN(new_n11007_));
  NOR3_X1    g08139(.A1(new_n11007_), .A2(new_n11005_), .A3(pi0172), .ZN(new_n11008_));
  NOR4_X1    g08140(.A1(new_n10638_), .A2(new_n3250_), .A3(pi0172), .A4(new_n10664_), .ZN(new_n11009_));
  NOR3_X1    g08141(.A1(new_n11009_), .A2(new_n7634_), .A3(new_n11008_), .ZN(new_n11010_));
  NOR2_X1    g08142(.A1(new_n10654_), .A2(new_n10896_), .ZN(new_n11011_));
  NAND2_X1   g08143(.A1(new_n7634_), .A2(new_n3250_), .ZN(new_n11012_));
  AOI21_X1   g08144(.A1(new_n10931_), .A2(new_n3250_), .B(new_n5340_), .ZN(new_n11013_));
  OAI21_X1   g08145(.A1(new_n11011_), .A2(new_n11012_), .B(new_n11013_), .ZN(new_n11014_));
  NOR2_X1    g08146(.A1(new_n5340_), .A2(pi0299), .ZN(new_n11015_));
  OAI21_X1   g08147(.A1(new_n10651_), .A2(new_n11014_), .B(new_n11015_), .ZN(new_n11016_));
  NOR2_X1    g08148(.A1(new_n10900_), .A2(new_n10504_), .ZN(new_n11017_));
  OAI22_X1   g08149(.A1(new_n11010_), .A2(new_n11016_), .B1(new_n7170_), .B2(new_n11017_), .ZN(new_n11018_));
  NOR2_X1    g08150(.A1(new_n10693_), .A2(new_n7634_), .ZN(new_n11019_));
  NOR2_X1    g08151(.A1(new_n11019_), .A2(new_n10505_), .ZN(new_n11020_));
  NAND2_X1   g08152(.A1(new_n3154_), .A2(pi0232), .ZN(new_n11021_));
  AOI21_X1   g08153(.A1(new_n11004_), .A2(new_n11018_), .B(new_n11021_), .ZN(new_n11022_));
  AOI21_X1   g08154(.A1(new_n10504_), .A2(new_n3172_), .B(pi0100), .ZN(new_n11023_));
  OAI21_X1   g08155(.A1(new_n11022_), .A2(new_n10980_), .B(new_n11023_), .ZN(new_n11024_));
  NOR2_X1    g08156(.A1(new_n10550_), .A2(new_n10754_), .ZN(new_n11025_));
  NOR2_X1    g08157(.A1(new_n10550_), .A2(new_n10559_), .ZN(new_n11026_));
  NOR4_X1    g08158(.A1(new_n11025_), .A2(new_n11026_), .A3(new_n3250_), .A4(pi0172), .ZN(new_n11027_));
  NOR2_X1    g08159(.A1(new_n10550_), .A2(new_n10755_), .ZN(new_n11028_));
  NAND2_X1   g08160(.A1(new_n11028_), .A2(pi0152), .ZN(new_n11029_));
  NAND3_X1   g08161(.A1(new_n11026_), .A2(new_n3250_), .A3(new_n10544_), .ZN(new_n11030_));
  NAND4_X1   g08162(.A1(new_n11030_), .A2(new_n11029_), .A3(new_n3707_), .A4(new_n5339_), .ZN(new_n11031_));
  NOR2_X1    g08163(.A1(new_n10897_), .A2(new_n3250_), .ZN(new_n11032_));
  OAI21_X1   g08164(.A1(new_n10550_), .A2(new_n11032_), .B(pi0172), .ZN(new_n11033_));
  NOR4_X1    g08165(.A1(new_n10551_), .A2(pi0172), .A3(new_n5339_), .A4(new_n10898_), .ZN(new_n11034_));
  NAND2_X1   g08166(.A1(new_n7640_), .A2(pi0299), .ZN(new_n11035_));
  AOI21_X1   g08167(.A1(new_n11034_), .A2(new_n11033_), .B(new_n11035_), .ZN(new_n11036_));
  OAI21_X1   g08168(.A1(new_n11027_), .A2(new_n11031_), .B(new_n11036_), .ZN(new_n11037_));
  NAND3_X1   g08169(.A1(new_n10604_), .A2(new_n3418_), .A3(new_n5109_), .ZN(new_n11038_));
  XOR2_X1    g08170(.A1(new_n11038_), .A2(new_n10738_), .Z(new_n11039_));
  NOR2_X1    g08171(.A1(new_n10737_), .A2(new_n10550_), .ZN(new_n11040_));
  OAI21_X1   g08172(.A1(new_n11039_), .A2(new_n11040_), .B(pi0152), .ZN(new_n11041_));
  NOR2_X1    g08173(.A1(new_n11041_), .A2(new_n3707_), .ZN(new_n11042_));
  OAI21_X1   g08174(.A1(new_n10549_), .A2(new_n10943_), .B(new_n3707_), .ZN(new_n11043_));
  NAND3_X1   g08175(.A1(new_n10730_), .A2(new_n3250_), .A3(new_n11043_), .ZN(new_n11044_));
  NAND2_X1   g08176(.A1(new_n11044_), .A2(new_n5339_), .ZN(new_n11045_));
  INV_X1     g08177(.I(new_n10550_), .ZN(new_n11046_));
  NAND2_X1   g08178(.A1(new_n10727_), .A2(new_n11046_), .ZN(new_n11047_));
  NAND2_X1   g08179(.A1(new_n11047_), .A2(new_n3250_), .ZN(new_n11048_));
  NAND2_X1   g08180(.A1(new_n11046_), .A2(new_n10579_), .ZN(new_n11049_));
  NAND2_X1   g08181(.A1(new_n11049_), .A2(pi0172), .ZN(new_n11050_));
  NOR2_X1    g08182(.A1(new_n10547_), .A2(new_n5108_), .ZN(new_n11051_));
  NOR2_X1    g08183(.A1(new_n11051_), .A2(new_n10546_), .ZN(new_n11052_));
  NAND2_X1   g08184(.A1(new_n10530_), .A2(new_n11052_), .ZN(new_n11053_));
  AOI21_X1   g08185(.A1(new_n11053_), .A2(new_n3707_), .B(pi0152), .ZN(new_n11054_));
  NAND3_X1   g08186(.A1(new_n10543_), .A2(new_n3707_), .A3(new_n5339_), .ZN(new_n11055_));
  AOI21_X1   g08187(.A1(new_n11050_), .A2(new_n11054_), .B(new_n11055_), .ZN(new_n11056_));
  NAND3_X1   g08188(.A1(new_n3172_), .A2(new_n7639_), .A3(pi0299), .ZN(new_n11057_));
  AOI21_X1   g08189(.A1(new_n11048_), .A2(new_n11056_), .B(new_n11057_), .ZN(new_n11058_));
  OAI21_X1   g08190(.A1(new_n11042_), .A2(new_n11045_), .B(new_n11058_), .ZN(new_n11059_));
  INV_X1     g08191(.I(new_n11039_), .ZN(new_n11060_));
  NOR2_X1    g08192(.A1(new_n11060_), .A2(new_n5323_), .ZN(new_n11061_));
  NOR2_X1    g08193(.A1(new_n11047_), .A2(new_n5323_), .ZN(new_n11062_));
  INV_X1     g08194(.I(new_n11040_), .ZN(new_n11063_));
  AOI21_X1   g08195(.A1(new_n5323_), .A2(new_n10548_), .B(new_n11053_), .ZN(new_n11064_));
  NAND4_X1   g08196(.A1(new_n11063_), .A2(new_n7151_), .A3(new_n3418_), .A4(new_n11064_), .ZN(new_n11065_));
  NAND3_X1   g08197(.A1(new_n11065_), .A2(new_n7151_), .A3(pi0193), .ZN(new_n11066_));
  NOR3_X1    g08198(.A1(new_n11061_), .A2(new_n11066_), .A3(new_n11062_), .ZN(new_n11067_));
  NOR3_X1    g08199(.A1(new_n11047_), .A2(pi0051), .A3(new_n5323_), .ZN(new_n11068_));
  NAND2_X1   g08200(.A1(new_n11046_), .A2(new_n5323_), .ZN(new_n11069_));
  OAI22_X1   g08201(.A1(new_n11068_), .A2(pi0174), .B1(new_n10730_), .B2(new_n11069_), .ZN(new_n11070_));
  NOR2_X1    g08202(.A1(new_n10550_), .A2(new_n10543_), .ZN(new_n11071_));
  INV_X1     g08203(.I(new_n11071_), .ZN(new_n11072_));
  NAND2_X1   g08204(.A1(new_n11028_), .A2(pi0174), .ZN(new_n11073_));
  AOI21_X1   g08205(.A1(new_n11073_), .A2(new_n11072_), .B(pi0193), .ZN(new_n11074_));
  NAND3_X1   g08206(.A1(new_n10753_), .A2(new_n5323_), .A3(pi0174), .ZN(new_n11075_));
  NAND2_X1   g08207(.A1(new_n10897_), .A2(pi0145), .ZN(new_n11076_));
  XOR2_X1    g08208(.A1(new_n11075_), .A2(new_n11076_), .Z(new_n11077_));
  OAI21_X1   g08209(.A1(new_n10560_), .A2(pi0145), .B(new_n7151_), .ZN(new_n11078_));
  NAND2_X1   g08210(.A1(new_n11046_), .A2(pi0193), .ZN(new_n11079_));
  AOI21_X1   g08211(.A1(new_n11077_), .A2(new_n11078_), .B(new_n11079_), .ZN(new_n11080_));
  OAI21_X1   g08212(.A1(new_n11080_), .A2(new_n11074_), .B(new_n7622_), .ZN(new_n11081_));
  NAND2_X1   g08213(.A1(new_n11064_), .A2(new_n7151_), .ZN(new_n11082_));
  NOR4_X1    g08214(.A1(pi0038), .A2(pi0177), .A3(pi0193), .A4(pi0299), .ZN(new_n11083_));
  NAND4_X1   g08215(.A1(new_n11070_), .A2(new_n11081_), .A3(new_n11082_), .A4(new_n11083_), .ZN(new_n11084_));
  NAND2_X1   g08216(.A1(pi0125), .A2(pi0133), .ZN(new_n11085_));
  NAND2_X1   g08217(.A1(new_n10500_), .A2(new_n10501_), .ZN(new_n11086_));
  NAND2_X1   g08218(.A1(new_n11086_), .A2(new_n11085_), .ZN(new_n11087_));
  NOR2_X1    g08219(.A1(new_n2587_), .A2(pi0162), .ZN(new_n11088_));
  NOR2_X1    g08220(.A1(pi0140), .A2(pi0299), .ZN(new_n11089_));
  NOR2_X1    g08221(.A1(new_n11088_), .A2(new_n11089_), .ZN(new_n11090_));
  AOI21_X1   g08222(.A1(new_n5988_), .A2(new_n11090_), .B(new_n3177_), .ZN(new_n11091_));
  NOR4_X1    g08223(.A1(new_n11087_), .A2(new_n7177_), .A3(new_n10723_), .A4(new_n11091_), .ZN(new_n11092_));
  OAI21_X1   g08224(.A1(new_n11084_), .A2(new_n11067_), .B(new_n11092_), .ZN(new_n11093_));
  AOI21_X1   g08225(.A1(new_n11037_), .A2(new_n11059_), .B(new_n11093_), .ZN(new_n11094_));
  OAI21_X1   g08226(.A1(new_n11087_), .A2(new_n10505_), .B(new_n3177_), .ZN(new_n11095_));
  AOI21_X1   g08227(.A1(new_n10900_), .A2(pi0232), .B(new_n11095_), .ZN(new_n11096_));
  NOR2_X1    g08228(.A1(new_n5989_), .A2(new_n3177_), .ZN(new_n11097_));
  NAND2_X1   g08229(.A1(new_n11097_), .A2(pi0162), .ZN(new_n11098_));
  OAI21_X1   g08230(.A1(new_n11096_), .A2(new_n11098_), .B(new_n6845_), .ZN(new_n11099_));
  AOI21_X1   g08231(.A1(new_n11094_), .A2(new_n11024_), .B(new_n11099_), .ZN(new_n11100_));
  OAI21_X1   g08232(.A1(new_n10977_), .A2(new_n2540_), .B(new_n11100_), .ZN(po0282));
  NOR3_X1    g08233(.A1(pi0121), .A2(pi0125), .A3(pi0133), .ZN(new_n11102_));
  OR4_X2     g08234(.A1(pi0126), .A2(new_n10498_), .A3(pi0132), .A4(new_n11102_), .Z(new_n11103_));
  NOR2_X1    g08235(.A1(new_n10683_), .A2(pi0051), .ZN(new_n11104_));
  INV_X1     g08236(.I(new_n11104_), .ZN(new_n11105_));
  AOI21_X1   g08237(.A1(new_n11105_), .A2(pi0232), .B(new_n11103_), .ZN(new_n11106_));
  OAI21_X1   g08238(.A1(new_n7928_), .A2(new_n10526_), .B(pi0051), .ZN(new_n11107_));
  NOR3_X1    g08239(.A1(new_n5109_), .A2(pi0051), .A3(new_n2526_), .ZN(new_n11108_));
  XOR2_X1    g08240(.A1(new_n11107_), .A2(new_n11108_), .Z(new_n11109_));
  INV_X1     g08241(.I(new_n11109_), .ZN(new_n11110_));
  NOR2_X1    g08242(.A1(new_n10504_), .A2(pi0232), .ZN(new_n11111_));
  OAI21_X1   g08243(.A1(new_n11106_), .A2(new_n11110_), .B(new_n11111_), .ZN(new_n11112_));
  OAI21_X1   g08244(.A1(new_n11112_), .A2(new_n10133_), .B(pi0087), .ZN(new_n11113_));
  NOR2_X1    g08245(.A1(new_n11113_), .A2(new_n6845_), .ZN(new_n11114_));
  NAND2_X1   g08246(.A1(new_n10940_), .A2(new_n8872_), .ZN(new_n11115_));
  NAND2_X1   g08247(.A1(new_n10935_), .A2(pi0189), .ZN(new_n11116_));
  NAND3_X1   g08248(.A1(new_n11116_), .A2(new_n11115_), .A3(new_n7345_), .ZN(new_n11117_));
  NOR3_X1    g08249(.A1(new_n10930_), .A2(new_n8872_), .A3(new_n10924_), .ZN(new_n11118_));
  AOI21_X1   g08250(.A1(pi0189), .A2(new_n10924_), .B(new_n10929_), .ZN(new_n11119_));
  OAI21_X1   g08251(.A1(new_n11118_), .A2(new_n11119_), .B(pi0178), .ZN(new_n11120_));
  INV_X1     g08252(.I(new_n10960_), .ZN(new_n11121_));
  NOR2_X1    g08253(.A1(new_n10538_), .A2(new_n8872_), .ZN(new_n11122_));
  INV_X1     g08254(.I(new_n11122_), .ZN(new_n11123_));
  NOR2_X1    g08255(.A1(new_n10543_), .A2(pi0178), .ZN(new_n11124_));
  AOI22_X1   g08256(.A1(new_n11121_), .A2(new_n8872_), .B1(new_n11123_), .B2(new_n11124_), .ZN(new_n11125_));
  AOI21_X1   g08257(.A1(new_n11120_), .A2(new_n11117_), .B(new_n5325_), .ZN(new_n11127_));
  NAND2_X1   g08258(.A1(new_n10543_), .A2(pi0153), .ZN(new_n11128_));
  AOI22_X1   g08259(.A1(new_n10940_), .A2(new_n10117_), .B1(new_n4549_), .B2(new_n11128_), .ZN(new_n11129_));
  OAI21_X1   g08260(.A1(new_n10930_), .A2(new_n10117_), .B(new_n11129_), .ZN(new_n11130_));
  NOR4_X1    g08261(.A1(new_n10926_), .A2(new_n2526_), .A3(pi0157), .A4(new_n10925_), .ZN(new_n11131_));
  INV_X1     g08262(.I(new_n10936_), .ZN(new_n11132_));
  NOR3_X1    g08263(.A1(new_n10935_), .A2(pi0153), .A3(new_n11132_), .ZN(new_n11133_));
  AOI21_X1   g08264(.A1(new_n10935_), .A2(new_n2526_), .B(new_n10936_), .ZN(new_n11134_));
  NOR4_X1    g08265(.A1(new_n11131_), .A2(pi0157), .A3(new_n11133_), .A4(new_n11134_), .ZN(new_n11135_));
  OAI21_X1   g08266(.A1(new_n11135_), .A2(new_n4549_), .B(new_n11130_), .ZN(new_n11136_));
  NOR2_X1    g08267(.A1(new_n11072_), .A2(pi0189), .ZN(new_n11137_));
  INV_X1     g08268(.I(new_n11137_), .ZN(new_n11138_));
  NAND2_X1   g08269(.A1(new_n10926_), .A2(new_n11138_), .ZN(new_n11139_));
  NOR3_X1    g08270(.A1(new_n10929_), .A2(pi0178), .A3(pi0189), .ZN(new_n11140_));
  NOR4_X1    g08271(.A1(new_n11115_), .A2(new_n8872_), .A3(new_n10543_), .A4(new_n11132_), .ZN(new_n11141_));
  OAI21_X1   g08272(.A1(new_n11141_), .A2(pi0178), .B(pi0181), .ZN(new_n11142_));
  AOI21_X1   g08273(.A1(new_n11139_), .A2(new_n11140_), .B(new_n11142_), .ZN(new_n11143_));
  NAND3_X1   g08274(.A1(new_n8915_), .A2(new_n7345_), .A3(pi0189), .ZN(new_n11144_));
  NOR4_X1    g08275(.A1(new_n10919_), .A2(pi0181), .A3(new_n11125_), .A4(new_n11144_), .ZN(new_n11145_));
  OAI21_X1   g08276(.A1(new_n10916_), .A2(new_n8872_), .B(new_n11145_), .ZN(new_n11146_));
  OR3_X2     g08277(.A1(new_n10913_), .A2(new_n2526_), .A3(new_n4549_), .Z(new_n11147_));
  NAND4_X1   g08278(.A1(new_n10916_), .A2(new_n10920_), .A3(new_n2526_), .A4(pi0166), .ZN(new_n11148_));
  AOI21_X1   g08279(.A1(new_n11147_), .A2(new_n11148_), .B(new_n10117_), .ZN(new_n11149_));
  MUX2_X1    g08280(.I0(new_n11121_), .I1(new_n10537_), .S(pi0166), .Z(new_n11150_));
  NAND2_X1   g08281(.A1(new_n11128_), .A2(new_n10117_), .ZN(new_n11151_));
  OAI21_X1   g08282(.A1(new_n11150_), .A2(new_n11151_), .B(new_n7401_), .ZN(new_n11152_));
  OAI22_X1   g08283(.A1(new_n11149_), .A2(new_n11152_), .B1(new_n11143_), .B2(new_n11146_), .ZN(new_n11153_));
  NAND3_X1   g08284(.A1(new_n11153_), .A2(new_n10658_), .A3(new_n11136_), .ZN(new_n11154_));
  OAI21_X1   g08285(.A1(new_n11154_), .A2(new_n11127_), .B(pi0232), .ZN(new_n11155_));
  OAI21_X1   g08286(.A1(new_n10854_), .A2(new_n10878_), .B(pi0189), .ZN(new_n11156_));
  NAND2_X1   g08287(.A1(new_n10880_), .A2(pi0189), .ZN(new_n11157_));
  NAND3_X1   g08288(.A1(new_n11156_), .A2(new_n5326_), .A3(new_n11157_), .ZN(new_n11159_));
  NAND2_X1   g08289(.A1(new_n11159_), .A2(new_n8871_), .ZN(new_n11160_));
  AOI22_X1   g08290(.A1(new_n10864_), .A2(new_n4549_), .B1(pi0051), .B2(new_n2526_), .ZN(new_n11161_));
  OAI21_X1   g08291(.A1(new_n4549_), .A2(new_n10872_), .B(new_n11161_), .ZN(new_n11162_));
  INV_X1     g08292(.I(new_n10886_), .ZN(new_n11163_));
  OAI21_X1   g08293(.A1(new_n11163_), .A2(new_n10869_), .B(pi0166), .ZN(new_n11164_));
  NOR2_X1    g08294(.A1(new_n10676_), .A2(new_n4549_), .ZN(new_n11165_));
  INV_X1     g08295(.I(new_n10782_), .ZN(new_n11166_));
  NOR2_X1    g08296(.A1(new_n11166_), .A2(new_n4549_), .ZN(new_n11167_));
  NOR4_X1    g08297(.A1(new_n11165_), .A2(pi0153), .A3(new_n5338_), .A4(new_n11167_), .ZN(new_n11168_));
  OAI21_X1   g08298(.A1(new_n2526_), .A2(new_n11164_), .B(new_n11168_), .ZN(new_n11169_));
  MUX2_X1    g08299(.I0(new_n11169_), .I1(new_n11162_), .S(new_n2562_), .Z(new_n11170_));
  NOR2_X1    g08300(.A1(new_n11170_), .A2(new_n5357_), .ZN(new_n11171_));
  NOR2_X1    g08301(.A1(new_n11110_), .A2(new_n11104_), .ZN(new_n11172_));
  NOR4_X1    g08302(.A1(new_n11172_), .A2(pi0160), .A3(new_n2562_), .A4(new_n5356_), .ZN(new_n11173_));
  OAI21_X1   g08303(.A1(new_n11171_), .A2(new_n11173_), .B(new_n2587_), .ZN(new_n11174_));
  NAND2_X1   g08304(.A1(new_n11174_), .A2(new_n11160_), .ZN(new_n11175_));
  NAND3_X1   g08305(.A1(new_n11156_), .A2(new_n5326_), .A3(new_n11157_), .ZN(new_n11176_));
  MUX2_X1    g08306(.I0(new_n10875_), .I1(new_n10867_), .S(pi0189), .Z(new_n11177_));
  AOI22_X1   g08307(.A1(new_n11177_), .A2(new_n5326_), .B1(new_n10544_), .B2(new_n11176_), .ZN(new_n11178_));
  NOR2_X1    g08308(.A1(new_n11178_), .A2(new_n8915_), .ZN(new_n11179_));
  NOR2_X1    g08309(.A1(new_n2491_), .A2(new_n10909_), .ZN(new_n11180_));
  INV_X1     g08310(.I(new_n11180_), .ZN(new_n11181_));
  OAI21_X1   g08311(.A1(new_n11181_), .A2(new_n3154_), .B(new_n5987_), .ZN(new_n11182_));
  NOR2_X1    g08312(.A1(new_n11179_), .A2(new_n11182_), .ZN(new_n11183_));
  AOI22_X1   g08313(.A1(new_n11155_), .A2(new_n10907_), .B1(new_n11175_), .B2(new_n11183_), .ZN(new_n11184_));
  MUX2_X1    g08314(.I0(new_n10727_), .I1(new_n10579_), .S(pi0189), .Z(new_n11185_));
  OAI21_X1   g08315(.A1(new_n11185_), .A2(pi0178), .B(new_n11046_), .ZN(new_n11186_));
  NOR4_X1    g08316(.A1(new_n10577_), .A2(new_n7345_), .A3(pi0181), .A4(new_n8896_), .ZN(new_n11187_));
  NOR2_X1    g08317(.A1(new_n11187_), .A2(new_n8914_), .ZN(new_n11188_));
  NAND3_X1   g08318(.A1(new_n11025_), .A2(new_n7345_), .A3(pi0189), .ZN(new_n11189_));
  OAI21_X1   g08319(.A1(new_n11063_), .A2(new_n8872_), .B(new_n7345_), .ZN(new_n11190_));
  AOI21_X1   g08320(.A1(new_n5325_), .A2(new_n11189_), .B(new_n11190_), .ZN(new_n11191_));
  OAI21_X1   g08321(.A1(new_n11060_), .A2(new_n8872_), .B(new_n11191_), .ZN(new_n11192_));
  AOI21_X1   g08322(.A1(new_n11186_), .A2(new_n11188_), .B(new_n11192_), .ZN(new_n11193_));
  AOI21_X1   g08323(.A1(new_n11060_), .A2(new_n11063_), .B(new_n4549_), .ZN(new_n11194_));
  OAI21_X1   g08324(.A1(new_n10549_), .A2(new_n7928_), .B(new_n2526_), .ZN(new_n11195_));
  NAND3_X1   g08325(.A1(new_n10730_), .A2(new_n4549_), .A3(new_n11195_), .ZN(new_n11196_));
  NAND2_X1   g08326(.A1(new_n11196_), .A2(new_n10117_), .ZN(new_n11197_));
  AOI21_X1   g08327(.A1(new_n11194_), .A2(pi0153), .B(new_n11197_), .ZN(new_n11198_));
  NAND2_X1   g08328(.A1(new_n11047_), .A2(new_n4549_), .ZN(new_n11199_));
  NOR3_X1    g08329(.A1(new_n10551_), .A2(pi0153), .A3(new_n11172_), .ZN(new_n11200_));
  AOI21_X1   g08330(.A1(pi0166), .A2(new_n10683_), .B(new_n10550_), .ZN(new_n11201_));
  OAI21_X1   g08331(.A1(new_n11201_), .A2(new_n2526_), .B(pi0157), .ZN(new_n11202_));
  OAI21_X1   g08332(.A1(new_n11202_), .A2(new_n11200_), .B(new_n7593_), .ZN(new_n11203_));
  NOR2_X1    g08333(.A1(new_n10543_), .A2(pi0166), .ZN(new_n11204_));
  INV_X1     g08334(.I(new_n11204_), .ZN(new_n11205_));
  OAI21_X1   g08335(.A1(new_n11053_), .A2(new_n4549_), .B(new_n11205_), .ZN(new_n11206_));
  NAND4_X1   g08336(.A1(new_n10530_), .A2(pi0166), .A3(new_n11052_), .A4(new_n11204_), .ZN(new_n11207_));
  NAND3_X1   g08337(.A1(new_n11206_), .A2(new_n2526_), .A3(new_n11207_), .ZN(new_n11208_));
  NAND3_X1   g08338(.A1(new_n11049_), .A2(pi0153), .A3(pi0166), .ZN(new_n11209_));
  AOI21_X1   g08339(.A1(new_n10117_), .A2(new_n11208_), .B(new_n11209_), .ZN(new_n11210_));
  NAND3_X1   g08340(.A1(new_n11199_), .A2(new_n11203_), .A3(new_n11210_), .ZN(new_n11211_));
  AOI21_X1   g08341(.A1(new_n11028_), .A2(pi0166), .B(new_n11204_), .ZN(new_n11212_));
  INV_X1     g08342(.I(new_n11028_), .ZN(new_n11213_));
  NOR3_X1    g08343(.A1(new_n11213_), .A2(new_n4549_), .A3(new_n11205_), .ZN(new_n11214_));
  NOR3_X1    g08344(.A1(new_n11214_), .A2(pi0153), .A3(new_n11212_), .ZN(new_n11215_));
  NOR2_X1    g08345(.A1(new_n11026_), .A2(pi0166), .ZN(new_n11216_));
  OR4_X2     g08346(.A1(new_n2526_), .A2(new_n7401_), .A3(pi0157), .A4(new_n4549_), .Z(new_n11217_));
  NOR4_X1    g08347(.A1(new_n11215_), .A2(new_n11025_), .A3(new_n11216_), .A4(new_n11217_), .ZN(new_n11218_));
  NAND2_X1   g08348(.A1(new_n11211_), .A2(new_n11218_), .ZN(new_n11219_));
  NOR3_X1    g08349(.A1(new_n11193_), .A2(new_n11198_), .A3(new_n11219_), .ZN(new_n11220_));
  AOI21_X1   g08350(.A1(new_n8011_), .A2(new_n10549_), .B(new_n10612_), .ZN(new_n11221_));
  NOR3_X1    g08351(.A1(new_n10611_), .A2(new_n8012_), .A3(new_n10549_), .ZN(new_n11222_));
  NAND2_X1   g08352(.A1(new_n7345_), .A2(pi0181), .ZN(new_n11225_));
  NOR3_X1    g08353(.A1(new_n11221_), .A2(new_n11222_), .A3(new_n11225_), .ZN(new_n11226_));
  OAI21_X1   g08354(.A1(new_n11053_), .A2(new_n8872_), .B(new_n7345_), .ZN(new_n11227_));
  NAND2_X1   g08355(.A1(new_n11072_), .A2(new_n11227_), .ZN(new_n11228_));
  AOI21_X1   g08356(.A1(new_n10727_), .A2(new_n8872_), .B(new_n11228_), .ZN(new_n11229_));
  NAND2_X1   g08357(.A1(new_n11138_), .A2(pi0178), .ZN(new_n11230_));
  NOR2_X1    g08358(.A1(new_n10552_), .A2(new_n8872_), .ZN(new_n11231_));
  OAI21_X1   g08359(.A1(new_n11230_), .A2(new_n11231_), .B(pi0181), .ZN(new_n11232_));
  NOR2_X1    g08360(.A1(new_n11232_), .A2(new_n11229_), .ZN(new_n11233_));
  OAI22_X1   g08361(.A1(new_n11226_), .A2(new_n11233_), .B1(pi0175), .B2(pi0299), .ZN(new_n11234_));
  OAI21_X1   g08362(.A1(new_n11220_), .A2(new_n11234_), .B(pi0232), .ZN(new_n11235_));
  INV_X1     g08363(.I(new_n10654_), .ZN(new_n11236_));
  NOR4_X1    g08364(.A1(new_n11236_), .A2(new_n5326_), .A3(pi0189), .A4(new_n10985_), .ZN(new_n11237_));
  INV_X1     g08365(.I(new_n10995_), .ZN(new_n11238_));
  NOR3_X1    g08366(.A1(new_n10993_), .A2(new_n8872_), .A3(new_n11238_), .ZN(new_n11239_));
  AOI21_X1   g08367(.A1(pi0189), .A2(new_n11238_), .B(new_n10994_), .ZN(new_n11240_));
  OAI21_X1   g08368(.A1(new_n11240_), .A2(new_n11239_), .B(new_n5326_), .ZN(new_n11241_));
  MUX2_X1    g08369(.I0(new_n10990_), .I1(new_n10984_), .S(new_n8872_), .Z(new_n11242_));
  OAI21_X1   g08370(.A1(new_n5326_), .A2(new_n11242_), .B(new_n11241_), .ZN(new_n11243_));
  AOI22_X1   g08371(.A1(new_n11243_), .A2(new_n8914_), .B1(new_n8871_), .B2(new_n11237_), .ZN(new_n11244_));
  MUX2_X1    g08372(.I0(new_n11020_), .I1(new_n10985_), .S(new_n2587_), .Z(new_n11245_));
  OAI21_X1   g08373(.A1(new_n11245_), .A2(pi0232), .B(pi0039), .ZN(new_n11246_));
  OAI21_X1   g08374(.A1(new_n10651_), .A2(pi0166), .B(new_n11236_), .ZN(new_n11247_));
  NAND3_X1   g08375(.A1(new_n10651_), .A2(new_n4549_), .A3(new_n10654_), .ZN(new_n11248_));
  NAND2_X1   g08376(.A1(new_n11128_), .A2(pi0160), .ZN(new_n11249_));
  AOI21_X1   g08377(.A1(new_n11247_), .A2(new_n11248_), .B(new_n11249_), .ZN(new_n11250_));
  NOR4_X1    g08378(.A1(new_n10638_), .A2(pi0153), .A3(new_n4549_), .A4(new_n10664_), .ZN(new_n11251_));
  AOI21_X1   g08379(.A1(new_n10633_), .A2(new_n7928_), .B(new_n10641_), .ZN(new_n11252_));
  NOR3_X1    g08380(.A1(new_n10633_), .A2(new_n8163_), .A3(new_n10640_), .ZN(new_n11253_));
  NOR3_X1    g08381(.A1(new_n11253_), .A2(new_n11252_), .A3(pi0153), .ZN(new_n11254_));
  OAI21_X1   g08382(.A1(new_n11251_), .A2(new_n11254_), .B(new_n5338_), .ZN(new_n11255_));
  AOI21_X1   g08383(.A1(new_n11110_), .A2(pi0299), .B(new_n7170_), .ZN(new_n11256_));
  OAI21_X1   g08384(.A1(new_n11250_), .A2(new_n11255_), .B(new_n11256_), .ZN(new_n11257_));
  NAND3_X1   g08385(.A1(new_n11257_), .A2(new_n5987_), .A3(new_n11246_), .ZN(new_n11258_));
  OAI21_X1   g08386(.A1(new_n11244_), .A2(new_n11258_), .B(new_n11103_), .ZN(new_n11259_));
  AOI21_X1   g08387(.A1(new_n11235_), .A2(new_n10979_), .B(new_n11259_), .ZN(new_n11260_));
  OAI21_X1   g08388(.A1(new_n11260_), .A2(new_n2622_), .B(new_n11103_), .ZN(new_n11261_));
  NAND2_X1   g08389(.A1(new_n10683_), .A2(new_n8872_), .ZN(new_n11262_));
  NAND2_X1   g08390(.A1(new_n10543_), .A2(pi0175), .ZN(new_n11263_));
  NAND4_X1   g08391(.A1(new_n11172_), .A2(new_n7348_), .A3(new_n11262_), .A4(new_n11263_), .ZN(new_n11264_));
  NAND2_X1   g08392(.A1(new_n2541_), .A2(new_n10505_), .ZN(new_n11265_));
  OAI21_X1   g08393(.A1(new_n11265_), .A2(new_n11103_), .B(new_n2622_), .ZN(new_n11266_));
  NOR2_X1    g08394(.A1(new_n11264_), .A2(new_n11266_), .ZN(new_n11267_));
  OAI21_X1   g08395(.A1(new_n11184_), .A2(new_n11261_), .B(new_n11267_), .ZN(new_n11268_));
  NAND2_X1   g08396(.A1(new_n11264_), .A2(new_n3230_), .ZN(new_n11269_));
  NAND2_X1   g08397(.A1(new_n11269_), .A2(new_n3177_), .ZN(new_n11270_));
  MUX2_X1    g08398(.I0(pi0185), .I1(pi0150), .S(pi0299), .Z(new_n11271_));
  AOI22_X1   g08399(.A1(new_n11103_), .A2(new_n10506_), .B1(new_n11097_), .B2(new_n11271_), .ZN(new_n11272_));
  AOI21_X1   g08400(.A1(new_n11270_), .A2(new_n11272_), .B(po1038), .ZN(new_n11273_));
  AOI21_X1   g08401(.A1(new_n11268_), .A2(new_n11273_), .B(new_n11114_), .ZN(po0283));
  NAND2_X1   g08402(.A1(new_n2548_), .A2(new_n7034_), .ZN(new_n11275_));
  NOR2_X1    g08403(.A1(new_n11275_), .A2(new_n3503_), .ZN(new_n11276_));
  NOR2_X1    g08404(.A1(new_n11276_), .A2(new_n5205_), .ZN(new_n11277_));
  NAND4_X1   g08405(.A1(new_n5875_), .A2(new_n3202_), .A3(pi0129), .A4(new_n5226_), .ZN(new_n11278_));
  INV_X1     g08406(.I(new_n8563_), .ZN(new_n11279_));
  NOR2_X1    g08407(.A1(new_n11279_), .A2(new_n3214_), .ZN(new_n11280_));
  AOI21_X1   g08408(.A1(new_n7034_), .A2(new_n11280_), .B(new_n6963_), .ZN(new_n11281_));
  NAND4_X1   g08409(.A1(new_n5875_), .A2(pi0055), .A3(pi0129), .A4(new_n3229_), .ZN(new_n11282_));
  NAND2_X1   g08410(.A1(new_n11282_), .A2(new_n2533_), .ZN(new_n11283_));
  AOI21_X1   g08411(.A1(new_n11278_), .A2(new_n11281_), .B(new_n11283_), .ZN(new_n11284_));
  XNOR2_X1   g08412(.A1(pi0056), .A2(pi0062), .ZN(new_n11285_));
  NOR2_X1    g08413(.A1(new_n11275_), .A2(new_n11285_), .ZN(new_n11286_));
  NOR2_X1    g08414(.A1(new_n11284_), .A2(new_n11286_), .ZN(new_n11287_));
  NAND2_X1   g08415(.A1(new_n11284_), .A2(new_n11286_), .ZN(new_n11288_));
  NAND2_X1   g08416(.A1(new_n11288_), .A2(pi0059), .ZN(new_n11289_));
  NOR2_X1    g08417(.A1(new_n11289_), .A2(new_n11287_), .ZN(new_n11290_));
  XOR2_X1    g08418(.A1(new_n11290_), .A2(new_n11276_), .Z(new_n11291_));
  NAND2_X1   g08419(.A1(new_n11291_), .A2(new_n5055_), .ZN(new_n11292_));
  XNOR2_X1   g08420(.A1(new_n11292_), .A2(new_n11277_), .ZN(po0284));
  INV_X1     g08421(.I(new_n5057_), .ZN(new_n11294_));
  NOR2_X1    g08422(.A1(new_n5889_), .A2(new_n5198_), .ZN(new_n11295_));
  NAND3_X1   g08423(.A1(new_n3379_), .A2(pi0038), .A3(new_n5153_), .ZN(new_n11296_));
  OAI21_X1   g08424(.A1(new_n3172_), .A2(new_n5153_), .B(new_n3524_), .ZN(new_n11297_));
  AOI21_X1   g08425(.A1(new_n11297_), .A2(new_n11296_), .B(pi0100), .ZN(new_n11298_));
  INV_X1     g08426(.I(new_n5192_), .ZN(new_n11299_));
  NAND2_X1   g08427(.A1(new_n5160_), .A2(new_n5185_), .ZN(new_n11300_));
  NAND4_X1   g08428(.A1(new_n11299_), .A2(new_n3177_), .A3(new_n5410_), .A4(new_n11300_), .ZN(new_n11301_));
  AOI21_X1   g08429(.A1(new_n5879_), .A2(new_n3203_), .B(new_n3214_), .ZN(new_n11302_));
  NOR2_X1    g08430(.A1(new_n11302_), .A2(new_n5880_), .ZN(new_n11303_));
  OAI21_X1   g08431(.A1(new_n11298_), .A2(new_n11301_), .B(new_n11303_), .ZN(new_n11304_));
  AOI21_X1   g08432(.A1(new_n11304_), .A2(new_n6962_), .B(new_n11295_), .ZN(new_n11305_));
  OAI21_X1   g08433(.A1(new_n11305_), .A2(pi0056), .B(new_n11294_), .ZN(new_n11306_));
  AOI21_X1   g08434(.A1(new_n5056_), .A2(new_n3341_), .B(new_n3240_), .ZN(new_n11307_));
  NOR2_X1    g08435(.A1(new_n11307_), .A2(pi0062), .ZN(new_n11308_));
  NAND2_X1   g08436(.A1(new_n5209_), .A2(new_n2571_), .ZN(new_n11309_));
  AOI21_X1   g08437(.A1(new_n11306_), .A2(new_n11308_), .B(new_n11309_), .ZN(po0286));
  AOI21_X1   g08438(.A1(new_n10683_), .A2(pi0169), .B(pi0051), .ZN(new_n11311_));
  NAND2_X1   g08439(.A1(new_n11311_), .A2(new_n3177_), .ZN(new_n11312_));
  INV_X1     g08440(.I(new_n11102_), .ZN(new_n11313_));
  NOR2_X1    g08441(.A1(new_n11313_), .A2(pi0126), .ZN(new_n11314_));
  INV_X1     g08442(.I(new_n11314_), .ZN(new_n11315_));
  NOR2_X1    g08443(.A1(new_n11315_), .A2(pi0132), .ZN(new_n11316_));
  INV_X1     g08444(.I(new_n11316_), .ZN(new_n11317_));
  NOR4_X1    g08445(.A1(new_n11317_), .A2(pi0130), .A3(pi0134), .A4(new_n10497_), .ZN(new_n11318_));
  NAND4_X1   g08446(.A1(new_n10577_), .A2(new_n3177_), .A3(pi0169), .A4(new_n5988_), .ZN(new_n11319_));
  NAND4_X1   g08447(.A1(new_n6845_), .A2(new_n3177_), .A3(pi0167), .A4(new_n5988_), .ZN(new_n11320_));
  NAND4_X1   g08448(.A1(new_n11312_), .A2(new_n11318_), .A3(new_n11319_), .A4(new_n11320_), .ZN(new_n11321_));
  INV_X1     g08449(.I(new_n11318_), .ZN(new_n11322_));
  INV_X1     g08450(.I(new_n10987_), .ZN(new_n11323_));
  NAND3_X1   g08451(.A1(new_n10643_), .A2(new_n2658_), .A3(new_n10649_), .ZN(new_n11324_));
  MUX2_X1    g08452(.I0(new_n11324_), .I1(new_n11323_), .S(new_n4272_), .Z(new_n11325_));
  NAND2_X1   g08453(.A1(new_n7170_), .A2(pi0162), .ZN(new_n11329_));
  NOR2_X1    g08454(.A1(new_n11325_), .A2(new_n11329_), .ZN(new_n11330_));
  OAI21_X1   g08455(.A1(new_n11245_), .A2(pi0051), .B(new_n5987_), .ZN(new_n11331_));
  INV_X1     g08456(.I(new_n11331_), .ZN(new_n11332_));
  NOR2_X1    g08457(.A1(new_n10985_), .A2(pi0051), .ZN(new_n11333_));
  NOR3_X1    g08458(.A1(new_n11333_), .A2(new_n7339_), .A3(new_n7137_), .ZN(new_n11334_));
  INV_X1     g08459(.I(new_n7138_), .ZN(new_n11335_));
  NOR2_X1    g08460(.A1(new_n5989_), .A2(new_n11335_), .ZN(new_n11336_));
  NOR3_X1    g08461(.A1(new_n11336_), .A2(new_n5525_), .A3(new_n10577_), .ZN(new_n11337_));
  AOI21_X1   g08462(.A1(pi0191), .A2(new_n2587_), .B(new_n7339_), .ZN(new_n11338_));
  AOI21_X1   g08463(.A1(new_n10648_), .A2(new_n11338_), .B(new_n5987_), .ZN(new_n11339_));
  OAI21_X1   g08464(.A1(new_n11337_), .A2(pi0100), .B(new_n11339_), .ZN(new_n11340_));
  AOI21_X1   g08465(.A1(new_n11334_), .A2(new_n10988_), .B(new_n11340_), .ZN(new_n11341_));
  OAI21_X1   g08466(.A1(new_n11332_), .A2(new_n8533_), .B(new_n11341_), .ZN(new_n11342_));
  NOR2_X1    g08467(.A1(new_n11336_), .A2(new_n10577_), .ZN(new_n11343_));
  NOR2_X1    g08468(.A1(new_n11104_), .A2(new_n11343_), .ZN(new_n11344_));
  AOI21_X1   g08469(.A1(new_n11344_), .A2(pi0100), .B(new_n2541_), .ZN(new_n11345_));
  NOR3_X1    g08470(.A1(new_n11345_), .A2(new_n3173_), .A3(new_n10505_), .ZN(new_n11346_));
  OAI21_X1   g08471(.A1(new_n11342_), .A2(new_n11330_), .B(new_n11346_), .ZN(new_n11347_));
  NOR2_X1    g08472(.A1(new_n11344_), .A2(new_n3229_), .ZN(new_n11348_));
  NOR2_X1    g08473(.A1(new_n11348_), .A2(pi0087), .ZN(new_n11349_));
  AOI21_X1   g08474(.A1(pi0087), .A2(new_n7358_), .B(new_n11349_), .ZN(new_n11350_));
  NAND2_X1   g08475(.A1(new_n11350_), .A2(new_n10507_), .ZN(new_n11351_));
  AOI21_X1   g08476(.A1(new_n11347_), .A2(new_n11322_), .B(new_n11351_), .ZN(new_n11352_));
  AOI21_X1   g08477(.A1(new_n5109_), .A2(new_n10640_), .B(new_n10862_), .ZN(new_n11353_));
  NOR2_X1    g08478(.A1(new_n11353_), .A2(pi0224), .ZN(new_n11354_));
  AOI21_X1   g08479(.A1(pi0051), .A2(new_n5109_), .B(new_n11163_), .ZN(new_n11355_));
  INV_X1     g08480(.I(new_n11355_), .ZN(new_n11356_));
  NOR2_X1    g08481(.A1(new_n11356_), .A2(new_n2595_), .ZN(new_n11357_));
  OAI21_X1   g08482(.A1(new_n11357_), .A2(new_n11354_), .B(new_n6050_), .ZN(new_n11358_));
  OAI21_X1   g08483(.A1(new_n6050_), .A2(new_n11105_), .B(new_n11358_), .ZN(new_n11359_));
  INV_X1     g08484(.I(new_n11359_), .ZN(new_n11360_));
  INV_X1     g08485(.I(pi0191), .ZN(new_n11361_));
  INV_X1     g08486(.I(new_n11353_), .ZN(new_n11362_));
  NOR2_X1    g08487(.A1(new_n11105_), .A2(new_n6462_), .ZN(new_n11363_));
  AOI21_X1   g08488(.A1(new_n11362_), .A2(new_n6462_), .B(new_n11363_), .ZN(new_n11364_));
  INV_X1     g08489(.I(new_n11364_), .ZN(new_n11365_));
  OAI22_X1   g08490(.A1(new_n11365_), .A2(pi0140), .B1(new_n11361_), .B2(pi0299), .ZN(new_n11366_));
  AOI21_X1   g08491(.A1(new_n11360_), .A2(pi0140), .B(new_n11366_), .ZN(new_n11367_));
  AOI21_X1   g08492(.A1(new_n7325_), .A2(pi0216), .B(new_n5357_), .ZN(new_n11368_));
  NOR2_X1    g08493(.A1(new_n11311_), .A2(new_n11368_), .ZN(new_n11369_));
  NOR2_X1    g08494(.A1(new_n11369_), .A2(new_n5356_), .ZN(new_n11370_));
  AOI21_X1   g08495(.A1(new_n10870_), .A2(new_n10639_), .B(pi0051), .ZN(new_n11371_));
  NOR2_X1    g08496(.A1(new_n11371_), .A2(new_n7339_), .ZN(new_n11372_));
  AOI21_X1   g08497(.A1(new_n10639_), .A2(new_n6462_), .B(pi0051), .ZN(new_n11373_));
  OAI22_X1   g08498(.A1(new_n11373_), .A2(pi0140), .B1(pi0191), .B2(pi0299), .ZN(new_n11374_));
  OAI22_X1   g08499(.A1(new_n11372_), .A2(new_n11374_), .B1(new_n2587_), .B2(new_n11370_), .ZN(new_n11375_));
  OAI21_X1   g08500(.A1(new_n11367_), .A2(new_n11375_), .B(pi0232), .ZN(new_n11376_));
  NOR2_X1    g08501(.A1(new_n10774_), .A2(new_n10909_), .ZN(new_n11377_));
  NOR2_X1    g08502(.A1(new_n11377_), .A2(pi0051), .ZN(new_n11378_));
  NOR2_X1    g08503(.A1(new_n11378_), .A2(new_n5864_), .ZN(new_n11379_));
  NAND2_X1   g08504(.A1(new_n11376_), .A2(new_n11379_), .ZN(new_n11380_));
  NOR2_X1    g08505(.A1(new_n10535_), .A2(new_n5109_), .ZN(new_n11381_));
  AOI21_X1   g08506(.A1(new_n10614_), .A2(new_n5109_), .B(new_n11381_), .ZN(new_n11382_));
  MUX2_X1    g08507(.I0(new_n11382_), .I1(new_n10613_), .S(new_n11335_), .Z(new_n11383_));
  AOI21_X1   g08508(.A1(new_n10614_), .A2(new_n5987_), .B(pi0039), .ZN(new_n11384_));
  OAI21_X1   g08509(.A1(new_n11383_), .A2(new_n5987_), .B(new_n11384_), .ZN(new_n11385_));
  NAND2_X1   g08510(.A1(new_n11385_), .A2(new_n11380_), .ZN(new_n11386_));
  MUX2_X1    g08511(.I0(new_n11386_), .I1(new_n11344_), .S(pi0038), .Z(new_n11387_));
  NOR2_X1    g08512(.A1(new_n2540_), .A2(pi0100), .ZN(new_n11388_));
  NAND2_X1   g08513(.A1(new_n11387_), .A2(new_n11388_), .ZN(new_n11389_));
  NOR2_X1    g08514(.A1(new_n11350_), .A2(new_n11322_), .ZN(new_n11390_));
  AOI21_X1   g08515(.A1(new_n11389_), .A2(new_n11390_), .B(new_n11352_), .ZN(new_n11391_));
  OAI21_X1   g08516(.A1(new_n11391_), .A2(po1038), .B(new_n11321_), .ZN(po0287));
  AND3_X2    g08517(.A1(new_n10246_), .A2(pi0100), .A3(new_n5872_), .Z(new_n11393_));
  AOI21_X1   g08518(.A1(pi0100), .A2(new_n5873_), .B(new_n10246_), .ZN(new_n11394_));
  OAI21_X1   g08519(.A1(new_n11393_), .A2(new_n11394_), .B(new_n2534_), .ZN(new_n11395_));
  AOI21_X1   g08520(.A1(new_n5875_), .A2(pi0075), .B(pi0092), .ZN(new_n11396_));
  OR3_X2     g08521(.A1(new_n5880_), .A2(pi0054), .A3(new_n6965_), .Z(new_n11397_));
  AOI21_X1   g08522(.A1(new_n11395_), .A2(new_n11396_), .B(new_n11397_), .ZN(po0288));
  INV_X1     g08523(.I(new_n10605_), .ZN(new_n11399_));
  NAND3_X1   g08524(.A1(new_n10592_), .A2(new_n5108_), .A3(new_n11399_), .ZN(new_n11400_));
  OAI21_X1   g08525(.A1(new_n5109_), .A2(new_n11399_), .B(new_n10591_), .ZN(new_n11401_));
  AOI21_X1   g08526(.A1(new_n11400_), .A2(new_n11401_), .B(new_n5326_), .ZN(new_n11402_));
  NAND2_X1   g08527(.A1(new_n10591_), .A2(new_n5109_), .ZN(new_n11403_));
  OAI21_X1   g08528(.A1(new_n10539_), .A2(new_n10597_), .B(new_n11403_), .ZN(new_n11404_));
  NAND2_X1   g08529(.A1(new_n11404_), .A2(pi0182), .ZN(new_n11405_));
  NOR2_X1    g08530(.A1(new_n10591_), .A2(new_n5108_), .ZN(new_n11406_));
  OAI21_X1   g08531(.A1(new_n10615_), .A2(new_n11406_), .B(pi0182), .ZN(new_n11407_));
  AOI21_X1   g08532(.A1(new_n11407_), .A2(new_n11405_), .B(new_n10056_), .ZN(new_n11408_));
  NOR2_X1    g08533(.A1(new_n10592_), .A2(pi0182), .ZN(new_n11409_));
  NOR2_X1    g08534(.A1(pi0190), .A2(pi0299), .ZN(new_n11410_));
  INV_X1     g08535(.I(new_n11410_), .ZN(new_n11411_));
  NAND2_X1   g08536(.A1(new_n11411_), .A2(new_n10056_), .ZN(new_n11412_));
  NOR4_X1    g08537(.A1(new_n11408_), .A2(new_n11402_), .A3(new_n11409_), .A4(new_n11412_), .ZN(new_n11413_));
  NAND2_X1   g08538(.A1(new_n11404_), .A2(new_n4413_), .ZN(new_n11414_));
  INV_X1     g08539(.I(new_n11406_), .ZN(new_n11415_));
  OAI21_X1   g08540(.A1(new_n11399_), .A2(pi0151), .B(new_n4413_), .ZN(new_n11416_));
  NOR2_X1    g08541(.A1(new_n2658_), .A2(pi0151), .ZN(new_n11417_));
  INV_X1     g08542(.I(new_n11417_), .ZN(new_n11418_));
  NAND2_X1   g08543(.A1(new_n5109_), .A2(new_n4413_), .ZN(new_n11419_));
  AOI21_X1   g08544(.A1(new_n10618_), .A2(new_n11418_), .B(new_n11419_), .ZN(new_n11420_));
  NOR3_X1    g08545(.A1(new_n11420_), .A2(new_n3417_), .A3(pi0160), .ZN(new_n11421_));
  NAND4_X1   g08546(.A1(new_n10613_), .A2(new_n11415_), .A3(new_n11416_), .A4(new_n11421_), .ZN(new_n11422_));
  NOR3_X1    g08547(.A1(new_n11406_), .A2(new_n4413_), .A3(new_n10918_), .ZN(new_n11423_));
  OAI21_X1   g08548(.A1(new_n10584_), .A2(new_n4413_), .B(new_n3417_), .ZN(new_n11424_));
  NAND3_X1   g08549(.A1(new_n10591_), .A2(new_n10089_), .A3(new_n11424_), .ZN(new_n11425_));
  NAND4_X1   g08550(.A1(new_n11425_), .A2(pi0151), .A3(new_n5338_), .A4(new_n2587_), .ZN(new_n11426_));
  NOR2_X1    g08551(.A1(new_n11426_), .A2(new_n11423_), .ZN(new_n11427_));
  NAND3_X1   g08552(.A1(new_n11427_), .A2(new_n11414_), .A3(new_n11422_), .ZN(new_n11428_));
  AOI21_X1   g08553(.A1(pi0051), .A2(new_n10056_), .B(new_n5109_), .ZN(new_n11429_));
  NOR3_X1    g08554(.A1(new_n10517_), .A2(new_n5326_), .A3(new_n11429_), .ZN(new_n11430_));
  AOI21_X1   g08555(.A1(new_n10534_), .A2(new_n11430_), .B(new_n10107_), .ZN(new_n11431_));
  AOI21_X1   g08556(.A1(new_n11403_), .A2(new_n11431_), .B(new_n5987_), .ZN(new_n11432_));
  NAND2_X1   g08557(.A1(new_n11428_), .A2(new_n11432_), .ZN(new_n11433_));
  OAI22_X1   g08558(.A1(new_n11413_), .A2(new_n11433_), .B1(pi0232), .B2(new_n10592_), .ZN(new_n11434_));
  NAND2_X1   g08559(.A1(new_n11434_), .A2(new_n3154_), .ZN(new_n11435_));
  OAI21_X1   g08560(.A1(pi0168), .A2(new_n10891_), .B(new_n10864_), .ZN(new_n11436_));
  NAND3_X1   g08561(.A1(new_n10863_), .A2(new_n4413_), .A3(new_n10891_), .ZN(new_n11437_));
  NAND3_X1   g08562(.A1(new_n11436_), .A2(new_n11418_), .A3(new_n11437_), .ZN(new_n11438_));
  NOR3_X1    g08563(.A1(new_n10676_), .A2(pi0168), .A3(new_n11166_), .ZN(new_n11439_));
  AOI21_X1   g08564(.A1(new_n4413_), .A2(new_n11166_), .B(new_n10677_), .ZN(new_n11440_));
  INV_X1     g08565(.I(new_n10869_), .ZN(new_n11441_));
  NOR4_X1    g08566(.A1(new_n11440_), .A2(new_n7067_), .A3(pi0151), .A4(new_n11439_), .ZN(new_n11443_));
  MUX2_X1    g08567(.I0(new_n11443_), .I1(new_n11438_), .S(new_n2562_), .Z(new_n11444_));
  AND2_X2    g08568(.A1(new_n11444_), .A2(new_n5356_), .Z(new_n11445_));
  AOI21_X1   g08569(.A1(new_n10089_), .A2(new_n10544_), .B(new_n11417_), .ZN(new_n11446_));
  NAND2_X1   g08570(.A1(new_n11446_), .A2(new_n10546_), .ZN(new_n11447_));
  INV_X1     g08571(.I(new_n11447_), .ZN(new_n11448_));
  NOR4_X1    g08572(.A1(new_n11448_), .A2(pi0149), .A3(new_n2562_), .A4(new_n5356_), .ZN(new_n11449_));
  AOI21_X1   g08573(.A1(new_n10853_), .A2(new_n7180_), .B(pi0173), .ZN(new_n11450_));
  OAI21_X1   g08574(.A1(new_n10856_), .A2(new_n7180_), .B(new_n11450_), .ZN(new_n11451_));
  OAI21_X1   g08575(.A1(new_n10863_), .A2(new_n6559_), .B(new_n7180_), .ZN(new_n11452_));
  NOR2_X1    g08576(.A1(new_n10867_), .A2(new_n10056_), .ZN(new_n11453_));
  NAND2_X1   g08577(.A1(new_n10878_), .A2(new_n7180_), .ZN(new_n11454_));
  NAND2_X1   g08578(.A1(new_n11454_), .A2(new_n10107_), .ZN(new_n11455_));
  AOI21_X1   g08579(.A1(new_n11453_), .A2(new_n11452_), .B(new_n11455_), .ZN(new_n11456_));
  NAND2_X1   g08580(.A1(new_n10056_), .A2(pi0183), .ZN(new_n11457_));
  AOI21_X1   g08581(.A1(new_n6559_), .A2(new_n7180_), .B(pi0173), .ZN(new_n11458_));
  AOI21_X1   g08582(.A1(new_n10859_), .A2(new_n11458_), .B(new_n11411_), .ZN(new_n11459_));
  OAI21_X1   g08583(.A1(new_n10874_), .A2(new_n11457_), .B(new_n11459_), .ZN(new_n11460_));
  AOI21_X1   g08584(.A1(new_n11451_), .A2(new_n11456_), .B(new_n11460_), .ZN(new_n11461_));
  OAI21_X1   g08585(.A1(new_n11445_), .A2(new_n11449_), .B(new_n11461_), .ZN(new_n11462_));
  NOR2_X1    g08586(.A1(new_n5987_), .A2(pi0039), .ZN(new_n11463_));
  AOI21_X1   g08587(.A1(new_n11462_), .A2(new_n11463_), .B(new_n2622_), .ZN(new_n11464_));
  INV_X1     g08588(.I(new_n7348_), .ZN(new_n11465_));
  NOR2_X1    g08589(.A1(new_n10897_), .A2(new_n10096_), .ZN(new_n11466_));
  NOR2_X1    g08590(.A1(new_n10544_), .A2(new_n10056_), .ZN(new_n11467_));
  NOR4_X1    g08591(.A1(new_n11466_), .A2(new_n11465_), .A3(new_n11447_), .A4(new_n11467_), .ZN(new_n11468_));
  INV_X1     g08592(.I(new_n11468_), .ZN(new_n11469_));
  NAND3_X1   g08593(.A1(new_n11469_), .A2(new_n2541_), .A3(new_n2621_), .ZN(new_n11470_));
  AOI21_X1   g08594(.A1(new_n11435_), .A2(new_n11464_), .B(new_n11470_), .ZN(new_n11471_));
  AND2_X2    g08595(.A1(new_n11316_), .A2(new_n10498_), .Z(new_n11472_));
  AOI21_X1   g08596(.A1(pi0132), .A2(new_n11315_), .B(new_n11472_), .ZN(new_n11473_));
  INV_X1     g08597(.I(new_n11473_), .ZN(new_n11474_));
  NAND2_X1   g08598(.A1(new_n7112_), .A2(pi0087), .ZN(new_n11475_));
  NAND2_X1   g08599(.A1(new_n11474_), .A2(new_n11475_), .ZN(new_n11476_));
  NAND3_X1   g08600(.A1(new_n11476_), .A2(new_n10800_), .A3(new_n11468_), .ZN(new_n11477_));
  OAI21_X1   g08601(.A1(new_n10544_), .A2(new_n10056_), .B(new_n11410_), .ZN(new_n11478_));
  NAND4_X1   g08602(.A1(new_n10986_), .A2(pi0183), .A3(new_n10654_), .A4(new_n11478_), .ZN(new_n11479_));
  NOR2_X1    g08603(.A1(new_n7180_), .A2(pi0173), .ZN(new_n11480_));
  AOI21_X1   g08604(.A1(new_n10993_), .A2(new_n10984_), .B(new_n7180_), .ZN(new_n11481_));
  AOI22_X1   g08605(.A1(new_n11481_), .A2(pi0173), .B1(new_n10650_), .B2(new_n11480_), .ZN(new_n11482_));
  OAI21_X1   g08606(.A1(new_n11482_), .A2(new_n10107_), .B(new_n11479_), .ZN(new_n11483_));
  MUX2_X1    g08607(.I0(new_n10663_), .I1(new_n10637_), .S(pi0168), .Z(new_n11484_));
  NOR3_X1    g08608(.A1(new_n10633_), .A2(new_n3417_), .A3(new_n10088_), .ZN(new_n11485_));
  NOR2_X1    g08609(.A1(new_n11485_), .A2(pi0149), .ZN(new_n11486_));
  OAI21_X1   g08610(.A1(new_n11484_), .A2(new_n3417_), .B(new_n11486_), .ZN(new_n11487_));
  AOI21_X1   g08611(.A1(new_n11441_), .A2(new_n11418_), .B(new_n10644_), .ZN(new_n11488_));
  NOR2_X1    g08612(.A1(new_n10654_), .A2(new_n11446_), .ZN(new_n11489_));
  NOR3_X1    g08613(.A1(new_n11489_), .A2(pi0149), .A3(pi0168), .ZN(new_n11490_));
  NOR4_X1    g08614(.A1(new_n11488_), .A2(new_n4413_), .A3(new_n7170_), .A4(new_n11490_), .ZN(new_n11491_));
  OAI21_X1   g08615(.A1(new_n11448_), .A2(new_n10504_), .B(new_n2587_), .ZN(new_n11492_));
  NAND2_X1   g08616(.A1(new_n11492_), .A2(new_n10180_), .ZN(new_n11493_));
  AOI21_X1   g08617(.A1(new_n11491_), .A2(new_n11487_), .B(new_n11493_), .ZN(new_n11494_));
  AOI21_X1   g08618(.A1(new_n11483_), .A2(new_n11494_), .B(new_n5987_), .ZN(new_n11495_));
  OAI21_X1   g08619(.A1(new_n11245_), .A2(pi0232), .B(new_n3154_), .ZN(new_n11496_));
  NAND2_X1   g08620(.A1(pi0151), .A2(pi0168), .ZN(new_n11497_));
  NOR2_X1    g08621(.A1(new_n10753_), .A2(new_n11497_), .ZN(new_n11498_));
  NAND3_X1   g08622(.A1(new_n10543_), .A2(new_n3417_), .A3(new_n4413_), .ZN(new_n11499_));
  OAI22_X1   g08623(.A1(new_n11051_), .A2(pi0160), .B1(new_n10559_), .B2(new_n11499_), .ZN(new_n11500_));
  NOR3_X1    g08624(.A1(new_n11052_), .A2(pi0151), .A3(new_n11448_), .ZN(new_n11501_));
  INV_X1     g08625(.I(new_n11051_), .ZN(new_n11502_));
  NAND2_X1   g08626(.A1(new_n10683_), .A2(new_n4413_), .ZN(new_n11503_));
  AOI21_X1   g08627(.A1(new_n11502_), .A2(new_n11503_), .B(new_n3417_), .ZN(new_n11504_));
  NOR4_X1    g08628(.A1(new_n11501_), .A2(new_n11504_), .A3(new_n5338_), .A4(pi0299), .ZN(new_n11505_));
  OAI21_X1   g08629(.A1(new_n11498_), .A2(new_n11500_), .B(new_n11505_), .ZN(new_n11506_));
  OAI21_X1   g08630(.A1(new_n2658_), .A2(pi0173), .B(new_n11502_), .ZN(new_n11507_));
  NOR3_X1    g08631(.A1(new_n10560_), .A2(pi0182), .A3(new_n10106_), .ZN(new_n11508_));
  NAND4_X1   g08632(.A1(new_n11052_), .A2(pi0182), .A3(new_n10548_), .A4(new_n11478_), .ZN(new_n11509_));
  NAND2_X1   g08633(.A1(new_n11509_), .A2(pi0232), .ZN(new_n11510_));
  AOI21_X1   g08634(.A1(new_n11507_), .A2(new_n11508_), .B(new_n11510_), .ZN(new_n11511_));
  OAI21_X1   g08635(.A1(new_n10548_), .A2(pi0232), .B(new_n3154_), .ZN(new_n11512_));
  AOI21_X1   g08636(.A1(new_n11506_), .A2(new_n11511_), .B(new_n11512_), .ZN(new_n11513_));
  OAI21_X1   g08637(.A1(new_n11495_), .A2(new_n11496_), .B(new_n11513_), .ZN(new_n11514_));
  NAND2_X1   g08638(.A1(new_n2541_), .A2(new_n2622_), .ZN(new_n11515_));
  AOI21_X1   g08639(.A1(new_n11469_), .A2(new_n10505_), .B(new_n11515_), .ZN(new_n11516_));
  NAND2_X1   g08640(.A1(new_n11473_), .A2(new_n11475_), .ZN(new_n11517_));
  AOI21_X1   g08641(.A1(new_n11469_), .A2(new_n10801_), .B(new_n11517_), .ZN(new_n11518_));
  NOR3_X1    g08642(.A1(new_n11518_), .A2(new_n11516_), .A3(new_n2621_), .ZN(new_n11519_));
  OAI21_X1   g08643(.A1(new_n11447_), .A2(new_n5987_), .B(new_n3177_), .ZN(new_n11520_));
  AOI21_X1   g08644(.A1(new_n11473_), .A2(new_n10504_), .B(new_n11520_), .ZN(new_n11521_));
  NAND2_X1   g08645(.A1(new_n11097_), .A2(pi0164), .ZN(new_n11522_));
  OAI21_X1   g08646(.A1(new_n11521_), .A2(new_n11522_), .B(new_n6845_), .ZN(new_n11523_));
  AOI21_X1   g08647(.A1(new_n11514_), .A2(new_n11519_), .B(new_n11523_), .ZN(new_n11524_));
  OAI21_X1   g08648(.A1(new_n11471_), .A2(new_n11477_), .B(new_n11524_), .ZN(po0289));
  INV_X1     g08649(.I(pi0133), .ZN(new_n11526_));
  OAI21_X1   g08650(.A1(new_n10500_), .A2(pi0125), .B(new_n11526_), .ZN(new_n11527_));
  NAND3_X1   g08651(.A1(new_n6845_), .A2(new_n11097_), .A3(pi0149), .ZN(new_n11528_));
  AOI21_X1   g08652(.A1(new_n11527_), .A2(new_n10506_), .B(new_n11528_), .ZN(new_n11529_));
  AOI21_X1   g08653(.A1(new_n5109_), .A2(new_n10562_), .B(new_n10606_), .ZN(new_n11530_));
  AND2_X2    g08654(.A1(new_n11530_), .A2(new_n7114_), .Z(new_n11531_));
  NOR3_X1    g08655(.A1(new_n3271_), .A2(new_n5987_), .A3(new_n2587_), .ZN(new_n11532_));
  INV_X1     g08656(.I(new_n11532_), .ZN(new_n11533_));
  NOR4_X1    g08657(.A1(new_n8625_), .A2(pi0039), .A3(pi0176), .A4(new_n11533_), .ZN(new_n11534_));
  OAI21_X1   g08658(.A1(new_n10563_), .A2(new_n11532_), .B(new_n11534_), .ZN(new_n11535_));
  AOI21_X1   g08659(.A1(new_n3154_), .A2(pi0176), .B(pi0087), .ZN(new_n11536_));
  NAND2_X1   g08660(.A1(new_n11527_), .A2(new_n11536_), .ZN(new_n11537_));
  AOI21_X1   g08661(.A1(new_n10563_), .A2(new_n7115_), .B(new_n11537_), .ZN(new_n11538_));
  OAI21_X1   g08662(.A1(new_n11530_), .A2(new_n11535_), .B(new_n11538_), .ZN(new_n11539_));
  MUX2_X1    g08663(.I0(pi0183), .I1(pi0149), .S(pi0299), .Z(new_n11540_));
  NAND2_X1   g08664(.A1(new_n5988_), .A2(new_n11540_), .ZN(new_n11541_));
  NAND3_X1   g08665(.A1(new_n10505_), .A2(pi0197), .A3(new_n10648_), .ZN(new_n11542_));
  OAI21_X1   g08666(.A1(new_n11019_), .A2(new_n11542_), .B(pi0299), .ZN(new_n11543_));
  NOR2_X1    g08667(.A1(new_n11236_), .A2(new_n5323_), .ZN(new_n11544_));
  NOR3_X1    g08668(.A1(new_n11544_), .A2(pi0299), .A3(new_n10985_), .ZN(new_n11545_));
  AOI21_X1   g08669(.A1(new_n11545_), .A2(new_n11543_), .B(new_n5987_), .ZN(new_n11546_));
  NOR2_X1    g08670(.A1(new_n11246_), .A2(new_n11546_), .ZN(new_n11547_));
  INV_X1     g08671(.I(new_n7117_), .ZN(new_n11548_));
  NAND2_X1   g08672(.A1(new_n11548_), .A2(new_n10697_), .ZN(new_n11549_));
  NOR4_X1    g08673(.A1(new_n2541_), .A2(pi0038), .A3(pi0100), .A4(new_n10504_), .ZN(new_n11550_));
  OAI21_X1   g08674(.A1(new_n10530_), .A2(new_n11549_), .B(new_n11550_), .ZN(new_n11551_));
  OAI22_X1   g08675(.A1(new_n11547_), .A2(new_n11551_), .B1(new_n10504_), .B2(new_n10800_), .ZN(new_n11552_));
  AOI22_X1   g08676(.A1(new_n11552_), .A2(new_n11527_), .B1(pi0087), .B2(new_n11541_), .ZN(new_n11553_));
  OAI21_X1   g08677(.A1(new_n11531_), .A2(new_n11539_), .B(new_n11553_), .ZN(new_n11554_));
  AOI21_X1   g08678(.A1(new_n11554_), .A2(new_n6845_), .B(new_n11529_), .ZN(po0290));
  INV_X1     g08679(.I(pi0134), .ZN(new_n11556_));
  NOR4_X1    g08680(.A1(new_n11315_), .A2(pi0130), .A3(pi0132), .A4(pi0136), .ZN(new_n11557_));
  INV_X1     g08681(.I(new_n11557_), .ZN(new_n11558_));
  NOR2_X1    g08682(.A1(new_n11558_), .A2(pi0135), .ZN(new_n11559_));
  NOR2_X1    g08683(.A1(new_n11559_), .A2(new_n11556_), .ZN(new_n11560_));
  NOR3_X1    g08684(.A1(new_n6845_), .A2(pi0051), .A3(pi0087), .ZN(new_n11561_));
  NOR2_X1    g08685(.A1(new_n5109_), .A2(new_n3842_), .ZN(new_n11562_));
  INV_X1     g08686(.I(new_n11562_), .ZN(new_n11563_));
  OAI21_X1   g08687(.A1(new_n11563_), .A2(new_n5987_), .B(new_n10492_), .ZN(new_n11564_));
  NOR2_X1    g08688(.A1(new_n11561_), .A2(new_n11564_), .ZN(new_n11565_));
  NOR4_X1    g08689(.A1(new_n10577_), .A2(pi0299), .A3(new_n7170_), .A4(new_n11562_), .ZN(new_n11567_));
  INV_X1     g08690(.I(new_n11567_), .ZN(new_n11568_));
  INV_X1     g08691(.I(new_n11333_), .ZN(new_n11569_));
  OAI21_X1   g08692(.A1(new_n11569_), .A2(pi0192), .B(new_n2587_), .ZN(new_n11570_));
  NAND3_X1   g08693(.A1(new_n11570_), .A2(new_n5987_), .A3(new_n11568_), .ZN(new_n11571_));
  INV_X1     g08694(.I(pi0192), .ZN(new_n11572_));
  MUX2_X1    g08695(.I0(new_n11572_), .I1(new_n3842_), .S(pi0299), .Z(new_n11573_));
  NOR2_X1    g08696(.A1(new_n5989_), .A2(new_n11573_), .ZN(new_n11574_));
  NOR2_X1    g08697(.A1(new_n11574_), .A2(new_n10577_), .ZN(new_n11575_));
  AOI21_X1   g08698(.A1(new_n7109_), .A2(pi0039), .B(pi0164), .ZN(new_n11576_));
  OAI21_X1   g08699(.A1(new_n11575_), .A2(pi0039), .B(new_n11576_), .ZN(new_n11577_));
  AOI21_X1   g08700(.A1(new_n11331_), .A2(new_n11571_), .B(new_n11577_), .ZN(new_n11578_));
  NOR2_X1    g08701(.A1(new_n10988_), .A2(new_n11569_), .ZN(new_n11579_));
  AOI21_X1   g08702(.A1(new_n11579_), .A2(new_n11572_), .B(pi0299), .ZN(new_n11580_));
  NOR3_X1    g08703(.A1(new_n11580_), .A2(pi0232), .A3(new_n11567_), .ZN(new_n11581_));
  NAND2_X1   g08704(.A1(pi0039), .A2(pi0186), .ZN(new_n11582_));
  NOR4_X1    g08705(.A1(new_n11578_), .A2(new_n11332_), .A3(new_n11581_), .A4(new_n11582_), .ZN(new_n11583_));
  NOR2_X1    g08706(.A1(new_n11562_), .A2(pi0299), .ZN(new_n11584_));
  NAND3_X1   g08707(.A1(new_n7634_), .A2(new_n10575_), .A3(new_n11584_), .ZN(new_n11587_));
  NAND3_X1   g08708(.A1(new_n11570_), .A2(new_n5987_), .A3(new_n11587_), .ZN(new_n11588_));
  AOI22_X1   g08709(.A1(new_n11331_), .A2(new_n11588_), .B1(pi0039), .B2(new_n7109_), .ZN(new_n11589_));
  NAND2_X1   g08710(.A1(new_n11587_), .A2(new_n5987_), .ZN(new_n11590_));
  NOR2_X1    g08711(.A1(new_n11580_), .A2(new_n11590_), .ZN(new_n11591_));
  NAND3_X1   g08712(.A1(new_n7058_), .A2(pi0039), .A3(pi0186), .ZN(new_n11592_));
  NOR4_X1    g08713(.A1(new_n11589_), .A2(new_n11332_), .A3(new_n11591_), .A4(new_n11592_), .ZN(new_n11593_));
  NOR2_X1    g08714(.A1(new_n11104_), .A2(new_n11575_), .ZN(new_n11594_));
  AOI21_X1   g08715(.A1(new_n11594_), .A2(new_n2622_), .B(new_n2541_), .ZN(new_n11595_));
  AOI21_X1   g08716(.A1(new_n11595_), .A2(new_n10505_), .B(new_n2621_), .ZN(new_n11596_));
  OAI21_X1   g08717(.A1(new_n11593_), .A2(new_n11583_), .B(new_n11596_), .ZN(new_n11597_));
  INV_X1     g08718(.I(new_n11382_), .ZN(new_n11598_));
  NOR2_X1    g08719(.A1(new_n11573_), .A2(new_n5987_), .ZN(new_n11599_));
  OAI21_X1   g08720(.A1(new_n10613_), .A2(new_n11599_), .B(new_n3154_), .ZN(new_n11600_));
  NAND3_X1   g08721(.A1(new_n11598_), .A2(new_n11600_), .A3(new_n11599_), .ZN(new_n11601_));
  NAND2_X1   g08722(.A1(new_n11360_), .A2(new_n2587_), .ZN(new_n11602_));
  NAND2_X1   g08723(.A1(new_n11572_), .A2(new_n2587_), .ZN(new_n11603_));
  OAI21_X1   g08724(.A1(new_n11371_), .A2(new_n11603_), .B(pi0186), .ZN(new_n11604_));
  NAND3_X1   g08725(.A1(new_n11602_), .A2(new_n11572_), .A3(new_n11604_), .ZN(new_n11605_));
  INV_X1     g08726(.I(new_n11373_), .ZN(new_n11606_));
  NAND3_X1   g08727(.A1(new_n11606_), .A2(new_n11572_), .A3(new_n2587_), .ZN(new_n11607_));
  AOI21_X1   g08728(.A1(new_n11607_), .A2(new_n11582_), .B(pi0192), .ZN(new_n11608_));
  OAI21_X1   g08729(.A1(new_n11365_), .A2(pi0299), .B(new_n11608_), .ZN(new_n11609_));
  NOR2_X1    g08730(.A1(new_n11594_), .A2(new_n10800_), .ZN(new_n11610_));
  NOR2_X1    g08731(.A1(new_n11563_), .A2(new_n10526_), .ZN(new_n11611_));
  NOR3_X1    g08732(.A1(new_n11611_), .A2(pi0051), .A3(new_n5356_), .ZN(new_n11613_));
  NOR3_X1    g08733(.A1(new_n11560_), .A2(pi0232), .A3(new_n2621_), .ZN(new_n11614_));
  OAI21_X1   g08734(.A1(new_n2587_), .A2(new_n11613_), .B(new_n11614_), .ZN(new_n11615_));
  OR4_X2     g08735(.A1(new_n11379_), .A2(new_n11615_), .A3(new_n11595_), .A4(new_n11610_), .Z(new_n11616_));
  AOI21_X1   g08736(.A1(new_n11605_), .A2(new_n11609_), .B(new_n11616_), .ZN(new_n11617_));
  NAND2_X1   g08737(.A1(new_n11575_), .A2(new_n10796_), .ZN(new_n11618_));
  NOR2_X1    g08738(.A1(new_n11560_), .A2(po1038), .ZN(new_n11619_));
  NAND2_X1   g08739(.A1(new_n11619_), .A2(new_n11618_), .ZN(new_n11620_));
  AOI21_X1   g08740(.A1(new_n11601_), .A2(new_n11617_), .B(new_n11620_), .ZN(new_n11621_));
  AOI22_X1   g08741(.A1(new_n11621_), .A2(new_n11597_), .B1(new_n11560_), .B2(new_n11565_), .ZN(po0291));
  NOR3_X1    g08742(.A1(new_n11558_), .A2(new_n11556_), .A3(pi0135), .ZN(new_n11623_));
  AOI21_X1   g08743(.A1(pi0135), .A2(new_n11558_), .B(new_n11623_), .ZN(new_n11624_));
  NOR2_X1    g08744(.A1(new_n11624_), .A2(new_n10492_), .ZN(new_n11625_));
  AOI21_X1   g08745(.A1(new_n5988_), .A2(pi0170), .B(new_n10526_), .ZN(new_n11626_));
  NOR3_X1    g08746(.A1(new_n11625_), .A2(new_n11561_), .A3(new_n11626_), .ZN(new_n11627_));
  INV_X1     g08747(.I(pi0194), .ZN(new_n11628_));
  NOR2_X1    g08748(.A1(new_n5109_), .A2(new_n3984_), .ZN(new_n11629_));
  INV_X1     g08749(.I(new_n11629_), .ZN(new_n11630_));
  NOR2_X1    g08750(.A1(new_n11630_), .A2(new_n8167_), .ZN(new_n11631_));
  NAND2_X1   g08751(.A1(new_n11631_), .A2(new_n10577_), .ZN(new_n11632_));
  INV_X1     g08752(.I(new_n11632_), .ZN(new_n11633_));
  OAI21_X1   g08753(.A1(new_n11633_), .A2(new_n11104_), .B(pi0038), .ZN(new_n11634_));
  INV_X1     g08754(.I(new_n11384_), .ZN(new_n11635_));
  OAI21_X1   g08755(.A1(new_n10614_), .A2(pi0170), .B(new_n8166_), .ZN(new_n11636_));
  NAND4_X1   g08756(.A1(new_n11635_), .A2(pi0170), .A3(new_n11382_), .A4(new_n11636_), .ZN(new_n11637_));
  INV_X1     g08757(.I(new_n11637_), .ZN(new_n11638_));
  OAI21_X1   g08758(.A1(pi0299), .A2(new_n10613_), .B(new_n11638_), .ZN(new_n11639_));
  OAI21_X1   g08759(.A1(pi0185), .A2(new_n11373_), .B(new_n11371_), .ZN(new_n11640_));
  NOR4_X1    g08760(.A1(new_n10633_), .A2(new_n3984_), .A3(new_n5109_), .A4(new_n6452_), .ZN(new_n11641_));
  AOI21_X1   g08761(.A1(new_n11629_), .A2(new_n10492_), .B(pi0051), .ZN(new_n11642_));
  INV_X1     g08762(.I(new_n11642_), .ZN(new_n11643_));
  NOR2_X1    g08763(.A1(new_n11643_), .A2(new_n6452_), .ZN(new_n11644_));
  NOR4_X1    g08764(.A1(new_n11641_), .A2(pi0150), .A3(new_n2587_), .A4(new_n11644_), .ZN(new_n11645_));
  NOR2_X1    g08765(.A1(new_n10868_), .A2(pi0051), .ZN(new_n11646_));
  NOR2_X1    g08766(.A1(new_n11646_), .A2(pi0170), .ZN(new_n11647_));
  OAI21_X1   g08767(.A1(new_n11355_), .A2(new_n3984_), .B(new_n2562_), .ZN(new_n11648_));
  OAI22_X1   g08768(.A1(new_n11648_), .A2(new_n11647_), .B1(new_n7170_), .B2(new_n11641_), .ZN(new_n11649_));
  NAND2_X1   g08769(.A1(pi0150), .A2(pi0299), .ZN(new_n11650_));
  AOI21_X1   g08770(.A1(new_n11642_), .A2(new_n5357_), .B(new_n11650_), .ZN(new_n11651_));
  AOI21_X1   g08771(.A1(new_n11649_), .A2(new_n11651_), .B(new_n11645_), .ZN(new_n11652_));
  OR3_X2     g08772(.A1(new_n11652_), .A2(new_n11465_), .A3(new_n11379_), .Z(new_n11653_));
  NOR3_X1    g08773(.A1(new_n11371_), .A2(pi0185), .A3(new_n11606_), .ZN(new_n11654_));
  NOR2_X1    g08774(.A1(new_n11653_), .A2(new_n11654_), .ZN(new_n11655_));
  AOI21_X1   g08775(.A1(new_n11655_), .A2(new_n11640_), .B(pi0038), .ZN(new_n11656_));
  AOI22_X1   g08776(.A1(new_n11639_), .A2(new_n11656_), .B1(new_n11628_), .B2(new_n11634_), .ZN(new_n11657_));
  OAI21_X1   g08777(.A1(pi0185), .A2(new_n11365_), .B(new_n11359_), .ZN(new_n11658_));
  NOR3_X1    g08778(.A1(new_n11359_), .A2(pi0185), .A3(new_n11364_), .ZN(new_n11659_));
  NOR2_X1    g08779(.A1(new_n11653_), .A2(new_n11659_), .ZN(new_n11660_));
  NOR3_X1    g08780(.A1(new_n11382_), .A2(new_n5987_), .A3(pi0299), .ZN(new_n11661_));
  AOI22_X1   g08781(.A1(new_n11637_), .A2(new_n11661_), .B1(new_n11658_), .B2(new_n11660_), .ZN(new_n11662_));
  NAND3_X1   g08782(.A1(new_n5989_), .A2(new_n3984_), .A3(pi0299), .ZN(new_n11663_));
  NOR2_X1    g08783(.A1(new_n11663_), .A2(new_n10575_), .ZN(new_n11664_));
  NOR2_X1    g08784(.A1(new_n11104_), .A2(new_n11664_), .ZN(new_n11665_));
  NAND2_X1   g08785(.A1(new_n11628_), .A2(pi0038), .ZN(new_n11666_));
  OAI21_X1   g08786(.A1(new_n11665_), .A2(new_n11666_), .B(new_n3172_), .ZN(new_n11667_));
  OAI21_X1   g08787(.A1(new_n11662_), .A2(new_n11667_), .B(new_n3173_), .ZN(new_n11668_));
  NOR4_X1    g08788(.A1(new_n11633_), .A2(new_n11628_), .A3(pi0299), .A4(new_n5989_), .ZN(new_n11669_));
  NOR2_X1    g08789(.A1(new_n11669_), .A2(new_n11104_), .ZN(new_n11670_));
  NAND2_X1   g08790(.A1(new_n2541_), .A2(new_n3173_), .ZN(new_n11671_));
  NOR4_X1    g08791(.A1(new_n11624_), .A2(new_n11670_), .A3(new_n10796_), .A4(new_n11671_), .ZN(new_n11672_));
  OAI21_X1   g08792(.A1(new_n11657_), .A2(new_n11668_), .B(new_n11672_), .ZN(new_n11673_));
  NOR2_X1    g08793(.A1(new_n11332_), .A2(new_n8533_), .ZN(new_n11674_));
  NAND2_X1   g08794(.A1(new_n11664_), .A2(new_n8533_), .ZN(new_n11675_));
  AOI21_X1   g08795(.A1(new_n11633_), .A2(new_n8533_), .B(pi0194), .ZN(new_n11676_));
  AOI21_X1   g08796(.A1(pi0194), .A2(new_n11675_), .B(new_n11676_), .ZN(new_n11677_));
  MUX2_X1    g08797(.I0(new_n11324_), .I1(new_n11323_), .S(new_n3984_), .Z(new_n11678_));
  OAI21_X1   g08798(.A1(new_n11678_), .A2(new_n7634_), .B(pi0150), .ZN(new_n11679_));
  NAND2_X1   g08799(.A1(new_n10674_), .A2(new_n11630_), .ZN(new_n11680_));
  NAND3_X1   g08800(.A1(new_n2491_), .A2(pi0170), .A3(new_n5108_), .ZN(new_n11681_));
  NAND3_X1   g08801(.A1(new_n11680_), .A2(new_n7170_), .A3(new_n11681_), .ZN(new_n11682_));
  AOI21_X1   g08802(.A1(new_n11682_), .A2(new_n10038_), .B(pi0299), .ZN(new_n11683_));
  NAND2_X1   g08803(.A1(new_n11675_), .A2(pi0194), .ZN(new_n11684_));
  NOR2_X1    g08804(.A1(new_n10649_), .A2(new_n10066_), .ZN(new_n11685_));
  OAI21_X1   g08805(.A1(new_n10989_), .A2(new_n10066_), .B(new_n11333_), .ZN(new_n11686_));
  AOI22_X1   g08806(.A1(new_n11686_), .A2(new_n11676_), .B1(new_n11684_), .B2(new_n11685_), .ZN(new_n11687_));
  NOR3_X1    g08807(.A1(new_n10577_), .A2(new_n7170_), .A3(new_n11629_), .ZN(new_n11688_));
  NOR2_X1    g08808(.A1(new_n11677_), .A2(new_n11688_), .ZN(new_n11689_));
  OAI21_X1   g08809(.A1(new_n11687_), .A2(pi0299), .B(new_n11689_), .ZN(new_n11690_));
  AOI21_X1   g08810(.A1(new_n11679_), .A2(new_n11683_), .B(new_n11690_), .ZN(new_n11691_));
  OAI22_X1   g08811(.A1(new_n11691_), .A2(new_n5987_), .B1(new_n11674_), .B2(new_n11677_), .ZN(new_n11692_));
  MUX2_X1    g08812(.I0(new_n11692_), .I1(new_n10504_), .S(pi0100), .Z(new_n11693_));
  OR3_X2     g08813(.A1(new_n11693_), .A2(new_n11670_), .A3(new_n11671_), .Z(new_n11694_));
  NAND2_X1   g08814(.A1(new_n11669_), .A2(new_n10796_), .ZN(new_n11695_));
  NOR2_X1    g08815(.A1(new_n11624_), .A2(new_n11695_), .ZN(new_n11696_));
  AOI21_X1   g08816(.A1(new_n11694_), .A2(new_n11696_), .B(po1038), .ZN(new_n11697_));
  AOI21_X1   g08817(.A1(new_n11673_), .A2(new_n11697_), .B(new_n11627_), .ZN(po0292));
  OAI21_X1   g08818(.A1(new_n5989_), .A2(new_n4130_), .B(new_n10492_), .ZN(new_n11699_));
  NOR3_X1    g08819(.A1(new_n11315_), .A2(pi0130), .A3(pi0132), .ZN(new_n11700_));
  NOR2_X1    g08820(.A1(pi0134), .A2(pi0135), .ZN(new_n11701_));
  NOR3_X1    g08821(.A1(new_n11700_), .A2(pi0136), .A3(new_n11701_), .ZN(new_n11702_));
  NAND2_X1   g08822(.A1(new_n11702_), .A2(new_n10577_), .ZN(new_n11703_));
  NAND2_X1   g08823(.A1(new_n11703_), .A2(new_n11699_), .ZN(new_n11704_));
  MUX2_X1    g08824(.I0(new_n10613_), .I1(new_n11382_), .S(new_n7658_), .Z(new_n11705_));
  INV_X1     g08825(.I(pi0141), .ZN(new_n11716_));
  NOR2_X1    g08826(.A1(new_n11716_), .A2(pi0299), .ZN(new_n11717_));
  INV_X1     g08827(.I(new_n11717_), .ZN(new_n11718_));
  NAND2_X1   g08828(.A1(new_n2622_), .A2(pi0232), .ZN(new_n11721_));
  NOR3_X1    g08829(.A1(new_n11705_), .A2(new_n11384_), .A3(new_n11721_), .ZN(new_n11722_));
  AOI21_X1   g08830(.A1(new_n7660_), .A2(new_n10492_), .B(pi0051), .ZN(new_n11723_));
  OAI21_X1   g08831(.A1(new_n11723_), .A2(new_n2621_), .B(new_n2540_), .ZN(new_n11724_));
  INV_X1     g08832(.I(new_n11723_), .ZN(new_n11725_));
  NOR3_X1    g08833(.A1(new_n11725_), .A2(new_n11702_), .A3(new_n10800_), .ZN(new_n11726_));
  OAI21_X1   g08834(.A1(new_n11722_), .A2(new_n11724_), .B(new_n11726_), .ZN(new_n11727_));
  NAND2_X1   g08835(.A1(new_n8534_), .A2(new_n10492_), .ZN(new_n11728_));
  NOR3_X1    g08836(.A1(new_n10577_), .A2(new_n5108_), .A3(new_n7170_), .ZN(new_n11729_));
  OAI21_X1   g08837(.A1(new_n11729_), .A2(new_n4130_), .B(new_n7634_), .ZN(new_n11730_));
  AOI21_X1   g08838(.A1(new_n10643_), .A2(new_n2658_), .B(new_n11730_), .ZN(new_n11731_));
  NAND2_X1   g08839(.A1(new_n11019_), .A2(new_n2658_), .ZN(new_n11732_));
  AOI22_X1   g08840(.A1(new_n11732_), .A2(new_n4130_), .B1(new_n8018_), .B2(new_n10041_), .ZN(new_n11733_));
  NOR2_X1    g08841(.A1(new_n10577_), .A2(pi0148), .ZN(new_n11734_));
  OAI21_X1   g08842(.A1(new_n11733_), .A2(new_n11734_), .B(new_n2587_), .ZN(new_n11735_));
  NOR2_X1    g08843(.A1(new_n11735_), .A2(new_n11731_), .ZN(new_n11736_));
  OR3_X2     g08844(.A1(new_n11333_), .A2(new_n8883_), .A3(new_n7657_), .Z(new_n11737_));
  NAND2_X1   g08845(.A1(new_n11718_), .A2(pi0184), .ZN(new_n11738_));
  OAI22_X1   g08846(.A1(new_n11737_), .A2(new_n10989_), .B1(new_n10649_), .B2(new_n11738_), .ZN(new_n11739_));
  NOR2_X1    g08847(.A1(pi0100), .A2(pi0232), .ZN(new_n11740_));
  OAI21_X1   g08848(.A1(new_n11736_), .A2(new_n11739_), .B(new_n11740_), .ZN(new_n11741_));
  OAI22_X1   g08849(.A1(new_n11674_), .A2(new_n11741_), .B1(new_n11723_), .B2(new_n11728_), .ZN(new_n11742_));
  NOR3_X1    g08850(.A1(new_n11725_), .A2(new_n10526_), .A3(new_n10800_), .ZN(new_n11743_));
  NOR3_X1    g08851(.A1(new_n11743_), .A2(new_n2541_), .A3(new_n11702_), .ZN(new_n11744_));
  AOI21_X1   g08852(.A1(new_n11742_), .A2(new_n11744_), .B(po1038), .ZN(new_n11745_));
  AOI22_X1   g08853(.A1(new_n11727_), .A2(new_n11745_), .B1(new_n11561_), .B2(new_n11704_), .ZN(po0293));
  NOR3_X1    g08854(.A1(new_n8163_), .A2(pi0210), .A3(new_n2575_), .ZN(new_n11747_));
  NAND2_X1   g08855(.A1(po1038), .A2(new_n11747_), .ZN(new_n11748_));
  NOR2_X1    g08856(.A1(po1038), .A2(pi0299), .ZN(new_n11749_));
  NOR2_X1    g08857(.A1(new_n8755_), .A2(pi0198), .ZN(new_n11750_));
  AOI22_X1   g08858(.A1(new_n11749_), .A2(new_n11750_), .B1(pi0299), .B2(new_n11747_), .ZN(new_n11751_));
  OAI21_X1   g08859(.A1(new_n8164_), .A2(new_n10843_), .B(new_n11751_), .ZN(new_n11752_));
  AOI21_X1   g08860(.A1(new_n11752_), .A2(new_n11748_), .B(new_n5987_), .ZN(new_n11753_));
  MUX2_X1    g08861(.I0(new_n11753_), .I1(pi0137), .S(new_n3154_), .Z(po0294));
  INV_X1     g08862(.I(pi0138), .ZN(new_n11755_));
  NOR4_X1    g08863(.A1(new_n7120_), .A2(pi0055), .A3(pi0092), .A4(new_n7147_), .ZN(new_n11756_));
  AOI21_X1   g08864(.A1(new_n7121_), .A2(new_n3177_), .B(pi0075), .ZN(new_n11757_));
  AOI21_X1   g08865(.A1(new_n5109_), .A2(new_n7519_), .B(new_n7511_), .ZN(new_n11758_));
  NAND3_X1   g08866(.A1(new_n7511_), .A2(new_n5109_), .A3(new_n7518_), .ZN(new_n11759_));
  NAND2_X1   g08867(.A1(new_n11759_), .A2(new_n2587_), .ZN(new_n11760_));
  NOR2_X1    g08868(.A1(new_n11760_), .A2(new_n11758_), .ZN(new_n11761_));
  INV_X1     g08869(.I(new_n11761_), .ZN(new_n11762_));
  NAND4_X1   g08870(.A1(new_n7519_), .A2(new_n11716_), .A3(new_n5987_), .A4(new_n2587_), .ZN(new_n11766_));
  NOR2_X1    g08871(.A1(new_n7518_), .A2(pi0299), .ZN(new_n11767_));
  INV_X1     g08872(.I(new_n11767_), .ZN(new_n11768_));
  AOI21_X1   g08873(.A1(new_n7453_), .A2(pi0299), .B(pi0232), .ZN(new_n11769_));
  AOI21_X1   g08874(.A1(new_n11769_), .A2(new_n11768_), .B(pi0039), .ZN(new_n11770_));
  INV_X1     g08875(.I(new_n11770_), .ZN(new_n11771_));
  NAND4_X1   g08876(.A1(new_n11762_), .A2(pi0141), .A3(new_n11766_), .A4(new_n11771_), .ZN(new_n11772_));
  AOI21_X1   g08877(.A1(new_n5094_), .A2(new_n9028_), .B(new_n7630_), .ZN(new_n11773_));
  OAI21_X1   g08878(.A1(new_n11773_), .A2(new_n7634_), .B(new_n7597_), .ZN(new_n11774_));
  NOR2_X1    g08879(.A1(new_n7630_), .A2(new_n9028_), .ZN(new_n11775_));
  NOR4_X1    g08880(.A1(new_n11775_), .A2(new_n7087_), .A3(new_n7154_), .A4(new_n7610_), .ZN(new_n11776_));
  NOR2_X1    g08881(.A1(new_n7605_), .A2(pi0299), .ZN(new_n11777_));
  INV_X1     g08882(.I(new_n11777_), .ZN(new_n11778_));
  NOR2_X1    g08883(.A1(new_n11776_), .A2(new_n11778_), .ZN(new_n11779_));
  INV_X1     g08884(.I(new_n11779_), .ZN(new_n11780_));
  AOI21_X1   g08885(.A1(new_n11780_), .A2(new_n11774_), .B(pi0232), .ZN(new_n11781_));
  INV_X1     g08886(.I(new_n11781_), .ZN(new_n11782_));
  NAND2_X1   g08887(.A1(new_n11776_), .A2(new_n7607_), .ZN(new_n11783_));
  NAND2_X1   g08888(.A1(new_n11783_), .A2(new_n11777_), .ZN(new_n11784_));
  INV_X1     g08889(.I(new_n11784_), .ZN(new_n11785_));
  NOR2_X1    g08890(.A1(new_n11785_), .A2(new_n11716_), .ZN(new_n11786_));
  NOR3_X1    g08891(.A1(new_n7606_), .A2(new_n11775_), .A3(new_n5094_), .ZN(new_n11787_));
  NOR2_X1    g08892(.A1(new_n4130_), .A2(pi0299), .ZN(new_n11788_));
  OAI21_X1   g08893(.A1(new_n11787_), .A2(new_n7596_), .B(new_n11788_), .ZN(new_n11789_));
  NAND2_X1   g08894(.A1(new_n11780_), .A2(pi0141), .ZN(new_n11790_));
  NAND3_X1   g08895(.A1(new_n11790_), .A2(pi0232), .A3(new_n11789_), .ZN(new_n11791_));
  OAI21_X1   g08896(.A1(new_n11791_), .A2(new_n11786_), .B(new_n11782_), .ZN(new_n11792_));
  AOI21_X1   g08897(.A1(new_n11792_), .A2(pi0039), .B(new_n2622_), .ZN(new_n11793_));
  AOI21_X1   g08898(.A1(new_n11772_), .A2(new_n11793_), .B(pi0087), .ZN(new_n11794_));
  NOR4_X1    g08899(.A1(new_n7119_), .A2(pi0092), .A3(new_n2538_), .A4(new_n7146_), .ZN(new_n11795_));
  INV_X1     g08900(.I(new_n11795_), .ZN(new_n11796_));
  NOR2_X1    g08901(.A1(new_n11796_), .A2(pi0092), .ZN(new_n11797_));
  OAI21_X1   g08902(.A1(new_n11794_), .A2(new_n11757_), .B(new_n11797_), .ZN(new_n11798_));
  AOI21_X1   g08903(.A1(new_n11798_), .A2(new_n3227_), .B(new_n11756_), .ZN(new_n11799_));
  OAI21_X1   g08904(.A1(new_n11799_), .A2(new_n3503_), .B(new_n7681_), .ZN(new_n11800_));
  NOR2_X1    g08905(.A1(new_n7252_), .A2(new_n2515_), .ZN(new_n11801_));
  INV_X1     g08906(.I(new_n11801_), .ZN(new_n11802_));
  NOR2_X1    g08907(.A1(new_n11802_), .A2(new_n7660_), .ZN(new_n11803_));
  NOR2_X1    g08908(.A1(new_n4130_), .A2(new_n2587_), .ZN(new_n11804_));
  NAND2_X1   g08909(.A1(new_n6548_), .A2(new_n11804_), .ZN(new_n11805_));
  NOR2_X1    g08910(.A1(new_n5370_), .A2(new_n6548_), .ZN(new_n11806_));
  NAND2_X1   g08911(.A1(new_n11806_), .A2(new_n7153_), .ZN(new_n11807_));
  NOR4_X1    g08912(.A1(new_n8690_), .A2(new_n5987_), .A3(new_n11717_), .A4(new_n11805_), .ZN(new_n11809_));
  MUX2_X1    g08913(.I0(new_n11809_), .I1(new_n11803_), .S(new_n3154_), .Z(new_n11810_));
  NAND2_X1   g08914(.A1(new_n11810_), .A2(new_n7855_), .ZN(new_n11811_));
  AOI21_X1   g08915(.A1(new_n11755_), .A2(new_n11811_), .B(new_n11800_), .ZN(new_n11812_));
  INV_X1     g08916(.I(new_n11811_), .ZN(new_n11813_));
  AND3_X2    g08917(.A1(new_n11800_), .A2(new_n11755_), .A3(new_n11813_), .Z(new_n11814_));
  NOR2_X1    g08918(.A1(new_n10213_), .A2(pi0118), .ZN(new_n11815_));
  INV_X1     g08919(.I(new_n11815_), .ZN(new_n11816_));
  NOR2_X1    g08920(.A1(new_n11816_), .A2(pi0139), .ZN(new_n11817_));
  INV_X1     g08921(.I(new_n11817_), .ZN(new_n11818_));
  INV_X1     g08922(.I(pi0195), .ZN(new_n11819_));
  INV_X1     g08923(.I(pi0196), .ZN(new_n11820_));
  AOI21_X1   g08924(.A1(new_n11819_), .A2(new_n11820_), .B(pi0138), .ZN(new_n11821_));
  AND2_X2    g08925(.A1(new_n11800_), .A2(new_n11821_), .Z(new_n11822_));
  NOR2_X1    g08926(.A1(new_n11813_), .A2(new_n11821_), .ZN(new_n11823_));
  OAI21_X1   g08927(.A1(new_n11822_), .A2(new_n11823_), .B(new_n11818_), .ZN(new_n11824_));
  NOR3_X1    g08928(.A1(new_n11824_), .A2(new_n11812_), .A3(new_n11814_), .ZN(po0295));
  INV_X1     g08929(.I(pi0139), .ZN(new_n11826_));
  NOR4_X1    g08930(.A1(new_n7518_), .A2(pi0191), .A3(pi0232), .A4(pi0299), .ZN(new_n11829_));
  NOR3_X1    g08931(.A1(new_n11770_), .A2(new_n11361_), .A3(new_n11829_), .ZN(new_n11830_));
  NOR2_X1    g08932(.A1(new_n11784_), .A2(new_n11361_), .ZN(new_n11831_));
  INV_X1     g08933(.I(new_n7630_), .ZN(new_n11832_));
  NOR2_X1    g08934(.A1(new_n11832_), .A2(pi0169), .ZN(new_n11833_));
  OAI21_X1   g08935(.A1(new_n11787_), .A2(new_n11833_), .B(new_n7170_), .ZN(new_n11834_));
  INV_X1     g08936(.I(new_n11834_), .ZN(new_n11835_));
  NOR2_X1    g08937(.A1(new_n11779_), .A2(pi0191), .ZN(new_n11836_));
  NAND2_X1   g08938(.A1(new_n7597_), .A2(new_n5987_), .ZN(new_n11837_));
  NOR4_X1    g08939(.A1(new_n11831_), .A2(new_n11835_), .A3(new_n11836_), .A4(new_n11837_), .ZN(new_n11838_));
  OAI21_X1   g08940(.A1(new_n11838_), .A2(new_n11781_), .B(new_n3319_), .ZN(new_n11839_));
  AOI21_X1   g08941(.A1(new_n11762_), .A2(new_n11830_), .B(new_n11839_), .ZN(new_n11840_));
  NOR2_X1    g08942(.A1(new_n11840_), .A2(pi0087), .ZN(new_n11841_));
  OAI21_X1   g08943(.A1(new_n11841_), .A2(new_n11757_), .B(new_n3203_), .ZN(new_n11842_));
  NAND2_X1   g08944(.A1(new_n11842_), .A2(new_n11795_), .ZN(new_n11843_));
  NOR2_X1    g08945(.A1(new_n11756_), .A2(pi0055), .ZN(new_n11844_));
  NAND2_X1   g08946(.A1(new_n11843_), .A2(new_n11844_), .ZN(new_n11845_));
  NOR2_X1    g08947(.A1(new_n3503_), .A2(new_n2571_), .ZN(new_n11846_));
  AND2_X2    g08948(.A1(new_n11845_), .A2(new_n11846_), .Z(new_n11847_));
  INV_X1     g08949(.I(new_n11847_), .ZN(new_n11848_));
  NOR2_X1    g08950(.A1(new_n11802_), .A2(new_n11336_), .ZN(new_n11849_));
  INV_X1     g08951(.I(new_n11849_), .ZN(new_n11850_));
  NOR3_X1    g08952(.A1(new_n5143_), .A2(new_n4272_), .A3(new_n2587_), .ZN(new_n11851_));
  NOR2_X1    g08953(.A1(new_n11807_), .A2(new_n11361_), .ZN(new_n11852_));
  INV_X1     g08954(.I(new_n8689_), .ZN(new_n11853_));
  OAI21_X1   g08955(.A1(new_n11853_), .A2(new_n11361_), .B(new_n2587_), .ZN(new_n11854_));
  OAI22_X1   g08956(.A1(new_n11854_), .A2(new_n11852_), .B1(new_n8688_), .B2(new_n11851_), .ZN(new_n11855_));
  MUX2_X1    g08957(.I0(new_n11855_), .I1(new_n8691_), .S(new_n5987_), .Z(new_n11856_));
  MUX2_X1    g08958(.I0(new_n11856_), .I1(new_n11850_), .S(new_n3154_), .Z(new_n11857_));
  NOR2_X1    g08959(.A1(new_n11857_), .A2(new_n7856_), .ZN(new_n11858_));
  INV_X1     g08960(.I(new_n11858_), .ZN(new_n11859_));
  AOI21_X1   g08961(.A1(new_n11826_), .A2(new_n11859_), .B(new_n11848_), .ZN(new_n11860_));
  NOR3_X1    g08962(.A1(new_n11847_), .A2(pi0139), .A3(new_n11859_), .ZN(new_n11861_));
  NOR2_X1    g08963(.A1(pi0138), .A2(pi0195), .ZN(new_n11862_));
  AOI21_X1   g08964(.A1(new_n11862_), .A2(new_n11820_), .B(pi0139), .ZN(new_n11863_));
  OAI21_X1   g08965(.A1(new_n11858_), .A2(new_n11863_), .B(new_n11816_), .ZN(new_n11864_));
  AOI21_X1   g08966(.A1(new_n11848_), .A2(new_n11863_), .B(new_n11864_), .ZN(new_n11865_));
  NOR4_X1    g08967(.A1(new_n11860_), .A2(new_n11815_), .A3(new_n11865_), .A4(new_n11861_), .ZN(po0296));
  INV_X1     g08968(.I(pi0790), .ZN(new_n11867_));
  INV_X1     g08969(.I(pi0792), .ZN(new_n11868_));
  INV_X1     g08970(.I(pi1159), .ZN(new_n11869_));
  INV_X1     g08971(.I(pi0785), .ZN(new_n11870_));
  NOR2_X1    g08972(.A1(new_n2925_), .A2(pi0140), .ZN(new_n11871_));
  INV_X1     g08973(.I(pi0621), .ZN(new_n11872_));
  NOR2_X1    g08974(.A1(new_n11872_), .A2(new_n2918_), .ZN(new_n11873_));
  NOR2_X1    g08975(.A1(new_n11873_), .A2(new_n5101_), .ZN(new_n11874_));
  INV_X1     g08976(.I(new_n11874_), .ZN(new_n11875_));
  NOR2_X1    g08977(.A1(new_n11875_), .A2(new_n2926_), .ZN(new_n11876_));
  INV_X1     g08978(.I(new_n11876_), .ZN(new_n11877_));
  NOR2_X1    g08979(.A1(new_n11877_), .A2(pi0761), .ZN(new_n11878_));
  NOR2_X1    g08980(.A1(new_n11878_), .A2(new_n11871_), .ZN(new_n11879_));
  INV_X1     g08981(.I(new_n11879_), .ZN(new_n11880_));
  INV_X1     g08982(.I(pi0738), .ZN(new_n11881_));
  INV_X1     g08983(.I(pi0665), .ZN(new_n11882_));
  NOR2_X1    g08984(.A1(new_n11882_), .A2(new_n2918_), .ZN(new_n11883_));
  NOR2_X1    g08985(.A1(new_n11883_), .A2(new_n5095_), .ZN(new_n11884_));
  INV_X1     g08986(.I(new_n11884_), .ZN(new_n11885_));
  NOR2_X1    g08987(.A1(new_n11885_), .A2(new_n2926_), .ZN(new_n11886_));
  AOI21_X1   g08988(.A1(new_n11886_), .A2(new_n11881_), .B(new_n11871_), .ZN(new_n11887_));
  NOR2_X1    g08989(.A1(new_n11887_), .A2(new_n11874_), .ZN(new_n11888_));
  NOR2_X1    g08990(.A1(new_n11880_), .A2(new_n11888_), .ZN(new_n11889_));
  NOR2_X1    g08991(.A1(new_n11889_), .A2(pi0778), .ZN(new_n11890_));
  INV_X1     g08992(.I(pi0778), .ZN(new_n11891_));
  NAND2_X1   g08993(.A1(new_n11888_), .A2(pi0625), .ZN(new_n11892_));
  INV_X1     g08994(.I(pi1153), .ZN(new_n11893_));
  INV_X1     g08995(.I(new_n11886_), .ZN(new_n11894_));
  NOR3_X1    g08996(.A1(new_n11894_), .A2(pi0625), .A3(pi0738), .ZN(new_n11895_));
  NOR4_X1    g08997(.A1(new_n11878_), .A2(pi0608), .A3(new_n11893_), .A4(new_n11871_), .ZN(new_n11896_));
  OAI21_X1   g08998(.A1(new_n11880_), .A2(new_n11888_), .B(new_n11892_), .ZN(new_n11897_));
  NOR3_X1    g08999(.A1(new_n11871_), .A2(pi0608), .A3(pi1153), .ZN(new_n11898_));
  AOI22_X1   g09000(.A1(new_n11897_), .A2(new_n11898_), .B1(new_n11892_), .B2(new_n11896_), .ZN(new_n11899_));
  NOR2_X1    g09001(.A1(new_n11899_), .A2(new_n11891_), .ZN(new_n11900_));
  XOR2_X1    g09002(.A1(new_n11900_), .A2(new_n11890_), .Z(new_n11901_));
  INV_X1     g09003(.I(new_n11901_), .ZN(new_n11902_));
  INV_X1     g09004(.I(pi0609), .ZN(new_n11903_));
  AOI21_X1   g09005(.A1(new_n11901_), .A2(new_n11903_), .B(pi1155), .ZN(new_n11904_));
  INV_X1     g09006(.I(new_n11887_), .ZN(new_n11905_));
  XOR2_X1    g09007(.A1(new_n11895_), .A2(pi1153), .Z(new_n11906_));
  NAND2_X1   g09008(.A1(new_n11906_), .A2(new_n11905_), .ZN(new_n11907_));
  OAI21_X1   g09009(.A1(new_n11895_), .A2(new_n11871_), .B(new_n11893_), .ZN(new_n11908_));
  AOI21_X1   g09010(.A1(new_n11907_), .A2(new_n11908_), .B(new_n11891_), .ZN(new_n11909_));
  NOR2_X1    g09011(.A1(new_n11887_), .A2(pi0778), .ZN(new_n11910_));
  OAI21_X1   g09012(.A1(new_n11909_), .A2(new_n11910_), .B(pi0609), .ZN(new_n11911_));
  INV_X1     g09013(.I(pi1155), .ZN(new_n11912_));
  XNOR2_X1   g09014(.A1(pi0608), .A2(pi1153), .ZN(new_n11913_));
  NOR2_X1    g09015(.A1(new_n11913_), .A2(new_n11891_), .ZN(new_n11914_));
  NOR2_X1    g09016(.A1(new_n11914_), .A2(new_n11903_), .ZN(new_n11915_));
  NOR2_X1    g09017(.A1(new_n11915_), .A2(new_n2926_), .ZN(new_n11916_));
  INV_X1     g09018(.I(new_n11916_), .ZN(new_n11917_));
  AOI21_X1   g09019(.A1(new_n11880_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n11918_));
  NOR2_X1    g09020(.A1(new_n11918_), .A2(pi0660), .ZN(new_n11919_));
  OAI21_X1   g09021(.A1(new_n11904_), .A2(new_n11911_), .B(new_n11919_), .ZN(new_n11920_));
  NOR2_X1    g09022(.A1(new_n11909_), .A2(new_n11910_), .ZN(new_n11921_));
  NAND4_X1   g09023(.A1(new_n11902_), .A2(pi0609), .A3(new_n11912_), .A4(new_n11921_), .ZN(new_n11922_));
  INV_X1     g09024(.I(pi0660), .ZN(new_n11923_));
  INV_X1     g09025(.I(new_n11914_), .ZN(new_n11924_));
  NOR2_X1    g09026(.A1(new_n11924_), .A2(new_n2926_), .ZN(new_n11925_));
  NOR2_X1    g09027(.A1(new_n11879_), .A2(new_n11925_), .ZN(new_n11926_));
  NOR2_X1    g09028(.A1(new_n2926_), .A2(new_n11903_), .ZN(new_n11927_));
  INV_X1     g09029(.I(new_n11927_), .ZN(new_n11928_));
  AOI21_X1   g09030(.A1(new_n11926_), .A2(new_n11928_), .B(pi1155), .ZN(new_n11929_));
  NOR2_X1    g09031(.A1(new_n11929_), .A2(new_n11923_), .ZN(new_n11930_));
  AOI21_X1   g09032(.A1(new_n11922_), .A2(new_n11930_), .B(new_n11870_), .ZN(new_n11931_));
  AOI22_X1   g09033(.A1(new_n11931_), .A2(new_n11920_), .B1(new_n11870_), .B2(new_n11902_), .ZN(new_n11932_));
  OR2_X2     g09034(.A1(new_n11932_), .A2(pi0781), .Z(new_n11933_));
  INV_X1     g09035(.I(pi0618), .ZN(new_n11934_));
  AOI21_X1   g09036(.A1(new_n11932_), .A2(new_n11934_), .B(pi1154), .ZN(new_n11935_));
  NOR2_X1    g09037(.A1(new_n11912_), .A2(pi0660), .ZN(new_n11936_));
  NOR2_X1    g09038(.A1(new_n11923_), .A2(pi1155), .ZN(new_n11937_));
  OAI21_X1   g09039(.A1(new_n11936_), .A2(new_n11937_), .B(pi0785), .ZN(new_n11938_));
  NOR2_X1    g09040(.A1(new_n11938_), .A2(new_n2926_), .ZN(new_n11939_));
  NOR2_X1    g09041(.A1(new_n11921_), .A2(new_n11939_), .ZN(new_n11940_));
  NAND2_X1   g09042(.A1(new_n11940_), .A2(pi0618), .ZN(new_n11941_));
  NOR2_X1    g09043(.A1(new_n11929_), .A2(new_n11918_), .ZN(new_n11942_));
  MUX2_X1    g09044(.I0(new_n11942_), .I1(new_n11926_), .S(new_n11870_), .Z(new_n11943_));
  NOR3_X1    g09045(.A1(new_n2926_), .A2(pi0618), .A3(pi1154), .ZN(new_n11944_));
  INV_X1     g09046(.I(new_n11944_), .ZN(new_n11945_));
  NOR2_X1    g09047(.A1(new_n11943_), .A2(new_n11945_), .ZN(new_n11946_));
  NOR2_X1    g09048(.A1(new_n11946_), .A2(pi0627), .ZN(new_n11947_));
  OAI21_X1   g09049(.A1(new_n11935_), .A2(new_n11941_), .B(new_n11947_), .ZN(new_n11948_));
  INV_X1     g09050(.I(pi0627), .ZN(new_n11949_));
  INV_X1     g09051(.I(pi1154), .ZN(new_n11950_));
  NOR2_X1    g09052(.A1(new_n2926_), .A2(new_n11934_), .ZN(new_n11951_));
  INV_X1     g09053(.I(new_n11951_), .ZN(new_n11952_));
  OAI21_X1   g09054(.A1(new_n11943_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n11953_));
  NOR4_X1    g09055(.A1(new_n11932_), .A2(new_n11934_), .A3(pi1154), .A4(new_n11940_), .ZN(new_n11954_));
  OAI21_X1   g09056(.A1(new_n11954_), .A2(new_n11953_), .B(new_n11949_), .ZN(new_n11955_));
  NAND2_X1   g09057(.A1(new_n11955_), .A2(new_n11948_), .ZN(new_n11956_));
  NAND2_X1   g09058(.A1(new_n11956_), .A2(pi0781), .ZN(new_n11957_));
  NAND2_X1   g09059(.A1(new_n11957_), .A2(new_n11933_), .ZN(new_n11958_));
  NOR2_X1    g09060(.A1(new_n11950_), .A2(pi0627), .ZN(new_n11959_));
  NOR2_X1    g09061(.A1(new_n11949_), .A2(pi1154), .ZN(new_n11960_));
  OAI21_X1   g09062(.A1(new_n11959_), .A2(new_n11960_), .B(pi0781), .ZN(new_n11961_));
  NOR2_X1    g09063(.A1(new_n11961_), .A2(new_n2926_), .ZN(new_n11962_));
  INV_X1     g09064(.I(new_n11962_), .ZN(new_n11963_));
  NAND2_X1   g09065(.A1(new_n11940_), .A2(new_n11963_), .ZN(new_n11964_));
  NAND4_X1   g09066(.A1(new_n11958_), .A2(pi0619), .A3(new_n11869_), .A4(new_n11964_), .ZN(new_n11965_));
  INV_X1     g09067(.I(pi0648), .ZN(new_n11966_));
  INV_X1     g09068(.I(pi0619), .ZN(new_n11967_));
  NOR2_X1    g09069(.A1(new_n11943_), .A2(pi0781), .ZN(new_n11968_));
  INV_X1     g09070(.I(pi0781), .ZN(new_n11969_));
  NOR2_X1    g09071(.A1(new_n11953_), .A2(new_n11946_), .ZN(new_n11970_));
  NOR2_X1    g09072(.A1(new_n11970_), .A2(new_n11969_), .ZN(new_n11971_));
  XOR2_X1    g09073(.A1(new_n11971_), .A2(new_n11968_), .Z(new_n11972_));
  INV_X1     g09074(.I(new_n11972_), .ZN(new_n11973_));
  NOR2_X1    g09075(.A1(new_n11973_), .A2(new_n11967_), .ZN(new_n11974_));
  INV_X1     g09076(.I(new_n11871_), .ZN(new_n11975_));
  OAI21_X1   g09077(.A1(new_n11975_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n11976_));
  NOR3_X1    g09078(.A1(new_n11974_), .A2(new_n11966_), .A3(new_n11976_), .ZN(new_n11977_));
  INV_X1     g09079(.I(new_n11964_), .ZN(new_n11978_));
  OAI21_X1   g09080(.A1(new_n11958_), .A2(pi0619), .B(new_n11869_), .ZN(new_n11979_));
  NAND3_X1   g09081(.A1(new_n11979_), .A2(pi0619), .A3(new_n11978_), .ZN(new_n11980_));
  INV_X1     g09082(.I(new_n11974_), .ZN(new_n11981_));
  AOI21_X1   g09083(.A1(new_n11975_), .A2(new_n11967_), .B(pi1159), .ZN(new_n11982_));
  AOI21_X1   g09084(.A1(new_n11981_), .A2(new_n11982_), .B(pi0648), .ZN(new_n11983_));
  AOI22_X1   g09085(.A1(new_n11980_), .A2(new_n11983_), .B1(new_n11965_), .B2(new_n11977_), .ZN(new_n11984_));
  INV_X1     g09086(.I(pi0789), .ZN(new_n11985_));
  INV_X1     g09087(.I(pi0788), .ZN(new_n11986_));
  INV_X1     g09088(.I(pi1158), .ZN(new_n11987_));
  NOR2_X1    g09089(.A1(new_n11987_), .A2(pi0641), .ZN(new_n11988_));
  INV_X1     g09090(.I(pi0641), .ZN(new_n11989_));
  NOR2_X1    g09091(.A1(new_n11989_), .A2(pi1158), .ZN(new_n11990_));
  NOR2_X1    g09092(.A1(new_n11988_), .A2(new_n11990_), .ZN(new_n11991_));
  NOR2_X1    g09093(.A1(new_n11991_), .A2(new_n11986_), .ZN(new_n11992_));
  NOR2_X1    g09094(.A1(new_n11987_), .A2(pi0626), .ZN(new_n11993_));
  INV_X1     g09095(.I(pi0626), .ZN(new_n11994_));
  NOR2_X1    g09096(.A1(new_n11994_), .A2(pi1158), .ZN(new_n11995_));
  NOR2_X1    g09097(.A1(new_n11993_), .A2(new_n11995_), .ZN(new_n11996_));
  NOR2_X1    g09098(.A1(new_n11996_), .A2(new_n11986_), .ZN(new_n11997_));
  NOR2_X1    g09099(.A1(new_n11992_), .A2(new_n11997_), .ZN(new_n11998_));
  INV_X1     g09100(.I(new_n11998_), .ZN(new_n11999_));
  OAI21_X1   g09101(.A1(new_n11958_), .A2(new_n11999_), .B(new_n11985_), .ZN(new_n12000_));
  NOR2_X1    g09102(.A1(new_n11984_), .A2(new_n12000_), .ZN(new_n12001_));
  INV_X1     g09103(.I(new_n11991_), .ZN(new_n12002_));
  INV_X1     g09104(.I(new_n11996_), .ZN(new_n12003_));
  NOR2_X1    g09105(.A1(new_n11973_), .A2(pi0789), .ZN(new_n12004_));
  NAND3_X1   g09106(.A1(new_n11975_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n12005_));
  NAND2_X1   g09107(.A1(new_n12005_), .A2(pi0789), .ZN(new_n12006_));
  XNOR2_X1   g09108(.A1(new_n12004_), .A2(new_n12006_), .ZN(new_n12007_));
  INV_X1     g09109(.I(new_n12007_), .ZN(new_n12008_));
  MUX2_X1    g09110(.I0(new_n12008_), .I1(new_n11871_), .S(new_n12003_), .Z(new_n12009_));
  NOR2_X1    g09111(.A1(new_n11869_), .A2(pi0648), .ZN(new_n12010_));
  NOR2_X1    g09112(.A1(new_n11966_), .A2(pi1159), .ZN(new_n12011_));
  NOR2_X1    g09113(.A1(new_n12010_), .A2(new_n12011_), .ZN(new_n12012_));
  NOR2_X1    g09114(.A1(new_n12012_), .A2(new_n11985_), .ZN(new_n12013_));
  INV_X1     g09115(.I(new_n12013_), .ZN(new_n12014_));
  NOR2_X1    g09116(.A1(new_n12014_), .A2(new_n2926_), .ZN(new_n12015_));
  NOR2_X1    g09117(.A1(new_n11989_), .A2(new_n11987_), .ZN(new_n12016_));
  NOR2_X1    g09118(.A1(pi0641), .A2(pi1158), .ZN(new_n12017_));
  INV_X1     g09119(.I(new_n12017_), .ZN(new_n12018_));
  NOR2_X1    g09120(.A1(new_n12018_), .A2(new_n11994_), .ZN(new_n12019_));
  AOI21_X1   g09121(.A1(new_n11994_), .A2(new_n12016_), .B(new_n12019_), .ZN(new_n12020_));
  NOR2_X1    g09122(.A1(new_n12015_), .A2(new_n12020_), .ZN(new_n12021_));
  INV_X1     g09123(.I(new_n12021_), .ZN(new_n12022_));
  OAI21_X1   g09124(.A1(new_n11964_), .A2(new_n12022_), .B(pi0788), .ZN(new_n12023_));
  AOI21_X1   g09125(.A1(new_n12009_), .A2(new_n12002_), .B(new_n12023_), .ZN(new_n12024_));
  NOR2_X1    g09126(.A1(new_n12001_), .A2(new_n12024_), .ZN(new_n12025_));
  INV_X1     g09127(.I(pi1156), .ZN(new_n12026_));
  NOR2_X1    g09128(.A1(new_n12007_), .A2(pi0788), .ZN(new_n12027_));
  AOI21_X1   g09129(.A1(new_n12009_), .A2(pi0788), .B(new_n12027_), .ZN(new_n12028_));
  NAND4_X1   g09130(.A1(new_n12025_), .A2(pi0628), .A3(new_n12026_), .A4(new_n12028_), .ZN(new_n12029_));
  INV_X1     g09131(.I(pi0629), .ZN(new_n12030_));
  INV_X1     g09132(.I(pi0628), .ZN(new_n12031_));
  NOR2_X1    g09133(.A1(new_n11992_), .A2(new_n12013_), .ZN(new_n12032_));
  NOR2_X1    g09134(.A1(new_n12032_), .A2(new_n2926_), .ZN(new_n12033_));
  INV_X1     g09135(.I(new_n12033_), .ZN(new_n12034_));
  NOR2_X1    g09136(.A1(new_n11978_), .A2(new_n12034_), .ZN(new_n12035_));
  OAI21_X1   g09137(.A1(new_n12031_), .A2(new_n2926_), .B(new_n12035_), .ZN(new_n12036_));
  AOI21_X1   g09138(.A1(new_n12036_), .A2(new_n12026_), .B(new_n12030_), .ZN(new_n12037_));
  NAND2_X1   g09139(.A1(new_n12029_), .A2(new_n12037_), .ZN(new_n12038_));
  NOR2_X1    g09140(.A1(new_n12025_), .A2(pi0628), .ZN(new_n12039_));
  NOR2_X1    g09141(.A1(new_n12039_), .A2(pi1156), .ZN(new_n12040_));
  OR2_X2     g09142(.A1(new_n12028_), .A2(new_n12031_), .Z(new_n12041_));
  AOI21_X1   g09143(.A1(new_n2925_), .A2(new_n12031_), .B(pi1156), .ZN(new_n12042_));
  AND2_X2    g09144(.A1(new_n12035_), .A2(new_n12042_), .Z(new_n12043_));
  OAI22_X1   g09145(.A1(new_n12040_), .A2(new_n12041_), .B1(pi0629), .B2(new_n12043_), .ZN(new_n12044_));
  AOI21_X1   g09146(.A1(new_n12044_), .A2(new_n12038_), .B(new_n11868_), .ZN(new_n12045_));
  AOI21_X1   g09147(.A1(new_n11868_), .A2(new_n12025_), .B(new_n12045_), .ZN(new_n12046_));
  NOR2_X1    g09148(.A1(new_n12046_), .A2(pi0787), .ZN(new_n12047_));
  INV_X1     g09149(.I(pi0787), .ZN(new_n12048_));
  INV_X1     g09150(.I(pi1157), .ZN(new_n12049_));
  NOR2_X1    g09151(.A1(new_n12026_), .A2(pi0629), .ZN(new_n12050_));
  NOR2_X1    g09152(.A1(new_n12030_), .A2(pi1156), .ZN(new_n12051_));
  NOR2_X1    g09153(.A1(new_n12050_), .A2(new_n12051_), .ZN(new_n12052_));
  NOR2_X1    g09154(.A1(new_n12052_), .A2(new_n11868_), .ZN(new_n12053_));
  INV_X1     g09155(.I(new_n12053_), .ZN(new_n12054_));
  NOR2_X1    g09156(.A1(new_n12054_), .A2(new_n11871_), .ZN(new_n12055_));
  AOI21_X1   g09157(.A1(new_n12028_), .A2(new_n12054_), .B(new_n12055_), .ZN(new_n12056_));
  XOR2_X1    g09158(.A1(new_n12046_), .A2(new_n12056_), .Z(new_n12057_));
  NAND2_X1   g09159(.A1(new_n12057_), .A2(pi0647), .ZN(new_n12058_));
  XOR2_X1    g09160(.A1(new_n12058_), .A2(new_n12046_), .Z(new_n12059_));
  INV_X1     g09161(.I(pi0630), .ZN(new_n12060_));
  INV_X1     g09162(.I(pi0647), .ZN(new_n12061_));
  INV_X1     g09163(.I(new_n12035_), .ZN(new_n12062_));
  NOR2_X1    g09164(.A1(new_n12031_), .A2(pi1156), .ZN(new_n12063_));
  NOR2_X1    g09165(.A1(new_n12026_), .A2(pi0628), .ZN(new_n12064_));
  NOR2_X1    g09166(.A1(new_n12063_), .A2(new_n12064_), .ZN(new_n12065_));
  NOR2_X1    g09167(.A1(new_n12065_), .A2(new_n11868_), .ZN(new_n12066_));
  INV_X1     g09168(.I(new_n12066_), .ZN(new_n12067_));
  NOR2_X1    g09169(.A1(new_n12067_), .A2(new_n2926_), .ZN(new_n12068_));
  NOR2_X1    g09170(.A1(new_n12062_), .A2(new_n12068_), .ZN(new_n12069_));
  NOR2_X1    g09171(.A1(new_n12069_), .A2(new_n12061_), .ZN(new_n12070_));
  OAI21_X1   g09172(.A1(new_n11871_), .A2(pi0647), .B(new_n12049_), .ZN(new_n12071_));
  OAI21_X1   g09173(.A1(new_n12070_), .A2(new_n12071_), .B(new_n12060_), .ZN(new_n12072_));
  AOI21_X1   g09174(.A1(new_n12059_), .A2(new_n12049_), .B(new_n12072_), .ZN(new_n12073_));
  XOR2_X1    g09175(.A1(new_n12058_), .A2(new_n12056_), .Z(new_n12074_));
  OAI21_X1   g09176(.A1(new_n11975_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n12075_));
  OR3_X2     g09177(.A1(new_n12070_), .A2(new_n12060_), .A3(new_n12075_), .Z(new_n12076_));
  AOI21_X1   g09178(.A1(new_n12074_), .A2(pi1157), .B(new_n12076_), .ZN(new_n12077_));
  NOR3_X1    g09179(.A1(new_n12073_), .A2(new_n12077_), .A3(new_n12048_), .ZN(new_n12078_));
  NOR2_X1    g09180(.A1(new_n12078_), .A2(new_n12047_), .ZN(new_n12079_));
  INV_X1     g09181(.I(new_n12079_), .ZN(new_n12080_));
  INV_X1     g09182(.I(pi1160), .ZN(new_n12081_));
  INV_X1     g09183(.I(pi0644), .ZN(new_n12082_));
  AOI21_X1   g09184(.A1(new_n12079_), .A2(new_n12082_), .B(pi0715), .ZN(new_n12083_));
  INV_X1     g09185(.I(new_n12069_), .ZN(new_n12084_));
  NAND3_X1   g09186(.A1(new_n11975_), .A2(new_n12061_), .A3(new_n12049_), .ZN(new_n12085_));
  MUX2_X1    g09187(.I0(new_n12085_), .I1(new_n12084_), .S(new_n12048_), .Z(new_n12086_));
  OR3_X2     g09188(.A1(new_n12083_), .A2(new_n12082_), .A3(new_n12086_), .Z(new_n12087_));
  NOR2_X1    g09189(.A1(new_n12049_), .A2(pi0630), .ZN(new_n12088_));
  NOR2_X1    g09190(.A1(new_n12060_), .A2(pi1157), .ZN(new_n12089_));
  NOR2_X1    g09191(.A1(new_n12088_), .A2(new_n12089_), .ZN(new_n12090_));
  NOR2_X1    g09192(.A1(new_n12090_), .A2(new_n12048_), .ZN(new_n12091_));
  INV_X1     g09193(.I(new_n12091_), .ZN(new_n12092_));
  NOR2_X1    g09194(.A1(new_n12092_), .A2(new_n11975_), .ZN(new_n12093_));
  AOI21_X1   g09195(.A1(new_n12056_), .A2(new_n12092_), .B(new_n12093_), .ZN(new_n12094_));
  NOR2_X1    g09196(.A1(new_n12082_), .A2(pi0715), .ZN(new_n12095_));
  INV_X1     g09197(.I(new_n12095_), .ZN(new_n12096_));
  AOI21_X1   g09198(.A1(new_n11871_), .A2(pi0644), .B(new_n12096_), .ZN(new_n12097_));
  AOI21_X1   g09199(.A1(new_n12094_), .A2(new_n12097_), .B(pi1160), .ZN(new_n12098_));
  INV_X1     g09200(.I(pi0715), .ZN(new_n12099_));
  NAND4_X1   g09201(.A1(new_n12080_), .A2(pi0644), .A3(new_n12099_), .A4(new_n12086_), .ZN(new_n12100_));
  INV_X1     g09202(.I(new_n12094_), .ZN(new_n12101_));
  OAI21_X1   g09203(.A1(pi0644), .A2(new_n11871_), .B(new_n12101_), .ZN(new_n12102_));
  NAND3_X1   g09204(.A1(new_n12094_), .A2(new_n12082_), .A3(new_n11871_), .ZN(new_n12103_));
  NAND4_X1   g09205(.A1(new_n12100_), .A2(new_n12099_), .A3(new_n12102_), .A4(new_n12103_), .ZN(new_n12104_));
  AOI22_X1   g09206(.A1(new_n12104_), .A2(new_n12081_), .B1(new_n12087_), .B2(new_n12098_), .ZN(new_n12105_));
  NOR3_X1    g09207(.A1(new_n12105_), .A2(new_n11867_), .A3(new_n12080_), .ZN(new_n12106_));
  AOI21_X1   g09208(.A1(new_n12105_), .A2(pi0790), .B(new_n12079_), .ZN(new_n12107_));
  OAI21_X1   g09209(.A1(new_n12106_), .A2(new_n12107_), .B(pi0832), .ZN(new_n12108_));
  NOR3_X1    g09210(.A1(new_n7945_), .A2(new_n2489_), .A3(new_n2926_), .ZN(new_n12109_));
  INV_X1     g09211(.I(new_n12109_), .ZN(new_n12110_));
  NOR2_X1    g09212(.A1(new_n11874_), .A2(new_n11883_), .ZN(new_n12111_));
  INV_X1     g09213(.I(new_n12111_), .ZN(new_n12112_));
  NOR2_X1    g09214(.A1(new_n12112_), .A2(new_n5095_), .ZN(new_n12113_));
  INV_X1     g09215(.I(new_n12113_), .ZN(new_n12114_));
  NOR2_X1    g09216(.A1(new_n12110_), .A2(new_n12114_), .ZN(new_n12115_));
  INV_X1     g09217(.I(pi0761), .ZN(new_n12116_));
  NOR3_X1    g09218(.A1(new_n12109_), .A2(pi0140), .A3(new_n12116_), .ZN(new_n12117_));
  NOR2_X1    g09219(.A1(new_n11894_), .A2(new_n11874_), .ZN(new_n12118_));
  OAI21_X1   g09220(.A1(new_n12118_), .A2(new_n11876_), .B(pi0140), .ZN(new_n12119_));
  OAI21_X1   g09221(.A1(new_n12119_), .A2(new_n2491_), .B(new_n12116_), .ZN(new_n12120_));
  NOR3_X1    g09222(.A1(new_n12110_), .A2(new_n11874_), .A3(new_n11884_), .ZN(new_n12121_));
  INV_X1     g09223(.I(new_n12121_), .ZN(new_n12122_));
  NAND2_X1   g09224(.A1(new_n12122_), .A2(new_n7339_), .ZN(new_n12123_));
  AOI22_X1   g09225(.A1(new_n12123_), .A2(new_n12120_), .B1(new_n12115_), .B2(new_n12117_), .ZN(new_n12124_));
  MUX2_X1    g09226(.I0(new_n12124_), .I1(pi0140), .S(pi0039), .Z(new_n12125_));
  INV_X1     g09227(.I(new_n12125_), .ZN(new_n12126_));
  NOR2_X1    g09228(.A1(pi0661), .A2(pi0681), .ZN(new_n12127_));
  INV_X1     g09229(.I(new_n12127_), .ZN(new_n12128_));
  NOR2_X1    g09230(.A1(new_n12128_), .A2(pi0662), .ZN(new_n12129_));
  NOR2_X1    g09231(.A1(new_n12129_), .A2(new_n5095_), .ZN(new_n12130_));
  NOR2_X1    g09232(.A1(new_n8648_), .A2(pi0287), .ZN(new_n12131_));
  NOR3_X1    g09233(.A1(new_n10267_), .A2(new_n2923_), .A3(new_n2924_), .ZN(new_n12132_));
  INV_X1     g09234(.I(new_n12132_), .ZN(new_n12133_));
  NOR2_X1    g09235(.A1(new_n12133_), .A2(new_n5108_), .ZN(new_n12134_));
  INV_X1     g09236(.I(new_n12134_), .ZN(new_n12135_));
  AOI21_X1   g09237(.A1(new_n12109_), .A2(new_n10267_), .B(pi1091), .ZN(new_n12136_));
  NAND3_X1   g09238(.A1(new_n7860_), .A2(new_n2488_), .A3(new_n8018_), .ZN(new_n12137_));
  NOR4_X1    g09239(.A1(new_n2459_), .A2(new_n2476_), .A3(new_n2482_), .A4(new_n12137_), .ZN(new_n12138_));
  NOR2_X1    g09240(.A1(new_n2928_), .A2(pi0824), .ZN(new_n12139_));
  OAI21_X1   g09241(.A1(new_n12138_), .A2(new_n12139_), .B(pi1092), .ZN(new_n12140_));
  INV_X1     g09242(.I(new_n12131_), .ZN(new_n12141_));
  OAI21_X1   g09243(.A1(new_n7945_), .A2(new_n2489_), .B(new_n12141_), .ZN(new_n12142_));
  NAND4_X1   g09244(.A1(new_n12140_), .A2(new_n5366_), .A3(new_n12142_), .A4(pi1093), .ZN(new_n12143_));
  AOI21_X1   g09245(.A1(new_n12143_), .A2(new_n10267_), .B(new_n12136_), .ZN(new_n12144_));
  INV_X1     g09246(.I(new_n12144_), .ZN(new_n12145_));
  NAND3_X1   g09247(.A1(new_n12140_), .A2(new_n5366_), .A3(new_n12142_), .ZN(new_n12146_));
  NOR3_X1    g09248(.A1(new_n6036_), .A2(pi0829), .A3(new_n2923_), .ZN(new_n12147_));
  AOI21_X1   g09249(.A1(new_n12138_), .A2(new_n12147_), .B(pi0829), .ZN(new_n12148_));
  NAND2_X1   g09250(.A1(new_n2490_), .A2(new_n12131_), .ZN(new_n12149_));
  NAND2_X1   g09251(.A1(new_n2925_), .A2(new_n2920_), .ZN(new_n12150_));
  NOR2_X1    g09252(.A1(new_n12149_), .A2(new_n12150_), .ZN(new_n12151_));
  AOI21_X1   g09253(.A1(new_n12146_), .A2(new_n12148_), .B(new_n12151_), .ZN(new_n12152_));
  NOR2_X1    g09254(.A1(new_n12109_), .A2(new_n10267_), .ZN(new_n12153_));
  NOR2_X1    g09255(.A1(new_n12153_), .A2(pi0120), .ZN(new_n12154_));
  OAI21_X1   g09256(.A1(new_n12152_), .A2(new_n2918_), .B(new_n12154_), .ZN(new_n12155_));
  NAND2_X1   g09257(.A1(new_n12155_), .A2(new_n12145_), .ZN(new_n12156_));
  OAI21_X1   g09258(.A1(new_n12156_), .A2(new_n5108_), .B(new_n12135_), .ZN(new_n12157_));
  INV_X1     g09259(.I(new_n12157_), .ZN(new_n12158_));
  NOR2_X1    g09260(.A1(new_n12133_), .A2(new_n11883_), .ZN(new_n12159_));
  INV_X1     g09261(.I(new_n12159_), .ZN(new_n12160_));
  OAI21_X1   g09262(.A1(new_n12155_), .A2(pi0665), .B(new_n12145_), .ZN(new_n12161_));
  NAND2_X1   g09263(.A1(new_n12161_), .A2(new_n12160_), .ZN(new_n12162_));
  NOR2_X1    g09264(.A1(new_n12162_), .A2(new_n11874_), .ZN(new_n12163_));
  NOR2_X1    g09265(.A1(new_n12163_), .A2(new_n12158_), .ZN(new_n12164_));
  INV_X1     g09266(.I(new_n12164_), .ZN(new_n12165_));
  INV_X1     g09267(.I(pi0616), .ZN(new_n12166_));
  NOR2_X1    g09268(.A1(pi0614), .A2(pi0642), .ZN(new_n12167_));
  NAND2_X1   g09269(.A1(new_n12167_), .A2(new_n12166_), .ZN(new_n12168_));
  NAND2_X1   g09270(.A1(new_n12162_), .A2(new_n12157_), .ZN(new_n12169_));
  OAI21_X1   g09271(.A1(new_n12155_), .A2(pi0621), .B(new_n12145_), .ZN(new_n12170_));
  NAND4_X1   g09272(.A1(new_n2483_), .A2(new_n2484_), .A3(new_n2486_), .A4(new_n8018_), .ZN(new_n12171_));
  NOR2_X1    g09273(.A1(new_n7861_), .A2(new_n12171_), .ZN(new_n12172_));
  NAND4_X1   g09274(.A1(new_n5268_), .A2(new_n2475_), .A3(new_n2481_), .A4(new_n12172_), .ZN(new_n12173_));
  INV_X1     g09275(.I(new_n12139_), .ZN(new_n12174_));
  AOI21_X1   g09276(.A1(new_n12173_), .A2(new_n12174_), .B(new_n2923_), .ZN(new_n12175_));
  OAI21_X1   g09277(.A1(new_n2490_), .A2(new_n12131_), .B(new_n5366_), .ZN(new_n12176_));
  OAI21_X1   g09278(.A1(new_n12175_), .A2(new_n12176_), .B(new_n12148_), .ZN(new_n12177_));
  NAND4_X1   g09279(.A1(new_n2490_), .A2(new_n2920_), .A3(new_n2925_), .A4(new_n12131_), .ZN(new_n12178_));
  NAND2_X1   g09280(.A1(new_n12177_), .A2(new_n12178_), .ZN(new_n12179_));
  INV_X1     g09281(.I(new_n12154_), .ZN(new_n12180_));
  AOI21_X1   g09282(.A1(new_n12179_), .A2(pi1091), .B(new_n12180_), .ZN(new_n12181_));
  NAND2_X1   g09283(.A1(new_n12181_), .A2(new_n11873_), .ZN(new_n12182_));
  NOR2_X1    g09284(.A1(new_n12182_), .A2(pi0665), .ZN(new_n12183_));
  NOR2_X1    g09285(.A1(new_n12183_), .A2(new_n12170_), .ZN(new_n12184_));
  MUX2_X1    g09286(.I0(new_n12184_), .I1(new_n12169_), .S(new_n5101_), .Z(new_n12185_));
  NOR3_X1    g09287(.A1(new_n12185_), .A2(new_n12165_), .A3(new_n12168_), .ZN(new_n12186_));
  INV_X1     g09288(.I(new_n12168_), .ZN(new_n12187_));
  AOI21_X1   g09289(.A1(new_n12185_), .A2(new_n12187_), .B(new_n12164_), .ZN(new_n12188_));
  OR2_X2     g09290(.A1(new_n12186_), .A2(new_n12188_), .Z(new_n12189_));
  INV_X1     g09291(.I(new_n5461_), .ZN(new_n12190_));
  NOR2_X1    g09292(.A1(new_n12181_), .A2(new_n12144_), .ZN(new_n12191_));
  NOR2_X1    g09293(.A1(new_n12190_), .A2(new_n12132_), .ZN(new_n12192_));
  NAND3_X1   g09294(.A1(new_n12191_), .A2(new_n12190_), .A3(new_n12192_), .ZN(new_n12193_));
  INV_X1     g09295(.I(new_n12192_), .ZN(new_n12194_));
  OAI21_X1   g09296(.A1(new_n12156_), .A2(new_n5461_), .B(new_n12194_), .ZN(new_n12195_));
  NAND2_X1   g09297(.A1(new_n12193_), .A2(new_n12195_), .ZN(new_n12196_));
  NOR2_X1    g09298(.A1(new_n12191_), .A2(new_n5217_), .ZN(new_n12197_));
  AOI21_X1   g09299(.A1(new_n12196_), .A2(new_n5217_), .B(new_n12197_), .ZN(new_n12198_));
  NOR2_X1    g09300(.A1(new_n12198_), .A2(new_n11875_), .ZN(new_n12199_));
  NOR2_X1    g09301(.A1(new_n12161_), .A2(new_n5217_), .ZN(new_n12200_));
  NOR3_X1    g09302(.A1(new_n12199_), .A2(new_n12130_), .A3(new_n12200_), .ZN(new_n12201_));
  INV_X1     g09303(.I(new_n12201_), .ZN(new_n12202_));
  AOI21_X1   g09304(.A1(new_n12189_), .A2(new_n12130_), .B(new_n12202_), .ZN(new_n12203_));
  AND2_X2    g09305(.A1(new_n12203_), .A2(new_n6460_), .Z(new_n12204_));
  MUX2_X1    g09306(.I0(new_n12156_), .I1(new_n12133_), .S(new_n5109_), .Z(new_n12205_));
  NOR2_X1    g09307(.A1(new_n12205_), .A2(new_n11874_), .ZN(new_n12206_));
  INV_X1     g09308(.I(new_n12206_), .ZN(new_n12207_));
  NOR2_X1    g09309(.A1(new_n11875_), .A2(new_n12133_), .ZN(new_n12208_));
  INV_X1     g09310(.I(new_n12208_), .ZN(new_n12209_));
  AOI21_X1   g09311(.A1(new_n12168_), .A2(new_n12209_), .B(new_n12207_), .ZN(new_n12210_));
  NOR3_X1    g09312(.A1(new_n11875_), .A2(new_n12133_), .A3(new_n12187_), .ZN(new_n12211_));
  INV_X1     g09313(.I(new_n11873_), .ZN(new_n12212_));
  NOR2_X1    g09314(.A1(new_n12155_), .A2(new_n12212_), .ZN(new_n12213_));
  NOR2_X1    g09315(.A1(new_n12133_), .A2(new_n12212_), .ZN(new_n12214_));
  NOR3_X1    g09316(.A1(new_n12214_), .A2(pi0603), .A3(new_n5109_), .ZN(new_n12215_));
  INV_X1     g09317(.I(new_n12215_), .ZN(new_n12216_));
  NOR2_X1    g09318(.A1(new_n12213_), .A2(new_n12216_), .ZN(new_n12217_));
  NOR2_X1    g09319(.A1(new_n5101_), .A2(pi0665), .ZN(new_n12218_));
  AOI21_X1   g09320(.A1(new_n12159_), .A2(new_n5101_), .B(new_n12218_), .ZN(new_n12219_));
  NOR2_X1    g09321(.A1(new_n12217_), .A2(new_n12219_), .ZN(new_n12220_));
  NOR2_X1    g09322(.A1(new_n12206_), .A2(new_n12220_), .ZN(new_n12221_));
  INV_X1     g09323(.I(new_n12130_), .ZN(new_n12222_));
  INV_X1     g09324(.I(new_n11883_), .ZN(new_n12223_));
  NOR2_X1    g09325(.A1(new_n5101_), .A2(pi0621), .ZN(new_n12224_));
  NOR2_X1    g09326(.A1(new_n12223_), .A2(new_n12224_), .ZN(new_n12225_));
  NOR2_X1    g09327(.A1(new_n12225_), .A2(new_n12133_), .ZN(new_n12226_));
  AOI21_X1   g09328(.A1(new_n12226_), .A2(new_n12168_), .B(new_n12222_), .ZN(new_n12227_));
  NOR3_X1    g09329(.A1(new_n12221_), .A2(new_n12168_), .A3(new_n12227_), .ZN(new_n12228_));
  NOR2_X1    g09330(.A1(new_n12133_), .A2(new_n5109_), .ZN(new_n12229_));
  AOI21_X1   g09331(.A1(new_n12155_), .A2(new_n12145_), .B(new_n5108_), .ZN(new_n12230_));
  NOR2_X1    g09332(.A1(new_n12230_), .A2(new_n12229_), .ZN(new_n12231_));
  NAND3_X1   g09333(.A1(new_n12163_), .A2(new_n5217_), .A3(new_n12231_), .ZN(new_n12232_));
  NAND2_X1   g09334(.A1(new_n12232_), .A2(new_n5095_), .ZN(new_n12233_));
  NOR4_X1    g09335(.A1(new_n12210_), .A2(new_n12228_), .A3(new_n12211_), .A4(new_n12233_), .ZN(new_n12234_));
  NAND3_X1   g09336(.A1(new_n2490_), .A2(new_n2925_), .A3(new_n12131_), .ZN(new_n12235_));
  NAND2_X1   g09337(.A1(new_n12235_), .A2(new_n10267_), .ZN(new_n12236_));
  NOR4_X1    g09338(.A1(new_n5125_), .A2(new_n10267_), .A3(new_n5366_), .A4(pi1091), .ZN(new_n12237_));
  INV_X1     g09339(.I(new_n12237_), .ZN(new_n12238_));
  NAND4_X1   g09340(.A1(new_n5124_), .A2(new_n10267_), .A3(new_n2958_), .A4(new_n8405_), .ZN(new_n12239_));
  AOI21_X1   g09341(.A1(new_n2490_), .A2(new_n2925_), .B(new_n12239_), .ZN(new_n12240_));
  OAI21_X1   g09342(.A1(new_n12240_), .A2(new_n2918_), .B(new_n12238_), .ZN(new_n12241_));
  NAND2_X1   g09343(.A1(new_n12241_), .A2(new_n12236_), .ZN(new_n12242_));
  NOR2_X1    g09344(.A1(new_n12242_), .A2(new_n5108_), .ZN(new_n12243_));
  AOI21_X1   g09345(.A1(new_n12243_), .A2(new_n5106_), .B(new_n12160_), .ZN(new_n12244_));
  NOR2_X1    g09346(.A1(new_n12243_), .A2(new_n12209_), .ZN(new_n12245_));
  NOR4_X1    g09347(.A1(new_n12244_), .A2(new_n12245_), .A3(new_n12187_), .A4(new_n12227_), .ZN(new_n12246_));
  NOR2_X1    g09348(.A1(new_n12132_), .A2(new_n5108_), .ZN(new_n12247_));
  INV_X1     g09349(.I(new_n12247_), .ZN(new_n12248_));
  OAI21_X1   g09350(.A1(new_n12242_), .A2(new_n5109_), .B(new_n12248_), .ZN(new_n12249_));
  NOR2_X1    g09351(.A1(new_n12249_), .A2(new_n12209_), .ZN(new_n12250_));
  NAND2_X1   g09352(.A1(new_n12243_), .A2(new_n12187_), .ZN(new_n12251_));
  AOI21_X1   g09353(.A1(new_n5217_), .A2(new_n12251_), .B(new_n12250_), .ZN(new_n12252_));
  NOR2_X1    g09354(.A1(new_n12252_), .A2(new_n12245_), .ZN(new_n12253_));
  OAI21_X1   g09355(.A1(new_n12243_), .A2(new_n12160_), .B(new_n12129_), .ZN(new_n12254_));
  NAND2_X1   g09356(.A1(new_n12254_), .A2(pi0680), .ZN(new_n12255_));
  INV_X1     g09357(.I(new_n12255_), .ZN(new_n12256_));
  AOI21_X1   g09358(.A1(new_n12253_), .A2(new_n12256_), .B(new_n12246_), .ZN(new_n12257_));
  NOR2_X1    g09359(.A1(new_n12249_), .A2(new_n12160_), .ZN(new_n12258_));
  NAND3_X1   g09360(.A1(new_n12256_), .A2(new_n12244_), .A3(new_n12258_), .ZN(new_n12259_));
  NAND2_X1   g09361(.A1(new_n12259_), .A2(new_n6460_), .ZN(new_n12260_));
  OAI21_X1   g09362(.A1(new_n12109_), .A2(new_n12239_), .B(pi1091), .ZN(new_n12261_));
  AOI22_X1   g09363(.A1(new_n12261_), .A2(new_n12238_), .B1(new_n10267_), .B2(new_n12235_), .ZN(new_n12262_));
  NOR2_X1    g09364(.A1(new_n12262_), .A2(new_n12209_), .ZN(new_n12263_));
  OR2_X2     g09365(.A1(new_n12252_), .A2(new_n12263_), .Z(new_n12264_));
  NOR2_X1    g09366(.A1(new_n12264_), .A2(pi0223), .ZN(new_n12265_));
  NAND2_X1   g09367(.A1(new_n12265_), .A2(new_n12260_), .ZN(new_n12266_));
  NAND3_X1   g09368(.A1(new_n12266_), .A2(new_n5141_), .A3(new_n12257_), .ZN(new_n12267_));
  NOR2_X1    g09369(.A1(new_n12118_), .A2(new_n11876_), .ZN(new_n12268_));
  NOR3_X1    g09370(.A1(new_n12268_), .A2(new_n2614_), .A3(new_n12133_), .ZN(new_n12269_));
  INV_X1     g09371(.I(new_n12269_), .ZN(new_n12270_));
  AND3_X2    g09372(.A1(new_n12267_), .A2(new_n10243_), .A3(new_n12270_), .Z(new_n12271_));
  OAI21_X1   g09373(.A1(new_n12234_), .A2(new_n6460_), .B(new_n12271_), .ZN(new_n12272_));
  OAI21_X1   g09374(.A1(new_n12118_), .A2(new_n11876_), .B(new_n3284_), .ZN(new_n12273_));
  OAI21_X1   g09375(.A1(new_n12273_), .A2(new_n12133_), .B(new_n2566_), .ZN(new_n12274_));
  AOI21_X1   g09376(.A1(new_n12274_), .A2(new_n3284_), .B(new_n2587_), .ZN(new_n12275_));
  INV_X1     g09377(.I(new_n12275_), .ZN(new_n12276_));
  OAI21_X1   g09378(.A1(new_n12204_), .A2(new_n12272_), .B(new_n12276_), .ZN(new_n12277_));
  NOR2_X1    g09379(.A1(new_n12240_), .A2(new_n2918_), .ZN(new_n12278_));
  NAND2_X1   g09380(.A1(new_n12278_), .A2(new_n12236_), .ZN(new_n12279_));
  NOR2_X1    g09381(.A1(new_n12279_), .A2(new_n11882_), .ZN(new_n12280_));
  NOR2_X1    g09382(.A1(new_n12133_), .A2(new_n12223_), .ZN(new_n12281_));
  INV_X1     g09383(.I(new_n12281_), .ZN(new_n12282_));
  NOR2_X1    g09384(.A1(new_n12282_), .A2(new_n5109_), .ZN(new_n12283_));
  AOI21_X1   g09385(.A1(new_n12280_), .A2(new_n5109_), .B(new_n12283_), .ZN(new_n12284_));
  NOR3_X1    g09386(.A1(new_n12284_), .A2(new_n5217_), .A3(new_n12224_), .ZN(new_n12285_));
  NOR2_X1    g09387(.A1(new_n12133_), .A2(new_n11874_), .ZN(new_n12286_));
  INV_X1     g09388(.I(new_n12286_), .ZN(new_n12287_));
  NOR2_X1    g09389(.A1(new_n12287_), .A2(new_n12187_), .ZN(new_n12288_));
  INV_X1     g09390(.I(new_n12288_), .ZN(new_n12289_));
  NAND3_X1   g09391(.A1(new_n12278_), .A2(new_n12236_), .A3(pi0621), .ZN(new_n12290_));
  NAND2_X1   g09392(.A1(new_n12290_), .A2(new_n5109_), .ZN(new_n12291_));
  INV_X1     g09393(.I(new_n12214_), .ZN(new_n12292_));
  AOI21_X1   g09394(.A1(new_n12292_), .A2(new_n5108_), .B(pi0603), .ZN(new_n12293_));
  NAND2_X1   g09395(.A1(new_n12291_), .A2(new_n12293_), .ZN(new_n12294_));
  NOR2_X1    g09396(.A1(new_n12132_), .A2(pi0603), .ZN(new_n12295_));
  NOR2_X1    g09397(.A1(new_n12295_), .A2(new_n12168_), .ZN(new_n12296_));
  NAND2_X1   g09398(.A1(new_n12294_), .A2(new_n12296_), .ZN(new_n12297_));
  NAND2_X1   g09399(.A1(new_n12297_), .A2(new_n12289_), .ZN(new_n12298_));
  NAND2_X1   g09400(.A1(new_n12298_), .A2(new_n5217_), .ZN(new_n12299_));
  NOR2_X1    g09401(.A1(new_n12299_), .A2(new_n11884_), .ZN(new_n12300_));
  NOR2_X1    g09402(.A1(new_n12300_), .A2(new_n12285_), .ZN(new_n12301_));
  INV_X1     g09403(.I(new_n12280_), .ZN(new_n12302_));
  NOR2_X1    g09404(.A1(new_n12135_), .A2(new_n12223_), .ZN(new_n12303_));
  INV_X1     g09405(.I(new_n12303_), .ZN(new_n12304_));
  NAND2_X1   g09406(.A1(new_n12302_), .A2(new_n12304_), .ZN(new_n12305_));
  AOI21_X1   g09407(.A1(new_n12298_), .A2(new_n12305_), .B(new_n12222_), .ZN(new_n12306_));
  NOR2_X1    g09408(.A1(new_n11874_), .A2(new_n2926_), .ZN(new_n12307_));
  INV_X1     g09409(.I(new_n12307_), .ZN(new_n12308_));
  NOR2_X1    g09410(.A1(new_n12249_), .A2(new_n12308_), .ZN(new_n12309_));
  INV_X1     g09411(.I(new_n12309_), .ZN(new_n12310_));
  INV_X1     g09412(.I(new_n12279_), .ZN(new_n12311_));
  NOR2_X1    g09413(.A1(new_n12311_), .A2(new_n5427_), .ZN(new_n12312_));
  NAND2_X1   g09414(.A1(new_n12310_), .A2(new_n12312_), .ZN(new_n12313_));
  AOI21_X1   g09415(.A1(new_n5217_), .A2(new_n12224_), .B(pi0680), .ZN(new_n12314_));
  NAND2_X1   g09416(.A1(new_n12313_), .A2(new_n12314_), .ZN(new_n12315_));
  NOR2_X1    g09417(.A1(new_n12306_), .A2(new_n12315_), .ZN(new_n12316_));
  NAND4_X1   g09418(.A1(new_n12301_), .A2(new_n2604_), .A3(new_n5141_), .A4(new_n12316_), .ZN(new_n12317_));
  NOR2_X1    g09419(.A1(new_n12155_), .A2(new_n12223_), .ZN(new_n12318_));
  NOR4_X1    g09420(.A1(new_n12318_), .A2(new_n5101_), .A3(pi0621), .A4(new_n5100_), .ZN(new_n12319_));
  INV_X1     g09421(.I(new_n12225_), .ZN(new_n12320_));
  INV_X1     g09422(.I(new_n12318_), .ZN(new_n12321_));
  OAI22_X1   g09423(.A1(new_n12321_), .A2(new_n5461_), .B1(new_n5427_), .B2(new_n12303_), .ZN(new_n12322_));
  NOR3_X1    g09424(.A1(new_n12322_), .A2(new_n12130_), .A3(new_n12320_), .ZN(new_n12323_));
  NOR3_X1    g09425(.A1(new_n12156_), .A2(new_n5461_), .A3(new_n12194_), .ZN(new_n12324_));
  AOI21_X1   g09426(.A1(new_n12191_), .A2(new_n12190_), .B(new_n12192_), .ZN(new_n12325_));
  NOR2_X1    g09427(.A1(new_n12325_), .A2(new_n12324_), .ZN(new_n12326_));
  NOR2_X1    g09428(.A1(new_n12326_), .A2(new_n11874_), .ZN(new_n12327_));
  OAI22_X1   g09429(.A1(pi0680), .A2(new_n12327_), .B1(new_n12323_), .B2(new_n12319_), .ZN(new_n12328_));
  AOI21_X1   g09430(.A1(new_n12318_), .A2(new_n5109_), .B(new_n12283_), .ZN(new_n12329_));
  NOR3_X1    g09431(.A1(new_n12329_), .A2(new_n5100_), .A3(new_n12320_), .ZN(new_n12330_));
  NOR2_X1    g09432(.A1(new_n12282_), .A2(new_n12224_), .ZN(new_n12331_));
  NOR4_X1    g09433(.A1(new_n12130_), .A2(new_n12223_), .A3(new_n12168_), .A4(new_n12295_), .ZN(new_n12332_));
  INV_X1     g09434(.I(new_n12332_), .ZN(new_n12333_));
  NOR2_X1    g09435(.A1(new_n12217_), .A2(new_n12333_), .ZN(new_n12334_));
  OAI21_X1   g09436(.A1(new_n12168_), .A2(new_n12295_), .B(new_n12217_), .ZN(new_n12335_));
  NAND3_X1   g09437(.A1(new_n12335_), .A2(new_n5095_), .A3(new_n12289_), .ZN(new_n12336_));
  NOR3_X1    g09438(.A1(new_n12336_), .A2(new_n12330_), .A3(new_n12334_), .ZN(new_n12337_));
  MUX2_X1    g09439(.I0(new_n12337_), .I1(new_n12328_), .S(new_n6460_), .Z(new_n12338_));
  INV_X1     g09440(.I(new_n12149_), .ZN(new_n12339_));
  NOR2_X1    g09441(.A1(new_n12339_), .A2(pi0120), .ZN(new_n12340_));
  NOR3_X1    g09442(.A1(new_n12122_), .A2(new_n12340_), .A3(new_n3155_), .ZN(new_n12341_));
  OAI22_X1   g09443(.A1(new_n12338_), .A2(new_n2614_), .B1(pi0223), .B2(new_n12341_), .ZN(new_n12342_));
  AOI21_X1   g09444(.A1(new_n12342_), .A2(new_n12317_), .B(pi0299), .ZN(new_n12343_));
  NAND4_X1   g09445(.A1(new_n12301_), .A2(new_n2566_), .A3(new_n5094_), .A4(new_n12316_), .ZN(new_n12344_));
  MUX2_X1    g09446(.I0(new_n12337_), .I1(new_n12328_), .S(new_n6445_), .Z(new_n12345_));
  NOR3_X1    g09447(.A1(new_n12122_), .A2(new_n12340_), .A3(new_n3285_), .ZN(new_n12346_));
  OAI22_X1   g09448(.A1(new_n12345_), .A2(new_n3284_), .B1(pi0215), .B2(new_n12346_), .ZN(new_n12347_));
  AOI21_X1   g09449(.A1(new_n12347_), .A2(new_n12344_), .B(new_n2587_), .ZN(new_n12348_));
  NOR2_X1    g09450(.A1(new_n12343_), .A2(new_n12348_), .ZN(new_n12349_));
  NOR3_X1    g09451(.A1(new_n12277_), .A2(new_n7339_), .A3(new_n12116_), .ZN(new_n12350_));
  NOR3_X1    g09452(.A1(new_n12263_), .A2(new_n12280_), .A3(new_n5217_), .ZN(new_n12351_));
  NOR3_X1    g09453(.A1(new_n12305_), .A2(new_n12187_), .A3(new_n12250_), .ZN(new_n12352_));
  NOR2_X1    g09454(.A1(new_n12304_), .A2(pi0603), .ZN(new_n12353_));
  NOR3_X1    g09455(.A1(new_n12263_), .A2(new_n12280_), .A3(new_n12353_), .ZN(new_n12354_));
  NOR2_X1    g09456(.A1(new_n12354_), .A2(new_n12168_), .ZN(new_n12355_));
  XOR2_X1    g09457(.A1(new_n12352_), .A2(new_n12355_), .Z(new_n12356_));
  NOR2_X1    g09458(.A1(new_n12356_), .A2(new_n12222_), .ZN(new_n12357_));
  NOR2_X1    g09459(.A1(new_n5103_), .A2(new_n5108_), .ZN(new_n12358_));
  INV_X1     g09460(.I(new_n12358_), .ZN(new_n12359_));
  MUX2_X1    g09461(.I0(new_n12242_), .I1(new_n12132_), .S(new_n12359_), .Z(new_n12360_));
  NOR3_X1    g09462(.A1(new_n12360_), .A2(pi0614), .A3(pi0616), .ZN(new_n12361_));
  NOR2_X1    g09463(.A1(new_n12361_), .A2(new_n12249_), .ZN(new_n12362_));
  OAI22_X1   g09464(.A1(new_n12357_), .A2(new_n12351_), .B1(pi0680), .B2(new_n12362_), .ZN(new_n12363_));
  AOI22_X1   g09465(.A1(new_n12241_), .A2(new_n12236_), .B1(new_n12133_), .B2(new_n12359_), .ZN(new_n12364_));
  INV_X1     g09466(.I(new_n12364_), .ZN(new_n12365_));
  NAND4_X1   g09467(.A1(new_n12241_), .A2(new_n12236_), .A3(new_n12132_), .A4(new_n12359_), .ZN(new_n12366_));
  NAND4_X1   g09468(.A1(new_n12365_), .A2(new_n5105_), .A3(new_n12133_), .A4(new_n12366_), .ZN(new_n12367_));
  NOR3_X1    g09469(.A1(new_n12262_), .A2(new_n12132_), .A3(new_n12359_), .ZN(new_n12368_));
  NAND4_X1   g09470(.A1(new_n12241_), .A2(new_n12236_), .A3(new_n12132_), .A4(new_n12358_), .ZN(new_n12369_));
  NAND2_X1   g09471(.A1(new_n12369_), .A2(new_n5105_), .ZN(new_n12370_));
  OAI21_X1   g09472(.A1(new_n12370_), .A2(new_n12368_), .B(new_n12132_), .ZN(new_n12371_));
  NAND2_X1   g09473(.A1(new_n12367_), .A2(new_n12371_), .ZN(new_n12372_));
  NOR2_X1    g09474(.A1(new_n12372_), .A2(pi0680), .ZN(new_n12373_));
  INV_X1     g09475(.I(new_n12373_), .ZN(new_n12374_));
  INV_X1     g09476(.I(new_n12245_), .ZN(new_n12375_));
  NAND3_X1   g09477(.A1(new_n12375_), .A2(new_n5100_), .A3(new_n12284_), .ZN(new_n12376_));
  NAND2_X1   g09478(.A1(new_n12374_), .A2(new_n12376_), .ZN(new_n12377_));
  NOR2_X1    g09479(.A1(new_n12111_), .A2(new_n12133_), .ZN(new_n12378_));
  NOR2_X1    g09480(.A1(new_n12378_), .A2(new_n12166_), .ZN(new_n12379_));
  INV_X1     g09481(.I(new_n12379_), .ZN(new_n12380_));
  NOR2_X1    g09482(.A1(new_n12245_), .A2(pi0642), .ZN(new_n12381_));
  INV_X1     g09483(.I(new_n12284_), .ZN(new_n12382_));
  NOR2_X1    g09484(.A1(new_n12382_), .A2(new_n12354_), .ZN(new_n12383_));
  INV_X1     g09485(.I(pi0642), .ZN(new_n12384_));
  OAI21_X1   g09486(.A1(new_n12378_), .A2(new_n12384_), .B(pi0614), .ZN(new_n12385_));
  AOI21_X1   g09487(.A1(new_n12383_), .A2(new_n12381_), .B(new_n12385_), .ZN(new_n12386_));
  NAND2_X1   g09488(.A1(new_n12378_), .A2(pi0614), .ZN(new_n12387_));
  INV_X1     g09489(.I(new_n12387_), .ZN(new_n12388_));
  NOR3_X1    g09490(.A1(new_n12386_), .A2(pi0616), .A3(new_n12388_), .ZN(new_n12389_));
  NAND2_X1   g09491(.A1(new_n12389_), .A2(new_n12380_), .ZN(new_n12390_));
  NAND3_X1   g09492(.A1(new_n12390_), .A2(new_n12130_), .A3(new_n12377_), .ZN(new_n12391_));
  INV_X1     g09493(.I(new_n12391_), .ZN(new_n12392_));
  NAND3_X1   g09494(.A1(new_n12392_), .A2(new_n5141_), .A3(new_n12363_), .ZN(new_n12393_));
  AOI21_X1   g09495(.A1(new_n5141_), .A2(new_n12391_), .B(new_n12363_), .ZN(new_n12394_));
  INV_X1     g09496(.I(new_n12394_), .ZN(new_n12395_));
  AOI21_X1   g09497(.A1(new_n12395_), .A2(new_n12393_), .B(new_n2604_), .ZN(new_n12396_));
  NOR2_X1    g09498(.A1(new_n5108_), .A2(new_n5101_), .ZN(new_n12397_));
  INV_X1     g09499(.I(new_n12397_), .ZN(new_n12398_));
  NOR4_X1    g09500(.A1(new_n12156_), .A2(new_n12384_), .A3(new_n12133_), .A4(new_n12398_), .ZN(new_n12399_));
  AOI22_X1   g09501(.A1(new_n12155_), .A2(new_n12145_), .B1(new_n12133_), .B2(new_n12398_), .ZN(new_n12400_));
  INV_X1     g09502(.I(new_n12400_), .ZN(new_n12401_));
  NAND4_X1   g09503(.A1(new_n12155_), .A2(new_n12145_), .A3(new_n12132_), .A4(new_n12398_), .ZN(new_n12402_));
  AOI22_X1   g09504(.A1(new_n12401_), .A2(new_n12402_), .B1(pi0642), .B2(new_n12133_), .ZN(new_n12403_));
  OAI21_X1   g09505(.A1(new_n12403_), .A2(new_n12399_), .B(new_n12112_), .ZN(new_n12404_));
  NAND2_X1   g09506(.A1(new_n12404_), .A2(pi0614), .ZN(new_n12405_));
  NAND4_X1   g09507(.A1(new_n12405_), .A2(new_n12166_), .A3(new_n12380_), .A4(new_n12387_), .ZN(new_n12406_));
  NOR4_X1    g09508(.A1(new_n12230_), .A2(new_n5103_), .A3(new_n12132_), .A4(new_n12229_), .ZN(new_n12407_));
  INV_X1     g09509(.I(new_n12229_), .ZN(new_n12408_));
  OAI21_X1   g09510(.A1(new_n12181_), .A2(new_n12144_), .B(new_n5109_), .ZN(new_n12409_));
  AOI22_X1   g09511(.A1(new_n12409_), .A2(new_n12408_), .B1(new_n5102_), .B2(new_n12132_), .ZN(new_n12410_));
  NOR2_X1    g09512(.A1(new_n12410_), .A2(new_n12407_), .ZN(new_n12411_));
  MUX2_X1    g09513(.I0(new_n12411_), .I1(new_n12132_), .S(new_n5104_), .Z(new_n12412_));
  AOI21_X1   g09514(.A1(new_n12156_), .A2(new_n5109_), .B(new_n12132_), .ZN(new_n12413_));
  NOR3_X1    g09515(.A1(new_n12156_), .A2(new_n5108_), .A3(new_n12133_), .ZN(new_n12414_));
  OAI21_X1   g09516(.A1(new_n12414_), .A2(new_n12413_), .B(pi0603), .ZN(new_n12415_));
  INV_X1     g09517(.I(new_n12283_), .ZN(new_n12416_));
  NAND2_X1   g09518(.A1(new_n11873_), .A2(new_n12218_), .ZN(new_n12417_));
  NAND3_X1   g09519(.A1(new_n12416_), .A2(new_n5101_), .A3(new_n12417_), .ZN(new_n12418_));
  AOI21_X1   g09520(.A1(new_n12321_), .A2(new_n5108_), .B(new_n12418_), .ZN(new_n12419_));
  AOI21_X1   g09521(.A1(new_n12415_), .A2(new_n12419_), .B(new_n5217_), .ZN(new_n12420_));
  INV_X1     g09522(.I(new_n12420_), .ZN(new_n12421_));
  OAI21_X1   g09523(.A1(new_n12412_), .A2(pi0680), .B(new_n12421_), .ZN(new_n12422_));
  AOI21_X1   g09524(.A1(new_n12130_), .A2(new_n12406_), .B(new_n12422_), .ZN(new_n12423_));
  NAND2_X1   g09525(.A1(new_n12326_), .A2(new_n5095_), .ZN(new_n12424_));
  NOR3_X1    g09526(.A1(new_n12145_), .A2(pi0603), .A3(pi0621), .ZN(new_n12425_));
  INV_X1     g09527(.I(new_n12425_), .ZN(new_n12426_));
  NAND2_X1   g09528(.A1(new_n12319_), .A2(new_n12426_), .ZN(new_n12427_));
  NAND2_X1   g09529(.A1(new_n12424_), .A2(new_n12427_), .ZN(new_n12428_));
  NAND4_X1   g09530(.A1(new_n12428_), .A2(new_n12112_), .A3(new_n12222_), .A4(new_n12196_), .ZN(new_n12429_));
  INV_X1     g09531(.I(new_n12429_), .ZN(new_n12430_));
  NOR2_X1    g09532(.A1(new_n6460_), .A2(new_n3155_), .ZN(new_n12431_));
  NOR2_X1    g09533(.A1(new_n12113_), .A2(new_n12133_), .ZN(new_n12432_));
  INV_X1     g09534(.I(new_n12432_), .ZN(new_n12433_));
  AOI21_X1   g09535(.A1(new_n12433_), .A2(new_n2614_), .B(pi0223), .ZN(new_n12434_));
  INV_X1     g09536(.I(new_n12434_), .ZN(new_n12435_));
  AOI21_X1   g09537(.A1(new_n12423_), .A2(new_n12431_), .B(new_n12435_), .ZN(new_n12436_));
  NOR2_X1    g09538(.A1(new_n12396_), .A2(new_n12436_), .ZN(new_n12437_));
  INV_X1     g09539(.I(new_n12363_), .ZN(new_n12438_));
  NOR3_X1    g09540(.A1(new_n12438_), .A2(new_n6445_), .A3(new_n12391_), .ZN(new_n12439_));
  AOI21_X1   g09541(.A1(new_n5094_), .A2(new_n12391_), .B(new_n12363_), .ZN(new_n12440_));
  OAI21_X1   g09542(.A1(new_n12439_), .A2(new_n12440_), .B(pi0215), .ZN(new_n12441_));
  AOI21_X1   g09543(.A1(new_n12432_), .A2(new_n3285_), .B(pi0215), .ZN(new_n12442_));
  INV_X1     g09544(.I(pi0614), .ZN(new_n12443_));
  INV_X1     g09545(.I(new_n12399_), .ZN(new_n12444_));
  INV_X1     g09546(.I(new_n12402_), .ZN(new_n12445_));
  OAI22_X1   g09547(.A1(new_n12445_), .A2(new_n12400_), .B1(new_n12384_), .B2(new_n12132_), .ZN(new_n12446_));
  NAND2_X1   g09548(.A1(new_n12446_), .A2(new_n12444_), .ZN(new_n12447_));
  AOI21_X1   g09549(.A1(new_n12447_), .A2(new_n12112_), .B(new_n12443_), .ZN(new_n12448_));
  NOR4_X1    g09550(.A1(new_n12448_), .A2(pi0616), .A3(new_n12379_), .A4(new_n12388_), .ZN(new_n12449_));
  NAND4_X1   g09551(.A1(new_n12409_), .A2(new_n5102_), .A3(new_n12133_), .A4(new_n12408_), .ZN(new_n12450_));
  OAI22_X1   g09552(.A1(new_n12230_), .A2(new_n12229_), .B1(new_n5103_), .B2(new_n12133_), .ZN(new_n12451_));
  NAND2_X1   g09553(.A1(new_n12450_), .A2(new_n12451_), .ZN(new_n12452_));
  MUX2_X1    g09554(.I0(new_n12452_), .I1(new_n12133_), .S(new_n5104_), .Z(new_n12453_));
  AOI21_X1   g09555(.A1(new_n12453_), .A2(new_n5095_), .B(new_n12420_), .ZN(new_n12454_));
  OAI21_X1   g09556(.A1(new_n12449_), .A2(new_n12222_), .B(new_n12454_), .ZN(new_n12455_));
  AOI21_X1   g09557(.A1(new_n6445_), .A2(new_n12429_), .B(new_n12455_), .ZN(new_n12456_));
  NOR3_X1    g09558(.A1(new_n12423_), .A2(new_n5094_), .A3(new_n12429_), .ZN(new_n12457_));
  NOR3_X1    g09559(.A1(new_n12456_), .A2(new_n12457_), .A3(new_n3284_), .ZN(new_n12458_));
  OAI21_X1   g09560(.A1(new_n12458_), .A2(new_n12442_), .B(new_n12441_), .ZN(new_n12459_));
  MUX2_X1    g09561(.I0(new_n12459_), .I1(new_n12437_), .S(new_n2587_), .Z(new_n12460_));
  INV_X1     g09562(.I(new_n12129_), .ZN(new_n12461_));
  NAND2_X1   g09563(.A1(new_n12242_), .A2(new_n12113_), .ZN(new_n12462_));
  INV_X1     g09564(.I(new_n12219_), .ZN(new_n12463_));
  AOI21_X1   g09565(.A1(new_n12262_), .A2(new_n5108_), .B(new_n12247_), .ZN(new_n12464_));
  NAND3_X1   g09566(.A1(new_n12464_), .A2(new_n12463_), .A3(new_n12307_), .ZN(new_n12465_));
  NAND2_X1   g09567(.A1(new_n12465_), .A2(pi0616), .ZN(new_n12466_));
  NAND2_X1   g09568(.A1(new_n12294_), .A2(new_n12463_), .ZN(new_n12467_));
  NAND2_X1   g09569(.A1(new_n12467_), .A2(new_n12384_), .ZN(new_n12468_));
  NAND2_X1   g09570(.A1(new_n12465_), .A2(new_n12443_), .ZN(new_n12469_));
  OAI21_X1   g09571(.A1(new_n12468_), .A2(new_n12469_), .B(new_n12166_), .ZN(new_n12470_));
  NAND2_X1   g09572(.A1(new_n12470_), .A2(new_n12466_), .ZN(new_n12471_));
  AOI22_X1   g09573(.A1(new_n12471_), .A2(new_n12461_), .B1(new_n12222_), .B2(new_n12462_), .ZN(new_n12472_));
  OAI21_X1   g09574(.A1(new_n12262_), .A2(new_n5108_), .B(new_n12408_), .ZN(new_n12473_));
  NAND3_X1   g09575(.A1(new_n12294_), .A2(new_n12473_), .A3(new_n5100_), .ZN(new_n12474_));
  AOI21_X1   g09576(.A1(new_n12297_), .A2(new_n12289_), .B(new_n11883_), .ZN(new_n12475_));
  NOR2_X1    g09577(.A1(new_n12475_), .A2(pi0616), .ZN(new_n12476_));
  NOR2_X1    g09578(.A1(new_n12287_), .A2(new_n11883_), .ZN(new_n12477_));
  INV_X1     g09579(.I(new_n12477_), .ZN(new_n12478_));
  AOI21_X1   g09580(.A1(new_n12478_), .A2(pi0616), .B(new_n12222_), .ZN(new_n12479_));
  INV_X1     g09581(.I(new_n12479_), .ZN(new_n12480_));
  OAI22_X1   g09582(.A1(new_n12476_), .A2(new_n12480_), .B1(new_n12219_), .B2(new_n12474_), .ZN(new_n12481_));
  MUX2_X1    g09583(.I0(new_n12481_), .I1(new_n12472_), .S(new_n5094_), .Z(new_n12482_));
  NAND2_X1   g09584(.A1(new_n12482_), .A2(new_n2566_), .ZN(new_n12483_));
  NOR2_X1    g09585(.A1(new_n12169_), .A2(pi0603), .ZN(new_n12484_));
  INV_X1     g09586(.I(new_n12183_), .ZN(new_n12485_));
  NOR2_X1    g09587(.A1(new_n12485_), .A2(new_n5101_), .ZN(new_n12486_));
  NOR2_X1    g09588(.A1(new_n12484_), .A2(new_n12486_), .ZN(new_n12487_));
  NOR2_X1    g09589(.A1(new_n5109_), .A2(pi0603), .ZN(new_n12488_));
  AOI22_X1   g09590(.A1(new_n12158_), .A2(new_n5101_), .B1(new_n12213_), .B2(new_n12488_), .ZN(new_n12489_));
  NAND2_X1   g09591(.A1(new_n12489_), .A2(new_n12162_), .ZN(new_n12490_));
  MUX2_X1    g09592(.I0(new_n12487_), .I1(new_n12490_), .S(new_n12187_), .Z(new_n12491_));
  NAND2_X1   g09593(.A1(new_n12485_), .A2(pi0603), .ZN(new_n12492_));
  OAI21_X1   g09594(.A1(new_n12492_), .A2(new_n12200_), .B(new_n12222_), .ZN(new_n12493_));
  AOI21_X1   g09595(.A1(new_n12491_), .A2(new_n12461_), .B(new_n12493_), .ZN(new_n12494_));
  NAND2_X1   g09596(.A1(new_n12409_), .A2(new_n12408_), .ZN(new_n12495_));
  NAND3_X1   g09597(.A1(new_n12220_), .A2(pi0616), .A3(new_n12167_), .ZN(new_n12496_));
  AOI22_X1   g09598(.A1(new_n12420_), .A2(new_n12495_), .B1(new_n12479_), .B2(new_n12496_), .ZN(new_n12497_));
  NOR3_X1    g09599(.A1(new_n5094_), .A2(new_n2566_), .A3(new_n3284_), .ZN(new_n12498_));
  OAI21_X1   g09600(.A1(new_n12497_), .A2(new_n6445_), .B(new_n12498_), .ZN(new_n12499_));
  OR2_X2     g09601(.A1(new_n12494_), .A2(new_n12499_), .Z(new_n12500_));
  AOI21_X1   g09602(.A1(new_n12500_), .A2(new_n12483_), .B(new_n2587_), .ZN(new_n12501_));
  NAND2_X1   g09603(.A1(new_n12497_), .A2(new_n5141_), .ZN(new_n12502_));
  NAND2_X1   g09604(.A1(new_n12502_), .A2(new_n3155_), .ZN(new_n12503_));
  NOR2_X1    g09605(.A1(new_n12133_), .A2(new_n3155_), .ZN(new_n12504_));
  INV_X1     g09606(.I(new_n12504_), .ZN(new_n12505_));
  NOR2_X1    g09607(.A1(new_n12505_), .A2(new_n11875_), .ZN(new_n12506_));
  NOR2_X1    g09608(.A1(new_n12506_), .A2(pi0223), .ZN(new_n12507_));
  INV_X1     g09609(.I(new_n12507_), .ZN(new_n12508_));
  NAND2_X1   g09610(.A1(new_n12269_), .A2(new_n12508_), .ZN(new_n12509_));
  NAND4_X1   g09611(.A1(new_n12494_), .A2(new_n6460_), .A3(new_n12503_), .A4(new_n12509_), .ZN(new_n12510_));
  INV_X1     g09612(.I(new_n12481_), .ZN(new_n12511_));
  MUX2_X1    g09613(.I0(new_n12511_), .I1(new_n12472_), .S(new_n6460_), .Z(new_n12512_));
  NAND2_X1   g09614(.A1(new_n12512_), .A2(pi0223), .ZN(new_n12513_));
  AOI21_X1   g09615(.A1(new_n12510_), .A2(new_n12513_), .B(pi0299), .ZN(new_n12514_));
  NOR2_X1    g09616(.A1(new_n12501_), .A2(new_n12514_), .ZN(new_n12515_));
  OAI21_X1   g09617(.A1(new_n12515_), .A2(new_n7339_), .B(pi0761), .ZN(new_n12516_));
  AOI21_X1   g09618(.A1(new_n12460_), .A2(new_n7339_), .B(new_n12516_), .ZN(new_n12517_));
  OAI21_X1   g09619(.A1(new_n12517_), .A2(new_n12350_), .B(pi0039), .ZN(new_n12518_));
  OAI21_X1   g09620(.A1(new_n2459_), .A2(pi0102), .B(new_n8394_), .ZN(new_n12519_));
  OAI21_X1   g09621(.A1(pi0102), .A2(new_n8572_), .B(new_n12519_), .ZN(new_n12520_));
  NAND2_X1   g09622(.A1(new_n12520_), .A2(new_n2710_), .ZN(new_n12521_));
  NOR2_X1    g09623(.A1(new_n8395_), .A2(new_n7843_), .ZN(new_n12522_));
  OR3_X2     g09624(.A1(new_n2681_), .A2(new_n5276_), .A3(new_n7903_), .Z(new_n12523_));
  OAI21_X1   g09625(.A1(new_n2664_), .A2(pi0091), .B(new_n2666_), .ZN(new_n12524_));
  NAND3_X1   g09626(.A1(new_n12523_), .A2(new_n12524_), .A3(new_n2661_), .ZN(new_n12525_));
  AOI21_X1   g09627(.A1(new_n12521_), .A2(new_n12522_), .B(new_n12525_), .ZN(new_n12526_));
  NOR3_X1    g09628(.A1(new_n8395_), .A2(pi0252), .A3(new_n7430_), .ZN(new_n12527_));
  NAND2_X1   g09629(.A1(new_n12521_), .A2(new_n12527_), .ZN(new_n12528_));
  NOR2_X1    g09630(.A1(new_n5240_), .A2(pi0035), .ZN(new_n12529_));
  NOR4_X1    g09631(.A1(new_n12529_), .A2(new_n3181_), .A3(new_n2507_), .A4(new_n2907_), .ZN(new_n12530_));
  NAND2_X1   g09632(.A1(new_n12530_), .A2(new_n12528_), .ZN(new_n12531_));
  NOR2_X1    g09633(.A1(new_n3365_), .A2(pi0032), .ZN(new_n12532_));
  OAI21_X1   g09634(.A1(new_n12531_), .A2(new_n12526_), .B(new_n12532_), .ZN(new_n12533_));
  NAND3_X1   g09635(.A1(new_n5241_), .A2(new_n2484_), .A3(new_n2955_), .ZN(new_n12534_));
  NOR2_X1    g09636(.A1(new_n12534_), .A2(new_n5366_), .ZN(new_n12535_));
  NOR2_X1    g09637(.A1(new_n7904_), .A2(new_n5276_), .ZN(new_n12536_));
  NOR2_X1    g09638(.A1(new_n8572_), .A2(pi0102), .ZN(new_n12537_));
  AOI21_X1   g09639(.A1(new_n5268_), .A2(new_n2462_), .B(pi0098), .ZN(new_n12538_));
  NOR3_X1    g09640(.A1(new_n6989_), .A2(new_n5956_), .A3(pi0088), .ZN(new_n12539_));
  INV_X1     g09641(.I(new_n12539_), .ZN(new_n12540_));
  NOR4_X1    g09642(.A1(new_n12538_), .A2(new_n12537_), .A3(new_n6987_), .A4(new_n12540_), .ZN(new_n12541_));
  NOR4_X1    g09643(.A1(new_n12536_), .A2(new_n12541_), .A3(new_n12524_), .A4(pi0047), .ZN(new_n12542_));
  NOR2_X1    g09644(.A1(new_n2506_), .A2(pi0040), .ZN(new_n12543_));
  NAND4_X1   g09645(.A1(new_n12542_), .A2(new_n2876_), .A3(new_n5970_), .A4(new_n12543_), .ZN(new_n12544_));
  NOR4_X1    g09646(.A1(new_n12520_), .A2(new_n7014_), .A3(new_n7250_), .A4(new_n12540_), .ZN(new_n12545_));
  NOR2_X1    g09647(.A1(new_n7194_), .A2(pi0040), .ZN(new_n12546_));
  INV_X1     g09648(.I(new_n12546_), .ZN(new_n12547_));
  OAI21_X1   g09649(.A1(new_n12545_), .A2(new_n12547_), .B(new_n3181_), .ZN(new_n12548_));
  INV_X1     g09650(.I(new_n12548_), .ZN(new_n12549_));
  NAND2_X1   g09651(.A1(new_n2858_), .A2(pi0252), .ZN(new_n12550_));
  INV_X1     g09652(.I(new_n12550_), .ZN(new_n12551_));
  NOR4_X1    g09653(.A1(new_n12549_), .A2(new_n12544_), .A3(new_n2484_), .A4(new_n12551_), .ZN(new_n12552_));
  NOR2_X1    g09654(.A1(new_n9157_), .A2(new_n2923_), .ZN(new_n12553_));
  AOI22_X1   g09655(.A1(new_n12552_), .A2(new_n12553_), .B1(new_n12533_), .B2(new_n12535_), .ZN(new_n12554_));
  NOR2_X1    g09656(.A1(new_n12554_), .A2(new_n9141_), .ZN(new_n12555_));
  INV_X1     g09657(.I(new_n12555_), .ZN(new_n12556_));
  NOR2_X1    g09658(.A1(new_n9859_), .A2(new_n2923_), .ZN(po1106));
  AOI21_X1   g09659(.A1(new_n12552_), .A2(po1106), .B(new_n2921_), .ZN(new_n12558_));
  INV_X1     g09660(.I(new_n12558_), .ZN(new_n12559_));
  AOI21_X1   g09661(.A1(new_n12544_), .A2(new_n12551_), .B(new_n12549_), .ZN(new_n12560_));
  NOR3_X1    g09662(.A1(new_n12534_), .A2(pi0824), .A3(new_n2927_), .ZN(new_n12561_));
  OAI21_X1   g09663(.A1(new_n12560_), .A2(pi0032), .B(new_n12561_), .ZN(new_n12562_));
  AOI21_X1   g09664(.A1(new_n12554_), .A2(new_n12562_), .B(new_n2924_), .ZN(new_n12563_));
  OAI21_X1   g09665(.A1(new_n12563_), .A2(new_n2920_), .B(new_n12559_), .ZN(new_n12564_));
  NAND2_X1   g09666(.A1(new_n12564_), .A2(new_n12556_), .ZN(new_n12565_));
  INV_X1     g09667(.I(new_n12524_), .ZN(new_n12566_));
  NOR3_X1    g09668(.A1(new_n12537_), .A2(new_n6987_), .A3(new_n12540_), .ZN(new_n12567_));
  NAND2_X1   g09669(.A1(new_n12567_), .A2(new_n12519_), .ZN(new_n12568_));
  NAND4_X1   g09670(.A1(new_n12568_), .A2(new_n12566_), .A3(new_n2661_), .A4(new_n12523_), .ZN(new_n12569_));
  NAND2_X1   g09671(.A1(new_n12529_), .A2(new_n12543_), .ZN(new_n12570_));
  AOI21_X1   g09672(.A1(new_n12569_), .A2(new_n2876_), .B(new_n12570_), .ZN(new_n12571_));
  NOR4_X1    g09673(.A1(new_n2511_), .A2(new_n3364_), .A3(new_n3181_), .A4(new_n2484_), .ZN(new_n12572_));
  NAND3_X1   g09674(.A1(new_n12571_), .A2(new_n12572_), .A3(new_n12553_), .ZN(new_n12573_));
  NAND2_X1   g09675(.A1(new_n12521_), .A2(new_n12522_), .ZN(new_n12574_));
  NAND4_X1   g09676(.A1(new_n12574_), .A2(new_n2661_), .A3(new_n12523_), .A4(new_n12524_), .ZN(new_n12575_));
  NAND2_X1   g09677(.A1(new_n7918_), .A2(new_n6004_), .ZN(new_n12576_));
  NAND4_X1   g09678(.A1(new_n12575_), .A2(new_n12528_), .A3(new_n12530_), .A4(new_n12576_), .ZN(new_n12577_));
  AOI21_X1   g09679(.A1(new_n12573_), .A2(new_n12577_), .B(new_n2924_), .ZN(new_n12578_));
  NOR2_X1    g09680(.A1(new_n12578_), .A2(new_n2920_), .ZN(new_n12579_));
  NOR2_X1    g09681(.A1(new_n12579_), .A2(new_n12558_), .ZN(new_n12580_));
  NAND2_X1   g09682(.A1(new_n12578_), .A2(new_n2918_), .ZN(new_n12581_));
  INV_X1     g09683(.I(new_n12581_), .ZN(new_n12582_));
  OAI21_X1   g09684(.A1(new_n12580_), .A2(new_n12582_), .B(new_n2601_), .ZN(new_n12583_));
  OAI21_X1   g09685(.A1(new_n12565_), .A2(new_n2601_), .B(new_n12583_), .ZN(new_n12584_));
  OAI21_X1   g09686(.A1(new_n2920_), .A2(new_n12578_), .B(new_n12559_), .ZN(new_n12585_));
  MUX2_X1    g09687(.I0(new_n12585_), .I1(new_n12564_), .S(pi0198), .Z(new_n12586_));
  NOR2_X1    g09688(.A1(new_n12586_), .A2(new_n11882_), .ZN(new_n12587_));
  NOR3_X1    g09689(.A1(new_n12587_), .A2(new_n5095_), .A3(new_n12584_), .ZN(new_n12588_));
  OAI21_X1   g09690(.A1(new_n12580_), .A2(new_n12582_), .B(new_n2631_), .ZN(new_n12589_));
  OAI21_X1   g09691(.A1(new_n12565_), .A2(new_n2631_), .B(new_n12589_), .ZN(new_n12590_));
  NAND2_X1   g09692(.A1(new_n12533_), .A2(new_n12535_), .ZN(new_n12591_));
  NAND2_X1   g09693(.A1(new_n12591_), .A2(new_n12573_), .ZN(new_n12592_));
  OAI21_X1   g09694(.A1(new_n12571_), .A2(new_n12550_), .B(new_n12548_), .ZN(new_n12593_));
  INV_X1     g09695(.I(new_n12561_), .ZN(new_n12594_));
  AOI21_X1   g09696(.A1(new_n12593_), .A2(new_n2632_), .B(new_n12594_), .ZN(new_n12595_));
  OAI21_X1   g09697(.A1(new_n12592_), .A2(new_n12595_), .B(pi1093), .ZN(new_n12596_));
  AOI21_X1   g09698(.A1(new_n12596_), .A2(new_n2958_), .B(new_n12558_), .ZN(new_n12597_));
  NAND3_X1   g09699(.A1(new_n12597_), .A2(pi0210), .A3(new_n12585_), .ZN(new_n12598_));
  OAI21_X1   g09700(.A1(new_n12597_), .A2(new_n2631_), .B(new_n12580_), .ZN(new_n12599_));
  AOI21_X1   g09701(.A1(new_n12599_), .A2(new_n12598_), .B(new_n11882_), .ZN(new_n12600_));
  NOR4_X1    g09702(.A1(new_n12600_), .A2(pi0299), .A3(new_n12590_), .A4(new_n5095_), .ZN(new_n12601_));
  NOR3_X1    g09703(.A1(new_n12588_), .A2(new_n12601_), .A3(pi0299), .ZN(new_n12602_));
  NOR3_X1    g09704(.A1(new_n12579_), .A2(pi0621), .A3(new_n12558_), .ZN(new_n12603_));
  OR3_X2     g09705(.A1(new_n12603_), .A2(pi0198), .A3(new_n12582_), .Z(new_n12604_));
  NOR3_X1    g09706(.A1(new_n12597_), .A2(pi0621), .A3(new_n12555_), .ZN(new_n12605_));
  NOR3_X1    g09707(.A1(new_n12604_), .A2(new_n12605_), .A3(new_n2601_), .ZN(new_n12606_));
  NOR3_X1    g09708(.A1(new_n12603_), .A2(pi0198), .A3(new_n12582_), .ZN(new_n12607_));
  NAND3_X1   g09709(.A1(new_n12564_), .A2(new_n11872_), .A3(new_n12556_), .ZN(new_n12608_));
  AOI21_X1   g09710(.A1(new_n12608_), .A2(pi0198), .B(new_n12607_), .ZN(new_n12609_));
  NOR3_X1    g09711(.A1(new_n12606_), .A2(new_n5101_), .A3(new_n12609_), .ZN(new_n12610_));
  NAND2_X1   g09712(.A1(new_n12610_), .A2(new_n2587_), .ZN(new_n12611_));
  OAI21_X1   g09713(.A1(new_n12603_), .A2(new_n12582_), .B(new_n2631_), .ZN(new_n12612_));
  OAI21_X1   g09714(.A1(new_n12608_), .A2(new_n2631_), .B(new_n12612_), .ZN(new_n12613_));
  NAND3_X1   g09715(.A1(new_n12613_), .A2(pi0299), .A3(pi0603), .ZN(new_n12614_));
  AOI21_X1   g09716(.A1(new_n12611_), .A2(new_n12614_), .B(new_n5095_), .ZN(new_n12615_));
  NOR2_X1    g09717(.A1(new_n12615_), .A2(new_n12602_), .ZN(new_n12616_));
  OAI21_X1   g09718(.A1(new_n12585_), .A2(new_n11872_), .B(new_n2601_), .ZN(new_n12617_));
  NAND3_X1   g09719(.A1(new_n12597_), .A2(new_n2601_), .A3(pi0621), .ZN(new_n12618_));
  NAND2_X1   g09720(.A1(new_n12618_), .A2(new_n12617_), .ZN(new_n12619_));
  NAND2_X1   g09721(.A1(new_n12619_), .A2(new_n11882_), .ZN(new_n12620_));
  AOI21_X1   g09722(.A1(new_n12580_), .A2(new_n11882_), .B(new_n12582_), .ZN(new_n12621_));
  NOR2_X1    g09723(.A1(new_n12621_), .A2(pi0198), .ZN(new_n12622_));
  OAI21_X1   g09724(.A1(new_n12564_), .A2(pi0665), .B(new_n12556_), .ZN(new_n12623_));
  AOI21_X1   g09725(.A1(pi0198), .A2(new_n12623_), .B(new_n12622_), .ZN(new_n12624_));
  MUX2_X1    g09726(.I0(new_n12624_), .I1(new_n12620_), .S(pi0603), .Z(new_n12625_));
  NOR3_X1    g09727(.A1(new_n12625_), .A2(pi0299), .A3(new_n5095_), .ZN(new_n12626_));
  AOI21_X1   g09728(.A1(new_n12599_), .A2(new_n12598_), .B(new_n11872_), .ZN(new_n12627_));
  NAND2_X1   g09729(.A1(new_n12627_), .A2(new_n11882_), .ZN(new_n12628_));
  NOR2_X1    g09730(.A1(new_n12621_), .A2(pi0210), .ZN(new_n12629_));
  AOI21_X1   g09731(.A1(pi0210), .A2(new_n12623_), .B(new_n12629_), .ZN(new_n12630_));
  MUX2_X1    g09732(.I0(new_n12630_), .I1(new_n12628_), .S(pi0603), .Z(new_n12631_));
  NOR3_X1    g09733(.A1(new_n12631_), .A2(new_n2587_), .A3(new_n5095_), .ZN(new_n12632_));
  NOR2_X1    g09734(.A1(new_n12632_), .A2(new_n12626_), .ZN(new_n12633_));
  AOI21_X1   g09735(.A1(new_n12633_), .A2(new_n12616_), .B(new_n7339_), .ZN(new_n12634_));
  NAND2_X1   g09736(.A1(new_n12634_), .A2(pi0761), .ZN(new_n12635_));
  INV_X1     g09737(.I(new_n12614_), .ZN(new_n12636_));
  AOI21_X1   g09738(.A1(new_n12610_), .A2(new_n2587_), .B(new_n12636_), .ZN(new_n12637_));
  INV_X1     g09739(.I(new_n12621_), .ZN(new_n12638_));
  NAND2_X1   g09740(.A1(new_n12638_), .A2(new_n2631_), .ZN(new_n12639_));
  NAND2_X1   g09741(.A1(new_n12623_), .A2(pi0210), .ZN(new_n12640_));
  NAND2_X1   g09742(.A1(new_n12639_), .A2(new_n12640_), .ZN(new_n12641_));
  OAI21_X1   g09743(.A1(new_n12641_), .A2(new_n12624_), .B(pi0299), .ZN(new_n12642_));
  NOR2_X1    g09744(.A1(new_n12642_), .A2(new_n5095_), .ZN(new_n12643_));
  INV_X1     g09745(.I(new_n12643_), .ZN(new_n12644_));
  NAND2_X1   g09746(.A1(new_n12644_), .A2(new_n12637_), .ZN(new_n12645_));
  INV_X1     g09747(.I(new_n12584_), .ZN(new_n12646_));
  MUX2_X1    g09748(.I0(new_n12580_), .I1(new_n12597_), .S(pi0198), .Z(new_n12647_));
  NAND2_X1   g09749(.A1(new_n12647_), .A2(pi0665), .ZN(new_n12648_));
  NAND3_X1   g09750(.A1(new_n12646_), .A2(new_n12648_), .A3(pi0680), .ZN(new_n12649_));
  NOR3_X1    g09751(.A1(new_n12597_), .A2(new_n2631_), .A3(new_n12555_), .ZN(new_n12650_));
  INV_X1     g09752(.I(new_n12589_), .ZN(new_n12651_));
  NOR2_X1    g09753(.A1(new_n12651_), .A2(new_n12650_), .ZN(new_n12652_));
  NOR3_X1    g09754(.A1(new_n12564_), .A2(new_n2631_), .A3(new_n12580_), .ZN(new_n12653_));
  AOI21_X1   g09755(.A1(new_n12564_), .A2(pi0210), .B(new_n12585_), .ZN(new_n12654_));
  OAI21_X1   g09756(.A1(new_n12653_), .A2(new_n12654_), .B(pi0665), .ZN(new_n12655_));
  NAND4_X1   g09757(.A1(new_n12655_), .A2(new_n12652_), .A3(new_n2587_), .A4(pi0680), .ZN(new_n12656_));
  NAND3_X1   g09758(.A1(new_n12649_), .A2(new_n12656_), .A3(new_n2587_), .ZN(new_n12657_));
  OAI21_X1   g09759(.A1(new_n12653_), .A2(new_n12654_), .B(pi0621), .ZN(new_n12658_));
  NAND4_X1   g09760(.A1(new_n12658_), .A2(new_n12652_), .A3(new_n2587_), .A4(pi0603), .ZN(new_n12659_));
  NAND3_X1   g09761(.A1(new_n12608_), .A2(new_n12607_), .A3(pi0198), .ZN(new_n12660_));
  OAI21_X1   g09762(.A1(new_n2601_), .A2(new_n12605_), .B(new_n12604_), .ZN(new_n12661_));
  NAND3_X1   g09763(.A1(new_n12618_), .A2(new_n12617_), .A3(new_n2587_), .ZN(new_n12662_));
  NAND4_X1   g09764(.A1(new_n12661_), .A2(new_n5101_), .A3(new_n12660_), .A4(new_n12662_), .ZN(new_n12663_));
  NAND2_X1   g09765(.A1(new_n12663_), .A2(new_n12659_), .ZN(new_n12664_));
  NOR2_X1    g09766(.A1(new_n12657_), .A2(new_n12664_), .ZN(new_n12665_));
  AOI21_X1   g09767(.A1(new_n7339_), .A2(new_n12665_), .B(new_n12645_), .ZN(new_n12666_));
  NAND2_X1   g09768(.A1(new_n12611_), .A2(new_n12614_), .ZN(new_n12667_));
  NOR2_X1    g09769(.A1(new_n12667_), .A2(new_n12643_), .ZN(new_n12668_));
  NOR3_X1    g09770(.A1(new_n12668_), .A2(pi0140), .A3(new_n12665_), .ZN(new_n12669_));
  NOR4_X1    g09771(.A1(new_n12666_), .A2(pi0039), .A3(pi0761), .A4(new_n12669_), .ZN(new_n12670_));
  AOI21_X1   g09772(.A1(new_n12670_), .A2(new_n12635_), .B(pi0038), .ZN(new_n12671_));
  AOI22_X1   g09773(.A1(new_n12518_), .A2(new_n12671_), .B1(pi0038), .B2(new_n12126_), .ZN(new_n12672_));
  NAND2_X1   g09774(.A1(new_n5217_), .A2(new_n12168_), .ZN(new_n12673_));
  MUX2_X1    g09775(.I0(new_n12206_), .I1(new_n12209_), .S(new_n12673_), .Z(new_n12674_));
  OAI21_X1   g09776(.A1(new_n12198_), .A2(new_n11875_), .B(new_n6445_), .ZN(new_n12675_));
  NOR2_X1    g09777(.A1(new_n12464_), .A2(new_n5094_), .ZN(new_n12676_));
  INV_X1     g09778(.I(new_n12676_), .ZN(new_n12677_));
  NAND2_X1   g09779(.A1(new_n12253_), .A2(new_n12677_), .ZN(new_n12678_));
  NAND2_X1   g09780(.A1(new_n12678_), .A2(pi0215), .ZN(new_n12679_));
  OAI21_X1   g09781(.A1(pi0120), .A2(new_n12131_), .B(new_n2490_), .ZN(new_n12680_));
  INV_X1     g09782(.I(new_n12680_), .ZN(new_n12681_));
  NAND3_X1   g09783(.A1(new_n12681_), .A2(new_n3284_), .A3(new_n11876_), .ZN(new_n12682_));
  NAND4_X1   g09784(.A1(new_n12679_), .A2(new_n4905_), .A3(new_n5094_), .A4(new_n12682_), .ZN(new_n12683_));
  AOI21_X1   g09785(.A1(new_n12675_), .A2(new_n3285_), .B(new_n12683_), .ZN(new_n12684_));
  NOR2_X1    g09786(.A1(new_n12464_), .A2(new_n5141_), .ZN(new_n12685_));
  INV_X1     g09787(.I(new_n12685_), .ZN(new_n12686_));
  NAND2_X1   g09788(.A1(new_n12253_), .A2(new_n12686_), .ZN(new_n12687_));
  AOI21_X1   g09789(.A1(new_n12687_), .A2(pi0223), .B(pi0299), .ZN(new_n12688_));
  INV_X1     g09790(.I(new_n12688_), .ZN(new_n12689_));
  NOR2_X1    g09791(.A1(new_n6460_), .A2(new_n3155_), .ZN(new_n12690_));
  NAND2_X1   g09792(.A1(new_n12674_), .A2(new_n12690_), .ZN(new_n12691_));
  NAND2_X1   g09793(.A1(new_n12691_), .A2(new_n12507_), .ZN(new_n12692_));
  AOI22_X1   g09794(.A1(new_n12684_), .A2(new_n12674_), .B1(new_n12692_), .B2(new_n12689_), .ZN(new_n12693_));
  MUX2_X1    g09795(.I0(new_n12693_), .I1(new_n12637_), .S(new_n3154_), .Z(new_n12694_));
  NOR3_X1    g09796(.A1(new_n12694_), .A2(new_n7339_), .A3(pi0761), .ZN(new_n12695_));
  NOR2_X1    g09797(.A1(new_n12652_), .A2(new_n2587_), .ZN(new_n12696_));
  AOI21_X1   g09798(.A1(new_n2587_), .A2(new_n12584_), .B(new_n12696_), .ZN(new_n12697_));
  NOR2_X1    g09799(.A1(new_n5096_), .A2(new_n5108_), .ZN(new_n12698_));
  NOR2_X1    g09800(.A1(new_n12242_), .A2(new_n12698_), .ZN(new_n12699_));
  NAND4_X1   g09801(.A1(new_n12367_), .A2(new_n12371_), .A3(new_n12698_), .A4(new_n12699_), .ZN(new_n12700_));
  INV_X1     g09802(.I(new_n12698_), .ZN(new_n12701_));
  INV_X1     g09803(.I(new_n12699_), .ZN(new_n12702_));
  OAI21_X1   g09804(.A1(new_n12372_), .A2(new_n12701_), .B(new_n12702_), .ZN(new_n12703_));
  NOR3_X1    g09805(.A1(new_n12361_), .A2(new_n12127_), .A3(new_n12249_), .ZN(new_n12704_));
  NAND4_X1   g09806(.A1(new_n12703_), .A2(new_n12127_), .A3(new_n12700_), .A4(new_n12704_), .ZN(new_n12705_));
  MUX2_X1    g09807(.I0(new_n12372_), .I1(new_n12242_), .S(new_n12701_), .Z(new_n12706_));
  INV_X1     g09808(.I(new_n12704_), .ZN(new_n12707_));
  OAI21_X1   g09809(.A1(new_n12706_), .A2(new_n12128_), .B(new_n12707_), .ZN(new_n12708_));
  AOI21_X1   g09810(.A1(new_n12708_), .A2(new_n12705_), .B(new_n5092_), .ZN(new_n12709_));
  NAND3_X1   g09811(.A1(new_n12708_), .A2(new_n5090_), .A3(new_n12705_), .ZN(new_n12710_));
  NOR2_X1    g09812(.A1(new_n12133_), .A2(new_n12129_), .ZN(new_n12711_));
  INV_X1     g09813(.I(new_n12711_), .ZN(new_n12712_));
  NOR2_X1    g09814(.A1(new_n12132_), .A2(pi0680), .ZN(new_n12713_));
  NOR3_X1    g09815(.A1(new_n12461_), .A2(new_n12166_), .A3(new_n12713_), .ZN(new_n12714_));
  INV_X1     g09816(.I(new_n12714_), .ZN(new_n12715_));
  NOR2_X1    g09817(.A1(new_n12473_), .A2(new_n5095_), .ZN(new_n12716_));
  OAI22_X1   g09818(.A1(new_n12716_), .A2(new_n12715_), .B1(new_n12166_), .B2(new_n12712_), .ZN(new_n12717_));
  NOR2_X1    g09819(.A1(new_n12129_), .A2(pi0616), .ZN(new_n12718_));
  INV_X1     g09820(.I(new_n12366_), .ZN(new_n12719_));
  NOR3_X1    g09821(.A1(new_n12719_), .A2(new_n12443_), .A3(new_n12364_), .ZN(new_n12720_));
  NOR2_X1    g09822(.A1(new_n12133_), .A2(new_n12443_), .ZN(new_n12721_));
  OAI21_X1   g09823(.A1(new_n12720_), .A2(new_n12721_), .B(new_n12718_), .ZN(new_n12722_));
  NOR2_X1    g09824(.A1(new_n12721_), .A2(pi0616), .ZN(new_n12723_));
  INV_X1     g09825(.I(new_n12723_), .ZN(new_n12724_));
  AOI21_X1   g09826(.A1(new_n12242_), .A2(new_n5109_), .B(new_n12229_), .ZN(new_n12725_));
  AOI21_X1   g09827(.A1(new_n12129_), .A2(new_n12166_), .B(pi0680), .ZN(new_n12726_));
  OAI21_X1   g09828(.A1(new_n12720_), .A2(new_n12724_), .B(new_n12726_), .ZN(new_n12727_));
  AOI21_X1   g09829(.A1(new_n12722_), .A2(new_n12727_), .B(new_n12717_), .ZN(new_n12728_));
  NAND2_X1   g09830(.A1(new_n12372_), .A2(pi0681), .ZN(new_n12729_));
  NOR3_X1    g09831(.A1(new_n12728_), .A2(pi0681), .A3(new_n12729_), .ZN(new_n12730_));
  INV_X1     g09832(.I(pi0681), .ZN(new_n12731_));
  NAND2_X1   g09833(.A1(new_n12725_), .A2(pi0680), .ZN(new_n12732_));
  AOI22_X1   g09834(.A1(new_n12732_), .A2(new_n12714_), .B1(pi0616), .B2(new_n12711_), .ZN(new_n12733_));
  INV_X1     g09835(.I(new_n12718_), .ZN(new_n12734_));
  NAND3_X1   g09836(.A1(new_n12365_), .A2(pi0614), .A3(new_n12366_), .ZN(new_n12735_));
  INV_X1     g09837(.I(new_n12721_), .ZN(new_n12736_));
  AOI21_X1   g09838(.A1(new_n12735_), .A2(new_n12736_), .B(new_n12734_), .ZN(new_n12737_));
  INV_X1     g09839(.I(new_n12726_), .ZN(new_n12738_));
  AOI21_X1   g09840(.A1(new_n12735_), .A2(new_n12723_), .B(new_n12738_), .ZN(new_n12739_));
  OAI21_X1   g09841(.A1(new_n12737_), .A2(new_n12739_), .B(new_n12733_), .ZN(new_n12740_));
  MUX2_X1    g09842(.I0(new_n12360_), .I1(new_n12133_), .S(new_n5104_), .Z(new_n12741_));
  NOR2_X1    g09843(.A1(new_n12741_), .A2(new_n12731_), .ZN(new_n12742_));
  AOI21_X1   g09844(.A1(new_n12731_), .A2(new_n12740_), .B(new_n12742_), .ZN(new_n12743_));
  OAI21_X1   g09845(.A1(new_n12743_), .A2(new_n12730_), .B(new_n5090_), .ZN(new_n12744_));
  AOI21_X1   g09846(.A1(new_n12710_), .A2(new_n12744_), .B(new_n5093_), .ZN(new_n12745_));
  NOR3_X1    g09847(.A1(new_n12745_), .A2(new_n2566_), .A3(new_n12709_), .ZN(new_n12746_));
  NAND3_X1   g09848(.A1(new_n12495_), .A2(new_n12443_), .A3(new_n5100_), .ZN(new_n12747_));
  NOR2_X1    g09849(.A1(new_n5100_), .A2(pi0614), .ZN(new_n12748_));
  OAI21_X1   g09850(.A1(pi0616), .A2(new_n12133_), .B(new_n12748_), .ZN(new_n12749_));
  NAND3_X1   g09851(.A1(new_n12450_), .A2(new_n12451_), .A3(new_n12166_), .ZN(new_n12750_));
  NAND2_X1   g09852(.A1(new_n12750_), .A2(new_n12749_), .ZN(new_n12751_));
  NOR2_X1    g09853(.A1(new_n12712_), .A2(new_n12443_), .ZN(new_n12752_));
  INV_X1     g09854(.I(new_n12752_), .ZN(new_n12753_));
  NOR3_X1    g09855(.A1(new_n12461_), .A2(new_n12443_), .A3(new_n12713_), .ZN(new_n12754_));
  INV_X1     g09856(.I(new_n12754_), .ZN(new_n12755_));
  NOR2_X1    g09857(.A1(new_n12495_), .A2(new_n5095_), .ZN(new_n12756_));
  OAI21_X1   g09858(.A1(new_n12756_), .A2(new_n12755_), .B(new_n12753_), .ZN(new_n12757_));
  AOI21_X1   g09859(.A1(new_n12751_), .A2(new_n12747_), .B(new_n12757_), .ZN(new_n12758_));
  MUX2_X1    g09860(.I0(new_n12758_), .I1(new_n12453_), .S(pi0681), .Z(new_n12759_));
  NOR4_X1    g09861(.A1(new_n12156_), .A2(new_n5098_), .A3(new_n12190_), .A4(new_n12133_), .ZN(new_n12760_));
  INV_X1     g09862(.I(new_n12760_), .ZN(new_n12761_));
  AOI21_X1   g09863(.A1(new_n5461_), .A2(new_n12132_), .B(new_n12156_), .ZN(new_n12762_));
  OAI22_X1   g09864(.A1(new_n12181_), .A2(new_n12144_), .B1(new_n12190_), .B2(new_n12132_), .ZN(new_n12763_));
  NAND2_X1   g09865(.A1(new_n12763_), .A2(new_n5099_), .ZN(new_n12764_));
  OAI21_X1   g09866(.A1(new_n12764_), .A2(new_n12762_), .B(new_n12156_), .ZN(new_n12765_));
  NAND3_X1   g09867(.A1(new_n12193_), .A2(new_n12195_), .A3(pi0681), .ZN(new_n12766_));
  NAND4_X1   g09868(.A1(new_n12765_), .A2(new_n12731_), .A3(new_n12766_), .A4(new_n12761_), .ZN(new_n12767_));
  AOI21_X1   g09869(.A1(new_n12767_), .A2(new_n5091_), .B(new_n5093_), .ZN(new_n12768_));
  NOR3_X1    g09870(.A1(new_n12768_), .A2(new_n3284_), .A3(new_n5090_), .ZN(new_n12769_));
  NOR2_X1    g09871(.A1(new_n12133_), .A2(new_n3285_), .ZN(new_n12770_));
  OAI21_X1   g09872(.A1(new_n12190_), .A2(new_n12133_), .B(new_n12191_), .ZN(new_n12771_));
  AOI22_X1   g09873(.A1(new_n12155_), .A2(new_n12145_), .B1(new_n5461_), .B2(new_n12133_), .ZN(new_n12772_));
  NOR2_X1    g09874(.A1(new_n12772_), .A2(new_n5098_), .ZN(new_n12773_));
  AOI21_X1   g09875(.A1(new_n12771_), .A2(new_n12773_), .B(new_n12191_), .ZN(new_n12774_));
  NOR3_X1    g09876(.A1(new_n12325_), .A2(new_n12324_), .A3(new_n12731_), .ZN(new_n12775_));
  NOR4_X1    g09877(.A1(new_n12774_), .A2(new_n12775_), .A3(pi0681), .A4(new_n12760_), .ZN(new_n12776_));
  AOI21_X1   g09878(.A1(new_n12776_), .A2(new_n5093_), .B(new_n3285_), .ZN(new_n12777_));
  NOR3_X1    g09879(.A1(new_n12777_), .A2(pi0215), .A3(new_n12770_), .ZN(new_n12778_));
  AOI21_X1   g09880(.A1(new_n12759_), .A2(new_n12769_), .B(new_n12778_), .ZN(new_n12779_));
  OAI21_X1   g09881(.A1(new_n12779_), .A2(new_n12746_), .B(pi0299), .ZN(new_n12780_));
  INV_X1     g09882(.I(new_n12705_), .ZN(new_n12781_));
  MUX2_X1    g09883(.I0(new_n12741_), .I1(new_n12262_), .S(new_n12701_), .Z(new_n12782_));
  AOI21_X1   g09884(.A1(new_n12782_), .A2(new_n12127_), .B(new_n12704_), .ZN(new_n12783_));
  NOR2_X1    g09885(.A1(new_n12783_), .A2(new_n12781_), .ZN(new_n12784_));
  NOR2_X1    g09886(.A1(new_n12784_), .A2(new_n5141_), .ZN(new_n12785_));
  NOR2_X1    g09887(.A1(new_n12743_), .A2(new_n12730_), .ZN(new_n12786_));
  NOR2_X1    g09888(.A1(new_n12786_), .A2(new_n6460_), .ZN(new_n12787_));
  NOR3_X1    g09889(.A1(new_n12785_), .A2(new_n2604_), .A3(new_n12787_), .ZN(new_n12788_));
  AOI21_X1   g09890(.A1(new_n12767_), .A2(new_n6460_), .B(new_n2614_), .ZN(new_n12789_));
  OAI21_X1   g09891(.A1(new_n12759_), .A2(new_n6460_), .B(new_n12789_), .ZN(new_n12790_));
  NOR2_X1    g09892(.A1(new_n12504_), .A2(pi0223), .ZN(new_n12791_));
  AOI21_X1   g09893(.A1(new_n12790_), .A2(new_n12791_), .B(new_n12788_), .ZN(new_n12792_));
  OAI21_X1   g09894(.A1(pi0299), .A2(new_n12792_), .B(new_n12780_), .ZN(new_n12793_));
  MUX2_X1    g09895(.I0(new_n12793_), .I1(new_n12697_), .S(new_n3154_), .Z(new_n12794_));
  NAND2_X1   g09896(.A1(new_n12299_), .A2(new_n12474_), .ZN(new_n12795_));
  NOR2_X1    g09897(.A1(new_n12312_), .A2(new_n5100_), .ZN(new_n12796_));
  NOR2_X1    g09898(.A1(new_n12262_), .A2(new_n12308_), .ZN(new_n12797_));
  AOI22_X1   g09899(.A1(new_n12796_), .A2(new_n12309_), .B1(new_n5100_), .B2(new_n12797_), .ZN(new_n12798_));
  INV_X1     g09900(.I(new_n12798_), .ZN(new_n12799_));
  OAI21_X1   g09901(.A1(new_n5094_), .A2(new_n12799_), .B(new_n12795_), .ZN(new_n12800_));
  INV_X1     g09902(.I(new_n12474_), .ZN(new_n12801_));
  AOI21_X1   g09903(.A1(new_n5217_), .A2(new_n12298_), .B(new_n12801_), .ZN(new_n12802_));
  NAND3_X1   g09904(.A1(new_n12802_), .A2(new_n6445_), .A3(new_n12799_), .ZN(new_n12803_));
  AOI21_X1   g09905(.A1(new_n12800_), .A2(new_n12803_), .B(new_n2566_), .ZN(new_n12804_));
  NAND3_X1   g09906(.A1(new_n12335_), .A2(new_n5217_), .A3(new_n12289_), .ZN(new_n12806_));
  NAND2_X1   g09907(.A1(new_n12806_), .A2(new_n5094_), .ZN(new_n12807_));
  INV_X1     g09908(.I(new_n12197_), .ZN(new_n12808_));
  OAI21_X1   g09909(.A1(new_n12326_), .A2(new_n5100_), .B(new_n12808_), .ZN(new_n12809_));
  INV_X1     g09910(.I(new_n12170_), .ZN(new_n12810_));
  NAND4_X1   g09911(.A1(new_n12158_), .A2(new_n5101_), .A3(new_n12810_), .A4(new_n12182_), .ZN(new_n12811_));
  NAND2_X1   g09912(.A1(new_n12809_), .A2(new_n12811_), .ZN(new_n12812_));
  AOI22_X1   g09913(.A1(new_n6445_), .A2(new_n12812_), .B1(new_n12807_), .B2(new_n3285_), .ZN(new_n12813_));
  OAI21_X1   g09914(.A1(new_n12287_), .A2(new_n3285_), .B(new_n2566_), .ZN(new_n12814_));
  OAI21_X1   g09915(.A1(new_n12813_), .A2(new_n12814_), .B(new_n2587_), .ZN(new_n12815_));
  NOR2_X1    g09916(.A1(new_n12815_), .A2(new_n12804_), .ZN(new_n12816_));
  MUX2_X1    g09917(.I0(new_n12798_), .I1(new_n12802_), .S(new_n5141_), .Z(new_n12817_));
  NAND2_X1   g09918(.A1(new_n12806_), .A2(new_n5141_), .ZN(new_n12818_));
  AOI22_X1   g09919(.A1(new_n6460_), .A2(new_n12812_), .B1(new_n12818_), .B2(new_n3155_), .ZN(new_n12819_));
  OAI21_X1   g09920(.A1(new_n12287_), .A2(new_n3155_), .B(new_n2604_), .ZN(new_n12820_));
  OAI22_X1   g09921(.A1(new_n12819_), .A2(new_n12820_), .B1(new_n2604_), .B2(new_n12817_), .ZN(new_n12821_));
  NAND2_X1   g09922(.A1(new_n12821_), .A2(new_n2587_), .ZN(new_n12822_));
  NOR2_X1    g09923(.A1(new_n12822_), .A2(new_n12816_), .ZN(new_n12823_));
  MUX2_X1    g09924(.I0(new_n12823_), .I1(new_n12664_), .S(new_n3154_), .Z(new_n12824_));
  NOR3_X1    g09925(.A1(new_n12794_), .A2(new_n7339_), .A3(new_n12116_), .ZN(new_n12825_));
  NOR2_X1    g09926(.A1(new_n12825_), .A2(new_n12695_), .ZN(new_n12826_));
  INV_X1     g09927(.I(new_n12826_), .ZN(new_n12827_));
  NOR2_X1    g09928(.A1(new_n5157_), .A2(new_n2926_), .ZN(new_n12828_));
  NOR2_X1    g09929(.A1(new_n5157_), .A2(new_n11877_), .ZN(new_n12829_));
  AOI21_X1   g09930(.A1(new_n12829_), .A2(new_n12116_), .B(new_n3172_), .ZN(new_n12830_));
  OAI21_X1   g09931(.A1(pi0140), .A2(new_n12828_), .B(new_n12830_), .ZN(new_n12831_));
  NAND3_X1   g09932(.A1(new_n12831_), .A2(pi0038), .A3(new_n11881_), .ZN(new_n12832_));
  OAI22_X1   g09933(.A1(new_n12672_), .A2(pi0738), .B1(new_n12827_), .B2(new_n12832_), .ZN(new_n12833_));
  MUX2_X1    g09934(.I0(new_n12833_), .I1(new_n7339_), .S(new_n3232_), .Z(new_n12834_));
  INV_X1     g09935(.I(new_n12834_), .ZN(new_n12835_));
  NOR2_X1    g09936(.A1(new_n3231_), .A2(pi0140), .ZN(new_n12836_));
  NAND3_X1   g09937(.A1(new_n12833_), .A2(new_n3231_), .A3(new_n12836_), .ZN(new_n12837_));
  INV_X1     g09938(.I(new_n12836_), .ZN(new_n12838_));
  NAND2_X1   g09939(.A1(new_n12126_), .A2(pi0038), .ZN(new_n12839_));
  NAND2_X1   g09940(.A1(new_n12518_), .A2(new_n12671_), .ZN(new_n12840_));
  NAND2_X1   g09941(.A1(new_n12840_), .A2(new_n12839_), .ZN(new_n12841_));
  NOR2_X1    g09942(.A1(new_n12827_), .A2(new_n12832_), .ZN(new_n12842_));
  AOI21_X1   g09943(.A1(new_n12841_), .A2(new_n11881_), .B(new_n12842_), .ZN(new_n12843_));
  OAI21_X1   g09944(.A1(new_n12843_), .A2(new_n3232_), .B(new_n12838_), .ZN(new_n12844_));
  NAND3_X1   g09945(.A1(new_n12844_), .A2(new_n12837_), .A3(pi0625), .ZN(new_n12845_));
  NOR2_X1    g09946(.A1(new_n12826_), .A2(pi0038), .ZN(new_n12846_));
  NAND2_X1   g09947(.A1(new_n12831_), .A2(new_n3231_), .ZN(new_n12847_));
  OAI21_X1   g09948(.A1(new_n12846_), .A2(new_n12847_), .B(new_n12838_), .ZN(new_n12848_));
  OAI21_X1   g09949(.A1(new_n12848_), .A2(pi0625), .B(new_n11893_), .ZN(new_n12849_));
  INV_X1     g09950(.I(new_n12849_), .ZN(new_n12850_));
  NAND2_X1   g09951(.A1(new_n12584_), .A2(new_n2587_), .ZN(new_n12851_));
  OAI21_X1   g09952(.A1(new_n2587_), .A2(new_n12652_), .B(new_n12851_), .ZN(new_n12852_));
  NOR2_X1    g09953(.A1(new_n12852_), .A2(pi0039), .ZN(new_n12853_));
  INV_X1     g09954(.I(new_n12853_), .ZN(new_n12854_));
  INV_X1     g09955(.I(new_n12709_), .ZN(new_n12855_));
  NOR3_X1    g09956(.A1(new_n12783_), .A2(new_n12781_), .A3(new_n5091_), .ZN(new_n12856_));
  NAND3_X1   g09957(.A1(new_n12740_), .A2(new_n12742_), .A3(new_n12731_), .ZN(new_n12857_));
  OAI21_X1   g09958(.A1(new_n12728_), .A2(pi0681), .B(new_n12729_), .ZN(new_n12858_));
  AOI21_X1   g09959(.A1(new_n12857_), .A2(new_n12858_), .B(new_n5091_), .ZN(new_n12859_));
  OAI21_X1   g09960(.A1(new_n12856_), .A2(new_n12859_), .B(new_n5092_), .ZN(new_n12860_));
  NAND3_X1   g09961(.A1(new_n12860_), .A2(pi0215), .A3(new_n12855_), .ZN(new_n12861_));
  NOR3_X1    g09962(.A1(new_n12231_), .A2(pi0614), .A3(new_n5217_), .ZN(new_n12862_));
  AOI21_X1   g09963(.A1(new_n12750_), .A2(new_n12749_), .B(new_n12862_), .ZN(new_n12863_));
  OAI21_X1   g09964(.A1(new_n12863_), .A2(new_n12757_), .B(new_n12731_), .ZN(new_n12864_));
  NOR4_X1    g09965(.A1(new_n12495_), .A2(new_n5102_), .A3(new_n5104_), .A4(new_n12132_), .ZN(new_n12865_));
  AOI21_X1   g09966(.A1(new_n12452_), .A2(new_n5105_), .B(new_n12133_), .ZN(new_n12866_));
  OAI21_X1   g09967(.A1(new_n12866_), .A2(new_n12865_), .B(pi0681), .ZN(new_n12867_));
  NOR2_X1    g09968(.A1(new_n12864_), .A2(new_n12867_), .ZN(new_n12868_));
  INV_X1     g09969(.I(new_n12749_), .ZN(new_n12869_));
  NOR3_X1    g09970(.A1(new_n12410_), .A2(new_n12407_), .A3(pi0616), .ZN(new_n12870_));
  OAI21_X1   g09971(.A1(new_n12870_), .A2(new_n12869_), .B(new_n12747_), .ZN(new_n12871_));
  NAND2_X1   g09972(.A1(new_n12231_), .A2(pi0680), .ZN(new_n12872_));
  AOI21_X1   g09973(.A1(new_n12872_), .A2(new_n12754_), .B(new_n12752_), .ZN(new_n12873_));
  AOI21_X1   g09974(.A1(new_n12871_), .A2(new_n12873_), .B(pi0681), .ZN(new_n12874_));
  INV_X1     g09975(.I(new_n12865_), .ZN(new_n12875_));
  OAI21_X1   g09976(.A1(new_n12411_), .A2(new_n5104_), .B(new_n12132_), .ZN(new_n12876_));
  AOI21_X1   g09977(.A1(new_n12876_), .A2(new_n12875_), .B(new_n12731_), .ZN(new_n12877_));
  NOR2_X1    g09978(.A1(new_n12874_), .A2(new_n12877_), .ZN(new_n12878_));
  NOR2_X1    g09979(.A1(new_n12878_), .A2(new_n12868_), .ZN(new_n12879_));
  INV_X1     g09980(.I(new_n12769_), .ZN(new_n12880_));
  INV_X1     g09981(.I(new_n12770_), .ZN(new_n12881_));
  OAI21_X1   g09982(.A1(new_n12767_), .A2(new_n5092_), .B(new_n3284_), .ZN(new_n12882_));
  NAND3_X1   g09983(.A1(new_n12882_), .A2(new_n2566_), .A3(new_n12881_), .ZN(new_n12883_));
  OAI21_X1   g09984(.A1(new_n12879_), .A2(new_n12880_), .B(new_n12883_), .ZN(new_n12884_));
  AOI21_X1   g09985(.A1(new_n12884_), .A2(new_n12861_), .B(new_n2587_), .ZN(new_n12885_));
  NAND2_X1   g09986(.A1(new_n12708_), .A2(new_n12705_), .ZN(new_n12886_));
  NAND2_X1   g09987(.A1(new_n12886_), .A2(new_n6460_), .ZN(new_n12887_));
  INV_X1     g09988(.I(new_n12787_), .ZN(new_n12888_));
  NAND3_X1   g09989(.A1(new_n12888_), .A2(pi0223), .A3(new_n12887_), .ZN(new_n12889_));
  NOR3_X1    g09990(.A1(new_n12878_), .A2(new_n12868_), .A3(new_n6460_), .ZN(new_n12890_));
  INV_X1     g09991(.I(new_n12789_), .ZN(new_n12891_));
  OAI21_X1   g09992(.A1(new_n12890_), .A2(new_n12891_), .B(new_n12791_), .ZN(new_n12892_));
  AOI21_X1   g09993(.A1(new_n12892_), .A2(new_n12889_), .B(pi0299), .ZN(new_n12893_));
  NOR2_X1    g09994(.A1(new_n12893_), .A2(new_n12885_), .ZN(new_n12894_));
  NOR3_X1    g09995(.A1(new_n12894_), .A2(new_n3154_), .A3(new_n12854_), .ZN(new_n12895_));
  AOI21_X1   g09996(.A1(new_n12793_), .A2(pi0039), .B(new_n12853_), .ZN(new_n12896_));
  OAI21_X1   g09997(.A1(new_n12895_), .A2(new_n12896_), .B(new_n3172_), .ZN(new_n12897_));
  NOR2_X1    g09998(.A1(new_n5154_), .A2(new_n2926_), .ZN(new_n12898_));
  INV_X1     g09999(.I(new_n12898_), .ZN(new_n12899_));
  NOR2_X1    g10000(.A1(new_n12899_), .A2(new_n3172_), .ZN(new_n12900_));
  INV_X1     g10001(.I(new_n12900_), .ZN(new_n12901_));
  NAND2_X1   g10002(.A1(new_n12897_), .A2(new_n12901_), .ZN(new_n12902_));
  NAND2_X1   g10003(.A1(new_n7339_), .A2(pi0738), .ZN(new_n12903_));
  OAI21_X1   g10004(.A1(new_n12602_), .A2(pi0140), .B(new_n3154_), .ZN(new_n12904_));
  NOR2_X1    g10005(.A1(new_n12644_), .A2(new_n7339_), .ZN(new_n12905_));
  AOI21_X1   g10006(.A1(new_n5427_), .A2(new_n12281_), .B(new_n5095_), .ZN(new_n12906_));
  INV_X1     g10007(.I(new_n12906_), .ZN(new_n12907_));
  AOI21_X1   g10008(.A1(new_n5217_), .A2(new_n12907_), .B(new_n12382_), .ZN(new_n12908_));
  AOI21_X1   g10009(.A1(new_n5427_), .A2(new_n12303_), .B(new_n12280_), .ZN(new_n12909_));
  NOR3_X1    g10010(.A1(new_n12362_), .A2(new_n5095_), .A3(new_n12909_), .ZN(new_n12910_));
  INV_X1     g10011(.I(new_n12362_), .ZN(new_n12911_));
  AOI21_X1   g10012(.A1(pi0680), .A2(new_n12909_), .B(new_n12911_), .ZN(new_n12912_));
  NOR2_X1    g10013(.A1(new_n12912_), .A2(new_n12910_), .ZN(new_n12913_));
  NOR2_X1    g10014(.A1(new_n12913_), .A2(new_n12908_), .ZN(new_n12914_));
  NOR2_X1    g10015(.A1(new_n12373_), .A2(new_n12908_), .ZN(new_n12915_));
  NOR4_X1    g10016(.A1(new_n12914_), .A2(pi0223), .A3(new_n6460_), .A4(new_n12915_), .ZN(new_n12916_));
  NAND2_X1   g10017(.A1(new_n12453_), .A2(new_n5095_), .ZN(new_n12917_));
  INV_X1     g10018(.I(new_n12329_), .ZN(new_n12918_));
  OAI21_X1   g10019(.A1(new_n12453_), .A2(new_n12918_), .B(pi0680), .ZN(new_n12919_));
  OAI21_X1   g10020(.A1(new_n12329_), .A2(new_n5427_), .B(new_n12906_), .ZN(new_n12920_));
  INV_X1     g10021(.I(new_n12920_), .ZN(new_n12921_));
  NOR2_X1    g10022(.A1(new_n12921_), .A2(new_n12129_), .ZN(new_n12922_));
  OAI22_X1   g10023(.A1(new_n12919_), .A2(new_n12461_), .B1(new_n12917_), .B2(new_n12922_), .ZN(new_n12923_));
  INV_X1     g10024(.I(new_n12424_), .ZN(new_n12924_));
  MUX2_X1    g10025(.I0(new_n12322_), .I1(new_n12321_), .S(new_n12129_), .Z(new_n12925_));
  AOI21_X1   g10026(.A1(new_n12925_), .A2(pi0680), .B(new_n12924_), .ZN(new_n12926_));
  AOI21_X1   g10027(.A1(new_n12926_), .A2(new_n3155_), .B(new_n5141_), .ZN(new_n12927_));
  NAND2_X1   g10028(.A1(new_n12923_), .A2(new_n12927_), .ZN(new_n12928_));
  AOI21_X1   g10029(.A1(new_n12504_), .A2(new_n11885_), .B(pi0223), .ZN(new_n12929_));
  AOI21_X1   g10030(.A1(new_n12928_), .A2(new_n12929_), .B(new_n12916_), .ZN(new_n12930_));
  NOR4_X1    g10031(.A1(new_n12914_), .A2(pi0215), .A3(new_n6445_), .A4(new_n12915_), .ZN(new_n12931_));
  AOI21_X1   g10032(.A1(new_n12926_), .A2(new_n3285_), .B(new_n5094_), .ZN(new_n12932_));
  NOR3_X1    g10033(.A1(new_n11884_), .A2(new_n2926_), .A3(new_n3285_), .ZN(new_n12933_));
  AOI21_X1   g10034(.A1(new_n12681_), .A2(new_n12933_), .B(pi0215), .ZN(new_n12934_));
  AOI21_X1   g10035(.A1(new_n12923_), .A2(new_n12932_), .B(new_n12934_), .ZN(new_n12935_));
  NOR2_X1    g10036(.A1(new_n12935_), .A2(new_n12931_), .ZN(new_n12936_));
  MUX2_X1    g10037(.I0(new_n12936_), .I1(new_n12930_), .S(new_n2587_), .Z(new_n12937_));
  INV_X1     g10038(.I(new_n12244_), .ZN(new_n12938_));
  NOR3_X1    g10039(.A1(new_n12938_), .A2(new_n5095_), .A3(new_n12685_), .ZN(new_n12939_));
  NAND3_X1   g10040(.A1(new_n12939_), .A2(pi0223), .A3(new_n12254_), .ZN(new_n12940_));
  NAND2_X1   g10041(.A1(new_n12495_), .A2(new_n12162_), .ZN(new_n12941_));
  AOI21_X1   g10042(.A1(new_n12941_), .A2(new_n12129_), .B(new_n5095_), .ZN(new_n12942_));
  NOR2_X1    g10043(.A1(new_n12159_), .A2(new_n5106_), .ZN(new_n12943_));
  AOI21_X1   g10044(.A1(new_n12941_), .A2(new_n5106_), .B(new_n12943_), .ZN(new_n12944_));
  OAI21_X1   g10045(.A1(new_n12129_), .A2(new_n12944_), .B(new_n12942_), .ZN(new_n12945_));
  NOR2_X1    g10046(.A1(new_n11885_), .A2(new_n12129_), .ZN(new_n12946_));
  AOI21_X1   g10047(.A1(new_n12196_), .A2(new_n12946_), .B(new_n12200_), .ZN(new_n12947_));
  AND3_X2    g10048(.A1(new_n12945_), .A2(new_n2614_), .A3(new_n5141_), .Z(new_n12948_));
  OAI21_X1   g10049(.A1(new_n12505_), .A2(new_n11885_), .B(new_n2604_), .ZN(new_n12949_));
  OAI21_X1   g10050(.A1(new_n12948_), .A2(new_n12949_), .B(new_n12940_), .ZN(new_n12950_));
  NOR3_X1    g10051(.A1(new_n12938_), .A2(new_n12677_), .A3(pi0680), .ZN(new_n12951_));
  AOI21_X1   g10052(.A1(new_n12951_), .A2(new_n12254_), .B(new_n2566_), .ZN(new_n12952_));
  NOR2_X1    g10053(.A1(new_n12952_), .A2(pi0299), .ZN(new_n12953_));
  NAND2_X1   g10054(.A1(new_n12950_), .A2(new_n12953_), .ZN(new_n12954_));
  INV_X1     g10055(.I(new_n12954_), .ZN(new_n12955_));
  MUX2_X1    g10056(.I0(new_n12955_), .I1(new_n12937_), .S(new_n7339_), .Z(new_n12956_));
  AOI22_X1   g10057(.A1(new_n12956_), .A2(pi0039), .B1(new_n12904_), .B2(new_n12905_), .ZN(new_n12957_));
  NAND2_X1   g10058(.A1(new_n3172_), .A2(new_n11881_), .ZN(new_n12959_));
  OAI22_X1   g10059(.A1(new_n12957_), .A2(new_n12959_), .B1(new_n12902_), .B2(new_n12903_), .ZN(new_n12960_));
  NAND3_X1   g10060(.A1(new_n12960_), .A2(new_n3231_), .A3(new_n12836_), .ZN(new_n12961_));
  AOI21_X1   g10061(.A1(new_n12960_), .A2(new_n3231_), .B(new_n12836_), .ZN(new_n12962_));
  INV_X1     g10062(.I(new_n12962_), .ZN(new_n12963_));
  NAND3_X1   g10063(.A1(new_n12963_), .A2(pi0625), .A3(new_n12961_), .ZN(new_n12964_));
  AOI21_X1   g10064(.A1(new_n12897_), .A2(new_n12901_), .B(new_n3232_), .ZN(new_n12965_));
  NOR2_X1    g10065(.A1(new_n12965_), .A2(pi0140), .ZN(new_n12966_));
  AOI21_X1   g10066(.A1(new_n12966_), .A2(pi0625), .B(pi1153), .ZN(new_n12967_));
  NAND3_X1   g10067(.A1(new_n12964_), .A2(pi0608), .A3(new_n12967_), .ZN(new_n12968_));
  AOI21_X1   g10068(.A1(new_n12845_), .A2(new_n12850_), .B(new_n12968_), .ZN(new_n12969_));
  INV_X1     g10069(.I(pi0625), .ZN(new_n12970_));
  NOR3_X1    g10070(.A1(new_n12843_), .A2(new_n3232_), .A3(new_n12838_), .ZN(new_n12971_));
  AOI21_X1   g10071(.A1(new_n12833_), .A2(new_n3231_), .B(new_n12836_), .ZN(new_n12972_));
  NOR3_X1    g10072(.A1(new_n12971_), .A2(new_n12970_), .A3(new_n12972_), .ZN(new_n12973_));
  INV_X1     g10073(.I(new_n12961_), .ZN(new_n12974_));
  NOR3_X1    g10074(.A1(new_n12974_), .A2(new_n12970_), .A3(new_n12962_), .ZN(new_n12975_));
  OAI21_X1   g10075(.A1(new_n12966_), .A2(pi0625), .B(new_n11893_), .ZN(new_n12976_));
  NOR2_X1    g10076(.A1(pi0608), .A2(pi1153), .ZN(new_n12977_));
  INV_X1     g10077(.I(new_n12977_), .ZN(new_n12978_));
  AOI21_X1   g10078(.A1(new_n12848_), .A2(pi0625), .B(new_n12978_), .ZN(new_n12979_));
  OAI21_X1   g10079(.A1(new_n12975_), .A2(new_n12976_), .B(new_n12979_), .ZN(new_n12980_));
  NOR2_X1    g10080(.A1(new_n12973_), .A2(new_n12980_), .ZN(new_n12981_));
  NOR2_X1    g10081(.A1(new_n12969_), .A2(new_n12981_), .ZN(new_n12982_));
  NOR3_X1    g10082(.A1(new_n12982_), .A2(new_n11891_), .A3(new_n12835_), .ZN(new_n12983_));
  AOI21_X1   g10083(.A1(new_n12982_), .A2(pi0778), .B(new_n12834_), .ZN(new_n12984_));
  NOR3_X1    g10084(.A1(new_n12983_), .A2(new_n12984_), .A3(pi0785), .ZN(new_n12985_));
  INV_X1     g10085(.I(new_n12985_), .ZN(new_n12986_));
  MUX2_X1    g10086(.I0(new_n12982_), .I1(new_n12834_), .S(new_n11891_), .Z(new_n12987_));
  NOR3_X1    g10087(.A1(new_n12974_), .A2(pi0778), .A3(new_n12962_), .ZN(new_n12988_));
  INV_X1     g10088(.I(new_n12988_), .ZN(new_n12989_));
  NOR4_X1    g10089(.A1(new_n12975_), .A2(pi0625), .A3(pi1153), .A4(new_n12966_), .ZN(new_n12990_));
  NOR3_X1    g10090(.A1(new_n12990_), .A2(new_n11891_), .A3(new_n12989_), .ZN(new_n12991_));
  NAND3_X1   g10091(.A1(new_n12964_), .A2(new_n12967_), .A3(new_n12976_), .ZN(new_n12992_));
  AOI21_X1   g10092(.A1(new_n12992_), .A2(pi0778), .B(new_n12988_), .ZN(new_n12993_));
  OAI21_X1   g10093(.A1(new_n12991_), .A2(new_n12993_), .B(new_n11903_), .ZN(new_n12994_));
  INV_X1     g10094(.I(new_n12966_), .ZN(new_n12995_));
  NOR2_X1    g10095(.A1(new_n11914_), .A2(pi0609), .ZN(new_n12996_));
  INV_X1     g10096(.I(new_n12996_), .ZN(new_n12997_));
  NAND2_X1   g10097(.A1(new_n12995_), .A2(new_n12997_), .ZN(new_n12998_));
  NOR2_X1    g10098(.A1(new_n12848_), .A2(new_n11914_), .ZN(new_n12999_));
  NAND2_X1   g10099(.A1(new_n12999_), .A2(new_n11903_), .ZN(new_n13000_));
  AOI21_X1   g10100(.A1(new_n13000_), .A2(new_n12998_), .B(pi1155), .ZN(new_n13001_));
  OAI21_X1   g10101(.A1(new_n13001_), .A2(new_n11923_), .B(pi0609), .ZN(new_n13002_));
  AOI21_X1   g10102(.A1(new_n12994_), .A2(pi1155), .B(new_n13002_), .ZN(new_n13003_));
  AOI21_X1   g10103(.A1(new_n12834_), .A2(pi0625), .B(new_n12849_), .ZN(new_n13004_));
  OAI22_X1   g10104(.A1(new_n13004_), .A2(new_n12968_), .B1(new_n12973_), .B2(new_n12980_), .ZN(new_n13005_));
  NAND3_X1   g10105(.A1(new_n13005_), .A2(pi0778), .A3(new_n12834_), .ZN(new_n13006_));
  OAI21_X1   g10106(.A1(new_n13005_), .A2(new_n11891_), .B(new_n12835_), .ZN(new_n13007_));
  NAND3_X1   g10107(.A1(new_n13007_), .A2(new_n13006_), .A3(new_n11903_), .ZN(new_n13008_));
  NOR2_X1    g10108(.A1(new_n12991_), .A2(new_n12993_), .ZN(new_n13009_));
  INV_X1     g10109(.I(new_n11915_), .ZN(new_n13010_));
  AOI22_X1   g10110(.A1(new_n12999_), .A2(pi0609), .B1(new_n13010_), .B2(new_n12995_), .ZN(new_n13011_));
  NOR2_X1    g10111(.A1(new_n11923_), .A2(pi1155), .ZN(new_n13012_));
  OAI21_X1   g10112(.A1(new_n13009_), .A2(new_n11903_), .B(new_n13012_), .ZN(new_n13013_));
  INV_X1     g10113(.I(new_n13013_), .ZN(new_n13014_));
  AOI22_X1   g10114(.A1(new_n13008_), .A2(new_n13014_), .B1(new_n12987_), .B2(new_n13003_), .ZN(new_n13015_));
  NOR3_X1    g10115(.A1(new_n13015_), .A2(new_n11870_), .A3(new_n12986_), .ZN(new_n13016_));
  NAND3_X1   g10116(.A1(new_n13003_), .A2(new_n13007_), .A3(new_n13006_), .ZN(new_n13017_));
  NOR3_X1    g10117(.A1(new_n12983_), .A2(new_n12984_), .A3(pi0609), .ZN(new_n13018_));
  OAI21_X1   g10118(.A1(new_n13018_), .A2(new_n13013_), .B(new_n13017_), .ZN(new_n13019_));
  AOI21_X1   g10119(.A1(new_n13019_), .A2(pi0785), .B(new_n12985_), .ZN(new_n13020_));
  NOR3_X1    g10120(.A1(new_n13020_), .A2(new_n13016_), .A3(pi0781), .ZN(new_n13021_));
  INV_X1     g10121(.I(new_n13021_), .ZN(new_n13022_));
  NOR2_X1    g10122(.A1(new_n13020_), .A2(new_n13016_), .ZN(new_n13023_));
  INV_X1     g10123(.I(new_n11938_), .ZN(new_n13024_));
  NAND2_X1   g10124(.A1(new_n12966_), .A2(new_n13024_), .ZN(new_n13025_));
  OAI21_X1   g10125(.A1(new_n13009_), .A2(new_n13024_), .B(new_n13025_), .ZN(new_n13026_));
  AOI21_X1   g10126(.A1(new_n13026_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n13027_));
  AOI21_X1   g10127(.A1(new_n12966_), .A2(new_n11914_), .B(pi0785), .ZN(new_n13028_));
  INV_X1     g10128(.I(new_n13028_), .ZN(new_n13029_));
  AOI21_X1   g10129(.A1(new_n12848_), .A2(new_n11924_), .B(new_n13029_), .ZN(new_n13030_));
  INV_X1     g10130(.I(new_n13030_), .ZN(new_n13031_));
  NOR2_X1    g10131(.A1(new_n13011_), .A2(new_n11912_), .ZN(new_n13032_));
  OAI21_X1   g10132(.A1(new_n13032_), .A2(new_n13001_), .B(pi0785), .ZN(new_n13033_));
  OR2_X2     g10133(.A1(new_n13033_), .A2(new_n13031_), .Z(new_n13034_));
  NAND2_X1   g10134(.A1(new_n13033_), .A2(new_n13031_), .ZN(new_n13035_));
  NAND3_X1   g10135(.A1(new_n13034_), .A2(pi0618), .A3(new_n13035_), .ZN(new_n13036_));
  NAND2_X1   g10136(.A1(new_n12966_), .A2(pi0618), .ZN(new_n13037_));
  NAND4_X1   g10137(.A1(new_n13036_), .A2(pi0627), .A3(new_n11950_), .A4(new_n13037_), .ZN(new_n13038_));
  NAND2_X1   g10138(.A1(new_n13038_), .A2(pi0618), .ZN(new_n13039_));
  NOR2_X1    g10139(.A1(new_n13039_), .A2(new_n13027_), .ZN(new_n13040_));
  NAND3_X1   g10140(.A1(new_n13019_), .A2(pi0785), .A3(new_n12985_), .ZN(new_n13041_));
  OAI21_X1   g10141(.A1(new_n13015_), .A2(new_n11870_), .B(new_n12986_), .ZN(new_n13042_));
  NAND3_X1   g10142(.A1(new_n13041_), .A2(new_n13042_), .A3(new_n11934_), .ZN(new_n13043_));
  INV_X1     g10143(.I(new_n13026_), .ZN(new_n13044_));
  NOR2_X1    g10144(.A1(new_n13044_), .A2(new_n11934_), .ZN(new_n13045_));
  AOI21_X1   g10145(.A1(new_n12995_), .A2(new_n11934_), .B(pi1154), .ZN(new_n13046_));
  AOI21_X1   g10146(.A1(new_n13036_), .A2(new_n13046_), .B(pi0627), .ZN(new_n13047_));
  NOR3_X1    g10147(.A1(new_n13045_), .A2(new_n13047_), .A3(pi1154), .ZN(new_n13048_));
  AOI22_X1   g10148(.A1(new_n13043_), .A2(new_n13048_), .B1(new_n13023_), .B2(new_n13040_), .ZN(new_n13049_));
  NOR3_X1    g10149(.A1(new_n13049_), .A2(new_n11969_), .A3(new_n13022_), .ZN(new_n13050_));
  NAND3_X1   g10150(.A1(new_n13041_), .A2(new_n13042_), .A3(new_n13040_), .ZN(new_n13051_));
  NOR3_X1    g10151(.A1(new_n13020_), .A2(new_n13016_), .A3(pi0618), .ZN(new_n13052_));
  INV_X1     g10152(.I(new_n13048_), .ZN(new_n13053_));
  OAI21_X1   g10153(.A1(new_n13052_), .A2(new_n13053_), .B(new_n13051_), .ZN(new_n13054_));
  AOI21_X1   g10154(.A1(new_n13054_), .A2(pi0781), .B(new_n13021_), .ZN(new_n13055_));
  NOR3_X1    g10155(.A1(new_n13050_), .A2(new_n13055_), .A3(pi0789), .ZN(new_n13056_));
  INV_X1     g10156(.I(new_n13056_), .ZN(new_n13057_));
  NOR2_X1    g10157(.A1(new_n13050_), .A2(new_n13055_), .ZN(new_n13058_));
  XOR2_X1    g10158(.A1(new_n13033_), .A2(new_n13031_), .Z(new_n13059_));
  NAND3_X1   g10159(.A1(new_n12995_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n13060_));
  MUX2_X1    g10160(.I0(new_n13060_), .I1(new_n13059_), .S(new_n11969_), .Z(new_n13061_));
  NAND2_X1   g10161(.A1(new_n13061_), .A2(pi0619), .ZN(new_n13062_));
  AOI21_X1   g10162(.A1(new_n12966_), .A2(pi0619), .B(pi1159), .ZN(new_n13063_));
  AND3_X2    g10163(.A1(new_n13062_), .A2(pi0648), .A3(new_n13063_), .Z(new_n13064_));
  NOR2_X1    g10164(.A1(new_n12966_), .A2(new_n11961_), .ZN(new_n13065_));
  AOI21_X1   g10165(.A1(new_n13044_), .A2(new_n11961_), .B(new_n13065_), .ZN(new_n13066_));
  NOR3_X1    g10166(.A1(new_n13064_), .A2(new_n11967_), .A3(pi1159), .ZN(new_n13067_));
  NAND3_X1   g10167(.A1(new_n13054_), .A2(pi0781), .A3(new_n13021_), .ZN(new_n13068_));
  OAI21_X1   g10168(.A1(new_n13049_), .A2(new_n11969_), .B(new_n13022_), .ZN(new_n13069_));
  NAND3_X1   g10169(.A1(new_n13069_), .A2(new_n13068_), .A3(new_n11967_), .ZN(new_n13070_));
  AOI21_X1   g10170(.A1(new_n12995_), .A2(new_n11967_), .B(pi1159), .ZN(new_n13071_));
  NAND2_X1   g10171(.A1(new_n13062_), .A2(new_n13071_), .ZN(new_n13072_));
  NAND2_X1   g10172(.A1(new_n13072_), .A2(new_n11966_), .ZN(new_n13073_));
  AOI21_X1   g10173(.A1(new_n13066_), .A2(pi0619), .B(pi1159), .ZN(new_n13074_));
  NAND2_X1   g10174(.A1(new_n13073_), .A2(new_n13074_), .ZN(new_n13075_));
  INV_X1     g10175(.I(new_n13075_), .ZN(new_n13076_));
  AOI22_X1   g10176(.A1(new_n13070_), .A2(new_n13076_), .B1(new_n13058_), .B2(new_n13067_), .ZN(new_n13077_));
  NOR3_X1    g10177(.A1(new_n13077_), .A2(new_n11985_), .A3(new_n13057_), .ZN(new_n13078_));
  NAND3_X1   g10178(.A1(new_n13069_), .A2(new_n13068_), .A3(new_n13067_), .ZN(new_n13079_));
  NOR3_X1    g10179(.A1(new_n13050_), .A2(new_n13055_), .A3(pi0619), .ZN(new_n13080_));
  OAI21_X1   g10180(.A1(new_n13080_), .A2(new_n13075_), .B(new_n13079_), .ZN(new_n13081_));
  AOI21_X1   g10181(.A1(new_n13081_), .A2(pi0789), .B(new_n13056_), .ZN(new_n13082_));
  NOR2_X1    g10182(.A1(new_n13078_), .A2(new_n13082_), .ZN(new_n13083_));
  INV_X1     g10183(.I(new_n13083_), .ZN(new_n13084_));
  NAND3_X1   g10184(.A1(new_n13081_), .A2(pi0789), .A3(new_n13056_), .ZN(new_n13085_));
  OAI21_X1   g10185(.A1(new_n13077_), .A2(new_n11985_), .B(new_n13057_), .ZN(new_n13086_));
  NOR2_X1    g10186(.A1(new_n12995_), .A2(new_n12014_), .ZN(new_n13087_));
  AOI21_X1   g10187(.A1(new_n13066_), .A2(new_n12014_), .B(new_n13087_), .ZN(new_n13088_));
  NOR2_X1    g10188(.A1(new_n11989_), .A2(pi0626), .ZN(new_n13089_));
  INV_X1     g10189(.I(new_n13089_), .ZN(new_n13090_));
  AOI21_X1   g10190(.A1(new_n13086_), .A2(new_n13085_), .B(new_n13090_), .ZN(new_n13091_));
  NOR2_X1    g10191(.A1(new_n11994_), .A2(pi0641), .ZN(new_n13092_));
  INV_X1     g10192(.I(new_n13092_), .ZN(new_n13093_));
  AOI21_X1   g10193(.A1(new_n13086_), .A2(new_n13085_), .B(new_n13093_), .ZN(new_n13094_));
  INV_X1     g10194(.I(new_n12016_), .ZN(new_n13095_));
  NAND3_X1   g10195(.A1(new_n12995_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n13096_));
  MUX2_X1    g10196(.I0(new_n13096_), .I1(new_n13061_), .S(new_n11985_), .Z(new_n13097_));
  NAND2_X1   g10197(.A1(new_n13097_), .A2(pi0626), .ZN(new_n13098_));
  AOI21_X1   g10198(.A1(new_n12995_), .A2(new_n11994_), .B(pi1158), .ZN(new_n13099_));
  NAND2_X1   g10199(.A1(new_n13098_), .A2(new_n13099_), .ZN(new_n13100_));
  AOI21_X1   g10200(.A1(new_n12966_), .A2(pi0626), .B(pi1158), .ZN(new_n13101_));
  NAND2_X1   g10201(.A1(new_n13098_), .A2(new_n13101_), .ZN(new_n13102_));
  INV_X1     g10202(.I(new_n13102_), .ZN(new_n13103_));
  AOI22_X1   g10203(.A1(new_n13103_), .A2(new_n12018_), .B1(new_n13100_), .B2(new_n13095_), .ZN(new_n13104_));
  INV_X1     g10204(.I(new_n13104_), .ZN(new_n13105_));
  NOR3_X1    g10205(.A1(new_n13091_), .A2(new_n13094_), .A3(new_n13105_), .ZN(new_n13106_));
  NOR3_X1    g10206(.A1(new_n13106_), .A2(new_n11986_), .A3(new_n13084_), .ZN(new_n13107_));
  AOI21_X1   g10207(.A1(new_n13106_), .A2(pi0788), .B(new_n13083_), .ZN(new_n13108_));
  NOR2_X1    g10208(.A1(new_n13107_), .A2(new_n13108_), .ZN(new_n13109_));
  NAND2_X1   g10209(.A1(new_n13097_), .A2(new_n11986_), .ZN(new_n13110_));
  AOI21_X1   g10210(.A1(new_n13103_), .A2(new_n13100_), .B(new_n11986_), .ZN(new_n13111_));
  XNOR2_X1   g10211(.A1(new_n13111_), .A2(new_n13110_), .ZN(new_n13112_));
  OR2_X2     g10212(.A1(new_n13112_), .A2(pi0628), .Z(new_n13113_));
  INV_X1     g10213(.I(new_n11992_), .ZN(new_n13114_));
  NOR2_X1    g10214(.A1(new_n12966_), .A2(new_n13114_), .ZN(new_n13115_));
  AOI21_X1   g10215(.A1(new_n13088_), .A2(new_n13114_), .B(new_n13115_), .ZN(new_n13116_));
  NOR3_X1    g10216(.A1(new_n12995_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n13117_));
  OAI21_X1   g10217(.A1(new_n13117_), .A2(new_n12030_), .B(pi0628), .ZN(new_n13118_));
  AOI21_X1   g10218(.A1(new_n13113_), .A2(pi1156), .B(new_n13118_), .ZN(new_n13119_));
  NOR2_X1    g10219(.A1(new_n13112_), .A2(new_n12031_), .ZN(new_n13120_));
  NOR2_X1    g10220(.A1(new_n12030_), .A2(pi0628), .ZN(new_n13121_));
  OAI21_X1   g10221(.A1(new_n13120_), .A2(pi1156), .B(new_n13121_), .ZN(new_n13122_));
  INV_X1     g10222(.I(new_n13122_), .ZN(new_n13123_));
  OAI22_X1   g10223(.A1(new_n13107_), .A2(new_n13108_), .B1(new_n13119_), .B2(new_n13123_), .ZN(new_n13124_));
  MUX2_X1    g10224(.I0(new_n13124_), .I1(new_n13109_), .S(new_n11868_), .Z(new_n13125_));
  OAI21_X1   g10225(.A1(new_n13078_), .A2(new_n13082_), .B(new_n13089_), .ZN(new_n13126_));
  OAI21_X1   g10226(.A1(new_n13078_), .A2(new_n13082_), .B(new_n13092_), .ZN(new_n13127_));
  NAND3_X1   g10227(.A1(new_n13126_), .A2(new_n13127_), .A3(new_n13104_), .ZN(new_n13128_));
  NAND3_X1   g10228(.A1(new_n13128_), .A2(pi0788), .A3(new_n13083_), .ZN(new_n13129_));
  OAI21_X1   g10229(.A1(new_n13128_), .A2(new_n11986_), .B(new_n13084_), .ZN(new_n13130_));
  INV_X1     g10230(.I(new_n13119_), .ZN(new_n13131_));
  AOI22_X1   g10231(.A1(new_n13130_), .A2(new_n13129_), .B1(new_n13131_), .B2(new_n13122_), .ZN(new_n13132_));
  NAND3_X1   g10232(.A1(new_n13132_), .A2(pi0792), .A3(new_n13109_), .ZN(new_n13133_));
  MUX2_X1    g10233(.I0(new_n13128_), .I1(new_n13084_), .S(new_n11986_), .Z(new_n13134_));
  OAI21_X1   g10234(.A1(new_n13132_), .A2(new_n11868_), .B(new_n13134_), .ZN(new_n13135_));
  NOR2_X1    g10235(.A1(new_n12966_), .A2(new_n12054_), .ZN(new_n13136_));
  AOI21_X1   g10236(.A1(new_n13112_), .A2(new_n12054_), .B(new_n13136_), .ZN(new_n13137_));
  AOI21_X1   g10237(.A1(new_n13137_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n13138_));
  NOR4_X1    g10238(.A1(new_n13116_), .A2(new_n12031_), .A3(pi1156), .A4(new_n12966_), .ZN(new_n13139_));
  NOR2_X1    g10239(.A1(new_n13139_), .A2(new_n13117_), .ZN(new_n13140_));
  MUX2_X1    g10240(.I0(new_n13140_), .I1(new_n13116_), .S(new_n11868_), .Z(new_n13141_));
  NAND2_X1   g10241(.A1(new_n13141_), .A2(pi0647), .ZN(new_n13142_));
  INV_X1     g10242(.I(new_n13142_), .ZN(new_n13143_));
  NOR2_X1    g10243(.A1(new_n12995_), .A2(new_n12061_), .ZN(new_n13144_));
  NOR4_X1    g10244(.A1(new_n13143_), .A2(new_n12060_), .A3(pi1157), .A4(new_n13144_), .ZN(new_n13145_));
  NOR3_X1    g10245(.A1(new_n13138_), .A2(new_n12061_), .A3(new_n13145_), .ZN(new_n13146_));
  NAND3_X1   g10246(.A1(new_n13135_), .A2(new_n13133_), .A3(new_n13146_), .ZN(new_n13147_));
  NOR3_X1    g10247(.A1(new_n13124_), .A2(new_n11868_), .A3(new_n13134_), .ZN(new_n13148_));
  AOI21_X1   g10248(.A1(new_n13124_), .A2(pi0792), .B(new_n13109_), .ZN(new_n13149_));
  NOR3_X1    g10249(.A1(new_n13148_), .A2(new_n13149_), .A3(pi0647), .ZN(new_n13150_));
  AND2_X2    g10250(.A1(new_n13137_), .A2(pi0647), .Z(new_n13151_));
  AOI21_X1   g10251(.A1(new_n12995_), .A2(new_n12061_), .B(pi1157), .ZN(new_n13152_));
  NAND2_X1   g10252(.A1(new_n13142_), .A2(new_n13152_), .ZN(new_n13153_));
  NAND2_X1   g10253(.A1(new_n13153_), .A2(new_n12060_), .ZN(new_n13154_));
  INV_X1     g10254(.I(new_n13154_), .ZN(new_n13155_));
  NOR3_X1    g10255(.A1(new_n13151_), .A2(pi1157), .A3(new_n13155_), .ZN(new_n13156_));
  INV_X1     g10256(.I(new_n13156_), .ZN(new_n13157_));
  OAI21_X1   g10257(.A1(new_n13150_), .A2(new_n13157_), .B(new_n13147_), .ZN(new_n13158_));
  MUX2_X1    g10258(.I0(new_n13158_), .I1(new_n13125_), .S(new_n12048_), .Z(new_n13159_));
  NAND2_X1   g10259(.A1(new_n13141_), .A2(new_n12048_), .ZN(new_n13160_));
  NAND3_X1   g10260(.A1(new_n12995_), .A2(new_n12061_), .A3(new_n12049_), .ZN(new_n13161_));
  NAND2_X1   g10261(.A1(new_n13161_), .A2(pi0787), .ZN(new_n13162_));
  XOR2_X1    g10262(.A1(new_n13160_), .A2(new_n13162_), .Z(new_n13163_));
  NOR2_X1    g10263(.A1(new_n12995_), .A2(new_n12092_), .ZN(new_n13164_));
  AOI21_X1   g10264(.A1(new_n13137_), .A2(new_n12092_), .B(new_n13164_), .ZN(new_n13165_));
  INV_X1     g10265(.I(new_n13165_), .ZN(new_n13166_));
  NOR2_X1    g10266(.A1(pi0644), .A2(pi0715), .ZN(new_n13167_));
  NOR2_X1    g10267(.A1(pi0715), .A2(pi1160), .ZN(new_n13168_));
  INV_X1     g10268(.I(new_n13168_), .ZN(new_n13169_));
  AOI21_X1   g10269(.A1(new_n13166_), .A2(new_n13167_), .B(new_n13169_), .ZN(new_n13170_));
  OAI21_X1   g10270(.A1(new_n12082_), .A2(new_n13163_), .B(new_n13170_), .ZN(new_n13171_));
  AOI21_X1   g10271(.A1(new_n13159_), .A2(new_n12082_), .B(new_n13171_), .ZN(new_n13172_));
  INV_X1     g10272(.I(new_n13125_), .ZN(new_n13173_));
  NAND3_X1   g10273(.A1(new_n13135_), .A2(new_n13133_), .A3(new_n12061_), .ZN(new_n13174_));
  AOI22_X1   g10274(.A1(new_n13174_), .A2(new_n13156_), .B1(new_n13125_), .B2(new_n13146_), .ZN(new_n13175_));
  MUX2_X1    g10275(.I0(new_n13175_), .I1(new_n13173_), .S(new_n12048_), .Z(new_n13176_));
  INV_X1     g10276(.I(new_n13163_), .ZN(new_n13177_));
  NAND3_X1   g10277(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n13178_));
  NOR2_X1    g10278(.A1(new_n12096_), .A2(pi0790), .ZN(new_n13179_));
  OAI21_X1   g10279(.A1(new_n13165_), .A2(new_n13178_), .B(new_n13179_), .ZN(new_n13180_));
  NOR2_X1    g10280(.A1(new_n13180_), .A2(new_n13177_), .ZN(new_n13181_));
  OAI21_X1   g10281(.A1(new_n13176_), .A2(new_n12082_), .B(new_n13181_), .ZN(new_n13182_));
  NOR2_X1    g10282(.A1(new_n13172_), .A2(new_n13182_), .ZN(new_n13183_));
  INV_X1     g10283(.I(pi0832), .ZN(new_n13184_));
  NAND2_X1   g10284(.A1(po1038), .A2(new_n7339_), .ZN(new_n13185_));
  AOI21_X1   g10285(.A1(new_n13185_), .A2(new_n13184_), .B(po1038), .ZN(new_n13186_));
  OAI21_X1   g10286(.A1(new_n13159_), .A2(pi0790), .B(new_n13186_), .ZN(new_n13187_));
  OAI21_X1   g10287(.A1(new_n13183_), .A2(new_n13187_), .B(new_n12108_), .ZN(po0297));
  NOR2_X1    g10288(.A1(new_n2925_), .A2(pi0141), .ZN(new_n13189_));
  INV_X1     g10289(.I(pi0749), .ZN(new_n13190_));
  NOR2_X1    g10290(.A1(new_n11877_), .A2(new_n13190_), .ZN(new_n13191_));
  NOR2_X1    g10291(.A1(new_n13191_), .A2(new_n13189_), .ZN(new_n13192_));
  INV_X1     g10292(.I(new_n13192_), .ZN(new_n13193_));
  AOI21_X1   g10293(.A1(new_n11886_), .A2(pi0706), .B(new_n13189_), .ZN(new_n13194_));
  NOR2_X1    g10294(.A1(new_n13194_), .A2(new_n11874_), .ZN(new_n13195_));
  NOR2_X1    g10295(.A1(new_n13193_), .A2(new_n13195_), .ZN(new_n13196_));
  NOR2_X1    g10296(.A1(new_n13196_), .A2(pi0778), .ZN(new_n13197_));
  NAND2_X1   g10297(.A1(new_n13195_), .A2(pi0625), .ZN(new_n13198_));
  INV_X1     g10298(.I(pi0706), .ZN(new_n13199_));
  NOR2_X1    g10299(.A1(new_n11894_), .A2(pi0625), .ZN(new_n13200_));
  INV_X1     g10300(.I(new_n13200_), .ZN(new_n13201_));
  NOR2_X1    g10301(.A1(new_n13201_), .A2(new_n13199_), .ZN(new_n13202_));
  NOR4_X1    g10302(.A1(new_n13191_), .A2(pi0608), .A3(new_n11893_), .A4(new_n13189_), .ZN(new_n13203_));
  OAI21_X1   g10303(.A1(new_n13193_), .A2(new_n13195_), .B(new_n13198_), .ZN(new_n13204_));
  NOR3_X1    g10304(.A1(new_n13189_), .A2(pi0608), .A3(pi1153), .ZN(new_n13205_));
  AOI22_X1   g10305(.A1(new_n13204_), .A2(new_n13205_), .B1(new_n13198_), .B2(new_n13203_), .ZN(new_n13206_));
  NOR2_X1    g10306(.A1(new_n13206_), .A2(new_n11891_), .ZN(new_n13207_));
  XOR2_X1    g10307(.A1(new_n13207_), .A2(new_n13197_), .Z(new_n13208_));
  INV_X1     g10308(.I(new_n13208_), .ZN(new_n13209_));
  NAND2_X1   g10309(.A1(new_n13209_), .A2(new_n11870_), .ZN(new_n13210_));
  AOI21_X1   g10310(.A1(new_n13208_), .A2(new_n11903_), .B(pi1155), .ZN(new_n13211_));
  INV_X1     g10311(.I(new_n13194_), .ZN(new_n13212_));
  XOR2_X1    g10312(.A1(new_n13202_), .A2(pi1153), .Z(new_n13213_));
  NAND2_X1   g10313(.A1(new_n13213_), .A2(new_n13212_), .ZN(new_n13214_));
  OAI21_X1   g10314(.A1(new_n13202_), .A2(new_n13189_), .B(new_n11893_), .ZN(new_n13215_));
  AOI21_X1   g10315(.A1(new_n13214_), .A2(new_n13215_), .B(new_n11891_), .ZN(new_n13216_));
  NOR2_X1    g10316(.A1(new_n13194_), .A2(pi0778), .ZN(new_n13217_));
  OAI21_X1   g10317(.A1(new_n13216_), .A2(new_n13217_), .B(pi0609), .ZN(new_n13218_));
  AOI21_X1   g10318(.A1(new_n13193_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n13219_));
  NOR2_X1    g10319(.A1(new_n13219_), .A2(pi0660), .ZN(new_n13220_));
  OAI21_X1   g10320(.A1(new_n13211_), .A2(new_n13218_), .B(new_n13220_), .ZN(new_n13221_));
  NOR2_X1    g10321(.A1(new_n13216_), .A2(new_n13217_), .ZN(new_n13222_));
  NAND4_X1   g10322(.A1(new_n13209_), .A2(pi0609), .A3(new_n11912_), .A4(new_n13222_), .ZN(new_n13223_));
  NOR2_X1    g10323(.A1(new_n13192_), .A2(new_n11925_), .ZN(new_n13224_));
  AOI21_X1   g10324(.A1(new_n13224_), .A2(new_n11928_), .B(pi1155), .ZN(new_n13225_));
  NOR2_X1    g10325(.A1(new_n13225_), .A2(new_n11923_), .ZN(new_n13226_));
  NAND2_X1   g10326(.A1(new_n13223_), .A2(new_n13226_), .ZN(new_n13227_));
  NAND3_X1   g10327(.A1(new_n13227_), .A2(pi0785), .A3(new_n13221_), .ZN(new_n13228_));
  NAND2_X1   g10328(.A1(new_n13228_), .A2(new_n13210_), .ZN(new_n13229_));
  INV_X1     g10329(.I(new_n13229_), .ZN(new_n13230_));
  NOR4_X1    g10330(.A1(new_n13222_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n13231_));
  NOR2_X1    g10331(.A1(new_n13224_), .A2(pi0785), .ZN(new_n13232_));
  OAI21_X1   g10332(.A1(new_n13225_), .A2(new_n13219_), .B(pi0785), .ZN(new_n13233_));
  XNOR2_X1   g10333(.A1(new_n13233_), .A2(new_n13232_), .ZN(new_n13234_));
  INV_X1     g10334(.I(new_n13234_), .ZN(new_n13235_));
  NOR2_X1    g10335(.A1(new_n13235_), .A2(new_n11945_), .ZN(new_n13236_));
  OR3_X2     g10336(.A1(new_n13231_), .A2(new_n13236_), .A3(pi0627), .Z(new_n13237_));
  OAI21_X1   g10337(.A1(new_n13235_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n13238_));
  NOR2_X1    g10338(.A1(new_n13222_), .A2(new_n11939_), .ZN(new_n13239_));
  NOR4_X1    g10339(.A1(new_n13230_), .A2(new_n11934_), .A3(pi1154), .A4(new_n13239_), .ZN(new_n13240_));
  OAI21_X1   g10340(.A1(new_n13240_), .A2(new_n13238_), .B(new_n11949_), .ZN(new_n13241_));
  AOI21_X1   g10341(.A1(new_n13241_), .A2(new_n13237_), .B(new_n11969_), .ZN(new_n13242_));
  AOI21_X1   g10342(.A1(new_n11969_), .A2(new_n13229_), .B(new_n13242_), .ZN(new_n13243_));
  INV_X1     g10343(.I(new_n13239_), .ZN(new_n13244_));
  NOR2_X1    g10344(.A1(new_n13244_), .A2(new_n11962_), .ZN(new_n13245_));
  NOR4_X1    g10345(.A1(new_n13243_), .A2(new_n11967_), .A3(pi1159), .A4(new_n13245_), .ZN(new_n13246_));
  NOR2_X1    g10346(.A1(new_n13235_), .A2(pi0781), .ZN(new_n13247_));
  NOR2_X1    g10347(.A1(new_n13238_), .A2(new_n13236_), .ZN(new_n13248_));
  NOR2_X1    g10348(.A1(new_n13248_), .A2(new_n11969_), .ZN(new_n13249_));
  XOR2_X1    g10349(.A1(new_n13249_), .A2(new_n13247_), .Z(new_n13250_));
  INV_X1     g10350(.I(new_n13250_), .ZN(new_n13251_));
  NOR2_X1    g10351(.A1(new_n13251_), .A2(new_n11967_), .ZN(new_n13252_));
  INV_X1     g10352(.I(new_n13189_), .ZN(new_n13253_));
  OAI21_X1   g10353(.A1(new_n13253_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n13254_));
  NOR4_X1    g10354(.A1(new_n13246_), .A2(new_n11966_), .A3(new_n13252_), .A4(new_n13254_), .ZN(new_n13255_));
  NOR4_X1    g10355(.A1(new_n13244_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n13256_));
  OAI21_X1   g10356(.A1(new_n13189_), .A2(pi0619), .B(new_n11869_), .ZN(new_n13257_));
  OAI21_X1   g10357(.A1(new_n13252_), .A2(new_n13257_), .B(new_n11966_), .ZN(new_n13258_));
  NOR2_X1    g10358(.A1(new_n13258_), .A2(new_n13256_), .ZN(new_n13259_));
  AOI21_X1   g10359(.A1(new_n13243_), .A2(new_n11998_), .B(pi0789), .ZN(new_n13260_));
  OAI21_X1   g10360(.A1(new_n13255_), .A2(new_n13259_), .B(new_n13260_), .ZN(new_n13261_));
  NOR2_X1    g10361(.A1(new_n13251_), .A2(pi0789), .ZN(new_n13262_));
  NOR3_X1    g10362(.A1(new_n13189_), .A2(pi0619), .A3(pi1159), .ZN(new_n13263_));
  NOR2_X1    g10363(.A1(new_n13263_), .A2(new_n11985_), .ZN(new_n13264_));
  XOR2_X1    g10364(.A1(new_n13262_), .A2(new_n13264_), .Z(new_n13265_));
  INV_X1     g10365(.I(new_n13265_), .ZN(new_n13266_));
  MUX2_X1    g10366(.I0(new_n13266_), .I1(new_n13189_), .S(new_n12003_), .Z(new_n13267_));
  NAND2_X1   g10367(.A1(new_n13267_), .A2(new_n12002_), .ZN(new_n13268_));
  AOI21_X1   g10368(.A1(new_n13245_), .A2(new_n12021_), .B(new_n11986_), .ZN(new_n13269_));
  NAND2_X1   g10369(.A1(new_n13268_), .A2(new_n13269_), .ZN(new_n13270_));
  NAND2_X1   g10370(.A1(new_n13261_), .A2(new_n13270_), .ZN(new_n13271_));
  NOR2_X1    g10371(.A1(new_n13271_), .A2(pi0792), .ZN(new_n13272_));
  NOR2_X1    g10372(.A1(new_n13265_), .A2(pi0788), .ZN(new_n13273_));
  AOI21_X1   g10373(.A1(new_n13267_), .A2(pi0788), .B(new_n13273_), .ZN(new_n13274_));
  INV_X1     g10374(.I(new_n13274_), .ZN(new_n13275_));
  NOR4_X1    g10375(.A1(new_n13271_), .A2(new_n12031_), .A3(pi1156), .A4(new_n13275_), .ZN(new_n13276_));
  NOR2_X1    g10376(.A1(new_n2926_), .A2(new_n12031_), .ZN(new_n13277_));
  NOR2_X1    g10377(.A1(new_n13245_), .A2(new_n12034_), .ZN(new_n13278_));
  INV_X1     g10378(.I(new_n13278_), .ZN(new_n13279_));
  OAI21_X1   g10379(.A1(new_n13279_), .A2(new_n13277_), .B(new_n12026_), .ZN(new_n13280_));
  NAND2_X1   g10380(.A1(new_n13280_), .A2(pi0629), .ZN(new_n13281_));
  AOI21_X1   g10381(.A1(new_n13271_), .A2(new_n12031_), .B(pi1156), .ZN(new_n13282_));
  NOR3_X1    g10382(.A1(new_n13282_), .A2(new_n12031_), .A3(new_n13274_), .ZN(new_n13283_));
  AOI21_X1   g10383(.A1(new_n13278_), .A2(new_n12042_), .B(pi0629), .ZN(new_n13284_));
  OAI22_X1   g10384(.A1(new_n13283_), .A2(new_n13284_), .B1(new_n13276_), .B2(new_n13281_), .ZN(new_n13285_));
  AOI21_X1   g10385(.A1(new_n13285_), .A2(pi0792), .B(new_n13272_), .ZN(new_n13286_));
  NOR2_X1    g10386(.A1(new_n12054_), .A2(new_n13189_), .ZN(new_n13287_));
  AOI21_X1   g10387(.A1(new_n13274_), .A2(new_n12054_), .B(new_n13287_), .ZN(new_n13288_));
  XNOR2_X1   g10388(.A1(new_n13286_), .A2(new_n13288_), .ZN(new_n13289_));
  NOR2_X1    g10389(.A1(new_n13289_), .A2(new_n12061_), .ZN(new_n13290_));
  XOR2_X1    g10390(.A1(new_n13290_), .A2(new_n13286_), .Z(new_n13291_));
  NOR2_X1    g10391(.A1(new_n13291_), .A2(pi1157), .ZN(new_n13292_));
  NOR2_X1    g10392(.A1(new_n13279_), .A2(new_n12068_), .ZN(new_n13293_));
  NOR2_X1    g10393(.A1(new_n13293_), .A2(new_n12061_), .ZN(new_n13294_));
  INV_X1     g10394(.I(new_n13294_), .ZN(new_n13295_));
  AOI21_X1   g10395(.A1(new_n13253_), .A2(new_n12061_), .B(pi1157), .ZN(new_n13296_));
  NAND2_X1   g10396(.A1(new_n13295_), .A2(new_n13296_), .ZN(new_n13297_));
  NAND2_X1   g10397(.A1(new_n13297_), .A2(new_n12060_), .ZN(new_n13298_));
  NOR2_X1    g10398(.A1(new_n13292_), .A2(new_n13298_), .ZN(new_n13299_));
  XOR2_X1    g10399(.A1(new_n13290_), .A2(new_n13288_), .Z(new_n13300_));
  NOR2_X1    g10400(.A1(new_n13300_), .A2(new_n12049_), .ZN(new_n13301_));
  NAND2_X1   g10401(.A1(new_n13189_), .A2(pi0647), .ZN(new_n13302_));
  NAND4_X1   g10402(.A1(new_n13295_), .A2(pi0630), .A3(new_n12049_), .A4(new_n13302_), .ZN(new_n13303_));
  OAI21_X1   g10403(.A1(new_n13301_), .A2(new_n13303_), .B(pi0787), .ZN(new_n13304_));
  OAI22_X1   g10404(.A1(new_n13304_), .A2(new_n13299_), .B1(pi0787), .B2(new_n13286_), .ZN(new_n13305_));
  OAI21_X1   g10405(.A1(new_n13305_), .A2(pi0644), .B(new_n12099_), .ZN(new_n13306_));
  INV_X1     g10406(.I(new_n13293_), .ZN(new_n13307_));
  NAND3_X1   g10407(.A1(new_n13253_), .A2(new_n12061_), .A3(new_n12049_), .ZN(new_n13308_));
  MUX2_X1    g10408(.I0(new_n13308_), .I1(new_n13307_), .S(new_n12048_), .Z(new_n13309_));
  NOR2_X1    g10409(.A1(new_n13309_), .A2(new_n12082_), .ZN(new_n13310_));
  NOR2_X1    g10410(.A1(new_n12092_), .A2(new_n13253_), .ZN(new_n13311_));
  AOI21_X1   g10411(.A1(new_n13288_), .A2(new_n12092_), .B(new_n13311_), .ZN(new_n13312_));
  NAND4_X1   g10412(.A1(new_n13312_), .A2(pi0644), .A3(new_n12099_), .A4(new_n13253_), .ZN(new_n13313_));
  NAND2_X1   g10413(.A1(new_n13313_), .A2(new_n12081_), .ZN(new_n13314_));
  AOI21_X1   g10414(.A1(new_n13306_), .A2(new_n13310_), .B(new_n13314_), .ZN(new_n13315_));
  NAND4_X1   g10415(.A1(new_n13305_), .A2(pi0644), .A3(new_n12099_), .A4(new_n13309_), .ZN(new_n13316_));
  AOI21_X1   g10416(.A1(new_n12082_), .A2(new_n13253_), .B(new_n13312_), .ZN(new_n13317_));
  NOR4_X1    g10417(.A1(new_n13288_), .A2(pi0644), .A3(new_n12091_), .A4(new_n13253_), .ZN(new_n13318_));
  NOR3_X1    g10418(.A1(new_n13317_), .A2(pi0715), .A3(new_n13318_), .ZN(new_n13319_));
  AOI21_X1   g10419(.A1(new_n13316_), .A2(new_n13319_), .B(pi1160), .ZN(new_n13320_));
  NOR2_X1    g10420(.A1(new_n13320_), .A2(new_n13315_), .ZN(new_n13321_));
  NOR3_X1    g10421(.A1(new_n13321_), .A2(new_n11867_), .A3(new_n13305_), .ZN(new_n13322_));
  INV_X1     g10422(.I(new_n13305_), .ZN(new_n13323_));
  AOI21_X1   g10423(.A1(new_n13321_), .A2(pi0790), .B(new_n13323_), .ZN(new_n13324_));
  OAI21_X1   g10424(.A1(new_n13322_), .A2(new_n13324_), .B(pi0832), .ZN(new_n13325_));
  NAND2_X1   g10425(.A1(new_n3232_), .A2(pi0141), .ZN(new_n13326_));
  INV_X1     g10426(.I(new_n12442_), .ZN(new_n13327_));
  NAND3_X1   g10427(.A1(new_n12455_), .A2(new_n6445_), .A3(new_n12430_), .ZN(new_n13328_));
  NAND2_X1   g10428(.A1(new_n13328_), .A2(new_n3285_), .ZN(new_n13329_));
  OAI21_X1   g10429(.A1(new_n13329_), .A2(new_n12456_), .B(new_n13327_), .ZN(new_n13330_));
  AOI21_X1   g10430(.A1(new_n13330_), .A2(new_n12441_), .B(new_n2587_), .ZN(new_n13331_));
  AOI21_X1   g10431(.A1(new_n2587_), .A2(new_n12437_), .B(new_n13331_), .ZN(new_n13332_));
  INV_X1     g10432(.I(new_n13332_), .ZN(new_n13333_));
  OAI21_X1   g10433(.A1(new_n12494_), .A2(new_n12499_), .B(new_n12483_), .ZN(new_n13334_));
  NAND2_X1   g10434(.A1(new_n13334_), .A2(pi0299), .ZN(new_n13335_));
  INV_X1     g10435(.I(new_n12514_), .ZN(new_n13336_));
  NAND2_X1   g10436(.A1(new_n13336_), .A2(new_n13335_), .ZN(new_n13337_));
  AOI21_X1   g10437(.A1(new_n13337_), .A2(pi0141), .B(pi0749), .ZN(new_n13338_));
  OAI21_X1   g10438(.A1(new_n13333_), .A2(new_n11716_), .B(new_n13338_), .ZN(new_n13339_));
  NAND3_X1   g10439(.A1(new_n12668_), .A2(pi0141), .A3(new_n12665_), .ZN(new_n13340_));
  NOR4_X1    g10440(.A1(new_n12627_), .A2(pi0299), .A3(new_n12590_), .A4(new_n5101_), .ZN(new_n13341_));
  AOI21_X1   g10441(.A1(new_n12580_), .A2(pi0621), .B(pi0198), .ZN(new_n13342_));
  NOR3_X1    g10442(.A1(new_n12564_), .A2(pi0198), .A3(new_n11872_), .ZN(new_n13343_));
  NOR3_X1    g10443(.A1(new_n13343_), .A2(pi0299), .A3(new_n13342_), .ZN(new_n13344_));
  NOR4_X1    g10444(.A1(new_n12606_), .A2(new_n13344_), .A3(new_n12609_), .A4(pi0603), .ZN(new_n13345_));
  NOR2_X1    g10445(.A1(new_n13345_), .A2(new_n13341_), .ZN(new_n13346_));
  NAND2_X1   g10446(.A1(new_n12602_), .A2(new_n13346_), .ZN(new_n13347_));
  OAI21_X1   g10447(.A1(new_n12668_), .A2(new_n11716_), .B(new_n13347_), .ZN(new_n13348_));
  NAND2_X1   g10448(.A1(new_n13348_), .A2(new_n13340_), .ZN(new_n13349_));
  NAND2_X1   g10449(.A1(new_n13349_), .A2(pi0749), .ZN(new_n13350_));
  NOR2_X1    g10450(.A1(new_n13343_), .A2(new_n13342_), .ZN(new_n13351_));
  NOR2_X1    g10451(.A1(new_n13351_), .A2(pi0665), .ZN(new_n13352_));
  NAND2_X1   g10452(.A1(new_n12623_), .A2(pi0198), .ZN(new_n13353_));
  OAI21_X1   g10453(.A1(pi0198), .A2(new_n12621_), .B(new_n13353_), .ZN(new_n13354_));
  MUX2_X1    g10454(.I0(new_n13354_), .I1(new_n13352_), .S(pi0603), .Z(new_n13355_));
  NAND3_X1   g10455(.A1(new_n13355_), .A2(new_n2587_), .A3(pi0680), .ZN(new_n13356_));
  NOR2_X1    g10456(.A1(new_n12658_), .A2(pi0665), .ZN(new_n13357_));
  MUX2_X1    g10457(.I0(new_n12641_), .I1(new_n13357_), .S(pi0603), .Z(new_n13358_));
  NAND3_X1   g10458(.A1(new_n13358_), .A2(pi0299), .A3(pi0680), .ZN(new_n13359_));
  NAND2_X1   g10459(.A1(new_n13356_), .A2(new_n13359_), .ZN(new_n13360_));
  NAND2_X1   g10460(.A1(new_n13360_), .A2(pi0141), .ZN(new_n13361_));
  OAI21_X1   g10461(.A1(new_n12637_), .A2(new_n5095_), .B(new_n12657_), .ZN(new_n13362_));
  NAND2_X1   g10462(.A1(new_n3154_), .A2(new_n13190_), .ZN(new_n13363_));
  AOI21_X1   g10463(.A1(new_n13362_), .A2(pi0141), .B(new_n13363_), .ZN(new_n13364_));
  NAND3_X1   g10464(.A1(new_n13350_), .A2(new_n13361_), .A3(new_n13364_), .ZN(new_n13365_));
  AOI21_X1   g10465(.A1(new_n13365_), .A2(new_n3172_), .B(pi0039), .ZN(new_n13366_));
  INV_X1     g10466(.I(new_n12829_), .ZN(new_n13367_));
  INV_X1     g10467(.I(new_n12828_), .ZN(new_n13368_));
  NAND2_X1   g10468(.A1(new_n13368_), .A2(new_n11716_), .ZN(new_n13369_));
  OAI21_X1   g10469(.A1(new_n13190_), .A2(new_n13367_), .B(new_n13369_), .ZN(new_n13370_));
  INV_X1     g10470(.I(new_n13370_), .ZN(new_n13371_));
  NOR2_X1    g10471(.A1(new_n12110_), .A2(pi0039), .ZN(new_n13372_));
  NAND3_X1   g10472(.A1(new_n13372_), .A2(new_n3172_), .A3(new_n12113_), .ZN(new_n13373_));
  INV_X1     g10473(.I(new_n13373_), .ZN(new_n13374_));
  AOI21_X1   g10474(.A1(new_n13371_), .A2(new_n13374_), .B(new_n13199_), .ZN(new_n13375_));
  INV_X1     g10475(.I(new_n13375_), .ZN(new_n13376_));
  AOI21_X1   g10476(.A1(new_n13366_), .A2(new_n13339_), .B(new_n13376_), .ZN(new_n13377_));
  NAND2_X1   g10477(.A1(new_n12693_), .A2(pi0141), .ZN(new_n13378_));
  NAND2_X1   g10478(.A1(new_n12894_), .A2(new_n13190_), .ZN(new_n13379_));
  AOI21_X1   g10479(.A1(new_n13379_), .A2(new_n13378_), .B(pi0039), .ZN(new_n13380_));
  INV_X1     g10480(.I(new_n12824_), .ZN(new_n13381_));
  NOR2_X1    g10481(.A1(new_n12667_), .A2(pi0039), .ZN(new_n13382_));
  NOR4_X1    g10482(.A1(new_n13381_), .A2(new_n11716_), .A3(pi0749), .A4(new_n13382_), .ZN(new_n13383_));
  NOR2_X1    g10483(.A1(new_n12697_), .A2(pi0039), .ZN(new_n13384_));
  NOR3_X1    g10484(.A1(new_n13384_), .A2(pi0141), .A3(pi0749), .ZN(new_n13385_));
  NOR2_X1    g10485(.A1(new_n13371_), .A2(new_n3172_), .ZN(new_n13386_));
  NOR2_X1    g10486(.A1(new_n13386_), .A2(pi0038), .ZN(new_n13387_));
  OAI21_X1   g10487(.A1(new_n13383_), .A2(new_n13385_), .B(new_n13387_), .ZN(new_n13388_));
  NOR2_X1    g10488(.A1(new_n13388_), .A2(new_n13380_), .ZN(new_n13389_));
  OAI21_X1   g10489(.A1(new_n13389_), .A2(pi0706), .B(new_n3231_), .ZN(new_n13390_));
  OAI21_X1   g10490(.A1(new_n13377_), .A2(new_n13390_), .B(new_n13326_), .ZN(new_n13391_));
  INV_X1     g10491(.I(new_n13391_), .ZN(new_n13392_));
  NAND2_X1   g10492(.A1(new_n11716_), .A2(new_n13199_), .ZN(new_n13393_));
  OAI21_X1   g10493(.A1(new_n12902_), .A2(new_n13393_), .B(new_n3231_), .ZN(new_n13394_));
  MUX2_X1    g10494(.I0(new_n12954_), .I1(new_n12643_), .S(new_n3154_), .Z(new_n13395_));
  INV_X1     g10495(.I(new_n13395_), .ZN(new_n13396_));
  OAI21_X1   g10496(.A1(new_n12935_), .A2(new_n12931_), .B(pi0299), .ZN(new_n13397_));
  OAI21_X1   g10497(.A1(pi0299), .A2(new_n12930_), .B(new_n13397_), .ZN(new_n13398_));
  MUX2_X1    g10498(.I0(new_n13398_), .I1(new_n12657_), .S(new_n3154_), .Z(new_n13399_));
  NOR3_X1    g10499(.A1(new_n13399_), .A2(pi0141), .A3(new_n13396_), .ZN(new_n13400_));
  AOI21_X1   g10500(.A1(new_n13399_), .A2(new_n11716_), .B(new_n13395_), .ZN(new_n13401_));
  NOR2_X1    g10501(.A1(new_n5157_), .A2(new_n11894_), .ZN(new_n13402_));
  NOR2_X1    g10502(.A1(new_n13402_), .A2(new_n3172_), .ZN(new_n13403_));
  NOR2_X1    g10503(.A1(pi0038), .A2(pi0706), .ZN(new_n13404_));
  NAND3_X1   g10504(.A1(new_n13369_), .A2(new_n13403_), .A3(new_n13404_), .ZN(new_n13405_));
  NOR3_X1    g10505(.A1(new_n13400_), .A2(new_n13401_), .A3(new_n13405_), .ZN(new_n13406_));
  AOI22_X1   g10506(.A1(new_n13406_), .A2(new_n13394_), .B1(pi0141), .B2(new_n3232_), .ZN(new_n13407_));
  NOR2_X1    g10507(.A1(new_n12965_), .A2(pi0141), .ZN(new_n13408_));
  INV_X1     g10508(.I(new_n13408_), .ZN(new_n13409_));
  NOR4_X1    g10509(.A1(new_n13407_), .A2(pi0625), .A3(new_n12978_), .A4(new_n13409_), .ZN(new_n13410_));
  NOR2_X1    g10510(.A1(new_n3231_), .A2(pi0141), .ZN(new_n13411_));
  INV_X1     g10511(.I(new_n13411_), .ZN(new_n13412_));
  NOR3_X1    g10512(.A1(new_n13389_), .A2(new_n3232_), .A3(new_n13412_), .ZN(new_n13413_));
  INV_X1     g10513(.I(new_n13413_), .ZN(new_n13414_));
  OAI21_X1   g10514(.A1(new_n13389_), .A2(new_n3232_), .B(new_n13412_), .ZN(new_n13415_));
  NAND2_X1   g10515(.A1(new_n13414_), .A2(new_n13415_), .ZN(new_n13416_));
  INV_X1     g10516(.I(new_n13416_), .ZN(new_n13417_));
  NAND3_X1   g10517(.A1(new_n13391_), .A2(pi0625), .A3(new_n11893_), .ZN(new_n13418_));
  NAND2_X1   g10518(.A1(new_n11716_), .A2(new_n12970_), .ZN(new_n13419_));
  OAI21_X1   g10519(.A1(new_n12965_), .A2(new_n13419_), .B(pi1153), .ZN(new_n13420_));
  NAND2_X1   g10520(.A1(new_n13420_), .A2(pi0625), .ZN(new_n13421_));
  NOR2_X1    g10521(.A1(new_n13407_), .A2(new_n13421_), .ZN(new_n13422_));
  NOR3_X1    g10522(.A1(new_n11893_), .A2(pi0608), .A3(pi0625), .ZN(new_n13423_));
  NAND2_X1   g10523(.A1(new_n13391_), .A2(new_n13423_), .ZN(new_n13424_));
  OAI22_X1   g10524(.A1(new_n13418_), .A2(new_n13410_), .B1(new_n13424_), .B2(new_n13422_), .ZN(new_n13425_));
  NAND3_X1   g10525(.A1(new_n13425_), .A2(pi0778), .A3(new_n13392_), .ZN(new_n13426_));
  OAI21_X1   g10526(.A1(new_n13425_), .A2(new_n11891_), .B(new_n13391_), .ZN(new_n13427_));
  NAND2_X1   g10527(.A1(new_n13427_), .A2(new_n13426_), .ZN(new_n13428_));
  NOR2_X1    g10528(.A1(new_n13428_), .A2(pi0785), .ZN(new_n13429_));
  INV_X1     g10529(.I(new_n13429_), .ZN(new_n13430_));
  NOR2_X1    g10530(.A1(new_n13407_), .A2(pi0778), .ZN(new_n13431_));
  INV_X1     g10531(.I(new_n13431_), .ZN(new_n13432_));
  NOR2_X1    g10532(.A1(new_n11893_), .A2(pi0625), .ZN(new_n13433_));
  NOR2_X1    g10533(.A1(new_n12970_), .A2(pi1153), .ZN(new_n13434_));
  NOR2_X1    g10534(.A1(new_n13433_), .A2(new_n13434_), .ZN(new_n13435_));
  MUX2_X1    g10535(.I0(new_n13409_), .I1(new_n13407_), .S(new_n13435_), .Z(new_n13436_));
  OAI21_X1   g10536(.A1(new_n13436_), .A2(new_n11891_), .B(new_n13432_), .ZN(new_n13437_));
  AOI21_X1   g10537(.A1(new_n13437_), .A2(new_n11903_), .B(new_n11912_), .ZN(new_n13438_));
  INV_X1     g10538(.I(new_n13438_), .ZN(new_n13439_));
  NOR2_X1    g10539(.A1(new_n13408_), .A2(new_n12996_), .ZN(new_n13440_));
  INV_X1     g10540(.I(new_n13415_), .ZN(new_n13441_));
  NOR4_X1    g10541(.A1(new_n13441_), .A2(pi0609), .A3(new_n13413_), .A4(new_n11914_), .ZN(new_n13442_));
  OAI21_X1   g10542(.A1(new_n13442_), .A2(new_n13440_), .B(new_n11912_), .ZN(new_n13443_));
  NAND2_X1   g10543(.A1(new_n13443_), .A2(pi0660), .ZN(new_n13444_));
  NAND2_X1   g10544(.A1(new_n13444_), .A2(pi0609), .ZN(new_n13445_));
  NOR2_X1    g10545(.A1(new_n13428_), .A2(new_n13445_), .ZN(new_n13446_));
  NAND3_X1   g10546(.A1(new_n13427_), .A2(new_n13426_), .A3(new_n11903_), .ZN(new_n13447_));
  NAND2_X1   g10547(.A1(new_n13437_), .A2(pi0609), .ZN(new_n13448_));
  NOR4_X1    g10548(.A1(new_n13441_), .A2(new_n11903_), .A3(new_n13413_), .A4(new_n11914_), .ZN(new_n13449_));
  AOI21_X1   g10549(.A1(new_n13010_), .A2(new_n13409_), .B(new_n13449_), .ZN(new_n13450_));
  NAND3_X1   g10550(.A1(new_n13448_), .A2(pi0660), .A3(new_n11912_), .ZN(new_n13451_));
  INV_X1     g10551(.I(new_n13451_), .ZN(new_n13452_));
  AOI22_X1   g10552(.A1(new_n13446_), .A2(new_n13439_), .B1(new_n13447_), .B2(new_n13452_), .ZN(new_n13453_));
  NOR3_X1    g10553(.A1(new_n13453_), .A2(new_n11870_), .A3(new_n13430_), .ZN(new_n13454_));
  OAI21_X1   g10554(.A1(new_n13453_), .A2(new_n11870_), .B(new_n13430_), .ZN(new_n13455_));
  INV_X1     g10555(.I(new_n13455_), .ZN(new_n13456_));
  NOR3_X1    g10556(.A1(new_n13456_), .A2(pi0781), .A3(new_n13454_), .ZN(new_n13457_));
  INV_X1     g10557(.I(new_n13457_), .ZN(new_n13458_));
  NOR2_X1    g10558(.A1(new_n13456_), .A2(new_n13454_), .ZN(new_n13459_));
  NAND2_X1   g10559(.A1(new_n13437_), .A2(new_n11938_), .ZN(new_n13460_));
  OAI21_X1   g10560(.A1(new_n11938_), .A2(new_n13409_), .B(new_n13460_), .ZN(new_n13461_));
  AOI21_X1   g10561(.A1(new_n13461_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n13462_));
  NOR2_X1    g10562(.A1(new_n13409_), .A2(new_n11924_), .ZN(new_n13463_));
  NOR2_X1    g10563(.A1(new_n13417_), .A2(new_n11914_), .ZN(new_n13464_));
  NOR3_X1    g10564(.A1(new_n13464_), .A2(pi0785), .A3(new_n13463_), .ZN(new_n13465_));
  OAI21_X1   g10565(.A1(new_n13450_), .A2(new_n11912_), .B(new_n13443_), .ZN(new_n13466_));
  AND3_X2    g10566(.A1(new_n13466_), .A2(new_n13465_), .A3(pi0785), .Z(new_n13467_));
  AOI21_X1   g10567(.A1(new_n13466_), .A2(pi0785), .B(new_n13465_), .ZN(new_n13468_));
  NOR3_X1    g10568(.A1(new_n13467_), .A2(new_n13468_), .A3(new_n11934_), .ZN(new_n13469_));
  NOR2_X1    g10569(.A1(new_n13409_), .A2(new_n11934_), .ZN(new_n13470_));
  NOR4_X1    g10570(.A1(new_n13469_), .A2(new_n11949_), .A3(pi1154), .A4(new_n13470_), .ZN(new_n13471_));
  NOR3_X1    g10571(.A1(new_n13471_), .A2(new_n11934_), .A3(new_n13462_), .ZN(new_n13472_));
  INV_X1     g10572(.I(new_n13454_), .ZN(new_n13473_));
  NAND3_X1   g10573(.A1(new_n13473_), .A2(new_n11934_), .A3(new_n13455_), .ZN(new_n13474_));
  INV_X1     g10574(.I(new_n13461_), .ZN(new_n13475_));
  NOR2_X1    g10575(.A1(new_n13475_), .A2(new_n11934_), .ZN(new_n13476_));
  INV_X1     g10576(.I(new_n13469_), .ZN(new_n13477_));
  AOI21_X1   g10577(.A1(new_n13409_), .A2(new_n11934_), .B(pi1154), .ZN(new_n13478_));
  AOI21_X1   g10578(.A1(new_n13477_), .A2(new_n13478_), .B(pi0627), .ZN(new_n13479_));
  NOR3_X1    g10579(.A1(new_n13479_), .A2(pi1154), .A3(new_n13476_), .ZN(new_n13480_));
  AOI22_X1   g10580(.A1(new_n13474_), .A2(new_n13480_), .B1(new_n13459_), .B2(new_n13472_), .ZN(new_n13481_));
  NOR3_X1    g10581(.A1(new_n13481_), .A2(new_n11969_), .A3(new_n13458_), .ZN(new_n13482_));
  NAND3_X1   g10582(.A1(new_n13473_), .A2(new_n13472_), .A3(new_n13455_), .ZN(new_n13483_));
  NOR3_X1    g10583(.A1(new_n13456_), .A2(pi0618), .A3(new_n13454_), .ZN(new_n13484_));
  INV_X1     g10584(.I(new_n13480_), .ZN(new_n13485_));
  OAI21_X1   g10585(.A1(new_n13484_), .A2(new_n13485_), .B(new_n13483_), .ZN(new_n13486_));
  AOI21_X1   g10586(.A1(new_n13486_), .A2(pi0781), .B(new_n13457_), .ZN(new_n13487_));
  NOR3_X1    g10587(.A1(new_n13482_), .A2(new_n13487_), .A3(pi0789), .ZN(new_n13488_));
  INV_X1     g10588(.I(new_n13488_), .ZN(new_n13489_));
  NOR2_X1    g10589(.A1(new_n13482_), .A2(new_n13487_), .ZN(new_n13490_));
  NOR2_X1    g10590(.A1(new_n13467_), .A2(new_n13468_), .ZN(new_n13491_));
  NAND3_X1   g10591(.A1(new_n13409_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n13492_));
  MUX2_X1    g10592(.I0(new_n13492_), .I1(new_n13491_), .S(new_n11969_), .Z(new_n13493_));
  NAND2_X1   g10593(.A1(new_n13493_), .A2(pi0619), .ZN(new_n13494_));
  AOI21_X1   g10594(.A1(new_n13408_), .A2(pi0619), .B(pi1159), .ZN(new_n13495_));
  AND3_X2    g10595(.A1(new_n13494_), .A2(pi0648), .A3(new_n13495_), .Z(new_n13496_));
  NOR2_X1    g10596(.A1(new_n13408_), .A2(new_n11961_), .ZN(new_n13497_));
  AOI21_X1   g10597(.A1(new_n13475_), .A2(new_n11961_), .B(new_n13497_), .ZN(new_n13498_));
  NOR3_X1    g10598(.A1(new_n13496_), .A2(new_n11967_), .A3(pi1159), .ZN(new_n13499_));
  NAND3_X1   g10599(.A1(new_n13486_), .A2(pi0781), .A3(new_n13457_), .ZN(new_n13500_));
  OAI21_X1   g10600(.A1(new_n13481_), .A2(new_n11969_), .B(new_n13458_), .ZN(new_n13501_));
  NAND3_X1   g10601(.A1(new_n13501_), .A2(new_n13500_), .A3(new_n11967_), .ZN(new_n13502_));
  AOI21_X1   g10602(.A1(new_n13409_), .A2(new_n11967_), .B(pi1159), .ZN(new_n13503_));
  NAND2_X1   g10603(.A1(new_n13494_), .A2(new_n13503_), .ZN(new_n13504_));
  NAND2_X1   g10604(.A1(new_n13504_), .A2(new_n11966_), .ZN(new_n13505_));
  AOI21_X1   g10605(.A1(new_n13498_), .A2(pi0619), .B(pi1159), .ZN(new_n13506_));
  NAND2_X1   g10606(.A1(new_n13505_), .A2(new_n13506_), .ZN(new_n13507_));
  INV_X1     g10607(.I(new_n13507_), .ZN(new_n13508_));
  AOI22_X1   g10608(.A1(new_n13502_), .A2(new_n13508_), .B1(new_n13490_), .B2(new_n13499_), .ZN(new_n13509_));
  NOR3_X1    g10609(.A1(new_n13509_), .A2(new_n11985_), .A3(new_n13489_), .ZN(new_n13510_));
  NAND3_X1   g10610(.A1(new_n13501_), .A2(new_n13500_), .A3(new_n13499_), .ZN(new_n13511_));
  NOR3_X1    g10611(.A1(new_n13482_), .A2(new_n13487_), .A3(pi0619), .ZN(new_n13512_));
  OAI21_X1   g10612(.A1(new_n13512_), .A2(new_n13507_), .B(new_n13511_), .ZN(new_n13513_));
  AOI21_X1   g10613(.A1(new_n13513_), .A2(pi0789), .B(new_n13488_), .ZN(new_n13514_));
  NOR2_X1    g10614(.A1(new_n13510_), .A2(new_n13514_), .ZN(new_n13515_));
  INV_X1     g10615(.I(new_n13515_), .ZN(new_n13516_));
  NAND3_X1   g10616(.A1(new_n13513_), .A2(pi0789), .A3(new_n13488_), .ZN(new_n13517_));
  OAI21_X1   g10617(.A1(new_n13509_), .A2(new_n11985_), .B(new_n13489_), .ZN(new_n13518_));
  NOR2_X1    g10618(.A1(new_n13409_), .A2(new_n12014_), .ZN(new_n13519_));
  AOI21_X1   g10619(.A1(new_n13498_), .A2(new_n12014_), .B(new_n13519_), .ZN(new_n13520_));
  NOR2_X1    g10620(.A1(new_n11989_), .A2(pi0626), .ZN(new_n13521_));
  INV_X1     g10621(.I(new_n13521_), .ZN(new_n13522_));
  AOI21_X1   g10622(.A1(new_n13518_), .A2(new_n13517_), .B(new_n13522_), .ZN(new_n13523_));
  NOR2_X1    g10623(.A1(new_n11994_), .A2(pi0641), .ZN(new_n13524_));
  INV_X1     g10624(.I(new_n13524_), .ZN(new_n13525_));
  AOI21_X1   g10625(.A1(new_n13518_), .A2(new_n13517_), .B(new_n13525_), .ZN(new_n13526_));
  NAND3_X1   g10626(.A1(new_n13409_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n13527_));
  MUX2_X1    g10627(.I0(new_n13527_), .I1(new_n13493_), .S(new_n11985_), .Z(new_n13528_));
  NAND2_X1   g10628(.A1(new_n13528_), .A2(pi0626), .ZN(new_n13529_));
  AOI21_X1   g10629(.A1(new_n13409_), .A2(new_n11994_), .B(pi1158), .ZN(new_n13530_));
  NAND2_X1   g10630(.A1(new_n13529_), .A2(new_n13530_), .ZN(new_n13531_));
  AOI21_X1   g10631(.A1(new_n13408_), .A2(pi0626), .B(pi1158), .ZN(new_n13532_));
  NAND2_X1   g10632(.A1(new_n13529_), .A2(new_n13532_), .ZN(new_n13533_));
  INV_X1     g10633(.I(new_n13533_), .ZN(new_n13534_));
  AOI22_X1   g10634(.A1(new_n13534_), .A2(new_n12018_), .B1(new_n13095_), .B2(new_n13531_), .ZN(new_n13535_));
  INV_X1     g10635(.I(new_n13535_), .ZN(new_n13536_));
  NOR3_X1    g10636(.A1(new_n13523_), .A2(new_n13526_), .A3(new_n13536_), .ZN(new_n13537_));
  NOR3_X1    g10637(.A1(new_n13537_), .A2(new_n11986_), .A3(new_n13516_), .ZN(new_n13538_));
  AOI21_X1   g10638(.A1(new_n13537_), .A2(pi0788), .B(new_n13515_), .ZN(new_n13539_));
  NOR2_X1    g10639(.A1(new_n13538_), .A2(new_n13539_), .ZN(new_n13540_));
  NAND2_X1   g10640(.A1(new_n13528_), .A2(new_n11986_), .ZN(new_n13541_));
  AOI21_X1   g10641(.A1(new_n13534_), .A2(new_n13531_), .B(new_n11986_), .ZN(new_n13542_));
  XNOR2_X1   g10642(.A1(new_n13542_), .A2(new_n13541_), .ZN(new_n13543_));
  OAI21_X1   g10643(.A1(new_n13543_), .A2(pi0628), .B(pi1156), .ZN(new_n13544_));
  NOR2_X1    g10644(.A1(new_n13408_), .A2(new_n13114_), .ZN(new_n13545_));
  AOI21_X1   g10645(.A1(new_n13520_), .A2(new_n13114_), .B(new_n13545_), .ZN(new_n13546_));
  NOR3_X1    g10646(.A1(new_n13409_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n13547_));
  NOR2_X1    g10647(.A1(new_n13547_), .A2(new_n12030_), .ZN(new_n13548_));
  NOR2_X1    g10648(.A1(new_n13548_), .A2(new_n12031_), .ZN(new_n13549_));
  NAND2_X1   g10649(.A1(new_n13544_), .A2(new_n13549_), .ZN(new_n13550_));
  INV_X1     g10650(.I(new_n13550_), .ZN(new_n13551_));
  NOR2_X1    g10651(.A1(new_n13543_), .A2(new_n12031_), .ZN(new_n13552_));
  NOR2_X1    g10652(.A1(new_n12030_), .A2(pi0628), .ZN(new_n13553_));
  OAI21_X1   g10653(.A1(new_n13552_), .A2(pi1156), .B(new_n13553_), .ZN(new_n13554_));
  INV_X1     g10654(.I(new_n13554_), .ZN(new_n13555_));
  OAI22_X1   g10655(.A1(new_n13538_), .A2(new_n13539_), .B1(new_n13551_), .B2(new_n13555_), .ZN(new_n13556_));
  MUX2_X1    g10656(.I0(new_n13556_), .I1(new_n13540_), .S(new_n11868_), .Z(new_n13557_));
  OAI21_X1   g10657(.A1(new_n13510_), .A2(new_n13514_), .B(new_n13521_), .ZN(new_n13558_));
  OAI21_X1   g10658(.A1(new_n13510_), .A2(new_n13514_), .B(new_n13524_), .ZN(new_n13559_));
  NAND3_X1   g10659(.A1(new_n13558_), .A2(new_n13559_), .A3(new_n13535_), .ZN(new_n13560_));
  NAND3_X1   g10660(.A1(new_n13560_), .A2(pi0788), .A3(new_n13515_), .ZN(new_n13561_));
  OAI21_X1   g10661(.A1(new_n13560_), .A2(new_n11986_), .B(new_n13516_), .ZN(new_n13562_));
  AOI22_X1   g10662(.A1(new_n13562_), .A2(new_n13561_), .B1(new_n13550_), .B2(new_n13554_), .ZN(new_n13563_));
  NAND3_X1   g10663(.A1(new_n13563_), .A2(pi0792), .A3(new_n13540_), .ZN(new_n13564_));
  NAND2_X1   g10664(.A1(new_n13562_), .A2(new_n13561_), .ZN(new_n13565_));
  OAI21_X1   g10665(.A1(new_n13563_), .A2(new_n11868_), .B(new_n13565_), .ZN(new_n13566_));
  NOR2_X1    g10666(.A1(new_n13408_), .A2(new_n12054_), .ZN(new_n13567_));
  AOI21_X1   g10667(.A1(new_n13543_), .A2(new_n12054_), .B(new_n13567_), .ZN(new_n13568_));
  AOI21_X1   g10668(.A1(new_n13568_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n13569_));
  NOR4_X1    g10669(.A1(new_n13546_), .A2(new_n12031_), .A3(pi1156), .A4(new_n13408_), .ZN(new_n13570_));
  NOR2_X1    g10670(.A1(new_n13570_), .A2(new_n13547_), .ZN(new_n13571_));
  MUX2_X1    g10671(.I0(new_n13571_), .I1(new_n13546_), .S(new_n11868_), .Z(new_n13572_));
  NAND2_X1   g10672(.A1(new_n13572_), .A2(pi0647), .ZN(new_n13573_));
  INV_X1     g10673(.I(new_n13573_), .ZN(new_n13574_));
  NOR2_X1    g10674(.A1(new_n13409_), .A2(new_n12061_), .ZN(new_n13575_));
  NOR4_X1    g10675(.A1(new_n13574_), .A2(new_n12060_), .A3(pi1157), .A4(new_n13575_), .ZN(new_n13576_));
  NOR3_X1    g10676(.A1(new_n13569_), .A2(new_n12061_), .A3(new_n13576_), .ZN(new_n13577_));
  NAND3_X1   g10677(.A1(new_n13566_), .A2(new_n13564_), .A3(new_n13577_), .ZN(new_n13578_));
  NOR3_X1    g10678(.A1(new_n13556_), .A2(new_n11868_), .A3(new_n13565_), .ZN(new_n13579_));
  AOI21_X1   g10679(.A1(new_n13556_), .A2(pi0792), .B(new_n13540_), .ZN(new_n13580_));
  NOR3_X1    g10680(.A1(new_n13579_), .A2(new_n13580_), .A3(pi0647), .ZN(new_n13581_));
  AOI21_X1   g10681(.A1(new_n13409_), .A2(new_n12061_), .B(pi1157), .ZN(new_n13582_));
  NAND2_X1   g10682(.A1(new_n13573_), .A2(new_n13582_), .ZN(new_n13583_));
  NAND2_X1   g10683(.A1(new_n13583_), .A2(new_n12060_), .ZN(new_n13584_));
  AOI21_X1   g10684(.A1(new_n13568_), .A2(pi0647), .B(pi1157), .ZN(new_n13585_));
  AND2_X2    g10685(.A1(new_n13585_), .A2(new_n13584_), .Z(new_n13586_));
  INV_X1     g10686(.I(new_n13586_), .ZN(new_n13587_));
  OAI21_X1   g10687(.A1(new_n13581_), .A2(new_n13587_), .B(new_n13578_), .ZN(new_n13588_));
  MUX2_X1    g10688(.I0(new_n13588_), .I1(new_n13557_), .S(new_n12048_), .Z(new_n13589_));
  NAND2_X1   g10689(.A1(new_n13572_), .A2(new_n12048_), .ZN(new_n13590_));
  NOR3_X1    g10690(.A1(new_n13408_), .A2(pi0647), .A3(pi1157), .ZN(new_n13591_));
  NOR2_X1    g10691(.A1(new_n13591_), .A2(new_n12048_), .ZN(new_n13592_));
  XNOR2_X1   g10692(.A1(new_n13590_), .A2(new_n13592_), .ZN(new_n13593_));
  NOR2_X1    g10693(.A1(new_n13409_), .A2(new_n12092_), .ZN(new_n13594_));
  AOI21_X1   g10694(.A1(new_n13568_), .A2(new_n12092_), .B(new_n13594_), .ZN(new_n13595_));
  INV_X1     g10695(.I(new_n13595_), .ZN(new_n13596_));
  NOR2_X1    g10696(.A1(pi0644), .A2(pi0715), .ZN(new_n13597_));
  AOI21_X1   g10697(.A1(new_n13596_), .A2(new_n13597_), .B(new_n13169_), .ZN(new_n13598_));
  OAI21_X1   g10698(.A1(new_n12082_), .A2(new_n13593_), .B(new_n13598_), .ZN(new_n13599_));
  AOI21_X1   g10699(.A1(new_n13589_), .A2(new_n12082_), .B(new_n13599_), .ZN(new_n13600_));
  INV_X1     g10700(.I(new_n13557_), .ZN(new_n13601_));
  NAND3_X1   g10701(.A1(new_n13566_), .A2(new_n13564_), .A3(new_n12061_), .ZN(new_n13602_));
  AOI22_X1   g10702(.A1(new_n13602_), .A2(new_n13586_), .B1(new_n13557_), .B2(new_n13577_), .ZN(new_n13603_));
  MUX2_X1    g10703(.I0(new_n13603_), .I1(new_n13601_), .S(new_n12048_), .Z(new_n13604_));
  INV_X1     g10704(.I(new_n13593_), .ZN(new_n13605_));
  NAND3_X1   g10705(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n13606_));
  OAI21_X1   g10706(.A1(new_n13595_), .A2(new_n13606_), .B(new_n13179_), .ZN(new_n13607_));
  NOR2_X1    g10707(.A1(new_n13607_), .A2(new_n13605_), .ZN(new_n13608_));
  OAI21_X1   g10708(.A1(new_n13604_), .A2(new_n12082_), .B(new_n13608_), .ZN(new_n13609_));
  NOR2_X1    g10709(.A1(new_n13600_), .A2(new_n13609_), .ZN(new_n13610_));
  NAND2_X1   g10710(.A1(po1038), .A2(new_n11716_), .ZN(new_n13611_));
  AOI21_X1   g10711(.A1(new_n13611_), .A2(new_n13184_), .B(po1038), .ZN(new_n13612_));
  OAI21_X1   g10712(.A1(new_n13589_), .A2(pi0790), .B(new_n13612_), .ZN(new_n13613_));
  OAI21_X1   g10713(.A1(new_n13610_), .A2(new_n13613_), .B(new_n13325_), .ZN(po0298));
  NOR2_X1    g10714(.A1(new_n2925_), .A2(new_n5460_), .ZN(new_n13615_));
  INV_X1     g10715(.I(pi0743), .ZN(new_n13616_));
  NOR2_X1    g10716(.A1(new_n11877_), .A2(new_n13616_), .ZN(new_n13617_));
  INV_X1     g10717(.I(new_n13617_), .ZN(new_n13618_));
  NOR3_X1    g10718(.A1(new_n13618_), .A2(pi0609), .A3(new_n11914_), .ZN(new_n13619_));
  NOR3_X1    g10719(.A1(new_n13619_), .A2(pi1155), .A3(new_n13615_), .ZN(new_n13620_));
  NOR2_X1    g10720(.A1(new_n11903_), .A2(pi1155), .ZN(new_n13621_));
  INV_X1     g10721(.I(new_n13615_), .ZN(new_n13622_));
  NOR2_X1    g10722(.A1(new_n13618_), .A2(new_n11914_), .ZN(new_n13623_));
  NAND3_X1   g10723(.A1(new_n13623_), .A2(new_n13621_), .A3(new_n13622_), .ZN(new_n13624_));
  NAND3_X1   g10724(.A1(new_n13620_), .A2(new_n13624_), .A3(pi0785), .ZN(new_n13625_));
  OAI21_X1   g10725(.A1(new_n13623_), .A2(new_n13615_), .B(new_n11870_), .ZN(new_n13626_));
  NAND2_X1   g10726(.A1(new_n13625_), .A2(new_n13626_), .ZN(new_n13627_));
  INV_X1     g10727(.I(new_n13627_), .ZN(new_n13628_));
  NAND2_X1   g10728(.A1(new_n13628_), .A2(new_n11969_), .ZN(new_n13629_));
  NAND3_X1   g10729(.A1(new_n13622_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n13630_));
  NAND2_X1   g10730(.A1(new_n13630_), .A2(pi0781), .ZN(new_n13631_));
  XOR2_X1    g10731(.A1(new_n13629_), .A2(new_n13631_), .Z(new_n13632_));
  NAND2_X1   g10732(.A1(new_n13632_), .A2(pi0619), .ZN(new_n13633_));
  INV_X1     g10733(.I(new_n13633_), .ZN(new_n13634_));
  NOR2_X1    g10734(.A1(new_n13622_), .A2(new_n11967_), .ZN(new_n13635_));
  NOR2_X1    g10735(.A1(new_n13435_), .A2(new_n11891_), .ZN(new_n13636_));
  INV_X1     g10736(.I(new_n13636_), .ZN(new_n13637_));
  INV_X1     g10737(.I(pi0735), .ZN(new_n13638_));
  NOR2_X1    g10738(.A1(new_n11894_), .A2(new_n13638_), .ZN(new_n13639_));
  AOI21_X1   g10739(.A1(new_n13639_), .A2(new_n13637_), .B(new_n13615_), .ZN(new_n13640_));
  NOR2_X1    g10740(.A1(new_n13640_), .A2(new_n13024_), .ZN(new_n13641_));
  AOI21_X1   g10741(.A1(new_n13641_), .A2(new_n11961_), .B(new_n13615_), .ZN(new_n13642_));
  INV_X1     g10742(.I(new_n13642_), .ZN(new_n13643_));
  INV_X1     g10743(.I(new_n12118_), .ZN(new_n13644_));
  NOR2_X1    g10744(.A1(new_n13644_), .A2(new_n13638_), .ZN(new_n13645_));
  NOR3_X1    g10745(.A1(new_n13645_), .A2(new_n13615_), .A3(new_n13617_), .ZN(new_n13646_));
  NOR2_X1    g10746(.A1(new_n13646_), .A2(pi0778), .ZN(new_n13647_));
  NOR2_X1    g10747(.A1(new_n13644_), .A2(new_n12970_), .ZN(new_n13648_));
  INV_X1     g10748(.I(new_n13648_), .ZN(new_n13649_));
  NOR2_X1    g10749(.A1(new_n13649_), .A2(new_n13638_), .ZN(new_n13650_));
  INV_X1     g10750(.I(new_n13650_), .ZN(new_n13651_));
  INV_X1     g10751(.I(new_n13639_), .ZN(new_n13652_));
  OAI21_X1   g10752(.A1(pi0625), .A2(pi1153), .B(new_n13652_), .ZN(new_n13653_));
  NAND4_X1   g10753(.A1(new_n13653_), .A2(pi0608), .A3(pi1153), .A4(new_n13622_), .ZN(new_n13654_));
  AOI21_X1   g10754(.A1(new_n13651_), .A2(new_n13618_), .B(new_n13654_), .ZN(new_n13655_));
  INV_X1     g10755(.I(new_n13655_), .ZN(new_n13656_));
  INV_X1     g10756(.I(pi0608), .ZN(new_n13657_));
  AOI21_X1   g10757(.A1(new_n13651_), .A2(new_n13646_), .B(pi1153), .ZN(new_n13658_));
  INV_X1     g10758(.I(new_n13434_), .ZN(new_n13659_));
  NOR3_X1    g10759(.A1(new_n13652_), .A2(new_n13659_), .A3(new_n13615_), .ZN(new_n13660_));
  OAI21_X1   g10760(.A1(new_n13658_), .A2(new_n13660_), .B(new_n13657_), .ZN(new_n13661_));
  AOI21_X1   g10761(.A1(new_n13661_), .A2(new_n13656_), .B(new_n11891_), .ZN(new_n13662_));
  NOR2_X1    g10762(.A1(new_n13662_), .A2(new_n13647_), .ZN(new_n13663_));
  INV_X1     g10763(.I(new_n13663_), .ZN(new_n13664_));
  NAND2_X1   g10764(.A1(new_n13664_), .A2(new_n11870_), .ZN(new_n13665_));
  XOR2_X1    g10765(.A1(new_n13663_), .A2(new_n13640_), .Z(new_n13666_));
  NOR2_X1    g10766(.A1(new_n13666_), .A2(new_n11903_), .ZN(new_n13667_));
  XOR2_X1    g10767(.A1(new_n13667_), .A2(new_n13664_), .Z(new_n13668_));
  NAND2_X1   g10768(.A1(new_n13624_), .A2(new_n11923_), .ZN(new_n13669_));
  AOI21_X1   g10769(.A1(new_n13668_), .A2(new_n11912_), .B(new_n13669_), .ZN(new_n13670_));
  NOR3_X1    g10770(.A1(new_n13619_), .A2(pi1155), .A3(new_n13615_), .ZN(new_n13671_));
  NOR2_X1    g10771(.A1(new_n13671_), .A2(pi0660), .ZN(new_n13672_));
  OAI21_X1   g10772(.A1(new_n13670_), .A2(new_n13672_), .B(pi0785), .ZN(new_n13673_));
  NAND2_X1   g10773(.A1(new_n13673_), .A2(new_n13665_), .ZN(new_n13674_));
  AOI21_X1   g10774(.A1(new_n13622_), .A2(new_n11934_), .B(pi1154), .ZN(new_n13675_));
  OAI21_X1   g10775(.A1(new_n13627_), .A2(new_n11934_), .B(new_n13675_), .ZN(new_n13676_));
  NOR2_X1    g10776(.A1(new_n13641_), .A2(new_n13615_), .ZN(new_n13677_));
  XNOR2_X1   g10777(.A1(new_n13674_), .A2(new_n13677_), .ZN(new_n13678_));
  NOR2_X1    g10778(.A1(new_n13678_), .A2(new_n11934_), .ZN(new_n13679_));
  XOR2_X1    g10779(.A1(new_n13679_), .A2(new_n13674_), .Z(new_n13680_));
  NAND2_X1   g10780(.A1(new_n13680_), .A2(new_n11950_), .ZN(new_n13681_));
  NAND3_X1   g10781(.A1(new_n13681_), .A2(new_n11949_), .A3(new_n13676_), .ZN(new_n13682_));
  NOR2_X1    g10782(.A1(new_n13627_), .A2(new_n11934_), .ZN(new_n13683_));
  NOR2_X1    g10783(.A1(new_n13622_), .A2(new_n11934_), .ZN(new_n13684_));
  NOR3_X1    g10784(.A1(new_n13683_), .A2(pi1154), .A3(new_n13684_), .ZN(new_n13685_));
  NOR2_X1    g10785(.A1(new_n13685_), .A2(pi0627), .ZN(new_n13686_));
  INV_X1     g10786(.I(new_n13686_), .ZN(new_n13687_));
  AOI21_X1   g10787(.A1(new_n13682_), .A2(new_n13687_), .B(new_n11969_), .ZN(new_n13688_));
  AOI21_X1   g10788(.A1(new_n11969_), .A2(new_n13674_), .B(new_n13688_), .ZN(new_n13689_));
  NOR4_X1    g10789(.A1(new_n13634_), .A2(new_n11966_), .A3(pi1159), .A4(new_n13635_), .ZN(new_n13691_));
  INV_X1     g10790(.I(new_n13691_), .ZN(new_n13692_));
  MUX2_X1    g10791(.I0(new_n13689_), .I1(new_n13643_), .S(pi0619), .Z(new_n13693_));
  NOR2_X1    g10792(.A1(new_n13693_), .A2(pi1159), .ZN(new_n13694_));
  OAI21_X1   g10793(.A1(new_n13615_), .A2(pi0619), .B(new_n11869_), .ZN(new_n13695_));
  OAI21_X1   g10794(.A1(new_n13634_), .A2(new_n13695_), .B(new_n11966_), .ZN(new_n13696_));
  OAI21_X1   g10795(.A1(new_n13694_), .A2(new_n13696_), .B(new_n13692_), .ZN(new_n13697_));
  AOI21_X1   g10796(.A1(new_n13689_), .A2(new_n11998_), .B(pi0789), .ZN(new_n13698_));
  INV_X1     g10797(.I(new_n13632_), .ZN(new_n13699_));
  NOR3_X1    g10798(.A1(new_n13615_), .A2(pi0619), .A3(pi1159), .ZN(new_n13700_));
  MUX2_X1    g10799(.I0(new_n13700_), .I1(new_n13699_), .S(new_n11985_), .Z(new_n13701_));
  MUX2_X1    g10800(.I0(new_n13701_), .I1(new_n13615_), .S(new_n12003_), .Z(new_n13702_));
  NAND4_X1   g10801(.A1(new_n13643_), .A2(new_n12014_), .A3(new_n12020_), .A4(new_n13615_), .ZN(new_n13703_));
  NAND2_X1   g10802(.A1(new_n13703_), .A2(pi0788), .ZN(new_n13704_));
  AOI21_X1   g10803(.A1(new_n13702_), .A2(new_n12002_), .B(new_n13704_), .ZN(new_n13705_));
  AOI21_X1   g10804(.A1(new_n13697_), .A2(new_n13698_), .B(new_n13705_), .ZN(new_n13706_));
  NAND2_X1   g10805(.A1(new_n13701_), .A2(new_n11986_), .ZN(new_n13707_));
  NAND2_X1   g10806(.A1(new_n13702_), .A2(pi0788), .ZN(new_n13708_));
  NAND2_X1   g10807(.A1(new_n13708_), .A2(new_n13707_), .ZN(new_n13709_));
  NAND3_X1   g10808(.A1(new_n13706_), .A2(new_n12031_), .A3(new_n13709_), .ZN(new_n13710_));
  INV_X1     g10809(.I(new_n13709_), .ZN(new_n13711_));
  OAI21_X1   g10810(.A1(new_n13706_), .A2(pi0628), .B(new_n13711_), .ZN(new_n13712_));
  INV_X1     g10811(.I(new_n12032_), .ZN(new_n13713_));
  INV_X1     g10812(.I(new_n11961_), .ZN(new_n13714_));
  NOR2_X1    g10813(.A1(new_n13024_), .A2(new_n13714_), .ZN(new_n13715_));
  INV_X1     g10814(.I(new_n13715_), .ZN(new_n13716_));
  NOR2_X1    g10815(.A1(new_n13713_), .A2(new_n13716_), .ZN(new_n13717_));
  NOR2_X1    g10816(.A1(new_n13640_), .A2(new_n13717_), .ZN(new_n13718_));
  INV_X1     g10817(.I(new_n13718_), .ZN(new_n13719_));
  OAI21_X1   g10818(.A1(new_n13719_), .A2(pi0628), .B(new_n13622_), .ZN(new_n13720_));
  NAND2_X1   g10819(.A1(new_n13720_), .A2(new_n12026_), .ZN(new_n13721_));
  NAND2_X1   g10820(.A1(new_n13721_), .A2(pi0629), .ZN(new_n13722_));
  NOR2_X1    g10821(.A1(new_n13615_), .A2(pi1156), .ZN(new_n13723_));
  OAI21_X1   g10822(.A1(new_n13719_), .A2(new_n12031_), .B(new_n13723_), .ZN(new_n13724_));
  AND4_X2    g10823(.A1(new_n12030_), .A2(new_n13722_), .A3(new_n12026_), .A4(new_n13724_), .Z(new_n13725_));
  NAND3_X1   g10824(.A1(new_n13712_), .A2(new_n13710_), .A3(new_n13725_), .ZN(new_n13726_));
  MUX2_X1    g10825(.I0(new_n13726_), .I1(new_n13706_), .S(new_n11868_), .Z(new_n13727_));
  INV_X1     g10826(.I(new_n13727_), .ZN(new_n13728_));
  NOR2_X1    g10827(.A1(new_n12054_), .A2(new_n13615_), .ZN(new_n13729_));
  AOI21_X1   g10828(.A1(new_n13711_), .A2(new_n12054_), .B(new_n13729_), .ZN(new_n13730_));
  INV_X1     g10829(.I(new_n13730_), .ZN(new_n13731_));
  NAND3_X1   g10830(.A1(new_n13727_), .A2(new_n12061_), .A3(new_n13731_), .ZN(new_n13732_));
  OAI21_X1   g10831(.A1(new_n13727_), .A2(pi0647), .B(new_n13730_), .ZN(new_n13733_));
  NOR2_X1    g10832(.A1(new_n13719_), .A2(new_n12066_), .ZN(new_n13734_));
  INV_X1     g10833(.I(new_n13734_), .ZN(new_n13735_));
  NOR2_X1    g10834(.A1(new_n12061_), .A2(pi1157), .ZN(new_n13736_));
  INV_X1     g10835(.I(new_n13736_), .ZN(new_n13737_));
  NOR3_X1    g10836(.A1(new_n13735_), .A2(new_n13615_), .A3(new_n13737_), .ZN(new_n13738_));
  NOR3_X1    g10837(.A1(new_n13738_), .A2(pi0630), .A3(pi1157), .ZN(new_n13739_));
  NAND3_X1   g10838(.A1(new_n13733_), .A2(new_n13732_), .A3(new_n13739_), .ZN(new_n13740_));
  NOR2_X1    g10839(.A1(new_n13735_), .A2(pi0647), .ZN(new_n13741_));
  INV_X1     g10840(.I(new_n13741_), .ZN(new_n13742_));
  INV_X1     g10841(.I(new_n12089_), .ZN(new_n13743_));
  NOR2_X1    g10842(.A1(new_n13615_), .A2(new_n13743_), .ZN(new_n13744_));
  AOI21_X1   g10843(.A1(new_n13742_), .A2(new_n13744_), .B(new_n12048_), .ZN(new_n13745_));
  AOI22_X1   g10844(.A1(new_n13740_), .A2(new_n13745_), .B1(new_n12048_), .B2(new_n13728_), .ZN(new_n13746_));
  NOR2_X1    g10845(.A1(new_n12049_), .A2(pi0647), .ZN(new_n13747_));
  OAI21_X1   g10846(.A1(new_n13736_), .A2(new_n13747_), .B(pi0787), .ZN(new_n13748_));
  AOI21_X1   g10847(.A1(new_n13734_), .A2(new_n13748_), .B(new_n13615_), .ZN(new_n13749_));
  INV_X1     g10848(.I(new_n13749_), .ZN(new_n13750_));
  XOR2_X1    g10849(.A1(new_n13746_), .A2(new_n13750_), .Z(new_n13751_));
  NAND2_X1   g10850(.A1(new_n13751_), .A2(pi0644), .ZN(new_n13752_));
  XOR2_X1    g10851(.A1(new_n13752_), .A2(new_n13746_), .Z(new_n13753_));
  NAND2_X1   g10852(.A1(new_n13753_), .A2(new_n12099_), .ZN(new_n13754_));
  NOR2_X1    g10853(.A1(new_n12092_), .A2(new_n13622_), .ZN(new_n13755_));
  AOI21_X1   g10854(.A1(new_n13730_), .A2(new_n12092_), .B(new_n13755_), .ZN(new_n13756_));
  AOI21_X1   g10855(.A1(new_n13615_), .A2(pi0644), .B(new_n12096_), .ZN(new_n13757_));
  AOI21_X1   g10856(.A1(new_n13756_), .A2(new_n13757_), .B(pi1160), .ZN(new_n13758_));
  XOR2_X1    g10857(.A1(new_n13752_), .A2(new_n13749_), .Z(new_n13759_));
  AOI21_X1   g10858(.A1(new_n12082_), .A2(new_n13622_), .B(new_n13756_), .ZN(new_n13760_));
  NOR4_X1    g10859(.A1(new_n13730_), .A2(pi0644), .A3(new_n12091_), .A4(new_n13622_), .ZN(new_n13761_));
  NOR3_X1    g10860(.A1(new_n13760_), .A2(pi0715), .A3(new_n13761_), .ZN(new_n13762_));
  OAI21_X1   g10861(.A1(new_n13759_), .A2(new_n12099_), .B(new_n13762_), .ZN(new_n13763_));
  AOI22_X1   g10862(.A1(new_n13763_), .A2(new_n12081_), .B1(new_n13754_), .B2(new_n13758_), .ZN(new_n13764_));
  MUX2_X1    g10863(.I0(new_n13764_), .I1(new_n13746_), .S(new_n11867_), .Z(new_n13765_));
  OR2_X2     g10864(.A1(new_n13765_), .A2(new_n13184_), .Z(new_n13766_));
  NOR2_X1    g10865(.A1(new_n3231_), .A2(new_n5460_), .ZN(new_n13767_));
  NOR2_X1    g10866(.A1(new_n12110_), .A2(pi0142), .ZN(new_n13768_));
  AOI21_X1   g10867(.A1(new_n2490_), .A2(new_n13617_), .B(new_n13768_), .ZN(new_n13769_));
  NAND3_X1   g10868(.A1(new_n13769_), .A2(pi0735), .A3(new_n12115_), .ZN(new_n13770_));
  NAND2_X1   g10869(.A1(pi0039), .A2(pi0142), .ZN(new_n13771_));
  NAND3_X1   g10870(.A1(new_n3232_), .A2(pi0038), .A3(new_n13771_), .ZN(new_n13772_));
  AOI21_X1   g10871(.A1(new_n13770_), .A2(new_n3154_), .B(new_n13772_), .ZN(new_n13773_));
  AOI21_X1   g10872(.A1(new_n5460_), .A2(new_n12511_), .B(new_n12391_), .ZN(new_n13774_));
  NAND3_X1   g10873(.A1(new_n12391_), .A2(new_n5460_), .A3(new_n12481_), .ZN(new_n13775_));
  NAND2_X1   g10874(.A1(new_n13775_), .A2(new_n13616_), .ZN(new_n13777_));
  OAI21_X1   g10875(.A1(new_n13777_), .A2(new_n13774_), .B(pi0735), .ZN(new_n13778_));
  NAND3_X1   g10876(.A1(new_n12438_), .A2(pi0142), .A3(pi0743), .ZN(new_n13779_));
  NAND2_X1   g10877(.A1(new_n12264_), .A2(new_n12259_), .ZN(new_n13780_));
  NAND4_X1   g10878(.A1(new_n13780_), .A2(new_n12316_), .A3(pi0142), .A4(new_n13616_), .ZN(new_n13781_));
  NAND2_X1   g10879(.A1(new_n13779_), .A2(new_n13781_), .ZN(new_n13782_));
  NAND2_X1   g10880(.A1(new_n13782_), .A2(pi0735), .ZN(new_n13783_));
  NAND4_X1   g10881(.A1(new_n13783_), .A2(new_n2604_), .A3(new_n5141_), .A4(new_n13778_), .ZN(new_n13784_));
  NOR4_X1    g10882(.A1(new_n12812_), .A2(new_n12199_), .A3(pi0142), .A4(pi0743), .ZN(new_n13785_));
  NAND2_X1   g10883(.A1(new_n12767_), .A2(pi0142), .ZN(new_n13786_));
  AOI21_X1   g10884(.A1(new_n13616_), .A2(new_n13786_), .B(new_n13785_), .ZN(new_n13787_));
  NOR3_X1    g10885(.A1(new_n12429_), .A2(new_n5460_), .A3(new_n13616_), .ZN(new_n13788_));
  MUX2_X1    g10886(.I0(new_n12328_), .I1(new_n12203_), .S(new_n5460_), .Z(new_n13789_));
  AOI21_X1   g10887(.A1(new_n13789_), .A2(pi0743), .B(new_n13788_), .ZN(new_n13790_));
  NOR3_X1    g10888(.A1(new_n13790_), .A2(new_n13638_), .A3(new_n13787_), .ZN(new_n13791_));
  INV_X1     g10889(.I(new_n13787_), .ZN(new_n13792_));
  AOI21_X1   g10890(.A1(new_n13790_), .A2(pi0735), .B(new_n13792_), .ZN(new_n13793_));
  NOR3_X1    g10891(.A1(new_n13791_), .A2(new_n13793_), .A3(new_n5141_), .ZN(new_n13794_));
  INV_X1     g10892(.I(new_n13794_), .ZN(new_n13795_));
  INV_X1     g10893(.I(new_n12337_), .ZN(new_n13796_));
  AOI21_X1   g10894(.A1(new_n12234_), .A2(new_n5460_), .B(new_n13796_), .ZN(new_n13797_));
  NOR3_X1    g10895(.A1(new_n12234_), .A2(pi0142), .A3(new_n12337_), .ZN(new_n13798_));
  OAI21_X1   g10896(.A1(new_n13798_), .A2(new_n13797_), .B(pi0743), .ZN(new_n13799_));
  NAND3_X1   g10897(.A1(new_n12423_), .A2(pi0142), .A3(pi0743), .ZN(new_n13800_));
  AOI21_X1   g10898(.A1(new_n13799_), .A2(new_n13800_), .B(new_n13638_), .ZN(new_n13801_));
  NAND3_X1   g10899(.A1(new_n12879_), .A2(pi0142), .A3(new_n13616_), .ZN(new_n13802_));
  OR2_X2     g10900(.A1(new_n12674_), .A2(pi0142), .Z(new_n13803_));
  NAND2_X1   g10901(.A1(new_n12806_), .A2(pi0142), .ZN(new_n13804_));
  XOR2_X1    g10902(.A1(new_n13803_), .A2(new_n13804_), .Z(new_n13805_));
  NOR2_X1    g10903(.A1(new_n13805_), .A2(new_n13616_), .ZN(new_n13806_));
  XOR2_X1    g10904(.A1(new_n13806_), .A2(new_n13802_), .Z(new_n13807_));
  AOI21_X1   g10905(.A1(new_n13807_), .A2(new_n13638_), .B(new_n13801_), .ZN(new_n13808_));
  AOI21_X1   g10906(.A1(new_n13808_), .A2(new_n5141_), .B(new_n2614_), .ZN(new_n13809_));
  NAND2_X1   g10907(.A1(new_n13809_), .A2(new_n13795_), .ZN(new_n13810_));
  NOR2_X1    g10908(.A1(new_n12132_), .A2(new_n5460_), .ZN(new_n13811_));
  AOI21_X1   g10909(.A1(new_n12208_), .A2(pi0743), .B(new_n13811_), .ZN(new_n13812_));
  INV_X1     g10910(.I(new_n13812_), .ZN(new_n13813_));
  AOI21_X1   g10911(.A1(new_n13769_), .A2(new_n12115_), .B(new_n12340_), .ZN(new_n13814_));
  OAI21_X1   g10912(.A1(new_n5460_), .A2(new_n12132_), .B(new_n13814_), .ZN(new_n13815_));
  MUX2_X1    g10913(.I0(new_n13815_), .I1(new_n13813_), .S(new_n13638_), .Z(new_n13816_));
  AOI21_X1   g10914(.A1(new_n13816_), .A2(new_n2614_), .B(pi0223), .ZN(new_n13817_));
  NAND2_X1   g10915(.A1(new_n13810_), .A2(new_n13817_), .ZN(new_n13818_));
  AOI21_X1   g10916(.A1(new_n13818_), .A2(new_n13784_), .B(pi0299), .ZN(new_n13819_));
  NOR2_X1    g10917(.A1(new_n2587_), .A2(pi0039), .ZN(new_n13820_));
  NAND4_X1   g10918(.A1(new_n13783_), .A2(new_n2566_), .A3(new_n5094_), .A4(new_n13778_), .ZN(new_n13821_));
  INV_X1     g10919(.I(new_n13821_), .ZN(new_n13822_));
  OR3_X2     g10920(.A1(new_n13791_), .A2(new_n13793_), .A3(new_n5094_), .Z(new_n13823_));
  NAND2_X1   g10921(.A1(new_n13816_), .A2(new_n3284_), .ZN(new_n13824_));
  AOI21_X1   g10922(.A1(new_n13824_), .A2(new_n2566_), .B(new_n6445_), .ZN(new_n13825_));
  NAND2_X1   g10923(.A1(new_n13808_), .A2(new_n13825_), .ZN(new_n13826_));
  AOI21_X1   g10924(.A1(new_n13823_), .A2(new_n3285_), .B(new_n13826_), .ZN(new_n13827_));
  OAI21_X1   g10925(.A1(new_n13827_), .A2(new_n13822_), .B(new_n13820_), .ZN(new_n13828_));
  NOR2_X1    g10926(.A1(new_n12631_), .A2(new_n5095_), .ZN(new_n13829_));
  NAND2_X1   g10927(.A1(new_n12613_), .A2(pi0603), .ZN(new_n13830_));
  INV_X1     g10928(.I(new_n13830_), .ZN(new_n13831_));
  AOI21_X1   g10929(.A1(new_n12655_), .A2(pi0680), .B(new_n12652_), .ZN(new_n13832_));
  OAI21_X1   g10930(.A1(new_n13831_), .A2(new_n13832_), .B(new_n5460_), .ZN(new_n13833_));
  NOR2_X1    g10931(.A1(pi0142), .A2(pi0299), .ZN(new_n13834_));
  AND3_X2    g10932(.A1(new_n13833_), .A2(new_n13616_), .A3(new_n13834_), .Z(new_n13835_));
  NAND2_X1   g10933(.A1(new_n13835_), .A2(new_n13829_), .ZN(new_n13836_));
  OAI21_X1   g10934(.A1(new_n12627_), .A2(new_n5101_), .B(new_n12590_), .ZN(new_n13837_));
  NOR2_X1    g10935(.A1(new_n13837_), .A2(new_n5460_), .ZN(new_n13838_));
  OAI21_X1   g10936(.A1(pi0680), .A2(new_n12655_), .B(new_n13838_), .ZN(new_n13839_));
  NOR2_X1    g10937(.A1(new_n13831_), .A2(pi0142), .ZN(new_n13840_));
  INV_X1     g10938(.I(new_n13840_), .ZN(new_n13841_));
  AOI21_X1   g10939(.A1(pi0680), .A2(new_n12641_), .B(new_n13841_), .ZN(new_n13842_));
  AOI21_X1   g10940(.A1(new_n13842_), .A2(new_n13839_), .B(new_n13616_), .ZN(new_n13843_));
  NOR2_X1    g10941(.A1(new_n12625_), .A2(new_n5095_), .ZN(new_n13844_));
  AOI21_X1   g10942(.A1(new_n12648_), .A2(pi0680), .B(new_n12646_), .ZN(new_n13845_));
  NOR2_X1    g10943(.A1(new_n13845_), .A2(new_n12610_), .ZN(new_n13846_));
  NAND4_X1   g10944(.A1(new_n13844_), .A2(new_n5460_), .A3(new_n13616_), .A4(new_n13846_), .ZN(new_n13847_));
  INV_X1     g10945(.I(new_n13845_), .ZN(new_n13848_));
  NOR2_X1    g10946(.A1(new_n12606_), .A2(new_n12609_), .ZN(new_n13849_));
  AOI21_X1   g10947(.A1(new_n13849_), .A2(new_n5101_), .B(new_n12619_), .ZN(new_n13850_));
  NOR3_X1    g10948(.A1(new_n13850_), .A2(new_n5460_), .A3(new_n13848_), .ZN(new_n13851_));
  NOR2_X1    g10949(.A1(new_n12624_), .A2(new_n5095_), .ZN(new_n13852_));
  NAND2_X1   g10950(.A1(new_n13834_), .A2(pi0743), .ZN(new_n13853_));
  NOR4_X1    g10951(.A1(new_n13851_), .A2(new_n12610_), .A3(new_n13852_), .A4(new_n13853_), .ZN(new_n13854_));
  AOI22_X1   g10952(.A1(new_n13843_), .A2(new_n13836_), .B1(new_n13847_), .B2(new_n13854_), .ZN(new_n13855_));
  AOI21_X1   g10953(.A1(new_n12652_), .A2(pi0142), .B(pi0743), .ZN(new_n13856_));
  NOR4_X1    g10954(.A1(new_n13840_), .A2(new_n2587_), .A3(new_n13838_), .A4(new_n13856_), .ZN(new_n13857_));
  NAND2_X1   g10955(.A1(new_n13849_), .A2(pi0603), .ZN(new_n13858_));
  INV_X1     g10956(.I(new_n13850_), .ZN(new_n13859_));
  MUX2_X1    g10957(.I0(new_n13859_), .I1(new_n13858_), .S(new_n5460_), .Z(new_n13860_));
  NAND3_X1   g10958(.A1(new_n12646_), .A2(pi0142), .A3(new_n13616_), .ZN(new_n13861_));
  OAI21_X1   g10959(.A1(new_n13860_), .A2(new_n13616_), .B(new_n13861_), .ZN(new_n13862_));
  AOI21_X1   g10960(.A1(new_n13862_), .A2(new_n2587_), .B(new_n13857_), .ZN(new_n13863_));
  NOR3_X1    g10961(.A1(new_n13863_), .A2(new_n13855_), .A3(pi0735), .ZN(new_n13864_));
  INV_X1     g10962(.I(new_n13855_), .ZN(new_n13865_));
  AOI21_X1   g10963(.A1(new_n13863_), .A2(new_n13638_), .B(new_n13865_), .ZN(new_n13866_));
  NOR3_X1    g10964(.A1(new_n13866_), .A2(pi0039), .A3(new_n13864_), .ZN(new_n13867_));
  OAI21_X1   g10965(.A1(new_n13819_), .A2(new_n13828_), .B(new_n13867_), .ZN(new_n13868_));
  NAND2_X1   g10966(.A1(new_n13868_), .A2(new_n3172_), .ZN(new_n13869_));
  AOI21_X1   g10967(.A1(new_n13869_), .A2(new_n13773_), .B(new_n13767_), .ZN(new_n13870_));
  INV_X1     g10968(.I(new_n13773_), .ZN(new_n13871_));
  NAND3_X1   g10969(.A1(new_n13868_), .A2(new_n3172_), .A3(new_n13871_), .ZN(new_n13872_));
  NOR2_X1    g10970(.A1(new_n13767_), .A2(pi0625), .ZN(new_n13873_));
  NOR2_X1    g10971(.A1(new_n6445_), .A2(pi0215), .ZN(new_n13874_));
  NAND2_X1   g10972(.A1(new_n13806_), .A2(new_n13802_), .ZN(new_n13875_));
  NAND2_X1   g10973(.A1(new_n12879_), .A2(pi0142), .ZN(new_n13876_));
  NOR2_X1    g10974(.A1(new_n13876_), .A2(pi0743), .ZN(new_n13877_));
  INV_X1     g10975(.I(new_n13877_), .ZN(new_n13878_));
  NAND3_X1   g10976(.A1(new_n13875_), .A2(new_n5094_), .A3(new_n13878_), .ZN(new_n13879_));
  NOR2_X1    g10977(.A1(new_n13787_), .A2(new_n5094_), .ZN(new_n13880_));
  INV_X1     g10978(.I(new_n13880_), .ZN(new_n13881_));
  NAND4_X1   g10979(.A1(new_n13879_), .A2(new_n3284_), .A3(new_n13812_), .A4(new_n13881_), .ZN(new_n13882_));
  AOI22_X1   g10980(.A1(new_n13879_), .A2(new_n13881_), .B1(new_n3284_), .B2(new_n13813_), .ZN(new_n13883_));
  INV_X1     g10981(.I(new_n13883_), .ZN(new_n13884_));
  AOI21_X1   g10982(.A1(new_n13884_), .A2(new_n13882_), .B(pi0215), .ZN(new_n13885_));
  NOR2_X1    g10983(.A1(new_n13885_), .A2(new_n13874_), .ZN(new_n13886_));
  AOI22_X1   g10984(.A1(new_n13875_), .A2(new_n13878_), .B1(new_n6460_), .B2(new_n13792_), .ZN(new_n13887_));
  NAND4_X1   g10985(.A1(new_n13875_), .A2(new_n6460_), .A3(new_n13787_), .A4(new_n13878_), .ZN(new_n13888_));
  NOR3_X1    g10986(.A1(new_n2614_), .A2(pi0223), .A3(pi0299), .ZN(new_n13889_));
  NAND2_X1   g10987(.A1(new_n13888_), .A2(new_n13889_), .ZN(new_n13890_));
  NOR2_X1    g10988(.A1(new_n13890_), .A2(new_n13887_), .ZN(new_n13891_));
  OAI21_X1   g10989(.A1(new_n13891_), .A2(new_n3154_), .B(pi0299), .ZN(new_n13892_));
  INV_X1     g10990(.I(new_n13863_), .ZN(new_n13893_));
  AOI21_X1   g10991(.A1(new_n13893_), .A2(new_n3154_), .B(pi0038), .ZN(new_n13894_));
  OAI21_X1   g10992(.A1(new_n13886_), .A2(new_n13892_), .B(new_n13894_), .ZN(new_n13895_));
  AOI21_X1   g10993(.A1(new_n13769_), .A2(new_n3154_), .B(new_n13772_), .ZN(new_n13896_));
  AOI21_X1   g10994(.A1(new_n13895_), .A2(new_n13896_), .B(new_n13767_), .ZN(new_n13897_));
  OAI21_X1   g10995(.A1(new_n13897_), .A2(pi0625), .B(new_n11893_), .ZN(new_n13898_));
  AOI21_X1   g10996(.A1(new_n13872_), .A2(new_n13873_), .B(new_n13898_), .ZN(new_n13899_));
  NOR2_X1    g10997(.A1(pi0608), .A2(pi0625), .ZN(new_n13900_));
  INV_X1     g10998(.I(new_n13767_), .ZN(new_n13901_));
  INV_X1     g10999(.I(new_n13873_), .ZN(new_n13902_));
  INV_X1     g11000(.I(new_n13875_), .ZN(new_n13903_));
  OAI22_X1   g11001(.A1(new_n13903_), .A2(new_n13877_), .B1(new_n5141_), .B2(new_n13787_), .ZN(new_n13904_));
  NAND3_X1   g11002(.A1(new_n13904_), .A2(new_n13888_), .A3(new_n13889_), .ZN(new_n13905_));
  AOI21_X1   g11003(.A1(new_n13905_), .A2(pi0039), .B(new_n2587_), .ZN(new_n13906_));
  OAI21_X1   g11004(.A1(new_n13874_), .A2(new_n13885_), .B(new_n13906_), .ZN(new_n13907_));
  INV_X1     g11005(.I(new_n13896_), .ZN(new_n13908_));
  AOI21_X1   g11006(.A1(new_n13907_), .A2(new_n13894_), .B(new_n13908_), .ZN(new_n13909_));
  OAI21_X1   g11007(.A1(new_n13909_), .A2(new_n13902_), .B(pi1153), .ZN(new_n13910_));
  NOR2_X1    g11008(.A1(new_n13876_), .A2(pi0735), .ZN(new_n13911_));
  NAND2_X1   g11009(.A1(new_n12945_), .A2(new_n5460_), .ZN(new_n13912_));
  INV_X1     g11010(.I(new_n13912_), .ZN(new_n13913_));
  AND2_X2    g11011(.A1(new_n12923_), .A2(pi0142), .Z(new_n13914_));
  XOR2_X1    g11012(.A1(new_n13914_), .A2(new_n13913_), .Z(new_n13915_));
  NOR3_X1    g11013(.A1(new_n13915_), .A2(new_n13638_), .A3(new_n13911_), .ZN(new_n13916_));
  NOR2_X1    g11014(.A1(new_n13876_), .A2(pi0735), .ZN(new_n13917_));
  NOR2_X1    g11015(.A1(new_n13786_), .A2(pi0735), .ZN(new_n13918_));
  NAND2_X1   g11016(.A1(new_n12947_), .A2(new_n5460_), .ZN(new_n13919_));
  OAI21_X1   g11017(.A1(new_n12926_), .A2(new_n5460_), .B(new_n13919_), .ZN(new_n13920_));
  NAND2_X1   g11018(.A1(new_n13920_), .A2(pi0735), .ZN(new_n13921_));
  XNOR2_X1   g11019(.A1(new_n13921_), .A2(new_n13918_), .ZN(new_n13922_));
  OAI22_X1   g11020(.A1(new_n13916_), .A2(new_n13917_), .B1(new_n5094_), .B2(new_n13922_), .ZN(new_n13923_));
  INV_X1     g11021(.I(new_n13922_), .ZN(new_n13924_));
  NOR4_X1    g11022(.A1(new_n13916_), .A2(new_n5094_), .A3(new_n13917_), .A4(new_n13924_), .ZN(new_n13925_));
  NOR2_X1    g11023(.A1(new_n13925_), .A2(new_n3284_), .ZN(new_n13926_));
  NOR2_X1    g11024(.A1(new_n12886_), .A2(new_n5460_), .ZN(new_n13927_));
  INV_X1     g11025(.I(new_n13927_), .ZN(new_n13928_));
  INV_X1     g11026(.I(new_n12914_), .ZN(new_n13929_));
  INV_X1     g11027(.I(new_n12254_), .ZN(new_n13930_));
  NOR4_X1    g11028(.A1(new_n12938_), .A2(new_n13930_), .A3(pi0142), .A4(new_n5095_), .ZN(new_n13931_));
  AOI22_X1   g11029(.A1(new_n13929_), .A2(pi0142), .B1(new_n12258_), .B2(new_n13931_), .ZN(new_n13932_));
  MUX2_X1    g11030(.I0(new_n13932_), .I1(new_n13928_), .S(new_n13638_), .Z(new_n13933_));
  NAND2_X1   g11031(.A1(new_n12786_), .A2(pi0142), .ZN(new_n13934_));
  NOR2_X1    g11032(.A1(new_n12915_), .A2(new_n5460_), .ZN(new_n13935_));
  NOR2_X1    g11033(.A1(new_n13935_), .A2(new_n13931_), .ZN(new_n13936_));
  MUX2_X1    g11034(.I0(new_n13936_), .I1(new_n13934_), .S(new_n13638_), .Z(new_n13937_));
  INV_X1     g11035(.I(new_n13937_), .ZN(new_n13938_));
  OAI21_X1   g11036(.A1(new_n13933_), .A2(new_n13938_), .B(new_n5094_), .ZN(new_n13939_));
  AOI21_X1   g11037(.A1(new_n12681_), .A2(new_n13639_), .B(new_n13811_), .ZN(new_n13940_));
  NAND2_X1   g11038(.A1(new_n13940_), .A2(new_n3284_), .ZN(new_n13941_));
  AOI21_X1   g11039(.A1(new_n13941_), .A2(new_n2566_), .B(pi0299), .ZN(new_n13942_));
  OAI21_X1   g11040(.A1(new_n13939_), .A2(new_n2566_), .B(new_n13942_), .ZN(new_n13943_));
  AOI21_X1   g11041(.A1(new_n13926_), .A2(new_n13923_), .B(new_n13943_), .ZN(new_n13944_));
  INV_X1     g11042(.I(new_n13911_), .ZN(new_n13945_));
  XOR2_X1    g11043(.A1(new_n13914_), .A2(new_n13912_), .Z(new_n13946_));
  NAND3_X1   g11044(.A1(new_n13946_), .A2(pi0735), .A3(new_n13945_), .ZN(new_n13947_));
  INV_X1     g11045(.I(new_n13917_), .ZN(new_n13948_));
  AOI22_X1   g11046(.A1(new_n13947_), .A2(new_n13948_), .B1(new_n6460_), .B2(new_n13924_), .ZN(new_n13949_));
  NAND4_X1   g11047(.A1(new_n13947_), .A2(new_n6460_), .A3(new_n13948_), .A4(new_n13922_), .ZN(new_n13950_));
  NOR3_X1    g11048(.A1(new_n2614_), .A2(pi0223), .A3(pi0299), .ZN(new_n13952_));
  NAND2_X1   g11049(.A1(new_n13950_), .A2(new_n13952_), .ZN(new_n13953_));
  OAI21_X1   g11050(.A1(new_n12852_), .A2(pi0735), .B(new_n5460_), .ZN(new_n13954_));
  NAND2_X1   g11051(.A1(new_n13954_), .A2(new_n3154_), .ZN(new_n13955_));
  OAI21_X1   g11052(.A1(new_n2491_), .A2(new_n13652_), .B(new_n3154_), .ZN(new_n13956_));
  NOR2_X1    g11053(.A1(new_n13768_), .A2(new_n13956_), .ZN(new_n13957_));
  OAI21_X1   g11054(.A1(new_n13957_), .A2(new_n13772_), .B(pi0039), .ZN(new_n13958_));
  AOI21_X1   g11055(.A1(new_n13955_), .A2(new_n3172_), .B(new_n13958_), .ZN(new_n13959_));
  OAI21_X1   g11056(.A1(new_n13953_), .A2(new_n13949_), .B(new_n13959_), .ZN(new_n13960_));
  OAI21_X1   g11057(.A1(new_n13944_), .A2(new_n13960_), .B(new_n13901_), .ZN(new_n13961_));
  AOI21_X1   g11058(.A1(new_n13927_), .A2(new_n13934_), .B(new_n6445_), .ZN(new_n13962_));
  NAND2_X1   g11059(.A1(new_n13962_), .A2(pi0215), .ZN(new_n13963_));
  INV_X1     g11060(.I(new_n13811_), .ZN(new_n13964_));
  AOI21_X1   g11061(.A1(new_n12767_), .A2(new_n6445_), .B(pi0142), .ZN(new_n13965_));
  OAI21_X1   g11062(.A1(new_n12759_), .A2(new_n6445_), .B(new_n13965_), .ZN(new_n13966_));
  MUX2_X1    g11063(.I0(new_n13966_), .I1(new_n13964_), .S(new_n3284_), .Z(new_n13967_));
  OAI21_X1   g11064(.A1(new_n13967_), .A2(pi0215), .B(new_n13963_), .ZN(new_n13968_));
  NAND3_X1   g11065(.A1(new_n13968_), .A2(pi0039), .A3(pi0299), .ZN(new_n13969_));
  NAND4_X1   g11066(.A1(new_n12893_), .A2(pi0039), .A3(new_n5460_), .A4(new_n12697_), .ZN(new_n13970_));
  AOI21_X1   g11067(.A1(new_n13969_), .A2(new_n13970_), .B(new_n10843_), .ZN(new_n13971_));
  AOI21_X1   g11068(.A1(new_n12899_), .A2(pi0038), .B(new_n3232_), .ZN(new_n13972_));
  NOR2_X1    g11069(.A1(new_n13972_), .A2(new_n5460_), .ZN(new_n13973_));
  NOR2_X1    g11070(.A1(new_n13971_), .A2(new_n13973_), .ZN(new_n13974_));
  AOI21_X1   g11071(.A1(new_n13974_), .A2(pi0625), .B(pi1153), .ZN(new_n13975_));
  OAI21_X1   g11072(.A1(new_n13961_), .A2(pi0625), .B(new_n13975_), .ZN(new_n13976_));
  NAND4_X1   g11073(.A1(new_n13910_), .A2(new_n13900_), .A3(new_n13976_), .A4(new_n13901_), .ZN(new_n13977_));
  INV_X1     g11074(.I(new_n13974_), .ZN(new_n13978_));
  AOI21_X1   g11075(.A1(new_n13978_), .A2(pi1153), .B(pi0625), .ZN(new_n13979_));
  AND2_X2    g11076(.A1(new_n13961_), .A2(new_n13979_), .Z(new_n13980_));
  NOR2_X1    g11077(.A1(new_n13980_), .A2(pi0608), .ZN(new_n13981_));
  OAI21_X1   g11078(.A1(new_n13977_), .A2(new_n13872_), .B(new_n13981_), .ZN(new_n13982_));
  NOR2_X1    g11079(.A1(new_n13982_), .A2(new_n13899_), .ZN(new_n13983_));
  NOR3_X1    g11080(.A1(new_n13983_), .A2(new_n11891_), .A3(new_n13870_), .ZN(new_n13984_));
  INV_X1     g11081(.I(new_n13870_), .ZN(new_n13985_));
  AOI21_X1   g11082(.A1(new_n13983_), .A2(pi0778), .B(new_n13985_), .ZN(new_n13986_));
  NOR2_X1    g11083(.A1(new_n13984_), .A2(new_n13986_), .ZN(new_n13987_));
  NAND2_X1   g11084(.A1(new_n13987_), .A2(new_n11870_), .ZN(new_n13988_));
  NAND2_X1   g11085(.A1(new_n13961_), .A2(new_n11891_), .ZN(new_n13989_));
  INV_X1     g11086(.I(new_n13976_), .ZN(new_n13990_));
  OAI21_X1   g11087(.A1(new_n13990_), .A2(new_n13980_), .B(pi0778), .ZN(new_n13991_));
  NOR2_X1    g11088(.A1(new_n13991_), .A2(new_n13989_), .ZN(new_n13992_));
  NAND2_X1   g11089(.A1(new_n13991_), .A2(new_n13989_), .ZN(new_n13993_));
  INV_X1     g11090(.I(new_n13993_), .ZN(new_n13994_));
  OAI21_X1   g11091(.A1(new_n13994_), .A2(new_n13992_), .B(new_n11903_), .ZN(new_n13995_));
  NOR2_X1    g11092(.A1(new_n13974_), .A2(new_n12996_), .ZN(new_n13996_));
  INV_X1     g11093(.I(new_n13996_), .ZN(new_n13997_));
  INV_X1     g11094(.I(new_n13874_), .ZN(new_n13998_));
  INV_X1     g11095(.I(new_n13882_), .ZN(new_n13999_));
  OAI21_X1   g11096(.A1(new_n13999_), .A2(new_n13883_), .B(new_n2566_), .ZN(new_n14000_));
  AOI21_X1   g11097(.A1(new_n13998_), .A2(new_n14000_), .B(new_n13892_), .ZN(new_n14001_));
  INV_X1     g11098(.I(new_n13894_), .ZN(new_n14002_));
  OAI21_X1   g11099(.A1(new_n14001_), .A2(new_n14002_), .B(new_n13896_), .ZN(new_n14003_));
  NAND2_X1   g11100(.A1(new_n14003_), .A2(new_n13901_), .ZN(new_n14004_));
  NAND3_X1   g11101(.A1(new_n14004_), .A2(new_n11903_), .A3(new_n11924_), .ZN(new_n14005_));
  AOI21_X1   g11102(.A1(new_n14005_), .A2(new_n13997_), .B(pi1155), .ZN(new_n14006_));
  OAI21_X1   g11103(.A1(new_n14006_), .A2(new_n11923_), .B(pi0609), .ZN(new_n14007_));
  AOI21_X1   g11104(.A1(new_n13995_), .A2(pi1155), .B(new_n14007_), .ZN(new_n14008_));
  INV_X1     g11105(.I(new_n13784_), .ZN(new_n14009_));
  INV_X1     g11106(.I(new_n13817_), .ZN(new_n14010_));
  AOI21_X1   g11107(.A1(new_n13809_), .A2(new_n13795_), .B(new_n14010_), .ZN(new_n14011_));
  OAI21_X1   g11108(.A1(new_n14011_), .A2(new_n14009_), .B(new_n2587_), .ZN(new_n14012_));
  INV_X1     g11109(.I(new_n13828_), .ZN(new_n14013_));
  INV_X1     g11110(.I(new_n13864_), .ZN(new_n14014_));
  OAI21_X1   g11111(.A1(new_n13893_), .A2(pi0735), .B(new_n13855_), .ZN(new_n14015_));
  NAND3_X1   g11112(.A1(new_n14014_), .A2(new_n14015_), .A3(new_n3154_), .ZN(new_n14016_));
  AOI21_X1   g11113(.A1(new_n14013_), .A2(new_n14012_), .B(new_n14016_), .ZN(new_n14017_));
  NOR3_X1    g11114(.A1(new_n14017_), .A2(pi0038), .A3(new_n13773_), .ZN(new_n14018_));
  AOI21_X1   g11115(.A1(new_n14004_), .A2(new_n12970_), .B(pi1153), .ZN(new_n14019_));
  OAI21_X1   g11116(.A1(new_n14018_), .A2(new_n13902_), .B(new_n14019_), .ZN(new_n14020_));
  NOR2_X1    g11117(.A1(new_n14017_), .A2(pi0038), .ZN(new_n14021_));
  NAND2_X1   g11118(.A1(new_n13901_), .A2(new_n13900_), .ZN(new_n14022_));
  NOR2_X1    g11119(.A1(new_n13990_), .A2(new_n14022_), .ZN(new_n14023_));
  NAND4_X1   g11120(.A1(new_n14023_), .A2(new_n14021_), .A3(new_n13871_), .A4(new_n13910_), .ZN(new_n14024_));
  NAND3_X1   g11121(.A1(new_n14024_), .A2(new_n14020_), .A3(new_n13981_), .ZN(new_n14025_));
  NAND3_X1   g11122(.A1(new_n14025_), .A2(pi0778), .A3(new_n13985_), .ZN(new_n14026_));
  OAI21_X1   g11123(.A1(new_n14025_), .A2(new_n11891_), .B(new_n13870_), .ZN(new_n14027_));
  NAND3_X1   g11124(.A1(new_n14027_), .A2(new_n14026_), .A3(new_n11903_), .ZN(new_n14028_));
  INV_X1     g11125(.I(new_n13992_), .ZN(new_n14029_));
  NAND2_X1   g11126(.A1(new_n14029_), .A2(new_n13993_), .ZN(new_n14030_));
  NOR2_X1    g11127(.A1(new_n13974_), .A2(new_n11915_), .ZN(new_n14031_));
  NAND2_X1   g11128(.A1(new_n14004_), .A2(new_n11924_), .ZN(new_n14032_));
  NOR2_X1    g11129(.A1(new_n14032_), .A2(new_n11903_), .ZN(new_n14033_));
  NOR2_X1    g11130(.A1(new_n11923_), .A2(pi1155), .ZN(new_n14034_));
  INV_X1     g11131(.I(new_n14034_), .ZN(new_n14035_));
  AOI21_X1   g11132(.A1(new_n14030_), .A2(pi0609), .B(new_n14035_), .ZN(new_n14036_));
  AOI22_X1   g11133(.A1(new_n14028_), .A2(new_n14036_), .B1(new_n13987_), .B2(new_n14008_), .ZN(new_n14037_));
  NOR3_X1    g11134(.A1(new_n14037_), .A2(new_n11870_), .A3(new_n13988_), .ZN(new_n14038_));
  MUX2_X1    g11135(.I0(new_n14025_), .I1(new_n13870_), .S(new_n11891_), .Z(new_n14039_));
  NOR2_X1    g11136(.A1(new_n14039_), .A2(pi0785), .ZN(new_n14040_));
  AOI21_X1   g11137(.A1(new_n14029_), .A2(new_n13993_), .B(pi0609), .ZN(new_n14041_));
  INV_X1     g11138(.I(new_n14007_), .ZN(new_n14042_));
  OAI21_X1   g11139(.A1(new_n14041_), .A2(new_n11912_), .B(new_n14042_), .ZN(new_n14043_));
  NOR3_X1    g11140(.A1(new_n13984_), .A2(new_n13986_), .A3(pi0609), .ZN(new_n14044_));
  NOR2_X1    g11141(.A1(new_n13994_), .A2(new_n13992_), .ZN(new_n14045_));
  OAI21_X1   g11142(.A1(new_n14045_), .A2(new_n11903_), .B(new_n14034_), .ZN(new_n14046_));
  OAI22_X1   g11143(.A1(new_n14044_), .A2(new_n14046_), .B1(new_n14039_), .B2(new_n14043_), .ZN(new_n14047_));
  AOI21_X1   g11144(.A1(new_n14047_), .A2(pi0785), .B(new_n14040_), .ZN(new_n14048_));
  NOR3_X1    g11145(.A1(new_n14038_), .A2(new_n14048_), .A3(pi0781), .ZN(new_n14049_));
  INV_X1     g11146(.I(new_n14049_), .ZN(new_n14050_));
  MUX2_X1    g11147(.I0(new_n14047_), .I1(new_n13987_), .S(new_n11870_), .Z(new_n14051_));
  OAI21_X1   g11148(.A1(new_n11924_), .A2(new_n13974_), .B(new_n14032_), .ZN(new_n14052_));
  INV_X1     g11149(.I(new_n14006_), .ZN(new_n14053_));
  OAI21_X1   g11150(.A1(new_n14033_), .A2(new_n14031_), .B(pi1155), .ZN(new_n14054_));
  NAND2_X1   g11151(.A1(new_n14054_), .A2(new_n14053_), .ZN(new_n14055_));
  MUX2_X1    g11152(.I0(new_n14055_), .I1(new_n14052_), .S(new_n11870_), .Z(new_n14056_));
  OAI21_X1   g11153(.A1(new_n13978_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n14057_));
  AOI21_X1   g11154(.A1(new_n14056_), .A2(pi0618), .B(new_n14057_), .ZN(new_n14058_));
  NOR2_X1    g11155(.A1(new_n13974_), .A2(new_n11938_), .ZN(new_n14059_));
  AOI21_X1   g11156(.A1(new_n14045_), .A2(new_n11938_), .B(new_n14059_), .ZN(new_n14060_));
  NAND2_X1   g11157(.A1(new_n11950_), .A2(pi0618), .ZN(new_n14061_));
  AOI21_X1   g11158(.A1(new_n14058_), .A2(pi0627), .B(new_n14061_), .ZN(new_n14062_));
  NAND3_X1   g11159(.A1(new_n14047_), .A2(pi0785), .A3(new_n14040_), .ZN(new_n14063_));
  OAI21_X1   g11160(.A1(new_n14037_), .A2(new_n11870_), .B(new_n13988_), .ZN(new_n14064_));
  NAND3_X1   g11161(.A1(new_n14064_), .A2(new_n14063_), .A3(new_n11934_), .ZN(new_n14065_));
  NAND2_X1   g11162(.A1(new_n14056_), .A2(pi0618), .ZN(new_n14066_));
  AOI21_X1   g11163(.A1(new_n13978_), .A2(new_n11934_), .B(pi1154), .ZN(new_n14067_));
  NAND2_X1   g11164(.A1(new_n14066_), .A2(new_n14067_), .ZN(new_n14068_));
  AOI21_X1   g11165(.A1(new_n14060_), .A2(pi0618), .B(pi1154), .ZN(new_n14069_));
  INV_X1     g11166(.I(new_n14069_), .ZN(new_n14070_));
  AOI21_X1   g11167(.A1(new_n14068_), .A2(new_n11949_), .B(new_n14070_), .ZN(new_n14071_));
  AOI22_X1   g11168(.A1(new_n14065_), .A2(new_n14071_), .B1(new_n14051_), .B2(new_n14062_), .ZN(new_n14072_));
  NOR3_X1    g11169(.A1(new_n14072_), .A2(new_n11969_), .A3(new_n14050_), .ZN(new_n14073_));
  NAND3_X1   g11170(.A1(new_n14064_), .A2(new_n14063_), .A3(new_n14062_), .ZN(new_n14074_));
  NOR3_X1    g11171(.A1(new_n14038_), .A2(new_n14048_), .A3(pi0618), .ZN(new_n14075_));
  INV_X1     g11172(.I(new_n14071_), .ZN(new_n14076_));
  OAI21_X1   g11173(.A1(new_n14075_), .A2(new_n14076_), .B(new_n14074_), .ZN(new_n14077_));
  AOI21_X1   g11174(.A1(new_n14077_), .A2(pi0781), .B(new_n14049_), .ZN(new_n14078_));
  NOR3_X1    g11175(.A1(new_n14078_), .A2(new_n14073_), .A3(pi0789), .ZN(new_n14079_));
  INV_X1     g11176(.I(new_n14079_), .ZN(new_n14080_));
  MUX2_X1    g11177(.I0(new_n14077_), .I1(new_n14051_), .S(new_n11969_), .Z(new_n14081_));
  NOR3_X1    g11178(.A1(new_n13974_), .A2(pi0618), .A3(pi1154), .ZN(new_n14082_));
  INV_X1     g11179(.I(new_n14082_), .ZN(new_n14083_));
  MUX2_X1    g11180(.I0(new_n14083_), .I1(new_n14056_), .S(new_n11969_), .Z(new_n14084_));
  OAI21_X1   g11181(.A1(new_n13978_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n14085_));
  AOI21_X1   g11182(.A1(new_n14084_), .A2(pi0619), .B(new_n14085_), .ZN(new_n14086_));
  NOR2_X1    g11183(.A1(new_n13978_), .A2(new_n11961_), .ZN(new_n14087_));
  AOI21_X1   g11184(.A1(new_n14060_), .A2(new_n11961_), .B(new_n14087_), .ZN(new_n14088_));
  NAND2_X1   g11185(.A1(new_n11869_), .A2(pi0619), .ZN(new_n14089_));
  AOI21_X1   g11186(.A1(new_n14086_), .A2(pi0648), .B(new_n14089_), .ZN(new_n14090_));
  NAND3_X1   g11187(.A1(new_n14077_), .A2(pi0781), .A3(new_n14049_), .ZN(new_n14091_));
  OAI21_X1   g11188(.A1(new_n14072_), .A2(new_n11969_), .B(new_n14050_), .ZN(new_n14092_));
  NAND3_X1   g11189(.A1(new_n14092_), .A2(new_n14091_), .A3(new_n11967_), .ZN(new_n14093_));
  AOI21_X1   g11190(.A1(new_n13978_), .A2(new_n11967_), .B(pi1159), .ZN(new_n14094_));
  INV_X1     g11191(.I(new_n14094_), .ZN(new_n14095_));
  AOI21_X1   g11192(.A1(new_n14084_), .A2(pi0619), .B(new_n14095_), .ZN(new_n14096_));
  OAI21_X1   g11193(.A1(new_n14088_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n14097_));
  INV_X1     g11194(.I(new_n14097_), .ZN(new_n14098_));
  OAI21_X1   g11195(.A1(new_n14096_), .A2(pi0648), .B(new_n14098_), .ZN(new_n14099_));
  INV_X1     g11196(.I(new_n14099_), .ZN(new_n14100_));
  AOI22_X1   g11197(.A1(new_n14093_), .A2(new_n14100_), .B1(new_n14081_), .B2(new_n14090_), .ZN(new_n14101_));
  NOR3_X1    g11198(.A1(new_n14101_), .A2(new_n11985_), .A3(new_n14080_), .ZN(new_n14102_));
  NAND3_X1   g11199(.A1(new_n14092_), .A2(new_n14091_), .A3(new_n14090_), .ZN(new_n14103_));
  NOR3_X1    g11200(.A1(new_n14078_), .A2(new_n14073_), .A3(pi0619), .ZN(new_n14104_));
  OAI21_X1   g11201(.A1(new_n14104_), .A2(new_n14099_), .B(new_n14103_), .ZN(new_n14105_));
  AOI21_X1   g11202(.A1(new_n14105_), .A2(pi0789), .B(new_n14079_), .ZN(new_n14106_));
  NOR2_X1    g11203(.A1(new_n14106_), .A2(new_n14102_), .ZN(new_n14107_));
  NAND3_X1   g11204(.A1(new_n14105_), .A2(pi0789), .A3(new_n14079_), .ZN(new_n14108_));
  OAI21_X1   g11205(.A1(new_n14101_), .A2(new_n11985_), .B(new_n14080_), .ZN(new_n14109_));
  NOR2_X1    g11206(.A1(new_n13974_), .A2(new_n12014_), .ZN(new_n14110_));
  AOI21_X1   g11207(.A1(new_n14088_), .A2(new_n12014_), .B(new_n14110_), .ZN(new_n14111_));
  NOR2_X1    g11208(.A1(new_n11989_), .A2(pi0626), .ZN(new_n14112_));
  INV_X1     g11209(.I(new_n14112_), .ZN(new_n14113_));
  AOI21_X1   g11210(.A1(new_n14109_), .A2(new_n14108_), .B(new_n14113_), .ZN(new_n14114_));
  NOR2_X1    g11211(.A1(new_n11994_), .A2(pi0641), .ZN(new_n14115_));
  INV_X1     g11212(.I(new_n14115_), .ZN(new_n14116_));
  AOI21_X1   g11213(.A1(new_n14109_), .A2(new_n14108_), .B(new_n14116_), .ZN(new_n14117_));
  AND2_X2    g11214(.A1(new_n14084_), .A2(new_n11985_), .Z(new_n14118_));
  INV_X1     g11215(.I(new_n14096_), .ZN(new_n14119_));
  AOI21_X1   g11216(.A1(new_n14119_), .A2(new_n14086_), .B(new_n11985_), .ZN(new_n14120_));
  XNOR2_X1   g11217(.A1(new_n14120_), .A2(new_n14118_), .ZN(new_n14121_));
  AOI21_X1   g11218(.A1(new_n13978_), .A2(new_n11994_), .B(pi1158), .ZN(new_n14122_));
  OAI21_X1   g11219(.A1(new_n14121_), .A2(new_n11994_), .B(new_n14122_), .ZN(new_n14123_));
  XOR2_X1    g11220(.A1(new_n14120_), .A2(new_n14118_), .Z(new_n14124_));
  AOI21_X1   g11221(.A1(new_n13974_), .A2(pi0626), .B(pi1158), .ZN(new_n14125_));
  INV_X1     g11222(.I(new_n14125_), .ZN(new_n14126_));
  AOI21_X1   g11223(.A1(new_n14124_), .A2(pi0626), .B(new_n14126_), .ZN(new_n14127_));
  AOI22_X1   g11224(.A1(new_n14123_), .A2(new_n13095_), .B1(new_n14127_), .B2(new_n12018_), .ZN(new_n14128_));
  INV_X1     g11225(.I(new_n14128_), .ZN(new_n14129_));
  NOR3_X1    g11226(.A1(new_n14114_), .A2(new_n14117_), .A3(new_n14129_), .ZN(new_n14130_));
  MUX2_X1    g11227(.I0(new_n14130_), .I1(new_n14107_), .S(new_n11986_), .Z(new_n14131_));
  INV_X1     g11228(.I(new_n14107_), .ZN(new_n14132_));
  NOR3_X1    g11229(.A1(new_n14130_), .A2(new_n11986_), .A3(new_n14132_), .ZN(new_n14133_));
  AOI21_X1   g11230(.A1(new_n14130_), .A2(pi0788), .B(new_n14107_), .ZN(new_n14134_));
  NOR3_X1    g11231(.A1(new_n13974_), .A2(pi0626), .A3(pi1158), .ZN(new_n14135_));
  NOR2_X1    g11232(.A1(new_n14135_), .A2(new_n11986_), .ZN(new_n14136_));
  NAND3_X1   g11233(.A1(new_n14124_), .A2(new_n11986_), .A3(new_n14136_), .ZN(new_n14137_));
  INV_X1     g11234(.I(new_n14136_), .ZN(new_n14138_));
  OAI21_X1   g11235(.A1(new_n14121_), .A2(pi0788), .B(new_n14138_), .ZN(new_n14139_));
  NAND2_X1   g11236(.A1(new_n14139_), .A2(new_n14137_), .ZN(new_n14140_));
  NAND2_X1   g11237(.A1(new_n14140_), .A2(new_n12031_), .ZN(new_n14141_));
  NOR2_X1    g11238(.A1(new_n14111_), .A2(new_n11992_), .ZN(new_n14142_));
  AOI21_X1   g11239(.A1(new_n11992_), .A2(new_n13978_), .B(new_n14142_), .ZN(new_n14143_));
  NOR3_X1    g11240(.A1(new_n13978_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n14144_));
  OAI21_X1   g11241(.A1(new_n14144_), .A2(new_n12030_), .B(pi0628), .ZN(new_n14145_));
  AOI21_X1   g11242(.A1(new_n14141_), .A2(pi1156), .B(new_n14145_), .ZN(new_n14146_));
  AOI21_X1   g11243(.A1(new_n14139_), .A2(new_n14137_), .B(new_n12031_), .ZN(new_n14147_));
  NOR2_X1    g11244(.A1(new_n12030_), .A2(pi0628), .ZN(new_n14148_));
  OAI21_X1   g11245(.A1(new_n14147_), .A2(pi1156), .B(new_n14148_), .ZN(new_n14149_));
  INV_X1     g11246(.I(new_n14149_), .ZN(new_n14150_));
  OAI22_X1   g11247(.A1(new_n14133_), .A2(new_n14134_), .B1(new_n14146_), .B2(new_n14150_), .ZN(new_n14151_));
  MUX2_X1    g11248(.I0(new_n14151_), .I1(new_n14131_), .S(new_n11868_), .Z(new_n14152_));
  INV_X1     g11249(.I(new_n14152_), .ZN(new_n14153_));
  NOR2_X1    g11250(.A1(new_n14140_), .A2(new_n12053_), .ZN(new_n14154_));
  AOI21_X1   g11251(.A1(new_n12053_), .A2(new_n13978_), .B(new_n14154_), .ZN(new_n14155_));
  AOI21_X1   g11252(.A1(new_n14155_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n14156_));
  NOR4_X1    g11253(.A1(new_n14143_), .A2(new_n12031_), .A3(pi1156), .A4(new_n13974_), .ZN(new_n14157_));
  NOR2_X1    g11254(.A1(new_n14157_), .A2(new_n14144_), .ZN(new_n14158_));
  MUX2_X1    g11255(.I0(new_n14158_), .I1(new_n14143_), .S(new_n11868_), .Z(new_n14159_));
  NAND2_X1   g11256(.A1(new_n14159_), .A2(pi0647), .ZN(new_n14160_));
  AOI21_X1   g11257(.A1(new_n13974_), .A2(pi0647), .B(pi1157), .ZN(new_n14161_));
  AND3_X2    g11258(.A1(new_n14160_), .A2(pi0630), .A3(new_n14161_), .Z(new_n14162_));
  NOR3_X1    g11259(.A1(new_n14156_), .A2(new_n12061_), .A3(new_n14162_), .ZN(new_n14163_));
  OAI21_X1   g11260(.A1(new_n14106_), .A2(new_n14102_), .B(new_n14112_), .ZN(new_n14164_));
  OAI21_X1   g11261(.A1(new_n14106_), .A2(new_n14102_), .B(new_n14115_), .ZN(new_n14165_));
  NAND3_X1   g11262(.A1(new_n14164_), .A2(new_n14165_), .A3(new_n14128_), .ZN(new_n14166_));
  NAND3_X1   g11263(.A1(new_n14166_), .A2(pi0788), .A3(new_n14107_), .ZN(new_n14167_));
  OAI21_X1   g11264(.A1(new_n14166_), .A2(new_n11986_), .B(new_n14132_), .ZN(new_n14168_));
  INV_X1     g11265(.I(new_n14146_), .ZN(new_n14169_));
  AOI21_X1   g11266(.A1(new_n14168_), .A2(new_n14167_), .B(new_n14169_), .ZN(new_n14170_));
  NAND3_X1   g11267(.A1(new_n14170_), .A2(pi0792), .A3(new_n14131_), .ZN(new_n14171_));
  NAND2_X1   g11268(.A1(new_n14168_), .A2(new_n14167_), .ZN(new_n14172_));
  AOI22_X1   g11269(.A1(new_n14168_), .A2(new_n14167_), .B1(new_n14169_), .B2(new_n14149_), .ZN(new_n14173_));
  OAI21_X1   g11270(.A1(new_n14173_), .A2(new_n11868_), .B(new_n14172_), .ZN(new_n14174_));
  NAND3_X1   g11271(.A1(new_n14174_), .A2(new_n14171_), .A3(new_n12061_), .ZN(new_n14175_));
  AOI21_X1   g11272(.A1(new_n13978_), .A2(new_n12061_), .B(pi1157), .ZN(new_n14176_));
  NAND2_X1   g11273(.A1(new_n14160_), .A2(new_n14176_), .ZN(new_n14177_));
  NAND2_X1   g11274(.A1(new_n14177_), .A2(new_n12060_), .ZN(new_n14178_));
  NAND2_X1   g11275(.A1(new_n14178_), .A2(new_n12049_), .ZN(new_n14179_));
  AOI21_X1   g11276(.A1(new_n14155_), .A2(pi0647), .B(new_n14179_), .ZN(new_n14180_));
  AOI22_X1   g11277(.A1(new_n14175_), .A2(new_n14180_), .B1(new_n14152_), .B2(new_n14163_), .ZN(new_n14181_));
  MUX2_X1    g11278(.I0(new_n14181_), .I1(new_n14153_), .S(new_n12048_), .Z(new_n14182_));
  NOR2_X1    g11279(.A1(new_n13978_), .A2(new_n12092_), .ZN(new_n14183_));
  AOI21_X1   g11280(.A1(new_n14155_), .A2(new_n12092_), .B(new_n14183_), .ZN(new_n14184_));
  NAND4_X1   g11281(.A1(new_n14184_), .A2(pi0644), .A3(new_n12099_), .A4(new_n13978_), .ZN(new_n14185_));
  NAND3_X1   g11282(.A1(new_n13978_), .A2(new_n12061_), .A3(new_n12049_), .ZN(new_n14186_));
  MUX2_X1    g11283(.I0(new_n14186_), .I1(new_n14159_), .S(new_n12048_), .Z(new_n14187_));
  OAI21_X1   g11284(.A1(new_n14187_), .A2(new_n12082_), .B(new_n12099_), .ZN(new_n14188_));
  AOI21_X1   g11285(.A1(new_n14185_), .A2(new_n12081_), .B(new_n14188_), .ZN(new_n14189_));
  OAI21_X1   g11286(.A1(new_n14182_), .A2(pi0644), .B(new_n14189_), .ZN(new_n14190_));
  NAND2_X1   g11287(.A1(new_n14152_), .A2(new_n12048_), .ZN(new_n14191_));
  OR3_X2     g11288(.A1(new_n14181_), .A2(new_n12048_), .A3(new_n14191_), .Z(new_n14192_));
  OAI21_X1   g11289(.A1(new_n14181_), .A2(new_n12048_), .B(new_n14191_), .ZN(new_n14193_));
  INV_X1     g11290(.I(new_n14184_), .ZN(new_n14194_));
  OAI21_X1   g11291(.A1(pi0644), .A2(new_n13974_), .B(new_n14194_), .ZN(new_n14195_));
  NAND3_X1   g11292(.A1(new_n14184_), .A2(new_n12082_), .A3(new_n13974_), .ZN(new_n14196_));
  NOR2_X1    g11293(.A1(new_n12081_), .A2(pi0715), .ZN(new_n14197_));
  NAND3_X1   g11294(.A1(new_n14195_), .A2(new_n14196_), .A3(new_n14197_), .ZN(new_n14198_));
  NOR2_X1    g11295(.A1(new_n12082_), .A2(pi0715), .ZN(new_n14199_));
  NAND4_X1   g11296(.A1(new_n14192_), .A2(new_n14193_), .A3(new_n14198_), .A4(new_n14199_), .ZN(new_n14200_));
  OAI21_X1   g11297(.A1(new_n14182_), .A2(new_n5223_), .B(new_n11867_), .ZN(new_n14201_));
  AOI21_X1   g11298(.A1(new_n14190_), .A2(new_n14200_), .B(new_n14201_), .ZN(new_n14202_));
  NAND2_X1   g11299(.A1(pi0057), .A2(pi0142), .ZN(new_n14203_));
  AOI21_X1   g11300(.A1(new_n14203_), .A2(new_n13184_), .B(pi0057), .ZN(new_n14204_));
  OAI21_X1   g11301(.A1(new_n5224_), .A2(pi0142), .B(new_n14204_), .ZN(new_n14205_));
  OAI21_X1   g11302(.A1(new_n14202_), .A2(new_n14205_), .B(new_n13766_), .ZN(po0299));
  NOR2_X1    g11303(.A1(new_n2925_), .A2(pi0143), .ZN(new_n14207_));
  NOR2_X1    g11304(.A1(new_n11877_), .A2(pi0774), .ZN(new_n14208_));
  NOR2_X1    g11305(.A1(new_n14208_), .A2(new_n14207_), .ZN(new_n14209_));
  INV_X1     g11306(.I(new_n14209_), .ZN(new_n14210_));
  AOI21_X1   g11307(.A1(new_n11886_), .A2(pi0687), .B(new_n14207_), .ZN(new_n14211_));
  NOR2_X1    g11308(.A1(new_n14211_), .A2(new_n11874_), .ZN(new_n14212_));
  NOR2_X1    g11309(.A1(new_n14210_), .A2(new_n14212_), .ZN(new_n14213_));
  NOR2_X1    g11310(.A1(new_n14213_), .A2(pi0778), .ZN(new_n14214_));
  NAND2_X1   g11311(.A1(new_n14212_), .A2(pi0625), .ZN(new_n14215_));
  INV_X1     g11312(.I(pi0687), .ZN(new_n14216_));
  NOR2_X1    g11313(.A1(new_n13201_), .A2(new_n14216_), .ZN(new_n14217_));
  NOR4_X1    g11314(.A1(new_n14208_), .A2(pi0608), .A3(new_n11893_), .A4(new_n14207_), .ZN(new_n14218_));
  OAI21_X1   g11315(.A1(new_n14210_), .A2(new_n14212_), .B(new_n14215_), .ZN(new_n14219_));
  NOR3_X1    g11316(.A1(new_n14207_), .A2(pi0608), .A3(pi1153), .ZN(new_n14220_));
  AOI22_X1   g11317(.A1(new_n14219_), .A2(new_n14220_), .B1(new_n14215_), .B2(new_n14218_), .ZN(new_n14221_));
  NOR2_X1    g11318(.A1(new_n14221_), .A2(new_n11891_), .ZN(new_n14222_));
  XOR2_X1    g11319(.A1(new_n14222_), .A2(new_n14214_), .Z(new_n14223_));
  INV_X1     g11320(.I(new_n14223_), .ZN(new_n14224_));
  NAND2_X1   g11321(.A1(new_n14224_), .A2(new_n11870_), .ZN(new_n14225_));
  AOI21_X1   g11322(.A1(new_n14223_), .A2(new_n11903_), .B(pi1155), .ZN(new_n14226_));
  INV_X1     g11323(.I(new_n14211_), .ZN(new_n14227_));
  XOR2_X1    g11324(.A1(new_n14217_), .A2(pi1153), .Z(new_n14228_));
  NAND2_X1   g11325(.A1(new_n14228_), .A2(new_n14227_), .ZN(new_n14229_));
  OAI21_X1   g11326(.A1(new_n14217_), .A2(new_n14207_), .B(new_n11893_), .ZN(new_n14230_));
  AOI21_X1   g11327(.A1(new_n14229_), .A2(new_n14230_), .B(new_n11891_), .ZN(new_n14231_));
  NOR2_X1    g11328(.A1(new_n14211_), .A2(pi0778), .ZN(new_n14232_));
  OAI21_X1   g11329(.A1(new_n14231_), .A2(new_n14232_), .B(pi0609), .ZN(new_n14233_));
  AOI21_X1   g11330(.A1(new_n14210_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n14234_));
  NOR2_X1    g11331(.A1(new_n14234_), .A2(pi0660), .ZN(new_n14235_));
  OAI21_X1   g11332(.A1(new_n14226_), .A2(new_n14233_), .B(new_n14235_), .ZN(new_n14236_));
  NOR2_X1    g11333(.A1(new_n14231_), .A2(new_n14232_), .ZN(new_n14237_));
  NAND4_X1   g11334(.A1(new_n14224_), .A2(pi0609), .A3(new_n11912_), .A4(new_n14237_), .ZN(new_n14238_));
  NOR2_X1    g11335(.A1(new_n14209_), .A2(new_n11925_), .ZN(new_n14239_));
  AOI21_X1   g11336(.A1(new_n14239_), .A2(new_n11928_), .B(pi1155), .ZN(new_n14240_));
  NOR2_X1    g11337(.A1(new_n14240_), .A2(new_n11923_), .ZN(new_n14241_));
  NAND2_X1   g11338(.A1(new_n14238_), .A2(new_n14241_), .ZN(new_n14242_));
  NAND3_X1   g11339(.A1(new_n14242_), .A2(pi0785), .A3(new_n14236_), .ZN(new_n14243_));
  NAND2_X1   g11340(.A1(new_n14243_), .A2(new_n14225_), .ZN(new_n14244_));
  INV_X1     g11341(.I(new_n14244_), .ZN(new_n14245_));
  NOR4_X1    g11342(.A1(new_n14237_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n14246_));
  NOR2_X1    g11343(.A1(new_n14239_), .A2(pi0785), .ZN(new_n14247_));
  OAI21_X1   g11344(.A1(new_n14240_), .A2(new_n14234_), .B(pi0785), .ZN(new_n14248_));
  XNOR2_X1   g11345(.A1(new_n14248_), .A2(new_n14247_), .ZN(new_n14249_));
  INV_X1     g11346(.I(new_n14249_), .ZN(new_n14250_));
  NOR2_X1    g11347(.A1(new_n14250_), .A2(new_n11945_), .ZN(new_n14251_));
  OR3_X2     g11348(.A1(new_n14246_), .A2(new_n14251_), .A3(pi0627), .Z(new_n14252_));
  OAI21_X1   g11349(.A1(new_n14250_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n14253_));
  NOR2_X1    g11350(.A1(new_n14237_), .A2(new_n11939_), .ZN(new_n14254_));
  NOR4_X1    g11351(.A1(new_n14245_), .A2(new_n11934_), .A3(pi1154), .A4(new_n14254_), .ZN(new_n14255_));
  OAI21_X1   g11352(.A1(new_n14255_), .A2(new_n14253_), .B(new_n11949_), .ZN(new_n14256_));
  AOI21_X1   g11353(.A1(new_n14256_), .A2(new_n14252_), .B(new_n11969_), .ZN(new_n14257_));
  AOI21_X1   g11354(.A1(new_n11969_), .A2(new_n14244_), .B(new_n14257_), .ZN(new_n14258_));
  INV_X1     g11355(.I(new_n14254_), .ZN(new_n14259_));
  NOR2_X1    g11356(.A1(new_n14259_), .A2(new_n11962_), .ZN(new_n14260_));
  NOR4_X1    g11357(.A1(new_n14258_), .A2(new_n11967_), .A3(pi1159), .A4(new_n14260_), .ZN(new_n14261_));
  NOR2_X1    g11358(.A1(new_n14250_), .A2(pi0781), .ZN(new_n14262_));
  NOR2_X1    g11359(.A1(new_n14253_), .A2(new_n14251_), .ZN(new_n14263_));
  NOR2_X1    g11360(.A1(new_n14263_), .A2(new_n11969_), .ZN(new_n14264_));
  XOR2_X1    g11361(.A1(new_n14264_), .A2(new_n14262_), .Z(new_n14265_));
  INV_X1     g11362(.I(new_n14265_), .ZN(new_n14266_));
  NOR2_X1    g11363(.A1(new_n14266_), .A2(new_n11967_), .ZN(new_n14267_));
  INV_X1     g11364(.I(new_n14207_), .ZN(new_n14268_));
  OAI21_X1   g11365(.A1(new_n14268_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n14269_));
  NOR4_X1    g11366(.A1(new_n14261_), .A2(new_n11966_), .A3(new_n14267_), .A4(new_n14269_), .ZN(new_n14270_));
  NOR4_X1    g11367(.A1(new_n14259_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n14271_));
  OAI21_X1   g11368(.A1(new_n14207_), .A2(pi0619), .B(new_n11869_), .ZN(new_n14272_));
  OAI21_X1   g11369(.A1(new_n14267_), .A2(new_n14272_), .B(new_n11966_), .ZN(new_n14273_));
  NOR2_X1    g11370(.A1(new_n14273_), .A2(new_n14271_), .ZN(new_n14274_));
  AOI21_X1   g11371(.A1(new_n14258_), .A2(new_n11998_), .B(pi0789), .ZN(new_n14275_));
  OAI21_X1   g11372(.A1(new_n14270_), .A2(new_n14274_), .B(new_n14275_), .ZN(new_n14276_));
  NOR2_X1    g11373(.A1(new_n14266_), .A2(pi0789), .ZN(new_n14277_));
  NOR3_X1    g11374(.A1(new_n14207_), .A2(pi0619), .A3(pi1159), .ZN(new_n14278_));
  NOR2_X1    g11375(.A1(new_n14278_), .A2(new_n11985_), .ZN(new_n14279_));
  XOR2_X1    g11376(.A1(new_n14277_), .A2(new_n14279_), .Z(new_n14280_));
  INV_X1     g11377(.I(new_n14280_), .ZN(new_n14281_));
  MUX2_X1    g11378(.I0(new_n14281_), .I1(new_n14207_), .S(new_n12003_), .Z(new_n14282_));
  NAND2_X1   g11379(.A1(new_n14282_), .A2(new_n12002_), .ZN(new_n14283_));
  AOI21_X1   g11380(.A1(new_n14260_), .A2(new_n12021_), .B(new_n11986_), .ZN(new_n14284_));
  NAND2_X1   g11381(.A1(new_n14283_), .A2(new_n14284_), .ZN(new_n14285_));
  NAND2_X1   g11382(.A1(new_n14276_), .A2(new_n14285_), .ZN(new_n14286_));
  NOR2_X1    g11383(.A1(new_n14286_), .A2(pi0792), .ZN(new_n14287_));
  NOR2_X1    g11384(.A1(new_n14280_), .A2(pi0788), .ZN(new_n14288_));
  AOI21_X1   g11385(.A1(new_n14282_), .A2(pi0788), .B(new_n14288_), .ZN(new_n14289_));
  INV_X1     g11386(.I(new_n14289_), .ZN(new_n14290_));
  NOR4_X1    g11387(.A1(new_n14286_), .A2(new_n12031_), .A3(pi1156), .A4(new_n14290_), .ZN(new_n14291_));
  NOR2_X1    g11388(.A1(new_n14260_), .A2(new_n12034_), .ZN(new_n14292_));
  INV_X1     g11389(.I(new_n14292_), .ZN(new_n14293_));
  OAI21_X1   g11390(.A1(new_n14293_), .A2(new_n13277_), .B(new_n12026_), .ZN(new_n14294_));
  NAND2_X1   g11391(.A1(new_n14294_), .A2(pi0629), .ZN(new_n14295_));
  AOI21_X1   g11392(.A1(new_n14286_), .A2(new_n12031_), .B(pi1156), .ZN(new_n14296_));
  NOR3_X1    g11393(.A1(new_n14296_), .A2(new_n12031_), .A3(new_n14289_), .ZN(new_n14297_));
  AOI21_X1   g11394(.A1(new_n14292_), .A2(new_n12042_), .B(pi0629), .ZN(new_n14298_));
  OAI22_X1   g11395(.A1(new_n14297_), .A2(new_n14298_), .B1(new_n14291_), .B2(new_n14295_), .ZN(new_n14299_));
  AOI21_X1   g11396(.A1(new_n14299_), .A2(pi0792), .B(new_n14287_), .ZN(new_n14300_));
  NOR2_X1    g11397(.A1(new_n12054_), .A2(new_n14207_), .ZN(new_n14301_));
  AOI21_X1   g11398(.A1(new_n14289_), .A2(new_n12054_), .B(new_n14301_), .ZN(new_n14302_));
  XNOR2_X1   g11399(.A1(new_n14300_), .A2(new_n14302_), .ZN(new_n14303_));
  NOR2_X1    g11400(.A1(new_n14303_), .A2(new_n12061_), .ZN(new_n14304_));
  XOR2_X1    g11401(.A1(new_n14304_), .A2(new_n14300_), .Z(new_n14305_));
  NOR2_X1    g11402(.A1(new_n14305_), .A2(pi1157), .ZN(new_n14306_));
  NOR2_X1    g11403(.A1(new_n14293_), .A2(new_n12068_), .ZN(new_n14307_));
  NOR2_X1    g11404(.A1(new_n14307_), .A2(new_n12061_), .ZN(new_n14308_));
  INV_X1     g11405(.I(new_n14308_), .ZN(new_n14309_));
  AOI21_X1   g11406(.A1(new_n14268_), .A2(new_n12061_), .B(pi1157), .ZN(new_n14310_));
  NAND2_X1   g11407(.A1(new_n14309_), .A2(new_n14310_), .ZN(new_n14311_));
  NAND2_X1   g11408(.A1(new_n14311_), .A2(new_n12060_), .ZN(new_n14312_));
  NOR2_X1    g11409(.A1(new_n14306_), .A2(new_n14312_), .ZN(new_n14313_));
  XOR2_X1    g11410(.A1(new_n14304_), .A2(new_n14302_), .Z(new_n14314_));
  NOR2_X1    g11411(.A1(new_n14314_), .A2(new_n12049_), .ZN(new_n14315_));
  NAND2_X1   g11412(.A1(new_n14207_), .A2(pi0647), .ZN(new_n14316_));
  NAND4_X1   g11413(.A1(new_n14309_), .A2(pi0630), .A3(new_n12049_), .A4(new_n14316_), .ZN(new_n14317_));
  OAI21_X1   g11414(.A1(new_n14315_), .A2(new_n14317_), .B(pi0787), .ZN(new_n14318_));
  OAI22_X1   g11415(.A1(new_n14318_), .A2(new_n14313_), .B1(pi0787), .B2(new_n14300_), .ZN(new_n14319_));
  OAI21_X1   g11416(.A1(new_n14319_), .A2(pi0644), .B(new_n12099_), .ZN(new_n14320_));
  INV_X1     g11417(.I(new_n14307_), .ZN(new_n14321_));
  NAND3_X1   g11418(.A1(new_n14268_), .A2(new_n12061_), .A3(new_n12049_), .ZN(new_n14322_));
  MUX2_X1    g11419(.I0(new_n14322_), .I1(new_n14321_), .S(new_n12048_), .Z(new_n14323_));
  NOR2_X1    g11420(.A1(new_n14323_), .A2(new_n12082_), .ZN(new_n14324_));
  NOR2_X1    g11421(.A1(new_n12092_), .A2(new_n14268_), .ZN(new_n14325_));
  AOI21_X1   g11422(.A1(new_n14302_), .A2(new_n12092_), .B(new_n14325_), .ZN(new_n14326_));
  NAND4_X1   g11423(.A1(new_n14326_), .A2(pi0644), .A3(new_n12099_), .A4(new_n14268_), .ZN(new_n14327_));
  NAND2_X1   g11424(.A1(new_n14327_), .A2(new_n12081_), .ZN(new_n14328_));
  AOI21_X1   g11425(.A1(new_n14320_), .A2(new_n14324_), .B(new_n14328_), .ZN(new_n14329_));
  NAND4_X1   g11426(.A1(new_n14319_), .A2(pi0644), .A3(new_n12099_), .A4(new_n14323_), .ZN(new_n14330_));
  AOI21_X1   g11427(.A1(new_n12082_), .A2(new_n14268_), .B(new_n14326_), .ZN(new_n14331_));
  NOR4_X1    g11428(.A1(new_n14302_), .A2(pi0644), .A3(new_n12091_), .A4(new_n14268_), .ZN(new_n14332_));
  NOR3_X1    g11429(.A1(new_n14331_), .A2(pi0715), .A3(new_n14332_), .ZN(new_n14333_));
  AOI21_X1   g11430(.A1(new_n14330_), .A2(new_n14333_), .B(pi1160), .ZN(new_n14334_));
  NOR2_X1    g11431(.A1(new_n14334_), .A2(new_n14329_), .ZN(new_n14335_));
  NOR3_X1    g11432(.A1(new_n14335_), .A2(new_n11867_), .A3(new_n14319_), .ZN(new_n14336_));
  INV_X1     g11433(.I(new_n14319_), .ZN(new_n14337_));
  AOI21_X1   g11434(.A1(new_n14335_), .A2(pi0790), .B(new_n14337_), .ZN(new_n14338_));
  OAI21_X1   g11435(.A1(new_n14336_), .A2(new_n14338_), .B(pi0832), .ZN(new_n14339_));
  NOR3_X1    g11436(.A1(new_n13368_), .A2(new_n3172_), .A3(new_n12113_), .ZN(new_n14340_));
  INV_X1     g11437(.I(new_n14340_), .ZN(new_n14341_));
  OAI21_X1   g11438(.A1(new_n12615_), .A2(new_n12602_), .B(new_n3154_), .ZN(new_n14342_));
  INV_X1     g11439(.I(new_n14342_), .ZN(new_n14343_));
  OAI21_X1   g11440(.A1(new_n12396_), .A2(new_n12436_), .B(new_n13820_), .ZN(new_n14344_));
  AOI21_X1   g11441(.A1(new_n12459_), .A2(pi0299), .B(new_n14344_), .ZN(new_n14345_));
  OAI21_X1   g11442(.A1(new_n14345_), .A2(new_n14343_), .B(new_n3172_), .ZN(new_n14346_));
  NAND2_X1   g11443(.A1(new_n14346_), .A2(new_n14341_), .ZN(new_n14347_));
  INV_X1     g11444(.I(pi0774), .ZN(new_n14348_));
  NOR3_X1    g11445(.A1(new_n12632_), .A2(pi0039), .A3(new_n12626_), .ZN(new_n14349_));
  NOR3_X1    g11446(.A1(new_n12501_), .A2(new_n3154_), .A3(new_n12514_), .ZN(new_n14350_));
  NOR3_X1    g11447(.A1(new_n14349_), .A2(pi0038), .A3(new_n14350_), .ZN(new_n14351_));
  NAND3_X1   g11448(.A1(new_n13372_), .A2(pi0038), .A3(new_n12113_), .ZN(new_n14352_));
  NAND4_X1   g11449(.A1(new_n14351_), .A2(pi0143), .A3(new_n14348_), .A4(new_n14352_), .ZN(new_n14353_));
  NAND3_X1   g11450(.A1(new_n14347_), .A2(new_n14353_), .A3(new_n10048_), .ZN(new_n14354_));
  NAND2_X1   g11451(.A1(new_n12794_), .A2(pi0038), .ZN(new_n14355_));
  NAND3_X1   g11452(.A1(new_n14355_), .A2(new_n10048_), .A3(new_n12901_), .ZN(new_n14356_));
  NAND2_X1   g11453(.A1(new_n14356_), .A2(new_n14348_), .ZN(new_n14357_));
  NOR2_X1    g11454(.A1(new_n5154_), .A2(new_n11877_), .ZN(new_n14358_));
  INV_X1     g11455(.I(new_n14358_), .ZN(new_n14359_));
  NOR2_X1    g11456(.A1(new_n14359_), .A2(new_n3172_), .ZN(new_n14360_));
  INV_X1     g11457(.I(new_n12693_), .ZN(new_n14361_));
  MUX2_X1    g11458(.I0(new_n14361_), .I1(new_n12667_), .S(new_n3154_), .Z(new_n14362_));
  NAND2_X1   g11459(.A1(new_n14362_), .A2(new_n3172_), .ZN(new_n14363_));
  AOI21_X1   g11460(.A1(new_n5156_), .A2(new_n12307_), .B(new_n3172_), .ZN(new_n14364_));
  AOI21_X1   g11461(.A1(new_n12824_), .A2(new_n3172_), .B(new_n14364_), .ZN(new_n14365_));
  NOR2_X1    g11462(.A1(pi0143), .A2(pi0774), .ZN(new_n14366_));
  AOI22_X1   g11463(.A1(new_n14363_), .A2(pi0143), .B1(new_n14365_), .B2(new_n14366_), .ZN(new_n14367_));
  NOR2_X1    g11464(.A1(new_n14367_), .A2(new_n14360_), .ZN(new_n14368_));
  NOR2_X1    g11465(.A1(new_n14368_), .A2(pi0687), .ZN(new_n14369_));
  NAND3_X1   g11466(.A1(new_n14369_), .A2(new_n14354_), .A3(new_n14357_), .ZN(new_n14370_));
  MUX2_X1    g11467(.I0(new_n14370_), .I1(new_n10048_), .S(new_n3232_), .Z(new_n14371_));
  INV_X1     g11468(.I(new_n14371_), .ZN(new_n14372_));
  NAND2_X1   g11469(.A1(new_n14371_), .A2(pi0625), .ZN(new_n14373_));
  NOR2_X1    g11470(.A1(new_n3231_), .A2(pi0143), .ZN(new_n14374_));
  INV_X1     g11471(.I(new_n14374_), .ZN(new_n14375_));
  NOR2_X1    g11472(.A1(new_n14356_), .A2(new_n14348_), .ZN(new_n14376_));
  OAI21_X1   g11473(.A1(new_n14367_), .A2(new_n14360_), .B(new_n3231_), .ZN(new_n14377_));
  OAI21_X1   g11474(.A1(new_n14376_), .A2(new_n14377_), .B(new_n14375_), .ZN(new_n14378_));
  INV_X1     g11475(.I(new_n14378_), .ZN(new_n14379_));
  AOI21_X1   g11476(.A1(new_n14379_), .A2(new_n12970_), .B(pi1153), .ZN(new_n14380_));
  NAND2_X1   g11477(.A1(new_n14373_), .A2(new_n14380_), .ZN(new_n14381_));
  MUX2_X1    g11478(.I0(new_n12937_), .I1(new_n12602_), .S(new_n3154_), .Z(new_n14382_));
  NAND3_X1   g11479(.A1(new_n14382_), .A2(new_n10048_), .A3(new_n13395_), .ZN(new_n14383_));
  AOI21_X1   g11480(.A1(new_n13399_), .A2(new_n10048_), .B(new_n13395_), .ZN(new_n14384_));
  NAND2_X1   g11481(.A1(new_n13368_), .A2(new_n10048_), .ZN(new_n14385_));
  NAND4_X1   g11482(.A1(new_n14385_), .A2(new_n3172_), .A3(new_n14216_), .A4(new_n13403_), .ZN(new_n14386_));
  NOR2_X1    g11483(.A1(new_n14384_), .A2(new_n14386_), .ZN(new_n14387_));
  AOI22_X1   g11484(.A1(new_n14387_), .A2(new_n14383_), .B1(new_n14216_), .B2(new_n14356_), .ZN(new_n14388_));
  NOR3_X1    g11485(.A1(new_n14388_), .A2(new_n3232_), .A3(new_n14375_), .ZN(new_n14389_));
  OAI21_X1   g11486(.A1(new_n14388_), .A2(new_n3232_), .B(new_n14375_), .ZN(new_n14390_));
  INV_X1     g11487(.I(new_n14390_), .ZN(new_n14391_));
  NOR3_X1    g11488(.A1(new_n14391_), .A2(new_n12970_), .A3(new_n14389_), .ZN(new_n14392_));
  NAND3_X1   g11489(.A1(new_n12793_), .A2(pi0039), .A3(new_n12853_), .ZN(new_n14393_));
  OAI21_X1   g11490(.A1(new_n12894_), .A2(new_n3154_), .B(new_n12854_), .ZN(new_n14394_));
  AOI21_X1   g11491(.A1(new_n14394_), .A2(new_n14393_), .B(pi0038), .ZN(new_n14395_));
  OAI21_X1   g11492(.A1(new_n14395_), .A2(new_n12900_), .B(new_n3231_), .ZN(new_n14396_));
  NAND2_X1   g11493(.A1(new_n14396_), .A2(new_n10048_), .ZN(new_n14397_));
  OAI21_X1   g11494(.A1(new_n14397_), .A2(new_n12970_), .B(new_n11893_), .ZN(new_n14398_));
  NOR3_X1    g11495(.A1(new_n14392_), .A2(new_n13657_), .A3(new_n14398_), .ZN(new_n14399_));
  NAND2_X1   g11496(.A1(new_n14387_), .A2(new_n14383_), .ZN(new_n14400_));
  NAND2_X1   g11497(.A1(new_n14356_), .A2(new_n14216_), .ZN(new_n14401_));
  NAND2_X1   g11498(.A1(new_n14400_), .A2(new_n14401_), .ZN(new_n14402_));
  NAND3_X1   g11499(.A1(new_n14402_), .A2(new_n3231_), .A3(new_n14374_), .ZN(new_n14403_));
  NAND3_X1   g11500(.A1(new_n14403_), .A2(pi0625), .A3(new_n14390_), .ZN(new_n14404_));
  AOI21_X1   g11501(.A1(new_n14397_), .A2(new_n12970_), .B(pi1153), .ZN(new_n14405_));
  OAI21_X1   g11502(.A1(new_n14379_), .A2(new_n12970_), .B(new_n12977_), .ZN(new_n14406_));
  AOI21_X1   g11503(.A1(new_n14404_), .A2(new_n14405_), .B(new_n14406_), .ZN(new_n14407_));
  AOI22_X1   g11504(.A1(new_n14381_), .A2(new_n14399_), .B1(new_n14373_), .B2(new_n14407_), .ZN(new_n14408_));
  NOR3_X1    g11505(.A1(new_n14408_), .A2(new_n11891_), .A3(new_n14372_), .ZN(new_n14409_));
  AOI21_X1   g11506(.A1(new_n14408_), .A2(pi0778), .B(new_n14371_), .ZN(new_n14410_));
  NOR2_X1    g11507(.A1(new_n14409_), .A2(new_n14410_), .ZN(new_n14411_));
  NAND2_X1   g11508(.A1(new_n14411_), .A2(new_n11870_), .ZN(new_n14412_));
  NOR3_X1    g11509(.A1(new_n14391_), .A2(pi0778), .A3(new_n14389_), .ZN(new_n14413_));
  INV_X1     g11510(.I(new_n14413_), .ZN(new_n14414_));
  NOR3_X1    g11511(.A1(new_n14392_), .A2(new_n14398_), .A3(new_n14405_), .ZN(new_n14415_));
  NOR3_X1    g11512(.A1(new_n14415_), .A2(new_n11891_), .A3(new_n14414_), .ZN(new_n14416_));
  NAND4_X1   g11513(.A1(new_n14404_), .A2(new_n12970_), .A3(new_n11893_), .A4(new_n14397_), .ZN(new_n14417_));
  AOI21_X1   g11514(.A1(new_n14417_), .A2(pi0778), .B(new_n14413_), .ZN(new_n14418_));
  OAI21_X1   g11515(.A1(new_n14416_), .A2(new_n14418_), .B(new_n11903_), .ZN(new_n14419_));
  NAND2_X1   g11516(.A1(new_n14397_), .A2(new_n12997_), .ZN(new_n14420_));
  NAND3_X1   g11517(.A1(new_n14379_), .A2(new_n11903_), .A3(new_n11924_), .ZN(new_n14421_));
  AOI21_X1   g11518(.A1(new_n14421_), .A2(new_n14420_), .B(pi1155), .ZN(new_n14422_));
  OAI21_X1   g11519(.A1(new_n14422_), .A2(new_n11923_), .B(pi0609), .ZN(new_n14423_));
  AOI21_X1   g11520(.A1(new_n14419_), .A2(pi1155), .B(new_n14423_), .ZN(new_n14424_));
  INV_X1     g11521(.I(new_n14380_), .ZN(new_n14425_));
  AOI21_X1   g11522(.A1(new_n14371_), .A2(pi0625), .B(new_n14425_), .ZN(new_n14426_));
  OR3_X2     g11523(.A1(new_n14392_), .A2(new_n13657_), .A3(new_n14398_), .Z(new_n14427_));
  NAND2_X1   g11524(.A1(new_n14407_), .A2(new_n14373_), .ZN(new_n14428_));
  OAI21_X1   g11525(.A1(new_n14427_), .A2(new_n14426_), .B(new_n14428_), .ZN(new_n14429_));
  NAND3_X1   g11526(.A1(new_n14429_), .A2(pi0778), .A3(new_n14371_), .ZN(new_n14430_));
  OAI21_X1   g11527(.A1(new_n14429_), .A2(new_n11891_), .B(new_n14372_), .ZN(new_n14431_));
  NAND3_X1   g11528(.A1(new_n14431_), .A2(new_n14430_), .A3(new_n11903_), .ZN(new_n14432_));
  NAND3_X1   g11529(.A1(new_n14417_), .A2(pi0778), .A3(new_n14413_), .ZN(new_n14433_));
  OAI21_X1   g11530(.A1(new_n14415_), .A2(new_n11891_), .B(new_n14414_), .ZN(new_n14434_));
  NAND2_X1   g11531(.A1(new_n14434_), .A2(new_n14433_), .ZN(new_n14435_));
  NOR2_X1    g11532(.A1(new_n14378_), .A2(new_n11914_), .ZN(new_n14436_));
  AOI22_X1   g11533(.A1(new_n14436_), .A2(pi0609), .B1(new_n13010_), .B2(new_n14397_), .ZN(new_n14437_));
  NOR2_X1    g11534(.A1(new_n11923_), .A2(pi1155), .ZN(new_n14438_));
  INV_X1     g11535(.I(new_n14438_), .ZN(new_n14439_));
  AOI21_X1   g11536(.A1(new_n14435_), .A2(pi0609), .B(new_n14439_), .ZN(new_n14440_));
  AOI22_X1   g11537(.A1(new_n14432_), .A2(new_n14440_), .B1(new_n14411_), .B2(new_n14424_), .ZN(new_n14441_));
  NOR3_X1    g11538(.A1(new_n14441_), .A2(new_n11870_), .A3(new_n14412_), .ZN(new_n14442_));
  NAND2_X1   g11539(.A1(new_n14431_), .A2(new_n14430_), .ZN(new_n14443_));
  NOR2_X1    g11540(.A1(new_n14443_), .A2(pi0785), .ZN(new_n14444_));
  INV_X1     g11541(.I(new_n14424_), .ZN(new_n14445_));
  NOR3_X1    g11542(.A1(new_n14409_), .A2(new_n14410_), .A3(pi0609), .ZN(new_n14446_));
  INV_X1     g11543(.I(new_n14440_), .ZN(new_n14447_));
  OAI22_X1   g11544(.A1(new_n14443_), .A2(new_n14445_), .B1(new_n14446_), .B2(new_n14447_), .ZN(new_n14448_));
  AOI21_X1   g11545(.A1(new_n14448_), .A2(pi0785), .B(new_n14444_), .ZN(new_n14449_));
  NOR3_X1    g11546(.A1(new_n14449_), .A2(new_n14442_), .A3(pi0781), .ZN(new_n14450_));
  INV_X1     g11547(.I(new_n14450_), .ZN(new_n14451_));
  NOR2_X1    g11548(.A1(new_n14449_), .A2(new_n14442_), .ZN(new_n14452_));
  NOR2_X1    g11549(.A1(new_n14397_), .A2(new_n11938_), .ZN(new_n14453_));
  AOI21_X1   g11550(.A1(new_n14435_), .A2(new_n11938_), .B(new_n14453_), .ZN(new_n14454_));
  OAI21_X1   g11551(.A1(new_n14454_), .A2(pi0618), .B(pi1154), .ZN(new_n14455_));
  INV_X1     g11552(.I(new_n14397_), .ZN(new_n14456_));
  AOI21_X1   g11553(.A1(new_n14456_), .A2(new_n11914_), .B(pi0785), .ZN(new_n14457_));
  OAI21_X1   g11554(.A1(new_n14379_), .A2(new_n11914_), .B(new_n14457_), .ZN(new_n14458_));
  NOR2_X1    g11555(.A1(new_n14437_), .A2(new_n11912_), .ZN(new_n14459_));
  OAI21_X1   g11556(.A1(new_n14459_), .A2(new_n14422_), .B(pi0785), .ZN(new_n14460_));
  OR2_X2     g11557(.A1(new_n14460_), .A2(new_n14458_), .Z(new_n14461_));
  NAND2_X1   g11558(.A1(new_n14460_), .A2(new_n14458_), .ZN(new_n14462_));
  NAND3_X1   g11559(.A1(new_n14461_), .A2(pi0618), .A3(new_n14462_), .ZN(new_n14463_));
  NAND2_X1   g11560(.A1(new_n14456_), .A2(pi0618), .ZN(new_n14464_));
  NAND4_X1   g11561(.A1(new_n14463_), .A2(pi0627), .A3(new_n11950_), .A4(new_n14464_), .ZN(new_n14465_));
  AND3_X2    g11562(.A1(new_n14465_), .A2(pi0618), .A3(new_n14455_), .Z(new_n14466_));
  NAND3_X1   g11563(.A1(new_n14448_), .A2(pi0785), .A3(new_n14444_), .ZN(new_n14467_));
  OAI21_X1   g11564(.A1(new_n14441_), .A2(new_n11870_), .B(new_n14412_), .ZN(new_n14468_));
  NAND3_X1   g11565(.A1(new_n14467_), .A2(new_n14468_), .A3(new_n11934_), .ZN(new_n14469_));
  NOR2_X1    g11566(.A1(new_n14454_), .A2(new_n11934_), .ZN(new_n14470_));
  AOI21_X1   g11567(.A1(new_n14397_), .A2(new_n11934_), .B(pi1154), .ZN(new_n14471_));
  AOI21_X1   g11568(.A1(new_n14463_), .A2(new_n14471_), .B(pi0627), .ZN(new_n14472_));
  NOR3_X1    g11569(.A1(new_n14472_), .A2(pi1154), .A3(new_n14470_), .ZN(new_n14473_));
  AOI22_X1   g11570(.A1(new_n14469_), .A2(new_n14473_), .B1(new_n14452_), .B2(new_n14466_), .ZN(new_n14474_));
  NOR3_X1    g11571(.A1(new_n14474_), .A2(new_n11969_), .A3(new_n14451_), .ZN(new_n14475_));
  NAND3_X1   g11572(.A1(new_n14467_), .A2(new_n14468_), .A3(new_n14466_), .ZN(new_n14476_));
  NOR3_X1    g11573(.A1(new_n14449_), .A2(new_n14442_), .A3(pi0618), .ZN(new_n14477_));
  INV_X1     g11574(.I(new_n14473_), .ZN(new_n14478_));
  OAI21_X1   g11575(.A1(new_n14477_), .A2(new_n14478_), .B(new_n14476_), .ZN(new_n14479_));
  AOI21_X1   g11576(.A1(new_n14479_), .A2(pi0781), .B(new_n14450_), .ZN(new_n14480_));
  NOR3_X1    g11577(.A1(new_n14475_), .A2(new_n14480_), .A3(pi0789), .ZN(new_n14481_));
  INV_X1     g11578(.I(new_n14481_), .ZN(new_n14482_));
  MUX2_X1    g11579(.I0(new_n14479_), .I1(new_n14452_), .S(new_n11969_), .Z(new_n14483_));
  NAND2_X1   g11580(.A1(new_n14461_), .A2(new_n14462_), .ZN(new_n14484_));
  INV_X1     g11581(.I(new_n14484_), .ZN(new_n14485_));
  NAND3_X1   g11582(.A1(new_n14397_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n14486_));
  MUX2_X1    g11583(.I0(new_n14486_), .I1(new_n14485_), .S(new_n11969_), .Z(new_n14487_));
  NAND2_X1   g11584(.A1(new_n14487_), .A2(pi0619), .ZN(new_n14488_));
  AOI21_X1   g11585(.A1(new_n14456_), .A2(pi0619), .B(pi1159), .ZN(new_n14489_));
  AND3_X2    g11586(.A1(new_n14488_), .A2(pi0648), .A3(new_n14489_), .Z(new_n14490_));
  NAND2_X1   g11587(.A1(new_n14454_), .A2(new_n11961_), .ZN(new_n14491_));
  OAI21_X1   g11588(.A1(new_n11961_), .A2(new_n14456_), .B(new_n14491_), .ZN(new_n14492_));
  INV_X1     g11589(.I(new_n14492_), .ZN(new_n14493_));
  NOR3_X1    g11590(.A1(new_n14490_), .A2(new_n11967_), .A3(pi1159), .ZN(new_n14494_));
  NAND3_X1   g11591(.A1(new_n14479_), .A2(pi0781), .A3(new_n14450_), .ZN(new_n14495_));
  OAI21_X1   g11592(.A1(new_n14474_), .A2(new_n11969_), .B(new_n14451_), .ZN(new_n14496_));
  NAND3_X1   g11593(.A1(new_n14496_), .A2(new_n14495_), .A3(new_n11967_), .ZN(new_n14497_));
  AOI21_X1   g11594(.A1(new_n14397_), .A2(new_n11967_), .B(pi1159), .ZN(new_n14498_));
  AOI21_X1   g11595(.A1(new_n14488_), .A2(new_n14498_), .B(pi0648), .ZN(new_n14499_));
  NOR2_X1    g11596(.A1(new_n14492_), .A2(new_n11967_), .ZN(new_n14500_));
  NOR3_X1    g11597(.A1(new_n14499_), .A2(pi1159), .A3(new_n14500_), .ZN(new_n14501_));
  AOI22_X1   g11598(.A1(new_n14497_), .A2(new_n14501_), .B1(new_n14483_), .B2(new_n14494_), .ZN(new_n14502_));
  NOR3_X1    g11599(.A1(new_n14502_), .A2(new_n11985_), .A3(new_n14482_), .ZN(new_n14503_));
  NAND3_X1   g11600(.A1(new_n14496_), .A2(new_n14495_), .A3(new_n14494_), .ZN(new_n14504_));
  NOR3_X1    g11601(.A1(new_n14475_), .A2(new_n14480_), .A3(pi0619), .ZN(new_n14505_));
  INV_X1     g11602(.I(new_n14501_), .ZN(new_n14506_));
  OAI21_X1   g11603(.A1(new_n14505_), .A2(new_n14506_), .B(new_n14504_), .ZN(new_n14507_));
  AOI21_X1   g11604(.A1(new_n14507_), .A2(pi0789), .B(new_n14481_), .ZN(new_n14508_));
  NOR2_X1    g11605(.A1(new_n14508_), .A2(new_n14503_), .ZN(new_n14509_));
  INV_X1     g11606(.I(new_n14509_), .ZN(new_n14510_));
  NAND3_X1   g11607(.A1(new_n14507_), .A2(pi0789), .A3(new_n14481_), .ZN(new_n14511_));
  OAI21_X1   g11608(.A1(new_n14502_), .A2(new_n11985_), .B(new_n14482_), .ZN(new_n14512_));
  NOR2_X1    g11609(.A1(new_n14397_), .A2(new_n12014_), .ZN(new_n14513_));
  AOI21_X1   g11610(.A1(new_n14493_), .A2(new_n12014_), .B(new_n14513_), .ZN(new_n14514_));
  NOR2_X1    g11611(.A1(new_n11989_), .A2(pi0626), .ZN(new_n14515_));
  INV_X1     g11612(.I(new_n14515_), .ZN(new_n14516_));
  AOI21_X1   g11613(.A1(new_n14512_), .A2(new_n14511_), .B(new_n14516_), .ZN(new_n14517_));
  NOR2_X1    g11614(.A1(new_n11994_), .A2(pi0641), .ZN(new_n14518_));
  INV_X1     g11615(.I(new_n14518_), .ZN(new_n14519_));
  AOI21_X1   g11616(.A1(new_n14512_), .A2(new_n14511_), .B(new_n14519_), .ZN(new_n14520_));
  NAND3_X1   g11617(.A1(new_n14397_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n14521_));
  MUX2_X1    g11618(.I0(new_n14521_), .I1(new_n14487_), .S(new_n11985_), .Z(new_n14522_));
  NAND2_X1   g11619(.A1(new_n14522_), .A2(pi0626), .ZN(new_n14523_));
  AOI21_X1   g11620(.A1(new_n14397_), .A2(new_n11994_), .B(pi1158), .ZN(new_n14524_));
  AOI21_X1   g11621(.A1(new_n14523_), .A2(new_n14524_), .B(new_n12016_), .ZN(new_n14525_));
  NAND2_X1   g11622(.A1(new_n14456_), .A2(pi0626), .ZN(new_n14526_));
  NAND4_X1   g11623(.A1(new_n14523_), .A2(pi0641), .A3(new_n11987_), .A4(new_n14526_), .ZN(new_n14527_));
  INV_X1     g11624(.I(new_n14527_), .ZN(new_n14528_));
  NOR2_X1    g11625(.A1(new_n14528_), .A2(new_n14525_), .ZN(new_n14529_));
  INV_X1     g11626(.I(new_n14529_), .ZN(new_n14530_));
  NOR3_X1    g11627(.A1(new_n14517_), .A2(new_n14520_), .A3(new_n14530_), .ZN(new_n14531_));
  NOR3_X1    g11628(.A1(new_n14531_), .A2(new_n11986_), .A3(new_n14510_), .ZN(new_n14532_));
  AOI21_X1   g11629(.A1(new_n14531_), .A2(pi0788), .B(new_n14509_), .ZN(new_n14533_));
  NOR2_X1    g11630(.A1(new_n14532_), .A2(new_n14533_), .ZN(new_n14534_));
  NAND3_X1   g11631(.A1(new_n14397_), .A2(new_n11994_), .A3(new_n11987_), .ZN(new_n14535_));
  MUX2_X1    g11632(.I0(new_n14535_), .I1(new_n14522_), .S(new_n11986_), .Z(new_n14536_));
  NOR2_X1    g11633(.A1(new_n14536_), .A2(pi0628), .ZN(new_n14537_));
  NOR2_X1    g11634(.A1(new_n14456_), .A2(new_n13114_), .ZN(new_n14538_));
  AOI21_X1   g11635(.A1(new_n14514_), .A2(new_n13114_), .B(new_n14538_), .ZN(new_n14539_));
  NOR3_X1    g11636(.A1(new_n14397_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n14540_));
  OAI21_X1   g11637(.A1(new_n14540_), .A2(new_n12030_), .B(pi0628), .ZN(new_n14541_));
  INV_X1     g11638(.I(new_n14541_), .ZN(new_n14542_));
  OAI21_X1   g11639(.A1(new_n14537_), .A2(new_n12026_), .B(new_n14542_), .ZN(new_n14543_));
  INV_X1     g11640(.I(new_n14543_), .ZN(new_n14544_));
  NOR2_X1    g11641(.A1(new_n14536_), .A2(new_n12031_), .ZN(new_n14545_));
  NOR2_X1    g11642(.A1(new_n12030_), .A2(pi0628), .ZN(new_n14546_));
  OAI21_X1   g11643(.A1(new_n14545_), .A2(pi1156), .B(new_n14546_), .ZN(new_n14547_));
  INV_X1     g11644(.I(new_n14547_), .ZN(new_n14548_));
  OAI22_X1   g11645(.A1(new_n14532_), .A2(new_n14533_), .B1(new_n14544_), .B2(new_n14548_), .ZN(new_n14549_));
  MUX2_X1    g11646(.I0(new_n14549_), .I1(new_n14534_), .S(new_n11868_), .Z(new_n14550_));
  OAI21_X1   g11647(.A1(new_n14508_), .A2(new_n14503_), .B(new_n14515_), .ZN(new_n14551_));
  OAI21_X1   g11648(.A1(new_n14508_), .A2(new_n14503_), .B(new_n14518_), .ZN(new_n14552_));
  NAND3_X1   g11649(.A1(new_n14551_), .A2(new_n14552_), .A3(new_n14529_), .ZN(new_n14553_));
  NAND3_X1   g11650(.A1(new_n14553_), .A2(pi0788), .A3(new_n14509_), .ZN(new_n14554_));
  OAI21_X1   g11651(.A1(new_n14553_), .A2(new_n11986_), .B(new_n14510_), .ZN(new_n14555_));
  AOI21_X1   g11652(.A1(new_n14555_), .A2(new_n14554_), .B(new_n14543_), .ZN(new_n14556_));
  NAND3_X1   g11653(.A1(new_n14556_), .A2(new_n14534_), .A3(pi0792), .ZN(new_n14557_));
  MUX2_X1    g11654(.I0(new_n14553_), .I1(new_n14510_), .S(new_n11986_), .Z(new_n14558_));
  AOI22_X1   g11655(.A1(new_n14555_), .A2(new_n14554_), .B1(new_n14543_), .B2(new_n14547_), .ZN(new_n14559_));
  OAI21_X1   g11656(.A1(new_n14559_), .A2(new_n11868_), .B(new_n14558_), .ZN(new_n14560_));
  NOR2_X1    g11657(.A1(new_n14456_), .A2(new_n12054_), .ZN(new_n14561_));
  AOI21_X1   g11658(.A1(new_n14536_), .A2(new_n12054_), .B(new_n14561_), .ZN(new_n14562_));
  AOI21_X1   g11659(.A1(new_n14562_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n14563_));
  NOR4_X1    g11660(.A1(new_n14539_), .A2(new_n12031_), .A3(pi1156), .A4(new_n14456_), .ZN(new_n14564_));
  NOR2_X1    g11661(.A1(new_n14564_), .A2(new_n14540_), .ZN(new_n14565_));
  MUX2_X1    g11662(.I0(new_n14565_), .I1(new_n14539_), .S(new_n11868_), .Z(new_n14566_));
  NAND2_X1   g11663(.A1(new_n14566_), .A2(pi0647), .ZN(new_n14567_));
  INV_X1     g11664(.I(new_n14567_), .ZN(new_n14568_));
  NOR2_X1    g11665(.A1(new_n14397_), .A2(new_n12061_), .ZN(new_n14569_));
  NOR4_X1    g11666(.A1(new_n14568_), .A2(new_n12060_), .A3(pi1157), .A4(new_n14569_), .ZN(new_n14570_));
  NOR3_X1    g11667(.A1(new_n14570_), .A2(new_n12061_), .A3(new_n14563_), .ZN(new_n14571_));
  NAND3_X1   g11668(.A1(new_n14560_), .A2(new_n14557_), .A3(new_n14571_), .ZN(new_n14572_));
  NOR3_X1    g11669(.A1(new_n14549_), .A2(new_n11868_), .A3(new_n14558_), .ZN(new_n14573_));
  AOI21_X1   g11670(.A1(new_n14549_), .A2(pi0792), .B(new_n14534_), .ZN(new_n14574_));
  NOR3_X1    g11671(.A1(new_n14573_), .A2(new_n14574_), .A3(pi0647), .ZN(new_n14575_));
  AOI21_X1   g11672(.A1(new_n14397_), .A2(new_n12061_), .B(pi1157), .ZN(new_n14576_));
  NAND2_X1   g11673(.A1(new_n14567_), .A2(new_n14576_), .ZN(new_n14577_));
  NAND2_X1   g11674(.A1(new_n14577_), .A2(new_n12060_), .ZN(new_n14578_));
  AOI21_X1   g11675(.A1(new_n14562_), .A2(pi0647), .B(pi1157), .ZN(new_n14579_));
  AND2_X2    g11676(.A1(new_n14578_), .A2(new_n14579_), .Z(new_n14580_));
  INV_X1     g11677(.I(new_n14580_), .ZN(new_n14581_));
  OAI21_X1   g11678(.A1(new_n14575_), .A2(new_n14581_), .B(new_n14572_), .ZN(new_n14582_));
  MUX2_X1    g11679(.I0(new_n14582_), .I1(new_n14550_), .S(new_n12048_), .Z(new_n14583_));
  NAND2_X1   g11680(.A1(new_n14566_), .A2(new_n12048_), .ZN(new_n14584_));
  NAND3_X1   g11681(.A1(new_n14397_), .A2(new_n12061_), .A3(new_n12049_), .ZN(new_n14585_));
  NAND2_X1   g11682(.A1(new_n14585_), .A2(pi0787), .ZN(new_n14586_));
  XOR2_X1    g11683(.A1(new_n14584_), .A2(new_n14586_), .Z(new_n14587_));
  NOR2_X1    g11684(.A1(new_n14397_), .A2(new_n12092_), .ZN(new_n14588_));
  AOI21_X1   g11685(.A1(new_n14562_), .A2(new_n12092_), .B(new_n14588_), .ZN(new_n14589_));
  INV_X1     g11686(.I(new_n14589_), .ZN(new_n14590_));
  NOR2_X1    g11687(.A1(pi0644), .A2(pi0715), .ZN(new_n14591_));
  AOI21_X1   g11688(.A1(new_n14590_), .A2(new_n14591_), .B(new_n13169_), .ZN(new_n14592_));
  OAI21_X1   g11689(.A1(new_n14587_), .A2(new_n12082_), .B(new_n14592_), .ZN(new_n14593_));
  AOI21_X1   g11690(.A1(new_n14583_), .A2(new_n12082_), .B(new_n14593_), .ZN(new_n14594_));
  INV_X1     g11691(.I(new_n14550_), .ZN(new_n14595_));
  NAND3_X1   g11692(.A1(new_n14560_), .A2(new_n14557_), .A3(new_n12061_), .ZN(new_n14596_));
  AOI22_X1   g11693(.A1(new_n14596_), .A2(new_n14580_), .B1(new_n14550_), .B2(new_n14571_), .ZN(new_n14597_));
  MUX2_X1    g11694(.I0(new_n14597_), .I1(new_n14595_), .S(new_n12048_), .Z(new_n14598_));
  INV_X1     g11695(.I(new_n14587_), .ZN(new_n14599_));
  NAND3_X1   g11696(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n14600_));
  OAI21_X1   g11697(.A1(new_n14589_), .A2(new_n14600_), .B(new_n13179_), .ZN(new_n14601_));
  NOR2_X1    g11698(.A1(new_n14599_), .A2(new_n14601_), .ZN(new_n14602_));
  OAI21_X1   g11699(.A1(new_n14598_), .A2(new_n12082_), .B(new_n14602_), .ZN(new_n14603_));
  NOR2_X1    g11700(.A1(new_n14594_), .A2(new_n14603_), .ZN(new_n14604_));
  NAND2_X1   g11701(.A1(po1038), .A2(new_n10048_), .ZN(new_n14605_));
  AOI21_X1   g11702(.A1(new_n14605_), .A2(new_n13184_), .B(po1038), .ZN(new_n14606_));
  OAI21_X1   g11703(.A1(new_n14583_), .A2(pi0790), .B(new_n14606_), .ZN(new_n14607_));
  OAI21_X1   g11704(.A1(new_n14604_), .A2(new_n14607_), .B(new_n14339_), .ZN(po0300));
  NOR2_X1    g11705(.A1(new_n2925_), .A2(new_n7504_), .ZN(new_n14609_));
  AOI21_X1   g11706(.A1(new_n11886_), .A2(pi0736), .B(new_n14609_), .ZN(new_n14610_));
  INV_X1     g11707(.I(pi0736), .ZN(new_n14611_));
  NOR3_X1    g11708(.A1(new_n11894_), .A2(new_n12970_), .A3(new_n14611_), .ZN(new_n14612_));
  NOR2_X1    g11709(.A1(new_n14609_), .A2(new_n11893_), .ZN(new_n14613_));
  INV_X1     g11710(.I(new_n14613_), .ZN(new_n14614_));
  OAI21_X1   g11711(.A1(new_n14612_), .A2(new_n14610_), .B(new_n11893_), .ZN(new_n14615_));
  OAI21_X1   g11712(.A1(new_n14612_), .A2(new_n14614_), .B(new_n14615_), .ZN(new_n14616_));
  MUX2_X1    g11713(.I0(new_n14616_), .I1(new_n14610_), .S(new_n11891_), .Z(new_n14617_));
  INV_X1     g11714(.I(new_n14617_), .ZN(new_n14618_));
  NOR2_X1    g11715(.A1(new_n14618_), .A2(new_n13717_), .ZN(new_n14619_));
  INV_X1     g11716(.I(new_n14619_), .ZN(new_n14620_));
  NOR2_X1    g11717(.A1(new_n14620_), .A2(new_n12066_), .ZN(new_n14621_));
  AOI21_X1   g11718(.A1(new_n14621_), .A2(new_n13748_), .B(new_n14609_), .ZN(new_n14622_));
  INV_X1     g11719(.I(new_n14622_), .ZN(new_n14623_));
  INV_X1     g11720(.I(new_n11997_), .ZN(new_n14624_));
  NOR2_X1    g11721(.A1(new_n11912_), .A2(pi0609), .ZN(new_n14625_));
  OAI21_X1   g11722(.A1(new_n13621_), .A2(new_n14625_), .B(pi0785), .ZN(new_n14626_));
  INV_X1     g11723(.I(new_n14626_), .ZN(new_n14627_));
  INV_X1     g11724(.I(pi0758), .ZN(new_n14628_));
  NOR2_X1    g11725(.A1(new_n11877_), .A2(new_n14628_), .ZN(new_n14629_));
  INV_X1     g11726(.I(new_n14629_), .ZN(new_n14630_));
  NOR2_X1    g11727(.A1(new_n14630_), .A2(new_n14627_), .ZN(new_n14631_));
  INV_X1     g11728(.I(new_n14631_), .ZN(new_n14632_));
  NOR2_X1    g11729(.A1(new_n11934_), .A2(pi1154), .ZN(new_n14633_));
  NOR2_X1    g11730(.A1(new_n11950_), .A2(pi0618), .ZN(new_n14634_));
  NOR2_X1    g11731(.A1(new_n14633_), .A2(new_n14634_), .ZN(new_n14635_));
  NOR2_X1    g11732(.A1(new_n14635_), .A2(new_n11969_), .ZN(new_n14636_));
  NOR2_X1    g11733(.A1(new_n14636_), .A2(new_n11914_), .ZN(new_n14637_));
  NOR2_X1    g11734(.A1(new_n11967_), .A2(pi1159), .ZN(new_n14638_));
  NOR2_X1    g11735(.A1(new_n11869_), .A2(pi0619), .ZN(new_n14639_));
  NOR2_X1    g11736(.A1(new_n14638_), .A2(new_n14639_), .ZN(new_n14640_));
  NOR2_X1    g11737(.A1(new_n14640_), .A2(new_n11985_), .ZN(new_n14641_));
  INV_X1     g11738(.I(new_n14641_), .ZN(new_n14642_));
  NOR2_X1    g11739(.A1(new_n14637_), .A2(new_n14642_), .ZN(new_n14643_));
  INV_X1     g11740(.I(new_n14643_), .ZN(new_n14644_));
  NOR2_X1    g11741(.A1(new_n14632_), .A2(new_n14644_), .ZN(new_n14645_));
  NAND2_X1   g11742(.A1(new_n14645_), .A2(new_n14624_), .ZN(new_n14646_));
  NOR2_X1    g11743(.A1(new_n14646_), .A2(new_n12053_), .ZN(new_n14647_));
  NOR2_X1    g11744(.A1(new_n14621_), .A2(new_n12060_), .ZN(new_n14648_));
  OAI22_X1   g11745(.A1(new_n14648_), .A2(pi0647), .B1(new_n12060_), .B2(new_n14647_), .ZN(new_n14649_));
  OAI21_X1   g11746(.A1(new_n14620_), .A2(new_n12066_), .B(new_n12060_), .ZN(new_n14650_));
  AOI22_X1   g11747(.A1(new_n14650_), .A2(pi0647), .B1(pi0630), .B2(new_n14647_), .ZN(new_n14651_));
  AOI21_X1   g11748(.A1(new_n14651_), .A2(pi1157), .B(new_n14649_), .ZN(new_n14652_));
  INV_X1     g11749(.I(new_n14649_), .ZN(new_n14653_));
  NOR3_X1    g11750(.A1(new_n14653_), .A2(new_n14651_), .A3(new_n12049_), .ZN(new_n14654_));
  NOR4_X1    g11751(.A1(new_n14654_), .A2(new_n14652_), .A3(new_n12048_), .A4(new_n14609_), .ZN(new_n14655_));
  INV_X1     g11752(.I(new_n14609_), .ZN(new_n14656_));
  NAND2_X1   g11753(.A1(new_n12118_), .A2(pi0736), .ZN(new_n14657_));
  AND3_X2    g11754(.A1(new_n14657_), .A2(new_n14656_), .A3(new_n14630_), .Z(new_n14658_));
  NOR2_X1    g11755(.A1(new_n13649_), .A2(new_n14611_), .ZN(new_n14659_));
  NOR3_X1    g11756(.A1(new_n14659_), .A2(new_n14614_), .A3(new_n14629_), .ZN(new_n14660_));
  NAND2_X1   g11757(.A1(new_n14615_), .A2(pi0608), .ZN(new_n14661_));
  INV_X1     g11758(.I(new_n14658_), .ZN(new_n14662_));
  NOR2_X1    g11759(.A1(new_n14662_), .A2(new_n14659_), .ZN(new_n14663_));
  NAND2_X1   g11760(.A1(new_n11893_), .A2(pi0608), .ZN(new_n14664_));
  OAI22_X1   g11761(.A1(new_n14660_), .A2(new_n14661_), .B1(new_n14663_), .B2(new_n14664_), .ZN(new_n14665_));
  MUX2_X1    g11762(.I0(new_n14665_), .I1(new_n14658_), .S(new_n11891_), .Z(new_n14666_));
  NOR3_X1    g11763(.A1(new_n14618_), .A2(new_n11903_), .A3(new_n11912_), .ZN(new_n14667_));
  NOR4_X1    g11764(.A1(new_n14630_), .A2(pi1155), .A3(new_n13010_), .A4(new_n14609_), .ZN(new_n14668_));
  NOR3_X1    g11765(.A1(new_n14667_), .A2(pi0660), .A3(new_n14668_), .ZN(new_n14669_));
  NOR4_X1    g11766(.A1(new_n14666_), .A2(new_n11903_), .A3(pi1155), .A4(new_n14617_), .ZN(new_n14670_));
  INV_X1     g11767(.I(new_n11937_), .ZN(new_n14671_));
  NOR2_X1    g11768(.A1(new_n14609_), .A2(new_n14671_), .ZN(new_n14672_));
  OAI21_X1   g11769(.A1(new_n14630_), .A2(new_n12997_), .B(new_n14672_), .ZN(new_n14673_));
  OAI21_X1   g11770(.A1(new_n14670_), .A2(new_n14673_), .B(pi0785), .ZN(new_n14674_));
  OAI22_X1   g11771(.A1(new_n14674_), .A2(new_n14669_), .B1(pi0785), .B2(new_n14666_), .ZN(new_n14675_));
  INV_X1     g11772(.I(new_n14675_), .ZN(new_n14676_));
  AOI21_X1   g11773(.A1(new_n14617_), .A2(new_n11938_), .B(new_n14609_), .ZN(new_n14677_));
  XOR2_X1    g11774(.A1(new_n14675_), .A2(new_n14677_), .Z(new_n14678_));
  NAND2_X1   g11775(.A1(new_n14678_), .A2(pi0618), .ZN(new_n14679_));
  XOR2_X1    g11776(.A1(new_n14679_), .A2(new_n14676_), .Z(new_n14680_));
  NAND4_X1   g11777(.A1(new_n11924_), .A2(pi0618), .A3(new_n11950_), .A4(new_n14656_), .ZN(new_n14681_));
  OAI21_X1   g11778(.A1(new_n14632_), .A2(new_n14681_), .B(new_n11949_), .ZN(new_n14682_));
  AOI21_X1   g11779(.A1(new_n14680_), .A2(new_n11950_), .B(new_n14682_), .ZN(new_n14683_));
  XOR2_X1    g11780(.A1(new_n14679_), .A2(new_n14677_), .Z(new_n14684_));
  NOR2_X1    g11781(.A1(new_n14684_), .A2(new_n11950_), .ZN(new_n14685_));
  NAND2_X1   g11782(.A1(new_n11924_), .A2(new_n11934_), .ZN(new_n14686_));
  INV_X1     g11783(.I(new_n11960_), .ZN(new_n14687_));
  NOR2_X1    g11784(.A1(new_n14609_), .A2(new_n14687_), .ZN(new_n14688_));
  OAI21_X1   g11785(.A1(new_n14632_), .A2(new_n14686_), .B(new_n14688_), .ZN(new_n14689_));
  OAI21_X1   g11786(.A1(new_n14685_), .A2(new_n14689_), .B(pi0781), .ZN(new_n14690_));
  OAI22_X1   g11787(.A1(new_n14690_), .A2(new_n14683_), .B1(pi0781), .B2(new_n14676_), .ZN(new_n14691_));
  AOI21_X1   g11788(.A1(new_n14618_), .A2(new_n13716_), .B(new_n14609_), .ZN(new_n14692_));
  INV_X1     g11789(.I(new_n14692_), .ZN(new_n14693_));
  XOR2_X1    g11790(.A1(new_n14691_), .A2(new_n14693_), .Z(new_n14694_));
  NAND2_X1   g11791(.A1(new_n14694_), .A2(pi0619), .ZN(new_n14695_));
  XNOR2_X1   g11792(.A1(new_n14695_), .A2(new_n14691_), .ZN(new_n14696_));
  NOR3_X1    g11793(.A1(new_n14636_), .A2(new_n11914_), .A3(new_n11967_), .ZN(new_n14697_));
  AND2_X2    g11794(.A1(new_n14631_), .A2(new_n14697_), .Z(new_n14698_));
  NAND2_X1   g11795(.A1(new_n14656_), .A2(pi1159), .ZN(new_n14699_));
  OAI21_X1   g11796(.A1(new_n14698_), .A2(new_n14699_), .B(new_n11966_), .ZN(new_n14700_));
  AOI21_X1   g11797(.A1(new_n14696_), .A2(new_n11869_), .B(new_n14700_), .ZN(new_n14701_));
  NOR3_X1    g11798(.A1(new_n14636_), .A2(new_n11914_), .A3(pi0619), .ZN(new_n14702_));
  NAND2_X1   g11799(.A1(new_n14656_), .A2(new_n11869_), .ZN(new_n14703_));
  AOI21_X1   g11800(.A1(new_n14631_), .A2(new_n14702_), .B(new_n14703_), .ZN(new_n14704_));
  XOR2_X1    g11801(.A1(new_n14695_), .A2(new_n14693_), .Z(new_n14705_));
  NOR2_X1    g11802(.A1(new_n14705_), .A2(new_n11869_), .ZN(new_n14706_));
  NOR2_X1    g11803(.A1(pi0648), .A2(pi0789), .ZN(new_n14707_));
  OAI21_X1   g11804(.A1(new_n14706_), .A2(new_n14704_), .B(new_n14707_), .ZN(new_n14708_));
  AOI21_X1   g11805(.A1(new_n14691_), .A2(new_n11985_), .B(new_n11999_), .ZN(new_n14709_));
  OAI21_X1   g11806(.A1(new_n14708_), .A2(new_n14701_), .B(new_n14709_), .ZN(new_n14710_));
  NOR2_X1    g11807(.A1(new_n12014_), .A2(new_n14609_), .ZN(new_n14711_));
  NOR3_X1    g11808(.A1(new_n11987_), .A2(pi0626), .A3(pi0641), .ZN(new_n14712_));
  NAND4_X1   g11809(.A1(new_n11986_), .A2(new_n11987_), .A3(pi0626), .A4(pi0641), .ZN(new_n14714_));
  NOR4_X1    g11810(.A1(new_n14693_), .A2(new_n14711_), .A3(new_n14712_), .A4(new_n14714_), .ZN(new_n14715_));
  INV_X1     g11811(.I(new_n14646_), .ZN(new_n14716_));
  OAI21_X1   g11812(.A1(new_n14716_), .A2(pi0628), .B(new_n12051_), .ZN(new_n14717_));
  AOI21_X1   g11813(.A1(new_n14619_), .A2(pi0628), .B(new_n14717_), .ZN(new_n14718_));
  NAND2_X1   g11814(.A1(new_n14620_), .A2(pi0628), .ZN(new_n14719_));
  OAI21_X1   g11815(.A1(new_n14716_), .A2(new_n12031_), .B(new_n12030_), .ZN(new_n14720_));
  AOI21_X1   g11816(.A1(new_n14719_), .A2(new_n14720_), .B(pi1156), .ZN(new_n14721_));
  OAI21_X1   g11817(.A1(new_n14721_), .A2(new_n14718_), .B(new_n14656_), .ZN(new_n14722_));
  AOI21_X1   g11818(.A1(new_n14722_), .A2(pi0792), .B(new_n14715_), .ZN(new_n14723_));
  XNOR2_X1   g11819(.A1(pi0630), .A2(pi0647), .ZN(new_n14724_));
  AOI21_X1   g11820(.A1(new_n12090_), .A2(new_n14724_), .B(new_n12048_), .ZN(new_n14725_));
  INV_X1     g11821(.I(new_n14725_), .ZN(new_n14726_));
  INV_X1     g11822(.I(new_n12065_), .ZN(new_n14727_));
  NOR2_X1    g11823(.A1(new_n12031_), .A2(pi0629), .ZN(new_n14728_));
  NOR2_X1    g11824(.A1(new_n12030_), .A2(pi0628), .ZN(new_n14729_));
  NOR3_X1    g11825(.A1(new_n14727_), .A2(new_n14728_), .A3(new_n14729_), .ZN(new_n14730_));
  NOR2_X1    g11826(.A1(new_n14730_), .A2(new_n11868_), .ZN(new_n14731_));
  INV_X1     g11827(.I(new_n14731_), .ZN(new_n14732_));
  OAI21_X1   g11828(.A1(new_n14722_), .A2(new_n14732_), .B(new_n14726_), .ZN(new_n14733_));
  AOI21_X1   g11829(.A1(new_n14710_), .A2(new_n14723_), .B(new_n14733_), .ZN(new_n14734_));
  NOR2_X1    g11830(.A1(new_n14734_), .A2(new_n14655_), .ZN(new_n14735_));
  NOR3_X1    g11831(.A1(new_n14735_), .A2(pi0644), .A3(new_n14623_), .ZN(new_n14736_));
  AOI21_X1   g11832(.A1(new_n14735_), .A2(new_n12082_), .B(new_n14622_), .ZN(new_n14737_));
  INV_X1     g11833(.I(new_n14647_), .ZN(new_n14738_));
  NOR2_X1    g11834(.A1(pi0644), .A2(pi0715), .ZN(new_n14739_));
  INV_X1     g11835(.I(new_n14739_), .ZN(new_n14740_));
  NOR4_X1    g11836(.A1(new_n14738_), .A2(new_n12091_), .A3(new_n14609_), .A4(new_n14740_), .ZN(new_n14741_));
  NOR4_X1    g11837(.A1(new_n14736_), .A2(new_n14737_), .A3(new_n13169_), .A4(new_n14741_), .ZN(new_n14742_));
  NOR3_X1    g11838(.A1(new_n14738_), .A2(new_n12082_), .A3(new_n12091_), .ZN(new_n14743_));
  NAND2_X1   g11839(.A1(new_n14656_), .A2(new_n12099_), .ZN(new_n14744_));
  OAI21_X1   g11840(.A1(new_n14743_), .A2(new_n14744_), .B(new_n12081_), .ZN(new_n14745_));
  NAND2_X1   g11841(.A1(new_n14745_), .A2(pi0790), .ZN(new_n14746_));
  NOR2_X1    g11842(.A1(new_n11867_), .A2(pi0832), .ZN(new_n14747_));
  INV_X1     g11843(.I(new_n14747_), .ZN(new_n14748_));
  NOR3_X1    g11844(.A1(new_n14734_), .A2(new_n14655_), .A3(new_n14748_), .ZN(new_n14749_));
  OAI21_X1   g11845(.A1(new_n14742_), .A2(new_n14746_), .B(new_n14749_), .ZN(new_n14750_));
  NAND2_X1   g11846(.A1(new_n3232_), .A2(pi0144), .ZN(new_n14751_));
  NOR2_X1    g11847(.A1(new_n11875_), .A2(new_n14628_), .ZN(new_n14752_));
  INV_X1     g11848(.I(new_n14752_), .ZN(new_n14753_));
  NOR3_X1    g11849(.A1(new_n13368_), .A2(pi0144), .A3(new_n14753_), .ZN(new_n14754_));
  AOI21_X1   g11850(.A1(new_n12828_), .A2(new_n14753_), .B(new_n7504_), .ZN(new_n14755_));
  OAI21_X1   g11851(.A1(new_n14754_), .A2(new_n14755_), .B(pi0038), .ZN(new_n14756_));
  NOR2_X1    g11852(.A1(new_n14628_), .A2(pi0144), .ZN(new_n14757_));
  NOR2_X1    g11853(.A1(new_n12894_), .A2(pi0758), .ZN(new_n14758_));
  INV_X1     g11854(.I(new_n12823_), .ZN(new_n14759_));
  OAI21_X1   g11855(.A1(new_n14759_), .A2(new_n14628_), .B(pi0039), .ZN(new_n14760_));
  AOI21_X1   g11856(.A1(new_n14628_), .A2(new_n12697_), .B(new_n12664_), .ZN(new_n14761_));
  NOR3_X1    g11857(.A1(new_n13346_), .A2(new_n12697_), .A3(pi0758), .ZN(new_n14762_));
  NOR3_X1    g11858(.A1(new_n14761_), .A2(pi0039), .A3(new_n14762_), .ZN(new_n14763_));
  OAI21_X1   g11859(.A1(new_n14760_), .A2(new_n14758_), .B(new_n14763_), .ZN(new_n14764_));
  AOI22_X1   g11860(.A1(new_n14764_), .A2(pi0144), .B1(new_n14362_), .B2(new_n14757_), .ZN(new_n14765_));
  OAI21_X1   g11861(.A1(new_n14765_), .A2(pi0038), .B(new_n14756_), .ZN(new_n14766_));
  INV_X1     g11862(.I(new_n12277_), .ZN(new_n14767_));
  NOR4_X1    g11863(.A1(new_n12349_), .A2(pi0039), .A3(pi0144), .A4(pi0758), .ZN(new_n14768_));
  OAI21_X1   g11864(.A1(pi0144), .A2(new_n14767_), .B(new_n14768_), .ZN(new_n14769_));
  NOR2_X1    g11865(.A1(new_n7504_), .A2(new_n14628_), .ZN(new_n14770_));
  NAND3_X1   g11866(.A1(new_n14769_), .A2(new_n13332_), .A3(new_n14770_), .ZN(new_n14771_));
  AOI21_X1   g11867(.A1(new_n13362_), .A2(pi0144), .B(pi0758), .ZN(new_n14772_));
  OAI21_X1   g11868(.A1(pi0144), .A2(new_n13360_), .B(new_n14772_), .ZN(new_n14773_));
  NOR4_X1    g11869(.A1(new_n12668_), .A2(new_n7504_), .A3(pi0758), .A4(new_n13347_), .ZN(new_n14774_));
  NOR2_X1    g11870(.A1(new_n14774_), .A2(pi0039), .ZN(new_n14775_));
  NAND2_X1   g11871(.A1(new_n14773_), .A2(new_n14775_), .ZN(new_n14776_));
  NAND3_X1   g11872(.A1(new_n14756_), .A2(pi0736), .A3(new_n14352_), .ZN(new_n14777_));
  NOR2_X1    g11873(.A1(new_n3231_), .A2(pi0038), .ZN(new_n14778_));
  NAND4_X1   g11874(.A1(new_n14776_), .A2(new_n14771_), .A3(new_n14777_), .A4(new_n14778_), .ZN(new_n14779_));
  NAND3_X1   g11875(.A1(new_n14779_), .A2(new_n14766_), .A3(new_n14611_), .ZN(new_n14780_));
  NAND2_X1   g11876(.A1(new_n14780_), .A2(new_n14751_), .ZN(new_n14781_));
  NAND3_X1   g11877(.A1(new_n14780_), .A2(pi0625), .A3(new_n14751_), .ZN(new_n14782_));
  NOR2_X1    g11878(.A1(new_n3231_), .A2(pi0144), .ZN(new_n14783_));
  AOI21_X1   g11879(.A1(new_n14766_), .A2(new_n3231_), .B(new_n14783_), .ZN(new_n14784_));
  AOI21_X1   g11880(.A1(new_n14784_), .A2(new_n12970_), .B(pi1153), .ZN(new_n14785_));
  NAND2_X1   g11881(.A1(new_n14782_), .A2(new_n14785_), .ZN(new_n14786_));
  NOR3_X1    g11882(.A1(new_n13399_), .A2(pi0144), .A3(new_n13396_), .ZN(new_n14787_));
  AOI21_X1   g11883(.A1(new_n7504_), .A2(new_n13396_), .B(new_n14382_), .ZN(new_n14788_));
  NOR3_X1    g11884(.A1(new_n3232_), .A2(pi0038), .A3(new_n14611_), .ZN(new_n14791_));
  INV_X1     g11885(.I(new_n14791_), .ZN(new_n14792_));
  NOR3_X1    g11886(.A1(new_n14788_), .A2(new_n14787_), .A3(new_n14792_), .ZN(new_n14793_));
  AOI22_X1   g11887(.A1(new_n14396_), .A2(pi0144), .B1(pi0736), .B2(new_n3231_), .ZN(new_n14794_));
  OAI21_X1   g11888(.A1(new_n14793_), .A2(new_n14794_), .B(new_n12970_), .ZN(new_n14795_));
  NOR2_X1    g11889(.A1(new_n12965_), .A2(new_n7504_), .ZN(new_n14796_));
  NOR2_X1    g11890(.A1(new_n14796_), .A2(new_n12970_), .ZN(new_n14797_));
  NOR2_X1    g11891(.A1(new_n14797_), .A2(pi1153), .ZN(new_n14798_));
  AOI21_X1   g11892(.A1(new_n14798_), .A2(new_n14795_), .B(new_n13657_), .ZN(new_n14799_));
  NOR3_X1    g11893(.A1(new_n14793_), .A2(new_n14794_), .A3(new_n12970_), .ZN(new_n14800_));
  OAI21_X1   g11894(.A1(new_n14800_), .A2(new_n14797_), .B(pi1153), .ZN(new_n14801_));
  INV_X1     g11895(.I(new_n14781_), .ZN(new_n14802_));
  OAI21_X1   g11896(.A1(new_n14784_), .A2(new_n12970_), .B(new_n12977_), .ZN(new_n14803_));
  AOI21_X1   g11897(.A1(new_n14802_), .A2(pi0625), .B(new_n14803_), .ZN(new_n14804_));
  AOI22_X1   g11898(.A1(new_n14804_), .A2(new_n14801_), .B1(new_n14786_), .B2(new_n14799_), .ZN(new_n14805_));
  NOR3_X1    g11899(.A1(new_n14805_), .A2(new_n11891_), .A3(new_n14781_), .ZN(new_n14806_));
  AOI21_X1   g11900(.A1(new_n14805_), .A2(pi0778), .B(new_n14802_), .ZN(new_n14807_));
  NOR3_X1    g11901(.A1(new_n14806_), .A2(new_n14807_), .A3(pi0785), .ZN(new_n14808_));
  INV_X1     g11902(.I(new_n14808_), .ZN(new_n14809_));
  NOR2_X1    g11903(.A1(new_n14793_), .A2(new_n14794_), .ZN(new_n14810_));
  INV_X1     g11904(.I(new_n14810_), .ZN(new_n14811_));
  NAND2_X1   g11905(.A1(new_n14798_), .A2(new_n14795_), .ZN(new_n14812_));
  NAND2_X1   g11906(.A1(new_n14801_), .A2(new_n14812_), .ZN(new_n14813_));
  NAND3_X1   g11907(.A1(new_n14813_), .A2(pi0778), .A3(new_n14811_), .ZN(new_n14814_));
  OAI21_X1   g11908(.A1(new_n14813_), .A2(new_n11891_), .B(new_n14810_), .ZN(new_n14815_));
  NAND2_X1   g11909(.A1(new_n14815_), .A2(new_n14814_), .ZN(new_n14816_));
  AOI21_X1   g11910(.A1(new_n14816_), .A2(new_n11903_), .B(new_n11912_), .ZN(new_n14817_));
  INV_X1     g11911(.I(new_n14817_), .ZN(new_n14818_));
  NAND2_X1   g11912(.A1(new_n14396_), .A2(pi0144), .ZN(new_n14819_));
  NOR2_X1    g11913(.A1(new_n14819_), .A2(new_n11924_), .ZN(new_n14820_));
  AOI21_X1   g11914(.A1(new_n14784_), .A2(new_n11924_), .B(new_n14820_), .ZN(new_n14821_));
  MUX2_X1    g11915(.I0(new_n14821_), .I1(new_n14819_), .S(pi0609), .Z(new_n14822_));
  NOR2_X1    g11916(.A1(new_n14822_), .A2(pi1155), .ZN(new_n14823_));
  OAI21_X1   g11917(.A1(new_n14823_), .A2(new_n11923_), .B(pi0609), .ZN(new_n14824_));
  NOR3_X1    g11918(.A1(new_n14806_), .A2(new_n14807_), .A3(new_n14824_), .ZN(new_n14825_));
  AND2_X2    g11919(.A1(new_n14782_), .A2(new_n14785_), .Z(new_n14826_));
  INV_X1     g11920(.I(new_n14799_), .ZN(new_n14827_));
  INV_X1     g11921(.I(new_n14801_), .ZN(new_n14828_));
  INV_X1     g11922(.I(new_n14756_), .ZN(new_n14829_));
  NAND2_X1   g11923(.A1(new_n14362_), .A2(new_n14757_), .ZN(new_n14830_));
  NAND2_X1   g11924(.A1(new_n14764_), .A2(pi0144), .ZN(new_n14831_));
  NAND2_X1   g11925(.A1(new_n14831_), .A2(new_n14830_), .ZN(new_n14832_));
  AOI21_X1   g11926(.A1(new_n14832_), .A2(new_n3172_), .B(new_n14829_), .ZN(new_n14833_));
  INV_X1     g11927(.I(new_n14783_), .ZN(new_n14834_));
  OAI21_X1   g11928(.A1(new_n14833_), .A2(new_n3232_), .B(new_n14834_), .ZN(new_n14835_));
  NAND2_X1   g11929(.A1(new_n14835_), .A2(pi0625), .ZN(new_n14836_));
  NAND3_X1   g11930(.A1(new_n14836_), .A2(new_n14782_), .A3(new_n12977_), .ZN(new_n14837_));
  OAI22_X1   g11931(.A1(new_n14826_), .A2(new_n14827_), .B1(new_n14837_), .B2(new_n14828_), .ZN(new_n14838_));
  NAND3_X1   g11932(.A1(new_n14838_), .A2(pi0778), .A3(new_n14802_), .ZN(new_n14839_));
  OAI21_X1   g11933(.A1(new_n14838_), .A2(new_n11891_), .B(new_n14781_), .ZN(new_n14840_));
  NAND3_X1   g11934(.A1(new_n14840_), .A2(new_n14839_), .A3(new_n11903_), .ZN(new_n14841_));
  NOR2_X1    g11935(.A1(new_n11923_), .A2(pi1155), .ZN(new_n14844_));
  INV_X1     g11936(.I(new_n14844_), .ZN(new_n14845_));
  AOI21_X1   g11937(.A1(new_n14816_), .A2(pi0609), .B(new_n14845_), .ZN(new_n14846_));
  AOI22_X1   g11938(.A1(new_n14825_), .A2(new_n14818_), .B1(new_n14841_), .B2(new_n14846_), .ZN(new_n14847_));
  NOR3_X1    g11939(.A1(new_n14847_), .A2(new_n11870_), .A3(new_n14809_), .ZN(new_n14848_));
  NOR4_X1    g11940(.A1(new_n14784_), .A2(new_n11903_), .A3(new_n11914_), .A4(new_n14819_), .ZN(new_n14849_));
  AOI21_X1   g11941(.A1(pi0609), .A2(new_n14819_), .B(new_n14821_), .ZN(new_n14850_));
  OAI21_X1   g11942(.A1(new_n14850_), .A2(new_n14849_), .B(new_n11912_), .ZN(new_n14851_));
  NAND2_X1   g11943(.A1(new_n14851_), .A2(pi0660), .ZN(new_n14852_));
  NAND4_X1   g11944(.A1(new_n14840_), .A2(new_n14839_), .A3(pi0609), .A4(new_n14852_), .ZN(new_n14853_));
  NOR3_X1    g11945(.A1(new_n14806_), .A2(new_n14807_), .A3(pi0609), .ZN(new_n14854_));
  INV_X1     g11946(.I(new_n14846_), .ZN(new_n14855_));
  OAI22_X1   g11947(.A1(new_n14854_), .A2(new_n14855_), .B1(new_n14853_), .B2(new_n14817_), .ZN(new_n14856_));
  AOI21_X1   g11948(.A1(new_n14856_), .A2(pi0785), .B(new_n14808_), .ZN(new_n14857_));
  NOR3_X1    g11949(.A1(new_n14857_), .A2(new_n14848_), .A3(pi0781), .ZN(new_n14858_));
  INV_X1     g11950(.I(new_n14858_), .ZN(new_n14859_));
  INV_X1     g11951(.I(new_n14820_), .ZN(new_n14860_));
  OAI21_X1   g11952(.A1(new_n14835_), .A2(new_n11914_), .B(new_n14860_), .ZN(new_n14861_));
  NOR3_X1    g11953(.A1(new_n14821_), .A2(new_n11903_), .A3(new_n14796_), .ZN(new_n14862_));
  AOI21_X1   g11954(.A1(new_n14821_), .A2(pi0609), .B(new_n14819_), .ZN(new_n14863_));
  OAI21_X1   g11955(.A1(new_n14862_), .A2(new_n14863_), .B(pi1155), .ZN(new_n14864_));
  NAND2_X1   g11956(.A1(new_n14851_), .A2(new_n14864_), .ZN(new_n14865_));
  MUX2_X1    g11957(.I0(new_n14865_), .I1(new_n14861_), .S(new_n11870_), .Z(new_n14866_));
  NAND3_X1   g11958(.A1(new_n14866_), .A2(new_n11934_), .A3(new_n14796_), .ZN(new_n14867_));
  OAI21_X1   g11959(.A1(new_n14866_), .A2(pi0618), .B(new_n14819_), .ZN(new_n14868_));
  NAND3_X1   g11960(.A1(new_n14868_), .A2(new_n14867_), .A3(new_n11950_), .ZN(new_n14869_));
  NOR2_X1    g11961(.A1(new_n14869_), .A2(new_n11949_), .ZN(new_n14870_));
  INV_X1     g11962(.I(new_n14870_), .ZN(new_n14871_));
  NOR2_X1    g11963(.A1(new_n14816_), .A2(new_n13024_), .ZN(new_n14872_));
  AOI21_X1   g11964(.A1(new_n13024_), .A2(new_n14796_), .B(new_n14872_), .ZN(new_n14873_));
  NOR4_X1    g11965(.A1(new_n14857_), .A2(new_n14848_), .A3(new_n11934_), .A4(pi1154), .ZN(new_n14874_));
  NAND3_X1   g11966(.A1(new_n14856_), .A2(pi0785), .A3(new_n14808_), .ZN(new_n14875_));
  OAI21_X1   g11967(.A1(new_n14847_), .A2(new_n11870_), .B(new_n14809_), .ZN(new_n14876_));
  NAND3_X1   g11968(.A1(new_n14875_), .A2(new_n14876_), .A3(new_n11934_), .ZN(new_n14877_));
  AOI21_X1   g11969(.A1(new_n14873_), .A2(pi0618), .B(new_n14687_), .ZN(new_n14878_));
  AOI22_X1   g11970(.A1(new_n14874_), .A2(new_n14871_), .B1(new_n14877_), .B2(new_n14878_), .ZN(new_n14879_));
  NOR3_X1    g11971(.A1(new_n14879_), .A2(new_n11969_), .A3(new_n14859_), .ZN(new_n14880_));
  NAND4_X1   g11972(.A1(new_n14875_), .A2(new_n14876_), .A3(pi0618), .A4(new_n11950_), .ZN(new_n14881_));
  NOR3_X1    g11973(.A1(new_n14857_), .A2(new_n14848_), .A3(pi0618), .ZN(new_n14882_));
  INV_X1     g11974(.I(new_n14878_), .ZN(new_n14883_));
  OAI22_X1   g11975(.A1(new_n14870_), .A2(new_n14881_), .B1(new_n14882_), .B2(new_n14883_), .ZN(new_n14884_));
  AOI21_X1   g11976(.A1(new_n14884_), .A2(pi0781), .B(new_n14858_), .ZN(new_n14885_));
  NOR3_X1    g11977(.A1(new_n14885_), .A2(new_n14880_), .A3(pi0789), .ZN(new_n14886_));
  INV_X1     g11978(.I(new_n14886_), .ZN(new_n14887_));
  NAND3_X1   g11979(.A1(new_n14861_), .A2(pi0609), .A3(new_n14819_), .ZN(new_n14888_));
  INV_X1     g11980(.I(new_n14863_), .ZN(new_n14889_));
  AOI21_X1   g11981(.A1(new_n14889_), .A2(new_n14888_), .B(new_n11912_), .ZN(new_n14890_));
  NOR2_X1    g11982(.A1(new_n14890_), .A2(new_n14823_), .ZN(new_n14891_));
  MUX2_X1    g11983(.I0(new_n14891_), .I1(new_n14821_), .S(new_n11870_), .Z(new_n14892_));
  MUX2_X1    g11984(.I0(new_n14869_), .I1(new_n14892_), .S(new_n11969_), .Z(new_n14893_));
  NOR3_X1    g11985(.A1(new_n14893_), .A2(pi0619), .A3(new_n14819_), .ZN(new_n14894_));
  AOI21_X1   g11986(.A1(new_n14893_), .A2(new_n11967_), .B(new_n14796_), .ZN(new_n14895_));
  NOR4_X1    g11987(.A1(new_n14894_), .A2(new_n14895_), .A3(new_n11966_), .A4(pi1159), .ZN(new_n14896_));
  INV_X1     g11988(.I(new_n14896_), .ZN(new_n14897_));
  NOR2_X1    g11989(.A1(new_n14796_), .A2(new_n11961_), .ZN(new_n14898_));
  AOI21_X1   g11990(.A1(new_n14873_), .A2(new_n11961_), .B(new_n14898_), .ZN(new_n14899_));
  NOR4_X1    g11991(.A1(new_n14885_), .A2(new_n14880_), .A3(new_n11967_), .A4(pi1159), .ZN(new_n14900_));
  NAND3_X1   g11992(.A1(new_n14884_), .A2(pi0781), .A3(new_n14858_), .ZN(new_n14901_));
  OAI21_X1   g11993(.A1(new_n14879_), .A2(new_n11969_), .B(new_n14859_), .ZN(new_n14902_));
  NAND3_X1   g11994(.A1(new_n14901_), .A2(new_n14902_), .A3(new_n11967_), .ZN(new_n14903_));
  INV_X1     g11995(.I(new_n12011_), .ZN(new_n14904_));
  INV_X1     g11996(.I(new_n14899_), .ZN(new_n14905_));
  AOI21_X1   g11997(.A1(new_n14905_), .A2(pi0619), .B(new_n14904_), .ZN(new_n14906_));
  AOI22_X1   g11998(.A1(new_n14900_), .A2(new_n14897_), .B1(new_n14903_), .B2(new_n14906_), .ZN(new_n14907_));
  NOR3_X1    g11999(.A1(new_n14907_), .A2(new_n11985_), .A3(new_n14887_), .ZN(new_n14908_));
  NOR2_X1    g12000(.A1(new_n11967_), .A2(pi1159), .ZN(new_n14909_));
  NAND3_X1   g12001(.A1(new_n14901_), .A2(new_n14902_), .A3(new_n14909_), .ZN(new_n14910_));
  NOR3_X1    g12002(.A1(new_n14885_), .A2(new_n14880_), .A3(pi0619), .ZN(new_n14911_));
  INV_X1     g12003(.I(new_n14906_), .ZN(new_n14912_));
  OAI22_X1   g12004(.A1(new_n14911_), .A2(new_n14912_), .B1(new_n14910_), .B2(new_n14896_), .ZN(new_n14913_));
  AOI21_X1   g12005(.A1(new_n14913_), .A2(pi0789), .B(new_n14886_), .ZN(new_n14914_));
  NOR2_X1    g12006(.A1(new_n14908_), .A2(new_n14914_), .ZN(new_n14915_));
  INV_X1     g12007(.I(new_n14915_), .ZN(new_n14916_));
  NOR3_X1    g12008(.A1(new_n14892_), .A2(pi0618), .A3(new_n14819_), .ZN(new_n14917_));
  AOI21_X1   g12009(.A1(new_n14892_), .A2(new_n11934_), .B(new_n14796_), .ZN(new_n14918_));
  NOR3_X1    g12010(.A1(new_n14917_), .A2(new_n14918_), .A3(pi1154), .ZN(new_n14919_));
  MUX2_X1    g12011(.I0(new_n14919_), .I1(new_n14866_), .S(new_n11969_), .Z(new_n14920_));
  NOR3_X1    g12012(.A1(new_n14894_), .A2(new_n14895_), .A3(pi1159), .ZN(new_n14921_));
  MUX2_X1    g12013(.I0(new_n14921_), .I1(new_n14920_), .S(new_n11985_), .Z(new_n14922_));
  NAND3_X1   g12014(.A1(new_n14922_), .A2(new_n11994_), .A3(new_n14796_), .ZN(new_n14923_));
  OAI21_X1   g12015(.A1(new_n14922_), .A2(pi0626), .B(new_n14819_), .ZN(new_n14924_));
  NAND4_X1   g12016(.A1(new_n14924_), .A2(new_n14923_), .A3(pi0641), .A4(new_n11987_), .ZN(new_n14925_));
  INV_X1     g12017(.I(new_n14925_), .ZN(new_n14926_));
  NAND3_X1   g12018(.A1(new_n14913_), .A2(pi0789), .A3(new_n14886_), .ZN(new_n14927_));
  OAI21_X1   g12019(.A1(new_n14907_), .A2(new_n11985_), .B(new_n14887_), .ZN(new_n14928_));
  NOR2_X1    g12020(.A1(new_n14819_), .A2(new_n12014_), .ZN(new_n14929_));
  AOI21_X1   g12021(.A1(new_n14899_), .A2(new_n12014_), .B(new_n14929_), .ZN(new_n14930_));
  NOR2_X1    g12022(.A1(new_n11989_), .A2(pi0626), .ZN(new_n14931_));
  INV_X1     g12023(.I(new_n14931_), .ZN(new_n14932_));
  AOI21_X1   g12024(.A1(new_n14928_), .A2(new_n14927_), .B(new_n14932_), .ZN(new_n14933_));
  NOR2_X1    g12025(.A1(new_n11994_), .A2(pi0641), .ZN(new_n14934_));
  INV_X1     g12026(.I(new_n14934_), .ZN(new_n14935_));
  AOI21_X1   g12027(.A1(new_n14928_), .A2(new_n14927_), .B(new_n14935_), .ZN(new_n14936_));
  NOR4_X1    g12028(.A1(new_n14933_), .A2(new_n14936_), .A3(new_n14926_), .A4(new_n13095_), .ZN(new_n14937_));
  NOR3_X1    g12029(.A1(new_n14937_), .A2(new_n11986_), .A3(new_n14916_), .ZN(new_n14938_));
  AOI21_X1   g12030(.A1(new_n14937_), .A2(pi0788), .B(new_n14915_), .ZN(new_n14939_));
  NOR2_X1    g12031(.A1(new_n14938_), .A2(new_n14939_), .ZN(new_n14940_));
  NAND3_X1   g12032(.A1(new_n14920_), .A2(new_n11967_), .A3(new_n14796_), .ZN(new_n14941_));
  OAI21_X1   g12033(.A1(new_n14920_), .A2(pi0619), .B(new_n14819_), .ZN(new_n14942_));
  NAND3_X1   g12034(.A1(new_n14942_), .A2(new_n14941_), .A3(new_n11869_), .ZN(new_n14943_));
  MUX2_X1    g12035(.I0(new_n14943_), .I1(new_n14893_), .S(new_n11985_), .Z(new_n14944_));
  NOR3_X1    g12036(.A1(new_n14944_), .A2(pi0626), .A3(new_n14819_), .ZN(new_n14945_));
  AOI21_X1   g12037(.A1(new_n14944_), .A2(new_n11994_), .B(new_n14796_), .ZN(new_n14946_));
  NOR3_X1    g12038(.A1(new_n14945_), .A2(new_n14946_), .A3(pi1158), .ZN(new_n14947_));
  NOR2_X1    g12039(.A1(new_n14922_), .A2(pi0788), .ZN(new_n14948_));
  INV_X1     g12040(.I(new_n14948_), .ZN(new_n14949_));
  NOR3_X1    g12041(.A1(new_n14947_), .A2(new_n11986_), .A3(new_n14949_), .ZN(new_n14950_));
  NAND3_X1   g12042(.A1(new_n14924_), .A2(new_n14923_), .A3(new_n11987_), .ZN(new_n14951_));
  AOI21_X1   g12043(.A1(new_n14951_), .A2(pi0788), .B(new_n14948_), .ZN(new_n14952_));
  OAI21_X1   g12044(.A1(new_n14950_), .A2(new_n14952_), .B(new_n12031_), .ZN(new_n14953_));
  NOR2_X1    g12045(.A1(new_n14796_), .A2(new_n13114_), .ZN(new_n14954_));
  AOI21_X1   g12046(.A1(new_n14930_), .A2(new_n13114_), .B(new_n14954_), .ZN(new_n14955_));
  INV_X1     g12047(.I(new_n14955_), .ZN(new_n14956_));
  NAND3_X1   g12048(.A1(new_n14956_), .A2(new_n12031_), .A3(new_n14796_), .ZN(new_n14957_));
  OAI21_X1   g12049(.A1(new_n14956_), .A2(pi0628), .B(new_n14819_), .ZN(new_n14958_));
  NAND3_X1   g12050(.A1(new_n14958_), .A2(new_n14957_), .A3(new_n12026_), .ZN(new_n14959_));
  INV_X1     g12051(.I(new_n14959_), .ZN(new_n14960_));
  AOI21_X1   g12052(.A1(new_n14960_), .A2(pi0629), .B(new_n12031_), .ZN(new_n14961_));
  INV_X1     g12053(.I(new_n14961_), .ZN(new_n14962_));
  AOI21_X1   g12054(.A1(new_n14953_), .A2(pi1156), .B(new_n14962_), .ZN(new_n14963_));
  NOR3_X1    g12055(.A1(new_n12030_), .A2(new_n12026_), .A3(pi0628), .ZN(new_n14965_));
  OAI22_X1   g12056(.A1(new_n14963_), .A2(new_n14965_), .B1(new_n14938_), .B2(new_n14939_), .ZN(new_n14966_));
  MUX2_X1    g12057(.I0(new_n14966_), .I1(new_n14940_), .S(new_n11868_), .Z(new_n14967_));
  INV_X1     g12058(.I(new_n14967_), .ZN(new_n14968_));
  OAI21_X1   g12059(.A1(new_n14950_), .A2(new_n14952_), .B(new_n12054_), .ZN(new_n14969_));
  OAI21_X1   g12060(.A1(new_n12054_), .A2(new_n14796_), .B(new_n14969_), .ZN(new_n14970_));
  NAND2_X1   g12061(.A1(new_n14970_), .A2(new_n12061_), .ZN(new_n14971_));
  MUX2_X1    g12062(.I0(new_n14960_), .I1(new_n14956_), .S(new_n11868_), .Z(new_n14972_));
  NAND3_X1   g12063(.A1(new_n14972_), .A2(new_n12061_), .A3(new_n14796_), .ZN(new_n14973_));
  OAI21_X1   g12064(.A1(new_n14972_), .A2(pi0647), .B(new_n14819_), .ZN(new_n14974_));
  NAND3_X1   g12065(.A1(new_n14974_), .A2(new_n14973_), .A3(new_n12049_), .ZN(new_n14975_));
  OAI21_X1   g12066(.A1(new_n14975_), .A2(new_n12060_), .B(pi0647), .ZN(new_n14976_));
  AOI21_X1   g12067(.A1(new_n14971_), .A2(pi1157), .B(new_n14976_), .ZN(new_n14977_));
  OAI21_X1   g12068(.A1(new_n14908_), .A2(new_n14914_), .B(new_n14931_), .ZN(new_n14978_));
  OAI21_X1   g12069(.A1(new_n14908_), .A2(new_n14914_), .B(new_n14934_), .ZN(new_n14979_));
  NAND4_X1   g12070(.A1(new_n14978_), .A2(new_n14979_), .A3(new_n12016_), .A4(new_n14925_), .ZN(new_n14980_));
  NAND3_X1   g12071(.A1(new_n14980_), .A2(pi0788), .A3(new_n14915_), .ZN(new_n14981_));
  OAI21_X1   g12072(.A1(new_n14980_), .A2(new_n11986_), .B(new_n14916_), .ZN(new_n14982_));
  NAND3_X1   g12073(.A1(new_n14951_), .A2(pi0788), .A3(new_n14948_), .ZN(new_n14983_));
  OAI21_X1   g12074(.A1(new_n14947_), .A2(new_n11986_), .B(new_n14949_), .ZN(new_n14984_));
  AOI21_X1   g12075(.A1(new_n14984_), .A2(new_n14983_), .B(pi0628), .ZN(new_n14985_));
  OAI21_X1   g12076(.A1(new_n14985_), .A2(new_n12026_), .B(new_n14961_), .ZN(new_n14986_));
  INV_X1     g12077(.I(new_n14965_), .ZN(new_n14987_));
  AOI22_X1   g12078(.A1(new_n14986_), .A2(new_n14987_), .B1(new_n14982_), .B2(new_n14981_), .ZN(new_n14988_));
  NAND3_X1   g12079(.A1(new_n14988_), .A2(pi0792), .A3(new_n14940_), .ZN(new_n14989_));
  NAND2_X1   g12080(.A1(new_n14982_), .A2(new_n14981_), .ZN(new_n14990_));
  OAI21_X1   g12081(.A1(new_n14988_), .A2(new_n11868_), .B(new_n14990_), .ZN(new_n14991_));
  NAND3_X1   g12082(.A1(new_n14991_), .A2(new_n14989_), .A3(new_n12061_), .ZN(new_n14992_));
  AOI21_X1   g12083(.A1(new_n14970_), .A2(pi0647), .B(new_n13743_), .ZN(new_n14993_));
  AOI22_X1   g12084(.A1(new_n14992_), .A2(new_n14993_), .B1(new_n14967_), .B2(new_n14977_), .ZN(new_n14994_));
  MUX2_X1    g12085(.I0(new_n14994_), .I1(new_n14968_), .S(new_n12048_), .Z(new_n14995_));
  NOR2_X1    g12086(.A1(new_n14970_), .A2(new_n12091_), .ZN(new_n14996_));
  AOI21_X1   g12087(.A1(new_n12091_), .A2(new_n14796_), .B(new_n14996_), .ZN(new_n14997_));
  NAND2_X1   g12088(.A1(new_n14997_), .A2(new_n12082_), .ZN(new_n14998_));
  AOI21_X1   g12089(.A1(new_n14819_), .A2(pi0644), .B(new_n12099_), .ZN(new_n14999_));
  NOR2_X1    g12090(.A1(new_n14972_), .A2(pi0787), .ZN(new_n15000_));
  NAND2_X1   g12091(.A1(new_n14975_), .A2(pi0787), .ZN(new_n15001_));
  XNOR2_X1   g12092(.A1(new_n15001_), .A2(new_n15000_), .ZN(new_n15002_));
  OAI21_X1   g12093(.A1(new_n15002_), .A2(new_n12082_), .B(new_n13168_), .ZN(new_n15003_));
  AOI21_X1   g12094(.A1(new_n14998_), .A2(new_n14999_), .B(new_n15003_), .ZN(new_n15004_));
  OAI21_X1   g12095(.A1(new_n14995_), .A2(pi0644), .B(new_n15004_), .ZN(new_n15005_));
  NAND2_X1   g12096(.A1(new_n14967_), .A2(new_n12048_), .ZN(new_n15006_));
  OR3_X2     g12097(.A1(new_n14994_), .A2(new_n12048_), .A3(new_n15006_), .Z(new_n15007_));
  OAI21_X1   g12098(.A1(new_n14994_), .A2(new_n12048_), .B(new_n15006_), .ZN(new_n15008_));
  NOR3_X1    g12099(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n15009_));
  NAND2_X1   g12100(.A1(new_n14997_), .A2(new_n15009_), .ZN(new_n15010_));
  NOR2_X1    g12101(.A1(new_n12082_), .A2(pi0715), .ZN(new_n15011_));
  NAND4_X1   g12102(.A1(new_n15007_), .A2(new_n15008_), .A3(new_n15010_), .A4(new_n15011_), .ZN(new_n15012_));
  OAI21_X1   g12103(.A1(new_n14995_), .A2(new_n5223_), .B(new_n11867_), .ZN(new_n15013_));
  AOI21_X1   g12104(.A1(new_n15005_), .A2(new_n15012_), .B(new_n15013_), .ZN(new_n15014_));
  NAND2_X1   g12105(.A1(pi0057), .A2(pi0144), .ZN(new_n15015_));
  AOI21_X1   g12106(.A1(new_n15015_), .A2(new_n13184_), .B(pi0057), .ZN(new_n15016_));
  OAI21_X1   g12107(.A1(new_n5224_), .A2(pi0144), .B(new_n15016_), .ZN(new_n15017_));
  OAI21_X1   g12108(.A1(new_n15014_), .A2(new_n15017_), .B(new_n14750_), .ZN(po0301));
  NOR2_X1    g12109(.A1(new_n2925_), .A2(pi0145), .ZN(new_n15019_));
  INV_X1     g12110(.I(new_n15019_), .ZN(new_n15020_));
  NAND2_X1   g12111(.A1(new_n12053_), .A2(new_n15020_), .ZN(new_n15021_));
  NOR2_X1    g12112(.A1(new_n11877_), .A2(pi0767), .ZN(new_n15022_));
  NOR2_X1    g12113(.A1(new_n15022_), .A2(new_n15019_), .ZN(new_n15023_));
  NOR2_X1    g12114(.A1(new_n15023_), .A2(new_n11925_), .ZN(new_n15024_));
  NOR2_X1    g12115(.A1(new_n15024_), .A2(pi0785), .ZN(new_n15025_));
  AOI21_X1   g12116(.A1(new_n15024_), .A2(new_n11928_), .B(pi1155), .ZN(new_n15026_));
  INV_X1     g12117(.I(new_n15023_), .ZN(new_n15027_));
  AOI21_X1   g12118(.A1(new_n15027_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n15028_));
  OAI21_X1   g12119(.A1(new_n15026_), .A2(new_n15028_), .B(pi0785), .ZN(new_n15029_));
  XNOR2_X1   g12120(.A1(new_n15029_), .A2(new_n15025_), .ZN(new_n15030_));
  NAND2_X1   g12121(.A1(new_n15030_), .A2(new_n11969_), .ZN(new_n15031_));
  INV_X1     g12122(.I(new_n15030_), .ZN(new_n15032_));
  OAI21_X1   g12123(.A1(new_n15032_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n15033_));
  NOR2_X1    g12124(.A1(new_n15032_), .A2(new_n11945_), .ZN(new_n15034_));
  OAI21_X1   g12125(.A1(new_n15033_), .A2(new_n15034_), .B(pi0781), .ZN(new_n15035_));
  XOR2_X1    g12126(.A1(new_n15035_), .A2(new_n15031_), .Z(new_n15036_));
  INV_X1     g12127(.I(new_n15036_), .ZN(new_n15037_));
  NOR2_X1    g12128(.A1(new_n15037_), .A2(pi0789), .ZN(new_n15038_));
  OAI21_X1   g12129(.A1(new_n15020_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n15039_));
  AOI21_X1   g12130(.A1(new_n15036_), .A2(pi0619), .B(new_n15039_), .ZN(new_n15040_));
  AOI21_X1   g12131(.A1(new_n15020_), .A2(new_n11967_), .B(pi1159), .ZN(new_n15041_));
  OAI21_X1   g12132(.A1(new_n15037_), .A2(new_n11967_), .B(new_n15041_), .ZN(new_n15042_));
  AOI21_X1   g12133(.A1(new_n15042_), .A2(new_n15040_), .B(new_n11985_), .ZN(new_n15043_));
  XOR2_X1    g12134(.A1(new_n15043_), .A2(new_n15038_), .Z(new_n15044_));
  INV_X1     g12135(.I(new_n15044_), .ZN(new_n15045_));
  MUX2_X1    g12136(.I0(new_n15045_), .I1(new_n15019_), .S(new_n12003_), .Z(new_n15046_));
  NAND2_X1   g12137(.A1(new_n15046_), .A2(pi0788), .ZN(new_n15047_));
  OAI21_X1   g12138(.A1(pi0788), .A2(new_n15044_), .B(new_n15047_), .ZN(new_n15048_));
  OAI21_X1   g12139(.A1(new_n15048_), .A2(new_n12053_), .B(new_n15021_), .ZN(new_n15049_));
  INV_X1     g12140(.I(new_n12068_), .ZN(new_n15050_));
  INV_X1     g12141(.I(pi0698), .ZN(new_n15051_));
  AOI21_X1   g12142(.A1(new_n11886_), .A2(new_n15051_), .B(new_n15019_), .ZN(new_n15052_));
  INV_X1     g12143(.I(new_n15052_), .ZN(new_n15053_));
  NOR3_X1    g12144(.A1(new_n11894_), .A2(pi0625), .A3(pi0698), .ZN(new_n15054_));
  XOR2_X1    g12145(.A1(new_n15054_), .A2(pi1153), .Z(new_n15055_));
  NAND2_X1   g12146(.A1(new_n15055_), .A2(new_n15053_), .ZN(new_n15056_));
  OAI21_X1   g12147(.A1(new_n15054_), .A2(new_n15019_), .B(new_n11893_), .ZN(new_n15057_));
  AOI21_X1   g12148(.A1(new_n15056_), .A2(new_n15057_), .B(new_n11891_), .ZN(new_n15058_));
  AOI21_X1   g12149(.A1(new_n11891_), .A2(new_n15053_), .B(new_n15058_), .ZN(new_n15059_));
  NOR2_X1    g12150(.A1(new_n15059_), .A2(new_n11939_), .ZN(new_n15060_));
  NAND2_X1   g12151(.A1(new_n15060_), .A2(new_n11963_), .ZN(new_n15061_));
  INV_X1     g12152(.I(new_n15061_), .ZN(new_n15062_));
  NOR2_X1    g12153(.A1(new_n15062_), .A2(new_n12034_), .ZN(new_n15063_));
  NAND2_X1   g12154(.A1(new_n15063_), .A2(new_n15050_), .ZN(new_n15064_));
  AOI21_X1   g12155(.A1(new_n15019_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n15065_));
  OAI21_X1   g12156(.A1(new_n15064_), .A2(new_n12061_), .B(new_n15065_), .ZN(new_n15066_));
  INV_X1     g12157(.I(new_n15066_), .ZN(new_n15067_));
  INV_X1     g12158(.I(new_n15064_), .ZN(new_n15068_));
  AOI21_X1   g12159(.A1(new_n15019_), .A2(pi0647), .B(pi1157), .ZN(new_n15069_));
  OAI21_X1   g12160(.A1(new_n15068_), .A2(new_n12061_), .B(new_n15069_), .ZN(new_n15070_));
  INV_X1     g12161(.I(new_n15070_), .ZN(new_n15071_));
  NAND2_X1   g12162(.A1(new_n15067_), .A2(new_n12060_), .ZN(new_n15072_));
  NOR2_X1    g12163(.A1(new_n15071_), .A2(new_n12060_), .ZN(new_n15073_));
  OAI21_X1   g12164(.A1(pi0630), .A2(new_n15066_), .B(new_n15073_), .ZN(new_n15074_));
  NAND2_X1   g12165(.A1(new_n13747_), .A2(pi0630), .ZN(new_n15075_));
  OAI21_X1   g12166(.A1(pi0630), .A2(new_n13737_), .B(new_n15075_), .ZN(new_n15076_));
  INV_X1     g12167(.I(new_n15076_), .ZN(new_n15077_));
  NOR2_X1    g12168(.A1(new_n15077_), .A2(pi0787), .ZN(new_n15078_));
  NAND4_X1   g12169(.A1(new_n15049_), .A2(new_n15072_), .A3(new_n15074_), .A4(new_n15078_), .ZN(new_n15079_));
  NOR2_X1    g12170(.A1(new_n13277_), .A2(pi1156), .ZN(new_n15080_));
  AOI22_X1   g12171(.A1(new_n15048_), .A2(new_n12064_), .B1(new_n15063_), .B2(new_n15080_), .ZN(new_n15081_));
  NOR2_X1    g12172(.A1(new_n15081_), .A2(new_n12030_), .ZN(new_n15082_));
  NAND2_X1   g12173(.A1(new_n15048_), .A2(new_n12063_), .ZN(new_n15083_));
  AOI21_X1   g12174(.A1(new_n2925_), .A2(new_n12031_), .B(new_n12026_), .ZN(new_n15084_));
  NOR2_X1    g12175(.A1(new_n12030_), .A2(pi0792), .ZN(new_n15085_));
  INV_X1     g12176(.I(new_n15085_), .ZN(new_n15086_));
  AOI21_X1   g12177(.A1(new_n15063_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n15087_));
  NAND2_X1   g12178(.A1(new_n15083_), .A2(new_n15087_), .ZN(new_n15088_));
  NOR2_X1    g12179(.A1(new_n15082_), .A2(new_n15088_), .ZN(new_n15089_));
  NOR2_X1    g12180(.A1(new_n15052_), .A2(new_n11874_), .ZN(new_n15090_));
  OAI21_X1   g12181(.A1(new_n15027_), .A2(new_n15090_), .B(new_n11891_), .ZN(new_n15091_));
  NAND2_X1   g12182(.A1(new_n15090_), .A2(pi0625), .ZN(new_n15092_));
  NOR4_X1    g12183(.A1(new_n15022_), .A2(pi0608), .A3(new_n11893_), .A4(new_n15019_), .ZN(new_n15093_));
  OAI21_X1   g12184(.A1(new_n15027_), .A2(new_n15090_), .B(new_n15092_), .ZN(new_n15094_));
  NOR3_X1    g12185(.A1(new_n15019_), .A2(pi0608), .A3(pi1153), .ZN(new_n15095_));
  AOI22_X1   g12186(.A1(new_n15094_), .A2(new_n15095_), .B1(new_n15092_), .B2(new_n15093_), .ZN(new_n15096_));
  NOR2_X1    g12187(.A1(new_n15096_), .A2(new_n11891_), .ZN(new_n15097_));
  XNOR2_X1   g12188(.A1(new_n15097_), .A2(new_n15091_), .ZN(new_n15098_));
  NOR2_X1    g12189(.A1(new_n15098_), .A2(pi0785), .ZN(new_n15099_));
  NOR3_X1    g12190(.A1(new_n15059_), .A2(new_n11903_), .A3(new_n11912_), .ZN(new_n15100_));
  NOR3_X1    g12191(.A1(new_n15100_), .A2(pi0660), .A3(new_n15028_), .ZN(new_n15101_));
  INV_X1     g12192(.I(new_n15059_), .ZN(new_n15102_));
  NOR4_X1    g12193(.A1(new_n15098_), .A2(new_n11903_), .A3(pi1155), .A4(new_n15102_), .ZN(new_n15103_));
  NOR3_X1    g12194(.A1(new_n15103_), .A2(new_n11923_), .A3(new_n15026_), .ZN(new_n15104_));
  NOR3_X1    g12195(.A1(new_n15104_), .A2(new_n11870_), .A3(new_n15101_), .ZN(new_n15105_));
  NOR2_X1    g12196(.A1(new_n15105_), .A2(new_n15099_), .ZN(new_n15106_));
  NOR2_X1    g12197(.A1(new_n15106_), .A2(pi0781), .ZN(new_n15107_));
  NOR4_X1    g12198(.A1(new_n15059_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n15108_));
  OAI21_X1   g12199(.A1(new_n15032_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n15109_));
  NOR4_X1    g12200(.A1(new_n15106_), .A2(new_n11934_), .A3(pi1154), .A4(new_n15060_), .ZN(new_n15110_));
  NOR2_X1    g12201(.A1(new_n15110_), .A2(new_n15033_), .ZN(new_n15111_));
  OAI22_X1   g12202(.A1(new_n15111_), .A2(pi0627), .B1(new_n15108_), .B2(new_n15109_), .ZN(new_n15112_));
  AOI21_X1   g12203(.A1(new_n15112_), .A2(pi0781), .B(new_n15107_), .ZN(new_n15113_));
  NOR4_X1    g12204(.A1(new_n15113_), .A2(new_n11967_), .A3(pi1159), .A4(new_n15062_), .ZN(new_n15114_));
  NAND2_X1   g12205(.A1(new_n15040_), .A2(pi0648), .ZN(new_n15115_));
  NOR3_X1    g12206(.A1(new_n15061_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n15116_));
  NAND2_X1   g12207(.A1(new_n15042_), .A2(new_n11966_), .ZN(new_n15117_));
  OAI22_X1   g12208(.A1(new_n15114_), .A2(new_n15115_), .B1(new_n15116_), .B2(new_n15117_), .ZN(new_n15118_));
  AOI21_X1   g12209(.A1(new_n15113_), .A2(new_n11998_), .B(pi0789), .ZN(new_n15119_));
  NAND2_X1   g12210(.A1(new_n15046_), .A2(new_n12002_), .ZN(new_n15120_));
  AOI21_X1   g12211(.A1(new_n15062_), .A2(new_n12021_), .B(new_n11986_), .ZN(new_n15121_));
  AOI22_X1   g12212(.A1(new_n15120_), .A2(new_n15121_), .B1(new_n15118_), .B2(new_n15119_), .ZN(new_n15122_));
  OAI21_X1   g12213(.A1(new_n15122_), .A2(new_n14731_), .B(new_n14726_), .ZN(new_n15123_));
  OAI21_X1   g12214(.A1(new_n15089_), .A2(new_n15123_), .B(new_n15079_), .ZN(new_n15124_));
  AND2_X2    g12215(.A1(new_n15124_), .A2(pi0644), .Z(new_n15125_));
  NOR2_X1    g12216(.A1(new_n15067_), .A2(new_n12048_), .ZN(new_n15126_));
  AOI22_X1   g12217(.A1(new_n15126_), .A2(new_n15071_), .B1(new_n12048_), .B2(new_n15068_), .ZN(new_n15127_));
  AND2_X2    g12218(.A1(new_n15127_), .A2(new_n12082_), .Z(new_n15128_));
  OAI21_X1   g12219(.A1(new_n15125_), .A2(new_n15128_), .B(new_n12099_), .ZN(new_n15129_));
  NOR2_X1    g12220(.A1(new_n12092_), .A2(new_n15019_), .ZN(new_n15130_));
  AOI21_X1   g12221(.A1(new_n15049_), .A2(new_n12092_), .B(new_n15130_), .ZN(new_n15131_));
  OAI21_X1   g12222(.A1(new_n15131_), .A2(new_n15019_), .B(new_n12082_), .ZN(new_n15132_));
  AOI21_X1   g12223(.A1(new_n15019_), .A2(new_n15131_), .B(new_n15132_), .ZN(new_n15133_));
  XOR2_X1    g12224(.A1(new_n15133_), .A2(new_n15131_), .Z(new_n15134_));
  OAI21_X1   g12225(.A1(new_n15134_), .A2(new_n15129_), .B(new_n12081_), .ZN(new_n15135_));
  XOR2_X1    g12226(.A1(new_n15133_), .A2(new_n15020_), .Z(new_n15136_));
  NAND2_X1   g12227(.A1(new_n15136_), .A2(pi0715), .ZN(new_n15137_));
  OAI21_X1   g12228(.A1(new_n15127_), .A2(new_n12082_), .B(new_n13168_), .ZN(new_n15138_));
  NOR2_X1    g12229(.A1(new_n15125_), .A2(new_n15138_), .ZN(new_n15139_));
  AOI21_X1   g12230(.A1(new_n15137_), .A2(new_n15139_), .B(new_n11867_), .ZN(new_n15140_));
  NAND2_X1   g12231(.A1(new_n15124_), .A2(new_n14747_), .ZN(new_n15141_));
  AOI21_X1   g12232(.A1(new_n15140_), .A2(new_n15135_), .B(new_n15141_), .ZN(new_n15142_));
  NOR2_X1    g12233(.A1(new_n12965_), .A2(pi0145), .ZN(new_n15143_));
  MUX2_X1    g12234(.I0(new_n12894_), .I1(new_n12852_), .S(new_n3154_), .Z(new_n15144_));
  INV_X1     g12235(.I(pi0767), .ZN(new_n15145_));
  AOI21_X1   g12236(.A1(new_n12694_), .A2(pi0145), .B(new_n15145_), .ZN(new_n15146_));
  OAI21_X1   g12237(.A1(pi0145), .A2(new_n15144_), .B(new_n15146_), .ZN(new_n15147_));
  NOR2_X1    g12238(.A1(new_n12828_), .A2(pi0145), .ZN(new_n15148_));
  AOI21_X1   g12239(.A1(new_n15145_), .A2(new_n12829_), .B(new_n15148_), .ZN(new_n15149_));
  MUX2_X1    g12240(.I0(new_n15149_), .I1(new_n15147_), .S(new_n3172_), .Z(new_n15150_));
  NOR2_X1    g12241(.A1(new_n15150_), .A2(new_n3232_), .ZN(new_n15151_));
  AOI21_X1   g12242(.A1(new_n5323_), .A2(new_n3232_), .B(new_n15151_), .ZN(new_n15152_));
  INV_X1     g12243(.I(new_n15152_), .ZN(new_n15153_));
  INV_X1     g12244(.I(new_n15143_), .ZN(new_n15154_));
  OAI21_X1   g12245(.A1(new_n15154_), .A2(new_n11924_), .B(new_n11870_), .ZN(new_n15155_));
  AOI21_X1   g12246(.A1(new_n15153_), .A2(new_n11924_), .B(new_n15155_), .ZN(new_n15156_));
  NAND2_X1   g12247(.A1(new_n15152_), .A2(new_n11924_), .ZN(new_n15157_));
  OAI22_X1   g12248(.A1(new_n15157_), .A2(pi0609), .B1(new_n12996_), .B2(new_n15143_), .ZN(new_n15158_));
  NAND2_X1   g12249(.A1(new_n15158_), .A2(new_n11912_), .ZN(new_n15159_));
  OAI22_X1   g12250(.A1(new_n15157_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n15143_), .ZN(new_n15160_));
  NAND2_X1   g12251(.A1(new_n15160_), .A2(pi1155), .ZN(new_n15161_));
  NAND2_X1   g12252(.A1(new_n15159_), .A2(new_n15161_), .ZN(new_n15162_));
  NAND2_X1   g12253(.A1(new_n15162_), .A2(pi0785), .ZN(new_n15163_));
  XOR2_X1    g12254(.A1(new_n15163_), .A2(new_n15156_), .Z(new_n15164_));
  NAND2_X1   g12255(.A1(new_n15164_), .A2(new_n11969_), .ZN(new_n15165_));
  INV_X1     g12256(.I(new_n14635_), .ZN(new_n15166_));
  MUX2_X1    g12257(.I0(new_n15164_), .I1(new_n15143_), .S(new_n15166_), .Z(new_n15167_));
  NAND2_X1   g12258(.A1(new_n15167_), .A2(pi0781), .ZN(new_n15168_));
  NAND2_X1   g12259(.A1(new_n15168_), .A2(new_n15165_), .ZN(new_n15169_));
  NAND2_X1   g12260(.A1(new_n15169_), .A2(new_n11985_), .ZN(new_n15170_));
  INV_X1     g12261(.I(new_n15169_), .ZN(new_n15171_));
  MUX2_X1    g12262(.I0(new_n15154_), .I1(new_n15171_), .S(new_n14640_), .Z(new_n15172_));
  OAI21_X1   g12263(.A1(new_n15172_), .A2(new_n11985_), .B(new_n15170_), .ZN(new_n15173_));
  AND2_X2    g12264(.A1(new_n15173_), .A2(new_n11986_), .Z(new_n15174_));
  MUX2_X1    g12265(.I0(new_n15173_), .I1(new_n15143_), .S(new_n12003_), .Z(new_n15175_));
  AOI21_X1   g12266(.A1(new_n15175_), .A2(pi0788), .B(new_n15174_), .ZN(new_n15176_));
  NAND2_X1   g12267(.A1(new_n15176_), .A2(new_n12054_), .ZN(new_n15177_));
  OAI21_X1   g12268(.A1(new_n12054_), .A2(new_n15143_), .B(new_n15177_), .ZN(new_n15178_));
  NOR2_X1    g12269(.A1(new_n15143_), .A2(new_n12092_), .ZN(new_n15179_));
  AOI21_X1   g12270(.A1(new_n15178_), .A2(new_n12092_), .B(new_n15179_), .ZN(new_n15180_));
  NOR3_X1    g12271(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n15181_));
  NAND2_X1   g12272(.A1(new_n15180_), .A2(new_n15181_), .ZN(new_n15182_));
  INV_X1     g12273(.I(new_n15078_), .ZN(new_n15183_));
  NOR2_X1    g12274(.A1(new_n15154_), .A2(pi0647), .ZN(new_n15184_));
  OAI21_X1   g12275(.A1(new_n13395_), .A2(new_n5323_), .B(new_n3172_), .ZN(new_n15185_));
  NAND2_X1   g12276(.A1(new_n15185_), .A2(new_n3231_), .ZN(new_n15186_));
  NOR2_X1    g12277(.A1(new_n13399_), .A2(pi0145), .ZN(new_n15187_));
  INV_X1     g12278(.I(new_n15187_), .ZN(new_n15188_));
  INV_X1     g12279(.I(new_n13403_), .ZN(new_n15189_));
  OAI21_X1   g12280(.A1(new_n15189_), .A2(new_n15148_), .B(new_n15051_), .ZN(new_n15190_));
  AOI21_X1   g12281(.A1(new_n15188_), .A2(new_n15186_), .B(new_n15190_), .ZN(new_n15191_));
  NOR2_X1    g12282(.A1(new_n3232_), .A2(pi0698), .ZN(new_n15192_));
  AOI21_X1   g12283(.A1(new_n15154_), .A2(new_n15192_), .B(new_n15191_), .ZN(new_n15193_));
  NOR3_X1    g12284(.A1(new_n15154_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n15194_));
  NOR4_X1    g12285(.A1(new_n15193_), .A2(new_n12970_), .A3(pi1153), .A4(new_n15143_), .ZN(new_n15195_));
  NOR2_X1    g12286(.A1(new_n15195_), .A2(new_n15194_), .ZN(new_n15196_));
  MUX2_X1    g12287(.I0(new_n15196_), .I1(new_n15193_), .S(new_n11891_), .Z(new_n15197_));
  NOR2_X1    g12288(.A1(new_n15197_), .A2(new_n13024_), .ZN(new_n15198_));
  AOI21_X1   g12289(.A1(new_n13024_), .A2(new_n15143_), .B(new_n15198_), .ZN(new_n15199_));
  INV_X1     g12290(.I(new_n15199_), .ZN(new_n15200_));
  NOR2_X1    g12291(.A1(new_n15200_), .A2(new_n13714_), .ZN(new_n15201_));
  AOI21_X1   g12292(.A1(new_n13714_), .A2(new_n15154_), .B(new_n15201_), .ZN(new_n15202_));
  NAND2_X1   g12293(.A1(new_n15202_), .A2(new_n12032_), .ZN(new_n15203_));
  NAND2_X1   g12294(.A1(new_n15143_), .A2(new_n13713_), .ZN(new_n15204_));
  XNOR2_X1   g12295(.A1(new_n15203_), .A2(new_n15204_), .ZN(new_n15205_));
  NOR3_X1    g12296(.A1(new_n15154_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n15207_));
  INV_X1     g12297(.I(new_n15207_), .ZN(new_n15208_));
  NAND4_X1   g12298(.A1(new_n15205_), .A2(pi0628), .A3(new_n12026_), .A4(new_n15154_), .ZN(new_n15209_));
  NAND2_X1   g12299(.A1(new_n15209_), .A2(new_n15208_), .ZN(new_n15210_));
  MUX2_X1    g12300(.I0(new_n15210_), .I1(new_n15205_), .S(new_n11868_), .Z(new_n15211_));
  AOI21_X1   g12301(.A1(new_n15211_), .A2(pi0647), .B(new_n15184_), .ZN(new_n15212_));
  NAND2_X1   g12302(.A1(new_n15212_), .A2(new_n12060_), .ZN(new_n15213_));
  INV_X1     g12303(.I(new_n12090_), .ZN(new_n15214_));
  NOR2_X1    g12304(.A1(new_n15154_), .A2(new_n12061_), .ZN(new_n15215_));
  AOI21_X1   g12305(.A1(new_n15211_), .A2(new_n12061_), .B(new_n15215_), .ZN(new_n15216_));
  AOI21_X1   g12306(.A1(new_n15216_), .A2(pi0630), .B(new_n15214_), .ZN(new_n15217_));
  AOI21_X1   g12307(.A1(new_n15217_), .A2(new_n15213_), .B(new_n15183_), .ZN(new_n15218_));
  NAND2_X1   g12308(.A1(new_n15178_), .A2(new_n15218_), .ZN(new_n15219_));
  INV_X1     g12309(.I(new_n14729_), .ZN(new_n15220_));
  NAND2_X1   g12310(.A1(new_n14728_), .A2(new_n12026_), .ZN(new_n15221_));
  OAI21_X1   g12311(.A1(new_n12026_), .A2(new_n15220_), .B(new_n15221_), .ZN(new_n15222_));
  NOR2_X1    g12312(.A1(new_n15207_), .A2(new_n12030_), .ZN(new_n15223_));
  AND2_X2    g12313(.A1(new_n15209_), .A2(new_n12030_), .Z(new_n15224_));
  OAI21_X1   g12314(.A1(new_n15224_), .A2(new_n15223_), .B(new_n11868_), .ZN(new_n15225_));
  AOI21_X1   g12315(.A1(new_n15176_), .A2(new_n15222_), .B(new_n15225_), .ZN(new_n15226_));
  INV_X1     g12316(.I(new_n15202_), .ZN(new_n15227_));
  NOR3_X1    g12317(.A1(new_n15227_), .A2(new_n12013_), .A3(new_n15154_), .ZN(new_n15228_));
  AOI21_X1   g12318(.A1(new_n12014_), .A2(new_n15154_), .B(new_n15202_), .ZN(new_n15229_));
  OAI21_X1   g12319(.A1(new_n15228_), .A2(new_n15229_), .B(new_n12020_), .ZN(new_n15230_));
  NAND2_X1   g12320(.A1(new_n15175_), .A2(new_n12002_), .ZN(new_n15231_));
  AOI21_X1   g12321(.A1(new_n15231_), .A2(new_n15230_), .B(pi0788), .ZN(new_n15232_));
  NOR3_X1    g12322(.A1(new_n15150_), .A2(new_n15051_), .A3(new_n3231_), .ZN(new_n15242_));
  AOI21_X1   g12323(.A1(pi0145), .A2(new_n3232_), .B(new_n15242_), .ZN(new_n15243_));
  INV_X1     g12324(.I(new_n15195_), .ZN(new_n15244_));
  NAND2_X1   g12325(.A1(new_n15243_), .A2(pi0625), .ZN(new_n15245_));
  NAND2_X1   g12326(.A1(new_n15153_), .A2(pi0625), .ZN(new_n15246_));
  NAND4_X1   g12327(.A1(new_n15246_), .A2(new_n12977_), .A3(new_n15244_), .A4(new_n15245_), .ZN(new_n15247_));
  NAND2_X1   g12328(.A1(new_n15152_), .A2(new_n12970_), .ZN(new_n15248_));
  AND3_X2    g12329(.A1(new_n15245_), .A2(new_n11893_), .A3(new_n15248_), .Z(new_n15249_));
  OAI21_X1   g12330(.A1(new_n15249_), .A2(new_n15194_), .B(new_n13657_), .ZN(new_n15250_));
  AOI21_X1   g12331(.A1(new_n15250_), .A2(new_n15247_), .B(new_n11891_), .ZN(new_n15251_));
  AOI21_X1   g12332(.A1(new_n11891_), .A2(new_n15243_), .B(new_n15251_), .ZN(new_n15252_));
  INV_X1     g12333(.I(new_n15197_), .ZN(new_n15253_));
  NOR4_X1    g12334(.A1(new_n15252_), .A2(new_n11903_), .A3(pi1155), .A4(new_n15253_), .ZN(new_n15254_));
  NAND2_X1   g12335(.A1(new_n15159_), .A2(pi0660), .ZN(new_n15255_));
  NOR3_X1    g12336(.A1(new_n15197_), .A2(new_n11903_), .A3(new_n11912_), .ZN(new_n15256_));
  NAND2_X1   g12337(.A1(new_n15161_), .A2(new_n11923_), .ZN(new_n15257_));
  OAI22_X1   g12338(.A1(new_n15254_), .A2(new_n15255_), .B1(new_n15256_), .B2(new_n15257_), .ZN(new_n15258_));
  MUX2_X1    g12339(.I0(new_n15258_), .I1(new_n15252_), .S(new_n11870_), .Z(new_n15259_));
  INV_X1     g12340(.I(new_n15259_), .ZN(new_n15260_));
  AOI21_X1   g12341(.A1(new_n15200_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n15261_));
  INV_X1     g12342(.I(new_n15164_), .ZN(new_n15262_));
  NAND3_X1   g12343(.A1(new_n11934_), .A2(new_n11949_), .A3(pi1154), .ZN(new_n15263_));
  OAI21_X1   g12344(.A1(new_n15262_), .A2(new_n15263_), .B(pi0618), .ZN(new_n15264_));
  NOR2_X1    g12345(.A1(new_n15264_), .A2(new_n15261_), .ZN(new_n15265_));
  NAND2_X1   g12346(.A1(new_n15259_), .A2(new_n11934_), .ZN(new_n15266_));
  NOR2_X1    g12347(.A1(new_n15199_), .A2(new_n11934_), .ZN(new_n15267_));
  NAND2_X1   g12348(.A1(new_n11950_), .A2(pi0618), .ZN(new_n15268_));
  NOR2_X1    g12349(.A1(new_n15262_), .A2(new_n15268_), .ZN(new_n15269_));
  NOR4_X1    g12350(.A1(new_n15269_), .A2(pi0627), .A3(pi1154), .A4(new_n15267_), .ZN(new_n15270_));
  AOI22_X1   g12351(.A1(new_n15266_), .A2(new_n15270_), .B1(new_n15259_), .B2(new_n15265_), .ZN(new_n15271_));
  MUX2_X1    g12352(.I0(new_n15271_), .I1(new_n15260_), .S(new_n11969_), .Z(new_n15272_));
  NAND3_X1   g12353(.A1(new_n11967_), .A2(new_n11966_), .A3(pi1159), .ZN(new_n15273_));
  NOR2_X1    g12354(.A1(new_n15171_), .A2(new_n15273_), .ZN(new_n15274_));
  NAND2_X1   g12355(.A1(new_n11869_), .A2(pi0619), .ZN(new_n15275_));
  OR3_X2     g12356(.A1(new_n15272_), .A2(new_n15274_), .A3(new_n15275_), .Z(new_n15276_));
  NOR2_X1    g12357(.A1(new_n11967_), .A2(pi1159), .ZN(new_n15277_));
  NOR2_X1    g12358(.A1(pi0648), .A2(pi1159), .ZN(new_n15278_));
  OAI21_X1   g12359(.A1(new_n15227_), .A2(new_n11967_), .B(new_n15278_), .ZN(new_n15279_));
  AOI21_X1   g12360(.A1(new_n15169_), .A2(new_n15277_), .B(new_n15279_), .ZN(new_n15280_));
  OAI21_X1   g12361(.A1(new_n15272_), .A2(pi0619), .B(new_n15280_), .ZN(new_n15281_));
  OAI21_X1   g12362(.A1(new_n15272_), .A2(new_n11999_), .B(new_n11985_), .ZN(new_n15282_));
  AOI21_X1   g12363(.A1(new_n15276_), .A2(new_n15281_), .B(new_n15282_), .ZN(new_n15283_));
  NOR4_X1    g12364(.A1(new_n15226_), .A2(new_n15232_), .A3(new_n14731_), .A4(new_n15283_), .ZN(new_n15284_));
  OAI21_X1   g12365(.A1(new_n15284_), .A2(new_n14725_), .B(new_n15219_), .ZN(new_n15285_));
  NOR4_X1    g12366(.A1(new_n15285_), .A2(new_n15182_), .A3(new_n12082_), .A4(pi0790), .ZN(new_n15286_));
  NAND2_X1   g12367(.A1(new_n15212_), .A2(pi1157), .ZN(new_n15287_));
  NAND2_X1   g12368(.A1(new_n15216_), .A2(new_n12049_), .ZN(new_n15288_));
  NAND2_X1   g12369(.A1(new_n15287_), .A2(new_n15288_), .ZN(new_n15289_));
  NOR2_X1    g12370(.A1(new_n15211_), .A2(pi0787), .ZN(new_n15290_));
  AOI21_X1   g12371(.A1(new_n15289_), .A2(pi0787), .B(new_n15290_), .ZN(new_n15291_));
  AOI21_X1   g12372(.A1(new_n15291_), .A2(new_n12082_), .B(new_n12099_), .ZN(new_n15292_));
  NAND2_X1   g12373(.A1(new_n15182_), .A2(new_n15292_), .ZN(new_n15293_));
  INV_X1     g12374(.I(new_n15291_), .ZN(new_n15294_));
  NAND3_X1   g12375(.A1(new_n15285_), .A2(new_n12082_), .A3(new_n15294_), .ZN(new_n15295_));
  OAI21_X1   g12376(.A1(new_n15285_), .A2(pi0644), .B(new_n15291_), .ZN(new_n15296_));
  NOR2_X1    g12377(.A1(new_n12081_), .A2(pi0715), .ZN(new_n15299_));
  NAND3_X1   g12378(.A1(new_n15296_), .A2(new_n15295_), .A3(new_n15299_), .ZN(new_n15300_));
  AOI21_X1   g12379(.A1(new_n15300_), .A2(new_n15293_), .B(new_n11867_), .ZN(new_n15301_));
  OAI21_X1   g12380(.A1(new_n15301_), .A2(new_n15286_), .B(new_n6845_), .ZN(new_n15302_));
  AOI21_X1   g12381(.A1(po1038), .A2(new_n5323_), .B(pi0832), .ZN(new_n15303_));
  AOI21_X1   g12382(.A1(new_n15302_), .A2(new_n15303_), .B(new_n15142_), .ZN(po0302));
  INV_X1     g12383(.I(pi0907), .ZN(new_n15305_));
  NOR2_X1    g12384(.A1(new_n13638_), .A2(new_n15305_), .ZN(new_n15306_));
  MUX2_X1    g12385(.I0(new_n15306_), .I1(pi0743), .S(pi0947), .Z(new_n15307_));
  INV_X1     g12386(.I(new_n15307_), .ZN(new_n15308_));
  NOR2_X1    g12387(.A1(new_n15308_), .A2(new_n2926_), .ZN(new_n15309_));
  NAND4_X1   g12388(.A1(new_n15309_), .A2(new_n3560_), .A3(pi0832), .A4(new_n2926_), .ZN(new_n15310_));
  NAND2_X1   g12389(.A1(new_n12886_), .A2(new_n15308_), .ZN(new_n15311_));
  AOI21_X1   g12390(.A1(new_n15311_), .A2(pi0215), .B(pi0146), .ZN(new_n15312_));
  OAI21_X1   g12391(.A1(new_n12709_), .A2(new_n12745_), .B(new_n15312_), .ZN(new_n15313_));
  NOR2_X1    g12392(.A1(new_n5091_), .A2(pi0907), .ZN(new_n15314_));
  INV_X1     g12393(.I(new_n15314_), .ZN(new_n15315_));
  NAND2_X1   g12394(.A1(new_n15315_), .A2(pi0146), .ZN(new_n15316_));
  OAI21_X1   g12395(.A1(new_n12767_), .A2(pi0743), .B(new_n5473_), .ZN(new_n15317_));
  AOI21_X1   g12396(.A1(new_n3560_), .A2(new_n12767_), .B(new_n15317_), .ZN(new_n15318_));
  NOR2_X1    g12397(.A1(new_n15315_), .A2(new_n3560_), .ZN(new_n15319_));
  NAND2_X1   g12398(.A1(new_n12776_), .A2(new_n15306_), .ZN(new_n15320_));
  AOI22_X1   g12399(.A1(new_n12879_), .A2(new_n15319_), .B1(new_n5473_), .B2(new_n15320_), .ZN(new_n15321_));
  OAI22_X1   g12400(.A1(new_n15321_), .A2(new_n15318_), .B1(new_n12776_), .B2(new_n15316_), .ZN(new_n15322_));
  NOR2_X1    g12401(.A1(new_n12132_), .A2(pi0146), .ZN(new_n15323_));
  AOI21_X1   g12402(.A1(new_n15307_), .A2(new_n12132_), .B(new_n15323_), .ZN(new_n15324_));
  MUX2_X1    g12403(.I0(new_n15322_), .I1(new_n15324_), .S(new_n3284_), .Z(new_n15325_));
  OAI21_X1   g12404(.A1(new_n15325_), .A2(pi0215), .B(new_n15313_), .ZN(new_n15326_));
  AOI21_X1   g12405(.A1(new_n12784_), .A2(new_n3560_), .B(new_n5141_), .ZN(new_n15327_));
  NOR4_X1    g12406(.A1(new_n15327_), .A2(new_n2604_), .A3(new_n12784_), .A4(new_n15308_), .ZN(new_n15328_));
  NOR2_X1    g12407(.A1(new_n15328_), .A2(pi0299), .ZN(new_n15329_));
  NAND4_X1   g12408(.A1(new_n12759_), .A2(new_n3560_), .A3(new_n6460_), .A4(new_n15307_), .ZN(new_n15330_));
  NAND3_X1   g12409(.A1(new_n12767_), .A2(pi0146), .A3(new_n15307_), .ZN(new_n15331_));
  OAI21_X1   g12410(.A1(new_n12776_), .A2(pi0146), .B(new_n15308_), .ZN(new_n15332_));
  NAND4_X1   g12411(.A1(new_n15330_), .A2(new_n6460_), .A3(new_n15331_), .A4(new_n15332_), .ZN(new_n15333_));
  OAI21_X1   g12412(.A1(new_n15324_), .A2(new_n3155_), .B(new_n2604_), .ZN(new_n15334_));
  AOI21_X1   g12413(.A1(new_n15333_), .A2(new_n3155_), .B(new_n15334_), .ZN(new_n15335_));
  AOI21_X1   g12414(.A1(new_n12646_), .A2(new_n3560_), .B(pi0299), .ZN(new_n15336_));
  NAND2_X1   g12415(.A1(new_n12584_), .A2(new_n15307_), .ZN(new_n15337_));
  OAI21_X1   g12416(.A1(new_n15336_), .A2(new_n15337_), .B(new_n3154_), .ZN(new_n15338_));
  NOR2_X1    g12417(.A1(new_n12828_), .A2(pi0146), .ZN(new_n15339_));
  NAND4_X1   g12418(.A1(new_n5156_), .A2(new_n3172_), .A3(new_n7833_), .A4(new_n15309_), .ZN(new_n15340_));
  OAI21_X1   g12419(.A1(new_n15339_), .A2(new_n15340_), .B(pi0039), .ZN(new_n15341_));
  AOI21_X1   g12420(.A1(new_n15338_), .A2(new_n3172_), .B(new_n15341_), .ZN(new_n15342_));
  OAI21_X1   g12421(.A1(new_n15335_), .A2(new_n15329_), .B(new_n15342_), .ZN(new_n15343_));
  AOI21_X1   g12422(.A1(new_n15326_), .A2(pi0299), .B(new_n15343_), .ZN(new_n15344_));
  OAI21_X1   g12423(.A1(new_n7832_), .A2(pi0146), .B(new_n13184_), .ZN(new_n15345_));
  OAI21_X1   g12424(.A1(new_n15344_), .A2(new_n15345_), .B(new_n15310_), .ZN(po0303));
  NAND2_X1   g12425(.A1(pi0726), .A2(pi0907), .ZN(new_n15347_));
  MUX2_X1    g12426(.I0(new_n15347_), .I1(pi0770), .S(pi0947), .Z(new_n15348_));
  MUX2_X1    g12427(.I0(new_n8836_), .I1(new_n15348_), .S(new_n2925_), .Z(new_n15349_));
  NOR2_X1    g12428(.A1(new_n15349_), .A2(new_n13184_), .ZN(new_n15350_));
  NOR2_X1    g12429(.A1(new_n15305_), .A2(pi0947), .ZN(new_n15351_));
  NOR3_X1    g12430(.A1(new_n12697_), .A2(pi0039), .A3(new_n15351_), .ZN(new_n15352_));
  NOR2_X1    g12431(.A1(new_n15351_), .A2(pi0299), .ZN(new_n15353_));
  NAND2_X1   g12432(.A1(new_n12792_), .A2(new_n15353_), .ZN(new_n15354_));
  INV_X1     g12433(.I(new_n12768_), .ZN(new_n15355_));
  AOI21_X1   g12434(.A1(new_n12879_), .A2(new_n5090_), .B(new_n15355_), .ZN(new_n15356_));
  NOR2_X1    g12435(.A1(new_n12767_), .A2(new_n5473_), .ZN(new_n15357_));
  NOR2_X1    g12436(.A1(new_n15356_), .A2(new_n15357_), .ZN(new_n15358_));
  NOR2_X1    g12437(.A1(new_n15358_), .A2(new_n3284_), .ZN(new_n15359_));
  INV_X1     g12438(.I(new_n15359_), .ZN(new_n15360_));
  NOR2_X1    g12439(.A1(new_n12881_), .A2(new_n15351_), .ZN(new_n15361_));
  INV_X1     g12440(.I(new_n15361_), .ZN(new_n15362_));
  AOI21_X1   g12441(.A1(new_n15360_), .A2(new_n15362_), .B(pi0215), .ZN(new_n15363_));
  AOI21_X1   g12442(.A1(pi0215), .A2(new_n12745_), .B(new_n15363_), .ZN(new_n15364_));
  INV_X1     g12443(.I(new_n15364_), .ZN(new_n15365_));
  NOR3_X1    g12444(.A1(new_n12784_), .A2(new_n2566_), .A3(new_n5473_), .ZN(new_n15366_));
  NOR2_X1    g12445(.A1(new_n15365_), .A2(new_n15366_), .ZN(new_n15367_));
  NOR2_X1    g12446(.A1(new_n15367_), .A2(new_n2587_), .ZN(new_n15368_));
  XOR2_X1    g12447(.A1(new_n15368_), .A2(new_n15354_), .Z(new_n15369_));
  NAND2_X1   g12448(.A1(new_n15369_), .A2(pi0039), .ZN(new_n15370_));
  XOR2_X1    g12449(.A1(new_n15370_), .A2(new_n15352_), .Z(new_n15371_));
  INV_X1     g12450(.I(new_n15351_), .ZN(new_n15372_));
  NOR2_X1    g12451(.A1(new_n12697_), .A2(new_n15372_), .ZN(new_n15373_));
  INV_X1     g12452(.I(new_n15373_), .ZN(new_n15374_));
  NOR2_X1    g12453(.A1(new_n15374_), .A2(pi0039), .ZN(new_n15375_));
  INV_X1     g12454(.I(new_n12792_), .ZN(new_n15376_));
  NOR2_X1    g12455(.A1(new_n15376_), .A2(new_n15372_), .ZN(new_n15377_));
  NOR2_X1    g12456(.A1(new_n15377_), .A2(pi0299), .ZN(new_n15378_));
  NOR2_X1    g12457(.A1(new_n15378_), .A2(pi0299), .ZN(new_n15379_));
  AOI21_X1   g12458(.A1(new_n15379_), .A2(pi0039), .B(new_n15375_), .ZN(new_n15380_));
  NOR2_X1    g12459(.A1(new_n13368_), .A2(new_n15372_), .ZN(new_n15381_));
  OAI21_X1   g12460(.A1(new_n15380_), .A2(new_n8836_), .B(new_n3172_), .ZN(new_n15383_));
  AOI21_X1   g12461(.A1(new_n15371_), .A2(pi0147), .B(new_n15383_), .ZN(new_n15384_));
  NOR3_X1    g12462(.A1(new_n12697_), .A2(pi0039), .A3(new_n5093_), .ZN(new_n15385_));
  OAI21_X1   g12463(.A1(new_n2491_), .A2(new_n12505_), .B(new_n12790_), .ZN(new_n15386_));
  AOI21_X1   g12464(.A1(new_n15386_), .A2(new_n5092_), .B(pi0223), .ZN(new_n15387_));
  INV_X1     g12465(.I(new_n15387_), .ZN(new_n15388_));
  NOR2_X1    g12466(.A1(new_n12785_), .A2(new_n12787_), .ZN(new_n15389_));
  NOR2_X1    g12467(.A1(new_n15389_), .A2(pi0947), .ZN(new_n15390_));
  NOR2_X1    g12468(.A1(new_n15390_), .A2(new_n2604_), .ZN(new_n15391_));
  INV_X1     g12469(.I(new_n15389_), .ZN(new_n15392_));
  AOI21_X1   g12470(.A1(new_n15392_), .A2(new_n15372_), .B(new_n2604_), .ZN(new_n15393_));
  NOR2_X1    g12471(.A1(new_n15391_), .A2(new_n15393_), .ZN(new_n15394_));
  AOI21_X1   g12472(.A1(new_n15388_), .A2(new_n15394_), .B(pi0299), .ZN(new_n15395_));
  INV_X1     g12473(.I(new_n15395_), .ZN(new_n15396_));
  NOR2_X1    g12474(.A1(pi0299), .A2(pi0947), .ZN(new_n15397_));
  NAND2_X1   g12475(.A1(new_n15365_), .A2(new_n15397_), .ZN(new_n15398_));
  NAND2_X1   g12476(.A1(new_n15398_), .A2(new_n15396_), .ZN(new_n15399_));
  INV_X1     g12477(.I(new_n15399_), .ZN(new_n15400_));
  NOR3_X1    g12478(.A1(new_n15400_), .A2(new_n3154_), .A3(new_n15385_), .ZN(new_n15401_));
  NOR3_X1    g12479(.A1(new_n12697_), .A2(pi0039), .A3(new_n5093_), .ZN(new_n15402_));
  NOR2_X1    g12480(.A1(new_n15401_), .A2(new_n15402_), .ZN(new_n15403_));
  INV_X1     g12481(.I(new_n15403_), .ZN(new_n15404_));
  NOR2_X1    g12482(.A1(new_n15404_), .A2(new_n8836_), .ZN(new_n15405_));
  NOR2_X1    g12483(.A1(new_n12697_), .A2(new_n5092_), .ZN(new_n15406_));
  INV_X1     g12484(.I(new_n15406_), .ZN(new_n15407_));
  NOR2_X1    g12485(.A1(new_n15407_), .A2(pi0039), .ZN(new_n15408_));
  NOR2_X1    g12486(.A1(new_n15376_), .A2(new_n5092_), .ZN(new_n15409_));
  NOR2_X1    g12487(.A1(new_n12709_), .A2(new_n2566_), .ZN(new_n15410_));
  NOR2_X1    g12488(.A1(new_n12133_), .A2(new_n5092_), .ZN(new_n15411_));
  NAND2_X1   g12489(.A1(new_n15411_), .A2(new_n3284_), .ZN(new_n15412_));
  NAND3_X1   g12490(.A1(new_n12882_), .A2(new_n2566_), .A3(new_n15412_), .ZN(new_n15413_));
  OAI21_X1   g12491(.A1(new_n15410_), .A2(new_n15413_), .B(pi0299), .ZN(new_n15414_));
  NOR3_X1    g12492(.A1(new_n15409_), .A2(pi0299), .A3(new_n15414_), .ZN(new_n15415_));
  NOR2_X1    g12493(.A1(new_n15409_), .A2(pi0299), .ZN(new_n15416_));
  INV_X1     g12494(.I(new_n15414_), .ZN(new_n15417_));
  NOR2_X1    g12495(.A1(new_n15416_), .A2(new_n15417_), .ZN(new_n15418_));
  NOR2_X1    g12496(.A1(new_n15418_), .A2(new_n15415_), .ZN(new_n15419_));
  AOI21_X1   g12497(.A1(new_n15419_), .A2(pi0039), .B(new_n15408_), .ZN(new_n15420_));
  NOR2_X1    g12498(.A1(new_n12899_), .A2(new_n5093_), .ZN(new_n15421_));
  NOR2_X1    g12499(.A1(pi0038), .A2(pi0770), .ZN(new_n15423_));
  OAI21_X1   g12500(.A1(new_n15420_), .A2(new_n8836_), .B(new_n15423_), .ZN(new_n15424_));
  NOR2_X1    g12501(.A1(pi0726), .A2(pi0770), .ZN(new_n15425_));
  OAI21_X1   g12502(.A1(new_n15405_), .A2(new_n15424_), .B(new_n15425_), .ZN(new_n15426_));
  INV_X1     g12503(.I(pi0770), .ZN(new_n15427_));
  NOR3_X1    g12504(.A1(new_n12899_), .A2(new_n3172_), .A3(pi0947), .ZN(new_n15428_));
  AOI21_X1   g12505(.A1(new_n12852_), .A2(new_n5473_), .B(pi0039), .ZN(new_n15429_));
  NAND2_X1   g12506(.A1(new_n12792_), .A2(new_n15397_), .ZN(new_n15430_));
  NOR2_X1    g12507(.A1(new_n12784_), .A2(new_n15372_), .ZN(new_n15431_));
  NOR2_X1    g12508(.A1(new_n12745_), .A2(new_n2566_), .ZN(new_n15432_));
  INV_X1     g12509(.I(new_n15432_), .ZN(new_n15433_));
  NOR2_X1    g12510(.A1(new_n15433_), .A2(new_n15431_), .ZN(new_n15434_));
  NOR2_X1    g12511(.A1(new_n12767_), .A2(new_n15372_), .ZN(new_n15435_));
  NOR2_X1    g12512(.A1(new_n15356_), .A2(new_n15435_), .ZN(new_n15436_));
  NOR2_X1    g12513(.A1(new_n15436_), .A2(new_n3284_), .ZN(new_n15437_));
  NOR2_X1    g12514(.A1(new_n15437_), .A2(pi0215), .ZN(new_n15438_));
  NOR3_X1    g12515(.A1(new_n15438_), .A2(pi0947), .A3(new_n12881_), .ZN(new_n15439_));
  NOR2_X1    g12516(.A1(new_n15439_), .A2(new_n15434_), .ZN(new_n15440_));
  NOR2_X1    g12517(.A1(new_n15440_), .A2(new_n2587_), .ZN(new_n15441_));
  XOR2_X1    g12518(.A1(new_n15441_), .A2(new_n15430_), .Z(new_n15442_));
  AOI21_X1   g12519(.A1(new_n15442_), .A2(pi0039), .B(new_n15429_), .ZN(new_n15443_));
  AOI21_X1   g12520(.A1(new_n15443_), .A2(new_n3172_), .B(new_n15428_), .ZN(new_n15444_));
  INV_X1     g12521(.I(new_n15444_), .ZN(new_n15445_));
  AOI21_X1   g12522(.A1(new_n15445_), .A2(new_n15427_), .B(pi0147), .ZN(new_n15446_));
  AOI21_X1   g12523(.A1(new_n12898_), .A2(pi0947), .B(new_n3172_), .ZN(new_n15447_));
  AOI21_X1   g12524(.A1(new_n12852_), .A2(pi0947), .B(pi0039), .ZN(new_n15448_));
  INV_X1     g12525(.I(new_n15448_), .ZN(new_n15449_));
  NOR2_X1    g12526(.A1(new_n15376_), .A2(new_n5473_), .ZN(new_n15450_));
  NOR2_X1    g12527(.A1(new_n15450_), .A2(pi0299), .ZN(new_n15451_));
  NOR2_X1    g12528(.A1(new_n12133_), .A2(new_n5473_), .ZN(new_n15452_));
  NOR2_X1    g12529(.A1(new_n15452_), .A2(new_n3285_), .ZN(new_n15453_));
  NOR2_X1    g12530(.A1(new_n15453_), .A2(pi0215), .ZN(new_n15454_));
  OAI21_X1   g12531(.A1(new_n15357_), .A2(new_n3284_), .B(new_n15454_), .ZN(new_n15455_));
  INV_X1     g12532(.I(new_n15455_), .ZN(new_n15456_));
  NOR3_X1    g12533(.A1(new_n15456_), .A2(new_n15366_), .A3(new_n2587_), .ZN(new_n15457_));
  NOR2_X1    g12534(.A1(new_n15451_), .A2(new_n15457_), .ZN(new_n15458_));
  OAI21_X1   g12535(.A1(new_n15458_), .A2(new_n3154_), .B(new_n15449_), .ZN(new_n15459_));
  AOI21_X1   g12536(.A1(new_n15459_), .A2(new_n3172_), .B(new_n15447_), .ZN(new_n15460_));
  INV_X1     g12537(.I(new_n15460_), .ZN(new_n15461_));
  NOR3_X1    g12538(.A1(new_n15461_), .A2(new_n8836_), .A3(pi0770), .ZN(new_n15462_));
  INV_X1     g12539(.I(pi0726), .ZN(new_n15463_));
  NAND4_X1   g12540(.A1(new_n12902_), .A2(new_n15463_), .A3(pi0770), .A4(new_n7833_), .ZN(new_n15464_));
  NOR3_X1    g12541(.A1(new_n15446_), .A2(new_n15462_), .A3(new_n15464_), .ZN(new_n15465_));
  OAI21_X1   g12542(.A1(new_n15384_), .A2(new_n15426_), .B(new_n15465_), .ZN(new_n15466_));
  AOI21_X1   g12543(.A1(new_n7833_), .A2(new_n8836_), .B(pi0832), .ZN(new_n15467_));
  AOI21_X1   g12544(.A1(new_n15466_), .A2(new_n15467_), .B(new_n15350_), .ZN(po0304));
  NOR2_X1    g12545(.A1(new_n13190_), .A2(new_n5473_), .ZN(new_n15469_));
  NOR4_X1    g12546(.A1(new_n15372_), .A2(new_n13199_), .A3(new_n2925_), .A4(new_n15469_), .ZN(new_n15470_));
  NAND3_X1   g12547(.A1(new_n2925_), .A2(new_n4130_), .A3(new_n13184_), .ZN(new_n15471_));
  NAND4_X1   g12548(.A1(new_n15400_), .A2(pi0148), .A3(new_n13190_), .A4(new_n15419_), .ZN(new_n15472_));
  INV_X1     g12549(.I(new_n15369_), .ZN(new_n15473_));
  NOR2_X1    g12550(.A1(new_n15473_), .A2(new_n11804_), .ZN(new_n15474_));
  NOR2_X1    g12551(.A1(new_n15376_), .A2(pi0299), .ZN(new_n15475_));
  OAI21_X1   g12552(.A1(new_n15475_), .A2(new_n4130_), .B(new_n13190_), .ZN(new_n15476_));
  OAI21_X1   g12553(.A1(new_n15474_), .A2(new_n15476_), .B(new_n15472_), .ZN(new_n15477_));
  AOI21_X1   g12554(.A1(new_n12697_), .A2(new_n4130_), .B(pi0039), .ZN(new_n15478_));
  INV_X1     g12555(.I(new_n15478_), .ZN(new_n15479_));
  AOI21_X1   g12556(.A1(new_n13190_), .A2(pi0947), .B(new_n15407_), .ZN(new_n15480_));
  AOI21_X1   g12557(.A1(new_n15480_), .A2(new_n15479_), .B(new_n2545_), .ZN(new_n15481_));
  AOI21_X1   g12558(.A1(new_n13190_), .A2(pi0947), .B(new_n5092_), .ZN(new_n15482_));
  NOR3_X1    g12559(.A1(new_n13368_), .A2(pi0148), .A3(new_n15482_), .ZN(new_n15483_));
  AOI21_X1   g12560(.A1(new_n12828_), .A2(new_n15482_), .B(new_n4130_), .ZN(new_n15484_));
  OAI21_X1   g12561(.A1(new_n15483_), .A2(new_n15484_), .B(new_n13404_), .ZN(new_n15485_));
  AOI21_X1   g12562(.A1(new_n15477_), .A2(new_n15481_), .B(new_n15485_), .ZN(new_n15486_));
  INV_X1     g12563(.I(new_n15440_), .ZN(new_n15487_));
  NOR2_X1    g12564(.A1(new_n15456_), .A2(new_n15366_), .ZN(new_n15488_));
  INV_X1     g12565(.I(new_n15488_), .ZN(new_n15489_));
  AOI21_X1   g12566(.A1(new_n15487_), .A2(new_n15489_), .B(new_n4130_), .ZN(new_n15490_));
  NAND2_X1   g12567(.A1(new_n15490_), .A2(pi0299), .ZN(new_n15491_));
  NAND2_X1   g12568(.A1(new_n4130_), .A2(new_n13190_), .ZN(new_n15492_));
  OAI21_X1   g12569(.A1(new_n12894_), .A2(new_n15492_), .B(pi0039), .ZN(new_n15493_));
  INV_X1     g12570(.I(new_n15451_), .ZN(new_n15494_));
  NOR2_X1    g12571(.A1(new_n12792_), .A2(pi0148), .ZN(new_n15495_));
  NOR4_X1    g12572(.A1(new_n15478_), .A2(new_n13190_), .A3(new_n5473_), .A4(new_n12697_), .ZN(new_n15496_));
  OAI21_X1   g12573(.A1(new_n13368_), .A2(new_n15469_), .B(pi0038), .ZN(new_n15497_));
  NAND3_X1   g12574(.A1(new_n12899_), .A2(pi0148), .A3(new_n15497_), .ZN(new_n15498_));
  NOR2_X1    g12575(.A1(new_n3232_), .A2(new_n5223_), .ZN(new_n15499_));
  INV_X1     g12576(.I(new_n15499_), .ZN(new_n15500_));
  NAND4_X1   g12577(.A1(new_n15498_), .A2(new_n13190_), .A3(new_n13404_), .A4(new_n15500_), .ZN(new_n15501_));
  NOR4_X1    g12578(.A1(new_n15494_), .A2(new_n15495_), .A3(new_n15496_), .A4(new_n15501_), .ZN(new_n15502_));
  NAND3_X1   g12579(.A1(new_n15491_), .A2(new_n15493_), .A3(new_n15502_), .ZN(new_n15503_));
  NOR2_X1    g12580(.A1(new_n5055_), .A2(new_n4130_), .ZN(new_n15504_));
  OAI21_X1   g12581(.A1(new_n15504_), .A2(pi0832), .B(new_n5055_), .ZN(new_n15505_));
  AOI21_X1   g12582(.A1(new_n15500_), .A2(new_n4130_), .B(new_n15505_), .ZN(new_n15506_));
  OAI21_X1   g12583(.A1(new_n15486_), .A2(new_n15503_), .B(new_n15506_), .ZN(new_n15507_));
  OAI21_X1   g12584(.A1(new_n15470_), .A2(new_n15471_), .B(new_n15507_), .ZN(po0305));
  INV_X1     g12585(.I(pi0755), .ZN(new_n15509_));
  NOR2_X1    g12586(.A1(new_n12792_), .A2(new_n15353_), .ZN(new_n15510_));
  NAND3_X1   g12587(.A1(new_n12792_), .A2(new_n7067_), .A3(new_n2587_), .ZN(new_n15511_));
  OAI21_X1   g12588(.A1(pi0149), .A2(new_n15475_), .B(new_n15368_), .ZN(new_n15512_));
  AOI22_X1   g12589(.A1(new_n15512_), .A2(new_n15511_), .B1(new_n15509_), .B2(new_n15510_), .ZN(new_n15513_));
  NAND2_X1   g12590(.A1(new_n15400_), .A2(pi0149), .ZN(new_n15514_));
  INV_X1     g12591(.I(new_n15419_), .ZN(new_n15515_));
  NAND2_X1   g12592(.A1(new_n15515_), .A2(pi0149), .ZN(new_n15516_));
  NAND4_X1   g12593(.A1(new_n15514_), .A2(pi0039), .A3(new_n15509_), .A4(new_n15516_), .ZN(new_n15517_));
  OAI21_X1   g12594(.A1(new_n12852_), .A2(pi0149), .B(new_n3154_), .ZN(new_n15518_));
  NOR2_X1    g12595(.A1(new_n5473_), .A2(pi0755), .ZN(new_n15519_));
  NAND3_X1   g12596(.A1(new_n15518_), .A2(new_n12852_), .A3(new_n15519_), .ZN(new_n15520_));
  OAI22_X1   g12597(.A1(new_n15517_), .A2(new_n15513_), .B1(new_n15373_), .B2(new_n15520_), .ZN(new_n15521_));
  NAND2_X1   g12598(.A1(new_n13368_), .A2(new_n7067_), .ZN(new_n15522_));
  NOR2_X1    g12599(.A1(new_n12110_), .A2(new_n5092_), .ZN(new_n15523_));
  NOR4_X1    g12600(.A1(new_n15523_), .A2(pi0039), .A3(new_n15509_), .A4(new_n5473_), .ZN(new_n15524_));
  NOR2_X1    g12601(.A1(new_n15524_), .A2(new_n3172_), .ZN(new_n15525_));
  AOI22_X1   g12602(.A1(new_n15521_), .A2(new_n3172_), .B1(new_n15522_), .B2(new_n15525_), .ZN(new_n15526_));
  AOI21_X1   g12603(.A1(pi0149), .A2(new_n2587_), .B(new_n15457_), .ZN(new_n15527_));
  AOI21_X1   g12604(.A1(new_n15440_), .A2(new_n7067_), .B(new_n15527_), .ZN(new_n15528_));
  AOI21_X1   g12605(.A1(new_n7067_), .A2(new_n15376_), .B(new_n15494_), .ZN(new_n15529_));
  NOR3_X1    g12606(.A1(new_n15528_), .A2(pi0755), .A3(new_n15529_), .ZN(new_n15530_));
  NOR2_X1    g12607(.A1(pi0039), .A2(pi0755), .ZN(new_n15531_));
  OAI21_X1   g12608(.A1(new_n12894_), .A2(pi0149), .B(new_n15531_), .ZN(new_n15532_));
  AND2_X2    g12609(.A1(new_n15520_), .A2(new_n3172_), .Z(new_n15533_));
  OAI21_X1   g12610(.A1(new_n15530_), .A2(new_n15532_), .B(new_n15533_), .ZN(new_n15534_));
  INV_X1     g12611(.I(pi0725), .ZN(new_n15535_));
  NAND2_X1   g12612(.A1(new_n12899_), .A2(pi0149), .ZN(new_n15536_));
  NOR2_X1    g12613(.A1(new_n13368_), .A2(new_n15519_), .ZN(new_n15537_));
  NOR2_X1    g12614(.A1(new_n15537_), .A2(new_n3172_), .ZN(new_n15538_));
  AOI21_X1   g12615(.A1(new_n15536_), .A2(new_n15538_), .B(new_n15535_), .ZN(new_n15539_));
  AOI21_X1   g12616(.A1(new_n15534_), .A2(new_n15539_), .B(new_n7833_), .ZN(new_n15540_));
  OAI21_X1   g12617(.A1(new_n15526_), .A2(pi0725), .B(new_n15540_), .ZN(new_n15541_));
  AOI21_X1   g12618(.A1(new_n7833_), .A2(new_n7067_), .B(pi0832), .ZN(new_n15542_));
  AOI21_X1   g12619(.A1(new_n15535_), .A2(new_n15351_), .B(new_n15519_), .ZN(new_n15543_));
  MUX2_X1    g12620(.I0(new_n15543_), .I1(pi0149), .S(new_n2926_), .Z(new_n15544_));
  AOI22_X1   g12621(.A1(new_n15541_), .A2(new_n15542_), .B1(pi0832), .B2(new_n15544_), .ZN(po0306));
  INV_X1     g12622(.I(pi0751), .ZN(new_n15546_));
  NAND4_X1   g12623(.A1(new_n15442_), .A2(new_n10038_), .A3(new_n15546_), .A4(new_n12793_), .ZN(new_n15547_));
  NAND2_X1   g12624(.A1(new_n12852_), .A2(new_n15546_), .ZN(new_n15548_));
  OAI21_X1   g12625(.A1(pi0150), .A2(new_n12852_), .B(new_n15548_), .ZN(new_n15549_));
  NOR2_X1    g12626(.A1(new_n12898_), .A2(new_n10038_), .ZN(new_n15550_));
  NOR2_X1    g12627(.A1(new_n5473_), .A2(pi0751), .ZN(new_n15551_));
  NOR2_X1    g12628(.A1(new_n13368_), .A2(new_n15551_), .ZN(new_n15552_));
  NOR4_X1    g12629(.A1(new_n15550_), .A2(pi0038), .A3(pi0701), .A4(new_n15552_), .ZN(new_n15553_));
  OAI21_X1   g12630(.A1(new_n15549_), .A2(new_n15429_), .B(new_n15553_), .ZN(new_n15554_));
  AOI21_X1   g12631(.A1(new_n15547_), .A2(new_n3154_), .B(new_n15554_), .ZN(new_n15555_));
  OAI21_X1   g12632(.A1(new_n15369_), .A2(new_n15379_), .B(pi0150), .ZN(new_n15556_));
  NOR2_X1    g12633(.A1(new_n15556_), .A2(new_n15546_), .ZN(new_n15557_));
  AOI21_X1   g12634(.A1(new_n15515_), .A2(pi0150), .B(pi0751), .ZN(new_n15558_));
  OAI21_X1   g12635(.A1(new_n15399_), .A2(new_n10038_), .B(new_n15558_), .ZN(new_n15559_));
  OAI21_X1   g12636(.A1(new_n15557_), .A2(new_n15559_), .B(pi0039), .ZN(new_n15560_));
  NOR4_X1    g12637(.A1(new_n12852_), .A2(new_n15546_), .A3(pi0907), .A4(new_n5473_), .ZN(new_n15561_));
  OAI21_X1   g12638(.A1(new_n12697_), .A2(pi0150), .B(new_n2544_), .ZN(new_n15562_));
  NOR2_X1    g12639(.A1(new_n15562_), .A2(new_n15561_), .ZN(new_n15563_));
  INV_X1     g12640(.I(pi0701), .ZN(new_n15564_));
  NOR2_X1    g12641(.A1(new_n12828_), .A2(pi0150), .ZN(new_n15565_));
  NAND3_X1   g12642(.A1(new_n3154_), .A2(pi0751), .A3(pi0947), .ZN(new_n15566_));
  OAI21_X1   g12643(.A1(new_n15523_), .A2(new_n15566_), .B(pi0038), .ZN(new_n15567_));
  OAI21_X1   g12644(.A1(new_n15565_), .A2(new_n15567_), .B(new_n15564_), .ZN(new_n15568_));
  AOI21_X1   g12645(.A1(new_n15560_), .A2(new_n15563_), .B(new_n15568_), .ZN(new_n15569_));
  OAI21_X1   g12646(.A1(new_n15569_), .A2(new_n15555_), .B(new_n7832_), .ZN(new_n15570_));
  AOI21_X1   g12647(.A1(new_n7833_), .A2(new_n10038_), .B(pi0832), .ZN(new_n15571_));
  NOR3_X1    g12648(.A1(new_n15305_), .A2(pi0701), .A3(pi0947), .ZN(new_n15572_));
  XOR2_X1    g12649(.A1(new_n15572_), .A2(new_n15551_), .Z(new_n15573_));
  MUX2_X1    g12650(.I0(new_n15573_), .I1(pi0150), .S(new_n2926_), .Z(new_n15574_));
  AOI22_X1   g12651(.A1(new_n15570_), .A2(new_n15571_), .B1(pi0832), .B2(new_n15574_), .ZN(po0307));
  AOI21_X1   g12652(.A1(pi0745), .A2(new_n12885_), .B(new_n12893_), .ZN(new_n15576_));
  NOR2_X1    g12653(.A1(new_n15576_), .A2(pi0151), .ZN(new_n15577_));
  INV_X1     g12654(.I(new_n15438_), .ZN(new_n15578_));
  NOR2_X1    g12655(.A1(new_n12745_), .A2(new_n15431_), .ZN(new_n15579_));
  AOI21_X1   g12656(.A1(new_n15579_), .A2(new_n3417_), .B(new_n12709_), .ZN(new_n15580_));
  NOR3_X1    g12657(.A1(new_n15580_), .A2(new_n2566_), .A3(new_n15431_), .ZN(new_n15581_));
  NOR2_X1    g12658(.A1(new_n12767_), .A2(new_n5092_), .ZN(new_n15582_));
  NOR2_X1    g12659(.A1(new_n15582_), .A2(new_n3417_), .ZN(new_n15583_));
  OAI21_X1   g12660(.A1(new_n15356_), .A2(new_n15583_), .B(new_n3285_), .ZN(new_n15584_));
  NAND2_X1   g12661(.A1(new_n12133_), .A2(new_n3417_), .ZN(new_n15585_));
  NAND4_X1   g12662(.A1(new_n15584_), .A2(new_n2587_), .A3(new_n15453_), .A4(new_n15585_), .ZN(new_n15586_));
  NOR3_X1    g12663(.A1(new_n15578_), .A2(new_n15581_), .A3(new_n15586_), .ZN(new_n15587_));
  NOR3_X1    g12664(.A1(new_n15587_), .A2(pi0745), .A3(new_n15451_), .ZN(new_n15588_));
  NOR4_X1    g12665(.A1(new_n15588_), .A2(pi0038), .A3(new_n3154_), .A4(new_n15577_), .ZN(new_n15589_));
  NOR2_X1    g12666(.A1(new_n12898_), .A2(new_n3417_), .ZN(new_n15590_));
  NOR2_X1    g12667(.A1(new_n5473_), .A2(pi0745), .ZN(new_n15591_));
  NOR2_X1    g12668(.A1(new_n13368_), .A2(new_n15591_), .ZN(new_n15592_));
  INV_X1     g12669(.I(pi0723), .ZN(new_n15593_));
  NAND2_X1   g12670(.A1(new_n3172_), .A2(new_n15593_), .ZN(new_n15594_));
  NOR4_X1    g12671(.A1(new_n15589_), .A2(new_n15590_), .A3(new_n15592_), .A4(new_n15594_), .ZN(new_n15595_));
  INV_X1     g12672(.I(pi0745), .ZN(new_n15596_));
  NOR2_X1    g12673(.A1(new_n15409_), .A2(new_n3417_), .ZN(new_n15597_));
  NOR2_X1    g12674(.A1(new_n12133_), .A2(new_n15372_), .ZN(new_n15598_));
  NOR2_X1    g12675(.A1(new_n15598_), .A2(new_n3285_), .ZN(new_n15599_));
  NAND2_X1   g12676(.A1(new_n15599_), .A2(new_n15585_), .ZN(new_n15600_));
  OAI21_X1   g12677(.A1(new_n15600_), .A2(new_n15411_), .B(new_n2566_), .ZN(new_n15601_));
  NOR2_X1    g12678(.A1(new_n15580_), .A2(new_n2566_), .ZN(new_n15602_));
  NOR3_X1    g12679(.A1(new_n15602_), .A2(new_n15584_), .A3(new_n15601_), .ZN(new_n15603_));
  NOR2_X1    g12680(.A1(new_n15584_), .A2(new_n15601_), .ZN(new_n15604_));
  INV_X1     g12681(.I(new_n15602_), .ZN(new_n15605_));
  OAI21_X1   g12682(.A1(new_n15605_), .A2(new_n15604_), .B(pi0299), .ZN(new_n15606_));
  OAI22_X1   g12683(.A1(new_n15396_), .A2(new_n15597_), .B1(new_n15603_), .B2(new_n15606_), .ZN(new_n15607_));
  INV_X1     g12684(.I(new_n15366_), .ZN(new_n15608_));
  NAND3_X1   g12685(.A1(new_n15360_), .A2(new_n2566_), .A3(new_n15600_), .ZN(new_n15609_));
  OAI21_X1   g12686(.A1(new_n15609_), .A2(new_n15584_), .B(new_n15605_), .ZN(new_n15610_));
  AOI21_X1   g12687(.A1(new_n15376_), .A2(new_n3417_), .B(pi0745), .ZN(new_n15611_));
  NAND2_X1   g12688(.A1(new_n15378_), .A2(new_n15611_), .ZN(new_n15612_));
  NAND4_X1   g12689(.A1(new_n15610_), .A2(new_n6593_), .A3(new_n15608_), .A4(new_n15612_), .ZN(new_n15613_));
  AOI21_X1   g12690(.A1(new_n15596_), .A2(new_n15607_), .B(new_n15613_), .ZN(new_n15614_));
  NOR2_X1    g12691(.A1(new_n12828_), .A2(pi0151), .ZN(new_n15615_));
  NAND3_X1   g12692(.A1(new_n3154_), .A2(pi0745), .A3(pi0947), .ZN(new_n15616_));
  OAI21_X1   g12693(.A1(new_n15523_), .A2(new_n15616_), .B(pi0038), .ZN(new_n15617_));
  OAI21_X1   g12694(.A1(new_n15615_), .A2(new_n15617_), .B(new_n15593_), .ZN(new_n15618_));
  AOI21_X1   g12695(.A1(new_n15614_), .A2(new_n3172_), .B(new_n15618_), .ZN(new_n15619_));
  OAI21_X1   g12696(.A1(new_n15619_), .A2(new_n15595_), .B(new_n7832_), .ZN(new_n15620_));
  AOI21_X1   g12697(.A1(new_n7833_), .A2(new_n3417_), .B(pi0832), .ZN(new_n15621_));
  NOR3_X1    g12698(.A1(new_n15305_), .A2(pi0723), .A3(pi0947), .ZN(new_n15622_));
  XOR2_X1    g12699(.A1(new_n15622_), .A2(new_n15591_), .Z(new_n15623_));
  MUX2_X1    g12700(.I0(new_n15623_), .I1(pi0151), .S(new_n2926_), .Z(new_n15624_));
  AOI22_X1   g12701(.A1(new_n15620_), .A2(new_n15621_), .B1(pi0832), .B2(new_n15624_), .ZN(po0308));
  AOI21_X1   g12702(.A1(new_n3250_), .A2(new_n12855_), .B(new_n15433_), .ZN(new_n15626_));
  INV_X1     g12703(.I(new_n15410_), .ZN(new_n15627_));
  NAND2_X1   g12704(.A1(new_n15627_), .A2(new_n15372_), .ZN(new_n15628_));
  NAND2_X1   g12705(.A1(new_n15626_), .A2(new_n15628_), .ZN(new_n15629_));
  NOR2_X1    g12706(.A1(new_n15435_), .A2(new_n3284_), .ZN(new_n15630_));
  INV_X1     g12707(.I(new_n15630_), .ZN(new_n15631_));
  AOI21_X1   g12708(.A1(new_n15358_), .A2(pi0152), .B(new_n15631_), .ZN(new_n15632_));
  NAND2_X1   g12709(.A1(new_n12133_), .A2(pi0152), .ZN(new_n15633_));
  OAI21_X1   g12710(.A1(new_n5092_), .A2(new_n12133_), .B(new_n15633_), .ZN(new_n15634_));
  AOI21_X1   g12711(.A1(new_n15634_), .A2(new_n3285_), .B(pi0215), .ZN(new_n15635_));
  OR3_X2     g12712(.A1(new_n15632_), .A2(new_n15361_), .A3(new_n15635_), .Z(new_n15636_));
  AOI21_X1   g12713(.A1(new_n15636_), .A2(new_n15629_), .B(pi0299), .ZN(new_n15637_));
  NOR2_X1    g12714(.A1(new_n12767_), .A2(new_n5141_), .ZN(new_n15638_));
  NOR2_X1    g12715(.A1(new_n12879_), .A2(new_n6460_), .ZN(new_n15639_));
  NOR2_X1    g12716(.A1(new_n15639_), .A2(new_n15638_), .ZN(new_n15640_));
  AOI21_X1   g12717(.A1(new_n15640_), .A2(new_n3250_), .B(new_n2614_), .ZN(new_n15641_));
  NOR2_X1    g12718(.A1(new_n15640_), .A2(new_n15351_), .ZN(new_n15642_));
  INV_X1     g12719(.I(new_n15642_), .ZN(new_n15643_));
  INV_X1     g12720(.I(new_n15598_), .ZN(new_n15644_));
  NAND2_X1   g12721(.A1(new_n15644_), .A2(new_n15633_), .ZN(new_n15645_));
  AOI22_X1   g12722(.A1(new_n15643_), .A2(new_n15641_), .B1(new_n2614_), .B2(new_n15645_), .ZN(new_n15646_));
  NAND2_X1   g12723(.A1(new_n15389_), .A2(new_n3250_), .ZN(new_n15647_));
  AOI21_X1   g12724(.A1(new_n15393_), .A2(new_n15647_), .B(pi0299), .ZN(new_n15648_));
  OAI21_X1   g12725(.A1(new_n15646_), .A2(pi0223), .B(new_n15648_), .ZN(new_n15649_));
  OAI21_X1   g12726(.A1(new_n15637_), .A2(pi0759), .B(new_n15649_), .ZN(new_n15650_));
  INV_X1     g12727(.I(new_n13820_), .ZN(new_n15651_));
  NOR2_X1    g12728(.A1(new_n15640_), .A2(pi0947), .ZN(new_n15652_));
  INV_X1     g12729(.I(new_n15652_), .ZN(new_n15653_));
  INV_X1     g12730(.I(new_n15640_), .ZN(new_n15654_));
  AOI21_X1   g12731(.A1(new_n15654_), .A2(new_n5093_), .B(new_n2614_), .ZN(new_n15655_));
  INV_X1     g12732(.I(new_n15655_), .ZN(new_n15656_));
  NAND3_X1   g12733(.A1(new_n15656_), .A2(new_n15641_), .A3(new_n15653_), .ZN(new_n15657_));
  OAI21_X1   g12734(.A1(new_n15634_), .A2(new_n3155_), .B(new_n2604_), .ZN(new_n15658_));
  AOI21_X1   g12735(.A1(new_n15393_), .A2(new_n15647_), .B(new_n15658_), .ZN(new_n15659_));
  INV_X1     g12736(.I(pi0759), .ZN(new_n15660_));
  AOI21_X1   g12737(.A1(new_n15391_), .A2(new_n15647_), .B(pi0299), .ZN(new_n15661_));
  NAND2_X1   g12738(.A1(new_n15661_), .A2(new_n15660_), .ZN(new_n15662_));
  AOI21_X1   g12739(.A1(new_n15657_), .A2(new_n15659_), .B(new_n15662_), .ZN(new_n15663_));
  INV_X1     g12740(.I(new_n15582_), .ZN(new_n15664_));
  AOI21_X1   g12741(.A1(new_n15632_), .A2(new_n15664_), .B(new_n15635_), .ZN(new_n15665_));
  NOR4_X1    g12742(.A1(new_n15663_), .A2(new_n15651_), .A3(new_n15626_), .A4(new_n15665_), .ZN(new_n15666_));
  NOR2_X1    g12743(.A1(new_n15660_), .A2(new_n5473_), .ZN(new_n15667_));
  OAI21_X1   g12744(.A1(new_n12852_), .A2(pi0152), .B(new_n15667_), .ZN(new_n15668_));
  OR3_X2     g12745(.A1(new_n12852_), .A2(new_n3250_), .A3(new_n15667_), .Z(new_n15669_));
  NAND4_X1   g12746(.A1(new_n15669_), .A2(new_n15668_), .A3(new_n15373_), .A4(new_n3154_), .ZN(new_n15670_));
  NOR2_X1    g12747(.A1(new_n12828_), .A2(pi0152), .ZN(new_n15671_));
  NOR2_X1    g12748(.A1(new_n12110_), .A2(new_n15351_), .ZN(new_n15672_));
  NOR2_X1    g12749(.A1(new_n15667_), .A2(pi0039), .ZN(new_n15673_));
  INV_X1     g12750(.I(pi0696), .ZN(new_n15674_));
  NAND2_X1   g12751(.A1(new_n3172_), .A2(new_n15674_), .ZN(new_n15675_));
  NOR4_X1    g12752(.A1(new_n15671_), .A2(new_n15672_), .A3(new_n15673_), .A4(new_n15675_), .ZN(new_n15676_));
  NAND2_X1   g12753(.A1(new_n15670_), .A2(new_n15676_), .ZN(new_n15677_));
  AOI21_X1   g12754(.A1(new_n15666_), .A2(new_n15650_), .B(new_n15677_), .ZN(new_n15678_));
  NOR2_X1    g12755(.A1(new_n12894_), .A2(pi0759), .ZN(new_n15679_));
  NOR3_X1    g12756(.A1(new_n15679_), .A2(pi0039), .A3(pi0152), .ZN(new_n15680_));
  INV_X1     g12757(.I(new_n15357_), .ZN(new_n15681_));
  OR2_X2     g12758(.A1(new_n15632_), .A2(new_n15437_), .Z(new_n15682_));
  NOR2_X1    g12759(.A1(new_n15366_), .A2(new_n2587_), .ZN(new_n15683_));
  INV_X1     g12760(.I(new_n15452_), .ZN(new_n15684_));
  NAND2_X1   g12761(.A1(new_n15684_), .A2(new_n15633_), .ZN(new_n15685_));
  NOR2_X1    g12762(.A1(new_n15685_), .A2(new_n3285_), .ZN(new_n15686_));
  NOR4_X1    g12763(.A1(new_n15683_), .A2(new_n3250_), .A3(pi0215), .A4(new_n15686_), .ZN(new_n15687_));
  NAND2_X1   g12764(.A1(new_n15434_), .A2(new_n15687_), .ZN(new_n15688_));
  AOI21_X1   g12765(.A1(new_n15682_), .A2(new_n15681_), .B(new_n15688_), .ZN(new_n15689_));
  AOI22_X1   g12766(.A1(new_n15653_), .A2(new_n15641_), .B1(new_n2614_), .B2(new_n15685_), .ZN(new_n15690_));
  NOR2_X1    g12767(.A1(new_n15661_), .A2(pi0759), .ZN(new_n15691_));
  OAI21_X1   g12768(.A1(new_n15690_), .A2(pi0223), .B(new_n15691_), .ZN(new_n15692_));
  NOR3_X1    g12769(.A1(new_n15692_), .A2(new_n15689_), .A3(new_n15680_), .ZN(new_n15693_));
  NOR2_X1    g12770(.A1(new_n15674_), .A2(pi0038), .ZN(new_n15695_));
  NAND4_X1   g12771(.A1(new_n15669_), .A2(new_n15668_), .A3(new_n3154_), .A4(new_n15695_), .ZN(new_n15696_));
  OAI21_X1   g12772(.A1(new_n15693_), .A2(new_n15696_), .B(new_n7832_), .ZN(new_n15697_));
  NOR2_X1    g12773(.A1(new_n15678_), .A2(new_n15697_), .ZN(new_n15698_));
  OAI21_X1   g12774(.A1(new_n7832_), .A2(pi0152), .B(new_n13184_), .ZN(new_n15699_));
  NOR4_X1    g12775(.A1(new_n15372_), .A2(new_n15674_), .A3(new_n2925_), .A4(new_n15667_), .ZN(new_n15700_));
  OAI21_X1   g12776(.A1(new_n2925_), .A2(pi0152), .B(pi0832), .ZN(new_n15701_));
  OAI22_X1   g12777(.A1(new_n15698_), .A2(new_n15699_), .B1(new_n15700_), .B2(new_n15701_), .ZN(po0309));
  OAI21_X1   g12778(.A1(new_n2925_), .A2(new_n2526_), .B(pi0832), .ZN(new_n15703_));
  AOI21_X1   g12779(.A1(pi0766), .A2(pi0947), .B(new_n2926_), .ZN(new_n15704_));
  INV_X1     g12780(.I(new_n15704_), .ZN(new_n15705_));
  NAND4_X1   g12781(.A1(new_n15705_), .A2(pi0700), .A3(new_n15703_), .A4(new_n15351_), .ZN(new_n15706_));
  INV_X1     g12782(.I(pi0766), .ZN(new_n15707_));
  NOR4_X1    g12783(.A1(new_n15523_), .A2(pi0039), .A3(new_n15707_), .A4(pi0947), .ZN(new_n15708_));
  NOR2_X1    g12784(.A1(new_n15708_), .A2(new_n3172_), .ZN(new_n15709_));
  OAI21_X1   g12785(.A1(pi0153), .A2(new_n12828_), .B(new_n15709_), .ZN(new_n15710_));
  NAND2_X1   g12786(.A1(new_n12855_), .A2(pi0153), .ZN(new_n15711_));
  NAND2_X1   g12787(.A1(new_n15432_), .A2(new_n15711_), .ZN(new_n15712_));
  NOR2_X1    g12788(.A1(new_n15582_), .A2(new_n2526_), .ZN(new_n15713_));
  OAI21_X1   g12789(.A1(new_n15356_), .A2(new_n15713_), .B(new_n3285_), .ZN(new_n15714_));
  OAI21_X1   g12790(.A1(pi0153), .A2(new_n12132_), .B(new_n15453_), .ZN(new_n15715_));
  NOR2_X1    g12791(.A1(new_n12133_), .A2(new_n15305_), .ZN(new_n15716_));
  AOI21_X1   g12792(.A1(new_n15715_), .A2(new_n15716_), .B(pi0215), .ZN(new_n15717_));
  OAI21_X1   g12793(.A1(new_n15714_), .A2(new_n15717_), .B(new_n15712_), .ZN(new_n15718_));
  NOR2_X1    g12794(.A1(new_n15409_), .A2(new_n2526_), .ZN(new_n15719_));
  AOI22_X1   g12795(.A1(new_n15396_), .A2(new_n15719_), .B1(pi0299), .B2(new_n15718_), .ZN(new_n15720_));
  INV_X1     g12796(.I(new_n15714_), .ZN(new_n15721_));
  INV_X1     g12797(.I(new_n15599_), .ZN(new_n15722_));
  AOI21_X1   g12798(.A1(new_n2526_), .A2(new_n12133_), .B(new_n15722_), .ZN(new_n15723_));
  OAI21_X1   g12799(.A1(new_n15359_), .A2(new_n15723_), .B(new_n15721_), .ZN(new_n15724_));
  NAND2_X1   g12800(.A1(new_n15712_), .A2(new_n15410_), .ZN(new_n15725_));
  NOR2_X1    g12801(.A1(new_n15366_), .A2(pi0299), .ZN(new_n15726_));
  NAND2_X1   g12802(.A1(new_n15725_), .A2(new_n15726_), .ZN(new_n15727_));
  AOI21_X1   g12803(.A1(new_n15724_), .A2(new_n2566_), .B(new_n15727_), .ZN(new_n15728_));
  INV_X1     g12804(.I(new_n15378_), .ZN(new_n15729_));
  NOR2_X1    g12805(.A1(new_n12792_), .A2(pi0153), .ZN(new_n15730_));
  NOR2_X1    g12806(.A1(pi0039), .A2(pi0766), .ZN(new_n15731_));
  OAI21_X1   g12807(.A1(new_n15729_), .A2(new_n15730_), .B(new_n15731_), .ZN(new_n15732_));
  NOR3_X1    g12808(.A1(new_n15720_), .A2(new_n15728_), .A3(new_n15732_), .ZN(new_n15733_));
  INV_X1     g12809(.I(new_n13384_), .ZN(new_n15734_));
  NOR2_X1    g12810(.A1(new_n15734_), .A2(pi0766), .ZN(new_n15735_));
  OAI22_X1   g12811(.A1(new_n15735_), .A2(new_n15448_), .B1(pi0153), .B2(new_n12852_), .ZN(new_n15736_));
  NOR2_X1    g12812(.A1(new_n15736_), .A2(new_n15373_), .ZN(new_n15737_));
  OAI21_X1   g12813(.A1(new_n15733_), .A2(new_n15737_), .B(new_n3172_), .ZN(new_n15738_));
  NAND2_X1   g12814(.A1(new_n2526_), .A2(new_n15707_), .ZN(new_n15739_));
  OAI21_X1   g12815(.A1(new_n12894_), .A2(new_n15739_), .B(pi0039), .ZN(new_n15740_));
  NOR3_X1    g12816(.A1(new_n15434_), .A2(pi0299), .A3(new_n15711_), .ZN(new_n15741_));
  NAND2_X1   g12817(.A1(new_n15715_), .A2(new_n15707_), .ZN(new_n15742_));
  NOR4_X1    g12818(.A1(new_n15578_), .A2(new_n15714_), .A3(new_n15741_), .A4(new_n15742_), .ZN(new_n15743_));
  NOR3_X1    g12819(.A1(new_n15743_), .A2(new_n15494_), .A3(new_n15730_), .ZN(new_n15744_));
  INV_X1     g12820(.I(pi0700), .ZN(new_n15745_));
  NAND2_X1   g12821(.A1(new_n5156_), .A2(new_n15704_), .ZN(new_n15746_));
  NAND4_X1   g12822(.A1(new_n12898_), .A2(new_n3172_), .A3(new_n2526_), .A4(new_n15746_), .ZN(new_n15747_));
  NAND4_X1   g12823(.A1(new_n15736_), .A2(new_n3172_), .A3(new_n15745_), .A4(new_n15747_), .ZN(new_n15748_));
  AOI21_X1   g12824(.A1(new_n15744_), .A2(new_n15740_), .B(new_n15748_), .ZN(new_n15749_));
  OAI21_X1   g12825(.A1(new_n15749_), .A2(new_n15500_), .B(pi0700), .ZN(new_n15750_));
  AOI21_X1   g12826(.A1(new_n15738_), .A2(new_n15710_), .B(new_n15750_), .ZN(new_n15751_));
  NAND2_X1   g12827(.A1(pi0057), .A2(pi0153), .ZN(new_n15752_));
  AOI21_X1   g12828(.A1(new_n15752_), .A2(new_n13184_), .B(pi0057), .ZN(new_n15753_));
  OAI21_X1   g12829(.A1(new_n15499_), .A2(pi0153), .B(new_n15753_), .ZN(new_n15754_));
  OAI21_X1   g12830(.A1(new_n15751_), .A2(new_n15754_), .B(new_n15706_), .ZN(po0310));
  INV_X1     g12831(.I(pi0704), .ZN(new_n15756_));
  NAND2_X1   g12832(.A1(new_n15756_), .A2(pi0907), .ZN(new_n15757_));
  MUX2_X1    g12833(.I0(new_n15757_), .I1(pi0742), .S(pi0947), .Z(new_n15758_));
  MUX2_X1    g12834(.I0(new_n15758_), .I1(new_n3271_), .S(new_n2926_), .Z(new_n15759_));
  XOR2_X1    g12835(.A1(new_n15442_), .A2(new_n15458_), .Z(new_n15760_));
  NAND2_X1   g12836(.A1(new_n15760_), .A2(new_n3271_), .ZN(new_n15761_));
  XOR2_X1    g12837(.A1(new_n15761_), .A2(new_n15458_), .Z(new_n15762_));
  NOR2_X1    g12838(.A1(new_n12852_), .A2(pi0154), .ZN(new_n15763_));
  INV_X1     g12839(.I(pi0742), .ZN(new_n15764_));
  NOR2_X1    g12840(.A1(new_n15764_), .A2(pi0038), .ZN(new_n15766_));
  OAI21_X1   g12841(.A1(new_n15449_), .A2(new_n15763_), .B(new_n15766_), .ZN(new_n15767_));
  AOI21_X1   g12842(.A1(new_n15762_), .A2(pi0039), .B(new_n15767_), .ZN(new_n15768_));
  NOR2_X1    g12843(.A1(new_n12902_), .A2(pi0154), .ZN(new_n15769_));
  NOR4_X1    g12844(.A1(new_n15768_), .A2(pi0704), .A3(pi0742), .A4(new_n15769_), .ZN(new_n15770_));
  OAI21_X1   g12845(.A1(new_n15400_), .A2(new_n15515_), .B(pi0154), .ZN(new_n15771_));
  NOR2_X1    g12846(.A1(new_n15771_), .A2(new_n3154_), .ZN(new_n15772_));
  NOR4_X1    g12847(.A1(new_n15373_), .A2(new_n15406_), .A3(new_n15763_), .A4(pi0039), .ZN(new_n15773_));
  NOR2_X1    g12848(.A1(new_n12828_), .A2(pi0154), .ZN(new_n15774_));
  NOR2_X1    g12849(.A1(pi0038), .A2(pi0742), .ZN(new_n15775_));
  OAI21_X1   g12850(.A1(new_n15772_), .A2(new_n15773_), .B(new_n15775_), .ZN(new_n15776_));
  NOR3_X1    g12851(.A1(new_n15373_), .A2(new_n15763_), .A3(pi0039), .ZN(new_n15777_));
  NOR4_X1    g12852(.A1(new_n15473_), .A2(pi0039), .A3(new_n3271_), .A4(new_n15379_), .ZN(new_n15778_));
  NOR2_X1    g12853(.A1(new_n15381_), .A2(new_n3172_), .ZN(new_n15779_));
  NOR2_X1    g12854(.A1(new_n15774_), .A2(pi0742), .ZN(new_n15780_));
  AOI21_X1   g12855(.A1(new_n15779_), .A2(new_n15780_), .B(pi0038), .ZN(new_n15781_));
  OAI21_X1   g12856(.A1(new_n15778_), .A2(new_n15777_), .B(new_n15781_), .ZN(new_n15782_));
  OAI21_X1   g12857(.A1(new_n7832_), .A2(pi0154), .B(new_n13184_), .ZN(new_n15783_));
  NOR2_X1    g12858(.A1(new_n7833_), .A2(pi0704), .ZN(new_n15784_));
  NAND4_X1   g12859(.A1(new_n15782_), .A2(new_n15776_), .A3(new_n15783_), .A4(new_n15784_), .ZN(new_n15785_));
  OAI22_X1   g12860(.A1(new_n15770_), .A2(new_n15785_), .B1(new_n13184_), .B2(new_n15759_), .ZN(po0311));
  INV_X1     g12861(.I(pi0757), .ZN(new_n15787_));
  NOR2_X1    g12862(.A1(new_n15305_), .A2(pi0686), .ZN(new_n15788_));
  MUX2_X1    g12863(.I0(new_n15788_), .I1(new_n15787_), .S(pi0947), .Z(new_n15789_));
  MUX2_X1    g12864(.I0(new_n15789_), .I1(pi0155), .S(new_n2926_), .Z(new_n15790_));
  NAND3_X1   g12865(.A1(new_n15445_), .A2(new_n15787_), .A3(new_n12902_), .ZN(new_n15791_));
  OAI21_X1   g12866(.A1(pi0757), .A2(new_n12902_), .B(new_n15444_), .ZN(new_n15792_));
  AOI21_X1   g12867(.A1(new_n15791_), .A2(new_n15792_), .B(pi0686), .ZN(new_n15793_));
  INV_X1     g12868(.I(pi0686), .ZN(new_n15794_));
  NOR2_X1    g12869(.A1(new_n15421_), .A2(new_n3172_), .ZN(new_n15795_));
  AOI21_X1   g12870(.A1(new_n15404_), .A2(new_n3172_), .B(new_n15795_), .ZN(new_n15796_));
  OAI21_X1   g12871(.A1(new_n15796_), .A2(pi0757), .B(new_n15794_), .ZN(new_n15797_));
  NOR2_X1    g12872(.A1(new_n7833_), .A2(pi0155), .ZN(new_n15798_));
  OAI21_X1   g12873(.A1(new_n15797_), .A2(new_n15793_), .B(new_n15798_), .ZN(new_n15799_));
  AOI21_X1   g12874(.A1(new_n12828_), .A2(new_n5093_), .B(new_n3172_), .ZN(new_n15800_));
  AOI21_X1   g12875(.A1(new_n15420_), .A2(new_n3172_), .B(new_n15800_), .ZN(new_n15801_));
  INV_X1     g12876(.I(new_n15801_), .ZN(new_n15802_));
  NAND2_X1   g12877(.A1(new_n15802_), .A2(pi0757), .ZN(new_n15803_));
  AOI21_X1   g12878(.A1(new_n15380_), .A2(new_n3172_), .B(new_n15779_), .ZN(new_n15804_));
  INV_X1     g12879(.I(new_n15804_), .ZN(new_n15805_));
  NOR2_X1    g12880(.A1(new_n15805_), .A2(new_n15787_), .ZN(new_n15806_));
  NAND4_X1   g12881(.A1(new_n7833_), .A2(new_n7639_), .A3(new_n15794_), .A4(new_n15787_), .ZN(new_n15807_));
  NOR3_X1    g12882(.A1(new_n15806_), .A2(new_n15461_), .A3(new_n15807_), .ZN(new_n15808_));
  AOI21_X1   g12883(.A1(new_n15808_), .A2(new_n15803_), .B(pi0832), .ZN(new_n15809_));
  AOI22_X1   g12884(.A1(new_n15799_), .A2(new_n15809_), .B1(pi0832), .B2(new_n15790_), .ZN(po0312));
  INV_X1     g12885(.I(pi0724), .ZN(new_n15811_));
  NAND2_X1   g12886(.A1(new_n15811_), .A2(pi0907), .ZN(new_n15812_));
  MUX2_X1    g12887(.I0(new_n15812_), .I1(pi0741), .S(pi0947), .Z(new_n15813_));
  MUX2_X1    g12888(.I0(new_n15813_), .I1(new_n8974_), .S(new_n2926_), .Z(new_n15814_));
  INV_X1     g12889(.I(pi0741), .ZN(new_n15815_));
  NOR3_X1    g12890(.A1(new_n15801_), .A2(new_n15805_), .A3(new_n15815_), .ZN(new_n15816_));
  AOI21_X1   g12891(.A1(pi0741), .A2(new_n15805_), .B(new_n15802_), .ZN(new_n15817_));
  OAI21_X1   g12892(.A1(new_n15817_), .A2(new_n15816_), .B(new_n15811_), .ZN(new_n15818_));
  NOR3_X1    g12893(.A1(new_n15461_), .A2(new_n15811_), .A3(pi0741), .ZN(new_n15819_));
  NOR3_X1    g12894(.A1(new_n15819_), .A2(new_n8974_), .A3(new_n7833_), .ZN(new_n15820_));
  AOI21_X1   g12895(.A1(new_n15818_), .A2(new_n15820_), .B(pi0832), .ZN(new_n15821_));
  AOI21_X1   g12896(.A1(new_n15445_), .A2(new_n15815_), .B(new_n12902_), .ZN(new_n15822_));
  AOI21_X1   g12897(.A1(new_n15144_), .A2(new_n3172_), .B(new_n12900_), .ZN(new_n15823_));
  NOR3_X1    g12898(.A1(new_n15445_), .A2(pi0741), .A3(new_n15823_), .ZN(new_n15824_));
  OAI21_X1   g12899(.A1(new_n15824_), .A2(new_n15822_), .B(pi0724), .ZN(new_n15825_));
  NOR3_X1    g12900(.A1(new_n15796_), .A2(pi0724), .A3(pi0741), .ZN(new_n15826_));
  NOR2_X1    g12901(.A1(new_n15826_), .A2(new_n7833_), .ZN(new_n15827_));
  AOI21_X1   g12902(.A1(new_n15827_), .A2(new_n15825_), .B(pi0156), .ZN(new_n15828_));
  OAI22_X1   g12903(.A1(new_n15828_), .A2(new_n15821_), .B1(new_n13184_), .B2(new_n15814_), .ZN(po0313));
  INV_X1     g12904(.I(pi0688), .ZN(new_n15830_));
  INV_X1     g12905(.I(pi0760), .ZN(new_n15831_));
  NAND3_X1   g12906(.A1(new_n15473_), .A2(new_n15831_), .A3(new_n15399_), .ZN(new_n15832_));
  OAI21_X1   g12907(.A1(pi0760), .A2(new_n15399_), .B(new_n15369_), .ZN(new_n15833_));
  INV_X1     g12908(.I(new_n15379_), .ZN(new_n15834_));
  NOR3_X1    g12909(.A1(new_n15515_), .A2(pi0760), .A3(new_n15834_), .ZN(new_n15835_));
  AOI21_X1   g12910(.A1(new_n15831_), .A2(new_n15834_), .B(new_n15419_), .ZN(new_n15836_));
  NOR4_X1    g12911(.A1(new_n15835_), .A2(new_n3154_), .A3(pi0157), .A4(new_n15836_), .ZN(new_n15837_));
  NAND3_X1   g12912(.A1(new_n15832_), .A2(new_n15833_), .A3(new_n15837_), .ZN(new_n15838_));
  OAI21_X1   g12913(.A1(new_n12852_), .A2(pi0157), .B(new_n3154_), .ZN(new_n15839_));
  NOR2_X1    g12914(.A1(new_n5473_), .A2(pi0760), .ZN(new_n15840_));
  AND3_X2    g12915(.A1(new_n15839_), .A2(new_n12852_), .A3(new_n15840_), .Z(new_n15841_));
  NAND2_X1   g12916(.A1(new_n15841_), .A2(new_n15374_), .ZN(new_n15842_));
  AOI21_X1   g12917(.A1(new_n15838_), .A2(new_n15842_), .B(pi0038), .ZN(new_n15843_));
  NOR2_X1    g12918(.A1(new_n12828_), .A2(pi0157), .ZN(new_n15844_));
  NOR4_X1    g12919(.A1(new_n15523_), .A2(pi0039), .A3(new_n15831_), .A4(new_n5473_), .ZN(new_n15845_));
  NOR3_X1    g12920(.A1(new_n15844_), .A2(new_n3172_), .A3(new_n15845_), .ZN(new_n15846_));
  OAI21_X1   g12921(.A1(new_n15843_), .A2(new_n15846_), .B(new_n15830_), .ZN(new_n15847_));
  AOI21_X1   g12922(.A1(pi0157), .A2(new_n2587_), .B(new_n15457_), .ZN(new_n15848_));
  AOI21_X1   g12923(.A1(new_n15440_), .A2(new_n10117_), .B(new_n15848_), .ZN(new_n15849_));
  AOI21_X1   g12924(.A1(new_n10117_), .A2(new_n15376_), .B(new_n15494_), .ZN(new_n15850_));
  NOR3_X1    g12925(.A1(new_n15849_), .A2(pi0760), .A3(new_n15850_), .ZN(new_n15851_));
  NOR2_X1    g12926(.A1(pi0039), .A2(pi0760), .ZN(new_n15852_));
  OAI21_X1   g12927(.A1(new_n12894_), .A2(pi0157), .B(new_n15852_), .ZN(new_n15853_));
  NOR2_X1    g12928(.A1(new_n15841_), .A2(pi0038), .ZN(new_n15854_));
  OAI21_X1   g12929(.A1(new_n15851_), .A2(new_n15853_), .B(new_n15854_), .ZN(new_n15855_));
  NAND2_X1   g12930(.A1(new_n12899_), .A2(pi0157), .ZN(new_n15856_));
  NOR2_X1    g12931(.A1(new_n13368_), .A2(new_n15840_), .ZN(new_n15857_));
  NOR2_X1    g12932(.A1(new_n15857_), .A2(new_n3172_), .ZN(new_n15858_));
  AOI21_X1   g12933(.A1(new_n15856_), .A2(new_n15858_), .B(new_n15830_), .ZN(new_n15859_));
  AOI21_X1   g12934(.A1(new_n15855_), .A2(new_n15859_), .B(new_n7833_), .ZN(new_n15860_));
  NAND2_X1   g12935(.A1(new_n15847_), .A2(new_n15860_), .ZN(new_n15861_));
  AOI21_X1   g12936(.A1(new_n7833_), .A2(new_n10117_), .B(pi0832), .ZN(new_n15862_));
  AOI21_X1   g12937(.A1(new_n15830_), .A2(new_n15351_), .B(new_n15840_), .ZN(new_n15863_));
  MUX2_X1    g12938(.I0(new_n15863_), .I1(pi0157), .S(new_n2926_), .Z(new_n15864_));
  AOI22_X1   g12939(.A1(new_n15861_), .A2(new_n15862_), .B1(pi0832), .B2(new_n15864_), .ZN(po0314));
  INV_X1     g12940(.I(pi0753), .ZN(new_n15866_));
  NAND4_X1   g12941(.A1(new_n15442_), .A2(new_n5340_), .A3(new_n15866_), .A4(new_n12793_), .ZN(new_n15867_));
  NAND2_X1   g12942(.A1(new_n12852_), .A2(new_n15866_), .ZN(new_n15868_));
  OAI21_X1   g12943(.A1(pi0158), .A2(new_n12852_), .B(new_n15868_), .ZN(new_n15869_));
  NOR2_X1    g12944(.A1(new_n12898_), .A2(new_n5340_), .ZN(new_n15870_));
  NOR2_X1    g12945(.A1(new_n5473_), .A2(pi0753), .ZN(new_n15871_));
  NOR2_X1    g12946(.A1(new_n13368_), .A2(new_n15871_), .ZN(new_n15872_));
  NOR4_X1    g12947(.A1(new_n15870_), .A2(pi0038), .A3(pi0702), .A4(new_n15872_), .ZN(new_n15873_));
  OAI21_X1   g12948(.A1(new_n15869_), .A2(new_n15429_), .B(new_n15873_), .ZN(new_n15874_));
  AOI21_X1   g12949(.A1(new_n15867_), .A2(new_n3154_), .B(new_n15874_), .ZN(new_n15875_));
  OAI21_X1   g12950(.A1(new_n15369_), .A2(new_n15379_), .B(pi0158), .ZN(new_n15876_));
  NOR2_X1    g12951(.A1(new_n15876_), .A2(new_n15866_), .ZN(new_n15877_));
  AOI21_X1   g12952(.A1(new_n15515_), .A2(pi0158), .B(pi0753), .ZN(new_n15878_));
  OAI21_X1   g12953(.A1(new_n15399_), .A2(new_n5340_), .B(new_n15878_), .ZN(new_n15879_));
  OAI21_X1   g12954(.A1(new_n15877_), .A2(new_n15879_), .B(pi0039), .ZN(new_n15880_));
  NOR4_X1    g12955(.A1(new_n12852_), .A2(new_n15866_), .A3(pi0907), .A4(new_n5473_), .ZN(new_n15881_));
  OAI21_X1   g12956(.A1(new_n12697_), .A2(pi0158), .B(new_n2544_), .ZN(new_n15882_));
  NOR2_X1    g12957(.A1(new_n15882_), .A2(new_n15881_), .ZN(new_n15883_));
  INV_X1     g12958(.I(pi0702), .ZN(new_n15884_));
  NOR2_X1    g12959(.A1(new_n12828_), .A2(pi0158), .ZN(new_n15885_));
  NAND3_X1   g12960(.A1(new_n3154_), .A2(pi0753), .A3(pi0947), .ZN(new_n15886_));
  OAI21_X1   g12961(.A1(new_n15523_), .A2(new_n15886_), .B(pi0038), .ZN(new_n15887_));
  OAI21_X1   g12962(.A1(new_n15885_), .A2(new_n15887_), .B(new_n15884_), .ZN(new_n15888_));
  AOI21_X1   g12963(.A1(new_n15880_), .A2(new_n15883_), .B(new_n15888_), .ZN(new_n15889_));
  OAI21_X1   g12964(.A1(new_n15889_), .A2(new_n15875_), .B(new_n7832_), .ZN(new_n15890_));
  AOI21_X1   g12965(.A1(new_n7833_), .A2(new_n5340_), .B(pi0832), .ZN(new_n15891_));
  NOR3_X1    g12966(.A1(new_n15305_), .A2(pi0702), .A3(pi0947), .ZN(new_n15892_));
  XOR2_X1    g12967(.A1(new_n15892_), .A2(new_n15871_), .Z(new_n15893_));
  MUX2_X1    g12968(.I0(new_n15893_), .I1(pi0158), .S(new_n2926_), .Z(new_n15894_));
  AOI22_X1   g12969(.A1(new_n15890_), .A2(new_n15891_), .B1(pi0832), .B2(new_n15894_), .ZN(po0315));
  INV_X1     g12970(.I(pi0754), .ZN(new_n15896_));
  NAND4_X1   g12971(.A1(new_n15442_), .A2(new_n5341_), .A3(new_n15896_), .A4(new_n12793_), .ZN(new_n15897_));
  NAND2_X1   g12972(.A1(new_n12852_), .A2(new_n15896_), .ZN(new_n15898_));
  OAI21_X1   g12973(.A1(pi0159), .A2(new_n12852_), .B(new_n15898_), .ZN(new_n15899_));
  NOR2_X1    g12974(.A1(new_n12898_), .A2(new_n5341_), .ZN(new_n15900_));
  NOR2_X1    g12975(.A1(new_n5473_), .A2(pi0754), .ZN(new_n15901_));
  NOR2_X1    g12976(.A1(new_n13368_), .A2(new_n15901_), .ZN(new_n15902_));
  NOR4_X1    g12977(.A1(new_n15900_), .A2(pi0038), .A3(pi0709), .A4(new_n15902_), .ZN(new_n15903_));
  OAI21_X1   g12978(.A1(new_n15899_), .A2(new_n15429_), .B(new_n15903_), .ZN(new_n15904_));
  AOI21_X1   g12979(.A1(new_n15897_), .A2(new_n3154_), .B(new_n15904_), .ZN(new_n15905_));
  OAI21_X1   g12980(.A1(new_n15369_), .A2(new_n15379_), .B(pi0159), .ZN(new_n15906_));
  NOR2_X1    g12981(.A1(new_n15906_), .A2(new_n15896_), .ZN(new_n15907_));
  AOI21_X1   g12982(.A1(new_n15515_), .A2(pi0159), .B(pi0754), .ZN(new_n15908_));
  OAI21_X1   g12983(.A1(new_n15399_), .A2(new_n5341_), .B(new_n15908_), .ZN(new_n15909_));
  OAI21_X1   g12984(.A1(new_n15907_), .A2(new_n15909_), .B(pi0039), .ZN(new_n15910_));
  NOR4_X1    g12985(.A1(new_n12852_), .A2(new_n15896_), .A3(pi0907), .A4(new_n5473_), .ZN(new_n15911_));
  OAI21_X1   g12986(.A1(new_n12697_), .A2(pi0159), .B(new_n2544_), .ZN(new_n15912_));
  NOR2_X1    g12987(.A1(new_n15912_), .A2(new_n15911_), .ZN(new_n15913_));
  INV_X1     g12988(.I(pi0709), .ZN(new_n15914_));
  NOR2_X1    g12989(.A1(new_n12828_), .A2(pi0159), .ZN(new_n15915_));
  NAND3_X1   g12990(.A1(new_n3154_), .A2(pi0754), .A3(pi0947), .ZN(new_n15916_));
  OAI21_X1   g12991(.A1(new_n15523_), .A2(new_n15916_), .B(pi0038), .ZN(new_n15917_));
  OAI21_X1   g12992(.A1(new_n15915_), .A2(new_n15917_), .B(new_n15914_), .ZN(new_n15918_));
  AOI21_X1   g12993(.A1(new_n15910_), .A2(new_n15913_), .B(new_n15918_), .ZN(new_n15919_));
  OAI21_X1   g12994(.A1(new_n15919_), .A2(new_n15905_), .B(new_n7832_), .ZN(new_n15920_));
  AOI21_X1   g12995(.A1(new_n7833_), .A2(new_n5341_), .B(pi0832), .ZN(new_n15921_));
  NOR3_X1    g12996(.A1(new_n15305_), .A2(pi0709), .A3(pi0947), .ZN(new_n15922_));
  XOR2_X1    g12997(.A1(new_n15922_), .A2(new_n15901_), .Z(new_n15923_));
  MUX2_X1    g12998(.I0(new_n15923_), .I1(pi0159), .S(new_n2926_), .Z(new_n15924_));
  AOI22_X1   g12999(.A1(new_n15920_), .A2(new_n15921_), .B1(pi0832), .B2(new_n15924_), .ZN(po0316));
  INV_X1     g13000(.I(pi0756), .ZN(new_n15926_));
  NAND3_X1   g13001(.A1(new_n12792_), .A2(new_n5338_), .A3(new_n2587_), .ZN(new_n15927_));
  OAI21_X1   g13002(.A1(pi0160), .A2(new_n15475_), .B(new_n15368_), .ZN(new_n15928_));
  AOI22_X1   g13003(.A1(new_n15928_), .A2(new_n15927_), .B1(new_n15926_), .B2(new_n15510_), .ZN(new_n15929_));
  NAND2_X1   g13004(.A1(new_n15400_), .A2(pi0160), .ZN(new_n15930_));
  NAND2_X1   g13005(.A1(new_n15515_), .A2(pi0160), .ZN(new_n15931_));
  NAND4_X1   g13006(.A1(new_n15930_), .A2(pi0039), .A3(new_n15926_), .A4(new_n15931_), .ZN(new_n15932_));
  OAI21_X1   g13007(.A1(new_n12852_), .A2(pi0160), .B(new_n3154_), .ZN(new_n15933_));
  NOR2_X1    g13008(.A1(new_n5473_), .A2(pi0756), .ZN(new_n15934_));
  NAND3_X1   g13009(.A1(new_n15933_), .A2(new_n12852_), .A3(new_n15934_), .ZN(new_n15935_));
  OAI22_X1   g13010(.A1(new_n15932_), .A2(new_n15929_), .B1(new_n15373_), .B2(new_n15935_), .ZN(new_n15936_));
  NAND2_X1   g13011(.A1(new_n13368_), .A2(new_n5338_), .ZN(new_n15937_));
  NOR4_X1    g13012(.A1(new_n15523_), .A2(pi0039), .A3(new_n15926_), .A4(new_n5473_), .ZN(new_n15938_));
  NOR2_X1    g13013(.A1(new_n15938_), .A2(new_n3172_), .ZN(new_n15939_));
  AOI22_X1   g13014(.A1(new_n15936_), .A2(new_n3172_), .B1(new_n15937_), .B2(new_n15939_), .ZN(new_n15940_));
  OAI21_X1   g13015(.A1(new_n15440_), .A2(new_n15488_), .B(pi0160), .ZN(new_n15941_));
  NOR2_X1    g13016(.A1(new_n15941_), .A2(new_n2587_), .ZN(new_n15942_));
  AOI21_X1   g13017(.A1(new_n5338_), .A2(new_n15376_), .B(new_n15494_), .ZN(new_n15943_));
  NOR3_X1    g13018(.A1(new_n15942_), .A2(pi0756), .A3(new_n15943_), .ZN(new_n15944_));
  NOR2_X1    g13019(.A1(pi0039), .A2(pi0756), .ZN(new_n15945_));
  OAI21_X1   g13020(.A1(new_n12894_), .A2(pi0160), .B(new_n15945_), .ZN(new_n15946_));
  AND2_X2    g13021(.A1(new_n15935_), .A2(new_n3172_), .Z(new_n15947_));
  OAI21_X1   g13022(.A1(new_n15944_), .A2(new_n15946_), .B(new_n15947_), .ZN(new_n15948_));
  INV_X1     g13023(.I(pi0734), .ZN(new_n15949_));
  NAND2_X1   g13024(.A1(new_n12899_), .A2(pi0160), .ZN(new_n15950_));
  NOR2_X1    g13025(.A1(new_n13368_), .A2(new_n15934_), .ZN(new_n15951_));
  NOR2_X1    g13026(.A1(new_n15951_), .A2(new_n3172_), .ZN(new_n15952_));
  AOI21_X1   g13027(.A1(new_n15950_), .A2(new_n15952_), .B(new_n15949_), .ZN(new_n15953_));
  AOI21_X1   g13028(.A1(new_n15948_), .A2(new_n15953_), .B(new_n7833_), .ZN(new_n15954_));
  OAI21_X1   g13029(.A1(new_n15940_), .A2(pi0734), .B(new_n15954_), .ZN(new_n15955_));
  AOI21_X1   g13030(.A1(new_n7833_), .A2(new_n5338_), .B(pi0832), .ZN(new_n15956_));
  AOI21_X1   g13031(.A1(new_n15949_), .A2(new_n15351_), .B(new_n15934_), .ZN(new_n15957_));
  MUX2_X1    g13032(.I0(new_n15957_), .I1(pi0160), .S(new_n2926_), .Z(new_n15958_));
  AOI22_X1   g13033(.A1(new_n15955_), .A2(new_n15956_), .B1(pi0832), .B2(new_n15958_), .ZN(po0317));
  AOI21_X1   g13034(.A1(new_n4701_), .A2(new_n12855_), .B(new_n15433_), .ZN(new_n15960_));
  NAND2_X1   g13035(.A1(new_n15960_), .A2(new_n15628_), .ZN(new_n15961_));
  AOI21_X1   g13036(.A1(new_n15358_), .A2(pi0161), .B(new_n15631_), .ZN(new_n15962_));
  NOR2_X1    g13037(.A1(new_n12132_), .A2(new_n4701_), .ZN(new_n15963_));
  NOR2_X1    g13038(.A1(new_n15411_), .A2(new_n15963_), .ZN(new_n15964_));
  INV_X1     g13039(.I(new_n15964_), .ZN(new_n15965_));
  AOI21_X1   g13040(.A1(new_n15965_), .A2(new_n3285_), .B(pi0215), .ZN(new_n15966_));
  OR3_X2     g13041(.A1(new_n15962_), .A2(new_n15361_), .A3(new_n15966_), .Z(new_n15967_));
  AOI21_X1   g13042(.A1(new_n15967_), .A2(new_n15961_), .B(pi0299), .ZN(new_n15968_));
  INV_X1     g13043(.I(new_n15963_), .ZN(new_n15969_));
  NAND2_X1   g13044(.A1(new_n15644_), .A2(new_n15969_), .ZN(new_n15970_));
  AOI21_X1   g13045(.A1(new_n15640_), .A2(new_n4701_), .B(new_n2614_), .ZN(new_n15971_));
  AOI22_X1   g13046(.A1(new_n15643_), .A2(new_n15971_), .B1(new_n2614_), .B2(new_n15970_), .ZN(new_n15972_));
  NAND2_X1   g13047(.A1(new_n15389_), .A2(new_n4701_), .ZN(new_n15973_));
  AOI21_X1   g13048(.A1(new_n15393_), .A2(new_n15973_), .B(pi0299), .ZN(new_n15974_));
  OAI21_X1   g13049(.A1(new_n15972_), .A2(pi0223), .B(new_n15974_), .ZN(new_n15975_));
  OAI21_X1   g13050(.A1(new_n15968_), .A2(pi0758), .B(new_n15975_), .ZN(new_n15976_));
  NAND2_X1   g13051(.A1(new_n15653_), .A2(new_n15971_), .ZN(new_n15977_));
  NAND2_X1   g13052(.A1(new_n15977_), .A2(new_n15655_), .ZN(new_n15978_));
  OAI21_X1   g13053(.A1(new_n15965_), .A2(new_n3155_), .B(new_n2604_), .ZN(new_n15979_));
  AOI21_X1   g13054(.A1(new_n15393_), .A2(new_n15973_), .B(new_n15979_), .ZN(new_n15980_));
  AOI21_X1   g13055(.A1(new_n15391_), .A2(new_n15973_), .B(pi0299), .ZN(new_n15981_));
  NAND2_X1   g13056(.A1(new_n15981_), .A2(new_n14628_), .ZN(new_n15982_));
  AOI21_X1   g13057(.A1(new_n15978_), .A2(new_n15980_), .B(new_n15982_), .ZN(new_n15983_));
  AOI21_X1   g13058(.A1(new_n15962_), .A2(new_n15664_), .B(new_n15966_), .ZN(new_n15984_));
  NOR4_X1    g13059(.A1(new_n15983_), .A2(new_n15651_), .A3(new_n15960_), .A4(new_n15984_), .ZN(new_n15985_));
  NOR2_X1    g13060(.A1(new_n14628_), .A2(new_n5473_), .ZN(new_n15986_));
  OAI21_X1   g13061(.A1(new_n12852_), .A2(pi0161), .B(new_n15986_), .ZN(new_n15987_));
  OR3_X2     g13062(.A1(new_n12852_), .A2(new_n4701_), .A3(new_n15986_), .Z(new_n15988_));
  NAND4_X1   g13063(.A1(new_n15988_), .A2(new_n15987_), .A3(new_n15373_), .A4(new_n3154_), .ZN(new_n15989_));
  NOR2_X1    g13064(.A1(new_n12828_), .A2(pi0161), .ZN(new_n15990_));
  NOR2_X1    g13065(.A1(new_n15986_), .A2(pi0039), .ZN(new_n15991_));
  NAND2_X1   g13066(.A1(new_n3172_), .A2(new_n14611_), .ZN(new_n15992_));
  NOR4_X1    g13067(.A1(new_n15990_), .A2(new_n15672_), .A3(new_n15991_), .A4(new_n15992_), .ZN(new_n15993_));
  NAND2_X1   g13068(.A1(new_n15989_), .A2(new_n15993_), .ZN(new_n15994_));
  AOI21_X1   g13069(.A1(new_n15985_), .A2(new_n15976_), .B(new_n15994_), .ZN(new_n15995_));
  NOR3_X1    g13070(.A1(new_n14758_), .A2(pi0039), .A3(pi0161), .ZN(new_n15996_));
  OR2_X2     g13071(.A1(new_n15962_), .A2(new_n15437_), .Z(new_n15997_));
  NAND2_X1   g13072(.A1(new_n15684_), .A2(new_n15969_), .ZN(new_n15998_));
  NOR2_X1    g13073(.A1(new_n15998_), .A2(new_n3285_), .ZN(new_n15999_));
  NOR4_X1    g13074(.A1(new_n15683_), .A2(new_n4701_), .A3(pi0215), .A4(new_n15999_), .ZN(new_n16000_));
  NAND2_X1   g13075(.A1(new_n15434_), .A2(new_n16000_), .ZN(new_n16001_));
  AOI21_X1   g13076(.A1(new_n15997_), .A2(new_n15681_), .B(new_n16001_), .ZN(new_n16002_));
  AOI22_X1   g13077(.A1(new_n15653_), .A2(new_n15971_), .B1(new_n2614_), .B2(new_n15998_), .ZN(new_n16003_));
  NOR2_X1    g13078(.A1(new_n15981_), .A2(pi0758), .ZN(new_n16004_));
  OAI21_X1   g13079(.A1(new_n16003_), .A2(pi0223), .B(new_n16004_), .ZN(new_n16005_));
  NOR3_X1    g13080(.A1(new_n16005_), .A2(new_n16002_), .A3(new_n15996_), .ZN(new_n16006_));
  NOR2_X1    g13081(.A1(new_n14611_), .A2(pi0038), .ZN(new_n16008_));
  NAND4_X1   g13082(.A1(new_n15988_), .A2(new_n15987_), .A3(new_n3154_), .A4(new_n16008_), .ZN(new_n16009_));
  OAI21_X1   g13083(.A1(new_n16006_), .A2(new_n16009_), .B(new_n7832_), .ZN(new_n16010_));
  NOR2_X1    g13084(.A1(new_n15995_), .A2(new_n16010_), .ZN(new_n16011_));
  OAI21_X1   g13085(.A1(new_n7832_), .A2(pi0161), .B(new_n13184_), .ZN(new_n16012_));
  NOR4_X1    g13086(.A1(new_n15372_), .A2(new_n14611_), .A3(new_n2925_), .A4(new_n15986_), .ZN(new_n16013_));
  OAI21_X1   g13087(.A1(new_n2925_), .A2(pi0161), .B(pi0832), .ZN(new_n16014_));
  OAI22_X1   g13088(.A1(new_n16011_), .A2(new_n16012_), .B1(new_n16013_), .B2(new_n16014_), .ZN(po0318));
  NOR2_X1    g13089(.A1(new_n7325_), .A2(new_n2587_), .ZN(new_n16016_));
  NOR2_X1    g13090(.A1(new_n15473_), .A2(new_n16016_), .ZN(new_n16017_));
  OAI21_X1   g13091(.A1(new_n15475_), .A2(new_n7325_), .B(pi0761), .ZN(new_n16018_));
  NOR2_X1    g13092(.A1(new_n16017_), .A2(new_n16018_), .ZN(new_n16019_));
  NAND2_X1   g13093(.A1(new_n15400_), .A2(pi0162), .ZN(new_n16020_));
  NAND2_X1   g13094(.A1(new_n15515_), .A2(pi0162), .ZN(new_n16021_));
  NAND4_X1   g13095(.A1(new_n16020_), .A2(pi0039), .A3(new_n12116_), .A4(new_n16021_), .ZN(new_n16022_));
  OAI21_X1   g13096(.A1(new_n12852_), .A2(pi0162), .B(new_n3154_), .ZN(new_n16023_));
  NOR2_X1    g13097(.A1(new_n5473_), .A2(pi0761), .ZN(new_n16024_));
  NAND3_X1   g13098(.A1(new_n16023_), .A2(new_n12852_), .A3(new_n16024_), .ZN(new_n16025_));
  OAI22_X1   g13099(.A1(new_n16019_), .A2(new_n16022_), .B1(new_n15373_), .B2(new_n16025_), .ZN(new_n16026_));
  NAND2_X1   g13100(.A1(new_n13368_), .A2(new_n7325_), .ZN(new_n16027_));
  NOR4_X1    g13101(.A1(new_n15523_), .A2(pi0039), .A3(new_n12116_), .A4(new_n5473_), .ZN(new_n16028_));
  NOR2_X1    g13102(.A1(new_n16028_), .A2(new_n3172_), .ZN(new_n16029_));
  AOI22_X1   g13103(.A1(new_n16026_), .A2(new_n3172_), .B1(new_n16027_), .B2(new_n16029_), .ZN(new_n16030_));
  NOR3_X1    g13104(.A1(new_n15441_), .A2(new_n12116_), .A3(new_n15475_), .ZN(new_n16031_));
  NAND2_X1   g13105(.A1(new_n12894_), .A2(pi0761), .ZN(new_n16032_));
  NAND2_X1   g13106(.A1(new_n15475_), .A2(pi0947), .ZN(new_n16033_));
  AOI21_X1   g13107(.A1(new_n15489_), .A2(new_n16016_), .B(pi0761), .ZN(new_n16034_));
  NAND2_X1   g13108(.A1(new_n16033_), .A2(new_n16034_), .ZN(new_n16035_));
  NAND4_X1   g13109(.A1(new_n16035_), .A2(pi0039), .A3(new_n7325_), .A4(new_n16032_), .ZN(new_n16036_));
  AND2_X2    g13110(.A1(new_n16025_), .A2(new_n3172_), .Z(new_n16037_));
  OAI21_X1   g13111(.A1(new_n16031_), .A2(new_n16036_), .B(new_n16037_), .ZN(new_n16038_));
  NAND2_X1   g13112(.A1(new_n12899_), .A2(pi0162), .ZN(new_n16039_));
  NOR2_X1    g13113(.A1(new_n13368_), .A2(new_n16024_), .ZN(new_n16040_));
  NOR2_X1    g13114(.A1(new_n16040_), .A2(new_n3172_), .ZN(new_n16041_));
  AOI21_X1   g13115(.A1(new_n16039_), .A2(new_n16041_), .B(new_n11881_), .ZN(new_n16042_));
  AOI21_X1   g13116(.A1(new_n16038_), .A2(new_n16042_), .B(new_n7833_), .ZN(new_n16043_));
  OAI21_X1   g13117(.A1(new_n16030_), .A2(pi0738), .B(new_n16043_), .ZN(new_n16044_));
  AOI21_X1   g13118(.A1(new_n7833_), .A2(new_n7325_), .B(pi0832), .ZN(new_n16045_));
  AOI21_X1   g13119(.A1(new_n11881_), .A2(new_n15351_), .B(new_n16024_), .ZN(new_n16046_));
  MUX2_X1    g13120(.I0(new_n16046_), .I1(pi0162), .S(new_n2926_), .Z(new_n16047_));
  AOI22_X1   g13121(.A1(new_n16044_), .A2(new_n16045_), .B1(pi0832), .B2(new_n16047_), .ZN(po0319));
  INV_X1     g13122(.I(pi0777), .ZN(new_n16049_));
  NAND3_X1   g13123(.A1(new_n12792_), .A2(new_n8826_), .A3(new_n2587_), .ZN(new_n16050_));
  OAI21_X1   g13124(.A1(pi0163), .A2(new_n15475_), .B(new_n15368_), .ZN(new_n16051_));
  AOI22_X1   g13125(.A1(new_n16051_), .A2(new_n16050_), .B1(new_n16049_), .B2(new_n15510_), .ZN(new_n16052_));
  NAND2_X1   g13126(.A1(new_n15400_), .A2(pi0163), .ZN(new_n16053_));
  NAND2_X1   g13127(.A1(new_n15515_), .A2(pi0163), .ZN(new_n16054_));
  NAND4_X1   g13128(.A1(new_n16053_), .A2(pi0039), .A3(new_n16049_), .A4(new_n16054_), .ZN(new_n16055_));
  OAI21_X1   g13129(.A1(new_n12852_), .A2(pi0163), .B(new_n3154_), .ZN(new_n16056_));
  NOR2_X1    g13130(.A1(new_n5473_), .A2(pi0777), .ZN(new_n16057_));
  NAND3_X1   g13131(.A1(new_n16056_), .A2(new_n12852_), .A3(new_n16057_), .ZN(new_n16058_));
  OAI22_X1   g13132(.A1(new_n16055_), .A2(new_n16052_), .B1(new_n15373_), .B2(new_n16058_), .ZN(new_n16059_));
  NAND2_X1   g13133(.A1(new_n13368_), .A2(new_n8826_), .ZN(new_n16060_));
  NOR4_X1    g13134(.A1(new_n15523_), .A2(pi0039), .A3(new_n16049_), .A4(new_n5473_), .ZN(new_n16061_));
  NOR2_X1    g13135(.A1(new_n16061_), .A2(new_n3172_), .ZN(new_n16062_));
  AOI22_X1   g13136(.A1(new_n16059_), .A2(new_n3172_), .B1(new_n16060_), .B2(new_n16062_), .ZN(new_n16063_));
  AOI21_X1   g13137(.A1(pi0163), .A2(new_n2587_), .B(new_n15457_), .ZN(new_n16064_));
  AOI21_X1   g13138(.A1(new_n15440_), .A2(new_n8826_), .B(new_n16064_), .ZN(new_n16065_));
  AOI21_X1   g13139(.A1(new_n8826_), .A2(new_n15376_), .B(new_n15494_), .ZN(new_n16066_));
  NOR3_X1    g13140(.A1(new_n16065_), .A2(pi0777), .A3(new_n16066_), .ZN(new_n16067_));
  NOR2_X1    g13141(.A1(pi0039), .A2(pi0777), .ZN(new_n16068_));
  OAI21_X1   g13142(.A1(new_n12894_), .A2(pi0163), .B(new_n16068_), .ZN(new_n16069_));
  AND2_X2    g13143(.A1(new_n16058_), .A2(new_n3172_), .Z(new_n16070_));
  OAI21_X1   g13144(.A1(new_n16067_), .A2(new_n16069_), .B(new_n16070_), .ZN(new_n16071_));
  INV_X1     g13145(.I(pi0737), .ZN(new_n16072_));
  NAND2_X1   g13146(.A1(new_n12899_), .A2(pi0163), .ZN(new_n16073_));
  NOR2_X1    g13147(.A1(new_n13368_), .A2(new_n16057_), .ZN(new_n16074_));
  NOR2_X1    g13148(.A1(new_n16074_), .A2(new_n3172_), .ZN(new_n16075_));
  AOI21_X1   g13149(.A1(new_n16073_), .A2(new_n16075_), .B(new_n16072_), .ZN(new_n16076_));
  AOI21_X1   g13150(.A1(new_n16071_), .A2(new_n16076_), .B(new_n7833_), .ZN(new_n16077_));
  OAI21_X1   g13151(.A1(new_n16063_), .A2(pi0737), .B(new_n16077_), .ZN(new_n16078_));
  AOI21_X1   g13152(.A1(new_n7833_), .A2(new_n8826_), .B(pi0832), .ZN(new_n16079_));
  AOI21_X1   g13153(.A1(new_n16072_), .A2(new_n15351_), .B(new_n16057_), .ZN(new_n16080_));
  MUX2_X1    g13154(.I0(new_n16080_), .I1(pi0163), .S(new_n2926_), .Z(new_n16081_));
  AOI22_X1   g13155(.A1(new_n16078_), .A2(new_n16079_), .B1(pi0832), .B2(new_n16081_), .ZN(po0320));
  INV_X1     g13156(.I(new_n15779_), .ZN(new_n16083_));
  NOR2_X1    g13157(.A1(new_n12828_), .A2(pi0164), .ZN(new_n16084_));
  NOR4_X1    g13158(.A1(new_n16083_), .A2(pi0038), .A3(pi0752), .A4(new_n16084_), .ZN(new_n16085_));
  OAI21_X1   g13159(.A1(new_n15380_), .A2(new_n7058_), .B(new_n16085_), .ZN(new_n16086_));
  AOI21_X1   g13160(.A1(new_n15371_), .A2(pi0164), .B(new_n16086_), .ZN(new_n16087_));
  NOR2_X1    g13161(.A1(new_n15404_), .A2(new_n7058_), .ZN(new_n16088_));
  INV_X1     g13162(.I(pi0752), .ZN(new_n16089_));
  NOR2_X1    g13163(.A1(new_n16089_), .A2(pi0038), .ZN(new_n16091_));
  OAI21_X1   g13164(.A1(new_n15420_), .A2(new_n7058_), .B(new_n16091_), .ZN(new_n16092_));
  OAI21_X1   g13165(.A1(new_n16088_), .A2(new_n16092_), .B(pi0703), .ZN(new_n16093_));
  INV_X1     g13166(.I(pi0703), .ZN(new_n16094_));
  OAI21_X1   g13167(.A1(new_n15823_), .A2(new_n16089_), .B(new_n16094_), .ZN(new_n16095_));
  INV_X1     g13168(.I(new_n15428_), .ZN(new_n16096_));
  NAND4_X1   g13169(.A1(new_n15460_), .A2(new_n7058_), .A3(new_n16089_), .A4(new_n16096_), .ZN(new_n16097_));
  NOR2_X1    g13170(.A1(new_n15444_), .A2(new_n16097_), .ZN(new_n16098_));
  AOI21_X1   g13171(.A1(new_n16098_), .A2(new_n16095_), .B(new_n7833_), .ZN(new_n16099_));
  OAI21_X1   g13172(.A1(new_n16087_), .A2(new_n16093_), .B(new_n16099_), .ZN(new_n16100_));
  AOI21_X1   g13173(.A1(new_n7833_), .A2(new_n7058_), .B(pi0832), .ZN(new_n16101_));
  NAND2_X1   g13174(.A1(pi0703), .A2(pi0907), .ZN(new_n16102_));
  MUX2_X1    g13175(.I0(new_n16102_), .I1(pi0752), .S(pi0947), .Z(new_n16103_));
  MUX2_X1    g13176(.I0(new_n7058_), .I1(new_n16103_), .S(new_n2925_), .Z(new_n16104_));
  NOR2_X1    g13177(.A1(new_n16104_), .A2(new_n13184_), .ZN(new_n16105_));
  AOI21_X1   g13178(.A1(new_n16100_), .A2(new_n16101_), .B(new_n16105_), .ZN(po0321));
  INV_X1     g13179(.I(pi0165), .ZN(new_n16107_));
  NOR2_X1    g13180(.A1(new_n12828_), .A2(pi0165), .ZN(new_n16108_));
  NOR4_X1    g13181(.A1(new_n16083_), .A2(pi0038), .A3(pi0774), .A4(new_n16108_), .ZN(new_n16109_));
  OAI21_X1   g13182(.A1(new_n15380_), .A2(new_n16107_), .B(new_n16109_), .ZN(new_n16110_));
  AOI21_X1   g13183(.A1(new_n15371_), .A2(pi0165), .B(new_n16110_), .ZN(new_n16111_));
  NOR2_X1    g13184(.A1(new_n15404_), .A2(new_n16107_), .ZN(new_n16112_));
  NOR2_X1    g13185(.A1(new_n14348_), .A2(pi0038), .ZN(new_n16114_));
  OAI21_X1   g13186(.A1(new_n15420_), .A2(new_n16107_), .B(new_n16114_), .ZN(new_n16115_));
  OAI21_X1   g13187(.A1(new_n16112_), .A2(new_n16115_), .B(pi0687), .ZN(new_n16116_));
  OAI21_X1   g13188(.A1(new_n15823_), .A2(new_n14348_), .B(new_n14216_), .ZN(new_n16117_));
  NAND4_X1   g13189(.A1(new_n15460_), .A2(new_n16107_), .A3(new_n14348_), .A4(new_n16096_), .ZN(new_n16118_));
  NOR2_X1    g13190(.A1(new_n15444_), .A2(new_n16118_), .ZN(new_n16119_));
  AOI21_X1   g13191(.A1(new_n16119_), .A2(new_n16117_), .B(new_n7833_), .ZN(new_n16120_));
  OAI21_X1   g13192(.A1(new_n16111_), .A2(new_n16116_), .B(new_n16120_), .ZN(new_n16121_));
  AOI21_X1   g13193(.A1(new_n7833_), .A2(new_n16107_), .B(pi0832), .ZN(new_n16122_));
  NAND2_X1   g13194(.A1(pi0687), .A2(pi0907), .ZN(new_n16123_));
  MUX2_X1    g13195(.I0(new_n16123_), .I1(pi0774), .S(pi0947), .Z(new_n16124_));
  MUX2_X1    g13196(.I0(new_n16107_), .I1(new_n16124_), .S(new_n2925_), .Z(new_n16125_));
  NOR2_X1    g13197(.A1(new_n16125_), .A2(new_n13184_), .ZN(new_n16126_));
  AOI21_X1   g13198(.A1(new_n16121_), .A2(new_n16122_), .B(new_n16126_), .ZN(po0322));
  INV_X1     g13199(.I(pi0727), .ZN(new_n16128_));
  INV_X1     g13200(.I(pi0772), .ZN(new_n16129_));
  AOI21_X1   g13201(.A1(new_n15358_), .A2(pi0166), .B(new_n15631_), .ZN(new_n16130_));
  NOR2_X1    g13202(.A1(new_n16130_), .A2(new_n15361_), .ZN(new_n16131_));
  OAI21_X1   g13203(.A1(pi0166), .A2(new_n12709_), .B(new_n15432_), .ZN(new_n16132_));
  NAND2_X1   g13204(.A1(new_n15628_), .A2(new_n2587_), .ZN(new_n16133_));
  NOR2_X1    g13205(.A1(new_n12132_), .A2(pi0166), .ZN(new_n16134_));
  AOI21_X1   g13206(.A1(new_n5092_), .A2(new_n12132_), .B(new_n16134_), .ZN(new_n16135_));
  OAI21_X1   g13207(.A1(new_n16135_), .A2(new_n3285_), .B(new_n2566_), .ZN(new_n16136_));
  OAI21_X1   g13208(.A1(new_n16133_), .A2(new_n16132_), .B(new_n16136_), .ZN(new_n16137_));
  NOR2_X1    g13209(.A1(new_n16131_), .A2(new_n16137_), .ZN(new_n16138_));
  OAI21_X1   g13210(.A1(new_n16135_), .A2(new_n3155_), .B(new_n2604_), .ZN(new_n16139_));
  AOI21_X1   g13211(.A1(new_n2614_), .A2(new_n15452_), .B(new_n16139_), .ZN(new_n16140_));
  AOI21_X1   g13212(.A1(new_n15640_), .A2(new_n4549_), .B(new_n15372_), .ZN(new_n16141_));
  NOR3_X1    g13213(.A1(new_n15654_), .A2(new_n4549_), .A3(new_n15351_), .ZN(new_n16142_));
  NOR3_X1    g13214(.A1(new_n16142_), .A2(new_n2614_), .A3(new_n16141_), .ZN(new_n16143_));
  OAI21_X1   g13215(.A1(new_n15389_), .A2(new_n5092_), .B(new_n4549_), .ZN(new_n16144_));
  NAND2_X1   g13216(.A1(new_n2587_), .A2(new_n16129_), .ZN(new_n16145_));
  AOI21_X1   g13217(.A1(new_n15393_), .A2(new_n16144_), .B(new_n16145_), .ZN(new_n16146_));
  OAI21_X1   g13218(.A1(new_n16143_), .A2(new_n16140_), .B(new_n16146_), .ZN(new_n16147_));
  OAI21_X1   g13219(.A1(new_n16147_), .A2(new_n16138_), .B(pi0039), .ZN(new_n16148_));
  AOI21_X1   g13220(.A1(new_n16130_), .A2(new_n15664_), .B(new_n16136_), .ZN(new_n16149_));
  NAND2_X1   g13221(.A1(new_n16132_), .A2(pi0299), .ZN(new_n16150_));
  INV_X1     g13222(.I(new_n15391_), .ZN(new_n16151_));
  NOR2_X1    g13223(.A1(new_n15392_), .A2(pi0166), .ZN(new_n16152_));
  OAI21_X1   g13224(.A1(new_n16151_), .A2(new_n16152_), .B(new_n2587_), .ZN(new_n16153_));
  NAND2_X1   g13225(.A1(new_n15640_), .A2(new_n4549_), .ZN(new_n16154_));
  AOI21_X1   g13226(.A1(new_n15393_), .A2(new_n16144_), .B(new_n15655_), .ZN(new_n16155_));
  NAND4_X1   g13227(.A1(new_n16155_), .A2(new_n15643_), .A3(new_n16139_), .A4(new_n16154_), .ZN(new_n16156_));
  OAI22_X1   g13228(.A1(new_n16156_), .A2(new_n16153_), .B1(new_n16149_), .B2(new_n16150_), .ZN(new_n16157_));
  NAND3_X1   g13229(.A1(new_n16157_), .A2(new_n16129_), .A3(new_n16148_), .ZN(new_n16158_));
  NOR2_X1    g13230(.A1(new_n16129_), .A2(new_n5473_), .ZN(new_n16159_));
  INV_X1     g13231(.I(new_n16159_), .ZN(new_n16160_));
  AOI21_X1   g13232(.A1(new_n12697_), .A2(new_n4549_), .B(new_n16160_), .ZN(new_n16161_));
  NOR3_X1    g13233(.A1(new_n12852_), .A2(new_n4549_), .A3(new_n16159_), .ZN(new_n16162_));
  NOR3_X1    g13234(.A1(new_n16161_), .A2(new_n16162_), .A3(pi0039), .ZN(new_n16163_));
  AOI21_X1   g13235(.A1(new_n16163_), .A2(new_n15373_), .B(pi0038), .ZN(new_n16166_));
  NAND2_X1   g13236(.A1(new_n16158_), .A2(new_n16166_), .ZN(new_n16167_));
  NAND2_X1   g13237(.A1(new_n12899_), .A2(new_n4549_), .ZN(new_n16168_));
  AOI21_X1   g13238(.A1(new_n12828_), .A2(new_n16160_), .B(new_n3172_), .ZN(new_n16169_));
  AOI21_X1   g13239(.A1(new_n16168_), .A2(new_n16169_), .B(pi0727), .ZN(new_n16170_));
  NOR2_X1    g13240(.A1(new_n15652_), .A2(new_n2614_), .ZN(new_n16171_));
  AOI21_X1   g13241(.A1(new_n5473_), .A2(new_n12132_), .B(new_n16134_), .ZN(new_n16172_));
  AOI22_X1   g13242(.A1(new_n16171_), .A2(new_n16154_), .B1(new_n2614_), .B2(new_n16172_), .ZN(new_n16173_));
  NAND2_X1   g13243(.A1(new_n2604_), .A2(new_n2587_), .ZN(new_n16174_));
  NOR2_X1    g13244(.A1(new_n16130_), .A2(new_n15437_), .ZN(new_n16175_));
  NOR2_X1    g13245(.A1(new_n16175_), .A2(new_n15357_), .ZN(new_n16176_));
  INV_X1     g13246(.I(new_n15434_), .ZN(new_n16177_));
  NOR2_X1    g13247(.A1(new_n4549_), .A2(pi0215), .ZN(new_n16178_));
  OAI21_X1   g13248(.A1(new_n16172_), .A2(new_n3285_), .B(new_n16178_), .ZN(new_n16179_));
  OR3_X2     g13249(.A1(new_n16177_), .A2(new_n15683_), .A3(new_n16179_), .Z(new_n16180_));
  OAI22_X1   g13250(.A1(new_n16173_), .A2(new_n16174_), .B1(new_n16176_), .B2(new_n16180_), .ZN(new_n16181_));
  NOR2_X1    g13251(.A1(pi0039), .A2(pi0166), .ZN(new_n16182_));
  AOI21_X1   g13252(.A1(new_n12894_), .A2(new_n16182_), .B(pi0772), .ZN(new_n16183_));
  NAND2_X1   g13253(.A1(new_n16163_), .A2(new_n3172_), .ZN(new_n16184_));
  AOI21_X1   g13254(.A1(new_n16181_), .A2(new_n16183_), .B(new_n16184_), .ZN(new_n16185_));
  OAI21_X1   g13255(.A1(new_n16185_), .A2(new_n16170_), .B(new_n7832_), .ZN(new_n16186_));
  AOI21_X1   g13256(.A1(new_n16167_), .A2(new_n16128_), .B(new_n16186_), .ZN(new_n16187_));
  OAI21_X1   g13257(.A1(new_n7832_), .A2(pi0166), .B(new_n13184_), .ZN(new_n16188_));
  NOR4_X1    g13258(.A1(new_n15372_), .A2(new_n16128_), .A3(new_n2925_), .A4(new_n16159_), .ZN(new_n16189_));
  OAI21_X1   g13259(.A1(new_n2925_), .A2(pi0166), .B(pi0832), .ZN(new_n16190_));
  OAI22_X1   g13260(.A1(new_n16187_), .A2(new_n16188_), .B1(new_n16189_), .B2(new_n16190_), .ZN(po0323));
  NAND2_X1   g13261(.A1(pi0705), .A2(pi0907), .ZN(new_n16192_));
  MUX2_X1    g13262(.I0(new_n16192_), .I1(pi0768), .S(pi0947), .Z(new_n16193_));
  MUX2_X1    g13263(.I0(new_n7334_), .I1(new_n16193_), .S(new_n2925_), .Z(new_n16194_));
  OAI21_X1   g13264(.A1(new_n15380_), .A2(new_n7334_), .B(new_n3172_), .ZN(new_n16196_));
  AOI21_X1   g13265(.A1(new_n15371_), .A2(pi0167), .B(new_n16196_), .ZN(new_n16197_));
  INV_X1     g13266(.I(pi0705), .ZN(new_n16198_));
  NAND2_X1   g13267(.A1(new_n15403_), .A2(pi0167), .ZN(new_n16199_));
  NOR2_X1    g13268(.A1(new_n15420_), .A2(new_n7334_), .ZN(new_n16200_));
  INV_X1     g13269(.I(pi0768), .ZN(new_n16201_));
  NAND2_X1   g13270(.A1(new_n3172_), .A2(new_n16201_), .ZN(new_n16203_));
  NOR2_X1    g13271(.A1(new_n16200_), .A2(new_n16203_), .ZN(new_n16204_));
  AOI21_X1   g13272(.A1(new_n16199_), .A2(new_n16204_), .B(new_n16198_), .ZN(new_n16205_));
  NOR3_X1    g13273(.A1(new_n16197_), .A2(pi0768), .A3(new_n16205_), .ZN(new_n16206_));
  OAI21_X1   g13274(.A1(new_n15443_), .A2(pi0167), .B(new_n3172_), .ZN(new_n16207_));
  NOR2_X1    g13275(.A1(new_n15459_), .A2(new_n7334_), .ZN(new_n16208_));
  NAND2_X1   g13276(.A1(new_n16207_), .A2(new_n16208_), .ZN(new_n16209_));
  NOR2_X1    g13277(.A1(new_n15144_), .A2(new_n3172_), .ZN(new_n16210_));
  NAND3_X1   g13278(.A1(new_n16210_), .A2(new_n16201_), .A3(new_n12901_), .ZN(new_n16211_));
  OAI21_X1   g13279(.A1(new_n16211_), .A2(pi0167), .B(new_n16198_), .ZN(new_n16212_));
  OAI21_X1   g13280(.A1(pi0167), .A2(new_n12898_), .B(new_n15447_), .ZN(new_n16213_));
  NAND2_X1   g13281(.A1(new_n16213_), .A2(new_n16201_), .ZN(new_n16214_));
  AOI21_X1   g13282(.A1(pi0167), .A2(new_n13184_), .B(new_n7832_), .ZN(new_n16215_));
  NAND4_X1   g13283(.A1(new_n16209_), .A2(new_n16212_), .A3(new_n16214_), .A4(new_n16215_), .ZN(new_n16216_));
  OAI22_X1   g13284(.A1(new_n16206_), .A2(new_n16216_), .B1(new_n13184_), .B2(new_n16194_), .ZN(po0324));
  OAI21_X1   g13285(.A1(new_n2925_), .A2(new_n4413_), .B(pi0832), .ZN(new_n16218_));
  AOI21_X1   g13286(.A1(pi0763), .A2(pi0947), .B(new_n2926_), .ZN(new_n16219_));
  INV_X1     g13287(.I(new_n16219_), .ZN(new_n16220_));
  NAND4_X1   g13288(.A1(new_n16220_), .A2(pi0699), .A3(new_n16218_), .A4(new_n15351_), .ZN(new_n16221_));
  INV_X1     g13289(.I(pi0763), .ZN(new_n16222_));
  NOR4_X1    g13290(.A1(new_n15523_), .A2(pi0039), .A3(new_n16222_), .A4(pi0947), .ZN(new_n16223_));
  NOR2_X1    g13291(.A1(new_n16223_), .A2(new_n3172_), .ZN(new_n16224_));
  OAI21_X1   g13292(.A1(pi0168), .A2(new_n12828_), .B(new_n16224_), .ZN(new_n16225_));
  NAND2_X1   g13293(.A1(new_n12855_), .A2(pi0168), .ZN(new_n16226_));
  NAND2_X1   g13294(.A1(new_n15432_), .A2(new_n16226_), .ZN(new_n16227_));
  NOR2_X1    g13295(.A1(new_n15582_), .A2(new_n4413_), .ZN(new_n16228_));
  OAI21_X1   g13296(.A1(new_n15356_), .A2(new_n16228_), .B(new_n3285_), .ZN(new_n16229_));
  OAI21_X1   g13297(.A1(pi0168), .A2(new_n12132_), .B(new_n15453_), .ZN(new_n16230_));
  AOI21_X1   g13298(.A1(new_n16230_), .A2(new_n15716_), .B(pi0215), .ZN(new_n16231_));
  OAI21_X1   g13299(.A1(new_n16229_), .A2(new_n16231_), .B(new_n16227_), .ZN(new_n16232_));
  NOR2_X1    g13300(.A1(new_n15409_), .A2(new_n4413_), .ZN(new_n16233_));
  AOI22_X1   g13301(.A1(new_n15396_), .A2(new_n16233_), .B1(pi0299), .B2(new_n16232_), .ZN(new_n16234_));
  INV_X1     g13302(.I(new_n16229_), .ZN(new_n16235_));
  AOI21_X1   g13303(.A1(new_n4413_), .A2(new_n12133_), .B(new_n15722_), .ZN(new_n16236_));
  OAI21_X1   g13304(.A1(new_n15359_), .A2(new_n16236_), .B(new_n16235_), .ZN(new_n16237_));
  NAND2_X1   g13305(.A1(new_n16227_), .A2(new_n15410_), .ZN(new_n16238_));
  NAND2_X1   g13306(.A1(new_n16238_), .A2(new_n15726_), .ZN(new_n16239_));
  AOI21_X1   g13307(.A1(new_n16237_), .A2(new_n2566_), .B(new_n16239_), .ZN(new_n16240_));
  NOR2_X1    g13308(.A1(new_n12792_), .A2(pi0168), .ZN(new_n16241_));
  NOR2_X1    g13309(.A1(pi0039), .A2(pi0763), .ZN(new_n16242_));
  OAI21_X1   g13310(.A1(new_n15729_), .A2(new_n16241_), .B(new_n16242_), .ZN(new_n16243_));
  NOR3_X1    g13311(.A1(new_n16234_), .A2(new_n16240_), .A3(new_n16243_), .ZN(new_n16244_));
  NOR2_X1    g13312(.A1(new_n15734_), .A2(pi0763), .ZN(new_n16245_));
  OAI22_X1   g13313(.A1(new_n16245_), .A2(new_n15448_), .B1(pi0168), .B2(new_n12852_), .ZN(new_n16246_));
  NOR2_X1    g13314(.A1(new_n16246_), .A2(new_n15373_), .ZN(new_n16247_));
  OAI21_X1   g13315(.A1(new_n16244_), .A2(new_n16247_), .B(new_n3172_), .ZN(new_n16248_));
  NAND2_X1   g13316(.A1(new_n4413_), .A2(new_n16222_), .ZN(new_n16249_));
  OAI21_X1   g13317(.A1(new_n12894_), .A2(new_n16249_), .B(pi0039), .ZN(new_n16250_));
  NOR3_X1    g13318(.A1(new_n15434_), .A2(pi0299), .A3(new_n16226_), .ZN(new_n16251_));
  NAND2_X1   g13319(.A1(new_n16230_), .A2(new_n16222_), .ZN(new_n16252_));
  NOR4_X1    g13320(.A1(new_n15578_), .A2(new_n16229_), .A3(new_n16251_), .A4(new_n16252_), .ZN(new_n16253_));
  NOR3_X1    g13321(.A1(new_n16253_), .A2(new_n15494_), .A3(new_n16241_), .ZN(new_n16254_));
  INV_X1     g13322(.I(pi0699), .ZN(new_n16255_));
  NAND2_X1   g13323(.A1(new_n5156_), .A2(new_n16219_), .ZN(new_n16256_));
  NAND4_X1   g13324(.A1(new_n12898_), .A2(new_n3172_), .A3(new_n4413_), .A4(new_n16256_), .ZN(new_n16257_));
  NAND4_X1   g13325(.A1(new_n16246_), .A2(new_n3172_), .A3(new_n16255_), .A4(new_n16257_), .ZN(new_n16258_));
  AOI21_X1   g13326(.A1(new_n16254_), .A2(new_n16250_), .B(new_n16258_), .ZN(new_n16259_));
  OAI21_X1   g13327(.A1(new_n16259_), .A2(new_n15500_), .B(pi0699), .ZN(new_n16260_));
  AOI21_X1   g13328(.A1(new_n16248_), .A2(new_n16225_), .B(new_n16260_), .ZN(new_n16261_));
  NAND2_X1   g13329(.A1(pi0057), .A2(pi0168), .ZN(new_n16262_));
  AOI21_X1   g13330(.A1(new_n16262_), .A2(new_n13184_), .B(pi0057), .ZN(new_n16263_));
  OAI21_X1   g13331(.A1(new_n15499_), .A2(pi0168), .B(new_n16263_), .ZN(new_n16264_));
  OAI21_X1   g13332(.A1(new_n16261_), .A2(new_n16264_), .B(new_n16221_), .ZN(po0325));
  OAI21_X1   g13333(.A1(new_n2925_), .A2(new_n4272_), .B(pi0832), .ZN(new_n16266_));
  AOI21_X1   g13334(.A1(pi0746), .A2(pi0947), .B(new_n2926_), .ZN(new_n16267_));
  INV_X1     g13335(.I(new_n16267_), .ZN(new_n16268_));
  NAND4_X1   g13336(.A1(new_n16268_), .A2(pi0729), .A3(new_n16266_), .A4(new_n15351_), .ZN(new_n16269_));
  INV_X1     g13337(.I(pi0746), .ZN(new_n16270_));
  NOR4_X1    g13338(.A1(new_n15523_), .A2(pi0039), .A3(new_n16270_), .A4(pi0947), .ZN(new_n16271_));
  NOR2_X1    g13339(.A1(new_n16271_), .A2(new_n3172_), .ZN(new_n16272_));
  OAI21_X1   g13340(.A1(pi0169), .A2(new_n12828_), .B(new_n16272_), .ZN(new_n16273_));
  NAND2_X1   g13341(.A1(new_n12855_), .A2(pi0169), .ZN(new_n16274_));
  NAND2_X1   g13342(.A1(new_n15432_), .A2(new_n16274_), .ZN(new_n16275_));
  NOR2_X1    g13343(.A1(new_n15582_), .A2(new_n4272_), .ZN(new_n16276_));
  OAI21_X1   g13344(.A1(new_n15356_), .A2(new_n16276_), .B(new_n3285_), .ZN(new_n16277_));
  OAI21_X1   g13345(.A1(pi0169), .A2(new_n12132_), .B(new_n15453_), .ZN(new_n16278_));
  AOI21_X1   g13346(.A1(new_n16278_), .A2(new_n15716_), .B(pi0215), .ZN(new_n16279_));
  OAI21_X1   g13347(.A1(new_n16277_), .A2(new_n16279_), .B(new_n16275_), .ZN(new_n16280_));
  NOR2_X1    g13348(.A1(new_n15409_), .A2(new_n4272_), .ZN(new_n16281_));
  AOI22_X1   g13349(.A1(new_n15396_), .A2(new_n16281_), .B1(pi0299), .B2(new_n16280_), .ZN(new_n16282_));
  INV_X1     g13350(.I(new_n16277_), .ZN(new_n16283_));
  AOI21_X1   g13351(.A1(new_n4272_), .A2(new_n12133_), .B(new_n15722_), .ZN(new_n16284_));
  OAI21_X1   g13352(.A1(new_n15359_), .A2(new_n16284_), .B(new_n16283_), .ZN(new_n16285_));
  NAND2_X1   g13353(.A1(new_n16275_), .A2(new_n15410_), .ZN(new_n16286_));
  NAND2_X1   g13354(.A1(new_n16286_), .A2(new_n15726_), .ZN(new_n16287_));
  AOI21_X1   g13355(.A1(new_n16285_), .A2(new_n2566_), .B(new_n16287_), .ZN(new_n16288_));
  NOR2_X1    g13356(.A1(new_n12792_), .A2(pi0169), .ZN(new_n16289_));
  NOR2_X1    g13357(.A1(pi0039), .A2(pi0746), .ZN(new_n16290_));
  OAI21_X1   g13358(.A1(new_n15729_), .A2(new_n16289_), .B(new_n16290_), .ZN(new_n16291_));
  NOR3_X1    g13359(.A1(new_n16282_), .A2(new_n16288_), .A3(new_n16291_), .ZN(new_n16292_));
  NOR2_X1    g13360(.A1(new_n15734_), .A2(pi0746), .ZN(new_n16293_));
  OAI22_X1   g13361(.A1(new_n16293_), .A2(new_n15448_), .B1(pi0169), .B2(new_n12852_), .ZN(new_n16294_));
  NOR2_X1    g13362(.A1(new_n16294_), .A2(new_n15373_), .ZN(new_n16295_));
  OAI21_X1   g13363(.A1(new_n16292_), .A2(new_n16295_), .B(new_n3172_), .ZN(new_n16296_));
  NAND2_X1   g13364(.A1(new_n4272_), .A2(new_n16270_), .ZN(new_n16297_));
  OAI21_X1   g13365(.A1(new_n12894_), .A2(new_n16297_), .B(pi0039), .ZN(new_n16298_));
  NOR3_X1    g13366(.A1(new_n15434_), .A2(pi0299), .A3(new_n16274_), .ZN(new_n16299_));
  NAND2_X1   g13367(.A1(new_n16278_), .A2(new_n16270_), .ZN(new_n16300_));
  NOR4_X1    g13368(.A1(new_n15578_), .A2(new_n16277_), .A3(new_n16299_), .A4(new_n16300_), .ZN(new_n16301_));
  NOR3_X1    g13369(.A1(new_n16301_), .A2(new_n15494_), .A3(new_n16289_), .ZN(new_n16302_));
  INV_X1     g13370(.I(pi0729), .ZN(new_n16303_));
  NAND2_X1   g13371(.A1(new_n5156_), .A2(new_n16267_), .ZN(new_n16304_));
  NAND4_X1   g13372(.A1(new_n12898_), .A2(new_n3172_), .A3(new_n4272_), .A4(new_n16304_), .ZN(new_n16305_));
  NAND4_X1   g13373(.A1(new_n16294_), .A2(new_n3172_), .A3(new_n16303_), .A4(new_n16305_), .ZN(new_n16306_));
  AOI21_X1   g13374(.A1(new_n16302_), .A2(new_n16298_), .B(new_n16306_), .ZN(new_n16307_));
  OAI21_X1   g13375(.A1(new_n16307_), .A2(new_n15500_), .B(pi0729), .ZN(new_n16308_));
  AOI21_X1   g13376(.A1(new_n16296_), .A2(new_n16273_), .B(new_n16308_), .ZN(new_n16309_));
  NAND2_X1   g13377(.A1(pi0057), .A2(pi0169), .ZN(new_n16310_));
  AOI21_X1   g13378(.A1(new_n16310_), .A2(new_n13184_), .B(pi0057), .ZN(new_n16311_));
  OAI21_X1   g13379(.A1(new_n15499_), .A2(pi0169), .B(new_n16311_), .ZN(new_n16312_));
  OAI21_X1   g13380(.A1(new_n16309_), .A2(new_n16312_), .B(new_n16269_), .ZN(po0326));
  OAI21_X1   g13381(.A1(new_n2925_), .A2(new_n3984_), .B(pi0832), .ZN(new_n16314_));
  INV_X1     g13382(.I(pi0748), .ZN(new_n16315_));
  OAI21_X1   g13383(.A1(new_n16315_), .A2(new_n5473_), .B(new_n2925_), .ZN(new_n16316_));
  NAND4_X1   g13384(.A1(new_n16316_), .A2(pi0730), .A3(new_n16314_), .A4(new_n15351_), .ZN(new_n16317_));
  INV_X1     g13385(.I(pi0730), .ZN(new_n16318_));
  NAND3_X1   g13386(.A1(new_n15823_), .A2(new_n3984_), .A3(new_n16315_), .ZN(new_n16319_));
  OAI21_X1   g13387(.A1(new_n12792_), .A2(pi0170), .B(new_n2587_), .ZN(new_n16320_));
  NAND2_X1   g13388(.A1(new_n15450_), .A2(new_n16320_), .ZN(new_n16321_));
  NAND4_X1   g13389(.A1(new_n16177_), .A2(pi0170), .A3(new_n2587_), .A4(new_n12855_), .ZN(new_n16322_));
  OAI21_X1   g13390(.A1(pi0170), .A2(new_n12132_), .B(new_n15453_), .ZN(new_n16323_));
  NOR2_X1    g13391(.A1(new_n15582_), .A2(new_n3984_), .ZN(new_n16324_));
  OAI21_X1   g13392(.A1(new_n15356_), .A2(new_n16324_), .B(new_n3285_), .ZN(new_n16325_));
  INV_X1     g13393(.I(new_n16325_), .ZN(new_n16326_));
  NAND4_X1   g13394(.A1(new_n16322_), .A2(new_n15438_), .A3(new_n16323_), .A4(new_n16326_), .ZN(new_n16327_));
  AOI21_X1   g13395(.A1(new_n16327_), .A2(new_n16321_), .B(new_n3154_), .ZN(new_n16328_));
  NOR2_X1    g13396(.A1(new_n12852_), .A2(pi0170), .ZN(new_n16329_));
  NOR2_X1    g13397(.A1(new_n15449_), .A2(new_n16329_), .ZN(new_n16330_));
  OAI21_X1   g13398(.A1(new_n16328_), .A2(new_n16330_), .B(new_n3172_), .ZN(new_n16331_));
  NAND2_X1   g13399(.A1(new_n12899_), .A2(new_n3984_), .ZN(new_n16332_));
  NOR2_X1    g13400(.A1(new_n15499_), .A2(pi0748), .ZN(new_n16333_));
  NAND4_X1   g13401(.A1(new_n16331_), .A2(new_n15447_), .A3(new_n16332_), .A4(new_n16333_), .ZN(new_n16334_));
  AOI21_X1   g13402(.A1(new_n16318_), .A2(new_n16319_), .B(new_n16334_), .ZN(new_n16335_));
  NAND2_X1   g13403(.A1(new_n15377_), .A2(new_n16320_), .ZN(new_n16336_));
  OAI21_X1   g13404(.A1(pi0170), .A2(new_n12132_), .B(new_n15599_), .ZN(new_n16337_));
  NAND2_X1   g13405(.A1(new_n15360_), .A2(new_n16337_), .ZN(new_n16338_));
  AOI21_X1   g13406(.A1(new_n16338_), .A2(new_n16326_), .B(pi0215), .ZN(new_n16339_));
  AOI21_X1   g13407(.A1(pi0170), .A2(new_n12855_), .B(new_n15433_), .ZN(new_n16340_));
  OAI21_X1   g13408(.A1(new_n16340_), .A2(new_n15627_), .B(new_n15608_), .ZN(new_n16341_));
  OAI21_X1   g13409(.A1(new_n16339_), .A2(new_n16341_), .B(pi0299), .ZN(new_n16342_));
  AOI21_X1   g13410(.A1(new_n16342_), .A2(new_n16336_), .B(new_n3154_), .ZN(new_n16343_));
  NOR3_X1    g13411(.A1(new_n15373_), .A2(new_n16329_), .A3(pi0039), .ZN(new_n16344_));
  OAI21_X1   g13412(.A1(new_n16343_), .A2(new_n16344_), .B(new_n3172_), .ZN(new_n16345_));
  AOI21_X1   g13413(.A1(new_n16323_), .A2(new_n15716_), .B(pi0215), .ZN(new_n16346_));
  NOR2_X1    g13414(.A1(new_n16325_), .A2(new_n16346_), .ZN(new_n16347_));
  OAI21_X1   g13415(.A1(new_n16347_), .A2(new_n16340_), .B(pi0299), .ZN(new_n16348_));
  OAI21_X1   g13416(.A1(new_n3984_), .A2(new_n15409_), .B(new_n15395_), .ZN(new_n16349_));
  AOI21_X1   g13417(.A1(new_n16349_), .A2(new_n16348_), .B(pi0039), .ZN(new_n16350_));
  NAND2_X1   g13418(.A1(new_n15407_), .A2(new_n3154_), .ZN(new_n16351_));
  OAI21_X1   g13419(.A1(new_n16351_), .A2(new_n16329_), .B(new_n3172_), .ZN(new_n16352_));
  INV_X1     g13420(.I(new_n15800_), .ZN(new_n16353_));
  NOR2_X1    g13421(.A1(new_n12828_), .A2(pi0170), .ZN(new_n16354_));
  NOR4_X1    g13422(.A1(new_n16353_), .A2(pi0730), .A3(pi0748), .A4(new_n16354_), .ZN(new_n16355_));
  OAI21_X1   g13423(.A1(new_n16350_), .A2(new_n16352_), .B(new_n16355_), .ZN(new_n16356_));
  OAI21_X1   g13424(.A1(new_n16083_), .A2(new_n16354_), .B(new_n16315_), .ZN(new_n16357_));
  NAND3_X1   g13425(.A1(new_n16345_), .A2(new_n16356_), .A3(new_n16357_), .ZN(new_n16358_));
  NOR2_X1    g13426(.A1(new_n5055_), .A2(new_n3984_), .ZN(new_n16359_));
  OAI21_X1   g13427(.A1(new_n16359_), .A2(pi0832), .B(new_n5055_), .ZN(new_n16360_));
  AOI21_X1   g13428(.A1(new_n15500_), .A2(new_n3984_), .B(new_n16360_), .ZN(new_n16361_));
  OAI21_X1   g13429(.A1(new_n16358_), .A2(new_n16335_), .B(new_n16361_), .ZN(new_n16362_));
  NAND2_X1   g13430(.A1(new_n16362_), .A2(new_n16317_), .ZN(po0327));
  OAI21_X1   g13431(.A1(new_n2925_), .A2(new_n3842_), .B(pi0832), .ZN(new_n16364_));
  AOI21_X1   g13432(.A1(pi0764), .A2(pi0947), .B(new_n2926_), .ZN(new_n16365_));
  INV_X1     g13433(.I(new_n16365_), .ZN(new_n16366_));
  NAND4_X1   g13434(.A1(new_n16366_), .A2(pi0691), .A3(new_n16364_), .A4(new_n15351_), .ZN(new_n16367_));
  INV_X1     g13435(.I(pi0764), .ZN(new_n16368_));
  NOR4_X1    g13436(.A1(new_n15523_), .A2(pi0039), .A3(new_n16368_), .A4(pi0947), .ZN(new_n16369_));
  NOR2_X1    g13437(.A1(new_n16369_), .A2(new_n3172_), .ZN(new_n16370_));
  OAI21_X1   g13438(.A1(pi0171), .A2(new_n12828_), .B(new_n16370_), .ZN(new_n16371_));
  NAND2_X1   g13439(.A1(new_n12855_), .A2(pi0171), .ZN(new_n16372_));
  NAND2_X1   g13440(.A1(new_n15432_), .A2(new_n16372_), .ZN(new_n16373_));
  NOR2_X1    g13441(.A1(new_n15582_), .A2(new_n3842_), .ZN(new_n16374_));
  OAI21_X1   g13442(.A1(new_n15356_), .A2(new_n16374_), .B(new_n3285_), .ZN(new_n16375_));
  OAI21_X1   g13443(.A1(pi0171), .A2(new_n12132_), .B(new_n15453_), .ZN(new_n16376_));
  AOI21_X1   g13444(.A1(new_n16376_), .A2(new_n15716_), .B(pi0215), .ZN(new_n16377_));
  OAI21_X1   g13445(.A1(new_n16375_), .A2(new_n16377_), .B(new_n16373_), .ZN(new_n16378_));
  NOR2_X1    g13446(.A1(new_n15409_), .A2(new_n3842_), .ZN(new_n16379_));
  AOI22_X1   g13447(.A1(new_n15396_), .A2(new_n16379_), .B1(pi0299), .B2(new_n16378_), .ZN(new_n16380_));
  INV_X1     g13448(.I(new_n16375_), .ZN(new_n16381_));
  AOI21_X1   g13449(.A1(new_n3842_), .A2(new_n12133_), .B(new_n15722_), .ZN(new_n16382_));
  OAI21_X1   g13450(.A1(new_n15359_), .A2(new_n16382_), .B(new_n16381_), .ZN(new_n16383_));
  NAND2_X1   g13451(.A1(new_n16373_), .A2(new_n15410_), .ZN(new_n16384_));
  NAND2_X1   g13452(.A1(new_n16384_), .A2(new_n15726_), .ZN(new_n16385_));
  AOI21_X1   g13453(.A1(new_n16383_), .A2(new_n2566_), .B(new_n16385_), .ZN(new_n16386_));
  NOR2_X1    g13454(.A1(new_n12792_), .A2(pi0171), .ZN(new_n16387_));
  NOR2_X1    g13455(.A1(pi0039), .A2(pi0764), .ZN(new_n16388_));
  OAI21_X1   g13456(.A1(new_n15729_), .A2(new_n16387_), .B(new_n16388_), .ZN(new_n16389_));
  NOR3_X1    g13457(.A1(new_n16380_), .A2(new_n16386_), .A3(new_n16389_), .ZN(new_n16390_));
  NOR2_X1    g13458(.A1(new_n15734_), .A2(pi0764), .ZN(new_n16391_));
  OAI22_X1   g13459(.A1(new_n16391_), .A2(new_n15448_), .B1(pi0171), .B2(new_n12852_), .ZN(new_n16392_));
  NOR2_X1    g13460(.A1(new_n16392_), .A2(new_n15373_), .ZN(new_n16393_));
  OAI21_X1   g13461(.A1(new_n16390_), .A2(new_n16393_), .B(new_n3172_), .ZN(new_n16394_));
  NAND2_X1   g13462(.A1(new_n3842_), .A2(new_n16368_), .ZN(new_n16395_));
  OAI21_X1   g13463(.A1(new_n12894_), .A2(new_n16395_), .B(pi0039), .ZN(new_n16396_));
  NOR3_X1    g13464(.A1(new_n15434_), .A2(pi0299), .A3(new_n16372_), .ZN(new_n16397_));
  NAND2_X1   g13465(.A1(new_n16376_), .A2(new_n16368_), .ZN(new_n16398_));
  NOR4_X1    g13466(.A1(new_n15578_), .A2(new_n16375_), .A3(new_n16397_), .A4(new_n16398_), .ZN(new_n16399_));
  NOR3_X1    g13467(.A1(new_n16399_), .A2(new_n15494_), .A3(new_n16387_), .ZN(new_n16400_));
  INV_X1     g13468(.I(pi0691), .ZN(new_n16401_));
  NAND2_X1   g13469(.A1(new_n5156_), .A2(new_n16365_), .ZN(new_n16402_));
  NAND4_X1   g13470(.A1(new_n12898_), .A2(new_n3172_), .A3(new_n3842_), .A4(new_n16402_), .ZN(new_n16403_));
  NAND4_X1   g13471(.A1(new_n16392_), .A2(new_n3172_), .A3(new_n16401_), .A4(new_n16403_), .ZN(new_n16404_));
  AOI21_X1   g13472(.A1(new_n16400_), .A2(new_n16396_), .B(new_n16404_), .ZN(new_n16405_));
  OAI21_X1   g13473(.A1(new_n16405_), .A2(new_n15500_), .B(pi0691), .ZN(new_n16406_));
  AOI21_X1   g13474(.A1(new_n16394_), .A2(new_n16371_), .B(new_n16406_), .ZN(new_n16407_));
  NAND2_X1   g13475(.A1(pi0057), .A2(pi0171), .ZN(new_n16408_));
  AOI21_X1   g13476(.A1(new_n16408_), .A2(new_n13184_), .B(pi0057), .ZN(new_n16409_));
  OAI21_X1   g13477(.A1(new_n15499_), .A2(pi0171), .B(new_n16409_), .ZN(new_n16410_));
  OAI21_X1   g13478(.A1(new_n16407_), .A2(new_n16410_), .B(new_n16367_), .ZN(po0328));
  NAND2_X1   g13479(.A1(pi0739), .A2(pi0947), .ZN(new_n16412_));
  NAND4_X1   g13480(.A1(new_n2926_), .A2(pi0690), .A3(new_n15351_), .A4(new_n16412_), .ZN(new_n16413_));
  NAND4_X1   g13481(.A1(new_n16413_), .A2(new_n3707_), .A3(new_n13184_), .A4(new_n2925_), .ZN(new_n16414_));
  INV_X1     g13482(.I(pi0739), .ZN(new_n16415_));
  NOR4_X1    g13483(.A1(new_n15523_), .A2(pi0039), .A3(new_n16415_), .A4(pi0947), .ZN(new_n16416_));
  NOR2_X1    g13484(.A1(new_n16416_), .A2(new_n3172_), .ZN(new_n16417_));
  OAI21_X1   g13485(.A1(pi0172), .A2(new_n12828_), .B(new_n16417_), .ZN(new_n16418_));
  NAND2_X1   g13486(.A1(new_n12855_), .A2(pi0172), .ZN(new_n16419_));
  NAND2_X1   g13487(.A1(new_n15432_), .A2(new_n16419_), .ZN(new_n16420_));
  NOR2_X1    g13488(.A1(new_n15582_), .A2(new_n3707_), .ZN(new_n16421_));
  OAI21_X1   g13489(.A1(new_n15356_), .A2(new_n16421_), .B(new_n3285_), .ZN(new_n16422_));
  OAI21_X1   g13490(.A1(pi0172), .A2(new_n12132_), .B(new_n15453_), .ZN(new_n16423_));
  AOI21_X1   g13491(.A1(new_n16423_), .A2(new_n15716_), .B(pi0215), .ZN(new_n16424_));
  OAI21_X1   g13492(.A1(new_n16422_), .A2(new_n16424_), .B(new_n16420_), .ZN(new_n16425_));
  NOR2_X1    g13493(.A1(new_n15409_), .A2(new_n3707_), .ZN(new_n16426_));
  AOI22_X1   g13494(.A1(new_n15396_), .A2(new_n16426_), .B1(pi0299), .B2(new_n16425_), .ZN(new_n16427_));
  INV_X1     g13495(.I(new_n16422_), .ZN(new_n16428_));
  AOI21_X1   g13496(.A1(new_n3707_), .A2(new_n12133_), .B(new_n15722_), .ZN(new_n16429_));
  OAI21_X1   g13497(.A1(new_n15359_), .A2(new_n16429_), .B(new_n16428_), .ZN(new_n16430_));
  NAND2_X1   g13498(.A1(new_n16420_), .A2(new_n15410_), .ZN(new_n16431_));
  NAND2_X1   g13499(.A1(new_n16431_), .A2(new_n15726_), .ZN(new_n16432_));
  AOI21_X1   g13500(.A1(new_n16430_), .A2(new_n2566_), .B(new_n16432_), .ZN(new_n16433_));
  NOR2_X1    g13501(.A1(new_n12792_), .A2(pi0172), .ZN(new_n16434_));
  NOR2_X1    g13502(.A1(new_n15729_), .A2(new_n16434_), .ZN(new_n16435_));
  NAND2_X1   g13503(.A1(new_n3154_), .A2(new_n16415_), .ZN(new_n16436_));
  NOR4_X1    g13504(.A1(new_n16427_), .A2(new_n16433_), .A3(new_n16435_), .A4(new_n16436_), .ZN(new_n16437_));
  AOI21_X1   g13505(.A1(new_n12697_), .A2(new_n3707_), .B(pi0039), .ZN(new_n16438_));
  OR3_X2     g13506(.A1(new_n16438_), .A2(new_n12697_), .A3(new_n16412_), .Z(new_n16439_));
  NOR2_X1    g13507(.A1(new_n16439_), .A2(new_n15373_), .ZN(new_n16440_));
  OAI21_X1   g13508(.A1(new_n16437_), .A2(new_n16440_), .B(new_n3172_), .ZN(new_n16441_));
  NAND2_X1   g13509(.A1(new_n3707_), .A2(new_n16415_), .ZN(new_n16442_));
  OAI21_X1   g13510(.A1(new_n12894_), .A2(new_n16442_), .B(pi0039), .ZN(new_n16443_));
  NOR3_X1    g13511(.A1(new_n15434_), .A2(pi0299), .A3(new_n16419_), .ZN(new_n16444_));
  NAND2_X1   g13512(.A1(new_n16423_), .A2(new_n16415_), .ZN(new_n16445_));
  NOR4_X1    g13513(.A1(new_n15578_), .A2(new_n16422_), .A3(new_n16444_), .A4(new_n16445_), .ZN(new_n16446_));
  NOR3_X1    g13514(.A1(new_n16446_), .A2(new_n15494_), .A3(new_n16434_), .ZN(new_n16447_));
  INV_X1     g13515(.I(pi0690), .ZN(new_n16448_));
  NAND3_X1   g13516(.A1(new_n5156_), .A2(new_n2925_), .A3(new_n16412_), .ZN(new_n16449_));
  NAND4_X1   g13517(.A1(new_n12898_), .A2(new_n3172_), .A3(new_n3707_), .A4(new_n16449_), .ZN(new_n16450_));
  NAND4_X1   g13518(.A1(new_n16439_), .A2(new_n3172_), .A3(new_n16448_), .A4(new_n16450_), .ZN(new_n16451_));
  AOI21_X1   g13519(.A1(new_n16447_), .A2(new_n16443_), .B(new_n16451_), .ZN(new_n16452_));
  OAI21_X1   g13520(.A1(new_n16452_), .A2(new_n15500_), .B(pi0690), .ZN(new_n16453_));
  AOI21_X1   g13521(.A1(new_n16441_), .A2(new_n16418_), .B(new_n16453_), .ZN(new_n16454_));
  NAND2_X1   g13522(.A1(pi0057), .A2(pi0172), .ZN(new_n16455_));
  AOI21_X1   g13523(.A1(new_n16455_), .A2(new_n13184_), .B(pi0057), .ZN(new_n16456_));
  OAI21_X1   g13524(.A1(new_n15499_), .A2(pi0172), .B(new_n16456_), .ZN(new_n16457_));
  OAI21_X1   g13525(.A1(new_n16454_), .A2(new_n16457_), .B(new_n16414_), .ZN(po0329));
  NOR2_X1    g13526(.A1(new_n2925_), .A2(pi0173), .ZN(new_n16459_));
  NOR2_X1    g13527(.A1(new_n12054_), .A2(new_n16459_), .ZN(new_n16460_));
  NOR2_X1    g13528(.A1(new_n11877_), .A2(pi0745), .ZN(new_n16461_));
  NOR2_X1    g13529(.A1(new_n16461_), .A2(new_n16459_), .ZN(new_n16462_));
  NOR2_X1    g13530(.A1(new_n16462_), .A2(new_n11925_), .ZN(new_n16463_));
  NOR2_X1    g13531(.A1(new_n16463_), .A2(pi0785), .ZN(new_n16464_));
  INV_X1     g13532(.I(new_n16461_), .ZN(new_n16465_));
  NOR4_X1    g13533(.A1(new_n16463_), .A2(pi1155), .A3(new_n12997_), .A4(new_n16465_), .ZN(new_n16466_));
  NOR2_X1    g13534(.A1(new_n16465_), .A2(new_n12997_), .ZN(new_n16467_));
  OR3_X2     g13535(.A1(new_n16467_), .A2(pi1155), .A3(new_n16459_), .Z(new_n16468_));
  OAI21_X1   g13536(.A1(new_n16468_), .A2(new_n16466_), .B(pi0785), .ZN(new_n16469_));
  XNOR2_X1   g13537(.A1(new_n16469_), .A2(new_n16464_), .ZN(new_n16470_));
  INV_X1     g13538(.I(new_n16470_), .ZN(new_n16471_));
  NOR2_X1    g13539(.A1(new_n16471_), .A2(pi0781), .ZN(new_n16472_));
  OAI21_X1   g13540(.A1(new_n16471_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n16473_));
  NOR2_X1    g13541(.A1(new_n16471_), .A2(new_n11945_), .ZN(new_n16474_));
  OAI21_X1   g13542(.A1(new_n16473_), .A2(new_n16474_), .B(pi0781), .ZN(new_n16475_));
  XNOR2_X1   g13543(.A1(new_n16475_), .A2(new_n16472_), .ZN(new_n16476_));
  INV_X1     g13544(.I(new_n16476_), .ZN(new_n16477_));
  NOR2_X1    g13545(.A1(new_n16477_), .A2(pi0789), .ZN(new_n16478_));
  NOR2_X1    g13546(.A1(new_n2926_), .A2(new_n11967_), .ZN(new_n16479_));
  NAND2_X1   g13547(.A1(new_n16476_), .A2(new_n16479_), .ZN(new_n16480_));
  NAND2_X1   g13548(.A1(new_n16480_), .A2(new_n11869_), .ZN(new_n16481_));
  NAND3_X1   g13549(.A1(new_n2925_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n16482_));
  NOR2_X1    g13550(.A1(new_n16477_), .A2(new_n16482_), .ZN(new_n16483_));
  OAI21_X1   g13551(.A1(new_n16481_), .A2(new_n16483_), .B(pi0789), .ZN(new_n16484_));
  XNOR2_X1   g13552(.A1(new_n16484_), .A2(new_n16478_), .ZN(new_n16485_));
  NOR2_X1    g13553(.A1(new_n16485_), .A2(pi0788), .ZN(new_n16486_));
  INV_X1     g13554(.I(new_n16459_), .ZN(new_n16487_));
  MUX2_X1    g13555(.I0(new_n16485_), .I1(new_n16487_), .S(new_n12003_), .Z(new_n16488_));
  NOR2_X1    g13556(.A1(new_n16488_), .A2(new_n11986_), .ZN(new_n16489_));
  NOR2_X1    g13557(.A1(new_n16489_), .A2(new_n16486_), .ZN(new_n16490_));
  AOI21_X1   g13558(.A1(new_n16490_), .A2(new_n12054_), .B(new_n16460_), .ZN(new_n16491_));
  AOI21_X1   g13559(.A1(new_n11886_), .A2(new_n15593_), .B(new_n16459_), .ZN(new_n16492_));
  NOR3_X1    g13560(.A1(new_n11894_), .A2(pi0625), .A3(pi0723), .ZN(new_n16493_));
  NOR2_X1    g13561(.A1(new_n16459_), .A2(pi1153), .ZN(new_n16494_));
  INV_X1     g13562(.I(new_n16494_), .ZN(new_n16495_));
  NOR2_X1    g13563(.A1(new_n16493_), .A2(new_n16495_), .ZN(new_n16496_));
  INV_X1     g13564(.I(new_n16496_), .ZN(new_n16497_));
  OAI21_X1   g13565(.A1(new_n16493_), .A2(new_n16492_), .B(pi1153), .ZN(new_n16498_));
  NAND2_X1   g13566(.A1(new_n16497_), .A2(new_n16498_), .ZN(new_n16499_));
  MUX2_X1    g13567(.I0(new_n16499_), .I1(new_n16492_), .S(new_n11891_), .Z(new_n16500_));
  NOR2_X1    g13568(.A1(new_n16500_), .A2(new_n11939_), .ZN(new_n16501_));
  NAND2_X1   g13569(.A1(new_n16501_), .A2(new_n11963_), .ZN(new_n16502_));
  INV_X1     g13570(.I(new_n16502_), .ZN(new_n16503_));
  NOR2_X1    g13571(.A1(new_n16503_), .A2(new_n12034_), .ZN(new_n16504_));
  NAND2_X1   g13572(.A1(new_n16504_), .A2(new_n15050_), .ZN(new_n16505_));
  AOI21_X1   g13573(.A1(new_n16459_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n16506_));
  OAI21_X1   g13574(.A1(new_n16505_), .A2(new_n12061_), .B(new_n16506_), .ZN(new_n16507_));
  INV_X1     g13575(.I(new_n16505_), .ZN(new_n16508_));
  AOI21_X1   g13576(.A1(new_n16459_), .A2(pi0647), .B(pi1157), .ZN(new_n16509_));
  OAI21_X1   g13577(.A1(new_n16508_), .A2(new_n12061_), .B(new_n16509_), .ZN(new_n16510_));
  INV_X1     g13578(.I(new_n16510_), .ZN(new_n16511_));
  NOR2_X1    g13579(.A1(new_n16507_), .A2(pi0630), .ZN(new_n16512_));
  NOR2_X1    g13580(.A1(new_n16507_), .A2(pi0630), .ZN(new_n16513_));
  NOR3_X1    g13581(.A1(new_n16511_), .A2(new_n12060_), .A3(new_n16513_), .ZN(new_n16514_));
  NOR4_X1    g13582(.A1(new_n16491_), .A2(new_n15183_), .A3(new_n16512_), .A4(new_n16514_), .ZN(new_n16515_));
  NOR2_X1    g13583(.A1(new_n16492_), .A2(new_n11874_), .ZN(new_n16516_));
  INV_X1     g13584(.I(new_n16516_), .ZN(new_n16517_));
  NAND2_X1   g13585(.A1(new_n16517_), .A2(new_n16462_), .ZN(new_n16518_));
  NAND2_X1   g13586(.A1(new_n16518_), .A2(new_n11891_), .ZN(new_n16519_));
  NOR2_X1    g13587(.A1(new_n16517_), .A2(new_n12970_), .ZN(new_n16520_));
  NOR4_X1    g13588(.A1(new_n16520_), .A2(new_n11893_), .A3(new_n16459_), .A4(new_n16461_), .ZN(new_n16521_));
  NAND2_X1   g13589(.A1(new_n16497_), .A2(pi0608), .ZN(new_n16522_));
  INV_X1     g13590(.I(new_n16520_), .ZN(new_n16523_));
  AOI21_X1   g13591(.A1(new_n16523_), .A2(new_n16518_), .B(new_n16495_), .ZN(new_n16524_));
  NAND2_X1   g13592(.A1(new_n16498_), .A2(new_n13657_), .ZN(new_n16525_));
  OAI22_X1   g13593(.A1(new_n16524_), .A2(new_n16525_), .B1(new_n16521_), .B2(new_n16522_), .ZN(new_n16526_));
  NAND2_X1   g13594(.A1(new_n16526_), .A2(pi0778), .ZN(new_n16527_));
  XOR2_X1    g13595(.A1(new_n16527_), .A2(new_n16519_), .Z(new_n16528_));
  INV_X1     g13596(.I(new_n16528_), .ZN(new_n16529_));
  XNOR2_X1   g13597(.A1(new_n16528_), .A2(new_n16500_), .ZN(new_n16530_));
  NAND2_X1   g13598(.A1(new_n16530_), .A2(pi0609), .ZN(new_n16531_));
  XOR2_X1    g13599(.A1(new_n16531_), .A2(new_n16529_), .Z(new_n16532_));
  NOR2_X1    g13600(.A1(new_n16466_), .A2(pi0660), .ZN(new_n16533_));
  OAI21_X1   g13601(.A1(new_n16532_), .A2(pi1155), .B(new_n16533_), .ZN(new_n16534_));
  NOR4_X1    g13602(.A1(new_n16467_), .A2(new_n11923_), .A3(pi1155), .A4(new_n16459_), .ZN(new_n16536_));
  NOR2_X1    g13603(.A1(new_n16536_), .A2(new_n11870_), .ZN(new_n16537_));
  AOI22_X1   g13604(.A1(new_n16534_), .A2(new_n16537_), .B1(new_n11870_), .B2(new_n16529_), .ZN(new_n16538_));
  NOR2_X1    g13605(.A1(new_n16538_), .A2(pi0781), .ZN(new_n16539_));
  NOR4_X1    g13606(.A1(new_n16500_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n16540_));
  OAI21_X1   g13607(.A1(new_n16471_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n16541_));
  NOR4_X1    g13608(.A1(new_n16538_), .A2(new_n11934_), .A3(pi1154), .A4(new_n16501_), .ZN(new_n16542_));
  NOR2_X1    g13609(.A1(new_n16542_), .A2(new_n16473_), .ZN(new_n16543_));
  OAI22_X1   g13610(.A1(new_n16543_), .A2(pi0627), .B1(new_n16540_), .B2(new_n16541_), .ZN(new_n16544_));
  AOI21_X1   g13611(.A1(new_n16544_), .A2(pi0781), .B(new_n16539_), .ZN(new_n16545_));
  INV_X1     g13612(.I(new_n16545_), .ZN(new_n16546_));
  NAND4_X1   g13613(.A1(new_n16546_), .A2(pi0619), .A3(new_n11869_), .A4(new_n16502_), .ZN(new_n16547_));
  NOR2_X1    g13614(.A1(new_n16481_), .A2(new_n11966_), .ZN(new_n16548_));
  NAND3_X1   g13615(.A1(new_n16503_), .A2(pi0619), .A3(pi1159), .ZN(new_n16549_));
  NOR2_X1    g13616(.A1(new_n16483_), .A2(pi0648), .ZN(new_n16550_));
  AOI22_X1   g13617(.A1(new_n16547_), .A2(new_n16548_), .B1(new_n16549_), .B2(new_n16550_), .ZN(new_n16551_));
  OAI21_X1   g13618(.A1(new_n16546_), .A2(new_n11999_), .B(new_n11985_), .ZN(new_n16552_));
  NOR2_X1    g13619(.A1(new_n16488_), .A2(new_n11991_), .ZN(new_n16553_));
  OAI21_X1   g13620(.A1(new_n16502_), .A2(new_n12022_), .B(pi0788), .ZN(new_n16554_));
  OAI22_X1   g13621(.A1(new_n16551_), .A2(new_n16552_), .B1(new_n16553_), .B2(new_n16554_), .ZN(new_n16555_));
  NAND2_X1   g13622(.A1(new_n16504_), .A2(new_n15080_), .ZN(new_n16556_));
  OAI21_X1   g13623(.A1(new_n16489_), .A2(new_n16486_), .B(new_n12064_), .ZN(new_n16557_));
  AOI21_X1   g13624(.A1(new_n16557_), .A2(new_n16556_), .B(new_n12030_), .ZN(new_n16558_));
  INV_X1     g13625(.I(new_n12063_), .ZN(new_n16559_));
  AOI21_X1   g13626(.A1(new_n16504_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n16560_));
  OAI21_X1   g13627(.A1(new_n16490_), .A2(new_n16559_), .B(new_n16560_), .ZN(new_n16561_));
  OAI21_X1   g13628(.A1(new_n16558_), .A2(new_n16561_), .B(new_n14726_), .ZN(new_n16562_));
  AOI21_X1   g13629(.A1(new_n16555_), .A2(new_n14732_), .B(new_n16562_), .ZN(new_n16563_));
  OR2_X2     g13630(.A1(new_n16563_), .A2(new_n16515_), .Z(new_n16564_));
  NAND2_X1   g13631(.A1(new_n16564_), .A2(pi0644), .ZN(new_n16565_));
  AND2_X2    g13632(.A1(new_n16507_), .A2(pi0787), .Z(new_n16566_));
  AOI22_X1   g13633(.A1(new_n16566_), .A2(new_n16511_), .B1(new_n12048_), .B2(new_n16508_), .ZN(new_n16567_));
  NAND2_X1   g13634(.A1(new_n16567_), .A2(new_n12082_), .ZN(new_n16568_));
  AND3_X2    g13635(.A1(new_n16565_), .A2(new_n12099_), .A3(new_n16568_), .Z(new_n16569_));
  NOR2_X1    g13636(.A1(new_n16491_), .A2(new_n12091_), .ZN(new_n16570_));
  NOR2_X1    g13637(.A1(new_n12092_), .A2(new_n16459_), .ZN(new_n16571_));
  NOR2_X1    g13638(.A1(new_n16570_), .A2(new_n16571_), .ZN(new_n16572_));
  OAI21_X1   g13639(.A1(new_n16572_), .A2(new_n16459_), .B(new_n12082_), .ZN(new_n16573_));
  AOI21_X1   g13640(.A1(new_n16459_), .A2(new_n16572_), .B(new_n16573_), .ZN(new_n16574_));
  OAI21_X1   g13641(.A1(new_n16570_), .A2(new_n16571_), .B(new_n16574_), .ZN(new_n16575_));
  OAI21_X1   g13642(.A1(pi0644), .A2(new_n16459_), .B(new_n16572_), .ZN(new_n16576_));
  NAND3_X1   g13643(.A1(new_n16575_), .A2(new_n12099_), .A3(new_n16576_), .ZN(new_n16577_));
  OAI21_X1   g13644(.A1(new_n16569_), .A2(new_n16577_), .B(new_n12081_), .ZN(new_n16578_));
  XOR2_X1    g13645(.A1(new_n16574_), .A2(new_n16487_), .Z(new_n16579_));
  OAI21_X1   g13646(.A1(new_n16567_), .A2(new_n12082_), .B(new_n13168_), .ZN(new_n16580_));
  AOI21_X1   g13647(.A1(new_n16579_), .A2(pi0715), .B(new_n16580_), .ZN(new_n16581_));
  AOI21_X1   g13648(.A1(new_n16581_), .A2(new_n16565_), .B(new_n11867_), .ZN(new_n16582_));
  NAND2_X1   g13649(.A1(new_n16564_), .A2(new_n14747_), .ZN(new_n16583_));
  AOI21_X1   g13650(.A1(new_n16578_), .A2(new_n16582_), .B(new_n16583_), .ZN(new_n16584_));
  NOR2_X1    g13651(.A1(new_n12965_), .A2(pi0173), .ZN(new_n16585_));
  AOI21_X1   g13652(.A1(new_n12694_), .A2(pi0173), .B(new_n15596_), .ZN(new_n16586_));
  OAI21_X1   g13653(.A1(pi0173), .A2(new_n15144_), .B(new_n16586_), .ZN(new_n16587_));
  NOR2_X1    g13654(.A1(new_n12828_), .A2(pi0173), .ZN(new_n16588_));
  AOI21_X1   g13655(.A1(new_n15596_), .A2(new_n12829_), .B(new_n16588_), .ZN(new_n16589_));
  MUX2_X1    g13656(.I0(new_n16589_), .I1(new_n16587_), .S(new_n3172_), .Z(new_n16590_));
  NOR2_X1    g13657(.A1(new_n16590_), .A2(new_n3232_), .ZN(new_n16591_));
  AOI21_X1   g13658(.A1(new_n10056_), .A2(new_n3232_), .B(new_n16591_), .ZN(new_n16592_));
  INV_X1     g13659(.I(new_n16592_), .ZN(new_n16593_));
  INV_X1     g13660(.I(new_n16585_), .ZN(new_n16594_));
  OAI21_X1   g13661(.A1(new_n16594_), .A2(new_n11924_), .B(new_n11870_), .ZN(new_n16595_));
  AOI21_X1   g13662(.A1(new_n16593_), .A2(new_n11924_), .B(new_n16595_), .ZN(new_n16596_));
  NAND2_X1   g13663(.A1(new_n16592_), .A2(new_n11924_), .ZN(new_n16597_));
  OAI22_X1   g13664(.A1(new_n16597_), .A2(pi0609), .B1(new_n12996_), .B2(new_n16585_), .ZN(new_n16598_));
  NAND2_X1   g13665(.A1(new_n16598_), .A2(new_n11912_), .ZN(new_n16599_));
  OAI22_X1   g13666(.A1(new_n16597_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n16585_), .ZN(new_n16600_));
  NAND2_X1   g13667(.A1(new_n16600_), .A2(pi1155), .ZN(new_n16601_));
  NAND2_X1   g13668(.A1(new_n16599_), .A2(new_n16601_), .ZN(new_n16602_));
  NAND2_X1   g13669(.A1(new_n16602_), .A2(pi0785), .ZN(new_n16603_));
  XOR2_X1    g13670(.A1(new_n16603_), .A2(new_n16596_), .Z(new_n16604_));
  NAND2_X1   g13671(.A1(new_n16604_), .A2(new_n11969_), .ZN(new_n16605_));
  MUX2_X1    g13672(.I0(new_n16604_), .I1(new_n16585_), .S(new_n15166_), .Z(new_n16606_));
  NAND2_X1   g13673(.A1(new_n16606_), .A2(pi0781), .ZN(new_n16607_));
  NAND2_X1   g13674(.A1(new_n16607_), .A2(new_n16605_), .ZN(new_n16608_));
  NAND2_X1   g13675(.A1(new_n16608_), .A2(new_n11985_), .ZN(new_n16609_));
  INV_X1     g13676(.I(new_n16608_), .ZN(new_n16610_));
  MUX2_X1    g13677(.I0(new_n16594_), .I1(new_n16610_), .S(new_n14640_), .Z(new_n16611_));
  OAI21_X1   g13678(.A1(new_n16611_), .A2(new_n11985_), .B(new_n16609_), .ZN(new_n16612_));
  AND2_X2    g13679(.A1(new_n16612_), .A2(new_n11986_), .Z(new_n16613_));
  MUX2_X1    g13680(.I0(new_n16612_), .I1(new_n16585_), .S(new_n12003_), .Z(new_n16614_));
  AOI21_X1   g13681(.A1(new_n16614_), .A2(pi0788), .B(new_n16613_), .ZN(new_n16615_));
  NAND2_X1   g13682(.A1(new_n16615_), .A2(new_n12054_), .ZN(new_n16616_));
  OAI21_X1   g13683(.A1(new_n12054_), .A2(new_n16585_), .B(new_n16616_), .ZN(new_n16617_));
  NOR2_X1    g13684(.A1(new_n16585_), .A2(new_n12092_), .ZN(new_n16618_));
  AOI21_X1   g13685(.A1(new_n16617_), .A2(new_n12092_), .B(new_n16618_), .ZN(new_n16619_));
  NOR3_X1    g13686(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n16620_));
  NAND2_X1   g13687(.A1(new_n16619_), .A2(new_n16620_), .ZN(new_n16621_));
  NOR2_X1    g13688(.A1(new_n16594_), .A2(pi0647), .ZN(new_n16622_));
  OAI21_X1   g13689(.A1(new_n13395_), .A2(new_n10056_), .B(new_n3172_), .ZN(new_n16623_));
  NAND2_X1   g13690(.A1(new_n16623_), .A2(new_n3231_), .ZN(new_n16624_));
  NOR2_X1    g13691(.A1(new_n13399_), .A2(pi0173), .ZN(new_n16625_));
  INV_X1     g13692(.I(new_n16625_), .ZN(new_n16626_));
  OAI21_X1   g13693(.A1(new_n15189_), .A2(new_n16588_), .B(new_n15593_), .ZN(new_n16627_));
  AOI21_X1   g13694(.A1(new_n16626_), .A2(new_n16624_), .B(new_n16627_), .ZN(new_n16628_));
  NOR2_X1    g13695(.A1(new_n3232_), .A2(pi0723), .ZN(new_n16629_));
  AOI21_X1   g13696(.A1(new_n16594_), .A2(new_n16629_), .B(new_n16628_), .ZN(new_n16630_));
  NOR3_X1    g13697(.A1(new_n16594_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n16631_));
  NOR4_X1    g13698(.A1(new_n16630_), .A2(new_n12970_), .A3(pi1153), .A4(new_n16585_), .ZN(new_n16632_));
  NOR2_X1    g13699(.A1(new_n16632_), .A2(new_n16631_), .ZN(new_n16633_));
  MUX2_X1    g13700(.I0(new_n16633_), .I1(new_n16630_), .S(new_n11891_), .Z(new_n16634_));
  NOR2_X1    g13701(.A1(new_n16634_), .A2(new_n13024_), .ZN(new_n16635_));
  AOI21_X1   g13702(.A1(new_n13024_), .A2(new_n16585_), .B(new_n16635_), .ZN(new_n16636_));
  INV_X1     g13703(.I(new_n16636_), .ZN(new_n16637_));
  NOR2_X1    g13704(.A1(new_n16637_), .A2(new_n13714_), .ZN(new_n16638_));
  AOI21_X1   g13705(.A1(new_n13714_), .A2(new_n16594_), .B(new_n16638_), .ZN(new_n16639_));
  NAND2_X1   g13706(.A1(new_n16639_), .A2(new_n12032_), .ZN(new_n16640_));
  NAND2_X1   g13707(.A1(new_n16585_), .A2(new_n13713_), .ZN(new_n16641_));
  XNOR2_X1   g13708(.A1(new_n16640_), .A2(new_n16641_), .ZN(new_n16642_));
  NOR3_X1    g13709(.A1(new_n16594_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n16644_));
  INV_X1     g13710(.I(new_n16644_), .ZN(new_n16645_));
  NAND4_X1   g13711(.A1(new_n16642_), .A2(pi0628), .A3(new_n12026_), .A4(new_n16594_), .ZN(new_n16646_));
  NAND2_X1   g13712(.A1(new_n16646_), .A2(new_n16645_), .ZN(new_n16647_));
  MUX2_X1    g13713(.I0(new_n16647_), .I1(new_n16642_), .S(new_n11868_), .Z(new_n16648_));
  AOI21_X1   g13714(.A1(new_n16648_), .A2(pi0647), .B(new_n16622_), .ZN(new_n16649_));
  NAND2_X1   g13715(.A1(new_n16649_), .A2(new_n12060_), .ZN(new_n16650_));
  NOR2_X1    g13716(.A1(new_n16594_), .A2(new_n12061_), .ZN(new_n16651_));
  AOI21_X1   g13717(.A1(new_n16648_), .A2(new_n12061_), .B(new_n16651_), .ZN(new_n16652_));
  AOI21_X1   g13718(.A1(new_n16652_), .A2(pi0630), .B(new_n15214_), .ZN(new_n16653_));
  AOI21_X1   g13719(.A1(new_n16653_), .A2(new_n16650_), .B(new_n15183_), .ZN(new_n16654_));
  NAND2_X1   g13720(.A1(new_n16617_), .A2(new_n16654_), .ZN(new_n16655_));
  NOR2_X1    g13721(.A1(new_n16644_), .A2(new_n12030_), .ZN(new_n16656_));
  AND2_X2    g13722(.A1(new_n16646_), .A2(new_n12030_), .Z(new_n16657_));
  OAI21_X1   g13723(.A1(new_n16657_), .A2(new_n16656_), .B(new_n11868_), .ZN(new_n16658_));
  AOI21_X1   g13724(.A1(new_n16615_), .A2(new_n15222_), .B(new_n16658_), .ZN(new_n16659_));
  INV_X1     g13725(.I(new_n16639_), .ZN(new_n16660_));
  NOR3_X1    g13726(.A1(new_n16660_), .A2(new_n12013_), .A3(new_n16594_), .ZN(new_n16661_));
  AOI21_X1   g13727(.A1(new_n12014_), .A2(new_n16594_), .B(new_n16639_), .ZN(new_n16662_));
  OAI21_X1   g13728(.A1(new_n16661_), .A2(new_n16662_), .B(new_n12020_), .ZN(new_n16663_));
  NAND2_X1   g13729(.A1(new_n16614_), .A2(new_n12002_), .ZN(new_n16664_));
  AOI21_X1   g13730(.A1(new_n16664_), .A2(new_n16663_), .B(pi0788), .ZN(new_n16665_));
  NOR3_X1    g13731(.A1(new_n16590_), .A2(new_n15593_), .A3(new_n3231_), .ZN(new_n16675_));
  AOI21_X1   g13732(.A1(pi0173), .A2(new_n3232_), .B(new_n16675_), .ZN(new_n16676_));
  INV_X1     g13733(.I(new_n16632_), .ZN(new_n16677_));
  NAND2_X1   g13734(.A1(new_n16676_), .A2(pi0625), .ZN(new_n16678_));
  NAND2_X1   g13735(.A1(new_n16593_), .A2(pi0625), .ZN(new_n16679_));
  NAND4_X1   g13736(.A1(new_n16679_), .A2(new_n12977_), .A3(new_n16677_), .A4(new_n16678_), .ZN(new_n16680_));
  NAND2_X1   g13737(.A1(new_n16592_), .A2(new_n12970_), .ZN(new_n16681_));
  AND3_X2    g13738(.A1(new_n16678_), .A2(new_n11893_), .A3(new_n16681_), .Z(new_n16682_));
  OAI21_X1   g13739(.A1(new_n16682_), .A2(new_n16631_), .B(new_n13657_), .ZN(new_n16683_));
  AOI21_X1   g13740(.A1(new_n16683_), .A2(new_n16680_), .B(new_n11891_), .ZN(new_n16684_));
  AOI21_X1   g13741(.A1(new_n11891_), .A2(new_n16676_), .B(new_n16684_), .ZN(new_n16685_));
  INV_X1     g13742(.I(new_n16634_), .ZN(new_n16686_));
  NOR4_X1    g13743(.A1(new_n16685_), .A2(new_n11903_), .A3(pi1155), .A4(new_n16686_), .ZN(new_n16687_));
  NAND2_X1   g13744(.A1(new_n16599_), .A2(pi0660), .ZN(new_n16688_));
  NOR3_X1    g13745(.A1(new_n16634_), .A2(new_n11903_), .A3(new_n11912_), .ZN(new_n16689_));
  NAND2_X1   g13746(.A1(new_n16601_), .A2(new_n11923_), .ZN(new_n16690_));
  OAI22_X1   g13747(.A1(new_n16687_), .A2(new_n16688_), .B1(new_n16689_), .B2(new_n16690_), .ZN(new_n16691_));
  MUX2_X1    g13748(.I0(new_n16691_), .I1(new_n16685_), .S(new_n11870_), .Z(new_n16692_));
  INV_X1     g13749(.I(new_n16692_), .ZN(new_n16693_));
  AOI21_X1   g13750(.A1(new_n16637_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n16694_));
  INV_X1     g13751(.I(new_n16604_), .ZN(new_n16695_));
  NAND3_X1   g13752(.A1(new_n11934_), .A2(new_n11949_), .A3(pi1154), .ZN(new_n16696_));
  OAI21_X1   g13753(.A1(new_n16695_), .A2(new_n16696_), .B(pi0618), .ZN(new_n16697_));
  NOR2_X1    g13754(.A1(new_n16697_), .A2(new_n16694_), .ZN(new_n16698_));
  NAND2_X1   g13755(.A1(new_n16692_), .A2(new_n11934_), .ZN(new_n16699_));
  NOR2_X1    g13756(.A1(new_n16636_), .A2(new_n11934_), .ZN(new_n16700_));
  NAND2_X1   g13757(.A1(new_n11950_), .A2(pi0618), .ZN(new_n16701_));
  NOR2_X1    g13758(.A1(new_n16695_), .A2(new_n16701_), .ZN(new_n16702_));
  NOR4_X1    g13759(.A1(new_n16702_), .A2(pi0627), .A3(pi1154), .A4(new_n16700_), .ZN(new_n16703_));
  AOI22_X1   g13760(.A1(new_n16699_), .A2(new_n16703_), .B1(new_n16692_), .B2(new_n16698_), .ZN(new_n16704_));
  MUX2_X1    g13761(.I0(new_n16704_), .I1(new_n16693_), .S(new_n11969_), .Z(new_n16705_));
  NAND3_X1   g13762(.A1(new_n11967_), .A2(new_n11966_), .A3(pi1159), .ZN(new_n16706_));
  NOR2_X1    g13763(.A1(new_n16610_), .A2(new_n16706_), .ZN(new_n16707_));
  NAND2_X1   g13764(.A1(new_n11869_), .A2(pi0619), .ZN(new_n16708_));
  OR3_X2     g13765(.A1(new_n16705_), .A2(new_n16707_), .A3(new_n16708_), .Z(new_n16709_));
  NOR2_X1    g13766(.A1(new_n11967_), .A2(pi1159), .ZN(new_n16710_));
  OAI21_X1   g13767(.A1(new_n16660_), .A2(new_n11967_), .B(new_n15278_), .ZN(new_n16711_));
  AOI21_X1   g13768(.A1(new_n16608_), .A2(new_n16710_), .B(new_n16711_), .ZN(new_n16712_));
  OAI21_X1   g13769(.A1(new_n16705_), .A2(pi0619), .B(new_n16712_), .ZN(new_n16713_));
  OAI21_X1   g13770(.A1(new_n16705_), .A2(new_n11999_), .B(new_n11985_), .ZN(new_n16714_));
  AOI21_X1   g13771(.A1(new_n16709_), .A2(new_n16713_), .B(new_n16714_), .ZN(new_n16715_));
  NOR4_X1    g13772(.A1(new_n16659_), .A2(new_n16665_), .A3(new_n14731_), .A4(new_n16715_), .ZN(new_n16716_));
  OAI21_X1   g13773(.A1(new_n16716_), .A2(new_n14725_), .B(new_n16655_), .ZN(new_n16717_));
  NOR4_X1    g13774(.A1(new_n16717_), .A2(new_n16621_), .A3(new_n12082_), .A4(pi0790), .ZN(new_n16718_));
  NAND2_X1   g13775(.A1(new_n16649_), .A2(pi1157), .ZN(new_n16719_));
  NAND2_X1   g13776(.A1(new_n16652_), .A2(new_n12049_), .ZN(new_n16720_));
  NAND2_X1   g13777(.A1(new_n16719_), .A2(new_n16720_), .ZN(new_n16721_));
  NOR2_X1    g13778(.A1(new_n16648_), .A2(pi0787), .ZN(new_n16722_));
  AOI21_X1   g13779(.A1(new_n16721_), .A2(pi0787), .B(new_n16722_), .ZN(new_n16723_));
  AOI21_X1   g13780(.A1(new_n16723_), .A2(new_n12082_), .B(new_n12099_), .ZN(new_n16724_));
  NAND2_X1   g13781(.A1(new_n16621_), .A2(new_n16724_), .ZN(new_n16725_));
  INV_X1     g13782(.I(new_n16723_), .ZN(new_n16726_));
  NAND3_X1   g13783(.A1(new_n16717_), .A2(new_n12082_), .A3(new_n16726_), .ZN(new_n16727_));
  OAI21_X1   g13784(.A1(new_n16717_), .A2(pi0644), .B(new_n16723_), .ZN(new_n16728_));
  NOR2_X1    g13785(.A1(new_n12081_), .A2(pi0715), .ZN(new_n16731_));
  NAND3_X1   g13786(.A1(new_n16728_), .A2(new_n16727_), .A3(new_n16731_), .ZN(new_n16732_));
  AOI21_X1   g13787(.A1(new_n16732_), .A2(new_n16725_), .B(new_n11867_), .ZN(new_n16733_));
  OAI21_X1   g13788(.A1(new_n16733_), .A2(new_n16718_), .B(new_n6845_), .ZN(new_n16734_));
  AOI21_X1   g13789(.A1(po1038), .A2(new_n10056_), .B(pi0832), .ZN(new_n16735_));
  AOI21_X1   g13790(.A1(new_n16734_), .A2(new_n16735_), .B(new_n16584_), .ZN(po0330));
  NOR2_X1    g13791(.A1(new_n2925_), .A2(new_n7151_), .ZN(new_n16737_));
  NOR2_X1    g13792(.A1(new_n11894_), .A2(new_n15674_), .ZN(new_n16738_));
  NOR2_X1    g13793(.A1(new_n16738_), .A2(new_n16737_), .ZN(new_n16739_));
  INV_X1     g13794(.I(new_n16739_), .ZN(new_n16740_));
  INV_X1     g13795(.I(new_n16738_), .ZN(new_n16741_));
  NOR3_X1    g13796(.A1(new_n16741_), .A2(new_n13659_), .A3(new_n16737_), .ZN(new_n16742_));
  INV_X1     g13797(.I(new_n16737_), .ZN(new_n16743_));
  NOR3_X1    g13798(.A1(new_n16738_), .A2(new_n12970_), .A3(new_n16743_), .ZN(new_n16744_));
  AOI21_X1   g13799(.A1(new_n16741_), .A2(new_n16743_), .B(pi0625), .ZN(new_n16745_));
  NOR3_X1    g13800(.A1(new_n16745_), .A2(pi1153), .A3(new_n16744_), .ZN(new_n16746_));
  INV_X1     g13801(.I(new_n16746_), .ZN(new_n16747_));
  NOR2_X1    g13802(.A1(new_n16747_), .A2(new_n16742_), .ZN(new_n16748_));
  MUX2_X1    g13803(.I0(new_n16748_), .I1(new_n16740_), .S(new_n11891_), .Z(new_n16749_));
  NOR2_X1    g13804(.A1(new_n16749_), .A2(new_n13717_), .ZN(new_n16750_));
  INV_X1     g13805(.I(new_n16750_), .ZN(new_n16751_));
  NOR2_X1    g13806(.A1(new_n16751_), .A2(new_n12066_), .ZN(new_n16752_));
  AOI21_X1   g13807(.A1(new_n16752_), .A2(new_n13748_), .B(new_n16737_), .ZN(new_n16753_));
  INV_X1     g13808(.I(new_n16753_), .ZN(new_n16754_));
  NOR2_X1    g13809(.A1(new_n11877_), .A2(new_n15660_), .ZN(new_n16755_));
  INV_X1     g13810(.I(new_n16755_), .ZN(new_n16756_));
  NOR2_X1    g13811(.A1(new_n16756_), .A2(new_n14627_), .ZN(new_n16757_));
  INV_X1     g13812(.I(new_n16757_), .ZN(new_n16758_));
  NOR2_X1    g13813(.A1(new_n16758_), .A2(new_n14644_), .ZN(new_n16759_));
  INV_X1     g13814(.I(new_n16759_), .ZN(new_n16760_));
  NOR2_X1    g13815(.A1(new_n16760_), .A2(new_n11997_), .ZN(new_n16761_));
  NOR3_X1    g13816(.A1(new_n12053_), .A2(new_n12060_), .A3(pi1157), .ZN(new_n16762_));
  AOI21_X1   g13817(.A1(new_n16761_), .A2(new_n16762_), .B(new_n12061_), .ZN(new_n16763_));
  OAI21_X1   g13818(.A1(new_n16752_), .A2(pi0630), .B(new_n16763_), .ZN(new_n16764_));
  OAI21_X1   g13819(.A1(new_n12053_), .A2(pi0630), .B(new_n12061_), .ZN(new_n16765_));
  OAI22_X1   g13820(.A1(new_n16752_), .A2(new_n12060_), .B1(new_n16761_), .B2(new_n16765_), .ZN(new_n16766_));
  NAND2_X1   g13821(.A1(new_n16766_), .A2(new_n12049_), .ZN(new_n16767_));
  NAND2_X1   g13822(.A1(new_n16767_), .A2(new_n16764_), .ZN(new_n16768_));
  NOR2_X1    g13823(.A1(new_n16737_), .A2(new_n12048_), .ZN(new_n16769_));
  NOR2_X1    g13824(.A1(new_n16750_), .A2(new_n12030_), .ZN(new_n16770_));
  OAI22_X1   g13825(.A1(new_n16770_), .A2(pi0628), .B1(new_n12030_), .B2(new_n16761_), .ZN(new_n16771_));
  INV_X1     g13826(.I(new_n16771_), .ZN(new_n16772_));
  NOR2_X1    g13827(.A1(new_n16761_), .A2(pi0628), .ZN(new_n16773_));
  OAI22_X1   g13828(.A1(new_n16751_), .A2(new_n12031_), .B1(new_n12030_), .B2(new_n16773_), .ZN(new_n16774_));
  OAI21_X1   g13829(.A1(new_n12026_), .A2(new_n16774_), .B(new_n16772_), .ZN(new_n16775_));
  NAND3_X1   g13830(.A1(new_n16771_), .A2(new_n16774_), .A3(pi1156), .ZN(new_n16776_));
  NAND4_X1   g13831(.A1(new_n16775_), .A2(pi0792), .A3(new_n16776_), .A4(new_n16743_), .ZN(new_n16777_));
  INV_X1     g13832(.I(new_n16749_), .ZN(new_n16778_));
  AOI21_X1   g13833(.A1(new_n16778_), .A2(new_n11938_), .B(new_n16737_), .ZN(new_n16779_));
  NAND2_X1   g13834(.A1(new_n12118_), .A2(pi0696), .ZN(new_n16780_));
  AND3_X2    g13835(.A1(new_n16780_), .A2(new_n16743_), .A3(new_n16756_), .Z(new_n16781_));
  NOR2_X1    g13836(.A1(new_n13649_), .A2(new_n15674_), .ZN(new_n16782_));
  NAND3_X1   g13837(.A1(new_n16756_), .A2(pi1153), .A3(new_n16743_), .ZN(new_n16783_));
  OAI21_X1   g13838(.A1(new_n16782_), .A2(new_n16783_), .B(pi0608), .ZN(new_n16784_));
  INV_X1     g13839(.I(new_n16781_), .ZN(new_n16785_));
  NOR2_X1    g13840(.A1(new_n16785_), .A2(new_n16782_), .ZN(new_n16786_));
  OAI21_X1   g13841(.A1(new_n16742_), .A2(pi0608), .B(new_n11893_), .ZN(new_n16787_));
  OAI22_X1   g13842(.A1(new_n16747_), .A2(new_n16784_), .B1(new_n16786_), .B2(new_n16787_), .ZN(new_n16788_));
  MUX2_X1    g13843(.I0(new_n16788_), .I1(new_n16781_), .S(new_n11891_), .Z(new_n16789_));
  NOR3_X1    g13844(.A1(new_n16749_), .A2(new_n11903_), .A3(new_n11912_), .ZN(new_n16790_));
  NOR4_X1    g13845(.A1(new_n16756_), .A2(pi1155), .A3(new_n13010_), .A4(new_n16737_), .ZN(new_n16791_));
  NOR3_X1    g13846(.A1(new_n16790_), .A2(pi0660), .A3(new_n16791_), .ZN(new_n16792_));
  NOR4_X1    g13847(.A1(new_n16789_), .A2(new_n11903_), .A3(pi1155), .A4(new_n16778_), .ZN(new_n16793_));
  NOR2_X1    g13848(.A1(new_n16737_), .A2(new_n14671_), .ZN(new_n16794_));
  OAI21_X1   g13849(.A1(new_n16756_), .A2(new_n12997_), .B(new_n16794_), .ZN(new_n16795_));
  OAI21_X1   g13850(.A1(new_n16793_), .A2(new_n16795_), .B(pi0785), .ZN(new_n16796_));
  OAI22_X1   g13851(.A1(new_n16796_), .A2(new_n16792_), .B1(pi0785), .B2(new_n16789_), .ZN(new_n16797_));
  MUX2_X1    g13852(.I0(new_n16797_), .I1(new_n16779_), .S(new_n11934_), .Z(new_n16798_));
  NOR2_X1    g13853(.A1(new_n16737_), .A2(new_n14687_), .ZN(new_n16799_));
  OAI21_X1   g13854(.A1(new_n16758_), .A2(new_n14686_), .B(new_n16799_), .ZN(new_n16800_));
  AOI21_X1   g13855(.A1(new_n16798_), .A2(pi1154), .B(new_n16800_), .ZN(new_n16801_));
  MUX2_X1    g13856(.I0(new_n16797_), .I1(new_n16779_), .S(pi0618), .Z(new_n16802_));
  NAND4_X1   g13857(.A1(new_n11924_), .A2(pi0618), .A3(new_n11950_), .A4(new_n16743_), .ZN(new_n16803_));
  OAI21_X1   g13858(.A1(new_n16758_), .A2(new_n16803_), .B(new_n11949_), .ZN(new_n16804_));
  AOI21_X1   g13859(.A1(new_n16802_), .A2(new_n11950_), .B(new_n16804_), .ZN(new_n16805_));
  OR2_X2     g13860(.A1(new_n16801_), .A2(new_n16805_), .Z(new_n16806_));
  NOR2_X1    g13861(.A1(new_n11967_), .A2(pi0648), .ZN(new_n16807_));
  NOR2_X1    g13862(.A1(new_n11966_), .A2(pi0619), .ZN(new_n16808_));
  NOR2_X1    g13863(.A1(new_n16807_), .A2(new_n16808_), .ZN(new_n16809_));
  AOI21_X1   g13864(.A1(new_n16809_), .A2(new_n14640_), .B(new_n11985_), .ZN(new_n16810_));
  INV_X1     g13865(.I(new_n16810_), .ZN(new_n16811_));
  OAI21_X1   g13866(.A1(new_n16797_), .A2(pi0781), .B(new_n16811_), .ZN(new_n16812_));
  AOI21_X1   g13867(.A1(new_n16806_), .A2(pi0781), .B(new_n16812_), .ZN(new_n16813_));
  NOR2_X1    g13868(.A1(new_n16749_), .A2(new_n13716_), .ZN(new_n16814_));
  AOI21_X1   g13869(.A1(new_n16757_), .A2(new_n14697_), .B(pi0648), .ZN(new_n16815_));
  INV_X1     g13870(.I(new_n14702_), .ZN(new_n16816_));
  OAI21_X1   g13871(.A1(new_n16758_), .A2(new_n16816_), .B(pi0648), .ZN(new_n16817_));
  NAND2_X1   g13872(.A1(new_n16817_), .A2(new_n12012_), .ZN(new_n16818_));
  NOR4_X1    g13873(.A1(new_n14640_), .A2(new_n16737_), .A3(new_n16809_), .A4(pi0789), .ZN(new_n16819_));
  OAI21_X1   g13874(.A1(new_n16818_), .A2(new_n16815_), .B(new_n16819_), .ZN(new_n16820_));
  NOR2_X1    g13875(.A1(new_n16814_), .A2(new_n16820_), .ZN(new_n16821_));
  INV_X1     g13876(.I(new_n11993_), .ZN(new_n16822_));
  AOI21_X1   g13877(.A1(new_n16814_), .A2(new_n12014_), .B(new_n16737_), .ZN(new_n16823_));
  OAI21_X1   g13878(.A1(new_n16760_), .A2(pi0626), .B(new_n16743_), .ZN(new_n16824_));
  NAND2_X1   g13879(.A1(new_n16824_), .A2(new_n11987_), .ZN(new_n16825_));
  NAND4_X1   g13880(.A1(new_n16823_), .A2(new_n11989_), .A3(new_n16822_), .A4(new_n16825_), .ZN(new_n16826_));
  INV_X1     g13881(.I(new_n11995_), .ZN(new_n16827_));
  NAND2_X1   g13882(.A1(new_n16823_), .A2(new_n16827_), .ZN(new_n16828_));
  OAI21_X1   g13883(.A1(new_n16760_), .A2(new_n11994_), .B(new_n16743_), .ZN(new_n16829_));
  NAND2_X1   g13884(.A1(new_n16829_), .A2(pi1158), .ZN(new_n16830_));
  NAND4_X1   g13885(.A1(new_n16826_), .A2(new_n11989_), .A3(new_n16828_), .A4(new_n16830_), .ZN(new_n16831_));
  NAND2_X1   g13886(.A1(new_n14732_), .A2(new_n11999_), .ZN(new_n16832_));
  AOI21_X1   g13887(.A1(new_n16831_), .A2(new_n11986_), .B(new_n16832_), .ZN(new_n16833_));
  OAI21_X1   g13888(.A1(new_n16813_), .A2(new_n16821_), .B(new_n16833_), .ZN(new_n16834_));
  NAND2_X1   g13889(.A1(new_n16834_), .A2(new_n16777_), .ZN(new_n16835_));
  AOI22_X1   g13890(.A1(new_n16835_), .A2(new_n14726_), .B1(new_n16768_), .B2(new_n16769_), .ZN(new_n16836_));
  NOR3_X1    g13891(.A1(new_n16836_), .A2(pi0644), .A3(new_n16754_), .ZN(new_n16837_));
  AOI21_X1   g13892(.A1(new_n16836_), .A2(new_n12082_), .B(new_n16753_), .ZN(new_n16838_));
  INV_X1     g13893(.I(new_n16761_), .ZN(new_n16839_));
  NOR2_X1    g13894(.A1(new_n12053_), .A2(new_n12091_), .ZN(new_n16840_));
  INV_X1     g13895(.I(new_n16840_), .ZN(new_n16841_));
  NOR4_X1    g13896(.A1(new_n16839_), .A2(new_n14740_), .A3(new_n16737_), .A4(new_n16841_), .ZN(new_n16842_));
  NOR4_X1    g13897(.A1(new_n16837_), .A2(new_n16838_), .A3(new_n13169_), .A4(new_n16842_), .ZN(new_n16843_));
  NOR3_X1    g13898(.A1(new_n16839_), .A2(new_n12082_), .A3(new_n16841_), .ZN(new_n16844_));
  NOR3_X1    g13899(.A1(new_n16844_), .A2(pi0715), .A3(new_n16737_), .ZN(new_n16845_));
  OAI21_X1   g13900(.A1(new_n16845_), .A2(pi1160), .B(pi0790), .ZN(new_n16846_));
  AND2_X2    g13901(.A1(new_n16836_), .A2(new_n14747_), .Z(new_n16847_));
  OAI21_X1   g13902(.A1(new_n16843_), .A2(new_n16846_), .B(new_n16847_), .ZN(new_n16848_));
  NOR2_X1    g13903(.A1(new_n11875_), .A2(new_n15660_), .ZN(new_n16849_));
  INV_X1     g13904(.I(new_n16849_), .ZN(new_n16850_));
  NOR3_X1    g13905(.A1(new_n13368_), .A2(pi0174), .A3(new_n16850_), .ZN(new_n16851_));
  AOI21_X1   g13906(.A1(new_n12828_), .A2(new_n16850_), .B(new_n7151_), .ZN(new_n16852_));
  OAI21_X1   g13907(.A1(new_n16851_), .A2(new_n16852_), .B(pi0038), .ZN(new_n16853_));
  NAND2_X1   g13908(.A1(new_n7151_), .A2(pi0759), .ZN(new_n16854_));
  OAI21_X1   g13909(.A1(new_n14759_), .A2(new_n15660_), .B(pi0039), .ZN(new_n16855_));
  NOR2_X1    g13910(.A1(new_n15679_), .A2(new_n16855_), .ZN(new_n16856_));
  OAI21_X1   g13911(.A1(pi0759), .A2(new_n12852_), .B(new_n13346_), .ZN(new_n16857_));
  NAND3_X1   g13912(.A1(new_n12664_), .A2(new_n15660_), .A3(new_n12852_), .ZN(new_n16858_));
  NAND3_X1   g13913(.A1(new_n16857_), .A2(new_n16858_), .A3(new_n3154_), .ZN(new_n16859_));
  NOR2_X1    g13914(.A1(new_n16856_), .A2(new_n16859_), .ZN(new_n16860_));
  OAI22_X1   g13915(.A1(new_n16860_), .A2(new_n7151_), .B1(new_n12694_), .B2(new_n16854_), .ZN(new_n16861_));
  NAND2_X1   g13916(.A1(new_n16861_), .A2(new_n3172_), .ZN(new_n16862_));
  NAND2_X1   g13917(.A1(new_n16862_), .A2(new_n16853_), .ZN(new_n16863_));
  NAND2_X1   g13918(.A1(new_n12277_), .A2(new_n7151_), .ZN(new_n16864_));
  NOR4_X1    g13919(.A1(new_n12349_), .A2(pi0039), .A3(pi0174), .A4(pi0759), .ZN(new_n16865_));
  NAND2_X1   g13920(.A1(pi0174), .A2(pi0759), .ZN(new_n16866_));
  AOI21_X1   g13921(.A1(new_n16864_), .A2(new_n16865_), .B(new_n16866_), .ZN(new_n16867_));
  NAND2_X1   g13922(.A1(new_n16867_), .A2(new_n13332_), .ZN(new_n16868_));
  AOI21_X1   g13923(.A1(new_n13362_), .A2(pi0174), .B(pi0759), .ZN(new_n16869_));
  OAI21_X1   g13924(.A1(pi0174), .A2(new_n13360_), .B(new_n16869_), .ZN(new_n16870_));
  NOR4_X1    g13925(.A1(new_n12668_), .A2(new_n7151_), .A3(pi0759), .A4(new_n13347_), .ZN(new_n16871_));
  NOR2_X1    g13926(.A1(new_n16871_), .A2(pi0039), .ZN(new_n16872_));
  NAND3_X1   g13927(.A1(new_n16853_), .A2(pi0696), .A3(new_n14352_), .ZN(new_n16873_));
  NAND2_X1   g13928(.A1(new_n16873_), .A2(new_n14778_), .ZN(new_n16874_));
  AOI21_X1   g13929(.A1(new_n16870_), .A2(new_n16872_), .B(new_n16874_), .ZN(new_n16875_));
  AOI21_X1   g13930(.A1(new_n16875_), .A2(new_n16868_), .B(pi0696), .ZN(new_n16876_));
  AOI22_X1   g13931(.A1(new_n16863_), .A2(new_n16876_), .B1(pi0174), .B2(new_n3232_), .ZN(new_n16877_));
  INV_X1     g13932(.I(new_n16877_), .ZN(new_n16878_));
  NOR2_X1    g13933(.A1(new_n3231_), .A2(pi0174), .ZN(new_n16879_));
  AOI21_X1   g13934(.A1(new_n16863_), .A2(new_n3231_), .B(new_n16879_), .ZN(new_n16880_));
  AOI21_X1   g13935(.A1(new_n16880_), .A2(new_n12970_), .B(pi1153), .ZN(new_n16881_));
  OAI21_X1   g13936(.A1(new_n12970_), .A2(new_n16878_), .B(new_n16881_), .ZN(new_n16882_));
  NAND3_X1   g13937(.A1(new_n14382_), .A2(new_n7151_), .A3(new_n13395_), .ZN(new_n16883_));
  OAI21_X1   g13938(.A1(pi0174), .A2(new_n13395_), .B(new_n13399_), .ZN(new_n16884_));
  NOR3_X1    g13939(.A1(new_n3232_), .A2(pi0038), .A3(new_n15674_), .ZN(new_n16887_));
  AND3_X2    g13940(.A1(new_n16883_), .A2(new_n16884_), .A3(new_n16887_), .Z(new_n16888_));
  AOI22_X1   g13941(.A1(new_n14396_), .A2(pi0174), .B1(pi0696), .B2(new_n3231_), .ZN(new_n16889_));
  NOR2_X1    g13942(.A1(new_n16888_), .A2(new_n16889_), .ZN(new_n16890_));
  INV_X1     g13943(.I(new_n16890_), .ZN(new_n16891_));
  NOR2_X1    g13944(.A1(new_n12965_), .A2(new_n7151_), .ZN(new_n16892_));
  INV_X1     g13945(.I(new_n16892_), .ZN(new_n16893_));
  NAND2_X1   g13946(.A1(new_n16893_), .A2(pi0625), .ZN(new_n16894_));
  NAND2_X1   g13947(.A1(new_n16894_), .A2(new_n11893_), .ZN(new_n16895_));
  AOI21_X1   g13948(.A1(new_n16891_), .A2(new_n12970_), .B(new_n16895_), .ZN(new_n16896_));
  NOR2_X1    g13949(.A1(new_n16896_), .A2(new_n13657_), .ZN(new_n16897_));
  NAND2_X1   g13950(.A1(new_n16882_), .A2(new_n16897_), .ZN(new_n16898_));
  NAND2_X1   g13951(.A1(new_n16890_), .A2(pi0625), .ZN(new_n16899_));
  AOI21_X1   g13952(.A1(new_n16899_), .A2(new_n16894_), .B(new_n11893_), .ZN(new_n16900_));
  INV_X1     g13953(.I(new_n16900_), .ZN(new_n16901_));
  OAI21_X1   g13954(.A1(new_n16880_), .A2(new_n12970_), .B(new_n12977_), .ZN(new_n16902_));
  AOI21_X1   g13955(.A1(pi0625), .A2(new_n16877_), .B(new_n16902_), .ZN(new_n16903_));
  NAND2_X1   g13956(.A1(new_n16903_), .A2(new_n16901_), .ZN(new_n16904_));
  NAND2_X1   g13957(.A1(new_n16904_), .A2(new_n16898_), .ZN(new_n16905_));
  MUX2_X1    g13958(.I0(new_n16905_), .I1(new_n16878_), .S(new_n11891_), .Z(new_n16906_));
  NOR2_X1    g13959(.A1(new_n16906_), .A2(pi0785), .ZN(new_n16907_));
  INV_X1     g13960(.I(new_n16907_), .ZN(new_n16908_));
  NOR2_X1    g13961(.A1(new_n16896_), .A2(new_n16900_), .ZN(new_n16909_));
  MUX2_X1    g13962(.I0(new_n16909_), .I1(new_n16891_), .S(new_n11891_), .Z(new_n16910_));
  OAI21_X1   g13963(.A1(new_n16910_), .A2(pi0609), .B(pi1155), .ZN(new_n16911_));
  NOR2_X1    g13964(.A1(new_n16893_), .A2(new_n11924_), .ZN(new_n16912_));
  AOI21_X1   g13965(.A1(new_n16880_), .A2(new_n11924_), .B(new_n16912_), .ZN(new_n16913_));
  NAND3_X1   g13966(.A1(new_n16913_), .A2(pi0609), .A3(new_n16892_), .ZN(new_n16914_));
  INV_X1     g13967(.I(new_n16914_), .ZN(new_n16915_));
  AOI21_X1   g13968(.A1(pi0609), .A2(new_n16893_), .B(new_n16913_), .ZN(new_n16916_));
  OAI21_X1   g13969(.A1(new_n16915_), .A2(new_n16916_), .B(new_n11912_), .ZN(new_n16917_));
  NAND2_X1   g13970(.A1(new_n16917_), .A2(pi0660), .ZN(new_n16918_));
  NAND2_X1   g13971(.A1(new_n16918_), .A2(pi0609), .ZN(new_n16919_));
  NOR2_X1    g13972(.A1(new_n16906_), .A2(new_n16919_), .ZN(new_n16920_));
  AOI22_X1   g13973(.A1(new_n16903_), .A2(new_n16901_), .B1(new_n16882_), .B2(new_n16897_), .ZN(new_n16921_));
  MUX2_X1    g13974(.I0(new_n16921_), .I1(new_n16877_), .S(new_n11891_), .Z(new_n16922_));
  NOR3_X1    g13975(.A1(new_n16913_), .A2(new_n11903_), .A3(new_n16892_), .ZN(new_n16923_));
  AOI21_X1   g13976(.A1(new_n16913_), .A2(pi0609), .B(new_n16893_), .ZN(new_n16924_));
  NOR2_X1    g13977(.A1(new_n11923_), .A2(pi1155), .ZN(new_n16925_));
  OAI21_X1   g13978(.A1(new_n16910_), .A2(new_n11903_), .B(new_n16925_), .ZN(new_n16926_));
  AOI21_X1   g13979(.A1(new_n16922_), .A2(new_n11903_), .B(new_n16926_), .ZN(new_n16927_));
  AOI21_X1   g13980(.A1(new_n16920_), .A2(new_n16911_), .B(new_n16927_), .ZN(new_n16928_));
  NOR3_X1    g13981(.A1(new_n16928_), .A2(new_n11870_), .A3(new_n16908_), .ZN(new_n16929_));
  NAND4_X1   g13982(.A1(new_n16922_), .A2(pi0609), .A3(new_n16911_), .A4(new_n16918_), .ZN(new_n16930_));
  NOR2_X1    g13983(.A1(new_n16906_), .A2(pi0609), .ZN(new_n16931_));
  OAI21_X1   g13984(.A1(new_n16931_), .A2(new_n16926_), .B(new_n16930_), .ZN(new_n16932_));
  AOI21_X1   g13985(.A1(new_n16932_), .A2(pi0785), .B(new_n16907_), .ZN(new_n16933_));
  NOR3_X1    g13986(.A1(new_n16933_), .A2(new_n16929_), .A3(pi0781), .ZN(new_n16934_));
  INV_X1     g13987(.I(new_n16934_), .ZN(new_n16935_));
  INV_X1     g13988(.I(new_n16913_), .ZN(new_n16936_));
  OAI21_X1   g13989(.A1(new_n16923_), .A2(new_n16924_), .B(pi1155), .ZN(new_n16937_));
  NAND2_X1   g13990(.A1(new_n16917_), .A2(new_n16937_), .ZN(new_n16938_));
  MUX2_X1    g13991(.I0(new_n16938_), .I1(new_n16936_), .S(new_n11870_), .Z(new_n16939_));
  NAND3_X1   g13992(.A1(new_n16939_), .A2(new_n11934_), .A3(new_n16892_), .ZN(new_n16940_));
  OAI21_X1   g13993(.A1(new_n16939_), .A2(pi0618), .B(new_n16893_), .ZN(new_n16941_));
  NAND3_X1   g13994(.A1(new_n16941_), .A2(new_n16940_), .A3(new_n11950_), .ZN(new_n16942_));
  NOR2_X1    g13995(.A1(new_n16942_), .A2(new_n11949_), .ZN(new_n16943_));
  INV_X1     g13996(.I(new_n16943_), .ZN(new_n16944_));
  NOR2_X1    g13997(.A1(new_n16893_), .A2(new_n11938_), .ZN(new_n16945_));
  AOI21_X1   g13998(.A1(new_n16910_), .A2(new_n11938_), .B(new_n16945_), .ZN(new_n16946_));
  NOR4_X1    g13999(.A1(new_n16933_), .A2(new_n16929_), .A3(new_n11934_), .A4(pi1154), .ZN(new_n16947_));
  NAND3_X1   g14000(.A1(new_n16932_), .A2(pi0785), .A3(new_n16907_), .ZN(new_n16948_));
  OAI21_X1   g14001(.A1(new_n16928_), .A2(new_n11870_), .B(new_n16908_), .ZN(new_n16949_));
  NAND3_X1   g14002(.A1(new_n16948_), .A2(new_n16949_), .A3(new_n11934_), .ZN(new_n16950_));
  AOI21_X1   g14003(.A1(new_n16946_), .A2(pi0618), .B(new_n14687_), .ZN(new_n16951_));
  AOI22_X1   g14004(.A1(new_n16947_), .A2(new_n16944_), .B1(new_n16950_), .B2(new_n16951_), .ZN(new_n16952_));
  NOR3_X1    g14005(.A1(new_n16952_), .A2(new_n11969_), .A3(new_n16935_), .ZN(new_n16953_));
  NAND4_X1   g14006(.A1(new_n16948_), .A2(new_n16949_), .A3(pi0618), .A4(new_n11950_), .ZN(new_n16954_));
  NOR3_X1    g14007(.A1(new_n16933_), .A2(new_n16929_), .A3(pi0618), .ZN(new_n16955_));
  INV_X1     g14008(.I(new_n16951_), .ZN(new_n16956_));
  OAI22_X1   g14009(.A1(new_n16943_), .A2(new_n16954_), .B1(new_n16955_), .B2(new_n16956_), .ZN(new_n16957_));
  AOI21_X1   g14010(.A1(new_n16957_), .A2(pi0781), .B(new_n16934_), .ZN(new_n16958_));
  NOR3_X1    g14011(.A1(new_n16958_), .A2(new_n16953_), .A3(pi0789), .ZN(new_n16959_));
  INV_X1     g14012(.I(new_n16959_), .ZN(new_n16960_));
  INV_X1     g14013(.I(new_n16916_), .ZN(new_n16961_));
  AOI21_X1   g14014(.A1(new_n16961_), .A2(new_n16914_), .B(pi1155), .ZN(new_n16962_));
  INV_X1     g14015(.I(new_n16937_), .ZN(new_n16963_));
  NOR2_X1    g14016(.A1(new_n16962_), .A2(new_n16963_), .ZN(new_n16964_));
  MUX2_X1    g14017(.I0(new_n16964_), .I1(new_n16913_), .S(new_n11870_), .Z(new_n16965_));
  MUX2_X1    g14018(.I0(new_n16942_), .I1(new_n16965_), .S(new_n11969_), .Z(new_n16966_));
  NOR3_X1    g14019(.A1(new_n16966_), .A2(pi0619), .A3(new_n16893_), .ZN(new_n16967_));
  AOI21_X1   g14020(.A1(new_n16966_), .A2(new_n11967_), .B(new_n16892_), .ZN(new_n16968_));
  NOR3_X1    g14021(.A1(new_n16967_), .A2(new_n16968_), .A3(pi1159), .ZN(new_n16969_));
  NAND2_X1   g14022(.A1(new_n16969_), .A2(pi0648), .ZN(new_n16970_));
  NOR2_X1    g14023(.A1(new_n16892_), .A2(new_n11961_), .ZN(new_n16971_));
  AOI21_X1   g14024(.A1(new_n16946_), .A2(new_n11961_), .B(new_n16971_), .ZN(new_n16972_));
  NOR4_X1    g14025(.A1(new_n16958_), .A2(new_n16953_), .A3(new_n11967_), .A4(pi1159), .ZN(new_n16973_));
  NAND3_X1   g14026(.A1(new_n16957_), .A2(pi0781), .A3(new_n16934_), .ZN(new_n16974_));
  OAI21_X1   g14027(.A1(new_n16952_), .A2(new_n11969_), .B(new_n16935_), .ZN(new_n16975_));
  NAND3_X1   g14028(.A1(new_n16974_), .A2(new_n16975_), .A3(new_n11967_), .ZN(new_n16976_));
  INV_X1     g14029(.I(new_n16972_), .ZN(new_n16977_));
  AOI21_X1   g14030(.A1(new_n16977_), .A2(pi0619), .B(new_n14904_), .ZN(new_n16978_));
  AOI22_X1   g14031(.A1(new_n16973_), .A2(new_n16970_), .B1(new_n16976_), .B2(new_n16978_), .ZN(new_n16979_));
  NOR3_X1    g14032(.A1(new_n16979_), .A2(new_n11985_), .A3(new_n16960_), .ZN(new_n16980_));
  INV_X1     g14033(.I(new_n16970_), .ZN(new_n16981_));
  NAND4_X1   g14034(.A1(new_n16974_), .A2(new_n16975_), .A3(pi0619), .A4(new_n11869_), .ZN(new_n16982_));
  NOR3_X1    g14035(.A1(new_n16958_), .A2(new_n16953_), .A3(pi0619), .ZN(new_n16983_));
  INV_X1     g14036(.I(new_n16978_), .ZN(new_n16984_));
  OAI22_X1   g14037(.A1(new_n16981_), .A2(new_n16982_), .B1(new_n16983_), .B2(new_n16984_), .ZN(new_n16985_));
  AOI21_X1   g14038(.A1(new_n16985_), .A2(pi0789), .B(new_n16959_), .ZN(new_n16986_));
  NOR2_X1    g14039(.A1(new_n16986_), .A2(new_n16980_), .ZN(new_n16987_));
  AND3_X2    g14040(.A1(new_n16941_), .A2(new_n16940_), .A3(new_n11950_), .Z(new_n16988_));
  MUX2_X1    g14041(.I0(new_n16988_), .I1(new_n16939_), .S(new_n11969_), .Z(new_n16989_));
  MUX2_X1    g14042(.I0(new_n16969_), .I1(new_n16989_), .S(new_n11985_), .Z(new_n16990_));
  NOR3_X1    g14043(.A1(new_n11994_), .A2(new_n11989_), .A3(pi1158), .ZN(new_n16991_));
  INV_X1     g14044(.I(new_n16991_), .ZN(new_n16992_));
  NOR2_X1    g14045(.A1(new_n16893_), .A2(new_n12014_), .ZN(new_n16993_));
  AOI21_X1   g14046(.A1(new_n16972_), .A2(new_n12014_), .B(new_n16993_), .ZN(new_n16994_));
  NOR2_X1    g14047(.A1(new_n11994_), .A2(pi0641), .ZN(new_n16995_));
  OAI21_X1   g14048(.A1(new_n16990_), .A2(new_n16992_), .B(new_n16995_), .ZN(new_n16996_));
  INV_X1     g14049(.I(new_n16996_), .ZN(new_n16997_));
  OR3_X2     g14050(.A1(new_n16967_), .A2(new_n16968_), .A3(pi1159), .Z(new_n16998_));
  NOR2_X1    g14051(.A1(new_n16989_), .A2(pi0789), .ZN(new_n16999_));
  NAND3_X1   g14052(.A1(new_n16998_), .A2(pi0789), .A3(new_n16999_), .ZN(new_n17000_));
  INV_X1     g14053(.I(new_n16999_), .ZN(new_n17001_));
  OAI21_X1   g14054(.A1(new_n16969_), .A2(new_n11985_), .B(new_n17001_), .ZN(new_n17002_));
  NAND3_X1   g14055(.A1(new_n17000_), .A2(new_n11994_), .A3(new_n17002_), .ZN(new_n17003_));
  AOI21_X1   g14056(.A1(new_n16892_), .A2(pi0626), .B(new_n11989_), .ZN(new_n17004_));
  NOR3_X1    g14057(.A1(new_n11989_), .A2(pi0626), .A3(pi1158), .ZN(new_n17005_));
  INV_X1     g14058(.I(new_n17005_), .ZN(new_n17006_));
  AOI21_X1   g14059(.A1(new_n17003_), .A2(new_n17004_), .B(new_n17006_), .ZN(new_n17007_));
  OAI22_X1   g14060(.A1(new_n16986_), .A2(new_n16980_), .B1(new_n17007_), .B2(new_n16997_), .ZN(new_n17008_));
  MUX2_X1    g14061(.I0(new_n17008_), .I1(new_n16987_), .S(new_n11986_), .Z(new_n17009_));
  NAND3_X1   g14062(.A1(new_n16985_), .A2(pi0789), .A3(new_n16959_), .ZN(new_n17010_));
  OAI21_X1   g14063(.A1(new_n16979_), .A2(new_n11985_), .B(new_n16960_), .ZN(new_n17011_));
  NAND2_X1   g14064(.A1(new_n17010_), .A2(new_n17011_), .ZN(new_n17012_));
  NOR3_X1    g14065(.A1(new_n17008_), .A2(new_n11986_), .A3(new_n17012_), .ZN(new_n17013_));
  AOI21_X1   g14066(.A1(new_n17008_), .A2(pi0788), .B(new_n16987_), .ZN(new_n17014_));
  NAND2_X1   g14067(.A1(new_n16990_), .A2(new_n14624_), .ZN(new_n17015_));
  NAND2_X1   g14068(.A1(new_n16893_), .A2(new_n11997_), .ZN(new_n17016_));
  AOI21_X1   g14069(.A1(new_n17015_), .A2(new_n17016_), .B(pi0628), .ZN(new_n17017_));
  NOR2_X1    g14070(.A1(new_n16892_), .A2(new_n13114_), .ZN(new_n17018_));
  AOI21_X1   g14071(.A1(new_n16994_), .A2(new_n13114_), .B(new_n17018_), .ZN(new_n17019_));
  INV_X1     g14072(.I(new_n17019_), .ZN(new_n17020_));
  NAND3_X1   g14073(.A1(new_n17020_), .A2(new_n12031_), .A3(new_n16892_), .ZN(new_n17021_));
  OAI21_X1   g14074(.A1(new_n17020_), .A2(pi0628), .B(new_n16893_), .ZN(new_n17022_));
  NAND3_X1   g14075(.A1(new_n17022_), .A2(new_n17021_), .A3(new_n12026_), .ZN(new_n17023_));
  INV_X1     g14076(.I(new_n17023_), .ZN(new_n17024_));
  AOI21_X1   g14077(.A1(new_n17024_), .A2(pi0629), .B(new_n12031_), .ZN(new_n17025_));
  OAI21_X1   g14078(.A1(new_n17017_), .A2(new_n12026_), .B(new_n17025_), .ZN(new_n17026_));
  INV_X1     g14079(.I(new_n17026_), .ZN(new_n17027_));
  AND2_X2    g14080(.A1(new_n17015_), .A2(new_n17016_), .Z(new_n17028_));
  NOR3_X1    g14081(.A1(new_n12030_), .A2(new_n12026_), .A3(pi0628), .ZN(new_n17029_));
  OAI22_X1   g14082(.A1(new_n17013_), .A2(new_n17014_), .B1(new_n17027_), .B2(new_n17029_), .ZN(new_n17030_));
  MUX2_X1    g14083(.I0(new_n17030_), .I1(new_n17009_), .S(new_n11868_), .Z(new_n17031_));
  INV_X1     g14084(.I(new_n17031_), .ZN(new_n17032_));
  NAND2_X1   g14085(.A1(new_n16893_), .A2(new_n12053_), .ZN(new_n17033_));
  OAI21_X1   g14086(.A1(new_n17028_), .A2(new_n12053_), .B(new_n17033_), .ZN(new_n17034_));
  AOI21_X1   g14087(.A1(new_n17034_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n17035_));
  MUX2_X1    g14088(.I0(new_n17024_), .I1(new_n17020_), .S(new_n11868_), .Z(new_n17036_));
  NAND3_X1   g14089(.A1(new_n17036_), .A2(new_n12061_), .A3(new_n16892_), .ZN(new_n17037_));
  OAI21_X1   g14090(.A1(new_n17036_), .A2(pi0647), .B(new_n16893_), .ZN(new_n17038_));
  NAND3_X1   g14091(.A1(new_n17038_), .A2(new_n17037_), .A3(new_n12049_), .ZN(new_n17039_));
  NOR2_X1    g14092(.A1(new_n17039_), .A2(new_n12060_), .ZN(new_n17040_));
  NOR3_X1    g14093(.A1(new_n17035_), .A2(new_n12061_), .A3(new_n17040_), .ZN(new_n17041_));
  AOI21_X1   g14094(.A1(new_n17010_), .A2(new_n17011_), .B(new_n16996_), .ZN(new_n17042_));
  NAND3_X1   g14095(.A1(new_n17042_), .A2(new_n16987_), .A3(pi0788), .ZN(new_n17043_));
  OAI21_X1   g14096(.A1(new_n16990_), .A2(pi0626), .B(new_n17004_), .ZN(new_n17044_));
  NAND2_X1   g14097(.A1(new_n17044_), .A2(new_n17005_), .ZN(new_n17045_));
  AOI22_X1   g14098(.A1(new_n17010_), .A2(new_n17011_), .B1(new_n17045_), .B2(new_n16996_), .ZN(new_n17046_));
  OAI21_X1   g14099(.A1(new_n17046_), .A2(new_n11986_), .B(new_n17012_), .ZN(new_n17047_));
  AOI21_X1   g14100(.A1(new_n17047_), .A2(new_n17043_), .B(new_n17026_), .ZN(new_n17048_));
  NAND3_X1   g14101(.A1(new_n17048_), .A2(pi0792), .A3(new_n17009_), .ZN(new_n17049_));
  NAND2_X1   g14102(.A1(new_n17047_), .A2(new_n17043_), .ZN(new_n17050_));
  INV_X1     g14103(.I(new_n17029_), .ZN(new_n17051_));
  AOI22_X1   g14104(.A1(new_n17047_), .A2(new_n17043_), .B1(new_n17026_), .B2(new_n17051_), .ZN(new_n17052_));
  OAI21_X1   g14105(.A1(new_n17052_), .A2(new_n11868_), .B(new_n17050_), .ZN(new_n17053_));
  NAND3_X1   g14106(.A1(new_n17053_), .A2(new_n17049_), .A3(new_n12061_), .ZN(new_n17054_));
  AOI21_X1   g14107(.A1(new_n17034_), .A2(pi0647), .B(new_n13743_), .ZN(new_n17055_));
  AOI22_X1   g14108(.A1(new_n17054_), .A2(new_n17055_), .B1(new_n17031_), .B2(new_n17041_), .ZN(new_n17056_));
  MUX2_X1    g14109(.I0(new_n17056_), .I1(new_n17032_), .S(new_n12048_), .Z(new_n17057_));
  NOR2_X1    g14110(.A1(new_n17034_), .A2(new_n12091_), .ZN(new_n17058_));
  AOI21_X1   g14111(.A1(new_n12091_), .A2(new_n16892_), .B(new_n17058_), .ZN(new_n17059_));
  NAND2_X1   g14112(.A1(new_n17059_), .A2(new_n12082_), .ZN(new_n17060_));
  AOI21_X1   g14113(.A1(new_n16893_), .A2(pi0644), .B(new_n12099_), .ZN(new_n17061_));
  NOR2_X1    g14114(.A1(new_n17036_), .A2(pi0787), .ZN(new_n17062_));
  NAND2_X1   g14115(.A1(new_n17039_), .A2(pi0787), .ZN(new_n17063_));
  XNOR2_X1   g14116(.A1(new_n17063_), .A2(new_n17062_), .ZN(new_n17064_));
  OAI21_X1   g14117(.A1(new_n17064_), .A2(new_n12082_), .B(new_n13168_), .ZN(new_n17065_));
  AOI21_X1   g14118(.A1(new_n17060_), .A2(new_n17061_), .B(new_n17065_), .ZN(new_n17066_));
  OAI21_X1   g14119(.A1(new_n17057_), .A2(pi0644), .B(new_n17066_), .ZN(new_n17067_));
  NAND2_X1   g14120(.A1(new_n17031_), .A2(new_n12048_), .ZN(new_n17068_));
  OR3_X2     g14121(.A1(new_n17056_), .A2(new_n12048_), .A3(new_n17068_), .Z(new_n17069_));
  OAI21_X1   g14122(.A1(new_n17056_), .A2(new_n12048_), .B(new_n17068_), .ZN(new_n17070_));
  NOR3_X1    g14123(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n17071_));
  NAND2_X1   g14124(.A1(new_n17059_), .A2(new_n17071_), .ZN(new_n17072_));
  NOR2_X1    g14125(.A1(new_n12082_), .A2(pi0715), .ZN(new_n17073_));
  NAND4_X1   g14126(.A1(new_n17069_), .A2(new_n17070_), .A3(new_n17072_), .A4(new_n17073_), .ZN(new_n17074_));
  OAI21_X1   g14127(.A1(new_n17057_), .A2(new_n5223_), .B(new_n11867_), .ZN(new_n17075_));
  AOI21_X1   g14128(.A1(new_n17067_), .A2(new_n17074_), .B(new_n17075_), .ZN(new_n17076_));
  NAND2_X1   g14129(.A1(pi0057), .A2(pi0174), .ZN(new_n17077_));
  AOI21_X1   g14130(.A1(new_n17077_), .A2(new_n13184_), .B(pi0057), .ZN(new_n17078_));
  OAI21_X1   g14131(.A1(new_n5224_), .A2(pi0174), .B(new_n17078_), .ZN(new_n17079_));
  OAI21_X1   g14132(.A1(new_n17076_), .A2(new_n17079_), .B(new_n16848_), .ZN(po0331));
  NOR2_X1    g14133(.A1(new_n2925_), .A2(pi0175), .ZN(new_n17081_));
  NOR2_X1    g14134(.A1(new_n11877_), .A2(new_n15707_), .ZN(new_n17082_));
  NOR2_X1    g14135(.A1(new_n17082_), .A2(new_n17081_), .ZN(new_n17083_));
  AOI21_X1   g14136(.A1(new_n11886_), .A2(pi0700), .B(new_n17081_), .ZN(new_n17084_));
  NOR2_X1    g14137(.A1(new_n17084_), .A2(new_n11874_), .ZN(new_n17085_));
  INV_X1     g14138(.I(new_n17085_), .ZN(new_n17086_));
  NAND2_X1   g14139(.A1(new_n17086_), .A2(new_n17083_), .ZN(new_n17087_));
  NAND2_X1   g14140(.A1(new_n17087_), .A2(new_n11891_), .ZN(new_n17088_));
  NOR2_X1    g14141(.A1(new_n17086_), .A2(new_n12970_), .ZN(new_n17089_));
  NOR4_X1    g14142(.A1(new_n17089_), .A2(new_n11893_), .A3(new_n17081_), .A4(new_n17082_), .ZN(new_n17090_));
  NOR2_X1    g14143(.A1(new_n13201_), .A2(new_n15745_), .ZN(new_n17091_));
  NOR2_X1    g14144(.A1(new_n17081_), .A2(pi1153), .ZN(new_n17092_));
  INV_X1     g14145(.I(new_n17092_), .ZN(new_n17093_));
  NOR2_X1    g14146(.A1(new_n17091_), .A2(new_n17093_), .ZN(new_n17094_));
  INV_X1     g14147(.I(new_n17094_), .ZN(new_n17095_));
  NAND2_X1   g14148(.A1(new_n17095_), .A2(pi0608), .ZN(new_n17096_));
  INV_X1     g14149(.I(new_n17089_), .ZN(new_n17097_));
  AOI21_X1   g14150(.A1(new_n17097_), .A2(new_n17087_), .B(new_n17093_), .ZN(new_n17098_));
  OAI21_X1   g14151(.A1(new_n17091_), .A2(new_n17084_), .B(pi1153), .ZN(new_n17099_));
  NAND2_X1   g14152(.A1(new_n17099_), .A2(new_n13657_), .ZN(new_n17100_));
  OAI22_X1   g14153(.A1(new_n17096_), .A2(new_n17090_), .B1(new_n17098_), .B2(new_n17100_), .ZN(new_n17101_));
  NAND2_X1   g14154(.A1(new_n17101_), .A2(pi0778), .ZN(new_n17102_));
  XOR2_X1    g14155(.A1(new_n17102_), .A2(new_n17088_), .Z(new_n17103_));
  INV_X1     g14156(.I(new_n17103_), .ZN(new_n17104_));
  NAND2_X1   g14157(.A1(new_n17095_), .A2(new_n17099_), .ZN(new_n17105_));
  MUX2_X1    g14158(.I0(new_n17105_), .I1(new_n17084_), .S(new_n11891_), .Z(new_n17106_));
  XNOR2_X1   g14159(.A1(new_n17103_), .A2(new_n17106_), .ZN(new_n17107_));
  NAND2_X1   g14160(.A1(new_n17107_), .A2(pi0609), .ZN(new_n17108_));
  XOR2_X1    g14161(.A1(new_n17108_), .A2(new_n17104_), .Z(new_n17109_));
  INV_X1     g14162(.I(new_n17082_), .ZN(new_n17110_));
  NOR2_X1    g14163(.A1(new_n17083_), .A2(new_n11925_), .ZN(new_n17111_));
  NOR4_X1    g14164(.A1(new_n17111_), .A2(pi1155), .A3(new_n12997_), .A4(new_n17110_), .ZN(new_n17112_));
  NOR2_X1    g14165(.A1(new_n17112_), .A2(pi0660), .ZN(new_n17113_));
  OAI21_X1   g14166(.A1(new_n17109_), .A2(pi1155), .B(new_n17113_), .ZN(new_n17114_));
  NOR2_X1    g14167(.A1(new_n17110_), .A2(new_n12997_), .ZN(new_n17115_));
  NOR4_X1    g14168(.A1(new_n17115_), .A2(new_n11923_), .A3(pi1155), .A4(new_n17081_), .ZN(new_n17117_));
  NOR2_X1    g14169(.A1(new_n17117_), .A2(new_n11870_), .ZN(new_n17118_));
  AOI22_X1   g14170(.A1(new_n17114_), .A2(new_n17118_), .B1(new_n11870_), .B2(new_n17104_), .ZN(new_n17119_));
  NOR2_X1    g14171(.A1(new_n17119_), .A2(pi0781), .ZN(new_n17120_));
  NOR4_X1    g14172(.A1(new_n17106_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n17121_));
  NOR2_X1    g14173(.A1(new_n17111_), .A2(pi0785), .ZN(new_n17122_));
  NOR4_X1    g14174(.A1(new_n17112_), .A2(pi1155), .A3(new_n17081_), .A4(new_n17115_), .ZN(new_n17123_));
  NOR2_X1    g14175(.A1(new_n17123_), .A2(new_n11870_), .ZN(new_n17124_));
  XOR2_X1    g14176(.A1(new_n17124_), .A2(new_n17122_), .Z(new_n17125_));
  INV_X1     g14177(.I(new_n17125_), .ZN(new_n17126_));
  OAI21_X1   g14178(.A1(new_n17126_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n17127_));
  OAI21_X1   g14179(.A1(new_n17126_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n17128_));
  NOR2_X1    g14180(.A1(new_n17106_), .A2(new_n11939_), .ZN(new_n17129_));
  NOR4_X1    g14181(.A1(new_n17119_), .A2(new_n11934_), .A3(pi1154), .A4(new_n17129_), .ZN(new_n17130_));
  NOR2_X1    g14182(.A1(new_n17130_), .A2(new_n17128_), .ZN(new_n17131_));
  OAI22_X1   g14183(.A1(new_n17131_), .A2(pi0627), .B1(new_n17121_), .B2(new_n17127_), .ZN(new_n17132_));
  AOI21_X1   g14184(.A1(new_n17132_), .A2(pi0781), .B(new_n17120_), .ZN(new_n17133_));
  INV_X1     g14185(.I(new_n17129_), .ZN(new_n17134_));
  NOR2_X1    g14186(.A1(new_n17134_), .A2(new_n11962_), .ZN(new_n17135_));
  NOR4_X1    g14187(.A1(new_n17133_), .A2(new_n11967_), .A3(pi1159), .A4(new_n17135_), .ZN(new_n17136_));
  NOR2_X1    g14188(.A1(new_n17126_), .A2(pi0781), .ZN(new_n17137_));
  AOI21_X1   g14189(.A1(new_n11944_), .A2(new_n17125_), .B(new_n17128_), .ZN(new_n17138_));
  NOR2_X1    g14190(.A1(new_n17138_), .A2(new_n11969_), .ZN(new_n17139_));
  XOR2_X1    g14191(.A1(new_n17139_), .A2(new_n17137_), .Z(new_n17140_));
  AOI21_X1   g14192(.A1(new_n17140_), .A2(new_n16479_), .B(pi1159), .ZN(new_n17141_));
  INV_X1     g14193(.I(new_n17141_), .ZN(new_n17142_));
  NOR3_X1    g14194(.A1(new_n17136_), .A2(new_n11966_), .A3(new_n17142_), .ZN(new_n17143_));
  NOR4_X1    g14195(.A1(new_n17134_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n17144_));
  INV_X1     g14196(.I(new_n17140_), .ZN(new_n17145_));
  NOR2_X1    g14197(.A1(new_n17145_), .A2(new_n16482_), .ZN(new_n17146_));
  NOR3_X1    g14198(.A1(new_n17146_), .A2(pi0648), .A3(new_n17144_), .ZN(new_n17147_));
  AOI21_X1   g14199(.A1(new_n17133_), .A2(new_n11998_), .B(pi0789), .ZN(new_n17148_));
  OAI21_X1   g14200(.A1(new_n17143_), .A2(new_n17147_), .B(new_n17148_), .ZN(new_n17149_));
  INV_X1     g14201(.I(new_n12064_), .ZN(new_n17150_));
  INV_X1     g14202(.I(new_n15080_), .ZN(new_n17151_));
  NOR3_X1    g14203(.A1(new_n17134_), .A2(new_n11962_), .A3(new_n12015_), .ZN(new_n17152_));
  NOR2_X1    g14204(.A1(new_n13114_), .A2(new_n2926_), .ZN(new_n17153_));
  INV_X1     g14205(.I(new_n17153_), .ZN(new_n17154_));
  NAND2_X1   g14206(.A1(new_n17152_), .A2(new_n17154_), .ZN(new_n17155_));
  NOR2_X1    g14207(.A1(new_n14624_), .A2(new_n17081_), .ZN(new_n17156_));
  OAI21_X1   g14208(.A1(new_n16482_), .A2(new_n17145_), .B(new_n17141_), .ZN(new_n17157_));
  MUX2_X1    g14209(.I0(new_n17157_), .I1(new_n17140_), .S(new_n11985_), .Z(new_n17158_));
  AOI21_X1   g14210(.A1(new_n17158_), .A2(new_n14624_), .B(new_n17156_), .ZN(new_n17159_));
  INV_X1     g14211(.I(new_n17159_), .ZN(new_n17160_));
  OAI22_X1   g14212(.A1(new_n17160_), .A2(new_n17150_), .B1(new_n17151_), .B2(new_n17155_), .ZN(new_n17161_));
  NAND2_X1   g14213(.A1(new_n17161_), .A2(pi0629), .ZN(new_n17162_));
  INV_X1     g14214(.I(new_n15084_), .ZN(new_n17163_));
  OAI21_X1   g14215(.A1(new_n17155_), .A2(new_n17163_), .B(new_n15085_), .ZN(new_n17164_));
  AOI21_X1   g14216(.A1(new_n17159_), .A2(new_n12063_), .B(new_n17164_), .ZN(new_n17165_));
  NAND2_X1   g14217(.A1(new_n17162_), .A2(new_n17165_), .ZN(new_n17166_));
  INV_X1     g14218(.I(new_n11988_), .ZN(new_n17167_));
  INV_X1     g14219(.I(new_n17081_), .ZN(new_n17168_));
  MUX2_X1    g14220(.I0(new_n17158_), .I1(new_n17168_), .S(new_n11994_), .Z(new_n17169_));
  NOR2_X1    g14221(.A1(new_n17169_), .A2(new_n17167_), .ZN(new_n17170_));
  INV_X1     g14222(.I(new_n11990_), .ZN(new_n17171_));
  OAI21_X1   g14223(.A1(new_n17158_), .A2(new_n17081_), .B(pi0626), .ZN(new_n17172_));
  INV_X1     g14224(.I(new_n12020_), .ZN(new_n17173_));
  AOI21_X1   g14225(.A1(new_n17152_), .A2(new_n17173_), .B(pi0788), .ZN(new_n17174_));
  OAI21_X1   g14226(.A1(new_n17172_), .A2(new_n17171_), .B(new_n17174_), .ZN(new_n17175_));
  OAI21_X1   g14227(.A1(new_n17170_), .A2(new_n17175_), .B(new_n14732_), .ZN(new_n17176_));
  AOI21_X1   g14228(.A1(new_n17166_), .A2(new_n14726_), .B(new_n17176_), .ZN(new_n17177_));
  NAND3_X1   g14229(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n17081_), .ZN(new_n17178_));
  NOR2_X1    g14230(.A1(new_n17155_), .A2(new_n12068_), .ZN(new_n17179_));
  AOI21_X1   g14231(.A1(new_n17081_), .A2(pi0647), .B(pi1157), .ZN(new_n17180_));
  OAI21_X1   g14232(.A1(new_n17179_), .A2(new_n12061_), .B(new_n17180_), .ZN(new_n17181_));
  NOR2_X1    g14233(.A1(new_n17168_), .A2(pi0647), .ZN(new_n17182_));
  AOI21_X1   g14234(.A1(new_n17179_), .A2(pi0647), .B(new_n17182_), .ZN(new_n17183_));
  NAND2_X1   g14235(.A1(new_n17183_), .A2(new_n12088_), .ZN(new_n17184_));
  NAND2_X1   g14236(.A1(new_n17184_), .A2(pi0787), .ZN(new_n17185_));
  AOI21_X1   g14237(.A1(pi0630), .A2(new_n17181_), .B(new_n17185_), .ZN(new_n17186_));
  AOI22_X1   g14238(.A1(new_n17149_), .A2(new_n17177_), .B1(new_n17178_), .B2(new_n17186_), .ZN(new_n17187_));
  OR2_X2     g14239(.A1(new_n17187_), .A2(new_n12082_), .Z(new_n17188_));
  MUX2_X1    g14240(.I0(new_n17160_), .I1(new_n17168_), .S(new_n16841_), .Z(new_n17189_));
  MUX2_X1    g14241(.I0(new_n17189_), .I1(new_n17168_), .S(pi0644), .Z(new_n17190_));
  NAND2_X1   g14242(.A1(new_n17183_), .A2(pi1157), .ZN(new_n17191_));
  NOR2_X1    g14243(.A1(new_n17181_), .A2(new_n12048_), .ZN(new_n17192_));
  AOI22_X1   g14244(.A1(new_n17192_), .A2(new_n17191_), .B1(new_n12048_), .B2(new_n17179_), .ZN(new_n17193_));
  OAI21_X1   g14245(.A1(new_n17193_), .A2(new_n12082_), .B(new_n13168_), .ZN(new_n17194_));
  AOI21_X1   g14246(.A1(new_n17190_), .A2(pi0715), .B(new_n17194_), .ZN(new_n17195_));
  AOI21_X1   g14247(.A1(new_n17193_), .A2(new_n12082_), .B(pi0715), .ZN(new_n17196_));
  NAND2_X1   g14248(.A1(new_n17188_), .A2(new_n17196_), .ZN(new_n17197_));
  NAND3_X1   g14249(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n17198_));
  NOR2_X1    g14250(.A1(new_n17189_), .A2(new_n17198_), .ZN(new_n17199_));
  AOI22_X1   g14251(.A1(new_n17197_), .A2(new_n17199_), .B1(new_n17188_), .B2(new_n17195_), .ZN(new_n17200_));
  AOI21_X1   g14252(.A1(new_n17187_), .A2(new_n11867_), .B(new_n13184_), .ZN(new_n17201_));
  OAI21_X1   g14253(.A1(new_n17200_), .A2(new_n11867_), .B(new_n17201_), .ZN(new_n17202_));
  NOR2_X1    g14254(.A1(new_n12965_), .A2(pi0175), .ZN(new_n17203_));
  INV_X1     g14255(.I(new_n17203_), .ZN(new_n17204_));
  NAND2_X1   g14256(.A1(new_n17204_), .A2(new_n11997_), .ZN(new_n17205_));
  NOR2_X1    g14257(.A1(new_n15707_), .A2(pi0175), .ZN(new_n17206_));
  OAI21_X1   g14258(.A1(new_n14361_), .A2(new_n8913_), .B(pi0039), .ZN(new_n17207_));
  AOI21_X1   g14259(.A1(new_n13381_), .A2(new_n17206_), .B(new_n17207_), .ZN(new_n17208_));
  OAI21_X1   g14260(.A1(pi0766), .A2(new_n12793_), .B(new_n17208_), .ZN(new_n17209_));
  NOR2_X1    g14261(.A1(new_n12828_), .A2(pi0175), .ZN(new_n17210_));
  AOI21_X1   g14262(.A1(new_n12829_), .A2(pi0766), .B(pi0038), .ZN(new_n17211_));
  AOI21_X1   g14263(.A1(new_n17209_), .A2(new_n17211_), .B(new_n3232_), .ZN(new_n17212_));
  AOI21_X1   g14264(.A1(new_n8913_), .A2(new_n3232_), .B(new_n17212_), .ZN(new_n17213_));
  OAI21_X1   g14265(.A1(new_n17213_), .A2(new_n11914_), .B(new_n11870_), .ZN(new_n17214_));
  AOI21_X1   g14266(.A1(new_n11914_), .A2(new_n17203_), .B(new_n17214_), .ZN(new_n17215_));
  NAND2_X1   g14267(.A1(new_n17213_), .A2(new_n11924_), .ZN(new_n17216_));
  OAI22_X1   g14268(.A1(new_n17216_), .A2(pi0609), .B1(new_n12996_), .B2(new_n17203_), .ZN(new_n17217_));
  NAND2_X1   g14269(.A1(new_n17217_), .A2(new_n11912_), .ZN(new_n17218_));
  OAI22_X1   g14270(.A1(new_n17216_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n17203_), .ZN(new_n17219_));
  NAND2_X1   g14271(.A1(new_n17219_), .A2(pi1155), .ZN(new_n17220_));
  NAND2_X1   g14272(.A1(new_n17218_), .A2(new_n17220_), .ZN(new_n17221_));
  NAND2_X1   g14273(.A1(new_n17221_), .A2(pi0785), .ZN(new_n17222_));
  XNOR2_X1   g14274(.A1(new_n17222_), .A2(new_n17215_), .ZN(new_n17223_));
  OAI21_X1   g14275(.A1(new_n17204_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n17224_));
  AOI21_X1   g14276(.A1(new_n17223_), .A2(pi0618), .B(new_n17224_), .ZN(new_n17225_));
  INV_X1     g14277(.I(new_n17223_), .ZN(new_n17226_));
  AOI21_X1   g14278(.A1(new_n17204_), .A2(new_n11934_), .B(pi1154), .ZN(new_n17227_));
  OAI21_X1   g14279(.A1(new_n17226_), .A2(new_n11934_), .B(new_n17227_), .ZN(new_n17228_));
  NAND2_X1   g14280(.A1(new_n17228_), .A2(new_n17225_), .ZN(new_n17229_));
  MUX2_X1    g14281(.I0(new_n17229_), .I1(new_n17223_), .S(new_n11969_), .Z(new_n17230_));
  NAND2_X1   g14282(.A1(new_n17230_), .A2(new_n11985_), .ZN(new_n17231_));
  NOR3_X1    g14283(.A1(new_n17203_), .A2(pi0619), .A3(pi1159), .ZN(new_n17232_));
  NOR2_X1    g14284(.A1(new_n17232_), .A2(new_n11985_), .ZN(new_n17233_));
  XOR2_X1    g14285(.A1(new_n17231_), .A2(new_n17233_), .Z(new_n17234_));
  OAI21_X1   g14286(.A1(new_n17234_), .A2(new_n11997_), .B(new_n17205_), .ZN(new_n17235_));
  NOR2_X1    g14287(.A1(new_n17203_), .A2(new_n12054_), .ZN(new_n17236_));
  AOI21_X1   g14288(.A1(new_n17235_), .A2(new_n12054_), .B(new_n17236_), .ZN(new_n17237_));
  INV_X1     g14289(.I(new_n17237_), .ZN(new_n17238_));
  NOR2_X1    g14290(.A1(new_n17203_), .A2(new_n12092_), .ZN(new_n17239_));
  AOI21_X1   g14291(.A1(new_n17238_), .A2(new_n12092_), .B(new_n17239_), .ZN(new_n17240_));
  NAND2_X1   g14292(.A1(new_n17240_), .A2(new_n12082_), .ZN(new_n17241_));
  AOI21_X1   g14293(.A1(new_n17203_), .A2(pi0644), .B(new_n12099_), .ZN(new_n17242_));
  AOI21_X1   g14294(.A1(new_n17241_), .A2(new_n17242_), .B(pi1160), .ZN(new_n17243_));
  NOR2_X1    g14295(.A1(new_n17203_), .A2(new_n13114_), .ZN(new_n17244_));
  NOR2_X1    g14296(.A1(new_n17204_), .A2(new_n12014_), .ZN(new_n17245_));
  NOR2_X1    g14297(.A1(new_n17203_), .A2(new_n11961_), .ZN(new_n17246_));
  NAND2_X1   g14298(.A1(new_n8913_), .A2(new_n15745_), .ZN(new_n17247_));
  OAI21_X1   g14299(.A1(new_n12902_), .A2(new_n17247_), .B(new_n3231_), .ZN(new_n17248_));
  NOR3_X1    g14300(.A1(new_n13399_), .A2(pi0175), .A3(new_n13396_), .ZN(new_n17249_));
  AOI21_X1   g14301(.A1(new_n13399_), .A2(new_n8913_), .B(new_n13395_), .ZN(new_n17250_));
  NAND3_X1   g14302(.A1(new_n13403_), .A2(new_n3172_), .A3(new_n15745_), .ZN(new_n17251_));
  NOR4_X1    g14303(.A1(new_n17249_), .A2(new_n17250_), .A3(new_n17210_), .A4(new_n17251_), .ZN(new_n17252_));
  AOI22_X1   g14304(.A1(new_n17252_), .A2(new_n17248_), .B1(pi0175), .B2(new_n3232_), .ZN(new_n17253_));
  NAND2_X1   g14305(.A1(new_n17253_), .A2(new_n11891_), .ZN(new_n17254_));
  AOI21_X1   g14306(.A1(new_n17253_), .A2(new_n12970_), .B(new_n17204_), .ZN(new_n17255_));
  NOR3_X1    g14307(.A1(new_n17253_), .A2(pi0625), .A3(new_n17203_), .ZN(new_n17256_));
  NOR3_X1    g14308(.A1(new_n17256_), .A2(new_n17255_), .A3(pi1153), .ZN(new_n17257_));
  NAND4_X1   g14309(.A1(new_n17253_), .A2(pi0625), .A3(new_n11893_), .A4(new_n17204_), .ZN(new_n17258_));
  NAND2_X1   g14310(.A1(new_n17257_), .A2(new_n17258_), .ZN(new_n17259_));
  NAND2_X1   g14311(.A1(new_n17259_), .A2(pi0778), .ZN(new_n17260_));
  XOR2_X1    g14312(.A1(new_n17260_), .A2(new_n17254_), .Z(new_n17261_));
  NOR2_X1    g14313(.A1(new_n17261_), .A2(new_n13024_), .ZN(new_n17262_));
  AOI21_X1   g14314(.A1(new_n13024_), .A2(new_n17203_), .B(new_n17262_), .ZN(new_n17263_));
  AOI21_X1   g14315(.A1(new_n17263_), .A2(new_n11961_), .B(new_n17246_), .ZN(new_n17264_));
  AOI21_X1   g14316(.A1(new_n17264_), .A2(new_n12014_), .B(new_n17245_), .ZN(new_n17265_));
  AOI21_X1   g14317(.A1(new_n17265_), .A2(new_n13114_), .B(new_n17244_), .ZN(new_n17266_));
  NOR2_X1    g14318(.A1(new_n17266_), .A2(pi0628), .ZN(new_n17267_));
  AOI21_X1   g14319(.A1(pi0628), .A2(new_n17204_), .B(new_n17267_), .ZN(new_n17268_));
  NOR2_X1    g14320(.A1(new_n17268_), .A2(pi1156), .ZN(new_n17269_));
  NOR2_X1    g14321(.A1(new_n17266_), .A2(new_n12031_), .ZN(new_n17270_));
  AOI21_X1   g14322(.A1(new_n12031_), .A2(new_n17204_), .B(new_n17270_), .ZN(new_n17271_));
  NOR2_X1    g14323(.A1(new_n17271_), .A2(new_n12026_), .ZN(new_n17272_));
  OAI21_X1   g14324(.A1(new_n17269_), .A2(new_n17272_), .B(pi0792), .ZN(new_n17273_));
  OAI21_X1   g14325(.A1(pi0792), .A2(new_n17266_), .B(new_n17273_), .ZN(new_n17274_));
  NOR2_X1    g14326(.A1(new_n17203_), .A2(new_n12061_), .ZN(new_n17275_));
  AOI21_X1   g14327(.A1(new_n17274_), .A2(new_n12061_), .B(new_n17275_), .ZN(new_n17276_));
  NOR2_X1    g14328(.A1(new_n17276_), .A2(pi1157), .ZN(new_n17277_));
  NOR2_X1    g14329(.A1(new_n17203_), .A2(pi0647), .ZN(new_n17278_));
  AOI21_X1   g14330(.A1(new_n17274_), .A2(pi0647), .B(new_n17278_), .ZN(new_n17279_));
  NOR2_X1    g14331(.A1(new_n17279_), .A2(new_n12049_), .ZN(new_n17280_));
  NOR2_X1    g14332(.A1(new_n17277_), .A2(new_n17280_), .ZN(new_n17281_));
  NOR2_X1    g14333(.A1(new_n17281_), .A2(new_n12048_), .ZN(new_n17282_));
  AOI21_X1   g14334(.A1(new_n12048_), .A2(new_n17274_), .B(new_n17282_), .ZN(new_n17283_));
  NAND2_X1   g14335(.A1(new_n17283_), .A2(pi0644), .ZN(new_n17284_));
  AOI21_X1   g14336(.A1(new_n17284_), .A2(new_n12099_), .B(new_n17243_), .ZN(new_n17285_));
  NOR3_X1    g14337(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n17286_));
  NAND2_X1   g14338(.A1(new_n17240_), .A2(new_n17286_), .ZN(new_n17287_));
  NAND2_X1   g14339(.A1(new_n17287_), .A2(pi0715), .ZN(new_n17288_));
  AOI21_X1   g14340(.A1(new_n17283_), .A2(new_n12082_), .B(new_n17288_), .ZN(new_n17289_));
  OAI21_X1   g14341(.A1(new_n17285_), .A2(new_n17289_), .B(pi0790), .ZN(new_n17290_));
  NAND2_X1   g14342(.A1(new_n17243_), .A2(new_n12082_), .ZN(new_n17291_));
  AOI21_X1   g14343(.A1(new_n17287_), .A2(pi0644), .B(pi0790), .ZN(new_n17292_));
  NAND2_X1   g14344(.A1(new_n17291_), .A2(new_n17292_), .ZN(new_n17293_));
  NAND2_X1   g14345(.A1(new_n17279_), .A2(new_n12060_), .ZN(new_n17294_));
  AOI21_X1   g14346(.A1(new_n17276_), .A2(pi0630), .B(new_n12090_), .ZN(new_n17295_));
  NAND2_X1   g14347(.A1(new_n17238_), .A2(new_n15078_), .ZN(new_n17296_));
  AOI21_X1   g14348(.A1(new_n17295_), .A2(new_n17294_), .B(new_n17296_), .ZN(new_n17297_));
  AND2_X2    g14349(.A1(new_n17271_), .A2(new_n12030_), .Z(new_n17298_));
  INV_X1     g14350(.I(new_n12052_), .ZN(new_n17299_));
  NAND2_X1   g14351(.A1(new_n17268_), .A2(pi0629), .ZN(new_n17300_));
  NAND2_X1   g14352(.A1(new_n17300_), .A2(new_n17299_), .ZN(new_n17301_));
  OR2_X2     g14353(.A1(new_n17301_), .A2(new_n17298_), .Z(new_n17302_));
  INV_X1     g14354(.I(new_n15222_), .ZN(new_n17303_));
  NOR2_X1    g14355(.A1(new_n17303_), .A2(pi0792), .ZN(new_n17304_));
  NAND3_X1   g14356(.A1(new_n17302_), .A2(new_n17235_), .A3(new_n17304_), .ZN(new_n17305_));
  NAND2_X1   g14357(.A1(new_n17230_), .A2(pi0619), .ZN(new_n17306_));
  NAND2_X1   g14358(.A1(new_n17203_), .A2(pi0619), .ZN(new_n17307_));
  INV_X1     g14359(.I(new_n17213_), .ZN(new_n17308_));
  NOR2_X1    g14360(.A1(new_n12110_), .A2(new_n12111_), .ZN(new_n17309_));
  NAND2_X1   g14361(.A1(new_n17309_), .A2(new_n15707_), .ZN(new_n17310_));
  AOI21_X1   g14362(.A1(new_n12122_), .A2(new_n17310_), .B(pi0039), .ZN(new_n17311_));
  AOI21_X1   g14363(.A1(new_n13644_), .A2(new_n17110_), .B(new_n8913_), .ZN(new_n17312_));
  AOI21_X1   g14364(.A1(new_n17312_), .A2(new_n5156_), .B(new_n3172_), .ZN(new_n17313_));
  OAI21_X1   g14365(.A1(new_n17311_), .A2(pi0175), .B(new_n17313_), .ZN(new_n17314_));
  NOR2_X1    g14366(.A1(new_n13333_), .A2(new_n8913_), .ZN(new_n17315_));
  OAI21_X1   g14367(.A1(new_n12515_), .A2(new_n8913_), .B(new_n15707_), .ZN(new_n17316_));
  NOR3_X1    g14368(.A1(new_n12645_), .A2(new_n8913_), .A3(new_n13347_), .ZN(new_n17317_));
  AOI21_X1   g14369(.A1(new_n12645_), .A2(pi0175), .B(new_n12665_), .ZN(new_n17318_));
  OAI21_X1   g14370(.A1(new_n17317_), .A2(new_n17318_), .B(pi0766), .ZN(new_n17319_));
  NAND2_X1   g14371(.A1(new_n13360_), .A2(pi0175), .ZN(new_n17320_));
  NAND2_X1   g14372(.A1(new_n13362_), .A2(pi0175), .ZN(new_n17321_));
  NAND4_X1   g14373(.A1(new_n17319_), .A2(new_n15731_), .A3(new_n17320_), .A4(new_n17321_), .ZN(new_n17322_));
  AOI21_X1   g14374(.A1(new_n17322_), .A2(new_n3172_), .B(pi0039), .ZN(new_n17323_));
  OAI21_X1   g14375(.A1(new_n17315_), .A2(new_n17316_), .B(new_n17323_), .ZN(new_n17324_));
  NAND2_X1   g14376(.A1(new_n3232_), .A2(new_n15745_), .ZN(new_n17325_));
  AOI21_X1   g14377(.A1(new_n17324_), .A2(new_n17314_), .B(new_n17325_), .ZN(new_n17326_));
  NAND2_X1   g14378(.A1(new_n17209_), .A2(new_n17211_), .ZN(new_n17327_));
  NAND2_X1   g14379(.A1(new_n17327_), .A2(new_n15745_), .ZN(new_n17328_));
  OAI22_X1   g14380(.A1(new_n17326_), .A2(new_n17328_), .B1(new_n8913_), .B2(new_n3231_), .ZN(new_n17329_));
  OAI21_X1   g14381(.A1(new_n17329_), .A2(pi0625), .B(new_n17308_), .ZN(new_n17330_));
  NAND3_X1   g14382(.A1(new_n17329_), .A2(new_n12970_), .A3(new_n17213_), .ZN(new_n17331_));
  NAND4_X1   g14383(.A1(new_n17330_), .A2(new_n17331_), .A3(new_n12977_), .A4(new_n17258_), .ZN(new_n17332_));
  INV_X1     g14384(.I(new_n17257_), .ZN(new_n17333_));
  NOR4_X1    g14385(.A1(new_n17329_), .A2(new_n12970_), .A3(pi1153), .A4(new_n17308_), .ZN(new_n17334_));
  OAI21_X1   g14386(.A1(new_n17334_), .A2(new_n17333_), .B(new_n13657_), .ZN(new_n17335_));
  NAND2_X1   g14387(.A1(new_n17332_), .A2(new_n17335_), .ZN(new_n17336_));
  NOR2_X1    g14388(.A1(new_n17329_), .A2(pi0778), .ZN(new_n17337_));
  AOI21_X1   g14389(.A1(new_n17336_), .A2(pi0778), .B(new_n17337_), .ZN(new_n17338_));
  NOR2_X1    g14390(.A1(new_n17338_), .A2(pi0785), .ZN(new_n17339_));
  INV_X1     g14391(.I(new_n17261_), .ZN(new_n17340_));
  NAND3_X1   g14392(.A1(new_n17340_), .A2(pi0609), .A3(pi1155), .ZN(new_n17341_));
  NAND3_X1   g14393(.A1(new_n17341_), .A2(new_n11923_), .A3(new_n17220_), .ZN(new_n17342_));
  NOR4_X1    g14394(.A1(new_n17338_), .A2(new_n11903_), .A3(new_n17340_), .A4(pi1155), .ZN(new_n17343_));
  NAND2_X1   g14395(.A1(new_n17218_), .A2(pi0660), .ZN(new_n17344_));
  NOR2_X1    g14396(.A1(new_n17343_), .A2(new_n17344_), .ZN(new_n17345_));
  NOR2_X1    g14397(.A1(new_n17345_), .A2(new_n11870_), .ZN(new_n17346_));
  AOI21_X1   g14398(.A1(new_n17346_), .A2(new_n17342_), .B(new_n17339_), .ZN(new_n17347_));
  INV_X1     g14399(.I(new_n17263_), .ZN(new_n17348_));
  NOR4_X1    g14400(.A1(new_n17347_), .A2(new_n11934_), .A3(pi1154), .A4(new_n17348_), .ZN(new_n17349_));
  NAND2_X1   g14401(.A1(new_n17225_), .A2(pi0627), .ZN(new_n17350_));
  NOR3_X1    g14402(.A1(new_n17263_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n17351_));
  NAND2_X1   g14403(.A1(new_n17228_), .A2(new_n11949_), .ZN(new_n17352_));
  OAI22_X1   g14404(.A1(new_n17349_), .A2(new_n17350_), .B1(new_n17351_), .B2(new_n17352_), .ZN(new_n17353_));
  MUX2_X1    g14405(.I0(new_n17353_), .I1(new_n17347_), .S(new_n11969_), .Z(new_n17354_));
  XNOR2_X1   g14406(.A1(new_n17354_), .A2(new_n17264_), .ZN(new_n17355_));
  NOR2_X1    g14407(.A1(new_n17355_), .A2(new_n11967_), .ZN(new_n17356_));
  NAND3_X1   g14408(.A1(new_n17306_), .A2(new_n11869_), .A3(new_n17307_), .ZN(new_n17357_));
  XOR2_X1    g14409(.A1(new_n17356_), .A2(new_n17354_), .Z(new_n17358_));
  AOI21_X1   g14410(.A1(new_n17204_), .A2(new_n11967_), .B(pi1159), .ZN(new_n17359_));
  AOI21_X1   g14411(.A1(new_n17306_), .A2(new_n17359_), .B(pi0648), .ZN(new_n17360_));
  OAI21_X1   g14412(.A1(new_n17358_), .A2(pi1159), .B(new_n17360_), .ZN(new_n17361_));
  OR2_X2     g14413(.A1(new_n17354_), .A2(pi0789), .Z(new_n17362_));
  NAND3_X1   g14414(.A1(new_n17234_), .A2(pi0626), .A3(new_n17204_), .ZN(new_n17363_));
  OAI21_X1   g14415(.A1(new_n17234_), .A2(new_n11994_), .B(new_n17203_), .ZN(new_n17364_));
  AOI21_X1   g14416(.A1(new_n17364_), .A2(new_n17363_), .B(new_n17167_), .ZN(new_n17365_));
  AOI21_X1   g14417(.A1(new_n17234_), .A2(new_n17204_), .B(new_n11994_), .ZN(new_n17366_));
  NAND2_X1   g14418(.A1(new_n17366_), .A2(new_n11990_), .ZN(new_n17367_));
  NOR2_X1    g14419(.A1(new_n17265_), .A2(new_n12020_), .ZN(new_n17368_));
  NOR2_X1    g14420(.A1(new_n17368_), .A2(pi0788), .ZN(new_n17369_));
  NAND2_X1   g14421(.A1(new_n17367_), .A2(new_n17369_), .ZN(new_n17370_));
  INV_X1     g14422(.I(new_n14707_), .ZN(new_n17371_));
  NOR2_X1    g14423(.A1(new_n14731_), .A2(new_n17371_), .ZN(new_n17372_));
  OAI21_X1   g14424(.A1(new_n17370_), .A2(new_n17365_), .B(new_n17372_), .ZN(new_n17373_));
  AOI21_X1   g14425(.A1(new_n11998_), .A2(new_n17362_), .B(new_n17373_), .ZN(new_n17374_));
  NAND3_X1   g14426(.A1(new_n17361_), .A2(new_n17357_), .A3(new_n17374_), .ZN(new_n17375_));
  AOI21_X1   g14427(.A1(new_n17375_), .A2(new_n17305_), .B(new_n14725_), .ZN(new_n17376_));
  OAI21_X1   g14428(.A1(new_n17376_), .A2(new_n17297_), .B(new_n17293_), .ZN(new_n17377_));
  AOI21_X1   g14429(.A1(new_n17290_), .A2(new_n17377_), .B(po1038), .ZN(new_n17378_));
  OAI21_X1   g14430(.A1(new_n6845_), .A2(pi0175), .B(new_n13184_), .ZN(new_n17379_));
  OAI21_X1   g14431(.A1(new_n17378_), .A2(new_n17379_), .B(new_n17202_), .ZN(po0332));
  NOR2_X1    g14432(.A1(new_n2925_), .A2(pi0176), .ZN(new_n17381_));
  NOR2_X1    g14433(.A1(new_n11877_), .A2(pi0742), .ZN(new_n17382_));
  NOR2_X1    g14434(.A1(new_n17382_), .A2(new_n17381_), .ZN(new_n17383_));
  INV_X1     g14435(.I(new_n17383_), .ZN(new_n17384_));
  AOI21_X1   g14436(.A1(new_n11886_), .A2(new_n15756_), .B(new_n17381_), .ZN(new_n17385_));
  NOR2_X1    g14437(.A1(new_n17385_), .A2(new_n11874_), .ZN(new_n17386_));
  NOR2_X1    g14438(.A1(new_n17384_), .A2(new_n17386_), .ZN(new_n17387_));
  NOR2_X1    g14439(.A1(new_n17387_), .A2(pi0778), .ZN(new_n17388_));
  NAND2_X1   g14440(.A1(new_n17386_), .A2(pi0625), .ZN(new_n17389_));
  NOR3_X1    g14441(.A1(new_n11894_), .A2(pi0625), .A3(pi0704), .ZN(new_n17390_));
  NOR4_X1    g14442(.A1(new_n17382_), .A2(pi0608), .A3(new_n11893_), .A4(new_n17381_), .ZN(new_n17391_));
  OAI21_X1   g14443(.A1(new_n17384_), .A2(new_n17386_), .B(new_n17389_), .ZN(new_n17392_));
  NOR3_X1    g14444(.A1(new_n17381_), .A2(pi0608), .A3(pi1153), .ZN(new_n17393_));
  AOI22_X1   g14445(.A1(new_n17392_), .A2(new_n17393_), .B1(new_n17389_), .B2(new_n17391_), .ZN(new_n17394_));
  NOR2_X1    g14446(.A1(new_n17394_), .A2(new_n11891_), .ZN(new_n17395_));
  XOR2_X1    g14447(.A1(new_n17395_), .A2(new_n17388_), .Z(new_n17396_));
  INV_X1     g14448(.I(new_n17396_), .ZN(new_n17397_));
  NAND2_X1   g14449(.A1(new_n17397_), .A2(new_n11870_), .ZN(new_n17398_));
  AOI21_X1   g14450(.A1(new_n17396_), .A2(new_n11903_), .B(pi1155), .ZN(new_n17399_));
  INV_X1     g14451(.I(new_n17385_), .ZN(new_n17400_));
  XOR2_X1    g14452(.A1(new_n17390_), .A2(pi1153), .Z(new_n17401_));
  NAND2_X1   g14453(.A1(new_n17401_), .A2(new_n17400_), .ZN(new_n17402_));
  OAI21_X1   g14454(.A1(new_n17390_), .A2(new_n17381_), .B(new_n11893_), .ZN(new_n17403_));
  AOI21_X1   g14455(.A1(new_n17402_), .A2(new_n17403_), .B(new_n11891_), .ZN(new_n17404_));
  NOR2_X1    g14456(.A1(new_n17385_), .A2(pi0778), .ZN(new_n17405_));
  OAI21_X1   g14457(.A1(new_n17404_), .A2(new_n17405_), .B(pi0609), .ZN(new_n17406_));
  AOI21_X1   g14458(.A1(new_n17384_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n17407_));
  NOR2_X1    g14459(.A1(new_n17407_), .A2(pi0660), .ZN(new_n17408_));
  OAI21_X1   g14460(.A1(new_n17399_), .A2(new_n17406_), .B(new_n17408_), .ZN(new_n17409_));
  NOR2_X1    g14461(.A1(new_n17404_), .A2(new_n17405_), .ZN(new_n17410_));
  NAND4_X1   g14462(.A1(new_n17397_), .A2(pi0609), .A3(new_n11912_), .A4(new_n17410_), .ZN(new_n17411_));
  NOR2_X1    g14463(.A1(new_n17383_), .A2(new_n11925_), .ZN(new_n17412_));
  AOI21_X1   g14464(.A1(new_n17412_), .A2(new_n11928_), .B(pi1155), .ZN(new_n17413_));
  NOR2_X1    g14465(.A1(new_n17413_), .A2(new_n11923_), .ZN(new_n17414_));
  NAND2_X1   g14466(.A1(new_n17411_), .A2(new_n17414_), .ZN(new_n17415_));
  NAND3_X1   g14467(.A1(new_n17415_), .A2(pi0785), .A3(new_n17409_), .ZN(new_n17416_));
  NAND2_X1   g14468(.A1(new_n17416_), .A2(new_n17398_), .ZN(new_n17417_));
  NOR4_X1    g14469(.A1(new_n17410_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n17419_));
  NOR2_X1    g14470(.A1(new_n17412_), .A2(pi0785), .ZN(new_n17420_));
  OAI21_X1   g14471(.A1(new_n17413_), .A2(new_n17407_), .B(pi0785), .ZN(new_n17421_));
  XNOR2_X1   g14472(.A1(new_n17421_), .A2(new_n17420_), .ZN(new_n17422_));
  INV_X1     g14473(.I(new_n17422_), .ZN(new_n17423_));
  NOR2_X1    g14474(.A1(new_n17423_), .A2(new_n11945_), .ZN(new_n17424_));
  NOR3_X1    g14475(.A1(new_n17424_), .A2(pi0627), .A3(new_n17419_), .ZN(new_n17425_));
  AOI21_X1   g14476(.A1(new_n17422_), .A2(new_n11951_), .B(pi1154), .ZN(new_n17426_));
  NOR2_X1    g14477(.A1(new_n17410_), .A2(new_n11939_), .ZN(new_n17427_));
  INV_X1     g14478(.I(new_n17427_), .ZN(new_n17428_));
  NAND4_X1   g14479(.A1(new_n17417_), .A2(pi0618), .A3(new_n11950_), .A4(new_n17428_), .ZN(new_n17429_));
  NAND2_X1   g14480(.A1(new_n17429_), .A2(new_n17426_), .ZN(new_n17430_));
  AOI21_X1   g14481(.A1(new_n17430_), .A2(new_n11949_), .B(new_n17425_), .ZN(new_n17431_));
  NOR2_X1    g14482(.A1(new_n17431_), .A2(new_n11969_), .ZN(new_n17432_));
  AOI21_X1   g14483(.A1(new_n11969_), .A2(new_n17417_), .B(new_n17432_), .ZN(new_n17433_));
  NOR2_X1    g14484(.A1(new_n17428_), .A2(new_n11962_), .ZN(new_n17434_));
  NOR4_X1    g14485(.A1(new_n17433_), .A2(new_n11967_), .A3(pi1159), .A4(new_n17434_), .ZN(new_n17435_));
  INV_X1     g14486(.I(new_n17424_), .ZN(new_n17436_));
  NAND2_X1   g14487(.A1(new_n17436_), .A2(new_n17426_), .ZN(new_n17437_));
  MUX2_X1    g14488(.I0(new_n17437_), .I1(new_n17422_), .S(new_n11969_), .Z(new_n17438_));
  NAND2_X1   g14489(.A1(new_n17438_), .A2(pi0619), .ZN(new_n17439_));
  INV_X1     g14490(.I(new_n17439_), .ZN(new_n17440_));
  INV_X1     g14491(.I(new_n17381_), .ZN(new_n17441_));
  OAI21_X1   g14492(.A1(new_n17441_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n17442_));
  NOR4_X1    g14493(.A1(new_n17435_), .A2(new_n11966_), .A3(new_n17440_), .A4(new_n17442_), .ZN(new_n17443_));
  NOR4_X1    g14494(.A1(new_n17428_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n17444_));
  OAI21_X1   g14495(.A1(new_n17381_), .A2(pi0619), .B(new_n11869_), .ZN(new_n17445_));
  OAI21_X1   g14496(.A1(new_n17440_), .A2(new_n17445_), .B(new_n11966_), .ZN(new_n17446_));
  NOR2_X1    g14497(.A1(new_n17446_), .A2(new_n17444_), .ZN(new_n17447_));
  AOI21_X1   g14498(.A1(new_n17433_), .A2(new_n11998_), .B(pi0789), .ZN(new_n17448_));
  OAI21_X1   g14499(.A1(new_n17443_), .A2(new_n17447_), .B(new_n17448_), .ZN(new_n17449_));
  INV_X1     g14500(.I(new_n12015_), .ZN(new_n17450_));
  NAND2_X1   g14501(.A1(new_n17434_), .A2(new_n17450_), .ZN(new_n17451_));
  NOR2_X1    g14502(.A1(new_n17451_), .A2(new_n17153_), .ZN(new_n17452_));
  INV_X1     g14503(.I(new_n17452_), .ZN(new_n17453_));
  NOR2_X1    g14504(.A1(new_n17453_), .A2(new_n17151_), .ZN(new_n17454_));
  NOR2_X1    g14505(.A1(new_n14624_), .A2(new_n17381_), .ZN(new_n17455_));
  NAND3_X1   g14506(.A1(new_n17441_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n17456_));
  MUX2_X1    g14507(.I0(new_n17456_), .I1(new_n17438_), .S(new_n11985_), .Z(new_n17457_));
  AOI21_X1   g14508(.A1(new_n17457_), .A2(new_n14624_), .B(new_n17455_), .ZN(new_n17458_));
  AND2_X2    g14509(.A1(new_n17458_), .A2(new_n12064_), .Z(new_n17459_));
  OAI21_X1   g14510(.A1(new_n17459_), .A2(new_n17454_), .B(pi0629), .ZN(new_n17460_));
  NAND2_X1   g14511(.A1(new_n17458_), .A2(new_n12063_), .ZN(new_n17461_));
  NAND2_X1   g14512(.A1(new_n17452_), .A2(new_n15084_), .ZN(new_n17462_));
  NAND4_X1   g14513(.A1(new_n17460_), .A2(new_n15085_), .A3(new_n17461_), .A4(new_n17462_), .ZN(new_n17463_));
  MUX2_X1    g14514(.I0(new_n17457_), .I1(new_n17441_), .S(new_n11994_), .Z(new_n17464_));
  NOR2_X1    g14515(.A1(new_n17464_), .A2(new_n17167_), .ZN(new_n17465_));
  OAI21_X1   g14516(.A1(new_n17457_), .A2(new_n17381_), .B(pi0626), .ZN(new_n17466_));
  NOR2_X1    g14517(.A1(new_n17451_), .A2(new_n12020_), .ZN(new_n17467_));
  NOR2_X1    g14518(.A1(new_n17467_), .A2(pi0788), .ZN(new_n17468_));
  OAI21_X1   g14519(.A1(new_n17466_), .A2(new_n17171_), .B(new_n17468_), .ZN(new_n17469_));
  OAI21_X1   g14520(.A1(new_n17465_), .A2(new_n17469_), .B(new_n14732_), .ZN(new_n17470_));
  AOI21_X1   g14521(.A1(new_n17463_), .A2(new_n14726_), .B(new_n17470_), .ZN(new_n17471_));
  NAND3_X1   g14522(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n17381_), .ZN(new_n17472_));
  NOR2_X1    g14523(.A1(new_n17453_), .A2(new_n12068_), .ZN(new_n17473_));
  INV_X1     g14524(.I(new_n17473_), .ZN(new_n17474_));
  NAND2_X1   g14525(.A1(new_n17474_), .A2(pi0647), .ZN(new_n17475_));
  NAND2_X1   g14526(.A1(new_n17381_), .A2(pi0647), .ZN(new_n17476_));
  NAND3_X1   g14527(.A1(new_n17475_), .A2(new_n12049_), .A3(new_n17476_), .ZN(new_n17477_));
  NOR2_X1    g14528(.A1(new_n17441_), .A2(pi0647), .ZN(new_n17478_));
  AOI21_X1   g14529(.A1(new_n17473_), .A2(pi0647), .B(new_n17478_), .ZN(new_n17479_));
  NAND2_X1   g14530(.A1(new_n17479_), .A2(new_n12088_), .ZN(new_n17480_));
  NAND2_X1   g14531(.A1(new_n17480_), .A2(pi0787), .ZN(new_n17481_));
  AOI21_X1   g14532(.A1(pi0630), .A2(new_n17477_), .B(new_n17481_), .ZN(new_n17482_));
  AOI22_X1   g14533(.A1(new_n17449_), .A2(new_n17471_), .B1(new_n17472_), .B2(new_n17482_), .ZN(new_n17483_));
  NOR2_X1    g14534(.A1(new_n17483_), .A2(new_n12082_), .ZN(new_n17484_));
  NAND4_X1   g14535(.A1(new_n17475_), .A2(pi0787), .A3(new_n12049_), .A4(new_n17476_), .ZN(new_n17485_));
  OAI21_X1   g14536(.A1(pi0787), .A2(new_n17474_), .B(new_n17485_), .ZN(new_n17486_));
  NOR2_X1    g14537(.A1(new_n17486_), .A2(pi0644), .ZN(new_n17487_));
  OR3_X2     g14538(.A1(new_n17484_), .A2(pi0715), .A3(new_n17487_), .Z(new_n17488_));
  MUX2_X1    g14539(.I0(new_n17458_), .I1(new_n17381_), .S(new_n16841_), .Z(new_n17489_));
  INV_X1     g14540(.I(new_n17489_), .ZN(new_n17490_));
  OAI21_X1   g14541(.A1(new_n17489_), .A2(new_n17381_), .B(new_n12082_), .ZN(new_n17491_));
  AOI21_X1   g14542(.A1(new_n17381_), .A2(new_n17489_), .B(new_n17491_), .ZN(new_n17492_));
  OAI21_X1   g14543(.A1(new_n17492_), .A2(new_n17490_), .B(new_n12099_), .ZN(new_n17493_));
  AOI21_X1   g14544(.A1(new_n17490_), .A2(new_n17492_), .B(new_n17493_), .ZN(new_n17494_));
  AOI21_X1   g14545(.A1(new_n17488_), .A2(new_n17494_), .B(pi1160), .ZN(new_n17495_));
  XOR2_X1    g14546(.A1(new_n17492_), .A2(new_n17381_), .Z(new_n17496_));
  AOI21_X1   g14547(.A1(new_n17486_), .A2(pi0644), .B(new_n13169_), .ZN(new_n17497_));
  OAI21_X1   g14548(.A1(new_n17496_), .A2(new_n12099_), .B(new_n17497_), .ZN(new_n17498_));
  OAI21_X1   g14549(.A1(new_n17484_), .A2(new_n17498_), .B(pi0790), .ZN(new_n17499_));
  NOR2_X1    g14550(.A1(new_n17483_), .A2(new_n14748_), .ZN(new_n17500_));
  OAI21_X1   g14551(.A1(new_n17495_), .A2(new_n17499_), .B(new_n17500_), .ZN(new_n17501_));
  NOR2_X1    g14552(.A1(new_n12965_), .A2(pi0176), .ZN(new_n17502_));
  INV_X1     g14553(.I(new_n17502_), .ZN(new_n17503_));
  NAND2_X1   g14554(.A1(new_n17503_), .A2(new_n11997_), .ZN(new_n17504_));
  NOR2_X1    g14555(.A1(new_n14358_), .A2(new_n3172_), .ZN(new_n17505_));
  AOI21_X1   g14556(.A1(new_n12694_), .A2(new_n3172_), .B(new_n17505_), .ZN(new_n17506_));
  OAI21_X1   g14557(.A1(new_n14365_), .A2(pi0176), .B(new_n15764_), .ZN(new_n17507_));
  AOI21_X1   g14558(.A1(pi0176), .A2(new_n17506_), .B(new_n17507_), .ZN(new_n17508_));
  AOI21_X1   g14559(.A1(new_n15823_), .A2(new_n7150_), .B(new_n15764_), .ZN(new_n17509_));
  XOR2_X1    g14560(.A1(new_n17508_), .A2(new_n17509_), .Z(new_n17510_));
  NOR2_X1    g14561(.A1(new_n17510_), .A2(new_n3232_), .ZN(new_n17511_));
  NOR2_X1    g14562(.A1(new_n3231_), .A2(pi0176), .ZN(new_n17512_));
  NOR2_X1    g14563(.A1(new_n17511_), .A2(new_n17512_), .ZN(new_n17513_));
  INV_X1     g14564(.I(new_n17513_), .ZN(new_n17514_));
  OAI21_X1   g14565(.A1(new_n17503_), .A2(new_n11924_), .B(new_n11870_), .ZN(new_n17515_));
  AOI21_X1   g14566(.A1(new_n17514_), .A2(new_n11924_), .B(new_n17515_), .ZN(new_n17516_));
  NAND2_X1   g14567(.A1(new_n17513_), .A2(new_n11924_), .ZN(new_n17517_));
  OAI22_X1   g14568(.A1(new_n17517_), .A2(pi0609), .B1(new_n12996_), .B2(new_n17502_), .ZN(new_n17518_));
  NAND2_X1   g14569(.A1(new_n17518_), .A2(new_n11912_), .ZN(new_n17519_));
  OAI22_X1   g14570(.A1(new_n17517_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n17502_), .ZN(new_n17520_));
  NAND2_X1   g14571(.A1(new_n17520_), .A2(pi1155), .ZN(new_n17521_));
  AOI21_X1   g14572(.A1(new_n17519_), .A2(new_n17521_), .B(new_n11870_), .ZN(new_n17522_));
  XNOR2_X1   g14573(.A1(new_n17522_), .A2(new_n17516_), .ZN(new_n17523_));
  NOR2_X1    g14574(.A1(new_n17523_), .A2(pi0781), .ZN(new_n17524_));
  NOR2_X1    g14575(.A1(new_n17523_), .A2(new_n11934_), .ZN(new_n17525_));
  OAI21_X1   g14576(.A1(new_n17503_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n17526_));
  NOR2_X1    g14577(.A1(new_n17525_), .A2(new_n17526_), .ZN(new_n17527_));
  AOI21_X1   g14578(.A1(new_n17503_), .A2(new_n11934_), .B(pi1154), .ZN(new_n17528_));
  OAI21_X1   g14579(.A1(new_n17523_), .A2(new_n11934_), .B(new_n17528_), .ZN(new_n17529_));
  AOI21_X1   g14580(.A1(new_n17527_), .A2(new_n17529_), .B(new_n11969_), .ZN(new_n17530_));
  XOR2_X1    g14581(.A1(new_n17530_), .A2(new_n17524_), .Z(new_n17531_));
  NOR2_X1    g14582(.A1(new_n17531_), .A2(pi0789), .ZN(new_n17532_));
  INV_X1     g14583(.I(new_n17531_), .ZN(new_n17533_));
  MUX2_X1    g14584(.I0(new_n17502_), .I1(new_n17533_), .S(new_n14640_), .Z(new_n17534_));
  AOI21_X1   g14585(.A1(new_n17534_), .A2(pi0789), .B(new_n17532_), .ZN(new_n17535_));
  NAND2_X1   g14586(.A1(new_n17535_), .A2(new_n14624_), .ZN(new_n17536_));
  AOI21_X1   g14587(.A1(new_n17536_), .A2(new_n17504_), .B(new_n12053_), .ZN(new_n17537_));
  NOR2_X1    g14588(.A1(new_n17502_), .A2(new_n12054_), .ZN(new_n17538_));
  OAI21_X1   g14589(.A1(new_n17537_), .A2(new_n17538_), .B(new_n12092_), .ZN(new_n17539_));
  NOR2_X1    g14590(.A1(new_n17502_), .A2(new_n12092_), .ZN(new_n17540_));
  INV_X1     g14591(.I(new_n17540_), .ZN(new_n17541_));
  NAND3_X1   g14592(.A1(new_n17539_), .A2(new_n12082_), .A3(new_n17541_), .ZN(new_n17542_));
  AOI21_X1   g14593(.A1(new_n17502_), .A2(pi0644), .B(new_n12099_), .ZN(new_n17543_));
  NAND2_X1   g14594(.A1(new_n17542_), .A2(new_n17543_), .ZN(new_n17544_));
  INV_X1     g14595(.I(new_n13402_), .ZN(new_n17545_));
  MUX2_X1    g14596(.I0(new_n13396_), .I1(new_n17545_), .S(new_n3172_), .Z(new_n17546_));
  NOR2_X1    g14597(.A1(new_n17546_), .A2(new_n3231_), .ZN(new_n17547_));
  NOR2_X1    g14598(.A1(new_n17547_), .A2(new_n7150_), .ZN(new_n17548_));
  NAND2_X1   g14599(.A1(new_n17548_), .A2(new_n11891_), .ZN(new_n17549_));
  NOR3_X1    g14600(.A1(new_n17502_), .A2(pi0625), .A3(pi1153), .ZN(new_n17550_));
  NOR2_X1    g14601(.A1(new_n17550_), .A2(new_n11891_), .ZN(new_n17551_));
  XNOR2_X1   g14602(.A1(new_n17551_), .A2(new_n17549_), .ZN(new_n17552_));
  NOR2_X1    g14603(.A1(new_n17552_), .A2(new_n13024_), .ZN(new_n17553_));
  AOI21_X1   g14604(.A1(new_n13024_), .A2(new_n17502_), .B(new_n17553_), .ZN(new_n17554_));
  INV_X1     g14605(.I(new_n17554_), .ZN(new_n17555_));
  NOR2_X1    g14606(.A1(new_n17555_), .A2(new_n13714_), .ZN(new_n17556_));
  AOI21_X1   g14607(.A1(new_n13714_), .A2(new_n17503_), .B(new_n17556_), .ZN(new_n17557_));
  INV_X1     g14608(.I(new_n17557_), .ZN(new_n17558_));
  MUX2_X1    g14609(.I0(new_n17558_), .I1(new_n17503_), .S(new_n13713_), .Z(new_n17559_));
  NAND2_X1   g14610(.A1(new_n17559_), .A2(new_n11868_), .ZN(new_n17560_));
  MUX2_X1    g14611(.I0(new_n17559_), .I1(new_n17503_), .S(new_n14727_), .Z(new_n17561_));
  NAND2_X1   g14612(.A1(new_n17561_), .A2(pi0792), .ZN(new_n17562_));
  NAND2_X1   g14613(.A1(new_n17562_), .A2(new_n17560_), .ZN(new_n17563_));
  INV_X1     g14614(.I(new_n17563_), .ZN(new_n17564_));
  NOR2_X1    g14615(.A1(new_n17564_), .A2(pi0787), .ZN(new_n17565_));
  NAND2_X1   g14616(.A1(new_n17503_), .A2(pi0647), .ZN(new_n17566_));
  OAI21_X1   g14617(.A1(new_n17564_), .A2(pi0647), .B(new_n17566_), .ZN(new_n17567_));
  NAND2_X1   g14618(.A1(new_n17567_), .A2(new_n12049_), .ZN(new_n17568_));
  NOR2_X1    g14619(.A1(new_n17502_), .A2(pi0647), .ZN(new_n17569_));
  AOI21_X1   g14620(.A1(new_n17563_), .A2(pi0647), .B(new_n17569_), .ZN(new_n17570_));
  OAI21_X1   g14621(.A1(new_n17570_), .A2(new_n12049_), .B(new_n17568_), .ZN(new_n17571_));
  AOI21_X1   g14622(.A1(new_n17571_), .A2(pi0787), .B(new_n17565_), .ZN(new_n17572_));
  NAND2_X1   g14623(.A1(new_n17572_), .A2(pi0644), .ZN(new_n17573_));
  AOI22_X1   g14624(.A1(new_n17544_), .A2(new_n12081_), .B1(new_n12099_), .B2(new_n17573_), .ZN(new_n17574_));
  NOR3_X1    g14625(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n17575_));
  NAND3_X1   g14626(.A1(new_n17539_), .A2(new_n17541_), .A3(new_n17575_), .ZN(new_n17576_));
  NAND2_X1   g14627(.A1(new_n17572_), .A2(new_n12082_), .ZN(new_n17577_));
  AND3_X2    g14628(.A1(new_n17576_), .A2(pi0715), .A3(new_n17577_), .Z(new_n17578_));
  OAI21_X1   g14629(.A1(new_n17574_), .A2(new_n17578_), .B(pi0790), .ZN(new_n17579_));
  NOR2_X1    g14630(.A1(new_n17510_), .A2(new_n15756_), .ZN(new_n17580_));
  INV_X1     g14631(.I(new_n14352_), .ZN(new_n17581_));
  NOR2_X1    g14632(.A1(new_n14351_), .A2(new_n17581_), .ZN(new_n17582_));
  MUX2_X1    g14633(.I0(new_n17582_), .I1(new_n14347_), .S(pi0176), .Z(new_n17583_));
  AOI21_X1   g14634(.A1(new_n17583_), .A2(new_n15764_), .B(pi0704), .ZN(new_n17584_));
  OAI21_X1   g14635(.A1(new_n17580_), .A2(new_n17584_), .B(new_n3231_), .ZN(new_n17585_));
  XNOR2_X1   g14636(.A1(new_n17585_), .A2(new_n17512_), .ZN(new_n17586_));
  AOI21_X1   g14637(.A1(new_n17548_), .A2(pi0625), .B(pi1153), .ZN(new_n17587_));
  OAI21_X1   g14638(.A1(pi0625), .A2(new_n17502_), .B(new_n17587_), .ZN(new_n17588_));
  INV_X1     g14639(.I(new_n17586_), .ZN(new_n17589_));
  NOR2_X1    g14640(.A1(new_n17589_), .A2(new_n12970_), .ZN(new_n17590_));
  INV_X1     g14641(.I(new_n17590_), .ZN(new_n17591_));
  NAND2_X1   g14642(.A1(new_n17514_), .A2(pi0625), .ZN(new_n17592_));
  NAND4_X1   g14643(.A1(new_n17591_), .A2(new_n12977_), .A3(new_n17588_), .A4(new_n17592_), .ZN(new_n17593_));
  OAI21_X1   g14644(.A1(new_n12970_), .A2(new_n17503_), .B(new_n17587_), .ZN(new_n17594_));
  OAI21_X1   g14645(.A1(new_n17514_), .A2(pi0625), .B(new_n11893_), .ZN(new_n17595_));
  NOR2_X1    g14646(.A1(new_n17590_), .A2(new_n17595_), .ZN(new_n17596_));
  OAI21_X1   g14647(.A1(new_n17596_), .A2(new_n17594_), .B(new_n13657_), .ZN(new_n17597_));
  AOI21_X1   g14648(.A1(new_n17597_), .A2(new_n17593_), .B(new_n11891_), .ZN(new_n17598_));
  AOI21_X1   g14649(.A1(new_n11891_), .A2(new_n17586_), .B(new_n17598_), .ZN(new_n17599_));
  NOR2_X1    g14650(.A1(new_n17599_), .A2(pi0785), .ZN(new_n17600_));
  INV_X1     g14651(.I(new_n17552_), .ZN(new_n17601_));
  NAND3_X1   g14652(.A1(new_n17601_), .A2(pi0609), .A3(pi1155), .ZN(new_n17602_));
  NAND3_X1   g14653(.A1(new_n17521_), .A2(new_n11923_), .A3(new_n17602_), .ZN(new_n17603_));
  NOR4_X1    g14654(.A1(new_n17599_), .A2(new_n11903_), .A3(pi1155), .A4(new_n17601_), .ZN(new_n17604_));
  NAND2_X1   g14655(.A1(new_n17519_), .A2(pi0660), .ZN(new_n17605_));
  NOR2_X1    g14656(.A1(new_n17604_), .A2(new_n17605_), .ZN(new_n17606_));
  NOR2_X1    g14657(.A1(new_n17606_), .A2(new_n11870_), .ZN(new_n17607_));
  AOI21_X1   g14658(.A1(new_n17607_), .A2(new_n17603_), .B(new_n17600_), .ZN(new_n17608_));
  NOR4_X1    g14659(.A1(new_n17608_), .A2(new_n11934_), .A3(pi1154), .A4(new_n17555_), .ZN(new_n17609_));
  NAND2_X1   g14660(.A1(new_n17527_), .A2(pi0627), .ZN(new_n17610_));
  NOR3_X1    g14661(.A1(new_n17554_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n17611_));
  NAND2_X1   g14662(.A1(new_n17529_), .A2(new_n11949_), .ZN(new_n17612_));
  OAI22_X1   g14663(.A1(new_n17609_), .A2(new_n17610_), .B1(new_n17611_), .B2(new_n17612_), .ZN(new_n17613_));
  MUX2_X1    g14664(.I0(new_n17613_), .I1(new_n17608_), .S(new_n11969_), .Z(new_n17614_));
  NOR3_X1    g14665(.A1(new_n11869_), .A2(pi0619), .A3(pi0648), .ZN(new_n17615_));
  NAND2_X1   g14666(.A1(new_n11869_), .A2(pi0619), .ZN(new_n17616_));
  AOI21_X1   g14667(.A1(new_n17533_), .A2(new_n17615_), .B(new_n17616_), .ZN(new_n17617_));
  NAND2_X1   g14668(.A1(new_n17614_), .A2(new_n17617_), .ZN(new_n17618_));
  AND2_X2    g14669(.A1(new_n17614_), .A2(new_n11967_), .Z(new_n17619_));
  NAND2_X1   g14670(.A1(new_n11869_), .A2(pi0619), .ZN(new_n17620_));
  INV_X1     g14671(.I(new_n15278_), .ZN(new_n17621_));
  AOI21_X1   g14672(.A1(new_n17557_), .A2(pi0619), .B(new_n17621_), .ZN(new_n17622_));
  OAI21_X1   g14673(.A1(new_n17531_), .A2(new_n17620_), .B(new_n17622_), .ZN(new_n17623_));
  OAI21_X1   g14674(.A1(new_n17619_), .A2(new_n17623_), .B(new_n17618_), .ZN(new_n17624_));
  AOI21_X1   g14675(.A1(new_n17614_), .A2(new_n11998_), .B(pi0789), .ZN(new_n17625_));
  MUX2_X1    g14676(.I0(new_n17535_), .I1(new_n17503_), .S(new_n11994_), .Z(new_n17626_));
  INV_X1     g14677(.I(new_n17535_), .ZN(new_n17627_));
  AOI21_X1   g14678(.A1(new_n17627_), .A2(new_n17503_), .B(new_n11994_), .ZN(new_n17628_));
  MUX2_X1    g14679(.I0(new_n17502_), .I1(new_n17558_), .S(new_n12013_), .Z(new_n17629_));
  AOI22_X1   g14680(.A1(new_n17628_), .A2(new_n11990_), .B1(new_n12020_), .B2(new_n17629_), .ZN(new_n17630_));
  OAI21_X1   g14681(.A1(new_n17167_), .A2(new_n17626_), .B(new_n17630_), .ZN(new_n17631_));
  AOI22_X1   g14682(.A1(new_n17624_), .A2(new_n17625_), .B1(new_n17631_), .B2(pi0788), .ZN(new_n17632_));
  NAND2_X1   g14683(.A1(new_n17536_), .A2(new_n17504_), .ZN(new_n17633_));
  NAND2_X1   g14684(.A1(new_n17633_), .A2(new_n15222_), .ZN(new_n17634_));
  MUX2_X1    g14685(.I0(new_n17559_), .I1(new_n17503_), .S(pi0628), .Z(new_n17635_));
  NAND2_X1   g14686(.A1(new_n17559_), .A2(pi0628), .ZN(new_n17636_));
  OAI21_X1   g14687(.A1(pi0628), .A2(new_n17502_), .B(new_n17636_), .ZN(new_n17637_));
  AOI22_X1   g14688(.A1(new_n17637_), .A2(new_n12050_), .B1(new_n12051_), .B2(new_n17635_), .ZN(new_n17638_));
  NAND2_X1   g14689(.A1(new_n17634_), .A2(new_n17638_), .ZN(new_n17639_));
  AOI21_X1   g14690(.A1(new_n17634_), .A2(new_n17638_), .B(new_n14732_), .ZN(new_n17640_));
  OAI22_X1   g14691(.A1(new_n17640_), .A2(new_n14725_), .B1(new_n17639_), .B2(new_n11868_), .ZN(new_n17641_));
  NOR2_X1    g14692(.A1(new_n17537_), .A2(new_n17538_), .ZN(new_n17642_));
  AND2_X2    g14693(.A1(new_n17570_), .A2(new_n12060_), .Z(new_n17643_));
  OAI21_X1   g14694(.A1(new_n17567_), .A2(new_n12060_), .B(new_n15214_), .ZN(new_n17644_));
  OAI21_X1   g14695(.A1(new_n17644_), .A2(new_n17643_), .B(new_n15078_), .ZN(new_n17645_));
  NOR2_X1    g14696(.A1(new_n17642_), .A2(new_n17645_), .ZN(new_n17646_));
  NAND3_X1   g14697(.A1(new_n17544_), .A2(new_n12082_), .A3(new_n12081_), .ZN(new_n17647_));
  AOI21_X1   g14698(.A1(new_n17576_), .A2(pi0644), .B(pi0790), .ZN(new_n17648_));
  AOI21_X1   g14699(.A1(new_n17647_), .A2(new_n17648_), .B(new_n17646_), .ZN(new_n17649_));
  OAI21_X1   g14700(.A1(new_n17632_), .A2(new_n17641_), .B(new_n17649_), .ZN(new_n17650_));
  AOI21_X1   g14701(.A1(new_n17650_), .A2(new_n17579_), .B(po1038), .ZN(new_n17651_));
  OAI21_X1   g14702(.A1(new_n6845_), .A2(pi0176), .B(new_n13184_), .ZN(new_n17652_));
  OAI21_X1   g14703(.A1(new_n17651_), .A2(new_n17652_), .B(new_n17501_), .ZN(po0333));
  NOR2_X1    g14704(.A1(new_n2925_), .A2(pi0177), .ZN(new_n17654_));
  NOR2_X1    g14705(.A1(new_n11877_), .A2(pi0757), .ZN(new_n17655_));
  NOR2_X1    g14706(.A1(new_n17655_), .A2(new_n17654_), .ZN(new_n17656_));
  INV_X1     g14707(.I(new_n17656_), .ZN(new_n17657_));
  AOI21_X1   g14708(.A1(new_n11886_), .A2(new_n15794_), .B(new_n17654_), .ZN(new_n17658_));
  NOR2_X1    g14709(.A1(new_n17658_), .A2(new_n11874_), .ZN(new_n17659_));
  NOR2_X1    g14710(.A1(new_n17657_), .A2(new_n17659_), .ZN(new_n17660_));
  NOR2_X1    g14711(.A1(new_n17660_), .A2(pi0778), .ZN(new_n17661_));
  NAND2_X1   g14712(.A1(new_n17659_), .A2(pi0625), .ZN(new_n17662_));
  NOR3_X1    g14713(.A1(new_n11894_), .A2(pi0625), .A3(pi0686), .ZN(new_n17663_));
  NOR4_X1    g14714(.A1(new_n17655_), .A2(pi0608), .A3(new_n11893_), .A4(new_n17654_), .ZN(new_n17664_));
  OAI21_X1   g14715(.A1(new_n17657_), .A2(new_n17659_), .B(new_n17662_), .ZN(new_n17665_));
  NOR3_X1    g14716(.A1(new_n17654_), .A2(pi0608), .A3(pi1153), .ZN(new_n17666_));
  AOI22_X1   g14717(.A1(new_n17665_), .A2(new_n17666_), .B1(new_n17662_), .B2(new_n17664_), .ZN(new_n17667_));
  NOR2_X1    g14718(.A1(new_n17667_), .A2(new_n11891_), .ZN(new_n17668_));
  XOR2_X1    g14719(.A1(new_n17668_), .A2(new_n17661_), .Z(new_n17669_));
  INV_X1     g14720(.I(new_n17669_), .ZN(new_n17670_));
  NAND2_X1   g14721(.A1(new_n17670_), .A2(new_n11870_), .ZN(new_n17671_));
  AOI21_X1   g14722(.A1(new_n17669_), .A2(new_n11903_), .B(pi1155), .ZN(new_n17672_));
  INV_X1     g14723(.I(new_n17658_), .ZN(new_n17673_));
  XOR2_X1    g14724(.A1(new_n17663_), .A2(pi1153), .Z(new_n17674_));
  NAND2_X1   g14725(.A1(new_n17674_), .A2(new_n17673_), .ZN(new_n17675_));
  OAI21_X1   g14726(.A1(new_n17663_), .A2(new_n17654_), .B(new_n11893_), .ZN(new_n17676_));
  AOI21_X1   g14727(.A1(new_n17675_), .A2(new_n17676_), .B(new_n11891_), .ZN(new_n17677_));
  NOR2_X1    g14728(.A1(new_n17658_), .A2(pi0778), .ZN(new_n17678_));
  OAI21_X1   g14729(.A1(new_n17677_), .A2(new_n17678_), .B(pi0609), .ZN(new_n17679_));
  AOI21_X1   g14730(.A1(new_n17657_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n17680_));
  NOR2_X1    g14731(.A1(new_n17680_), .A2(pi0660), .ZN(new_n17681_));
  OAI21_X1   g14732(.A1(new_n17672_), .A2(new_n17679_), .B(new_n17681_), .ZN(new_n17682_));
  NOR2_X1    g14733(.A1(new_n17677_), .A2(new_n17678_), .ZN(new_n17683_));
  NAND4_X1   g14734(.A1(new_n17670_), .A2(pi0609), .A3(new_n11912_), .A4(new_n17683_), .ZN(new_n17684_));
  NOR2_X1    g14735(.A1(new_n17656_), .A2(new_n11925_), .ZN(new_n17685_));
  AOI21_X1   g14736(.A1(new_n17685_), .A2(new_n11928_), .B(pi1155), .ZN(new_n17686_));
  NOR2_X1    g14737(.A1(new_n17686_), .A2(new_n11923_), .ZN(new_n17687_));
  NAND2_X1   g14738(.A1(new_n17684_), .A2(new_n17687_), .ZN(new_n17688_));
  NAND3_X1   g14739(.A1(new_n17688_), .A2(pi0785), .A3(new_n17682_), .ZN(new_n17689_));
  NAND2_X1   g14740(.A1(new_n17689_), .A2(new_n17671_), .ZN(new_n17690_));
  NOR4_X1    g14741(.A1(new_n17683_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n17692_));
  NOR2_X1    g14742(.A1(new_n17685_), .A2(pi0785), .ZN(new_n17693_));
  OAI21_X1   g14743(.A1(new_n17686_), .A2(new_n17680_), .B(pi0785), .ZN(new_n17694_));
  XNOR2_X1   g14744(.A1(new_n17694_), .A2(new_n17693_), .ZN(new_n17695_));
  INV_X1     g14745(.I(new_n17695_), .ZN(new_n17696_));
  NOR2_X1    g14746(.A1(new_n17696_), .A2(new_n11945_), .ZN(new_n17697_));
  NOR3_X1    g14747(.A1(new_n17697_), .A2(pi0627), .A3(new_n17692_), .ZN(new_n17698_));
  AOI21_X1   g14748(.A1(new_n17695_), .A2(new_n11951_), .B(pi1154), .ZN(new_n17699_));
  NOR2_X1    g14749(.A1(new_n17683_), .A2(new_n11939_), .ZN(new_n17700_));
  INV_X1     g14750(.I(new_n17700_), .ZN(new_n17701_));
  NAND4_X1   g14751(.A1(new_n17690_), .A2(pi0618), .A3(new_n11950_), .A4(new_n17701_), .ZN(new_n17702_));
  NAND2_X1   g14752(.A1(new_n17702_), .A2(new_n17699_), .ZN(new_n17703_));
  AOI21_X1   g14753(.A1(new_n17703_), .A2(new_n11949_), .B(new_n17698_), .ZN(new_n17704_));
  NOR2_X1    g14754(.A1(new_n17704_), .A2(new_n11969_), .ZN(new_n17705_));
  AOI21_X1   g14755(.A1(new_n11969_), .A2(new_n17690_), .B(new_n17705_), .ZN(new_n17706_));
  NOR2_X1    g14756(.A1(new_n17701_), .A2(new_n11962_), .ZN(new_n17707_));
  NOR4_X1    g14757(.A1(new_n17706_), .A2(new_n11967_), .A3(pi1159), .A4(new_n17707_), .ZN(new_n17708_));
  INV_X1     g14758(.I(new_n17697_), .ZN(new_n17709_));
  NAND2_X1   g14759(.A1(new_n17709_), .A2(new_n17699_), .ZN(new_n17710_));
  MUX2_X1    g14760(.I0(new_n17710_), .I1(new_n17695_), .S(new_n11969_), .Z(new_n17711_));
  NAND2_X1   g14761(.A1(new_n17711_), .A2(pi0619), .ZN(new_n17712_));
  INV_X1     g14762(.I(new_n17712_), .ZN(new_n17713_));
  INV_X1     g14763(.I(new_n17654_), .ZN(new_n17714_));
  OAI21_X1   g14764(.A1(new_n17714_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n17715_));
  NOR4_X1    g14765(.A1(new_n17708_), .A2(new_n11966_), .A3(new_n17713_), .A4(new_n17715_), .ZN(new_n17716_));
  NOR4_X1    g14766(.A1(new_n17701_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n17717_));
  OAI21_X1   g14767(.A1(new_n17654_), .A2(pi0619), .B(new_n11869_), .ZN(new_n17718_));
  OAI21_X1   g14768(.A1(new_n17713_), .A2(new_n17718_), .B(new_n11966_), .ZN(new_n17719_));
  NOR2_X1    g14769(.A1(new_n17719_), .A2(new_n17717_), .ZN(new_n17720_));
  AOI21_X1   g14770(.A1(new_n17706_), .A2(new_n11998_), .B(pi0789), .ZN(new_n17721_));
  OAI21_X1   g14771(.A1(new_n17716_), .A2(new_n17720_), .B(new_n17721_), .ZN(new_n17722_));
  NAND2_X1   g14772(.A1(new_n17707_), .A2(new_n17450_), .ZN(new_n17723_));
  NOR2_X1    g14773(.A1(new_n17723_), .A2(new_n17153_), .ZN(new_n17724_));
  INV_X1     g14774(.I(new_n17724_), .ZN(new_n17725_));
  NOR2_X1    g14775(.A1(new_n17725_), .A2(new_n17151_), .ZN(new_n17726_));
  NOR2_X1    g14776(.A1(new_n14624_), .A2(new_n17654_), .ZN(new_n17727_));
  NAND3_X1   g14777(.A1(new_n17714_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n17728_));
  MUX2_X1    g14778(.I0(new_n17728_), .I1(new_n17711_), .S(new_n11985_), .Z(new_n17729_));
  AOI21_X1   g14779(.A1(new_n17729_), .A2(new_n14624_), .B(new_n17727_), .ZN(new_n17730_));
  AND2_X2    g14780(.A1(new_n17730_), .A2(new_n12064_), .Z(new_n17731_));
  OAI21_X1   g14781(.A1(new_n17731_), .A2(new_n17726_), .B(pi0629), .ZN(new_n17732_));
  NAND2_X1   g14782(.A1(new_n17730_), .A2(new_n12063_), .ZN(new_n17733_));
  NAND2_X1   g14783(.A1(new_n17724_), .A2(new_n15084_), .ZN(new_n17734_));
  NAND4_X1   g14784(.A1(new_n17732_), .A2(new_n15085_), .A3(new_n17733_), .A4(new_n17734_), .ZN(new_n17735_));
  MUX2_X1    g14785(.I0(new_n17729_), .I1(new_n17714_), .S(new_n11994_), .Z(new_n17736_));
  NOR2_X1    g14786(.A1(new_n17736_), .A2(new_n17167_), .ZN(new_n17737_));
  OAI21_X1   g14787(.A1(new_n17729_), .A2(new_n17654_), .B(pi0626), .ZN(new_n17738_));
  NOR2_X1    g14788(.A1(new_n17723_), .A2(new_n12020_), .ZN(new_n17739_));
  NOR2_X1    g14789(.A1(new_n17739_), .A2(pi0788), .ZN(new_n17740_));
  OAI21_X1   g14790(.A1(new_n17738_), .A2(new_n17171_), .B(new_n17740_), .ZN(new_n17741_));
  OAI21_X1   g14791(.A1(new_n17737_), .A2(new_n17741_), .B(new_n14732_), .ZN(new_n17742_));
  AOI21_X1   g14792(.A1(new_n17735_), .A2(new_n14726_), .B(new_n17742_), .ZN(new_n17743_));
  NAND3_X1   g14793(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n17654_), .ZN(new_n17744_));
  NOR2_X1    g14794(.A1(new_n17725_), .A2(new_n12068_), .ZN(new_n17745_));
  INV_X1     g14795(.I(new_n17745_), .ZN(new_n17746_));
  NAND2_X1   g14796(.A1(new_n17746_), .A2(pi0647), .ZN(new_n17747_));
  NAND2_X1   g14797(.A1(new_n17654_), .A2(pi0647), .ZN(new_n17748_));
  NAND3_X1   g14798(.A1(new_n17747_), .A2(new_n12049_), .A3(new_n17748_), .ZN(new_n17749_));
  NOR2_X1    g14799(.A1(new_n17714_), .A2(pi0647), .ZN(new_n17750_));
  AOI21_X1   g14800(.A1(new_n17745_), .A2(pi0647), .B(new_n17750_), .ZN(new_n17751_));
  NAND2_X1   g14801(.A1(new_n17751_), .A2(new_n12088_), .ZN(new_n17752_));
  NAND2_X1   g14802(.A1(new_n17752_), .A2(pi0787), .ZN(new_n17753_));
  AOI21_X1   g14803(.A1(pi0630), .A2(new_n17749_), .B(new_n17753_), .ZN(new_n17754_));
  AOI22_X1   g14804(.A1(new_n17722_), .A2(new_n17743_), .B1(new_n17744_), .B2(new_n17754_), .ZN(new_n17755_));
  NOR2_X1    g14805(.A1(new_n17755_), .A2(new_n12082_), .ZN(new_n17756_));
  NAND4_X1   g14806(.A1(new_n17747_), .A2(pi0787), .A3(new_n12049_), .A4(new_n17748_), .ZN(new_n17757_));
  OAI21_X1   g14807(.A1(pi0787), .A2(new_n17746_), .B(new_n17757_), .ZN(new_n17758_));
  NOR2_X1    g14808(.A1(new_n17758_), .A2(pi0644), .ZN(new_n17759_));
  OR3_X2     g14809(.A1(new_n17756_), .A2(pi0715), .A3(new_n17759_), .Z(new_n17760_));
  MUX2_X1    g14810(.I0(new_n17730_), .I1(new_n17654_), .S(new_n16841_), .Z(new_n17761_));
  INV_X1     g14811(.I(new_n17761_), .ZN(new_n17762_));
  OAI21_X1   g14812(.A1(new_n17761_), .A2(new_n17654_), .B(new_n12082_), .ZN(new_n17763_));
  AOI21_X1   g14813(.A1(new_n17654_), .A2(new_n17761_), .B(new_n17763_), .ZN(new_n17764_));
  OAI21_X1   g14814(.A1(new_n17764_), .A2(new_n17762_), .B(new_n12099_), .ZN(new_n17765_));
  AOI21_X1   g14815(.A1(new_n17762_), .A2(new_n17764_), .B(new_n17765_), .ZN(new_n17766_));
  AOI21_X1   g14816(.A1(new_n17760_), .A2(new_n17766_), .B(pi1160), .ZN(new_n17767_));
  XOR2_X1    g14817(.A1(new_n17764_), .A2(new_n17654_), .Z(new_n17768_));
  AOI21_X1   g14818(.A1(new_n17758_), .A2(pi0644), .B(new_n13169_), .ZN(new_n17769_));
  OAI21_X1   g14819(.A1(new_n17768_), .A2(new_n12099_), .B(new_n17769_), .ZN(new_n17770_));
  OAI21_X1   g14820(.A1(new_n17756_), .A2(new_n17770_), .B(pi0790), .ZN(new_n17771_));
  NOR2_X1    g14821(.A1(new_n17755_), .A2(new_n14748_), .ZN(new_n17772_));
  OAI21_X1   g14822(.A1(new_n17767_), .A2(new_n17771_), .B(new_n17772_), .ZN(new_n17773_));
  NOR2_X1    g14823(.A1(new_n3231_), .A2(pi0686), .ZN(new_n17774_));
  INV_X1     g14824(.I(new_n17774_), .ZN(new_n17775_));
  NOR2_X1    g14825(.A1(new_n12665_), .A2(pi0039), .ZN(new_n17776_));
  AOI21_X1   g14826(.A1(pi0039), .A2(new_n12349_), .B(new_n17776_), .ZN(new_n17777_));
  AOI21_X1   g14827(.A1(new_n17777_), .A2(new_n7620_), .B(pi0038), .ZN(new_n17778_));
  NAND2_X1   g14828(.A1(new_n12277_), .A2(pi0039), .ZN(new_n17779_));
  NAND2_X1   g14829(.A1(new_n12668_), .A2(new_n3154_), .ZN(new_n17780_));
  NAND3_X1   g14830(.A1(new_n17779_), .A2(pi0177), .A3(new_n17780_), .ZN(new_n17781_));
  NOR2_X1    g14831(.A1(new_n5157_), .A2(new_n12268_), .ZN(new_n17782_));
  INV_X1     g14832(.I(new_n17782_), .ZN(new_n17783_));
  NOR2_X1    g14833(.A1(new_n12122_), .A2(pi0039), .ZN(new_n17784_));
  MUX2_X1    g14834(.I0(new_n17784_), .I1(new_n17783_), .S(pi0177), .Z(new_n17785_));
  AOI21_X1   g14835(.A1(new_n17785_), .A2(pi0038), .B(pi0757), .ZN(new_n17786_));
  OAI21_X1   g14836(.A1(new_n17778_), .A2(new_n17781_), .B(new_n17786_), .ZN(new_n17787_));
  OAI21_X1   g14837(.A1(new_n13331_), .A2(new_n14344_), .B(new_n14342_), .ZN(new_n17788_));
  INV_X1     g14838(.I(new_n17788_), .ZN(new_n17789_));
  NOR2_X1    g14839(.A1(new_n12633_), .A2(pi0039), .ZN(new_n17790_));
  NOR2_X1    g14840(.A1(new_n12515_), .A2(new_n3154_), .ZN(new_n17791_));
  OAI21_X1   g14841(.A1(new_n17790_), .A2(new_n17791_), .B(pi0177), .ZN(new_n17792_));
  NAND2_X1   g14842(.A1(new_n13374_), .A2(new_n15787_), .ZN(new_n17793_));
  OAI21_X1   g14843(.A1(new_n17793_), .A2(new_n13368_), .B(new_n7620_), .ZN(new_n17794_));
  AOI21_X1   g14844(.A1(new_n17792_), .A2(new_n3172_), .B(new_n17794_), .ZN(new_n17795_));
  NAND2_X1   g14845(.A1(new_n17795_), .A2(new_n17789_), .ZN(new_n17796_));
  AOI21_X1   g14846(.A1(new_n17796_), .A2(new_n17787_), .B(new_n17775_), .ZN(new_n17797_));
  INV_X1     g14847(.I(new_n14360_), .ZN(new_n17798_));
  OAI21_X1   g14848(.A1(new_n14363_), .A2(new_n7620_), .B(new_n17798_), .ZN(new_n17799_));
  NAND2_X1   g14849(.A1(new_n12901_), .A2(new_n15787_), .ZN(new_n17800_));
  OAI22_X1   g14850(.A1(new_n14355_), .A2(new_n17800_), .B1(pi0757), .B2(new_n14365_), .ZN(new_n17801_));
  AOI22_X1   g14851(.A1(new_n17801_), .A2(new_n7620_), .B1(new_n15787_), .B2(new_n17799_), .ZN(new_n17802_));
  NAND2_X1   g14852(.A1(new_n17802_), .A2(pi0686), .ZN(new_n17803_));
  OAI22_X1   g14853(.A1(new_n17803_), .A2(new_n17797_), .B1(new_n7620_), .B2(new_n3231_), .ZN(new_n17804_));
  NOR2_X1    g14854(.A1(new_n3231_), .A2(pi0177), .ZN(new_n17805_));
  AOI21_X1   g14855(.A1(new_n17802_), .A2(new_n3231_), .B(new_n17805_), .ZN(new_n17806_));
  OAI21_X1   g14856(.A1(new_n17806_), .A2(pi0625), .B(pi1153), .ZN(new_n17807_));
  NOR2_X1    g14857(.A1(new_n3231_), .A2(new_n7620_), .ZN(new_n17808_));
  OAI21_X1   g14858(.A1(new_n12902_), .A2(pi0177), .B(new_n17774_), .ZN(new_n17809_));
  NOR3_X1    g14859(.A1(new_n13399_), .A2(pi0177), .A3(new_n13396_), .ZN(new_n17810_));
  AOI21_X1   g14860(.A1(new_n13399_), .A2(new_n7620_), .B(new_n13395_), .ZN(new_n17811_));
  NAND2_X1   g14861(.A1(new_n3172_), .A2(pi0686), .ZN(new_n17813_));
  NOR3_X1    g14862(.A1(new_n17810_), .A2(new_n17811_), .A3(new_n17813_), .ZN(new_n17814_));
  AOI21_X1   g14863(.A1(new_n17814_), .A2(new_n17809_), .B(new_n17808_), .ZN(new_n17815_));
  INV_X1     g14864(.I(new_n17815_), .ZN(new_n17816_));
  NOR2_X1    g14865(.A1(new_n12965_), .A2(pi0177), .ZN(new_n17817_));
  INV_X1     g14866(.I(new_n17817_), .ZN(new_n17818_));
  NOR4_X1    g14867(.A1(new_n17818_), .A2(pi0608), .A3(pi0625), .A4(pi1153), .ZN(new_n17819_));
  NAND2_X1   g14868(.A1(new_n17804_), .A2(pi0625), .ZN(new_n17820_));
  AOI21_X1   g14869(.A1(new_n17816_), .A2(new_n17819_), .B(new_n17820_), .ZN(new_n17821_));
  OAI21_X1   g14870(.A1(new_n17806_), .A2(new_n12970_), .B(new_n11893_), .ZN(new_n17822_));
  INV_X1     g14871(.I(new_n17804_), .ZN(new_n17823_));
  NOR3_X1    g14872(.A1(new_n17823_), .A2(pi0608), .A3(pi0625), .ZN(new_n17826_));
  AOI22_X1   g14873(.A1(new_n17821_), .A2(new_n17807_), .B1(new_n17826_), .B2(new_n17822_), .ZN(new_n17827_));
  NOR3_X1    g14874(.A1(new_n17827_), .A2(new_n11891_), .A3(new_n17804_), .ZN(new_n17828_));
  AOI21_X1   g14875(.A1(new_n17827_), .A2(pi0778), .B(new_n17823_), .ZN(new_n17829_));
  NOR2_X1    g14876(.A1(new_n17828_), .A2(new_n17829_), .ZN(new_n17830_));
  INV_X1     g14877(.I(new_n17830_), .ZN(new_n17831_));
  MUX2_X1    g14878(.I0(new_n17818_), .I1(new_n17815_), .S(new_n13435_), .Z(new_n17832_));
  NOR2_X1    g14879(.A1(new_n17832_), .A2(new_n11891_), .ZN(new_n17833_));
  AOI21_X1   g14880(.A1(new_n11891_), .A2(new_n17816_), .B(new_n17833_), .ZN(new_n17834_));
  OAI21_X1   g14881(.A1(new_n17834_), .A2(pi0609), .B(pi1155), .ZN(new_n17835_));
  NOR2_X1    g14882(.A1(new_n17817_), .A2(new_n12996_), .ZN(new_n17836_));
  INV_X1     g14883(.I(new_n17806_), .ZN(new_n17837_));
  NOR3_X1    g14884(.A1(new_n17837_), .A2(pi0609), .A3(new_n11914_), .ZN(new_n17838_));
  OAI21_X1   g14885(.A1(new_n17838_), .A2(new_n17836_), .B(new_n11912_), .ZN(new_n17839_));
  NAND2_X1   g14886(.A1(new_n17839_), .A2(pi0660), .ZN(new_n17840_));
  NAND3_X1   g14887(.A1(new_n17835_), .A2(pi0609), .A3(new_n17840_), .ZN(new_n17841_));
  NOR3_X1    g14888(.A1(new_n17828_), .A2(new_n17829_), .A3(pi0609), .ZN(new_n17842_));
  NOR2_X1    g14889(.A1(new_n17817_), .A2(new_n11915_), .ZN(new_n17843_));
  NOR3_X1    g14890(.A1(new_n17837_), .A2(new_n11903_), .A3(new_n11914_), .ZN(new_n17844_));
  NOR2_X1    g14891(.A1(new_n11923_), .A2(pi1155), .ZN(new_n17845_));
  OAI21_X1   g14892(.A1(new_n17834_), .A2(new_n11903_), .B(new_n17845_), .ZN(new_n17846_));
  OAI22_X1   g14893(.A1(new_n17831_), .A2(new_n17841_), .B1(new_n17842_), .B2(new_n17846_), .ZN(new_n17847_));
  MUX2_X1    g14894(.I0(new_n17847_), .I1(new_n17830_), .S(new_n11870_), .Z(new_n17848_));
  NAND2_X1   g14895(.A1(new_n17848_), .A2(new_n11969_), .ZN(new_n17849_));
  INV_X1     g14896(.I(new_n17834_), .ZN(new_n17850_));
  NOR2_X1    g14897(.A1(new_n17818_), .A2(new_n11938_), .ZN(new_n17851_));
  AOI21_X1   g14898(.A1(new_n17850_), .A2(new_n11938_), .B(new_n17851_), .ZN(new_n17852_));
  INV_X1     g14899(.I(new_n17852_), .ZN(new_n17853_));
  AOI21_X1   g14900(.A1(new_n17853_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n17854_));
  AOI21_X1   g14901(.A1(new_n17817_), .A2(new_n11914_), .B(pi0785), .ZN(new_n17855_));
  OAI21_X1   g14902(.A1(new_n17806_), .A2(new_n11914_), .B(new_n17855_), .ZN(new_n17856_));
  INV_X1     g14903(.I(new_n17856_), .ZN(new_n17857_));
  OAI21_X1   g14904(.A1(new_n17844_), .A2(new_n17843_), .B(pi1155), .ZN(new_n17858_));
  NAND2_X1   g14905(.A1(new_n17839_), .A2(new_n17858_), .ZN(new_n17859_));
  AND3_X2    g14906(.A1(new_n17859_), .A2(pi0785), .A3(new_n17857_), .Z(new_n17860_));
  AOI21_X1   g14907(.A1(new_n17859_), .A2(pi0785), .B(new_n17857_), .ZN(new_n17861_));
  NOR3_X1    g14908(.A1(new_n17860_), .A2(new_n11934_), .A3(new_n17861_), .ZN(new_n17862_));
  NOR2_X1    g14909(.A1(new_n17818_), .A2(new_n11934_), .ZN(new_n17863_));
  NOR4_X1    g14910(.A1(new_n17862_), .A2(new_n11949_), .A3(pi1154), .A4(new_n17863_), .ZN(new_n17864_));
  NOR3_X1    g14911(.A1(new_n17864_), .A2(new_n11934_), .A3(new_n17854_), .ZN(new_n17865_));
  NAND2_X1   g14912(.A1(new_n17848_), .A2(new_n11934_), .ZN(new_n17866_));
  NOR2_X1    g14913(.A1(new_n17817_), .A2(pi0618), .ZN(new_n17867_));
  OR3_X2     g14914(.A1(new_n17862_), .A2(pi1154), .A3(new_n17867_), .Z(new_n17868_));
  NAND2_X1   g14915(.A1(new_n17868_), .A2(new_n11949_), .ZN(new_n17869_));
  AOI21_X1   g14916(.A1(new_n17853_), .A2(pi0618), .B(pi1154), .ZN(new_n17870_));
  AND2_X2    g14917(.A1(new_n17869_), .A2(new_n17870_), .Z(new_n17871_));
  AOI22_X1   g14918(.A1(new_n17866_), .A2(new_n17871_), .B1(new_n17848_), .B2(new_n17865_), .ZN(new_n17872_));
  NOR3_X1    g14919(.A1(new_n17872_), .A2(new_n11969_), .A3(new_n17849_), .ZN(new_n17873_));
  INV_X1     g14920(.I(new_n17849_), .ZN(new_n17874_));
  NAND2_X1   g14921(.A1(new_n17848_), .A2(new_n17865_), .ZN(new_n17875_));
  NOR2_X1    g14922(.A1(new_n17831_), .A2(pi0785), .ZN(new_n17876_));
  NAND3_X1   g14923(.A1(new_n17847_), .A2(pi0785), .A3(new_n17876_), .ZN(new_n17877_));
  INV_X1     g14924(.I(new_n17877_), .ZN(new_n17878_));
  AOI21_X1   g14925(.A1(new_n17847_), .A2(pi0785), .B(new_n17876_), .ZN(new_n17879_));
  NOR3_X1    g14926(.A1(new_n17878_), .A2(new_n17879_), .A3(pi0618), .ZN(new_n17880_));
  INV_X1     g14927(.I(new_n17871_), .ZN(new_n17881_));
  OAI21_X1   g14928(.A1(new_n17881_), .A2(new_n17880_), .B(new_n17875_), .ZN(new_n17882_));
  AOI21_X1   g14929(.A1(new_n17882_), .A2(pi0781), .B(new_n17874_), .ZN(new_n17883_));
  NOR3_X1    g14930(.A1(new_n17883_), .A2(new_n17873_), .A3(pi0789), .ZN(new_n17884_));
  INV_X1     g14931(.I(new_n17884_), .ZN(new_n17885_));
  NOR2_X1    g14932(.A1(new_n17883_), .A2(new_n17873_), .ZN(new_n17886_));
  NOR2_X1    g14933(.A1(new_n17860_), .A2(new_n17861_), .ZN(new_n17887_));
  NAND3_X1   g14934(.A1(new_n17818_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n17888_));
  MUX2_X1    g14935(.I0(new_n17888_), .I1(new_n17887_), .S(new_n11969_), .Z(new_n17889_));
  NAND2_X1   g14936(.A1(new_n17889_), .A2(pi0619), .ZN(new_n17890_));
  AOI21_X1   g14937(.A1(new_n17817_), .A2(pi0619), .B(pi1159), .ZN(new_n17891_));
  AND3_X2    g14938(.A1(new_n17890_), .A2(pi0648), .A3(new_n17891_), .Z(new_n17892_));
  NOR2_X1    g14939(.A1(new_n17817_), .A2(new_n11961_), .ZN(new_n17893_));
  AOI21_X1   g14940(.A1(new_n17852_), .A2(new_n11961_), .B(new_n17893_), .ZN(new_n17894_));
  NOR3_X1    g14941(.A1(new_n17892_), .A2(new_n11967_), .A3(pi1159), .ZN(new_n17895_));
  NAND3_X1   g14942(.A1(new_n17882_), .A2(pi0781), .A3(new_n17874_), .ZN(new_n17896_));
  OAI21_X1   g14943(.A1(new_n17872_), .A2(new_n11969_), .B(new_n17849_), .ZN(new_n17897_));
  NAND3_X1   g14944(.A1(new_n17896_), .A2(new_n17897_), .A3(new_n11967_), .ZN(new_n17898_));
  AOI21_X1   g14945(.A1(new_n17818_), .A2(new_n11967_), .B(pi1159), .ZN(new_n17899_));
  NAND2_X1   g14946(.A1(new_n17890_), .A2(new_n17899_), .ZN(new_n17900_));
  NAND2_X1   g14947(.A1(new_n17900_), .A2(new_n11966_), .ZN(new_n17901_));
  AOI21_X1   g14948(.A1(new_n17894_), .A2(pi0619), .B(pi1159), .ZN(new_n17902_));
  NAND2_X1   g14949(.A1(new_n17901_), .A2(new_n17902_), .ZN(new_n17903_));
  INV_X1     g14950(.I(new_n17903_), .ZN(new_n17904_));
  AOI22_X1   g14951(.A1(new_n17898_), .A2(new_n17904_), .B1(new_n17886_), .B2(new_n17895_), .ZN(new_n17905_));
  NOR3_X1    g14952(.A1(new_n17905_), .A2(new_n11985_), .A3(new_n17885_), .ZN(new_n17906_));
  NAND3_X1   g14953(.A1(new_n17896_), .A2(new_n17897_), .A3(new_n17895_), .ZN(new_n17907_));
  NOR3_X1    g14954(.A1(new_n17883_), .A2(new_n17873_), .A3(pi0619), .ZN(new_n17908_));
  OAI21_X1   g14955(.A1(new_n17908_), .A2(new_n17903_), .B(new_n17907_), .ZN(new_n17909_));
  AOI21_X1   g14956(.A1(new_n17909_), .A2(pi0789), .B(new_n17884_), .ZN(new_n17910_));
  NOR2_X1    g14957(.A1(new_n17906_), .A2(new_n17910_), .ZN(new_n17911_));
  NAND3_X1   g14958(.A1(new_n17909_), .A2(pi0789), .A3(new_n17884_), .ZN(new_n17912_));
  OAI21_X1   g14959(.A1(new_n17905_), .A2(new_n11985_), .B(new_n17885_), .ZN(new_n17913_));
  NAND2_X1   g14960(.A1(new_n17889_), .A2(new_n11985_), .ZN(new_n17914_));
  NOR3_X1    g14961(.A1(new_n17817_), .A2(pi0619), .A3(pi1159), .ZN(new_n17915_));
  NOR2_X1    g14962(.A1(new_n17915_), .A2(new_n11985_), .ZN(new_n17916_));
  XNOR2_X1   g14963(.A1(new_n17914_), .A2(new_n17916_), .ZN(new_n17917_));
  NOR3_X1    g14964(.A1(new_n11994_), .A2(new_n11989_), .A3(pi1158), .ZN(new_n17918_));
  NAND2_X1   g14965(.A1(new_n17917_), .A2(new_n17918_), .ZN(new_n17919_));
  NOR2_X1    g14966(.A1(new_n17818_), .A2(new_n12014_), .ZN(new_n17920_));
  AOI21_X1   g14967(.A1(new_n17894_), .A2(new_n12014_), .B(new_n17920_), .ZN(new_n17921_));
  NOR2_X1    g14968(.A1(new_n11994_), .A2(pi0641), .ZN(new_n17922_));
  NAND2_X1   g14969(.A1(new_n17919_), .A2(new_n17922_), .ZN(new_n17923_));
  INV_X1     g14970(.I(new_n17917_), .ZN(new_n17924_));
  NOR2_X1    g14971(.A1(new_n17924_), .A2(pi0626), .ZN(new_n17925_));
  OAI21_X1   g14972(.A1(new_n17817_), .A2(new_n11994_), .B(pi0641), .ZN(new_n17926_));
  NOR3_X1    g14973(.A1(new_n11989_), .A2(pi0626), .A3(pi1158), .ZN(new_n17927_));
  OAI21_X1   g14974(.A1(new_n17925_), .A2(new_n17926_), .B(new_n17927_), .ZN(new_n17928_));
  AOI22_X1   g14975(.A1(new_n17913_), .A2(new_n17912_), .B1(new_n17923_), .B2(new_n17928_), .ZN(new_n17929_));
  NAND3_X1   g14976(.A1(new_n17929_), .A2(pi0788), .A3(new_n17911_), .ZN(new_n17930_));
  NAND2_X1   g14977(.A1(new_n17913_), .A2(new_n17912_), .ZN(new_n17931_));
  OAI21_X1   g14978(.A1(new_n17929_), .A2(new_n11986_), .B(new_n17931_), .ZN(new_n17932_));
  NAND2_X1   g14979(.A1(new_n17932_), .A2(new_n17930_), .ZN(new_n17933_));
  INV_X1     g14980(.I(new_n17923_), .ZN(new_n17934_));
  INV_X1     g14981(.I(new_n17928_), .ZN(new_n17935_));
  OAI22_X1   g14982(.A1(new_n17906_), .A2(new_n17910_), .B1(new_n17934_), .B2(new_n17935_), .ZN(new_n17936_));
  NOR3_X1    g14983(.A1(new_n17936_), .A2(new_n11986_), .A3(new_n17931_), .ZN(new_n17937_));
  AOI21_X1   g14984(.A1(new_n17936_), .A2(pi0788), .B(new_n17911_), .ZN(new_n17938_));
  NOR2_X1    g14985(.A1(new_n17924_), .A2(new_n11997_), .ZN(new_n17939_));
  AOI21_X1   g14986(.A1(new_n11997_), .A2(new_n17818_), .B(new_n17939_), .ZN(new_n17940_));
  INV_X1     g14987(.I(new_n17940_), .ZN(new_n17941_));
  OAI21_X1   g14988(.A1(new_n17941_), .A2(pi0628), .B(pi1156), .ZN(new_n17942_));
  NOR2_X1    g14989(.A1(new_n17817_), .A2(new_n13114_), .ZN(new_n17943_));
  AOI21_X1   g14990(.A1(new_n17921_), .A2(new_n13114_), .B(new_n17943_), .ZN(new_n17944_));
  NOR3_X1    g14991(.A1(new_n17818_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n17945_));
  NOR2_X1    g14992(.A1(new_n17945_), .A2(new_n12030_), .ZN(new_n17946_));
  NOR2_X1    g14993(.A1(new_n17946_), .A2(new_n12031_), .ZN(new_n17947_));
  NAND2_X1   g14994(.A1(new_n17942_), .A2(new_n17947_), .ZN(new_n17948_));
  INV_X1     g14995(.I(new_n17948_), .ZN(new_n17949_));
  NOR2_X1    g14996(.A1(new_n17941_), .A2(new_n12031_), .ZN(new_n17950_));
  NOR2_X1    g14997(.A1(new_n12030_), .A2(pi0628), .ZN(new_n17951_));
  OAI21_X1   g14998(.A1(new_n17950_), .A2(pi1156), .B(new_n17951_), .ZN(new_n17952_));
  INV_X1     g14999(.I(new_n17952_), .ZN(new_n17953_));
  OAI22_X1   g15000(.A1(new_n17937_), .A2(new_n17938_), .B1(new_n17949_), .B2(new_n17953_), .ZN(new_n17954_));
  NOR3_X1    g15001(.A1(new_n17954_), .A2(new_n11868_), .A3(new_n17933_), .ZN(new_n17955_));
  NOR2_X1    g15002(.A1(new_n17937_), .A2(new_n17938_), .ZN(new_n17956_));
  AOI21_X1   g15003(.A1(new_n17954_), .A2(pi0792), .B(new_n17956_), .ZN(new_n17957_));
  NOR2_X1    g15004(.A1(new_n17955_), .A2(new_n17957_), .ZN(new_n17958_));
  AOI22_X1   g15005(.A1(new_n17932_), .A2(new_n17930_), .B1(new_n17948_), .B2(new_n17952_), .ZN(new_n17959_));
  NAND3_X1   g15006(.A1(new_n17959_), .A2(pi0792), .A3(new_n17956_), .ZN(new_n17960_));
  OAI21_X1   g15007(.A1(new_n17959_), .A2(new_n11868_), .B(new_n17933_), .ZN(new_n17961_));
  NAND2_X1   g15008(.A1(new_n17961_), .A2(new_n17960_), .ZN(new_n17962_));
  NOR4_X1    g15009(.A1(new_n17944_), .A2(new_n12031_), .A3(pi1156), .A4(new_n17817_), .ZN(new_n17963_));
  NOR2_X1    g15010(.A1(new_n17963_), .A2(new_n17945_), .ZN(new_n17964_));
  MUX2_X1    g15011(.I0(new_n17964_), .I1(new_n17944_), .S(new_n11868_), .Z(new_n17965_));
  NAND2_X1   g15012(.A1(new_n17965_), .A2(pi0647), .ZN(new_n17966_));
  AOI21_X1   g15013(.A1(new_n17817_), .A2(pi0647), .B(pi1157), .ZN(new_n17967_));
  NAND2_X1   g15014(.A1(new_n17966_), .A2(new_n17967_), .ZN(new_n17968_));
  NOR2_X1    g15015(.A1(new_n17817_), .A2(new_n12054_), .ZN(new_n17969_));
  AOI21_X1   g15016(.A1(new_n17941_), .A2(new_n12054_), .B(new_n17969_), .ZN(new_n17970_));
  NOR2_X1    g15017(.A1(new_n12061_), .A2(pi1157), .ZN(new_n17971_));
  OAI21_X1   g15018(.A1(new_n17968_), .A2(new_n12060_), .B(new_n17971_), .ZN(new_n17972_));
  NOR3_X1    g15019(.A1(new_n17955_), .A2(new_n17957_), .A3(pi0647), .ZN(new_n17973_));
  AOI21_X1   g15020(.A1(new_n17818_), .A2(new_n12061_), .B(pi1157), .ZN(new_n17974_));
  NAND2_X1   g15021(.A1(new_n17966_), .A2(new_n17974_), .ZN(new_n17975_));
  NAND2_X1   g15022(.A1(new_n17975_), .A2(new_n12060_), .ZN(new_n17976_));
  AOI21_X1   g15023(.A1(new_n17970_), .A2(pi0647), .B(pi1157), .ZN(new_n17977_));
  AND2_X2    g15024(.A1(new_n17977_), .A2(new_n17976_), .Z(new_n17978_));
  INV_X1     g15025(.I(new_n17978_), .ZN(new_n17979_));
  OAI22_X1   g15026(.A1(new_n17973_), .A2(new_n17979_), .B1(new_n17962_), .B2(new_n17972_), .ZN(new_n17980_));
  MUX2_X1    g15027(.I0(new_n17980_), .I1(new_n17958_), .S(new_n12048_), .Z(new_n17981_));
  INV_X1     g15028(.I(new_n17965_), .ZN(new_n17982_));
  NOR3_X1    g15029(.A1(new_n17817_), .A2(pi0647), .A3(pi1157), .ZN(new_n17983_));
  MUX2_X1    g15030(.I0(new_n17983_), .I1(new_n17982_), .S(new_n12048_), .Z(new_n17984_));
  NAND2_X1   g15031(.A1(new_n17984_), .A2(pi0644), .ZN(new_n17985_));
  NOR2_X1    g15032(.A1(new_n17818_), .A2(new_n12092_), .ZN(new_n17986_));
  AOI21_X1   g15033(.A1(new_n17970_), .A2(new_n12092_), .B(new_n17986_), .ZN(new_n17987_));
  NAND2_X1   g15034(.A1(new_n12082_), .A2(new_n12099_), .ZN(new_n17988_));
  OR2_X2     g15035(.A1(new_n17987_), .A2(new_n17988_), .Z(new_n17989_));
  NAND3_X1   g15036(.A1(new_n17989_), .A2(new_n13168_), .A3(new_n17985_), .ZN(new_n17990_));
  AOI21_X1   g15037(.A1(new_n17981_), .A2(new_n12082_), .B(new_n17990_), .ZN(new_n17991_));
  INV_X1     g15038(.I(new_n17972_), .ZN(new_n17992_));
  NAND3_X1   g15039(.A1(new_n17961_), .A2(new_n17960_), .A3(new_n12061_), .ZN(new_n17993_));
  AOI22_X1   g15040(.A1(new_n17993_), .A2(new_n17978_), .B1(new_n17958_), .B2(new_n17992_), .ZN(new_n17994_));
  MUX2_X1    g15041(.I0(new_n17994_), .I1(new_n17962_), .S(new_n12048_), .Z(new_n17995_));
  NAND3_X1   g15042(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n17996_));
  OAI21_X1   g15043(.A1(new_n17987_), .A2(new_n17996_), .B(new_n13179_), .ZN(new_n17997_));
  NOR2_X1    g15044(.A1(new_n17997_), .A2(new_n17984_), .ZN(new_n17998_));
  OAI21_X1   g15045(.A1(new_n17995_), .A2(new_n12082_), .B(new_n17998_), .ZN(new_n17999_));
  NOR2_X1    g15046(.A1(new_n17999_), .A2(new_n17991_), .ZN(new_n18000_));
  NAND2_X1   g15047(.A1(po1038), .A2(new_n7620_), .ZN(new_n18001_));
  AOI21_X1   g15048(.A1(new_n18001_), .A2(new_n13184_), .B(po1038), .ZN(new_n18002_));
  OAI21_X1   g15049(.A1(new_n17981_), .A2(pi0790), .B(new_n18002_), .ZN(new_n18003_));
  OAI21_X1   g15050(.A1(new_n18000_), .A2(new_n18003_), .B(new_n17773_), .ZN(po0334));
  NOR2_X1    g15051(.A1(new_n2925_), .A2(pi0178), .ZN(new_n18005_));
  NOR2_X1    g15052(.A1(new_n11877_), .A2(pi0760), .ZN(new_n18006_));
  NOR2_X1    g15053(.A1(new_n18006_), .A2(new_n18005_), .ZN(new_n18007_));
  AOI21_X1   g15054(.A1(new_n11886_), .A2(new_n15830_), .B(new_n18005_), .ZN(new_n18008_));
  NOR2_X1    g15055(.A1(new_n18008_), .A2(new_n11874_), .ZN(new_n18009_));
  INV_X1     g15056(.I(new_n18009_), .ZN(new_n18010_));
  NAND2_X1   g15057(.A1(new_n18010_), .A2(new_n18007_), .ZN(new_n18011_));
  NAND2_X1   g15058(.A1(new_n18011_), .A2(new_n11891_), .ZN(new_n18012_));
  NOR2_X1    g15059(.A1(new_n18010_), .A2(new_n12970_), .ZN(new_n18013_));
  NOR4_X1    g15060(.A1(new_n18013_), .A2(new_n11893_), .A3(new_n18005_), .A4(new_n18006_), .ZN(new_n18014_));
  NOR3_X1    g15061(.A1(new_n11894_), .A2(pi0625), .A3(pi0688), .ZN(new_n18015_));
  NOR2_X1    g15062(.A1(new_n18005_), .A2(pi1153), .ZN(new_n18016_));
  INV_X1     g15063(.I(new_n18016_), .ZN(new_n18017_));
  NOR2_X1    g15064(.A1(new_n18015_), .A2(new_n18017_), .ZN(new_n18018_));
  INV_X1     g15065(.I(new_n18018_), .ZN(new_n18019_));
  NAND2_X1   g15066(.A1(new_n18019_), .A2(pi0608), .ZN(new_n18020_));
  INV_X1     g15067(.I(new_n18013_), .ZN(new_n18021_));
  AOI21_X1   g15068(.A1(new_n18021_), .A2(new_n18011_), .B(new_n18017_), .ZN(new_n18022_));
  OAI21_X1   g15069(.A1(new_n18015_), .A2(new_n18008_), .B(pi1153), .ZN(new_n18023_));
  NAND2_X1   g15070(.A1(new_n18023_), .A2(new_n13657_), .ZN(new_n18024_));
  OAI22_X1   g15071(.A1(new_n18022_), .A2(new_n18024_), .B1(new_n18014_), .B2(new_n18020_), .ZN(new_n18025_));
  NAND2_X1   g15072(.A1(new_n18025_), .A2(pi0778), .ZN(new_n18026_));
  XOR2_X1    g15073(.A1(new_n18026_), .A2(new_n18012_), .Z(new_n18027_));
  INV_X1     g15074(.I(new_n18027_), .ZN(new_n18028_));
  NAND2_X1   g15075(.A1(new_n18019_), .A2(new_n18023_), .ZN(new_n18029_));
  MUX2_X1    g15076(.I0(new_n18029_), .I1(new_n18008_), .S(new_n11891_), .Z(new_n18030_));
  XNOR2_X1   g15077(.A1(new_n18027_), .A2(new_n18030_), .ZN(new_n18031_));
  NAND2_X1   g15078(.A1(new_n18031_), .A2(pi0609), .ZN(new_n18032_));
  XOR2_X1    g15079(.A1(new_n18032_), .A2(new_n18027_), .Z(new_n18033_));
  NAND2_X1   g15080(.A1(new_n18033_), .A2(new_n11912_), .ZN(new_n18034_));
  NOR2_X1    g15081(.A1(new_n18007_), .A2(new_n11925_), .ZN(new_n18035_));
  INV_X1     g15082(.I(new_n18035_), .ZN(new_n18036_));
  NOR3_X1    g15083(.A1(new_n12997_), .A2(new_n11877_), .A3(pi0760), .ZN(new_n18037_));
  NAND3_X1   g15084(.A1(new_n18036_), .A2(new_n11912_), .A3(new_n18037_), .ZN(new_n18038_));
  NAND3_X1   g15085(.A1(new_n18034_), .A2(new_n11923_), .A3(new_n18038_), .ZN(new_n18039_));
  NOR4_X1    g15086(.A1(new_n18037_), .A2(new_n11923_), .A3(pi1155), .A4(new_n18005_), .ZN(new_n18041_));
  NOR2_X1    g15087(.A1(new_n18041_), .A2(new_n11870_), .ZN(new_n18042_));
  AOI22_X1   g15088(.A1(new_n18039_), .A2(new_n18042_), .B1(new_n11870_), .B2(new_n18028_), .ZN(new_n18043_));
  NOR2_X1    g15089(.A1(new_n18043_), .A2(pi0781), .ZN(new_n18044_));
  NOR4_X1    g15090(.A1(new_n18030_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n18045_));
  NOR3_X1    g15091(.A1(new_n18037_), .A2(pi1155), .A3(new_n18005_), .ZN(new_n18046_));
  NAND2_X1   g15092(.A1(new_n18038_), .A2(new_n18046_), .ZN(new_n18047_));
  MUX2_X1    g15093(.I0(new_n18047_), .I1(new_n18036_), .S(new_n11870_), .Z(new_n18048_));
  INV_X1     g15094(.I(new_n18048_), .ZN(new_n18049_));
  OAI21_X1   g15095(.A1(new_n18049_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n18050_));
  OAI21_X1   g15096(.A1(new_n18049_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n18051_));
  NOR2_X1    g15097(.A1(new_n18030_), .A2(new_n11939_), .ZN(new_n18052_));
  NOR4_X1    g15098(.A1(new_n18043_), .A2(new_n11934_), .A3(pi1154), .A4(new_n18052_), .ZN(new_n18053_));
  NOR2_X1    g15099(.A1(new_n18053_), .A2(new_n18051_), .ZN(new_n18054_));
  OAI22_X1   g15100(.A1(new_n18054_), .A2(pi0627), .B1(new_n18045_), .B2(new_n18050_), .ZN(new_n18055_));
  AOI21_X1   g15101(.A1(new_n18055_), .A2(pi0781), .B(new_n18044_), .ZN(new_n18056_));
  INV_X1     g15102(.I(new_n18052_), .ZN(new_n18057_));
  NOR2_X1    g15103(.A1(new_n18057_), .A2(new_n11962_), .ZN(new_n18058_));
  NOR4_X1    g15104(.A1(new_n18056_), .A2(new_n11967_), .A3(pi1159), .A4(new_n18058_), .ZN(new_n18059_));
  NOR2_X1    g15105(.A1(new_n18049_), .A2(pi0781), .ZN(new_n18060_));
  AOI21_X1   g15106(.A1(new_n11944_), .A2(new_n18048_), .B(new_n18051_), .ZN(new_n18061_));
  NOR2_X1    g15107(.A1(new_n18061_), .A2(new_n11969_), .ZN(new_n18062_));
  XOR2_X1    g15108(.A1(new_n18062_), .A2(new_n18060_), .Z(new_n18063_));
  AOI21_X1   g15109(.A1(new_n18063_), .A2(new_n16479_), .B(pi1159), .ZN(new_n18064_));
  INV_X1     g15110(.I(new_n18064_), .ZN(new_n18065_));
  NOR3_X1    g15111(.A1(new_n18059_), .A2(new_n11966_), .A3(new_n18065_), .ZN(new_n18066_));
  NOR4_X1    g15112(.A1(new_n18057_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n18067_));
  INV_X1     g15113(.I(new_n18063_), .ZN(new_n18068_));
  NOR2_X1    g15114(.A1(new_n18068_), .A2(new_n16482_), .ZN(new_n18069_));
  NOR3_X1    g15115(.A1(new_n18069_), .A2(pi0648), .A3(new_n18067_), .ZN(new_n18070_));
  AOI21_X1   g15116(.A1(new_n18056_), .A2(new_n11998_), .B(pi0789), .ZN(new_n18071_));
  OAI21_X1   g15117(.A1(new_n18066_), .A2(new_n18070_), .B(new_n18071_), .ZN(new_n18072_));
  NAND2_X1   g15118(.A1(new_n18058_), .A2(new_n17450_), .ZN(new_n18073_));
  NOR2_X1    g15119(.A1(new_n18073_), .A2(new_n17153_), .ZN(new_n18074_));
  NOR2_X1    g15120(.A1(new_n14624_), .A2(new_n18005_), .ZN(new_n18075_));
  NOR2_X1    g15121(.A1(new_n18068_), .A2(pi0789), .ZN(new_n18076_));
  NOR2_X1    g15122(.A1(new_n18065_), .A2(new_n18069_), .ZN(new_n18077_));
  NOR2_X1    g15123(.A1(new_n18077_), .A2(new_n11985_), .ZN(new_n18078_));
  XOR2_X1    g15124(.A1(new_n18078_), .A2(new_n18076_), .Z(new_n18079_));
  AOI21_X1   g15125(.A1(new_n18079_), .A2(new_n14624_), .B(new_n18075_), .ZN(new_n18080_));
  AOI22_X1   g15126(.A1(new_n18080_), .A2(new_n12064_), .B1(new_n15080_), .B2(new_n18074_), .ZN(new_n18081_));
  NOR2_X1    g15127(.A1(new_n18081_), .A2(new_n12030_), .ZN(new_n18082_));
  NAND2_X1   g15128(.A1(new_n18080_), .A2(new_n12063_), .ZN(new_n18083_));
  AOI21_X1   g15129(.A1(new_n18074_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n18084_));
  NAND2_X1   g15130(.A1(new_n18083_), .A2(new_n18084_), .ZN(new_n18085_));
  OAI21_X1   g15131(.A1(new_n18082_), .A2(new_n18085_), .B(new_n14726_), .ZN(new_n18086_));
  INV_X1     g15132(.I(new_n18005_), .ZN(new_n18087_));
  MUX2_X1    g15133(.I0(new_n18079_), .I1(new_n18087_), .S(new_n11994_), .Z(new_n18088_));
  INV_X1     g15134(.I(new_n18079_), .ZN(new_n18089_));
  AOI21_X1   g15135(.A1(new_n18089_), .A2(new_n18087_), .B(new_n11994_), .ZN(new_n18090_));
  OAI21_X1   g15136(.A1(new_n18073_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n18091_));
  AOI21_X1   g15137(.A1(new_n18090_), .A2(new_n11990_), .B(new_n18091_), .ZN(new_n18092_));
  OAI21_X1   g15138(.A1(new_n17167_), .A2(new_n18088_), .B(new_n18092_), .ZN(new_n18093_));
  NAND4_X1   g15139(.A1(new_n18072_), .A2(new_n14732_), .A3(new_n18086_), .A4(new_n18093_), .ZN(new_n18094_));
  NAND3_X1   g15140(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n18005_), .ZN(new_n18095_));
  NAND2_X1   g15141(.A1(new_n18074_), .A2(new_n15050_), .ZN(new_n18096_));
  NAND2_X1   g15142(.A1(new_n18096_), .A2(pi0647), .ZN(new_n18097_));
  NAND2_X1   g15143(.A1(new_n18005_), .A2(pi0647), .ZN(new_n18098_));
  NAND3_X1   g15144(.A1(new_n18097_), .A2(new_n12049_), .A3(new_n18098_), .ZN(new_n18099_));
  NAND2_X1   g15145(.A1(new_n18099_), .A2(pi0630), .ZN(new_n18100_));
  NOR2_X1    g15146(.A1(new_n18096_), .A2(new_n12061_), .ZN(new_n18101_));
  AOI21_X1   g15147(.A1(new_n12061_), .A2(new_n18005_), .B(new_n18101_), .ZN(new_n18102_));
  NAND2_X1   g15148(.A1(new_n18102_), .A2(new_n12088_), .ZN(new_n18103_));
  NAND4_X1   g15149(.A1(new_n18103_), .A2(new_n18100_), .A3(pi0787), .A4(new_n18095_), .ZN(new_n18104_));
  AND2_X2    g15150(.A1(new_n18094_), .A2(new_n18104_), .Z(new_n18105_));
  NOR2_X1    g15151(.A1(new_n18105_), .A2(new_n12082_), .ZN(new_n18106_));
  NAND4_X1   g15152(.A1(new_n18097_), .A2(pi0787), .A3(new_n12049_), .A4(new_n18098_), .ZN(new_n18107_));
  OAI21_X1   g15153(.A1(pi0787), .A2(new_n18096_), .B(new_n18107_), .ZN(new_n18108_));
  NOR2_X1    g15154(.A1(new_n18108_), .A2(pi0644), .ZN(new_n18109_));
  OR3_X2     g15155(.A1(new_n18106_), .A2(pi0715), .A3(new_n18109_), .Z(new_n18110_));
  MUX2_X1    g15156(.I0(new_n18080_), .I1(new_n18005_), .S(new_n16841_), .Z(new_n18111_));
  INV_X1     g15157(.I(new_n18111_), .ZN(new_n18112_));
  OAI21_X1   g15158(.A1(new_n18111_), .A2(new_n18005_), .B(new_n12082_), .ZN(new_n18113_));
  AOI21_X1   g15159(.A1(new_n18005_), .A2(new_n18111_), .B(new_n18113_), .ZN(new_n18114_));
  OAI21_X1   g15160(.A1(new_n18114_), .A2(new_n18112_), .B(new_n12099_), .ZN(new_n18115_));
  AOI21_X1   g15161(.A1(new_n18112_), .A2(new_n18114_), .B(new_n18115_), .ZN(new_n18116_));
  AOI21_X1   g15162(.A1(new_n18110_), .A2(new_n18116_), .B(pi1160), .ZN(new_n18117_));
  XOR2_X1    g15163(.A1(new_n18114_), .A2(new_n18005_), .Z(new_n18118_));
  AOI21_X1   g15164(.A1(new_n18108_), .A2(pi0644), .B(new_n13169_), .ZN(new_n18119_));
  OAI21_X1   g15165(.A1(new_n18118_), .A2(new_n12099_), .B(new_n18119_), .ZN(new_n18120_));
  OAI21_X1   g15166(.A1(new_n18106_), .A2(new_n18120_), .B(pi0790), .ZN(new_n18121_));
  NOR2_X1    g15167(.A1(new_n18105_), .A2(new_n14748_), .ZN(new_n18122_));
  OAI21_X1   g15168(.A1(new_n18117_), .A2(new_n18121_), .B(new_n18122_), .ZN(new_n18123_));
  NOR2_X1    g15169(.A1(new_n12965_), .A2(pi0178), .ZN(new_n18124_));
  INV_X1     g15170(.I(new_n18124_), .ZN(new_n18125_));
  NAND2_X1   g15171(.A1(new_n18125_), .A2(new_n11997_), .ZN(new_n18126_));
  AOI21_X1   g15172(.A1(new_n12794_), .A2(new_n7345_), .B(pi0760), .ZN(new_n18127_));
  NAND3_X1   g15173(.A1(new_n13381_), .A2(new_n7345_), .A3(new_n14362_), .ZN(new_n18128_));
  OAI21_X1   g15174(.A1(new_n13381_), .A2(pi0178), .B(new_n12694_), .ZN(new_n18129_));
  NAND3_X1   g15175(.A1(new_n18129_), .A2(new_n18128_), .A3(new_n15831_), .ZN(new_n18130_));
  NOR2_X1    g15176(.A1(new_n18130_), .A2(new_n18127_), .ZN(new_n18131_));
  NOR2_X1    g15177(.A1(new_n12828_), .A2(pi0178), .ZN(new_n18132_));
  OAI21_X1   g15178(.A1(new_n13367_), .A2(pi0760), .B(pi0038), .ZN(new_n18133_));
  OAI22_X1   g15179(.A1(new_n18131_), .A2(pi0038), .B1(new_n18132_), .B2(new_n18133_), .ZN(new_n18134_));
  NOR2_X1    g15180(.A1(new_n18134_), .A2(new_n3232_), .ZN(new_n18135_));
  AOI21_X1   g15181(.A1(new_n7345_), .A2(new_n3232_), .B(new_n18135_), .ZN(new_n18136_));
  INV_X1     g15182(.I(new_n18136_), .ZN(new_n18137_));
  OAI21_X1   g15183(.A1(new_n18125_), .A2(new_n11924_), .B(new_n11870_), .ZN(new_n18138_));
  AOI21_X1   g15184(.A1(new_n18137_), .A2(new_n11924_), .B(new_n18138_), .ZN(new_n18139_));
  NAND2_X1   g15185(.A1(new_n18136_), .A2(new_n11924_), .ZN(new_n18140_));
  OAI22_X1   g15186(.A1(new_n18140_), .A2(pi0609), .B1(new_n12996_), .B2(new_n18124_), .ZN(new_n18141_));
  NAND2_X1   g15187(.A1(new_n18141_), .A2(new_n11912_), .ZN(new_n18142_));
  OAI22_X1   g15188(.A1(new_n18140_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n18124_), .ZN(new_n18143_));
  NAND2_X1   g15189(.A1(new_n18143_), .A2(pi1155), .ZN(new_n18144_));
  AOI21_X1   g15190(.A1(new_n18142_), .A2(new_n18144_), .B(new_n11870_), .ZN(new_n18145_));
  XOR2_X1    g15191(.A1(new_n18145_), .A2(new_n18139_), .Z(new_n18146_));
  OAI21_X1   g15192(.A1(new_n18125_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n18147_));
  AOI21_X1   g15193(.A1(new_n18146_), .A2(pi0618), .B(new_n18147_), .ZN(new_n18148_));
  NAND2_X1   g15194(.A1(new_n18146_), .A2(pi0618), .ZN(new_n18149_));
  AOI21_X1   g15195(.A1(new_n18125_), .A2(new_n11934_), .B(pi1154), .ZN(new_n18150_));
  NAND2_X1   g15196(.A1(new_n18149_), .A2(new_n18150_), .ZN(new_n18151_));
  NAND2_X1   g15197(.A1(new_n18151_), .A2(new_n18148_), .ZN(new_n18152_));
  MUX2_X1    g15198(.I0(new_n18152_), .I1(new_n18146_), .S(new_n11969_), .Z(new_n18153_));
  NAND2_X1   g15199(.A1(new_n18153_), .A2(new_n11985_), .ZN(new_n18154_));
  NOR3_X1    g15200(.A1(new_n18124_), .A2(pi0619), .A3(pi1159), .ZN(new_n18155_));
  NOR2_X1    g15201(.A1(new_n18155_), .A2(new_n11985_), .ZN(new_n18156_));
  XOR2_X1    g15202(.A1(new_n18154_), .A2(new_n18156_), .Z(new_n18157_));
  OAI21_X1   g15203(.A1(new_n18157_), .A2(new_n11997_), .B(new_n18126_), .ZN(new_n18158_));
  NOR2_X1    g15204(.A1(new_n18124_), .A2(new_n12054_), .ZN(new_n18159_));
  AOI21_X1   g15205(.A1(new_n18158_), .A2(new_n12054_), .B(new_n18159_), .ZN(new_n18160_));
  NAND2_X1   g15206(.A1(new_n18125_), .A2(new_n12091_), .ZN(new_n18161_));
  OAI21_X1   g15207(.A1(new_n18160_), .A2(new_n12091_), .B(new_n18161_), .ZN(new_n18162_));
  AOI21_X1   g15208(.A1(new_n18124_), .A2(pi0644), .B(new_n12099_), .ZN(new_n18163_));
  OAI21_X1   g15209(.A1(new_n18162_), .A2(pi0644), .B(new_n18163_), .ZN(new_n18164_));
  AND2_X2    g15210(.A1(new_n18164_), .A2(new_n12081_), .Z(new_n18165_));
  NOR2_X1    g15211(.A1(new_n18125_), .A2(pi0647), .ZN(new_n18166_));
  NOR2_X1    g15212(.A1(new_n18124_), .A2(new_n13114_), .ZN(new_n18167_));
  NOR2_X1    g15213(.A1(new_n18125_), .A2(new_n12014_), .ZN(new_n18168_));
  NOR2_X1    g15214(.A1(new_n18124_), .A2(new_n11961_), .ZN(new_n18169_));
  OAI21_X1   g15215(.A1(new_n15189_), .A2(new_n18132_), .B(new_n15830_), .ZN(new_n18170_));
  NOR2_X1    g15216(.A1(new_n13395_), .A2(new_n7345_), .ZN(new_n18171_));
  NOR2_X1    g15217(.A1(new_n18171_), .A2(pi0038), .ZN(new_n18172_));
  OAI22_X1   g15218(.A1(new_n18172_), .A2(new_n3232_), .B1(pi0178), .B2(new_n13399_), .ZN(new_n18173_));
  NOR2_X1    g15219(.A1(new_n3232_), .A2(pi0688), .ZN(new_n18174_));
  AOI22_X1   g15220(.A1(new_n18125_), .A2(new_n18174_), .B1(new_n18170_), .B2(new_n18173_), .ZN(new_n18175_));
  NOR3_X1    g15221(.A1(new_n18125_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n18176_));
  NOR4_X1    g15222(.A1(new_n18175_), .A2(new_n12970_), .A3(pi1153), .A4(new_n18124_), .ZN(new_n18177_));
  NOR2_X1    g15223(.A1(new_n18177_), .A2(new_n18176_), .ZN(new_n18178_));
  MUX2_X1    g15224(.I0(new_n18178_), .I1(new_n18175_), .S(new_n11891_), .Z(new_n18179_));
  NOR2_X1    g15225(.A1(new_n18179_), .A2(new_n13024_), .ZN(new_n18180_));
  AOI21_X1   g15226(.A1(new_n13024_), .A2(new_n18124_), .B(new_n18180_), .ZN(new_n18181_));
  AOI21_X1   g15227(.A1(new_n18181_), .A2(new_n11961_), .B(new_n18169_), .ZN(new_n18182_));
  AOI21_X1   g15228(.A1(new_n18182_), .A2(new_n12014_), .B(new_n18168_), .ZN(new_n18183_));
  AOI21_X1   g15229(.A1(new_n18183_), .A2(new_n13114_), .B(new_n18167_), .ZN(new_n18184_));
  INV_X1     g15230(.I(new_n18184_), .ZN(new_n18185_));
  NAND3_X1   g15231(.A1(new_n18124_), .A2(pi0628), .A3(pi1156), .ZN(new_n18186_));
  NOR4_X1    g15232(.A1(new_n18184_), .A2(new_n12031_), .A3(pi1156), .A4(new_n18124_), .ZN(new_n18187_));
  INV_X1     g15233(.I(new_n18187_), .ZN(new_n18188_));
  NAND2_X1   g15234(.A1(new_n18188_), .A2(new_n18186_), .ZN(new_n18189_));
  MUX2_X1    g15235(.I0(new_n18189_), .I1(new_n18185_), .S(new_n11868_), .Z(new_n18190_));
  AOI21_X1   g15236(.A1(new_n18190_), .A2(pi0647), .B(new_n18166_), .ZN(new_n18191_));
  NAND2_X1   g15237(.A1(new_n18191_), .A2(pi1157), .ZN(new_n18192_));
  NOR2_X1    g15238(.A1(new_n18125_), .A2(new_n12061_), .ZN(new_n18193_));
  AOI21_X1   g15239(.A1(new_n18190_), .A2(new_n12061_), .B(new_n18193_), .ZN(new_n18194_));
  NAND2_X1   g15240(.A1(new_n18194_), .A2(new_n12049_), .ZN(new_n18195_));
  NAND2_X1   g15241(.A1(new_n18192_), .A2(new_n18195_), .ZN(new_n18196_));
  NOR2_X1    g15242(.A1(new_n18190_), .A2(pi0787), .ZN(new_n18197_));
  AOI21_X1   g15243(.A1(new_n18196_), .A2(pi0787), .B(new_n18197_), .ZN(new_n18198_));
  AOI21_X1   g15244(.A1(new_n18198_), .A2(pi0644), .B(pi0715), .ZN(new_n18199_));
  NOR2_X1    g15245(.A1(new_n18165_), .A2(new_n18199_), .ZN(new_n18200_));
  NAND3_X1   g15246(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n18201_));
  OR2_X2     g15247(.A1(new_n18162_), .A2(new_n18201_), .Z(new_n18202_));
  NAND2_X1   g15248(.A1(new_n18202_), .A2(pi0715), .ZN(new_n18203_));
  AOI21_X1   g15249(.A1(new_n12082_), .A2(new_n18198_), .B(new_n18203_), .ZN(new_n18204_));
  OAI21_X1   g15250(.A1(new_n18204_), .A2(new_n18200_), .B(pi0790), .ZN(new_n18205_));
  NAND2_X1   g15251(.A1(new_n18153_), .A2(pi0619), .ZN(new_n18206_));
  NAND2_X1   g15252(.A1(new_n18124_), .A2(pi0619), .ZN(new_n18207_));
  NOR3_X1    g15253(.A1(new_n18134_), .A2(new_n15830_), .A3(new_n3231_), .ZN(new_n18217_));
  AOI21_X1   g15254(.A1(pi0178), .A2(new_n3232_), .B(new_n18217_), .ZN(new_n18218_));
  INV_X1     g15255(.I(new_n18177_), .ZN(new_n18219_));
  NAND2_X1   g15256(.A1(new_n18218_), .A2(pi0625), .ZN(new_n18220_));
  NAND2_X1   g15257(.A1(new_n18137_), .A2(pi0625), .ZN(new_n18221_));
  NAND4_X1   g15258(.A1(new_n18221_), .A2(new_n12977_), .A3(new_n18219_), .A4(new_n18220_), .ZN(new_n18222_));
  NAND2_X1   g15259(.A1(new_n18136_), .A2(new_n12970_), .ZN(new_n18223_));
  AND3_X2    g15260(.A1(new_n18220_), .A2(new_n11893_), .A3(new_n18223_), .Z(new_n18224_));
  OAI21_X1   g15261(.A1(new_n18224_), .A2(new_n18176_), .B(new_n13657_), .ZN(new_n18225_));
  AOI21_X1   g15262(.A1(new_n18225_), .A2(new_n18222_), .B(new_n11891_), .ZN(new_n18226_));
  AOI21_X1   g15263(.A1(new_n11891_), .A2(new_n18218_), .B(new_n18226_), .ZN(new_n18227_));
  NOR2_X1    g15264(.A1(new_n18227_), .A2(pi0785), .ZN(new_n18228_));
  INV_X1     g15265(.I(new_n18179_), .ZN(new_n18229_));
  NAND3_X1   g15266(.A1(new_n18229_), .A2(pi0609), .A3(pi1155), .ZN(new_n18230_));
  NAND3_X1   g15267(.A1(new_n18230_), .A2(new_n11923_), .A3(new_n18144_), .ZN(new_n18231_));
  NOR4_X1    g15268(.A1(new_n18227_), .A2(new_n11903_), .A3(pi1155), .A4(new_n18229_), .ZN(new_n18232_));
  NAND2_X1   g15269(.A1(new_n18142_), .A2(pi0660), .ZN(new_n18233_));
  NOR2_X1    g15270(.A1(new_n18232_), .A2(new_n18233_), .ZN(new_n18234_));
  NOR2_X1    g15271(.A1(new_n18234_), .A2(new_n11870_), .ZN(new_n18235_));
  AOI21_X1   g15272(.A1(new_n18235_), .A2(new_n18231_), .B(new_n18228_), .ZN(new_n18236_));
  INV_X1     g15273(.I(new_n18181_), .ZN(new_n18237_));
  NOR4_X1    g15274(.A1(new_n18236_), .A2(new_n11934_), .A3(pi1154), .A4(new_n18237_), .ZN(new_n18238_));
  NAND2_X1   g15275(.A1(new_n18148_), .A2(pi0627), .ZN(new_n18239_));
  NOR3_X1    g15276(.A1(new_n18181_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n18240_));
  NAND2_X1   g15277(.A1(new_n18151_), .A2(new_n11949_), .ZN(new_n18241_));
  OAI22_X1   g15278(.A1(new_n18238_), .A2(new_n18239_), .B1(new_n18240_), .B2(new_n18241_), .ZN(new_n18242_));
  MUX2_X1    g15279(.I0(new_n18242_), .I1(new_n18236_), .S(new_n11969_), .Z(new_n18243_));
  XNOR2_X1   g15280(.A1(new_n18243_), .A2(new_n18182_), .ZN(new_n18244_));
  NOR2_X1    g15281(.A1(new_n18244_), .A2(new_n11967_), .ZN(new_n18245_));
  NAND3_X1   g15282(.A1(new_n18206_), .A2(new_n11869_), .A3(new_n18207_), .ZN(new_n18246_));
  XNOR2_X1   g15283(.A1(new_n18245_), .A2(new_n18243_), .ZN(new_n18247_));
  NAND2_X1   g15284(.A1(new_n18247_), .A2(new_n11869_), .ZN(new_n18248_));
  AOI21_X1   g15285(.A1(new_n18125_), .A2(new_n11967_), .B(pi1159), .ZN(new_n18249_));
  AOI21_X1   g15286(.A1(new_n18206_), .A2(new_n18249_), .B(pi0648), .ZN(new_n18250_));
  INV_X1     g15287(.I(new_n18157_), .ZN(new_n18251_));
  MUX2_X1    g15288(.I0(new_n18251_), .I1(new_n18125_), .S(new_n11994_), .Z(new_n18252_));
  AOI21_X1   g15289(.A1(new_n18157_), .A2(new_n18125_), .B(new_n11994_), .ZN(new_n18253_));
  OAI21_X1   g15290(.A1(new_n18183_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n18254_));
  AOI21_X1   g15291(.A1(new_n18253_), .A2(new_n11990_), .B(new_n18254_), .ZN(new_n18255_));
  OAI21_X1   g15292(.A1(new_n18252_), .A2(new_n17167_), .B(new_n18255_), .ZN(new_n18256_));
  OAI21_X1   g15293(.A1(new_n18243_), .A2(pi0789), .B(new_n11998_), .ZN(new_n18257_));
  NAND3_X1   g15294(.A1(new_n18256_), .A2(new_n17372_), .A3(new_n18257_), .ZN(new_n18258_));
  AOI21_X1   g15295(.A1(new_n18248_), .A2(new_n18250_), .B(new_n18258_), .ZN(new_n18259_));
  NAND2_X1   g15296(.A1(new_n18186_), .A2(pi0629), .ZN(new_n18260_));
  OAI21_X1   g15297(.A1(new_n18187_), .A2(pi0629), .B(new_n18260_), .ZN(new_n18261_));
  NAND2_X1   g15298(.A1(new_n18158_), .A2(new_n15222_), .ZN(new_n18262_));
  NAND2_X1   g15299(.A1(new_n18262_), .A2(new_n18261_), .ZN(new_n18263_));
  AOI22_X1   g15300(.A1(new_n18259_), .A2(new_n18246_), .B1(pi0792), .B2(new_n18263_), .ZN(new_n18264_));
  NAND2_X1   g15301(.A1(new_n18191_), .A2(new_n12060_), .ZN(new_n18265_));
  AOI21_X1   g15302(.A1(new_n18194_), .A2(pi0630), .B(new_n15214_), .ZN(new_n18266_));
  NAND2_X1   g15303(.A1(new_n18266_), .A2(new_n18265_), .ZN(new_n18267_));
  NOR2_X1    g15304(.A1(new_n18160_), .A2(new_n15183_), .ZN(new_n18268_));
  NAND2_X1   g15305(.A1(new_n18165_), .A2(new_n12082_), .ZN(new_n18269_));
  AOI21_X1   g15306(.A1(new_n18202_), .A2(pi0644), .B(pi0790), .ZN(new_n18270_));
  AOI22_X1   g15307(.A1(new_n18269_), .A2(new_n18270_), .B1(new_n18267_), .B2(new_n18268_), .ZN(new_n18271_));
  OAI21_X1   g15308(.A1(new_n18264_), .A2(new_n14725_), .B(new_n18271_), .ZN(new_n18272_));
  AOI21_X1   g15309(.A1(new_n18272_), .A2(new_n18205_), .B(po1038), .ZN(new_n18273_));
  OAI21_X1   g15310(.A1(new_n6845_), .A2(pi0178), .B(new_n13184_), .ZN(new_n18274_));
  OAI21_X1   g15311(.A1(new_n18273_), .A2(new_n18274_), .B(new_n18123_), .ZN(po0335));
  NOR2_X1    g15312(.A1(new_n2925_), .A2(pi0179), .ZN(new_n18276_));
  NOR2_X1    g15313(.A1(new_n11877_), .A2(pi0741), .ZN(new_n18277_));
  NOR2_X1    g15314(.A1(new_n18277_), .A2(new_n18276_), .ZN(new_n18278_));
  INV_X1     g15315(.I(new_n18278_), .ZN(new_n18279_));
  AOI21_X1   g15316(.A1(new_n11886_), .A2(new_n15811_), .B(new_n18276_), .ZN(new_n18280_));
  NOR2_X1    g15317(.A1(new_n18280_), .A2(new_n11874_), .ZN(new_n18281_));
  NOR2_X1    g15318(.A1(new_n18279_), .A2(new_n18281_), .ZN(new_n18282_));
  NOR2_X1    g15319(.A1(new_n18282_), .A2(pi0778), .ZN(new_n18283_));
  NAND2_X1   g15320(.A1(new_n18281_), .A2(pi0625), .ZN(new_n18284_));
  NOR3_X1    g15321(.A1(new_n11894_), .A2(pi0625), .A3(pi0724), .ZN(new_n18285_));
  NOR4_X1    g15322(.A1(new_n18277_), .A2(pi0608), .A3(new_n11893_), .A4(new_n18276_), .ZN(new_n18286_));
  OAI21_X1   g15323(.A1(new_n18279_), .A2(new_n18281_), .B(new_n18284_), .ZN(new_n18287_));
  NOR3_X1    g15324(.A1(new_n18276_), .A2(pi0608), .A3(pi1153), .ZN(new_n18288_));
  AOI22_X1   g15325(.A1(new_n18287_), .A2(new_n18288_), .B1(new_n18284_), .B2(new_n18286_), .ZN(new_n18289_));
  NOR2_X1    g15326(.A1(new_n18289_), .A2(new_n11891_), .ZN(new_n18290_));
  XOR2_X1    g15327(.A1(new_n18290_), .A2(new_n18283_), .Z(new_n18291_));
  INV_X1     g15328(.I(new_n18291_), .ZN(new_n18292_));
  NAND2_X1   g15329(.A1(new_n18292_), .A2(new_n11870_), .ZN(new_n18293_));
  AOI21_X1   g15330(.A1(new_n18291_), .A2(new_n11903_), .B(pi1155), .ZN(new_n18294_));
  INV_X1     g15331(.I(new_n18280_), .ZN(new_n18295_));
  XOR2_X1    g15332(.A1(new_n18285_), .A2(pi1153), .Z(new_n18296_));
  NAND2_X1   g15333(.A1(new_n18296_), .A2(new_n18295_), .ZN(new_n18297_));
  OAI21_X1   g15334(.A1(new_n18285_), .A2(new_n18276_), .B(new_n11893_), .ZN(new_n18298_));
  AOI21_X1   g15335(.A1(new_n18297_), .A2(new_n18298_), .B(new_n11891_), .ZN(new_n18299_));
  NOR2_X1    g15336(.A1(new_n18280_), .A2(pi0778), .ZN(new_n18300_));
  OAI21_X1   g15337(.A1(new_n18299_), .A2(new_n18300_), .B(pi0609), .ZN(new_n18301_));
  AOI21_X1   g15338(.A1(new_n18279_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n18302_));
  NOR2_X1    g15339(.A1(new_n18302_), .A2(pi0660), .ZN(new_n18303_));
  OAI21_X1   g15340(.A1(new_n18294_), .A2(new_n18301_), .B(new_n18303_), .ZN(new_n18304_));
  NOR2_X1    g15341(.A1(new_n18299_), .A2(new_n18300_), .ZN(new_n18305_));
  NAND4_X1   g15342(.A1(new_n18292_), .A2(pi0609), .A3(new_n11912_), .A4(new_n18305_), .ZN(new_n18306_));
  NOR2_X1    g15343(.A1(new_n18278_), .A2(new_n11925_), .ZN(new_n18307_));
  AOI21_X1   g15344(.A1(new_n18307_), .A2(new_n11928_), .B(pi1155), .ZN(new_n18308_));
  NOR2_X1    g15345(.A1(new_n18308_), .A2(new_n11923_), .ZN(new_n18309_));
  NAND2_X1   g15346(.A1(new_n18306_), .A2(new_n18309_), .ZN(new_n18310_));
  NAND3_X1   g15347(.A1(new_n18310_), .A2(pi0785), .A3(new_n18304_), .ZN(new_n18311_));
  NAND2_X1   g15348(.A1(new_n18311_), .A2(new_n18293_), .ZN(new_n18312_));
  NOR4_X1    g15349(.A1(new_n18305_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n18314_));
  NOR2_X1    g15350(.A1(new_n18307_), .A2(pi0785), .ZN(new_n18315_));
  OAI21_X1   g15351(.A1(new_n18308_), .A2(new_n18302_), .B(pi0785), .ZN(new_n18316_));
  XNOR2_X1   g15352(.A1(new_n18316_), .A2(new_n18315_), .ZN(new_n18317_));
  INV_X1     g15353(.I(new_n18317_), .ZN(new_n18318_));
  NOR2_X1    g15354(.A1(new_n18318_), .A2(new_n11945_), .ZN(new_n18319_));
  NOR3_X1    g15355(.A1(new_n18319_), .A2(pi0627), .A3(new_n18314_), .ZN(new_n18320_));
  AOI21_X1   g15356(.A1(new_n18317_), .A2(new_n11951_), .B(pi1154), .ZN(new_n18321_));
  NOR2_X1    g15357(.A1(new_n18305_), .A2(new_n11939_), .ZN(new_n18322_));
  INV_X1     g15358(.I(new_n18322_), .ZN(new_n18323_));
  NAND4_X1   g15359(.A1(new_n18312_), .A2(pi0618), .A3(new_n11950_), .A4(new_n18323_), .ZN(new_n18324_));
  NAND2_X1   g15360(.A1(new_n18324_), .A2(new_n18321_), .ZN(new_n18325_));
  AOI21_X1   g15361(.A1(new_n18325_), .A2(new_n11949_), .B(new_n18320_), .ZN(new_n18326_));
  NOR2_X1    g15362(.A1(new_n18326_), .A2(new_n11969_), .ZN(new_n18327_));
  AOI21_X1   g15363(.A1(new_n11969_), .A2(new_n18312_), .B(new_n18327_), .ZN(new_n18328_));
  NOR2_X1    g15364(.A1(new_n18323_), .A2(new_n11962_), .ZN(new_n18329_));
  NOR4_X1    g15365(.A1(new_n18328_), .A2(new_n11967_), .A3(pi1159), .A4(new_n18329_), .ZN(new_n18330_));
  INV_X1     g15366(.I(new_n18319_), .ZN(new_n18331_));
  NAND2_X1   g15367(.A1(new_n18331_), .A2(new_n18321_), .ZN(new_n18332_));
  MUX2_X1    g15368(.I0(new_n18332_), .I1(new_n18317_), .S(new_n11969_), .Z(new_n18333_));
  NAND2_X1   g15369(.A1(new_n18333_), .A2(pi0619), .ZN(new_n18334_));
  INV_X1     g15370(.I(new_n18334_), .ZN(new_n18335_));
  INV_X1     g15371(.I(new_n18276_), .ZN(new_n18336_));
  OAI21_X1   g15372(.A1(new_n18336_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n18337_));
  NOR4_X1    g15373(.A1(new_n18330_), .A2(new_n11966_), .A3(new_n18335_), .A4(new_n18337_), .ZN(new_n18338_));
  NOR4_X1    g15374(.A1(new_n18323_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n18339_));
  OAI21_X1   g15375(.A1(new_n18276_), .A2(pi0619), .B(new_n11869_), .ZN(new_n18340_));
  OAI21_X1   g15376(.A1(new_n18335_), .A2(new_n18340_), .B(new_n11966_), .ZN(new_n18341_));
  NOR2_X1    g15377(.A1(new_n18341_), .A2(new_n18339_), .ZN(new_n18342_));
  AOI21_X1   g15378(.A1(new_n18328_), .A2(new_n11998_), .B(pi0789), .ZN(new_n18343_));
  OAI21_X1   g15379(.A1(new_n18338_), .A2(new_n18342_), .B(new_n18343_), .ZN(new_n18344_));
  NAND2_X1   g15380(.A1(new_n18329_), .A2(new_n17450_), .ZN(new_n18345_));
  NOR2_X1    g15381(.A1(new_n18345_), .A2(new_n17153_), .ZN(new_n18346_));
  INV_X1     g15382(.I(new_n18346_), .ZN(new_n18347_));
  NOR2_X1    g15383(.A1(new_n18347_), .A2(new_n17151_), .ZN(new_n18348_));
  NOR2_X1    g15384(.A1(new_n14624_), .A2(new_n18276_), .ZN(new_n18349_));
  NAND3_X1   g15385(.A1(new_n18336_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n18350_));
  MUX2_X1    g15386(.I0(new_n18350_), .I1(new_n18333_), .S(new_n11985_), .Z(new_n18351_));
  AOI21_X1   g15387(.A1(new_n18351_), .A2(new_n14624_), .B(new_n18349_), .ZN(new_n18352_));
  AND2_X2    g15388(.A1(new_n18352_), .A2(new_n12064_), .Z(new_n18353_));
  OAI21_X1   g15389(.A1(new_n18353_), .A2(new_n18348_), .B(pi0629), .ZN(new_n18354_));
  NAND2_X1   g15390(.A1(new_n18352_), .A2(new_n12063_), .ZN(new_n18355_));
  NAND2_X1   g15391(.A1(new_n18346_), .A2(new_n15084_), .ZN(new_n18356_));
  NAND4_X1   g15392(.A1(new_n18354_), .A2(new_n15085_), .A3(new_n18355_), .A4(new_n18356_), .ZN(new_n18357_));
  MUX2_X1    g15393(.I0(new_n18351_), .I1(new_n18336_), .S(new_n11994_), .Z(new_n18358_));
  NOR2_X1    g15394(.A1(new_n18358_), .A2(new_n17167_), .ZN(new_n18359_));
  OAI21_X1   g15395(.A1(new_n18351_), .A2(new_n18276_), .B(pi0626), .ZN(new_n18360_));
  NOR2_X1    g15396(.A1(new_n18345_), .A2(new_n12020_), .ZN(new_n18361_));
  NOR2_X1    g15397(.A1(new_n18361_), .A2(pi0788), .ZN(new_n18362_));
  OAI21_X1   g15398(.A1(new_n18360_), .A2(new_n17171_), .B(new_n18362_), .ZN(new_n18363_));
  OAI21_X1   g15399(.A1(new_n18359_), .A2(new_n18363_), .B(new_n14732_), .ZN(new_n18364_));
  AOI21_X1   g15400(.A1(new_n18357_), .A2(new_n14726_), .B(new_n18364_), .ZN(new_n18365_));
  NAND3_X1   g15401(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n18276_), .ZN(new_n18366_));
  NOR2_X1    g15402(.A1(new_n18347_), .A2(new_n12068_), .ZN(new_n18367_));
  INV_X1     g15403(.I(new_n18367_), .ZN(new_n18368_));
  NAND2_X1   g15404(.A1(new_n18368_), .A2(pi0647), .ZN(new_n18369_));
  NAND2_X1   g15405(.A1(new_n18276_), .A2(pi0647), .ZN(new_n18370_));
  NAND3_X1   g15406(.A1(new_n18369_), .A2(new_n12049_), .A3(new_n18370_), .ZN(new_n18371_));
  NOR2_X1    g15407(.A1(new_n18336_), .A2(pi0647), .ZN(new_n18372_));
  AOI21_X1   g15408(.A1(new_n18367_), .A2(pi0647), .B(new_n18372_), .ZN(new_n18373_));
  NAND2_X1   g15409(.A1(new_n18373_), .A2(new_n12088_), .ZN(new_n18374_));
  NAND2_X1   g15410(.A1(new_n18374_), .A2(pi0787), .ZN(new_n18375_));
  AOI21_X1   g15411(.A1(pi0630), .A2(new_n18371_), .B(new_n18375_), .ZN(new_n18376_));
  AOI22_X1   g15412(.A1(new_n18344_), .A2(new_n18365_), .B1(new_n18366_), .B2(new_n18376_), .ZN(new_n18377_));
  NOR2_X1    g15413(.A1(new_n18377_), .A2(new_n12082_), .ZN(new_n18378_));
  NAND4_X1   g15414(.A1(new_n18369_), .A2(pi0787), .A3(new_n12049_), .A4(new_n18370_), .ZN(new_n18379_));
  OAI21_X1   g15415(.A1(pi0787), .A2(new_n18368_), .B(new_n18379_), .ZN(new_n18380_));
  NOR2_X1    g15416(.A1(new_n18380_), .A2(pi0644), .ZN(new_n18381_));
  OR3_X2     g15417(.A1(new_n18378_), .A2(pi0715), .A3(new_n18381_), .Z(new_n18382_));
  MUX2_X1    g15418(.I0(new_n18352_), .I1(new_n18276_), .S(new_n16841_), .Z(new_n18383_));
  INV_X1     g15419(.I(new_n18383_), .ZN(new_n18384_));
  OAI21_X1   g15420(.A1(new_n18383_), .A2(new_n18276_), .B(new_n12082_), .ZN(new_n18385_));
  AOI21_X1   g15421(.A1(new_n18276_), .A2(new_n18383_), .B(new_n18385_), .ZN(new_n18386_));
  OAI21_X1   g15422(.A1(new_n18386_), .A2(new_n18384_), .B(new_n12099_), .ZN(new_n18387_));
  AOI21_X1   g15423(.A1(new_n18384_), .A2(new_n18386_), .B(new_n18387_), .ZN(new_n18388_));
  AOI21_X1   g15424(.A1(new_n18382_), .A2(new_n18388_), .B(pi1160), .ZN(new_n18389_));
  XOR2_X1    g15425(.A1(new_n18386_), .A2(new_n18276_), .Z(new_n18390_));
  AOI21_X1   g15426(.A1(new_n18380_), .A2(pi0644), .B(new_n13169_), .ZN(new_n18391_));
  OAI21_X1   g15427(.A1(new_n18390_), .A2(new_n12099_), .B(new_n18391_), .ZN(new_n18392_));
  OAI21_X1   g15428(.A1(new_n18378_), .A2(new_n18392_), .B(pi0790), .ZN(new_n18393_));
  NOR2_X1    g15429(.A1(new_n18377_), .A2(new_n14748_), .ZN(new_n18394_));
  OAI21_X1   g15430(.A1(new_n18389_), .A2(new_n18393_), .B(new_n18394_), .ZN(new_n18395_));
  NOR3_X1    g15431(.A1(new_n13337_), .A2(pi0039), .A3(new_n8983_), .ZN(new_n18396_));
  NAND2_X1   g15432(.A1(new_n13332_), .A2(new_n18396_), .ZN(new_n18397_));
  OAI21_X1   g15433(.A1(new_n12616_), .A2(new_n8983_), .B(new_n3154_), .ZN(new_n18398_));
  AOI21_X1   g15434(.A1(pi0179), .A2(new_n13360_), .B(new_n18398_), .ZN(new_n18399_));
  NAND2_X1   g15435(.A1(new_n18397_), .A2(new_n18399_), .ZN(new_n18400_));
  NAND2_X1   g15436(.A1(new_n18400_), .A2(new_n3172_), .ZN(new_n18401_));
  NOR2_X1    g15437(.A1(new_n12828_), .A2(pi0179), .ZN(new_n18402_));
  INV_X1     g15438(.I(new_n18402_), .ZN(new_n18403_));
  AOI21_X1   g15439(.A1(new_n18403_), .A2(new_n13374_), .B(new_n15815_), .ZN(new_n18404_));
  NAND2_X1   g15440(.A1(new_n18401_), .A2(new_n18404_), .ZN(new_n18405_));
  AOI22_X1   g15441(.A1(new_n18405_), .A2(new_n15811_), .B1(pi0179), .B2(new_n3232_), .ZN(new_n18410_));
  INV_X1     g15442(.I(new_n18410_), .ZN(new_n18411_));
  AOI21_X1   g15443(.A1(new_n18403_), .A2(new_n13403_), .B(pi0724), .ZN(new_n18412_));
  INV_X1     g15444(.I(new_n18412_), .ZN(new_n18413_));
  OAI21_X1   g15445(.A1(new_n13395_), .A2(new_n8983_), .B(new_n3172_), .ZN(new_n18414_));
  NAND2_X1   g15446(.A1(new_n18414_), .A2(new_n3231_), .ZN(new_n18415_));
  NAND2_X1   g15447(.A1(new_n14382_), .A2(new_n8983_), .ZN(new_n18416_));
  NAND2_X1   g15448(.A1(new_n18416_), .A2(new_n18415_), .ZN(new_n18417_));
  AOI21_X1   g15449(.A1(new_n3231_), .A2(new_n15811_), .B(pi0179), .ZN(new_n18418_));
  AOI22_X1   g15450(.A1(new_n18417_), .A2(new_n18413_), .B1(new_n14396_), .B2(new_n18418_), .ZN(new_n18419_));
  NOR2_X1    g15451(.A1(new_n18419_), .A2(pi0625), .ZN(new_n18420_));
  NOR2_X1    g15452(.A1(new_n12965_), .A2(pi0179), .ZN(new_n18421_));
  INV_X1     g15453(.I(new_n18421_), .ZN(new_n18422_));
  AOI21_X1   g15454(.A1(new_n18422_), .A2(new_n12970_), .B(pi1153), .ZN(new_n18423_));
  OR3_X2     g15455(.A1(new_n18420_), .A2(pi0608), .A3(new_n18423_), .Z(new_n18424_));
  NOR2_X1    g15456(.A1(new_n18410_), .A2(new_n13659_), .ZN(new_n18425_));
  NOR3_X1    g15457(.A1(new_n11893_), .A2(pi0608), .A3(pi0625), .ZN(new_n18427_));
  AOI22_X1   g15458(.A1(new_n18424_), .A2(new_n18425_), .B1(new_n18411_), .B2(new_n18427_), .ZN(new_n18428_));
  MUX2_X1    g15459(.I0(new_n18428_), .I1(new_n18410_), .S(new_n11891_), .Z(new_n18429_));
  NAND2_X1   g15460(.A1(new_n18429_), .A2(new_n11870_), .ZN(new_n18430_));
  NOR3_X1    g15461(.A1(new_n18419_), .A2(new_n13433_), .A3(new_n13434_), .ZN(new_n18431_));
  NOR2_X1    g15462(.A1(new_n18422_), .A2(new_n13435_), .ZN(new_n18432_));
  XOR2_X1    g15463(.A1(new_n18431_), .A2(new_n18432_), .Z(new_n18433_));
  NOR2_X1    g15464(.A1(new_n18419_), .A2(pi0778), .ZN(new_n18434_));
  INV_X1     g15465(.I(new_n18434_), .ZN(new_n18435_));
  OAI21_X1   g15466(.A1(new_n18433_), .A2(new_n11891_), .B(new_n18435_), .ZN(new_n18436_));
  NAND2_X1   g15467(.A1(new_n18436_), .A2(new_n11903_), .ZN(new_n18437_));
  OAI21_X1   g15468(.A1(new_n18422_), .A2(new_n12996_), .B(new_n11912_), .ZN(new_n18438_));
  AOI21_X1   g15469(.A1(new_n18438_), .A2(pi0660), .B(new_n11903_), .ZN(new_n18439_));
  INV_X1     g15470(.I(new_n18439_), .ZN(new_n18440_));
  AOI21_X1   g15471(.A1(new_n18437_), .A2(pi1155), .B(new_n18440_), .ZN(new_n18441_));
  NAND2_X1   g15472(.A1(new_n18429_), .A2(new_n11903_), .ZN(new_n18442_));
  NOR2_X1    g15473(.A1(new_n11923_), .A2(pi1155), .ZN(new_n18443_));
  INV_X1     g15474(.I(new_n18443_), .ZN(new_n18444_));
  AOI21_X1   g15475(.A1(new_n18436_), .A2(pi0609), .B(new_n18444_), .ZN(new_n18445_));
  AOI22_X1   g15476(.A1(new_n18442_), .A2(new_n18445_), .B1(new_n18441_), .B2(new_n18429_), .ZN(new_n18446_));
  OR3_X2     g15477(.A1(new_n18446_), .A2(new_n11870_), .A3(new_n18430_), .Z(new_n18447_));
  OAI21_X1   g15478(.A1(new_n18446_), .A2(new_n11870_), .B(new_n18430_), .ZN(new_n18448_));
  NAND2_X1   g15479(.A1(new_n18447_), .A2(new_n18448_), .ZN(new_n18449_));
  NOR2_X1    g15480(.A1(new_n18449_), .A2(pi0781), .ZN(new_n18450_));
  INV_X1     g15481(.I(new_n18450_), .ZN(new_n18451_));
  INV_X1     g15482(.I(new_n18449_), .ZN(new_n18452_));
  NOR2_X1    g15483(.A1(new_n18422_), .A2(new_n11938_), .ZN(new_n18453_));
  AOI21_X1   g15484(.A1(new_n18436_), .A2(new_n11938_), .B(new_n18453_), .ZN(new_n18454_));
  INV_X1     g15485(.I(new_n18454_), .ZN(new_n18455_));
  AOI21_X1   g15486(.A1(new_n18455_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n18456_));
  OAI21_X1   g15487(.A1(new_n18422_), .A2(new_n11924_), .B(new_n11870_), .ZN(new_n18457_));
  OAI21_X1   g15488(.A1(new_n18422_), .A2(new_n11915_), .B(pi1155), .ZN(new_n18458_));
  AOI21_X1   g15489(.A1(new_n18438_), .A2(new_n18458_), .B(new_n11870_), .ZN(new_n18459_));
  XOR2_X1    g15490(.A1(new_n18459_), .A2(new_n18457_), .Z(new_n18460_));
  NOR2_X1    g15491(.A1(new_n18460_), .A2(new_n11934_), .ZN(new_n18461_));
  NOR2_X1    g15492(.A1(new_n18422_), .A2(new_n11934_), .ZN(new_n18462_));
  NOR4_X1    g15493(.A1(new_n18461_), .A2(new_n11949_), .A3(pi1154), .A4(new_n18462_), .ZN(new_n18463_));
  NOR3_X1    g15494(.A1(new_n18456_), .A2(new_n11934_), .A3(new_n18463_), .ZN(new_n18464_));
  NAND3_X1   g15495(.A1(new_n18447_), .A2(new_n18448_), .A3(new_n11934_), .ZN(new_n18465_));
  OAI21_X1   g15496(.A1(new_n18421_), .A2(pi0618), .B(new_n11950_), .ZN(new_n18466_));
  OAI21_X1   g15497(.A1(new_n18461_), .A2(new_n18466_), .B(new_n11949_), .ZN(new_n18467_));
  NAND2_X1   g15498(.A1(new_n18455_), .A2(pi0618), .ZN(new_n18468_));
  AND3_X2    g15499(.A1(new_n18468_), .A2(new_n11950_), .A3(new_n18467_), .Z(new_n18469_));
  AOI22_X1   g15500(.A1(new_n18452_), .A2(new_n18464_), .B1(new_n18465_), .B2(new_n18469_), .ZN(new_n18470_));
  NOR3_X1    g15501(.A1(new_n18470_), .A2(new_n11969_), .A3(new_n18451_), .ZN(new_n18471_));
  OAI21_X1   g15502(.A1(new_n18470_), .A2(new_n11969_), .B(new_n18451_), .ZN(new_n18472_));
  INV_X1     g15503(.I(new_n18472_), .ZN(new_n18473_));
  NOR2_X1    g15504(.A1(new_n18473_), .A2(new_n18471_), .ZN(new_n18474_));
  NAND2_X1   g15505(.A1(new_n18474_), .A2(new_n11985_), .ZN(new_n18475_));
  INV_X1     g15506(.I(new_n18475_), .ZN(new_n18476_));
  NOR2_X1    g15507(.A1(new_n18460_), .A2(pi0781), .ZN(new_n18477_));
  NOR4_X1    g15508(.A1(new_n18461_), .A2(pi0618), .A3(pi1154), .A4(new_n18421_), .ZN(new_n18478_));
  NOR2_X1    g15509(.A1(new_n18478_), .A2(new_n11969_), .ZN(new_n18479_));
  XNOR2_X1   g15510(.A1(new_n18479_), .A2(new_n18477_), .ZN(new_n18480_));
  NOR2_X1    g15511(.A1(new_n18480_), .A2(new_n11967_), .ZN(new_n18481_));
  NOR2_X1    g15512(.A1(new_n18422_), .A2(new_n11967_), .ZN(new_n18482_));
  NOR4_X1    g15513(.A1(new_n18481_), .A2(new_n11966_), .A3(pi1159), .A4(new_n18482_), .ZN(new_n18483_));
  NOR2_X1    g15514(.A1(new_n18421_), .A2(new_n11961_), .ZN(new_n18484_));
  AOI21_X1   g15515(.A1(new_n18454_), .A2(new_n11961_), .B(new_n18484_), .ZN(new_n18485_));
  NOR3_X1    g15516(.A1(new_n18483_), .A2(new_n11967_), .A3(pi1159), .ZN(new_n18486_));
  INV_X1     g15517(.I(new_n18471_), .ZN(new_n18487_));
  NAND3_X1   g15518(.A1(new_n18487_), .A2(new_n11967_), .A3(new_n18472_), .ZN(new_n18488_));
  AOI21_X1   g15519(.A1(new_n18422_), .A2(new_n11967_), .B(pi1159), .ZN(new_n18489_));
  OAI21_X1   g15520(.A1(new_n18480_), .A2(new_n11967_), .B(new_n18489_), .ZN(new_n18490_));
  AOI21_X1   g15521(.A1(new_n18485_), .A2(pi0619), .B(pi1159), .ZN(new_n18491_));
  INV_X1     g15522(.I(new_n18491_), .ZN(new_n18492_));
  AOI21_X1   g15523(.A1(new_n18490_), .A2(new_n11966_), .B(new_n18492_), .ZN(new_n18493_));
  AOI22_X1   g15524(.A1(new_n18488_), .A2(new_n18493_), .B1(new_n18474_), .B2(new_n18486_), .ZN(new_n18494_));
  INV_X1     g15525(.I(new_n18494_), .ZN(new_n18495_));
  NAND3_X1   g15526(.A1(new_n18495_), .A2(pi0789), .A3(new_n18476_), .ZN(new_n18496_));
  OAI21_X1   g15527(.A1(new_n18494_), .A2(new_n11985_), .B(new_n18475_), .ZN(new_n18497_));
  NAND2_X1   g15528(.A1(new_n18496_), .A2(new_n18497_), .ZN(new_n18498_));
  NOR3_X1    g15529(.A1(new_n18494_), .A2(new_n11985_), .A3(new_n18475_), .ZN(new_n18499_));
  INV_X1     g15530(.I(new_n18497_), .ZN(new_n18500_));
  INV_X1     g15531(.I(new_n18480_), .ZN(new_n18501_));
  NAND2_X1   g15532(.A1(new_n18501_), .A2(new_n11985_), .ZN(new_n18502_));
  NOR3_X1    g15533(.A1(new_n18421_), .A2(pi0619), .A3(pi1159), .ZN(new_n18503_));
  NOR2_X1    g15534(.A1(new_n18503_), .A2(new_n11985_), .ZN(new_n18504_));
  XOR2_X1    g15535(.A1(new_n18502_), .A2(new_n18504_), .Z(new_n18505_));
  INV_X1     g15536(.I(new_n18505_), .ZN(new_n18506_));
  NOR3_X1    g15537(.A1(new_n11994_), .A2(new_n11989_), .A3(pi1158), .ZN(new_n18507_));
  NAND2_X1   g15538(.A1(new_n18506_), .A2(new_n18507_), .ZN(new_n18508_));
  NOR2_X1    g15539(.A1(new_n18422_), .A2(new_n12014_), .ZN(new_n18509_));
  AOI21_X1   g15540(.A1(new_n18485_), .A2(new_n12014_), .B(new_n18509_), .ZN(new_n18510_));
  NOR2_X1    g15541(.A1(new_n11994_), .A2(pi0641), .ZN(new_n18511_));
  NAND2_X1   g15542(.A1(new_n18508_), .A2(new_n18511_), .ZN(new_n18512_));
  INV_X1     g15543(.I(new_n18512_), .ZN(new_n18513_));
  NOR2_X1    g15544(.A1(new_n18505_), .A2(pi0626), .ZN(new_n18514_));
  OAI21_X1   g15545(.A1(new_n18421_), .A2(new_n11994_), .B(pi0641), .ZN(new_n18515_));
  NOR3_X1    g15546(.A1(new_n11989_), .A2(pi0626), .A3(pi1158), .ZN(new_n18516_));
  OAI21_X1   g15547(.A1(new_n18514_), .A2(new_n18515_), .B(new_n18516_), .ZN(new_n18517_));
  INV_X1     g15548(.I(new_n18517_), .ZN(new_n18518_));
  OAI22_X1   g15549(.A1(new_n18500_), .A2(new_n18499_), .B1(new_n18513_), .B2(new_n18518_), .ZN(new_n18519_));
  NOR3_X1    g15550(.A1(new_n18519_), .A2(new_n11986_), .A3(new_n18498_), .ZN(new_n18520_));
  NOR2_X1    g15551(.A1(new_n18500_), .A2(new_n18499_), .ZN(new_n18521_));
  AOI21_X1   g15552(.A1(new_n18519_), .A2(pi0788), .B(new_n18521_), .ZN(new_n18522_));
  NOR2_X1    g15553(.A1(new_n18520_), .A2(new_n18522_), .ZN(new_n18523_));
  NOR2_X1    g15554(.A1(new_n18505_), .A2(new_n11997_), .ZN(new_n18524_));
  AOI21_X1   g15555(.A1(new_n11997_), .A2(new_n18422_), .B(new_n18524_), .ZN(new_n18525_));
  NAND2_X1   g15556(.A1(new_n18525_), .A2(new_n12031_), .ZN(new_n18526_));
  NOR2_X1    g15557(.A1(new_n18421_), .A2(new_n13114_), .ZN(new_n18527_));
  AOI21_X1   g15558(.A1(new_n18510_), .A2(new_n13114_), .B(new_n18527_), .ZN(new_n18528_));
  NOR3_X1    g15559(.A1(new_n18422_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n18529_));
  OAI21_X1   g15560(.A1(new_n18529_), .A2(new_n12030_), .B(pi0628), .ZN(new_n18530_));
  AOI21_X1   g15561(.A1(new_n18526_), .A2(pi1156), .B(new_n18530_), .ZN(new_n18531_));
  INV_X1     g15562(.I(new_n18525_), .ZN(new_n18532_));
  NOR2_X1    g15563(.A1(new_n18532_), .A2(new_n12031_), .ZN(new_n18533_));
  NOR2_X1    g15564(.A1(new_n12030_), .A2(pi0628), .ZN(new_n18534_));
  OAI21_X1   g15565(.A1(new_n18533_), .A2(pi1156), .B(new_n18534_), .ZN(new_n18535_));
  INV_X1     g15566(.I(new_n18535_), .ZN(new_n18536_));
  OAI22_X1   g15567(.A1(new_n18520_), .A2(new_n18522_), .B1(new_n18531_), .B2(new_n18536_), .ZN(new_n18537_));
  MUX2_X1    g15568(.I0(new_n18537_), .I1(new_n18523_), .S(new_n11868_), .Z(new_n18538_));
  AOI22_X1   g15569(.A1(new_n18496_), .A2(new_n18497_), .B1(new_n18512_), .B2(new_n18517_), .ZN(new_n18539_));
  NAND3_X1   g15570(.A1(new_n18539_), .A2(pi0788), .A3(new_n18521_), .ZN(new_n18540_));
  OAI21_X1   g15571(.A1(new_n18539_), .A2(new_n11986_), .B(new_n18498_), .ZN(new_n18541_));
  INV_X1     g15572(.I(new_n18531_), .ZN(new_n18542_));
  AOI22_X1   g15573(.A1(new_n18541_), .A2(new_n18540_), .B1(new_n18542_), .B2(new_n18535_), .ZN(new_n18543_));
  NAND3_X1   g15574(.A1(new_n18543_), .A2(pi0792), .A3(new_n18523_), .ZN(new_n18544_));
  NAND2_X1   g15575(.A1(new_n18541_), .A2(new_n18540_), .ZN(new_n18545_));
  OAI21_X1   g15576(.A1(new_n18543_), .A2(new_n11868_), .B(new_n18545_), .ZN(new_n18546_));
  NAND2_X1   g15577(.A1(new_n18546_), .A2(new_n18544_), .ZN(new_n18547_));
  NOR4_X1    g15578(.A1(new_n18528_), .A2(new_n12031_), .A3(pi1156), .A4(new_n18421_), .ZN(new_n18548_));
  NOR2_X1    g15579(.A1(new_n18548_), .A2(new_n18529_), .ZN(new_n18549_));
  MUX2_X1    g15580(.I0(new_n18549_), .I1(new_n18528_), .S(new_n11868_), .Z(new_n18550_));
  NAND2_X1   g15581(.A1(new_n18550_), .A2(pi0647), .ZN(new_n18551_));
  AOI21_X1   g15582(.A1(new_n18421_), .A2(pi0647), .B(pi1157), .ZN(new_n18552_));
  NAND2_X1   g15583(.A1(new_n18551_), .A2(new_n18552_), .ZN(new_n18553_));
  NOR2_X1    g15584(.A1(new_n18421_), .A2(new_n12054_), .ZN(new_n18554_));
  AOI21_X1   g15585(.A1(new_n18532_), .A2(new_n12054_), .B(new_n18554_), .ZN(new_n18555_));
  NOR2_X1    g15586(.A1(new_n12061_), .A2(pi1157), .ZN(new_n18556_));
  OAI21_X1   g15587(.A1(new_n18553_), .A2(new_n12060_), .B(new_n18556_), .ZN(new_n18557_));
  NOR3_X1    g15588(.A1(new_n18537_), .A2(new_n11868_), .A3(new_n18545_), .ZN(new_n18558_));
  AOI21_X1   g15589(.A1(new_n18537_), .A2(pi0792), .B(new_n18523_), .ZN(new_n18559_));
  NOR3_X1    g15590(.A1(new_n18558_), .A2(new_n18559_), .A3(pi0647), .ZN(new_n18560_));
  AOI21_X1   g15591(.A1(new_n18422_), .A2(new_n12061_), .B(pi1157), .ZN(new_n18561_));
  NAND2_X1   g15592(.A1(new_n18551_), .A2(new_n18561_), .ZN(new_n18562_));
  NAND2_X1   g15593(.A1(new_n18562_), .A2(new_n12060_), .ZN(new_n18563_));
  AOI21_X1   g15594(.A1(new_n18555_), .A2(pi0647), .B(pi1157), .ZN(new_n18564_));
  AND2_X2    g15595(.A1(new_n18564_), .A2(new_n18563_), .Z(new_n18565_));
  INV_X1     g15596(.I(new_n18565_), .ZN(new_n18566_));
  OAI22_X1   g15597(.A1(new_n18560_), .A2(new_n18566_), .B1(new_n18547_), .B2(new_n18557_), .ZN(new_n18567_));
  MUX2_X1    g15598(.I0(new_n18567_), .I1(new_n18538_), .S(new_n12048_), .Z(new_n18568_));
  NAND2_X1   g15599(.A1(new_n18550_), .A2(new_n12048_), .ZN(new_n18569_));
  INV_X1     g15600(.I(new_n18562_), .ZN(new_n18570_));
  OAI21_X1   g15601(.A1(new_n18570_), .A2(new_n18553_), .B(pi0787), .ZN(new_n18571_));
  XOR2_X1    g15602(.A1(new_n18571_), .A2(new_n18569_), .Z(new_n18572_));
  NOR2_X1    g15603(.A1(new_n18422_), .A2(new_n12092_), .ZN(new_n18573_));
  AOI21_X1   g15604(.A1(new_n18555_), .A2(new_n12092_), .B(new_n18573_), .ZN(new_n18574_));
  INV_X1     g15605(.I(new_n18574_), .ZN(new_n18575_));
  NOR2_X1    g15606(.A1(pi0644), .A2(pi0715), .ZN(new_n18576_));
  AOI21_X1   g15607(.A1(new_n18575_), .A2(new_n18576_), .B(new_n13169_), .ZN(new_n18577_));
  OAI21_X1   g15608(.A1(new_n12082_), .A2(new_n18572_), .B(new_n18577_), .ZN(new_n18578_));
  AOI21_X1   g15609(.A1(new_n18568_), .A2(new_n12082_), .B(new_n18578_), .ZN(new_n18579_));
  INV_X1     g15610(.I(new_n18557_), .ZN(new_n18580_));
  NAND3_X1   g15611(.A1(new_n18546_), .A2(new_n18544_), .A3(new_n12061_), .ZN(new_n18581_));
  AOI22_X1   g15612(.A1(new_n18581_), .A2(new_n18565_), .B1(new_n18538_), .B2(new_n18580_), .ZN(new_n18582_));
  MUX2_X1    g15613(.I0(new_n18582_), .I1(new_n18547_), .S(new_n12048_), .Z(new_n18583_));
  INV_X1     g15614(.I(new_n18572_), .ZN(new_n18584_));
  NAND3_X1   g15615(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n18585_));
  OAI21_X1   g15616(.A1(new_n18574_), .A2(new_n18585_), .B(new_n13179_), .ZN(new_n18586_));
  NOR2_X1    g15617(.A1(new_n18586_), .A2(new_n18584_), .ZN(new_n18587_));
  OAI21_X1   g15618(.A1(new_n18583_), .A2(new_n12082_), .B(new_n18587_), .ZN(new_n18588_));
  NOR2_X1    g15619(.A1(new_n18579_), .A2(new_n18588_), .ZN(new_n18589_));
  NAND2_X1   g15620(.A1(po1038), .A2(new_n8983_), .ZN(new_n18590_));
  AOI21_X1   g15621(.A1(new_n18590_), .A2(new_n13184_), .B(po1038), .ZN(new_n18591_));
  OAI21_X1   g15622(.A1(new_n18568_), .A2(pi0790), .B(new_n18591_), .ZN(new_n18592_));
  OAI21_X1   g15623(.A1(new_n18589_), .A2(new_n18592_), .B(new_n18395_), .ZN(po0336));
  NOR2_X1    g15624(.A1(new_n2925_), .A2(pi0180), .ZN(new_n18594_));
  NOR2_X1    g15625(.A1(new_n11877_), .A2(pi0753), .ZN(new_n18595_));
  NOR2_X1    g15626(.A1(new_n18595_), .A2(new_n18594_), .ZN(new_n18596_));
  AOI21_X1   g15627(.A1(new_n11886_), .A2(new_n15884_), .B(new_n18594_), .ZN(new_n18597_));
  NOR2_X1    g15628(.A1(new_n18597_), .A2(new_n11874_), .ZN(new_n18598_));
  INV_X1     g15629(.I(new_n18598_), .ZN(new_n18599_));
  NAND2_X1   g15630(.A1(new_n18599_), .A2(new_n18596_), .ZN(new_n18600_));
  NAND2_X1   g15631(.A1(new_n18600_), .A2(new_n11891_), .ZN(new_n18601_));
  NOR2_X1    g15632(.A1(new_n18599_), .A2(new_n12970_), .ZN(new_n18602_));
  NOR4_X1    g15633(.A1(new_n18602_), .A2(new_n11893_), .A3(new_n18594_), .A4(new_n18595_), .ZN(new_n18603_));
  NOR3_X1    g15634(.A1(new_n11894_), .A2(pi0625), .A3(pi0702), .ZN(new_n18604_));
  NOR2_X1    g15635(.A1(new_n18594_), .A2(pi1153), .ZN(new_n18605_));
  INV_X1     g15636(.I(new_n18605_), .ZN(new_n18606_));
  NOR2_X1    g15637(.A1(new_n18604_), .A2(new_n18606_), .ZN(new_n18607_));
  INV_X1     g15638(.I(new_n18607_), .ZN(new_n18608_));
  NAND2_X1   g15639(.A1(new_n18608_), .A2(pi0608), .ZN(new_n18609_));
  INV_X1     g15640(.I(new_n18602_), .ZN(new_n18610_));
  AOI21_X1   g15641(.A1(new_n18610_), .A2(new_n18600_), .B(new_n18606_), .ZN(new_n18611_));
  OAI21_X1   g15642(.A1(new_n18604_), .A2(new_n18597_), .B(pi1153), .ZN(new_n18612_));
  NAND2_X1   g15643(.A1(new_n18612_), .A2(new_n13657_), .ZN(new_n18613_));
  OAI22_X1   g15644(.A1(new_n18611_), .A2(new_n18613_), .B1(new_n18603_), .B2(new_n18609_), .ZN(new_n18614_));
  NAND2_X1   g15645(.A1(new_n18614_), .A2(pi0778), .ZN(new_n18615_));
  XOR2_X1    g15646(.A1(new_n18615_), .A2(new_n18601_), .Z(new_n18616_));
  INV_X1     g15647(.I(new_n18616_), .ZN(new_n18617_));
  NAND2_X1   g15648(.A1(new_n18608_), .A2(new_n18612_), .ZN(new_n18618_));
  MUX2_X1    g15649(.I0(new_n18618_), .I1(new_n18597_), .S(new_n11891_), .Z(new_n18619_));
  XNOR2_X1   g15650(.A1(new_n18616_), .A2(new_n18619_), .ZN(new_n18620_));
  NAND2_X1   g15651(.A1(new_n18620_), .A2(pi0609), .ZN(new_n18621_));
  XOR2_X1    g15652(.A1(new_n18621_), .A2(new_n18616_), .Z(new_n18622_));
  NAND2_X1   g15653(.A1(new_n18622_), .A2(new_n11912_), .ZN(new_n18623_));
  NOR2_X1    g15654(.A1(new_n18596_), .A2(new_n11925_), .ZN(new_n18624_));
  INV_X1     g15655(.I(new_n18624_), .ZN(new_n18625_));
  NOR3_X1    g15656(.A1(new_n12997_), .A2(new_n11877_), .A3(pi0753), .ZN(new_n18626_));
  NAND3_X1   g15657(.A1(new_n18625_), .A2(new_n11912_), .A3(new_n18626_), .ZN(new_n18627_));
  NAND3_X1   g15658(.A1(new_n18623_), .A2(new_n11923_), .A3(new_n18627_), .ZN(new_n18628_));
  NOR4_X1    g15659(.A1(new_n18626_), .A2(new_n11923_), .A3(pi1155), .A4(new_n18594_), .ZN(new_n18630_));
  NOR2_X1    g15660(.A1(new_n18630_), .A2(new_n11870_), .ZN(new_n18631_));
  AOI22_X1   g15661(.A1(new_n18628_), .A2(new_n18631_), .B1(new_n11870_), .B2(new_n18617_), .ZN(new_n18632_));
  NOR2_X1    g15662(.A1(new_n18632_), .A2(pi0781), .ZN(new_n18633_));
  NOR4_X1    g15663(.A1(new_n18619_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n18634_));
  NOR3_X1    g15664(.A1(new_n18626_), .A2(pi1155), .A3(new_n18594_), .ZN(new_n18635_));
  NAND2_X1   g15665(.A1(new_n18627_), .A2(new_n18635_), .ZN(new_n18636_));
  MUX2_X1    g15666(.I0(new_n18636_), .I1(new_n18625_), .S(new_n11870_), .Z(new_n18637_));
  INV_X1     g15667(.I(new_n18637_), .ZN(new_n18638_));
  OAI21_X1   g15668(.A1(new_n18638_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n18639_));
  OAI21_X1   g15669(.A1(new_n18638_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n18640_));
  NOR2_X1    g15670(.A1(new_n18619_), .A2(new_n11939_), .ZN(new_n18641_));
  NOR4_X1    g15671(.A1(new_n18632_), .A2(new_n11934_), .A3(pi1154), .A4(new_n18641_), .ZN(new_n18642_));
  NOR2_X1    g15672(.A1(new_n18642_), .A2(new_n18640_), .ZN(new_n18643_));
  OAI22_X1   g15673(.A1(new_n18643_), .A2(pi0627), .B1(new_n18634_), .B2(new_n18639_), .ZN(new_n18644_));
  AOI21_X1   g15674(.A1(new_n18644_), .A2(pi0781), .B(new_n18633_), .ZN(new_n18645_));
  INV_X1     g15675(.I(new_n18641_), .ZN(new_n18646_));
  NOR2_X1    g15676(.A1(new_n18646_), .A2(new_n11962_), .ZN(new_n18647_));
  NOR4_X1    g15677(.A1(new_n18645_), .A2(new_n11967_), .A3(pi1159), .A4(new_n18647_), .ZN(new_n18648_));
  NOR2_X1    g15678(.A1(new_n18638_), .A2(pi0781), .ZN(new_n18649_));
  AOI21_X1   g15679(.A1(new_n11944_), .A2(new_n18637_), .B(new_n18640_), .ZN(new_n18650_));
  NOR2_X1    g15680(.A1(new_n18650_), .A2(new_n11969_), .ZN(new_n18651_));
  XOR2_X1    g15681(.A1(new_n18651_), .A2(new_n18649_), .Z(new_n18652_));
  AOI21_X1   g15682(.A1(new_n18652_), .A2(new_n16479_), .B(pi1159), .ZN(new_n18653_));
  INV_X1     g15683(.I(new_n18653_), .ZN(new_n18654_));
  NOR3_X1    g15684(.A1(new_n18648_), .A2(new_n11966_), .A3(new_n18654_), .ZN(new_n18655_));
  NOR4_X1    g15685(.A1(new_n18646_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n18656_));
  INV_X1     g15686(.I(new_n18652_), .ZN(new_n18657_));
  NOR2_X1    g15687(.A1(new_n18657_), .A2(new_n16482_), .ZN(new_n18658_));
  NOR3_X1    g15688(.A1(new_n18658_), .A2(pi0648), .A3(new_n18656_), .ZN(new_n18659_));
  AOI21_X1   g15689(.A1(new_n18645_), .A2(new_n11998_), .B(pi0789), .ZN(new_n18660_));
  OAI21_X1   g15690(.A1(new_n18655_), .A2(new_n18659_), .B(new_n18660_), .ZN(new_n18661_));
  NAND2_X1   g15691(.A1(new_n18647_), .A2(new_n17450_), .ZN(new_n18662_));
  NOR2_X1    g15692(.A1(new_n18662_), .A2(new_n17153_), .ZN(new_n18663_));
  NOR2_X1    g15693(.A1(new_n14624_), .A2(new_n18594_), .ZN(new_n18664_));
  NOR2_X1    g15694(.A1(new_n18657_), .A2(pi0789), .ZN(new_n18665_));
  NOR2_X1    g15695(.A1(new_n18654_), .A2(new_n18658_), .ZN(new_n18666_));
  NOR2_X1    g15696(.A1(new_n18666_), .A2(new_n11985_), .ZN(new_n18667_));
  XOR2_X1    g15697(.A1(new_n18667_), .A2(new_n18665_), .Z(new_n18668_));
  AOI21_X1   g15698(.A1(new_n18668_), .A2(new_n14624_), .B(new_n18664_), .ZN(new_n18669_));
  AOI22_X1   g15699(.A1(new_n18669_), .A2(new_n12064_), .B1(new_n15080_), .B2(new_n18663_), .ZN(new_n18670_));
  NOR2_X1    g15700(.A1(new_n18670_), .A2(new_n12030_), .ZN(new_n18671_));
  NAND2_X1   g15701(.A1(new_n18669_), .A2(new_n12063_), .ZN(new_n18672_));
  AOI21_X1   g15702(.A1(new_n18663_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n18673_));
  NAND2_X1   g15703(.A1(new_n18672_), .A2(new_n18673_), .ZN(new_n18674_));
  OAI21_X1   g15704(.A1(new_n18671_), .A2(new_n18674_), .B(new_n14726_), .ZN(new_n18675_));
  INV_X1     g15705(.I(new_n18594_), .ZN(new_n18676_));
  MUX2_X1    g15706(.I0(new_n18668_), .I1(new_n18676_), .S(new_n11994_), .Z(new_n18677_));
  INV_X1     g15707(.I(new_n18668_), .ZN(new_n18678_));
  AOI21_X1   g15708(.A1(new_n18678_), .A2(new_n18676_), .B(new_n11994_), .ZN(new_n18679_));
  OAI21_X1   g15709(.A1(new_n18662_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n18680_));
  AOI21_X1   g15710(.A1(new_n18679_), .A2(new_n11990_), .B(new_n18680_), .ZN(new_n18681_));
  OAI21_X1   g15711(.A1(new_n17167_), .A2(new_n18677_), .B(new_n18681_), .ZN(new_n18682_));
  NAND4_X1   g15712(.A1(new_n18661_), .A2(new_n14732_), .A3(new_n18675_), .A4(new_n18682_), .ZN(new_n18683_));
  NAND3_X1   g15713(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n18594_), .ZN(new_n18684_));
  NAND2_X1   g15714(.A1(new_n18663_), .A2(new_n15050_), .ZN(new_n18685_));
  NAND2_X1   g15715(.A1(new_n18685_), .A2(pi0647), .ZN(new_n18686_));
  NAND2_X1   g15716(.A1(new_n18594_), .A2(pi0647), .ZN(new_n18687_));
  NAND3_X1   g15717(.A1(new_n18686_), .A2(new_n12049_), .A3(new_n18687_), .ZN(new_n18688_));
  NAND2_X1   g15718(.A1(new_n18688_), .A2(pi0630), .ZN(new_n18689_));
  NOR2_X1    g15719(.A1(new_n18685_), .A2(new_n12061_), .ZN(new_n18690_));
  AOI21_X1   g15720(.A1(new_n12061_), .A2(new_n18594_), .B(new_n18690_), .ZN(new_n18691_));
  NAND2_X1   g15721(.A1(new_n18691_), .A2(new_n12088_), .ZN(new_n18692_));
  NAND4_X1   g15722(.A1(new_n18692_), .A2(new_n18689_), .A3(pi0787), .A4(new_n18684_), .ZN(new_n18693_));
  AND2_X2    g15723(.A1(new_n18683_), .A2(new_n18693_), .Z(new_n18694_));
  NOR2_X1    g15724(.A1(new_n18694_), .A2(new_n12082_), .ZN(new_n18695_));
  NAND4_X1   g15725(.A1(new_n18686_), .A2(pi0787), .A3(new_n12049_), .A4(new_n18687_), .ZN(new_n18696_));
  OAI21_X1   g15726(.A1(pi0787), .A2(new_n18685_), .B(new_n18696_), .ZN(new_n18697_));
  NOR2_X1    g15727(.A1(new_n18697_), .A2(pi0644), .ZN(new_n18698_));
  OR3_X2     g15728(.A1(new_n18695_), .A2(pi0715), .A3(new_n18698_), .Z(new_n18699_));
  MUX2_X1    g15729(.I0(new_n18669_), .I1(new_n18594_), .S(new_n16841_), .Z(new_n18700_));
  INV_X1     g15730(.I(new_n18700_), .ZN(new_n18701_));
  OAI21_X1   g15731(.A1(new_n18700_), .A2(new_n18594_), .B(new_n12082_), .ZN(new_n18702_));
  AOI21_X1   g15732(.A1(new_n18594_), .A2(new_n18700_), .B(new_n18702_), .ZN(new_n18703_));
  OAI21_X1   g15733(.A1(new_n18703_), .A2(new_n18701_), .B(new_n12099_), .ZN(new_n18704_));
  AOI21_X1   g15734(.A1(new_n18701_), .A2(new_n18703_), .B(new_n18704_), .ZN(new_n18705_));
  AOI21_X1   g15735(.A1(new_n18699_), .A2(new_n18705_), .B(pi1160), .ZN(new_n18706_));
  XOR2_X1    g15736(.A1(new_n18703_), .A2(new_n18594_), .Z(new_n18707_));
  AOI21_X1   g15737(.A1(new_n18697_), .A2(pi0644), .B(new_n13169_), .ZN(new_n18708_));
  OAI21_X1   g15738(.A1(new_n18707_), .A2(new_n12099_), .B(new_n18708_), .ZN(new_n18709_));
  OAI21_X1   g15739(.A1(new_n18695_), .A2(new_n18709_), .B(pi0790), .ZN(new_n18710_));
  NOR2_X1    g15740(.A1(new_n18694_), .A2(new_n14748_), .ZN(new_n18711_));
  OAI21_X1   g15741(.A1(new_n18706_), .A2(new_n18710_), .B(new_n18711_), .ZN(new_n18712_));
  NOR2_X1    g15742(.A1(new_n12965_), .A2(pi0180), .ZN(new_n18713_));
  INV_X1     g15743(.I(new_n18713_), .ZN(new_n18714_));
  NAND2_X1   g15744(.A1(new_n18714_), .A2(new_n11997_), .ZN(new_n18715_));
  NAND2_X1   g15745(.A1(new_n12894_), .A2(pi0753), .ZN(new_n18716_));
  NOR2_X1    g15746(.A1(new_n15866_), .A2(pi0180), .ZN(new_n18717_));
  OAI21_X1   g15747(.A1(new_n14361_), .A2(new_n5324_), .B(pi0039), .ZN(new_n18720_));
  AOI21_X1   g15748(.A1(new_n12824_), .A2(new_n18717_), .B(new_n18720_), .ZN(new_n18721_));
  NOR2_X1    g15749(.A1(new_n12828_), .A2(pi0180), .ZN(new_n18722_));
  AOI21_X1   g15750(.A1(new_n12829_), .A2(new_n15866_), .B(pi0038), .ZN(new_n18723_));
  INV_X1     g15751(.I(new_n18723_), .ZN(new_n18724_));
  AOI21_X1   g15752(.A1(new_n18721_), .A2(new_n18716_), .B(new_n18724_), .ZN(new_n18725_));
  NOR2_X1    g15753(.A1(new_n18725_), .A2(new_n3232_), .ZN(new_n18726_));
  AOI21_X1   g15754(.A1(new_n5324_), .A2(new_n3232_), .B(new_n18726_), .ZN(new_n18727_));
  OAI21_X1   g15755(.A1(new_n18727_), .A2(new_n11914_), .B(new_n11870_), .ZN(new_n18728_));
  AOI21_X1   g15756(.A1(new_n11914_), .A2(new_n18713_), .B(new_n18728_), .ZN(new_n18729_));
  NAND2_X1   g15757(.A1(new_n18727_), .A2(new_n11924_), .ZN(new_n18730_));
  OAI22_X1   g15758(.A1(new_n18730_), .A2(pi0609), .B1(new_n12996_), .B2(new_n18713_), .ZN(new_n18731_));
  NAND2_X1   g15759(.A1(new_n18731_), .A2(new_n11912_), .ZN(new_n18732_));
  OAI22_X1   g15760(.A1(new_n18730_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n18713_), .ZN(new_n18733_));
  NAND2_X1   g15761(.A1(new_n18733_), .A2(pi1155), .ZN(new_n18734_));
  AOI21_X1   g15762(.A1(new_n18732_), .A2(new_n18734_), .B(new_n11870_), .ZN(new_n18735_));
  XNOR2_X1   g15763(.A1(new_n18735_), .A2(new_n18729_), .ZN(new_n18736_));
  NOR2_X1    g15764(.A1(new_n18736_), .A2(pi0781), .ZN(new_n18737_));
  NOR3_X1    g15765(.A1(new_n18713_), .A2(pi0618), .A3(pi1154), .ZN(new_n18738_));
  NOR2_X1    g15766(.A1(new_n18738_), .A2(new_n11969_), .ZN(new_n18739_));
  XOR2_X1    g15767(.A1(new_n18737_), .A2(new_n18739_), .Z(new_n18740_));
  NAND2_X1   g15768(.A1(new_n18740_), .A2(new_n11985_), .ZN(new_n18741_));
  NAND3_X1   g15769(.A1(new_n18714_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n18742_));
  NAND2_X1   g15770(.A1(new_n18742_), .A2(pi0789), .ZN(new_n18743_));
  XNOR2_X1   g15771(.A1(new_n18741_), .A2(new_n18743_), .ZN(new_n18744_));
  OAI21_X1   g15772(.A1(new_n18744_), .A2(new_n11997_), .B(new_n18715_), .ZN(new_n18745_));
  NOR2_X1    g15773(.A1(new_n18713_), .A2(new_n12054_), .ZN(new_n18746_));
  AOI21_X1   g15774(.A1(new_n18745_), .A2(new_n12054_), .B(new_n18746_), .ZN(new_n18747_));
  NAND2_X1   g15775(.A1(new_n18714_), .A2(new_n12091_), .ZN(new_n18748_));
  OAI21_X1   g15776(.A1(new_n18747_), .A2(new_n12091_), .B(new_n18748_), .ZN(new_n18749_));
  OR2_X2     g15777(.A1(new_n18749_), .A2(pi0644), .Z(new_n18750_));
  AOI21_X1   g15778(.A1(new_n18713_), .A2(pi0644), .B(new_n12099_), .ZN(new_n18751_));
  AOI21_X1   g15779(.A1(new_n18750_), .A2(new_n18751_), .B(pi1160), .ZN(new_n18752_));
  NOR2_X1    g15780(.A1(new_n18713_), .A2(new_n13114_), .ZN(new_n18753_));
  NOR2_X1    g15781(.A1(new_n18714_), .A2(new_n12014_), .ZN(new_n18754_));
  NOR2_X1    g15782(.A1(new_n18713_), .A2(new_n11961_), .ZN(new_n18755_));
  OAI21_X1   g15783(.A1(new_n15189_), .A2(new_n18722_), .B(new_n15884_), .ZN(new_n18756_));
  NOR2_X1    g15784(.A1(new_n13395_), .A2(new_n5324_), .ZN(new_n18757_));
  NOR2_X1    g15785(.A1(new_n18757_), .A2(pi0038), .ZN(new_n18758_));
  OAI22_X1   g15786(.A1(new_n18758_), .A2(new_n3232_), .B1(pi0180), .B2(new_n13399_), .ZN(new_n18759_));
  NOR2_X1    g15787(.A1(new_n3232_), .A2(pi0702), .ZN(new_n18760_));
  AOI22_X1   g15788(.A1(new_n18714_), .A2(new_n18760_), .B1(new_n18756_), .B2(new_n18759_), .ZN(new_n18761_));
  NOR3_X1    g15789(.A1(new_n18714_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n18762_));
  NOR4_X1    g15790(.A1(new_n18761_), .A2(new_n12970_), .A3(pi1153), .A4(new_n18713_), .ZN(new_n18763_));
  NOR2_X1    g15791(.A1(new_n18763_), .A2(new_n18762_), .ZN(new_n18764_));
  MUX2_X1    g15792(.I0(new_n18764_), .I1(new_n18761_), .S(new_n11891_), .Z(new_n18765_));
  INV_X1     g15793(.I(new_n18765_), .ZN(new_n18766_));
  NOR2_X1    g15794(.A1(new_n18714_), .A2(new_n11938_), .ZN(new_n18767_));
  AOI21_X1   g15795(.A1(new_n18766_), .A2(new_n11938_), .B(new_n18767_), .ZN(new_n18768_));
  AOI21_X1   g15796(.A1(new_n18768_), .A2(new_n11961_), .B(new_n18755_), .ZN(new_n18769_));
  AOI21_X1   g15797(.A1(new_n18769_), .A2(new_n12014_), .B(new_n18754_), .ZN(new_n18770_));
  AOI21_X1   g15798(.A1(new_n18770_), .A2(new_n13114_), .B(new_n18753_), .ZN(new_n18771_));
  NOR3_X1    g15799(.A1(new_n18714_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n18772_));
  NOR4_X1    g15800(.A1(new_n18771_), .A2(new_n12031_), .A3(pi1156), .A4(new_n18713_), .ZN(new_n18773_));
  NOR2_X1    g15801(.A1(new_n18773_), .A2(new_n18772_), .ZN(new_n18774_));
  MUX2_X1    g15802(.I0(new_n18774_), .I1(new_n18771_), .S(new_n11868_), .Z(new_n18775_));
  NOR2_X1    g15803(.A1(new_n18775_), .A2(new_n12061_), .ZN(new_n18776_));
  AOI21_X1   g15804(.A1(new_n12061_), .A2(new_n18713_), .B(new_n18776_), .ZN(new_n18777_));
  NAND2_X1   g15805(.A1(new_n18777_), .A2(pi1157), .ZN(new_n18778_));
  NOR2_X1    g15806(.A1(new_n18775_), .A2(pi0647), .ZN(new_n18779_));
  AOI21_X1   g15807(.A1(pi0647), .A2(new_n18713_), .B(new_n18779_), .ZN(new_n18780_));
  NAND2_X1   g15808(.A1(new_n18780_), .A2(new_n12049_), .ZN(new_n18781_));
  AOI21_X1   g15809(.A1(new_n18781_), .A2(new_n18778_), .B(new_n12048_), .ZN(new_n18782_));
  AOI21_X1   g15810(.A1(new_n12048_), .A2(new_n18775_), .B(new_n18782_), .ZN(new_n18783_));
  NAND2_X1   g15811(.A1(new_n18783_), .A2(pi0644), .ZN(new_n18784_));
  AOI21_X1   g15812(.A1(new_n18784_), .A2(new_n12099_), .B(new_n18752_), .ZN(new_n18785_));
  NAND3_X1   g15813(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n18786_));
  OAI21_X1   g15814(.A1(new_n18749_), .A2(new_n18786_), .B(pi0715), .ZN(new_n18787_));
  AOI21_X1   g15815(.A1(new_n18783_), .A2(new_n12082_), .B(new_n18787_), .ZN(new_n18788_));
  OAI21_X1   g15816(.A1(new_n18785_), .A2(new_n18788_), .B(pi0790), .ZN(new_n18789_));
  NAND2_X1   g15817(.A1(new_n18740_), .A2(pi0619), .ZN(new_n18790_));
  NAND2_X1   g15818(.A1(new_n18713_), .A2(pi0619), .ZN(new_n18791_));
  INV_X1     g15819(.I(new_n18763_), .ZN(new_n18792_));
  INV_X1     g15820(.I(new_n18727_), .ZN(new_n18793_));
  OR3_X2     g15821(.A1(new_n18725_), .A2(new_n15884_), .A3(new_n3231_), .Z(new_n18803_));
  OAI21_X1   g15822(.A1(new_n5324_), .A2(new_n3231_), .B(new_n18803_), .ZN(new_n18804_));
  OAI21_X1   g15823(.A1(new_n18804_), .A2(pi0625), .B(new_n18793_), .ZN(new_n18805_));
  NAND3_X1   g15824(.A1(new_n18804_), .A2(new_n12970_), .A3(new_n18727_), .ZN(new_n18806_));
  NAND4_X1   g15825(.A1(new_n18792_), .A2(new_n12977_), .A3(new_n18805_), .A4(new_n18806_), .ZN(new_n18807_));
  NOR4_X1    g15826(.A1(new_n18804_), .A2(new_n18793_), .A3(new_n12970_), .A4(pi1153), .ZN(new_n18808_));
  OAI21_X1   g15827(.A1(new_n18808_), .A2(new_n18762_), .B(new_n13657_), .ZN(new_n18809_));
  NAND2_X1   g15828(.A1(new_n18807_), .A2(new_n18809_), .ZN(new_n18810_));
  NOR2_X1    g15829(.A1(new_n18804_), .A2(pi0778), .ZN(new_n18811_));
  AOI21_X1   g15830(.A1(new_n18810_), .A2(pi0778), .B(new_n18811_), .ZN(new_n18812_));
  NOR2_X1    g15831(.A1(new_n18812_), .A2(pi0785), .ZN(new_n18813_));
  NAND3_X1   g15832(.A1(new_n18766_), .A2(pi0609), .A3(pi1155), .ZN(new_n18814_));
  NAND3_X1   g15833(.A1(new_n18814_), .A2(new_n11923_), .A3(new_n18734_), .ZN(new_n18815_));
  NAND2_X1   g15834(.A1(new_n18812_), .A2(pi0609), .ZN(new_n18816_));
  NAND3_X1   g15835(.A1(new_n18816_), .A2(new_n13621_), .A3(new_n18765_), .ZN(new_n18817_));
  NAND3_X1   g15836(.A1(new_n18817_), .A2(pi0660), .A3(new_n18732_), .ZN(new_n18818_));
  AND3_X2    g15837(.A1(new_n18818_), .A2(pi0785), .A3(new_n18815_), .Z(new_n18819_));
  NOR2_X1    g15838(.A1(new_n18819_), .A2(new_n18813_), .ZN(new_n18820_));
  NAND2_X1   g15839(.A1(new_n18820_), .A2(new_n11969_), .ZN(new_n18821_));
  NAND2_X1   g15840(.A1(new_n18820_), .A2(pi0618), .ZN(new_n18822_));
  AND2_X2    g15841(.A1(new_n18768_), .A2(new_n14633_), .Z(new_n18823_));
  NOR2_X1    g15842(.A1(new_n18736_), .A2(new_n11934_), .ZN(new_n18824_));
  OAI21_X1   g15843(.A1(new_n18714_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n18825_));
  OR3_X2     g15844(.A1(new_n18824_), .A2(new_n11949_), .A3(new_n18825_), .Z(new_n18826_));
  AOI21_X1   g15845(.A1(new_n18822_), .A2(new_n18823_), .B(new_n18826_), .ZN(new_n18827_));
  NOR3_X1    g15846(.A1(new_n18768_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n18828_));
  OAI21_X1   g15847(.A1(new_n18713_), .A2(pi0618), .B(new_n11950_), .ZN(new_n18829_));
  OAI21_X1   g15848(.A1(new_n18824_), .A2(new_n18829_), .B(new_n11949_), .ZN(new_n18830_));
  NOR2_X1    g15849(.A1(new_n18830_), .A2(new_n18828_), .ZN(new_n18831_));
  OAI21_X1   g15850(.A1(new_n18827_), .A2(new_n18831_), .B(pi0781), .ZN(new_n18832_));
  XOR2_X1    g15851(.A1(new_n18832_), .A2(new_n18821_), .Z(new_n18833_));
  XNOR2_X1   g15852(.A1(new_n18833_), .A2(new_n18769_), .ZN(new_n18834_));
  NOR2_X1    g15853(.A1(new_n18834_), .A2(new_n11967_), .ZN(new_n18835_));
  NAND3_X1   g15854(.A1(new_n18790_), .A2(new_n11869_), .A3(new_n18791_), .ZN(new_n18836_));
  XNOR2_X1   g15855(.A1(new_n18835_), .A2(new_n18833_), .ZN(new_n18837_));
  NAND2_X1   g15856(.A1(new_n18837_), .A2(new_n11869_), .ZN(new_n18838_));
  AOI21_X1   g15857(.A1(new_n18714_), .A2(new_n11967_), .B(pi1159), .ZN(new_n18839_));
  AOI21_X1   g15858(.A1(new_n18790_), .A2(new_n18839_), .B(pi0648), .ZN(new_n18840_));
  OAI21_X1   g15859(.A1(new_n18833_), .A2(pi0789), .B(new_n11998_), .ZN(new_n18841_));
  INV_X1     g15860(.I(new_n17372_), .ZN(new_n18842_));
  MUX2_X1    g15861(.I0(new_n18744_), .I1(new_n18713_), .S(new_n11994_), .Z(new_n18843_));
  NAND2_X1   g15862(.A1(new_n18843_), .A2(new_n11988_), .ZN(new_n18844_));
  AOI21_X1   g15863(.A1(new_n18744_), .A2(new_n18714_), .B(new_n11994_), .ZN(new_n18845_));
  OAI21_X1   g15864(.A1(new_n18770_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n18846_));
  AOI21_X1   g15865(.A1(new_n18845_), .A2(new_n11990_), .B(new_n18846_), .ZN(new_n18847_));
  AOI21_X1   g15866(.A1(new_n18844_), .A2(new_n18847_), .B(new_n18842_), .ZN(new_n18848_));
  NAND2_X1   g15867(.A1(new_n18841_), .A2(new_n18848_), .ZN(new_n18849_));
  AOI21_X1   g15868(.A1(new_n18838_), .A2(new_n18840_), .B(new_n18849_), .ZN(new_n18850_));
  NOR2_X1    g15869(.A1(new_n18772_), .A2(new_n12030_), .ZN(new_n18851_));
  NOR2_X1    g15870(.A1(new_n18773_), .A2(pi0629), .ZN(new_n18852_));
  NAND2_X1   g15871(.A1(new_n18745_), .A2(new_n15222_), .ZN(new_n18853_));
  OAI21_X1   g15872(.A1(new_n18851_), .A2(new_n18852_), .B(new_n18853_), .ZN(new_n18854_));
  AOI22_X1   g15873(.A1(new_n18850_), .A2(new_n18836_), .B1(pi0792), .B2(new_n18854_), .ZN(new_n18855_));
  NAND2_X1   g15874(.A1(new_n18777_), .A2(new_n12060_), .ZN(new_n18856_));
  AOI21_X1   g15875(.A1(new_n18780_), .A2(pi0630), .B(new_n15214_), .ZN(new_n18857_));
  NAND2_X1   g15876(.A1(new_n18857_), .A2(new_n18856_), .ZN(new_n18858_));
  NOR2_X1    g15877(.A1(new_n18747_), .A2(new_n15183_), .ZN(new_n18859_));
  OAI21_X1   g15878(.A1(new_n18749_), .A2(new_n18786_), .B(pi0644), .ZN(new_n18860_));
  NAND2_X1   g15879(.A1(new_n18860_), .A2(new_n11867_), .ZN(new_n18861_));
  AOI21_X1   g15880(.A1(new_n18752_), .A2(new_n12082_), .B(new_n18861_), .ZN(new_n18862_));
  AOI21_X1   g15881(.A1(new_n18858_), .A2(new_n18859_), .B(new_n18862_), .ZN(new_n18863_));
  OAI21_X1   g15882(.A1(new_n18855_), .A2(new_n14725_), .B(new_n18863_), .ZN(new_n18864_));
  AOI21_X1   g15883(.A1(new_n18864_), .A2(new_n18789_), .B(po1038), .ZN(new_n18865_));
  OAI21_X1   g15884(.A1(new_n6845_), .A2(pi0180), .B(new_n13184_), .ZN(new_n18866_));
  OAI21_X1   g15885(.A1(new_n18865_), .A2(new_n18866_), .B(new_n18712_), .ZN(po0337));
  NOR2_X1    g15886(.A1(new_n2925_), .A2(pi0181), .ZN(new_n18868_));
  NOR2_X1    g15887(.A1(new_n11877_), .A2(pi0754), .ZN(new_n18869_));
  NOR2_X1    g15888(.A1(new_n18869_), .A2(new_n18868_), .ZN(new_n18870_));
  AOI21_X1   g15889(.A1(new_n11886_), .A2(new_n15914_), .B(new_n18868_), .ZN(new_n18871_));
  NOR2_X1    g15890(.A1(new_n18871_), .A2(new_n11874_), .ZN(new_n18872_));
  INV_X1     g15891(.I(new_n18872_), .ZN(new_n18873_));
  NAND2_X1   g15892(.A1(new_n18873_), .A2(new_n18870_), .ZN(new_n18874_));
  NAND2_X1   g15893(.A1(new_n18874_), .A2(new_n11891_), .ZN(new_n18875_));
  NOR2_X1    g15894(.A1(new_n18873_), .A2(new_n12970_), .ZN(new_n18876_));
  NOR4_X1    g15895(.A1(new_n18876_), .A2(new_n11893_), .A3(new_n18868_), .A4(new_n18869_), .ZN(new_n18877_));
  NOR3_X1    g15896(.A1(new_n11894_), .A2(pi0625), .A3(pi0709), .ZN(new_n18878_));
  NOR2_X1    g15897(.A1(new_n18868_), .A2(pi1153), .ZN(new_n18879_));
  INV_X1     g15898(.I(new_n18879_), .ZN(new_n18880_));
  NOR2_X1    g15899(.A1(new_n18878_), .A2(new_n18880_), .ZN(new_n18881_));
  INV_X1     g15900(.I(new_n18881_), .ZN(new_n18882_));
  NAND2_X1   g15901(.A1(new_n18882_), .A2(pi0608), .ZN(new_n18883_));
  INV_X1     g15902(.I(new_n18876_), .ZN(new_n18884_));
  AOI21_X1   g15903(.A1(new_n18884_), .A2(new_n18874_), .B(new_n18880_), .ZN(new_n18885_));
  OAI21_X1   g15904(.A1(new_n18878_), .A2(new_n18871_), .B(pi1153), .ZN(new_n18886_));
  NAND2_X1   g15905(.A1(new_n18886_), .A2(new_n13657_), .ZN(new_n18887_));
  OAI22_X1   g15906(.A1(new_n18885_), .A2(new_n18887_), .B1(new_n18877_), .B2(new_n18883_), .ZN(new_n18888_));
  NAND2_X1   g15907(.A1(new_n18888_), .A2(pi0778), .ZN(new_n18889_));
  XOR2_X1    g15908(.A1(new_n18889_), .A2(new_n18875_), .Z(new_n18890_));
  INV_X1     g15909(.I(new_n18890_), .ZN(new_n18891_));
  NAND2_X1   g15910(.A1(new_n18882_), .A2(new_n18886_), .ZN(new_n18892_));
  MUX2_X1    g15911(.I0(new_n18892_), .I1(new_n18871_), .S(new_n11891_), .Z(new_n18893_));
  XNOR2_X1   g15912(.A1(new_n18890_), .A2(new_n18893_), .ZN(new_n18894_));
  NAND2_X1   g15913(.A1(new_n18894_), .A2(pi0609), .ZN(new_n18895_));
  XOR2_X1    g15914(.A1(new_n18895_), .A2(new_n18890_), .Z(new_n18896_));
  NAND2_X1   g15915(.A1(new_n18896_), .A2(new_n11912_), .ZN(new_n18897_));
  NOR2_X1    g15916(.A1(new_n18870_), .A2(new_n11925_), .ZN(new_n18898_));
  INV_X1     g15917(.I(new_n18898_), .ZN(new_n18899_));
  NOR3_X1    g15918(.A1(new_n12997_), .A2(new_n11877_), .A3(pi0754), .ZN(new_n18900_));
  NAND3_X1   g15919(.A1(new_n18899_), .A2(new_n11912_), .A3(new_n18900_), .ZN(new_n18901_));
  NAND3_X1   g15920(.A1(new_n18897_), .A2(new_n11923_), .A3(new_n18901_), .ZN(new_n18902_));
  NOR4_X1    g15921(.A1(new_n18900_), .A2(new_n11923_), .A3(pi1155), .A4(new_n18868_), .ZN(new_n18904_));
  NOR2_X1    g15922(.A1(new_n18904_), .A2(new_n11870_), .ZN(new_n18905_));
  AOI22_X1   g15923(.A1(new_n18902_), .A2(new_n18905_), .B1(new_n11870_), .B2(new_n18891_), .ZN(new_n18906_));
  NOR2_X1    g15924(.A1(new_n18906_), .A2(pi0781), .ZN(new_n18907_));
  NOR4_X1    g15925(.A1(new_n18893_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n18908_));
  NOR3_X1    g15926(.A1(new_n18900_), .A2(pi1155), .A3(new_n18868_), .ZN(new_n18909_));
  NAND2_X1   g15927(.A1(new_n18901_), .A2(new_n18909_), .ZN(new_n18910_));
  MUX2_X1    g15928(.I0(new_n18910_), .I1(new_n18899_), .S(new_n11870_), .Z(new_n18911_));
  INV_X1     g15929(.I(new_n18911_), .ZN(new_n18912_));
  OAI21_X1   g15930(.A1(new_n18912_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n18913_));
  OAI21_X1   g15931(.A1(new_n18912_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n18914_));
  NOR2_X1    g15932(.A1(new_n18893_), .A2(new_n11939_), .ZN(new_n18915_));
  NOR4_X1    g15933(.A1(new_n18906_), .A2(new_n11934_), .A3(pi1154), .A4(new_n18915_), .ZN(new_n18916_));
  NOR2_X1    g15934(.A1(new_n18916_), .A2(new_n18914_), .ZN(new_n18917_));
  OAI22_X1   g15935(.A1(new_n18917_), .A2(pi0627), .B1(new_n18908_), .B2(new_n18913_), .ZN(new_n18918_));
  AOI21_X1   g15936(.A1(new_n18918_), .A2(pi0781), .B(new_n18907_), .ZN(new_n18919_));
  INV_X1     g15937(.I(new_n18915_), .ZN(new_n18920_));
  NOR2_X1    g15938(.A1(new_n18920_), .A2(new_n11962_), .ZN(new_n18921_));
  NOR4_X1    g15939(.A1(new_n18919_), .A2(new_n11967_), .A3(pi1159), .A4(new_n18921_), .ZN(new_n18922_));
  NOR2_X1    g15940(.A1(new_n18912_), .A2(pi0781), .ZN(new_n18923_));
  AOI21_X1   g15941(.A1(new_n11944_), .A2(new_n18911_), .B(new_n18914_), .ZN(new_n18924_));
  NOR2_X1    g15942(.A1(new_n18924_), .A2(new_n11969_), .ZN(new_n18925_));
  XOR2_X1    g15943(.A1(new_n18925_), .A2(new_n18923_), .Z(new_n18926_));
  AOI21_X1   g15944(.A1(new_n18926_), .A2(new_n16479_), .B(pi1159), .ZN(new_n18927_));
  INV_X1     g15945(.I(new_n18927_), .ZN(new_n18928_));
  NOR3_X1    g15946(.A1(new_n18922_), .A2(new_n11966_), .A3(new_n18928_), .ZN(new_n18929_));
  NOR4_X1    g15947(.A1(new_n18920_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n18930_));
  INV_X1     g15948(.I(new_n18926_), .ZN(new_n18931_));
  NOR2_X1    g15949(.A1(new_n18931_), .A2(new_n16482_), .ZN(new_n18932_));
  NOR3_X1    g15950(.A1(new_n18932_), .A2(pi0648), .A3(new_n18930_), .ZN(new_n18933_));
  AOI21_X1   g15951(.A1(new_n18919_), .A2(new_n11998_), .B(pi0789), .ZN(new_n18934_));
  OAI21_X1   g15952(.A1(new_n18929_), .A2(new_n18933_), .B(new_n18934_), .ZN(new_n18935_));
  NAND2_X1   g15953(.A1(new_n18921_), .A2(new_n17450_), .ZN(new_n18936_));
  NOR2_X1    g15954(.A1(new_n18936_), .A2(new_n17153_), .ZN(new_n18937_));
  NOR2_X1    g15955(.A1(new_n14624_), .A2(new_n18868_), .ZN(new_n18938_));
  NOR2_X1    g15956(.A1(new_n18931_), .A2(pi0789), .ZN(new_n18939_));
  NOR2_X1    g15957(.A1(new_n18928_), .A2(new_n18932_), .ZN(new_n18940_));
  NOR2_X1    g15958(.A1(new_n18940_), .A2(new_n11985_), .ZN(new_n18941_));
  XOR2_X1    g15959(.A1(new_n18941_), .A2(new_n18939_), .Z(new_n18942_));
  AOI21_X1   g15960(.A1(new_n18942_), .A2(new_n14624_), .B(new_n18938_), .ZN(new_n18943_));
  AOI22_X1   g15961(.A1(new_n18943_), .A2(new_n12064_), .B1(new_n15080_), .B2(new_n18937_), .ZN(new_n18944_));
  NOR2_X1    g15962(.A1(new_n18944_), .A2(new_n12030_), .ZN(new_n18945_));
  NAND2_X1   g15963(.A1(new_n18943_), .A2(new_n12063_), .ZN(new_n18946_));
  AOI21_X1   g15964(.A1(new_n18937_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n18947_));
  NAND2_X1   g15965(.A1(new_n18946_), .A2(new_n18947_), .ZN(new_n18948_));
  OAI21_X1   g15966(.A1(new_n18945_), .A2(new_n18948_), .B(new_n14726_), .ZN(new_n18949_));
  INV_X1     g15967(.I(new_n18868_), .ZN(new_n18950_));
  MUX2_X1    g15968(.I0(new_n18942_), .I1(new_n18950_), .S(new_n11994_), .Z(new_n18951_));
  INV_X1     g15969(.I(new_n18942_), .ZN(new_n18952_));
  AOI21_X1   g15970(.A1(new_n18952_), .A2(new_n18950_), .B(new_n11994_), .ZN(new_n18953_));
  OAI21_X1   g15971(.A1(new_n18936_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n18954_));
  AOI21_X1   g15972(.A1(new_n18953_), .A2(new_n11990_), .B(new_n18954_), .ZN(new_n18955_));
  OAI21_X1   g15973(.A1(new_n17167_), .A2(new_n18951_), .B(new_n18955_), .ZN(new_n18956_));
  NAND4_X1   g15974(.A1(new_n18935_), .A2(new_n14732_), .A3(new_n18949_), .A4(new_n18956_), .ZN(new_n18957_));
  NAND3_X1   g15975(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n18868_), .ZN(new_n18958_));
  NAND2_X1   g15976(.A1(new_n18937_), .A2(new_n15050_), .ZN(new_n18959_));
  NAND2_X1   g15977(.A1(new_n18959_), .A2(pi0647), .ZN(new_n18960_));
  NAND2_X1   g15978(.A1(new_n18868_), .A2(pi0647), .ZN(new_n18961_));
  NAND3_X1   g15979(.A1(new_n18960_), .A2(new_n12049_), .A3(new_n18961_), .ZN(new_n18962_));
  NAND2_X1   g15980(.A1(new_n18962_), .A2(pi0630), .ZN(new_n18963_));
  NOR2_X1    g15981(.A1(new_n18959_), .A2(new_n12061_), .ZN(new_n18964_));
  AOI21_X1   g15982(.A1(new_n12061_), .A2(new_n18868_), .B(new_n18964_), .ZN(new_n18965_));
  NAND2_X1   g15983(.A1(new_n18965_), .A2(new_n12088_), .ZN(new_n18966_));
  NAND4_X1   g15984(.A1(new_n18966_), .A2(new_n18963_), .A3(pi0787), .A4(new_n18958_), .ZN(new_n18967_));
  AND2_X2    g15985(.A1(new_n18957_), .A2(new_n18967_), .Z(new_n18968_));
  NOR2_X1    g15986(.A1(new_n18968_), .A2(new_n12082_), .ZN(new_n18969_));
  NAND4_X1   g15987(.A1(new_n18960_), .A2(pi0787), .A3(new_n12049_), .A4(new_n18961_), .ZN(new_n18970_));
  OAI21_X1   g15988(.A1(pi0787), .A2(new_n18959_), .B(new_n18970_), .ZN(new_n18971_));
  NOR2_X1    g15989(.A1(new_n18971_), .A2(pi0644), .ZN(new_n18972_));
  OR3_X2     g15990(.A1(new_n18969_), .A2(pi0715), .A3(new_n18972_), .Z(new_n18973_));
  MUX2_X1    g15991(.I0(new_n18943_), .I1(new_n18868_), .S(new_n16841_), .Z(new_n18974_));
  INV_X1     g15992(.I(new_n18974_), .ZN(new_n18975_));
  OAI21_X1   g15993(.A1(new_n18974_), .A2(new_n18868_), .B(new_n12082_), .ZN(new_n18976_));
  AOI21_X1   g15994(.A1(new_n18868_), .A2(new_n18974_), .B(new_n18976_), .ZN(new_n18977_));
  OAI21_X1   g15995(.A1(new_n18977_), .A2(new_n18975_), .B(new_n12099_), .ZN(new_n18978_));
  AOI21_X1   g15996(.A1(new_n18975_), .A2(new_n18977_), .B(new_n18978_), .ZN(new_n18979_));
  AOI21_X1   g15997(.A1(new_n18973_), .A2(new_n18979_), .B(pi1160), .ZN(new_n18980_));
  XOR2_X1    g15998(.A1(new_n18977_), .A2(new_n18868_), .Z(new_n18981_));
  AOI21_X1   g15999(.A1(new_n18971_), .A2(pi0644), .B(new_n13169_), .ZN(new_n18982_));
  OAI21_X1   g16000(.A1(new_n18981_), .A2(new_n12099_), .B(new_n18982_), .ZN(new_n18983_));
  OAI21_X1   g16001(.A1(new_n18969_), .A2(new_n18983_), .B(pi0790), .ZN(new_n18984_));
  NOR2_X1    g16002(.A1(new_n18968_), .A2(new_n14748_), .ZN(new_n18985_));
  OAI21_X1   g16003(.A1(new_n18980_), .A2(new_n18984_), .B(new_n18985_), .ZN(new_n18986_));
  NOR2_X1    g16004(.A1(new_n12965_), .A2(pi0181), .ZN(new_n18987_));
  INV_X1     g16005(.I(new_n18987_), .ZN(new_n18988_));
  NAND2_X1   g16006(.A1(new_n18988_), .A2(new_n11997_), .ZN(new_n18989_));
  NAND2_X1   g16007(.A1(new_n12894_), .A2(pi0754), .ZN(new_n18990_));
  NOR2_X1    g16008(.A1(new_n15896_), .A2(pi0181), .ZN(new_n18991_));
  OAI21_X1   g16009(.A1(new_n14361_), .A2(new_n5325_), .B(pi0039), .ZN(new_n18994_));
  AOI21_X1   g16010(.A1(new_n12824_), .A2(new_n18991_), .B(new_n18994_), .ZN(new_n18995_));
  NOR2_X1    g16011(.A1(new_n12828_), .A2(pi0181), .ZN(new_n18996_));
  AOI21_X1   g16012(.A1(new_n12829_), .A2(new_n15896_), .B(pi0038), .ZN(new_n18997_));
  INV_X1     g16013(.I(new_n18997_), .ZN(new_n18998_));
  AOI21_X1   g16014(.A1(new_n18995_), .A2(new_n18990_), .B(new_n18998_), .ZN(new_n18999_));
  NOR2_X1    g16015(.A1(new_n18999_), .A2(new_n3232_), .ZN(new_n19000_));
  AOI21_X1   g16016(.A1(new_n5325_), .A2(new_n3232_), .B(new_n19000_), .ZN(new_n19001_));
  OAI21_X1   g16017(.A1(new_n19001_), .A2(new_n11914_), .B(new_n11870_), .ZN(new_n19002_));
  AOI21_X1   g16018(.A1(new_n11914_), .A2(new_n18987_), .B(new_n19002_), .ZN(new_n19003_));
  NAND2_X1   g16019(.A1(new_n19001_), .A2(new_n11924_), .ZN(new_n19004_));
  OAI22_X1   g16020(.A1(new_n19004_), .A2(pi0609), .B1(new_n12996_), .B2(new_n18987_), .ZN(new_n19005_));
  NAND2_X1   g16021(.A1(new_n19005_), .A2(new_n11912_), .ZN(new_n19006_));
  OAI22_X1   g16022(.A1(new_n19004_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n18987_), .ZN(new_n19007_));
  NAND2_X1   g16023(.A1(new_n19007_), .A2(pi1155), .ZN(new_n19008_));
  AOI21_X1   g16024(.A1(new_n19006_), .A2(new_n19008_), .B(new_n11870_), .ZN(new_n19009_));
  XNOR2_X1   g16025(.A1(new_n19009_), .A2(new_n19003_), .ZN(new_n19010_));
  NOR2_X1    g16026(.A1(new_n19010_), .A2(pi0781), .ZN(new_n19011_));
  NOR3_X1    g16027(.A1(new_n18987_), .A2(pi0618), .A3(pi1154), .ZN(new_n19012_));
  NOR2_X1    g16028(.A1(new_n19012_), .A2(new_n11969_), .ZN(new_n19013_));
  XOR2_X1    g16029(.A1(new_n19011_), .A2(new_n19013_), .Z(new_n19014_));
  NAND2_X1   g16030(.A1(new_n19014_), .A2(new_n11985_), .ZN(new_n19015_));
  NAND3_X1   g16031(.A1(new_n18988_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n19016_));
  NAND2_X1   g16032(.A1(new_n19016_), .A2(pi0789), .ZN(new_n19017_));
  XNOR2_X1   g16033(.A1(new_n19015_), .A2(new_n19017_), .ZN(new_n19018_));
  OAI21_X1   g16034(.A1(new_n19018_), .A2(new_n11997_), .B(new_n18989_), .ZN(new_n19019_));
  NOR2_X1    g16035(.A1(new_n18987_), .A2(new_n12054_), .ZN(new_n19020_));
  AOI21_X1   g16036(.A1(new_n19019_), .A2(new_n12054_), .B(new_n19020_), .ZN(new_n19021_));
  NAND2_X1   g16037(.A1(new_n18988_), .A2(new_n12091_), .ZN(new_n19022_));
  OAI21_X1   g16038(.A1(new_n19021_), .A2(new_n12091_), .B(new_n19022_), .ZN(new_n19023_));
  OR2_X2     g16039(.A1(new_n19023_), .A2(pi0644), .Z(new_n19024_));
  AOI21_X1   g16040(.A1(new_n18987_), .A2(pi0644), .B(new_n12099_), .ZN(new_n19025_));
  AOI21_X1   g16041(.A1(new_n19024_), .A2(new_n19025_), .B(pi1160), .ZN(new_n19026_));
  NOR2_X1    g16042(.A1(new_n18987_), .A2(new_n13114_), .ZN(new_n19027_));
  NOR2_X1    g16043(.A1(new_n18988_), .A2(new_n12014_), .ZN(new_n19028_));
  NOR2_X1    g16044(.A1(new_n18987_), .A2(new_n11961_), .ZN(new_n19029_));
  OAI21_X1   g16045(.A1(new_n15189_), .A2(new_n18996_), .B(new_n15914_), .ZN(new_n19030_));
  NOR2_X1    g16046(.A1(new_n13395_), .A2(new_n5325_), .ZN(new_n19031_));
  NOR2_X1    g16047(.A1(new_n19031_), .A2(pi0038), .ZN(new_n19032_));
  OAI22_X1   g16048(.A1(new_n19032_), .A2(new_n3232_), .B1(pi0181), .B2(new_n13399_), .ZN(new_n19033_));
  NOR2_X1    g16049(.A1(new_n3232_), .A2(pi0709), .ZN(new_n19034_));
  AOI22_X1   g16050(.A1(new_n18988_), .A2(new_n19034_), .B1(new_n19030_), .B2(new_n19033_), .ZN(new_n19035_));
  NOR3_X1    g16051(.A1(new_n18988_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n19036_));
  NOR4_X1    g16052(.A1(new_n19035_), .A2(new_n12970_), .A3(pi1153), .A4(new_n18987_), .ZN(new_n19037_));
  NOR2_X1    g16053(.A1(new_n19037_), .A2(new_n19036_), .ZN(new_n19038_));
  MUX2_X1    g16054(.I0(new_n19038_), .I1(new_n19035_), .S(new_n11891_), .Z(new_n19039_));
  INV_X1     g16055(.I(new_n19039_), .ZN(new_n19040_));
  NOR2_X1    g16056(.A1(new_n18988_), .A2(new_n11938_), .ZN(new_n19041_));
  AOI21_X1   g16057(.A1(new_n19040_), .A2(new_n11938_), .B(new_n19041_), .ZN(new_n19042_));
  AOI21_X1   g16058(.A1(new_n19042_), .A2(new_n11961_), .B(new_n19029_), .ZN(new_n19043_));
  AOI21_X1   g16059(.A1(new_n19043_), .A2(new_n12014_), .B(new_n19028_), .ZN(new_n19044_));
  AOI21_X1   g16060(.A1(new_n19044_), .A2(new_n13114_), .B(new_n19027_), .ZN(new_n19045_));
  NOR3_X1    g16061(.A1(new_n18988_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n19046_));
  NOR4_X1    g16062(.A1(new_n19045_), .A2(new_n12031_), .A3(pi1156), .A4(new_n18987_), .ZN(new_n19047_));
  NOR2_X1    g16063(.A1(new_n19047_), .A2(new_n19046_), .ZN(new_n19048_));
  MUX2_X1    g16064(.I0(new_n19048_), .I1(new_n19045_), .S(new_n11868_), .Z(new_n19049_));
  NOR2_X1    g16065(.A1(new_n19049_), .A2(new_n12061_), .ZN(new_n19050_));
  AOI21_X1   g16066(.A1(new_n12061_), .A2(new_n18987_), .B(new_n19050_), .ZN(new_n19051_));
  NAND2_X1   g16067(.A1(new_n19051_), .A2(pi1157), .ZN(new_n19052_));
  NOR2_X1    g16068(.A1(new_n19049_), .A2(pi0647), .ZN(new_n19053_));
  AOI21_X1   g16069(.A1(pi0647), .A2(new_n18987_), .B(new_n19053_), .ZN(new_n19054_));
  NAND2_X1   g16070(.A1(new_n19054_), .A2(new_n12049_), .ZN(new_n19055_));
  AOI21_X1   g16071(.A1(new_n19055_), .A2(new_n19052_), .B(new_n12048_), .ZN(new_n19056_));
  AOI21_X1   g16072(.A1(new_n12048_), .A2(new_n19049_), .B(new_n19056_), .ZN(new_n19057_));
  NAND2_X1   g16073(.A1(new_n19057_), .A2(pi0644), .ZN(new_n19058_));
  AOI21_X1   g16074(.A1(new_n19058_), .A2(new_n12099_), .B(new_n19026_), .ZN(new_n19059_));
  NAND3_X1   g16075(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n19060_));
  OAI21_X1   g16076(.A1(new_n19023_), .A2(new_n19060_), .B(pi0715), .ZN(new_n19061_));
  AOI21_X1   g16077(.A1(new_n19057_), .A2(new_n12082_), .B(new_n19061_), .ZN(new_n19062_));
  OAI21_X1   g16078(.A1(new_n19059_), .A2(new_n19062_), .B(pi0790), .ZN(new_n19063_));
  NAND2_X1   g16079(.A1(new_n19014_), .A2(pi0619), .ZN(new_n19064_));
  NAND2_X1   g16080(.A1(new_n18987_), .A2(pi0619), .ZN(new_n19065_));
  INV_X1     g16081(.I(new_n19037_), .ZN(new_n19066_));
  INV_X1     g16082(.I(new_n19001_), .ZN(new_n19067_));
  OR3_X2     g16083(.A1(new_n18999_), .A2(new_n15914_), .A3(new_n3231_), .Z(new_n19077_));
  OAI21_X1   g16084(.A1(new_n5325_), .A2(new_n3231_), .B(new_n19077_), .ZN(new_n19078_));
  OAI21_X1   g16085(.A1(new_n19078_), .A2(pi0625), .B(new_n19067_), .ZN(new_n19079_));
  NAND3_X1   g16086(.A1(new_n19078_), .A2(new_n12970_), .A3(new_n19001_), .ZN(new_n19080_));
  NAND4_X1   g16087(.A1(new_n19066_), .A2(new_n12977_), .A3(new_n19079_), .A4(new_n19080_), .ZN(new_n19081_));
  NOR4_X1    g16088(.A1(new_n19078_), .A2(new_n19067_), .A3(new_n12970_), .A4(pi1153), .ZN(new_n19082_));
  OAI21_X1   g16089(.A1(new_n19082_), .A2(new_n19036_), .B(new_n13657_), .ZN(new_n19083_));
  NAND2_X1   g16090(.A1(new_n19081_), .A2(new_n19083_), .ZN(new_n19084_));
  NOR2_X1    g16091(.A1(new_n19078_), .A2(pi0778), .ZN(new_n19085_));
  AOI21_X1   g16092(.A1(new_n19084_), .A2(pi0778), .B(new_n19085_), .ZN(new_n19086_));
  NOR2_X1    g16093(.A1(new_n19086_), .A2(pi0785), .ZN(new_n19087_));
  NAND3_X1   g16094(.A1(new_n19040_), .A2(pi0609), .A3(pi1155), .ZN(new_n19088_));
  NAND3_X1   g16095(.A1(new_n19088_), .A2(new_n11923_), .A3(new_n19008_), .ZN(new_n19089_));
  NAND2_X1   g16096(.A1(new_n19086_), .A2(pi0609), .ZN(new_n19090_));
  NAND3_X1   g16097(.A1(new_n19090_), .A2(new_n13621_), .A3(new_n19039_), .ZN(new_n19091_));
  NAND3_X1   g16098(.A1(new_n19091_), .A2(pi0660), .A3(new_n19006_), .ZN(new_n19092_));
  AND3_X2    g16099(.A1(new_n19092_), .A2(pi0785), .A3(new_n19089_), .Z(new_n19093_));
  NOR2_X1    g16100(.A1(new_n19093_), .A2(new_n19087_), .ZN(new_n19094_));
  NAND2_X1   g16101(.A1(new_n19094_), .A2(new_n11969_), .ZN(new_n19095_));
  NAND2_X1   g16102(.A1(new_n19094_), .A2(pi0618), .ZN(new_n19096_));
  AND2_X2    g16103(.A1(new_n19042_), .A2(new_n14633_), .Z(new_n19097_));
  NOR2_X1    g16104(.A1(new_n19010_), .A2(new_n11934_), .ZN(new_n19098_));
  OAI21_X1   g16105(.A1(new_n18988_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n19099_));
  OR3_X2     g16106(.A1(new_n19098_), .A2(new_n11949_), .A3(new_n19099_), .Z(new_n19100_));
  AOI21_X1   g16107(.A1(new_n19096_), .A2(new_n19097_), .B(new_n19100_), .ZN(new_n19101_));
  NOR3_X1    g16108(.A1(new_n19042_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n19102_));
  OAI21_X1   g16109(.A1(new_n18987_), .A2(pi0618), .B(new_n11950_), .ZN(new_n19103_));
  OAI21_X1   g16110(.A1(new_n19098_), .A2(new_n19103_), .B(new_n11949_), .ZN(new_n19104_));
  NOR2_X1    g16111(.A1(new_n19104_), .A2(new_n19102_), .ZN(new_n19105_));
  OAI21_X1   g16112(.A1(new_n19101_), .A2(new_n19105_), .B(pi0781), .ZN(new_n19106_));
  XOR2_X1    g16113(.A1(new_n19106_), .A2(new_n19095_), .Z(new_n19107_));
  XNOR2_X1   g16114(.A1(new_n19107_), .A2(new_n19043_), .ZN(new_n19108_));
  NOR2_X1    g16115(.A1(new_n19108_), .A2(new_n11967_), .ZN(new_n19109_));
  NAND3_X1   g16116(.A1(new_n19064_), .A2(new_n11869_), .A3(new_n19065_), .ZN(new_n19110_));
  XNOR2_X1   g16117(.A1(new_n19109_), .A2(new_n19107_), .ZN(new_n19111_));
  NAND2_X1   g16118(.A1(new_n19111_), .A2(new_n11869_), .ZN(new_n19112_));
  AOI21_X1   g16119(.A1(new_n18988_), .A2(new_n11967_), .B(pi1159), .ZN(new_n19113_));
  AOI21_X1   g16120(.A1(new_n19064_), .A2(new_n19113_), .B(pi0648), .ZN(new_n19114_));
  OAI21_X1   g16121(.A1(new_n19107_), .A2(pi0789), .B(new_n11998_), .ZN(new_n19115_));
  MUX2_X1    g16122(.I0(new_n19018_), .I1(new_n18987_), .S(new_n11994_), .Z(new_n19116_));
  NAND2_X1   g16123(.A1(new_n19116_), .A2(new_n11988_), .ZN(new_n19117_));
  AOI21_X1   g16124(.A1(new_n19018_), .A2(new_n18988_), .B(new_n11994_), .ZN(new_n19118_));
  OAI21_X1   g16125(.A1(new_n19044_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n19119_));
  AOI21_X1   g16126(.A1(new_n19118_), .A2(new_n11990_), .B(new_n19119_), .ZN(new_n19120_));
  AOI21_X1   g16127(.A1(new_n19117_), .A2(new_n19120_), .B(new_n18842_), .ZN(new_n19121_));
  NAND2_X1   g16128(.A1(new_n19115_), .A2(new_n19121_), .ZN(new_n19122_));
  AOI21_X1   g16129(.A1(new_n19112_), .A2(new_n19114_), .B(new_n19122_), .ZN(new_n19123_));
  NOR2_X1    g16130(.A1(new_n19046_), .A2(new_n12030_), .ZN(new_n19124_));
  NOR2_X1    g16131(.A1(new_n19047_), .A2(pi0629), .ZN(new_n19125_));
  NAND2_X1   g16132(.A1(new_n19019_), .A2(new_n15222_), .ZN(new_n19126_));
  OAI21_X1   g16133(.A1(new_n19124_), .A2(new_n19125_), .B(new_n19126_), .ZN(new_n19127_));
  AOI22_X1   g16134(.A1(new_n19123_), .A2(new_n19110_), .B1(pi0792), .B2(new_n19127_), .ZN(new_n19128_));
  NAND2_X1   g16135(.A1(new_n19051_), .A2(new_n12060_), .ZN(new_n19129_));
  AOI21_X1   g16136(.A1(new_n19054_), .A2(pi0630), .B(new_n15214_), .ZN(new_n19130_));
  NAND2_X1   g16137(.A1(new_n19130_), .A2(new_n19129_), .ZN(new_n19131_));
  NOR2_X1    g16138(.A1(new_n19021_), .A2(new_n15183_), .ZN(new_n19132_));
  OAI21_X1   g16139(.A1(new_n19023_), .A2(new_n19060_), .B(pi0644), .ZN(new_n19133_));
  NAND2_X1   g16140(.A1(new_n19133_), .A2(new_n11867_), .ZN(new_n19134_));
  AOI21_X1   g16141(.A1(new_n19026_), .A2(new_n12082_), .B(new_n19134_), .ZN(new_n19135_));
  AOI21_X1   g16142(.A1(new_n19131_), .A2(new_n19132_), .B(new_n19135_), .ZN(new_n19136_));
  OAI21_X1   g16143(.A1(new_n19128_), .A2(new_n14725_), .B(new_n19136_), .ZN(new_n19137_));
  AOI21_X1   g16144(.A1(new_n19137_), .A2(new_n19063_), .B(po1038), .ZN(new_n19138_));
  OAI21_X1   g16145(.A1(new_n6845_), .A2(pi0181), .B(new_n13184_), .ZN(new_n19139_));
  OAI21_X1   g16146(.A1(new_n19138_), .A2(new_n19139_), .B(new_n18986_), .ZN(po0338));
  NOR2_X1    g16147(.A1(new_n2925_), .A2(pi0182), .ZN(new_n19141_));
  NOR2_X1    g16148(.A1(new_n11877_), .A2(pi0756), .ZN(new_n19142_));
  NOR2_X1    g16149(.A1(new_n19142_), .A2(new_n19141_), .ZN(new_n19143_));
  AOI21_X1   g16150(.A1(new_n11886_), .A2(new_n15949_), .B(new_n19141_), .ZN(new_n19144_));
  NOR2_X1    g16151(.A1(new_n19144_), .A2(new_n11874_), .ZN(new_n19145_));
  INV_X1     g16152(.I(new_n19145_), .ZN(new_n19146_));
  NAND2_X1   g16153(.A1(new_n19146_), .A2(new_n19143_), .ZN(new_n19147_));
  NAND2_X1   g16154(.A1(new_n19147_), .A2(new_n11891_), .ZN(new_n19148_));
  NOR2_X1    g16155(.A1(new_n19146_), .A2(new_n12970_), .ZN(new_n19149_));
  NOR4_X1    g16156(.A1(new_n19149_), .A2(new_n11893_), .A3(new_n19141_), .A4(new_n19142_), .ZN(new_n19150_));
  NOR3_X1    g16157(.A1(new_n11894_), .A2(pi0625), .A3(pi0734), .ZN(new_n19151_));
  NOR2_X1    g16158(.A1(new_n19141_), .A2(pi1153), .ZN(new_n19152_));
  INV_X1     g16159(.I(new_n19152_), .ZN(new_n19153_));
  NOR2_X1    g16160(.A1(new_n19151_), .A2(new_n19153_), .ZN(new_n19154_));
  INV_X1     g16161(.I(new_n19154_), .ZN(new_n19155_));
  NAND2_X1   g16162(.A1(new_n19155_), .A2(pi0608), .ZN(new_n19156_));
  INV_X1     g16163(.I(new_n19149_), .ZN(new_n19157_));
  AOI21_X1   g16164(.A1(new_n19157_), .A2(new_n19147_), .B(new_n19153_), .ZN(new_n19158_));
  OAI21_X1   g16165(.A1(new_n19151_), .A2(new_n19144_), .B(pi1153), .ZN(new_n19159_));
  NAND2_X1   g16166(.A1(new_n19159_), .A2(new_n13657_), .ZN(new_n19160_));
  OAI22_X1   g16167(.A1(new_n19158_), .A2(new_n19160_), .B1(new_n19150_), .B2(new_n19156_), .ZN(new_n19161_));
  NAND2_X1   g16168(.A1(new_n19161_), .A2(pi0778), .ZN(new_n19162_));
  XOR2_X1    g16169(.A1(new_n19162_), .A2(new_n19148_), .Z(new_n19163_));
  INV_X1     g16170(.I(new_n19163_), .ZN(new_n19164_));
  NAND2_X1   g16171(.A1(new_n19155_), .A2(new_n19159_), .ZN(new_n19165_));
  MUX2_X1    g16172(.I0(new_n19165_), .I1(new_n19144_), .S(new_n11891_), .Z(new_n19166_));
  XNOR2_X1   g16173(.A1(new_n19163_), .A2(new_n19166_), .ZN(new_n19167_));
  NAND2_X1   g16174(.A1(new_n19167_), .A2(pi0609), .ZN(new_n19168_));
  XOR2_X1    g16175(.A1(new_n19168_), .A2(new_n19163_), .Z(new_n19169_));
  NAND2_X1   g16176(.A1(new_n19169_), .A2(new_n11912_), .ZN(new_n19170_));
  NOR2_X1    g16177(.A1(new_n19143_), .A2(new_n11925_), .ZN(new_n19171_));
  INV_X1     g16178(.I(new_n19171_), .ZN(new_n19172_));
  NOR3_X1    g16179(.A1(new_n12997_), .A2(new_n11877_), .A3(pi0756), .ZN(new_n19173_));
  NAND3_X1   g16180(.A1(new_n19172_), .A2(new_n11912_), .A3(new_n19173_), .ZN(new_n19174_));
  NAND3_X1   g16181(.A1(new_n19170_), .A2(new_n11923_), .A3(new_n19174_), .ZN(new_n19175_));
  NOR4_X1    g16182(.A1(new_n19173_), .A2(new_n11923_), .A3(pi1155), .A4(new_n19141_), .ZN(new_n19177_));
  NOR2_X1    g16183(.A1(new_n19177_), .A2(new_n11870_), .ZN(new_n19178_));
  AOI22_X1   g16184(.A1(new_n19175_), .A2(new_n19178_), .B1(new_n11870_), .B2(new_n19164_), .ZN(new_n19179_));
  NOR2_X1    g16185(.A1(new_n19179_), .A2(pi0781), .ZN(new_n19180_));
  NOR4_X1    g16186(.A1(new_n19166_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n19181_));
  NOR3_X1    g16187(.A1(new_n19173_), .A2(pi1155), .A3(new_n19141_), .ZN(new_n19182_));
  NAND2_X1   g16188(.A1(new_n19174_), .A2(new_n19182_), .ZN(new_n19183_));
  MUX2_X1    g16189(.I0(new_n19183_), .I1(new_n19172_), .S(new_n11870_), .Z(new_n19184_));
  INV_X1     g16190(.I(new_n19184_), .ZN(new_n19185_));
  OAI21_X1   g16191(.A1(new_n19185_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n19186_));
  OAI21_X1   g16192(.A1(new_n19185_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n19187_));
  NOR2_X1    g16193(.A1(new_n19166_), .A2(new_n11939_), .ZN(new_n19188_));
  NOR4_X1    g16194(.A1(new_n19179_), .A2(new_n11934_), .A3(pi1154), .A4(new_n19188_), .ZN(new_n19189_));
  NOR2_X1    g16195(.A1(new_n19189_), .A2(new_n19187_), .ZN(new_n19190_));
  OAI22_X1   g16196(.A1(new_n19190_), .A2(pi0627), .B1(new_n19181_), .B2(new_n19186_), .ZN(new_n19191_));
  AOI21_X1   g16197(.A1(new_n19191_), .A2(pi0781), .B(new_n19180_), .ZN(new_n19192_));
  INV_X1     g16198(.I(new_n19188_), .ZN(new_n19193_));
  NOR2_X1    g16199(.A1(new_n19193_), .A2(new_n11962_), .ZN(new_n19194_));
  NOR4_X1    g16200(.A1(new_n19192_), .A2(new_n11967_), .A3(pi1159), .A4(new_n19194_), .ZN(new_n19195_));
  NOR2_X1    g16201(.A1(new_n19185_), .A2(pi0781), .ZN(new_n19196_));
  AOI21_X1   g16202(.A1(new_n11944_), .A2(new_n19184_), .B(new_n19187_), .ZN(new_n19197_));
  NOR2_X1    g16203(.A1(new_n19197_), .A2(new_n11969_), .ZN(new_n19198_));
  XOR2_X1    g16204(.A1(new_n19198_), .A2(new_n19196_), .Z(new_n19199_));
  AOI21_X1   g16205(.A1(new_n19199_), .A2(new_n16479_), .B(pi1159), .ZN(new_n19200_));
  INV_X1     g16206(.I(new_n19200_), .ZN(new_n19201_));
  NOR3_X1    g16207(.A1(new_n19195_), .A2(new_n11966_), .A3(new_n19201_), .ZN(new_n19202_));
  NOR4_X1    g16208(.A1(new_n19193_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n19203_));
  INV_X1     g16209(.I(new_n19199_), .ZN(new_n19204_));
  NOR2_X1    g16210(.A1(new_n19204_), .A2(new_n16482_), .ZN(new_n19205_));
  NOR3_X1    g16211(.A1(new_n19205_), .A2(pi0648), .A3(new_n19203_), .ZN(new_n19206_));
  AOI21_X1   g16212(.A1(new_n19192_), .A2(new_n11998_), .B(pi0789), .ZN(new_n19207_));
  OAI21_X1   g16213(.A1(new_n19202_), .A2(new_n19206_), .B(new_n19207_), .ZN(new_n19208_));
  NAND2_X1   g16214(.A1(new_n19194_), .A2(new_n17450_), .ZN(new_n19209_));
  NOR2_X1    g16215(.A1(new_n19209_), .A2(new_n17153_), .ZN(new_n19210_));
  NOR2_X1    g16216(.A1(new_n14624_), .A2(new_n19141_), .ZN(new_n19211_));
  NOR2_X1    g16217(.A1(new_n19204_), .A2(pi0789), .ZN(new_n19212_));
  NOR2_X1    g16218(.A1(new_n19201_), .A2(new_n19205_), .ZN(new_n19213_));
  NOR2_X1    g16219(.A1(new_n19213_), .A2(new_n11985_), .ZN(new_n19214_));
  XOR2_X1    g16220(.A1(new_n19214_), .A2(new_n19212_), .Z(new_n19215_));
  AOI21_X1   g16221(.A1(new_n19215_), .A2(new_n14624_), .B(new_n19211_), .ZN(new_n19216_));
  AOI22_X1   g16222(.A1(new_n19216_), .A2(new_n12064_), .B1(new_n15080_), .B2(new_n19210_), .ZN(new_n19217_));
  NOR2_X1    g16223(.A1(new_n19217_), .A2(new_n12030_), .ZN(new_n19218_));
  NAND2_X1   g16224(.A1(new_n19216_), .A2(new_n12063_), .ZN(new_n19219_));
  AOI21_X1   g16225(.A1(new_n19210_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n19220_));
  NAND2_X1   g16226(.A1(new_n19219_), .A2(new_n19220_), .ZN(new_n19221_));
  OAI21_X1   g16227(.A1(new_n19218_), .A2(new_n19221_), .B(new_n14726_), .ZN(new_n19222_));
  INV_X1     g16228(.I(new_n19141_), .ZN(new_n19223_));
  MUX2_X1    g16229(.I0(new_n19215_), .I1(new_n19223_), .S(new_n11994_), .Z(new_n19224_));
  INV_X1     g16230(.I(new_n19215_), .ZN(new_n19225_));
  AOI21_X1   g16231(.A1(new_n19225_), .A2(new_n19223_), .B(new_n11994_), .ZN(new_n19226_));
  OAI21_X1   g16232(.A1(new_n19209_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n19227_));
  AOI21_X1   g16233(.A1(new_n19226_), .A2(new_n11990_), .B(new_n19227_), .ZN(new_n19228_));
  OAI21_X1   g16234(.A1(new_n17167_), .A2(new_n19224_), .B(new_n19228_), .ZN(new_n19229_));
  NAND4_X1   g16235(.A1(new_n19208_), .A2(new_n14732_), .A3(new_n19222_), .A4(new_n19229_), .ZN(new_n19230_));
  NAND3_X1   g16236(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n19141_), .ZN(new_n19231_));
  NAND2_X1   g16237(.A1(new_n19210_), .A2(new_n15050_), .ZN(new_n19232_));
  NAND2_X1   g16238(.A1(new_n19232_), .A2(pi0647), .ZN(new_n19233_));
  NAND2_X1   g16239(.A1(new_n19141_), .A2(pi0647), .ZN(new_n19234_));
  NAND3_X1   g16240(.A1(new_n19233_), .A2(new_n12049_), .A3(new_n19234_), .ZN(new_n19235_));
  NAND2_X1   g16241(.A1(new_n19235_), .A2(pi0630), .ZN(new_n19236_));
  NOR2_X1    g16242(.A1(new_n19232_), .A2(new_n12061_), .ZN(new_n19237_));
  AOI21_X1   g16243(.A1(new_n12061_), .A2(new_n19141_), .B(new_n19237_), .ZN(new_n19238_));
  NAND2_X1   g16244(.A1(new_n19238_), .A2(new_n12088_), .ZN(new_n19239_));
  NAND4_X1   g16245(.A1(new_n19239_), .A2(new_n19236_), .A3(pi0787), .A4(new_n19231_), .ZN(new_n19240_));
  AND2_X2    g16246(.A1(new_n19230_), .A2(new_n19240_), .Z(new_n19241_));
  NOR2_X1    g16247(.A1(new_n19241_), .A2(new_n12082_), .ZN(new_n19242_));
  NAND4_X1   g16248(.A1(new_n19233_), .A2(pi0787), .A3(new_n12049_), .A4(new_n19234_), .ZN(new_n19243_));
  OAI21_X1   g16249(.A1(pi0787), .A2(new_n19232_), .B(new_n19243_), .ZN(new_n19244_));
  NOR2_X1    g16250(.A1(new_n19244_), .A2(pi0644), .ZN(new_n19245_));
  OR3_X2     g16251(.A1(new_n19242_), .A2(pi0715), .A3(new_n19245_), .Z(new_n19246_));
  MUX2_X1    g16252(.I0(new_n19216_), .I1(new_n19141_), .S(new_n16841_), .Z(new_n19247_));
  INV_X1     g16253(.I(new_n19247_), .ZN(new_n19248_));
  OAI21_X1   g16254(.A1(new_n19247_), .A2(new_n19141_), .B(new_n12082_), .ZN(new_n19249_));
  AOI21_X1   g16255(.A1(new_n19141_), .A2(new_n19247_), .B(new_n19249_), .ZN(new_n19250_));
  OAI21_X1   g16256(.A1(new_n19250_), .A2(new_n19248_), .B(new_n12099_), .ZN(new_n19251_));
  AOI21_X1   g16257(.A1(new_n19248_), .A2(new_n19250_), .B(new_n19251_), .ZN(new_n19252_));
  AOI21_X1   g16258(.A1(new_n19246_), .A2(new_n19252_), .B(pi1160), .ZN(new_n19253_));
  XOR2_X1    g16259(.A1(new_n19250_), .A2(new_n19141_), .Z(new_n19254_));
  AOI21_X1   g16260(.A1(new_n19244_), .A2(pi0644), .B(new_n13169_), .ZN(new_n19255_));
  OAI21_X1   g16261(.A1(new_n19254_), .A2(new_n12099_), .B(new_n19255_), .ZN(new_n19256_));
  OAI21_X1   g16262(.A1(new_n19242_), .A2(new_n19256_), .B(pi0790), .ZN(new_n19257_));
  NOR2_X1    g16263(.A1(new_n19241_), .A2(new_n14748_), .ZN(new_n19258_));
  OAI21_X1   g16264(.A1(new_n19253_), .A2(new_n19257_), .B(new_n19258_), .ZN(new_n19259_));
  NOR2_X1    g16265(.A1(new_n12965_), .A2(pi0182), .ZN(new_n19260_));
  INV_X1     g16266(.I(new_n19260_), .ZN(new_n19261_));
  NAND2_X1   g16267(.A1(new_n19261_), .A2(new_n11997_), .ZN(new_n19262_));
  AOI21_X1   g16268(.A1(new_n12794_), .A2(new_n5326_), .B(pi0756), .ZN(new_n19263_));
  NAND3_X1   g16269(.A1(new_n13381_), .A2(new_n5326_), .A3(new_n14362_), .ZN(new_n19264_));
  OAI21_X1   g16270(.A1(new_n13381_), .A2(pi0182), .B(new_n12694_), .ZN(new_n19265_));
  NAND3_X1   g16271(.A1(new_n19265_), .A2(new_n19264_), .A3(new_n15926_), .ZN(new_n19266_));
  NOR2_X1    g16272(.A1(new_n19266_), .A2(new_n19263_), .ZN(new_n19267_));
  NOR2_X1    g16273(.A1(new_n12828_), .A2(pi0182), .ZN(new_n19268_));
  OAI21_X1   g16274(.A1(new_n13367_), .A2(pi0756), .B(pi0038), .ZN(new_n19269_));
  OAI22_X1   g16275(.A1(new_n19267_), .A2(pi0038), .B1(new_n19268_), .B2(new_n19269_), .ZN(new_n19270_));
  NOR2_X1    g16276(.A1(new_n19270_), .A2(new_n3232_), .ZN(new_n19271_));
  AOI21_X1   g16277(.A1(new_n5326_), .A2(new_n3232_), .B(new_n19271_), .ZN(new_n19272_));
  INV_X1     g16278(.I(new_n19272_), .ZN(new_n19273_));
  OAI21_X1   g16279(.A1(new_n19261_), .A2(new_n11924_), .B(new_n11870_), .ZN(new_n19274_));
  AOI21_X1   g16280(.A1(new_n19273_), .A2(new_n11924_), .B(new_n19274_), .ZN(new_n19275_));
  NAND2_X1   g16281(.A1(new_n19272_), .A2(new_n11924_), .ZN(new_n19276_));
  OAI22_X1   g16282(.A1(new_n19276_), .A2(pi0609), .B1(new_n12996_), .B2(new_n19260_), .ZN(new_n19277_));
  NAND2_X1   g16283(.A1(new_n19277_), .A2(new_n11912_), .ZN(new_n19278_));
  OAI22_X1   g16284(.A1(new_n19276_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n19260_), .ZN(new_n19279_));
  NAND2_X1   g16285(.A1(new_n19279_), .A2(pi1155), .ZN(new_n19280_));
  AOI21_X1   g16286(.A1(new_n19278_), .A2(new_n19280_), .B(new_n11870_), .ZN(new_n19281_));
  XOR2_X1    g16287(.A1(new_n19281_), .A2(new_n19275_), .Z(new_n19282_));
  OAI21_X1   g16288(.A1(new_n19261_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n19283_));
  AOI21_X1   g16289(.A1(new_n19282_), .A2(pi0618), .B(new_n19283_), .ZN(new_n19284_));
  NAND2_X1   g16290(.A1(new_n19282_), .A2(pi0618), .ZN(new_n19285_));
  AOI21_X1   g16291(.A1(new_n19261_), .A2(new_n11934_), .B(pi1154), .ZN(new_n19286_));
  NAND2_X1   g16292(.A1(new_n19285_), .A2(new_n19286_), .ZN(new_n19287_));
  NAND2_X1   g16293(.A1(new_n19287_), .A2(new_n19284_), .ZN(new_n19288_));
  MUX2_X1    g16294(.I0(new_n19288_), .I1(new_n19282_), .S(new_n11969_), .Z(new_n19289_));
  NAND2_X1   g16295(.A1(new_n19289_), .A2(new_n11985_), .ZN(new_n19290_));
  NOR3_X1    g16296(.A1(new_n19260_), .A2(pi0619), .A3(pi1159), .ZN(new_n19291_));
  NOR2_X1    g16297(.A1(new_n19291_), .A2(new_n11985_), .ZN(new_n19292_));
  XOR2_X1    g16298(.A1(new_n19290_), .A2(new_n19292_), .Z(new_n19293_));
  OAI21_X1   g16299(.A1(new_n19293_), .A2(new_n11997_), .B(new_n19262_), .ZN(new_n19294_));
  NOR2_X1    g16300(.A1(new_n19260_), .A2(new_n12054_), .ZN(new_n19295_));
  AOI21_X1   g16301(.A1(new_n19294_), .A2(new_n12054_), .B(new_n19295_), .ZN(new_n19296_));
  NAND2_X1   g16302(.A1(new_n19261_), .A2(new_n12091_), .ZN(new_n19297_));
  OAI21_X1   g16303(.A1(new_n19296_), .A2(new_n12091_), .B(new_n19297_), .ZN(new_n19298_));
  AOI21_X1   g16304(.A1(new_n19260_), .A2(pi0644), .B(new_n12099_), .ZN(new_n19299_));
  OAI21_X1   g16305(.A1(new_n19298_), .A2(pi0644), .B(new_n19299_), .ZN(new_n19300_));
  AND2_X2    g16306(.A1(new_n19300_), .A2(new_n12081_), .Z(new_n19301_));
  NOR2_X1    g16307(.A1(new_n19261_), .A2(pi0647), .ZN(new_n19302_));
  NOR2_X1    g16308(.A1(new_n19260_), .A2(new_n13114_), .ZN(new_n19303_));
  NOR2_X1    g16309(.A1(new_n19261_), .A2(new_n12014_), .ZN(new_n19304_));
  NOR2_X1    g16310(.A1(new_n19260_), .A2(new_n11961_), .ZN(new_n19305_));
  OAI21_X1   g16311(.A1(new_n15189_), .A2(new_n19268_), .B(new_n15949_), .ZN(new_n19306_));
  NOR2_X1    g16312(.A1(new_n13395_), .A2(new_n5326_), .ZN(new_n19307_));
  NOR2_X1    g16313(.A1(new_n19307_), .A2(pi0038), .ZN(new_n19308_));
  OAI22_X1   g16314(.A1(new_n19308_), .A2(new_n3232_), .B1(pi0182), .B2(new_n13399_), .ZN(new_n19309_));
  NOR2_X1    g16315(.A1(new_n3232_), .A2(pi0734), .ZN(new_n19310_));
  AOI22_X1   g16316(.A1(new_n19261_), .A2(new_n19310_), .B1(new_n19306_), .B2(new_n19309_), .ZN(new_n19311_));
  NOR3_X1    g16317(.A1(new_n19261_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n19312_));
  NOR4_X1    g16318(.A1(new_n19311_), .A2(new_n12970_), .A3(pi1153), .A4(new_n19260_), .ZN(new_n19313_));
  NOR2_X1    g16319(.A1(new_n19313_), .A2(new_n19312_), .ZN(new_n19314_));
  MUX2_X1    g16320(.I0(new_n19314_), .I1(new_n19311_), .S(new_n11891_), .Z(new_n19315_));
  NOR2_X1    g16321(.A1(new_n19315_), .A2(new_n13024_), .ZN(new_n19316_));
  AOI21_X1   g16322(.A1(new_n13024_), .A2(new_n19260_), .B(new_n19316_), .ZN(new_n19317_));
  AOI21_X1   g16323(.A1(new_n19317_), .A2(new_n11961_), .B(new_n19305_), .ZN(new_n19318_));
  AOI21_X1   g16324(.A1(new_n19318_), .A2(new_n12014_), .B(new_n19304_), .ZN(new_n19319_));
  AOI21_X1   g16325(.A1(new_n19319_), .A2(new_n13114_), .B(new_n19303_), .ZN(new_n19320_));
  INV_X1     g16326(.I(new_n19320_), .ZN(new_n19321_));
  NAND3_X1   g16327(.A1(new_n19260_), .A2(pi0628), .A3(pi1156), .ZN(new_n19322_));
  NOR4_X1    g16328(.A1(new_n19320_), .A2(new_n12031_), .A3(pi1156), .A4(new_n19260_), .ZN(new_n19323_));
  INV_X1     g16329(.I(new_n19323_), .ZN(new_n19324_));
  NAND2_X1   g16330(.A1(new_n19324_), .A2(new_n19322_), .ZN(new_n19325_));
  MUX2_X1    g16331(.I0(new_n19325_), .I1(new_n19321_), .S(new_n11868_), .Z(new_n19326_));
  AOI21_X1   g16332(.A1(new_n19326_), .A2(pi0647), .B(new_n19302_), .ZN(new_n19327_));
  NAND2_X1   g16333(.A1(new_n19327_), .A2(pi1157), .ZN(new_n19328_));
  NOR2_X1    g16334(.A1(new_n19261_), .A2(new_n12061_), .ZN(new_n19329_));
  AOI21_X1   g16335(.A1(new_n19326_), .A2(new_n12061_), .B(new_n19329_), .ZN(new_n19330_));
  NAND2_X1   g16336(.A1(new_n19330_), .A2(new_n12049_), .ZN(new_n19331_));
  NAND2_X1   g16337(.A1(new_n19328_), .A2(new_n19331_), .ZN(new_n19332_));
  NOR2_X1    g16338(.A1(new_n19326_), .A2(pi0787), .ZN(new_n19333_));
  AOI21_X1   g16339(.A1(new_n19332_), .A2(pi0787), .B(new_n19333_), .ZN(new_n19334_));
  AOI21_X1   g16340(.A1(new_n19334_), .A2(pi0644), .B(pi0715), .ZN(new_n19335_));
  NOR2_X1    g16341(.A1(new_n19301_), .A2(new_n19335_), .ZN(new_n19336_));
  NAND3_X1   g16342(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n19337_));
  OR2_X2     g16343(.A1(new_n19298_), .A2(new_n19337_), .Z(new_n19338_));
  NAND2_X1   g16344(.A1(new_n19338_), .A2(pi0715), .ZN(new_n19339_));
  AOI21_X1   g16345(.A1(new_n12082_), .A2(new_n19334_), .B(new_n19339_), .ZN(new_n19340_));
  OAI21_X1   g16346(.A1(new_n19340_), .A2(new_n19336_), .B(pi0790), .ZN(new_n19341_));
  NAND2_X1   g16347(.A1(new_n19289_), .A2(pi0619), .ZN(new_n19342_));
  NAND2_X1   g16348(.A1(new_n19260_), .A2(pi0619), .ZN(new_n19343_));
  NOR3_X1    g16349(.A1(new_n19270_), .A2(new_n15949_), .A3(new_n3231_), .ZN(new_n19353_));
  AOI21_X1   g16350(.A1(pi0182), .A2(new_n3232_), .B(new_n19353_), .ZN(new_n19354_));
  INV_X1     g16351(.I(new_n19313_), .ZN(new_n19355_));
  NAND2_X1   g16352(.A1(new_n19354_), .A2(pi0625), .ZN(new_n19356_));
  NAND2_X1   g16353(.A1(new_n19273_), .A2(pi0625), .ZN(new_n19357_));
  NAND4_X1   g16354(.A1(new_n19357_), .A2(new_n12977_), .A3(new_n19355_), .A4(new_n19356_), .ZN(new_n19358_));
  NAND2_X1   g16355(.A1(new_n19272_), .A2(new_n12970_), .ZN(new_n19359_));
  AND3_X2    g16356(.A1(new_n19356_), .A2(new_n11893_), .A3(new_n19359_), .Z(new_n19360_));
  OAI21_X1   g16357(.A1(new_n19360_), .A2(new_n19312_), .B(new_n13657_), .ZN(new_n19361_));
  AOI21_X1   g16358(.A1(new_n19361_), .A2(new_n19358_), .B(new_n11891_), .ZN(new_n19362_));
  AOI21_X1   g16359(.A1(new_n11891_), .A2(new_n19354_), .B(new_n19362_), .ZN(new_n19363_));
  NOR2_X1    g16360(.A1(new_n19363_), .A2(pi0785), .ZN(new_n19364_));
  INV_X1     g16361(.I(new_n19315_), .ZN(new_n19365_));
  NAND3_X1   g16362(.A1(new_n19365_), .A2(pi0609), .A3(pi1155), .ZN(new_n19366_));
  NAND3_X1   g16363(.A1(new_n19366_), .A2(new_n11923_), .A3(new_n19280_), .ZN(new_n19367_));
  NOR4_X1    g16364(.A1(new_n19363_), .A2(new_n11903_), .A3(pi1155), .A4(new_n19365_), .ZN(new_n19368_));
  NAND2_X1   g16365(.A1(new_n19278_), .A2(pi0660), .ZN(new_n19369_));
  NOR2_X1    g16366(.A1(new_n19368_), .A2(new_n19369_), .ZN(new_n19370_));
  NOR2_X1    g16367(.A1(new_n19370_), .A2(new_n11870_), .ZN(new_n19371_));
  AOI21_X1   g16368(.A1(new_n19371_), .A2(new_n19367_), .B(new_n19364_), .ZN(new_n19372_));
  INV_X1     g16369(.I(new_n19317_), .ZN(new_n19373_));
  NOR4_X1    g16370(.A1(new_n19372_), .A2(new_n11934_), .A3(pi1154), .A4(new_n19373_), .ZN(new_n19374_));
  NAND2_X1   g16371(.A1(new_n19284_), .A2(pi0627), .ZN(new_n19375_));
  NOR3_X1    g16372(.A1(new_n19317_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n19376_));
  NAND2_X1   g16373(.A1(new_n19287_), .A2(new_n11949_), .ZN(new_n19377_));
  OAI22_X1   g16374(.A1(new_n19374_), .A2(new_n19375_), .B1(new_n19376_), .B2(new_n19377_), .ZN(new_n19378_));
  MUX2_X1    g16375(.I0(new_n19378_), .I1(new_n19372_), .S(new_n11969_), .Z(new_n19379_));
  XNOR2_X1   g16376(.A1(new_n19379_), .A2(new_n19318_), .ZN(new_n19380_));
  NOR2_X1    g16377(.A1(new_n19380_), .A2(new_n11967_), .ZN(new_n19381_));
  NAND3_X1   g16378(.A1(new_n19342_), .A2(new_n11869_), .A3(new_n19343_), .ZN(new_n19382_));
  XNOR2_X1   g16379(.A1(new_n19381_), .A2(new_n19379_), .ZN(new_n19383_));
  NAND2_X1   g16380(.A1(new_n19383_), .A2(new_n11869_), .ZN(new_n19384_));
  AOI21_X1   g16381(.A1(new_n19261_), .A2(new_n11967_), .B(pi1159), .ZN(new_n19385_));
  AOI21_X1   g16382(.A1(new_n19342_), .A2(new_n19385_), .B(pi0648), .ZN(new_n19386_));
  INV_X1     g16383(.I(new_n19293_), .ZN(new_n19387_));
  MUX2_X1    g16384(.I0(new_n19387_), .I1(new_n19261_), .S(new_n11994_), .Z(new_n19388_));
  AOI21_X1   g16385(.A1(new_n19293_), .A2(new_n19261_), .B(new_n11994_), .ZN(new_n19389_));
  OAI21_X1   g16386(.A1(new_n19319_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n19390_));
  AOI21_X1   g16387(.A1(new_n19389_), .A2(new_n11990_), .B(new_n19390_), .ZN(new_n19391_));
  OAI21_X1   g16388(.A1(new_n19388_), .A2(new_n17167_), .B(new_n19391_), .ZN(new_n19392_));
  OAI21_X1   g16389(.A1(new_n19379_), .A2(pi0789), .B(new_n11998_), .ZN(new_n19393_));
  NAND3_X1   g16390(.A1(new_n19392_), .A2(new_n17372_), .A3(new_n19393_), .ZN(new_n19394_));
  AOI21_X1   g16391(.A1(new_n19384_), .A2(new_n19386_), .B(new_n19394_), .ZN(new_n19395_));
  NAND2_X1   g16392(.A1(new_n19322_), .A2(pi0629), .ZN(new_n19396_));
  OAI21_X1   g16393(.A1(new_n19323_), .A2(pi0629), .B(new_n19396_), .ZN(new_n19397_));
  NAND2_X1   g16394(.A1(new_n19294_), .A2(new_n15222_), .ZN(new_n19398_));
  NAND2_X1   g16395(.A1(new_n19398_), .A2(new_n19397_), .ZN(new_n19399_));
  AOI22_X1   g16396(.A1(new_n19395_), .A2(new_n19382_), .B1(pi0792), .B2(new_n19399_), .ZN(new_n19400_));
  NAND2_X1   g16397(.A1(new_n19327_), .A2(new_n12060_), .ZN(new_n19401_));
  AOI21_X1   g16398(.A1(new_n19330_), .A2(pi0630), .B(new_n15214_), .ZN(new_n19402_));
  NAND2_X1   g16399(.A1(new_n19402_), .A2(new_n19401_), .ZN(new_n19403_));
  NOR2_X1    g16400(.A1(new_n19296_), .A2(new_n15183_), .ZN(new_n19404_));
  NAND2_X1   g16401(.A1(new_n19301_), .A2(new_n12082_), .ZN(new_n19405_));
  AOI21_X1   g16402(.A1(new_n19338_), .A2(pi0644), .B(pi0790), .ZN(new_n19406_));
  AOI22_X1   g16403(.A1(new_n19405_), .A2(new_n19406_), .B1(new_n19403_), .B2(new_n19404_), .ZN(new_n19407_));
  OAI21_X1   g16404(.A1(new_n19400_), .A2(new_n14725_), .B(new_n19407_), .ZN(new_n19408_));
  AOI21_X1   g16405(.A1(new_n19408_), .A2(new_n19341_), .B(po1038), .ZN(new_n19409_));
  OAI21_X1   g16406(.A1(new_n6845_), .A2(pi0182), .B(new_n13184_), .ZN(new_n19410_));
  OAI21_X1   g16407(.A1(new_n19409_), .A2(new_n19410_), .B(new_n19259_), .ZN(po0339));
  NOR2_X1    g16408(.A1(new_n2925_), .A2(pi0183), .ZN(new_n19412_));
  NOR2_X1    g16409(.A1(new_n11877_), .A2(pi0755), .ZN(new_n19413_));
  NOR2_X1    g16410(.A1(new_n19413_), .A2(new_n19412_), .ZN(new_n19414_));
  AOI21_X1   g16411(.A1(new_n11886_), .A2(new_n15535_), .B(new_n19412_), .ZN(new_n19415_));
  NOR2_X1    g16412(.A1(new_n19415_), .A2(new_n11874_), .ZN(new_n19416_));
  INV_X1     g16413(.I(new_n19416_), .ZN(new_n19417_));
  NAND2_X1   g16414(.A1(new_n19417_), .A2(new_n19414_), .ZN(new_n19418_));
  NAND2_X1   g16415(.A1(new_n19418_), .A2(new_n11891_), .ZN(new_n19419_));
  NOR2_X1    g16416(.A1(new_n19417_), .A2(new_n12970_), .ZN(new_n19420_));
  NOR4_X1    g16417(.A1(new_n19420_), .A2(new_n11893_), .A3(new_n19412_), .A4(new_n19413_), .ZN(new_n19421_));
  NOR3_X1    g16418(.A1(new_n11894_), .A2(pi0625), .A3(pi0725), .ZN(new_n19422_));
  NOR2_X1    g16419(.A1(new_n19412_), .A2(pi1153), .ZN(new_n19423_));
  INV_X1     g16420(.I(new_n19423_), .ZN(new_n19424_));
  NOR2_X1    g16421(.A1(new_n19422_), .A2(new_n19424_), .ZN(new_n19425_));
  INV_X1     g16422(.I(new_n19425_), .ZN(new_n19426_));
  NAND2_X1   g16423(.A1(new_n19426_), .A2(pi0608), .ZN(new_n19427_));
  INV_X1     g16424(.I(new_n19420_), .ZN(new_n19428_));
  AOI21_X1   g16425(.A1(new_n19428_), .A2(new_n19418_), .B(new_n19424_), .ZN(new_n19429_));
  OAI21_X1   g16426(.A1(new_n19422_), .A2(new_n19415_), .B(pi1153), .ZN(new_n19430_));
  NAND2_X1   g16427(.A1(new_n19430_), .A2(new_n13657_), .ZN(new_n19431_));
  OAI22_X1   g16428(.A1(new_n19429_), .A2(new_n19431_), .B1(new_n19421_), .B2(new_n19427_), .ZN(new_n19432_));
  NAND2_X1   g16429(.A1(new_n19432_), .A2(pi0778), .ZN(new_n19433_));
  XOR2_X1    g16430(.A1(new_n19433_), .A2(new_n19419_), .Z(new_n19434_));
  INV_X1     g16431(.I(new_n19434_), .ZN(new_n19435_));
  NAND2_X1   g16432(.A1(new_n19426_), .A2(new_n19430_), .ZN(new_n19436_));
  MUX2_X1    g16433(.I0(new_n19436_), .I1(new_n19415_), .S(new_n11891_), .Z(new_n19437_));
  XNOR2_X1   g16434(.A1(new_n19434_), .A2(new_n19437_), .ZN(new_n19438_));
  NAND2_X1   g16435(.A1(new_n19438_), .A2(pi0609), .ZN(new_n19439_));
  XOR2_X1    g16436(.A1(new_n19439_), .A2(new_n19434_), .Z(new_n19440_));
  NAND2_X1   g16437(.A1(new_n19440_), .A2(new_n11912_), .ZN(new_n19441_));
  NOR2_X1    g16438(.A1(new_n19414_), .A2(new_n11925_), .ZN(new_n19442_));
  INV_X1     g16439(.I(new_n19442_), .ZN(new_n19443_));
  NOR3_X1    g16440(.A1(new_n12997_), .A2(new_n11877_), .A3(pi0755), .ZN(new_n19444_));
  NAND3_X1   g16441(.A1(new_n19443_), .A2(new_n11912_), .A3(new_n19444_), .ZN(new_n19445_));
  NAND3_X1   g16442(.A1(new_n19441_), .A2(new_n11923_), .A3(new_n19445_), .ZN(new_n19446_));
  NOR4_X1    g16443(.A1(new_n19444_), .A2(new_n11923_), .A3(pi1155), .A4(new_n19412_), .ZN(new_n19448_));
  NOR2_X1    g16444(.A1(new_n19448_), .A2(new_n11870_), .ZN(new_n19449_));
  AOI22_X1   g16445(.A1(new_n19446_), .A2(new_n19449_), .B1(new_n11870_), .B2(new_n19435_), .ZN(new_n19450_));
  NOR2_X1    g16446(.A1(new_n19450_), .A2(pi0781), .ZN(new_n19451_));
  NOR4_X1    g16447(.A1(new_n19437_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n19452_));
  NOR3_X1    g16448(.A1(new_n19444_), .A2(pi1155), .A3(new_n19412_), .ZN(new_n19453_));
  NAND2_X1   g16449(.A1(new_n19445_), .A2(new_n19453_), .ZN(new_n19454_));
  MUX2_X1    g16450(.I0(new_n19454_), .I1(new_n19443_), .S(new_n11870_), .Z(new_n19455_));
  INV_X1     g16451(.I(new_n19455_), .ZN(new_n19456_));
  OAI21_X1   g16452(.A1(new_n19456_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n19457_));
  OAI21_X1   g16453(.A1(new_n19456_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n19458_));
  NOR2_X1    g16454(.A1(new_n19437_), .A2(new_n11939_), .ZN(new_n19459_));
  NOR4_X1    g16455(.A1(new_n19450_), .A2(new_n11934_), .A3(pi1154), .A4(new_n19459_), .ZN(new_n19460_));
  NOR2_X1    g16456(.A1(new_n19460_), .A2(new_n19458_), .ZN(new_n19461_));
  OAI22_X1   g16457(.A1(new_n19461_), .A2(pi0627), .B1(new_n19452_), .B2(new_n19457_), .ZN(new_n19462_));
  AOI21_X1   g16458(.A1(new_n19462_), .A2(pi0781), .B(new_n19451_), .ZN(new_n19463_));
  INV_X1     g16459(.I(new_n19459_), .ZN(new_n19464_));
  NOR2_X1    g16460(.A1(new_n19464_), .A2(new_n11962_), .ZN(new_n19465_));
  NOR4_X1    g16461(.A1(new_n19463_), .A2(new_n11967_), .A3(pi1159), .A4(new_n19465_), .ZN(new_n19466_));
  NOR2_X1    g16462(.A1(new_n19456_), .A2(pi0781), .ZN(new_n19467_));
  AOI21_X1   g16463(.A1(new_n11944_), .A2(new_n19455_), .B(new_n19458_), .ZN(new_n19468_));
  NOR2_X1    g16464(.A1(new_n19468_), .A2(new_n11969_), .ZN(new_n19469_));
  XOR2_X1    g16465(.A1(new_n19469_), .A2(new_n19467_), .Z(new_n19470_));
  AOI21_X1   g16466(.A1(new_n19470_), .A2(new_n16479_), .B(pi1159), .ZN(new_n19471_));
  INV_X1     g16467(.I(new_n19471_), .ZN(new_n19472_));
  NOR3_X1    g16468(.A1(new_n19466_), .A2(new_n11966_), .A3(new_n19472_), .ZN(new_n19473_));
  NOR4_X1    g16469(.A1(new_n19464_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n19474_));
  INV_X1     g16470(.I(new_n19470_), .ZN(new_n19475_));
  NOR2_X1    g16471(.A1(new_n19475_), .A2(new_n16482_), .ZN(new_n19476_));
  NOR3_X1    g16472(.A1(new_n19476_), .A2(pi0648), .A3(new_n19474_), .ZN(new_n19477_));
  AOI21_X1   g16473(.A1(new_n19463_), .A2(new_n11998_), .B(pi0789), .ZN(new_n19478_));
  OAI21_X1   g16474(.A1(new_n19473_), .A2(new_n19477_), .B(new_n19478_), .ZN(new_n19479_));
  NAND2_X1   g16475(.A1(new_n19465_), .A2(new_n17450_), .ZN(new_n19480_));
  NOR2_X1    g16476(.A1(new_n19480_), .A2(new_n17153_), .ZN(new_n19481_));
  NOR2_X1    g16477(.A1(new_n14624_), .A2(new_n19412_), .ZN(new_n19482_));
  NOR2_X1    g16478(.A1(new_n19475_), .A2(pi0789), .ZN(new_n19483_));
  NOR2_X1    g16479(.A1(new_n19472_), .A2(new_n19476_), .ZN(new_n19484_));
  NOR2_X1    g16480(.A1(new_n19484_), .A2(new_n11985_), .ZN(new_n19485_));
  XOR2_X1    g16481(.A1(new_n19485_), .A2(new_n19483_), .Z(new_n19486_));
  AOI21_X1   g16482(.A1(new_n19486_), .A2(new_n14624_), .B(new_n19482_), .ZN(new_n19487_));
  AOI22_X1   g16483(.A1(new_n19487_), .A2(new_n12064_), .B1(new_n15080_), .B2(new_n19481_), .ZN(new_n19488_));
  NOR2_X1    g16484(.A1(new_n19488_), .A2(new_n12030_), .ZN(new_n19489_));
  NAND2_X1   g16485(.A1(new_n19487_), .A2(new_n12063_), .ZN(new_n19490_));
  AOI21_X1   g16486(.A1(new_n19481_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n19491_));
  NAND2_X1   g16487(.A1(new_n19490_), .A2(new_n19491_), .ZN(new_n19492_));
  OAI21_X1   g16488(.A1(new_n19489_), .A2(new_n19492_), .B(new_n14726_), .ZN(new_n19493_));
  INV_X1     g16489(.I(new_n19412_), .ZN(new_n19494_));
  MUX2_X1    g16490(.I0(new_n19486_), .I1(new_n19494_), .S(new_n11994_), .Z(new_n19495_));
  INV_X1     g16491(.I(new_n19486_), .ZN(new_n19496_));
  AOI21_X1   g16492(.A1(new_n19496_), .A2(new_n19494_), .B(new_n11994_), .ZN(new_n19497_));
  OAI21_X1   g16493(.A1(new_n19480_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n19498_));
  AOI21_X1   g16494(.A1(new_n19497_), .A2(new_n11990_), .B(new_n19498_), .ZN(new_n19499_));
  OAI21_X1   g16495(.A1(new_n17167_), .A2(new_n19495_), .B(new_n19499_), .ZN(new_n19500_));
  NAND4_X1   g16496(.A1(new_n19479_), .A2(new_n14732_), .A3(new_n19493_), .A4(new_n19500_), .ZN(new_n19501_));
  NAND3_X1   g16497(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n19412_), .ZN(new_n19502_));
  NAND2_X1   g16498(.A1(new_n19481_), .A2(new_n15050_), .ZN(new_n19503_));
  NAND2_X1   g16499(.A1(new_n19503_), .A2(pi0647), .ZN(new_n19504_));
  NAND2_X1   g16500(.A1(new_n19412_), .A2(pi0647), .ZN(new_n19505_));
  NAND3_X1   g16501(.A1(new_n19504_), .A2(new_n12049_), .A3(new_n19505_), .ZN(new_n19506_));
  NAND2_X1   g16502(.A1(new_n19506_), .A2(pi0630), .ZN(new_n19507_));
  NOR2_X1    g16503(.A1(new_n19503_), .A2(new_n12061_), .ZN(new_n19508_));
  AOI21_X1   g16504(.A1(new_n12061_), .A2(new_n19412_), .B(new_n19508_), .ZN(new_n19509_));
  NAND2_X1   g16505(.A1(new_n19509_), .A2(new_n12088_), .ZN(new_n19510_));
  NAND4_X1   g16506(.A1(new_n19510_), .A2(new_n19507_), .A3(pi0787), .A4(new_n19502_), .ZN(new_n19511_));
  AND2_X2    g16507(.A1(new_n19501_), .A2(new_n19511_), .Z(new_n19512_));
  NOR2_X1    g16508(.A1(new_n19512_), .A2(new_n12082_), .ZN(new_n19513_));
  NAND4_X1   g16509(.A1(new_n19504_), .A2(pi0787), .A3(new_n12049_), .A4(new_n19505_), .ZN(new_n19514_));
  OAI21_X1   g16510(.A1(pi0787), .A2(new_n19503_), .B(new_n19514_), .ZN(new_n19515_));
  NOR2_X1    g16511(.A1(new_n19515_), .A2(pi0644), .ZN(new_n19516_));
  OR3_X2     g16512(.A1(new_n19513_), .A2(pi0715), .A3(new_n19516_), .Z(new_n19517_));
  MUX2_X1    g16513(.I0(new_n19487_), .I1(new_n19412_), .S(new_n16841_), .Z(new_n19518_));
  INV_X1     g16514(.I(new_n19518_), .ZN(new_n19519_));
  OAI21_X1   g16515(.A1(new_n19518_), .A2(new_n19412_), .B(new_n12082_), .ZN(new_n19520_));
  AOI21_X1   g16516(.A1(new_n19412_), .A2(new_n19518_), .B(new_n19520_), .ZN(new_n19521_));
  OAI21_X1   g16517(.A1(new_n19521_), .A2(new_n19519_), .B(new_n12099_), .ZN(new_n19522_));
  AOI21_X1   g16518(.A1(new_n19519_), .A2(new_n19521_), .B(new_n19522_), .ZN(new_n19523_));
  AOI21_X1   g16519(.A1(new_n19517_), .A2(new_n19523_), .B(pi1160), .ZN(new_n19524_));
  XOR2_X1    g16520(.A1(new_n19521_), .A2(new_n19412_), .Z(new_n19525_));
  AOI21_X1   g16521(.A1(new_n19515_), .A2(pi0644), .B(new_n13169_), .ZN(new_n19526_));
  OAI21_X1   g16522(.A1(new_n19525_), .A2(new_n12099_), .B(new_n19526_), .ZN(new_n19527_));
  OAI21_X1   g16523(.A1(new_n19513_), .A2(new_n19527_), .B(pi0790), .ZN(new_n19528_));
  NOR2_X1    g16524(.A1(new_n19512_), .A2(new_n14748_), .ZN(new_n19529_));
  OAI21_X1   g16525(.A1(new_n19524_), .A2(new_n19528_), .B(new_n19529_), .ZN(new_n19530_));
  NOR2_X1    g16526(.A1(new_n12965_), .A2(pi0183), .ZN(new_n19531_));
  INV_X1     g16527(.I(new_n19531_), .ZN(new_n19532_));
  NAND2_X1   g16528(.A1(new_n19532_), .A2(new_n11997_), .ZN(new_n19533_));
  AOI21_X1   g16529(.A1(new_n12794_), .A2(new_n7180_), .B(pi0755), .ZN(new_n19534_));
  NAND3_X1   g16530(.A1(new_n13381_), .A2(new_n7180_), .A3(new_n14362_), .ZN(new_n19535_));
  OAI21_X1   g16531(.A1(new_n13381_), .A2(pi0183), .B(new_n12694_), .ZN(new_n19536_));
  NAND3_X1   g16532(.A1(new_n19536_), .A2(new_n19535_), .A3(new_n15509_), .ZN(new_n19537_));
  NOR2_X1    g16533(.A1(new_n19537_), .A2(new_n19534_), .ZN(new_n19538_));
  NOR2_X1    g16534(.A1(new_n12828_), .A2(pi0183), .ZN(new_n19539_));
  OAI21_X1   g16535(.A1(new_n13367_), .A2(pi0755), .B(pi0038), .ZN(new_n19540_));
  OAI22_X1   g16536(.A1(new_n19538_), .A2(pi0038), .B1(new_n19539_), .B2(new_n19540_), .ZN(new_n19541_));
  NOR2_X1    g16537(.A1(new_n19541_), .A2(new_n3232_), .ZN(new_n19542_));
  AOI21_X1   g16538(.A1(new_n7180_), .A2(new_n3232_), .B(new_n19542_), .ZN(new_n19543_));
  INV_X1     g16539(.I(new_n19543_), .ZN(new_n19544_));
  OAI21_X1   g16540(.A1(new_n19532_), .A2(new_n11924_), .B(new_n11870_), .ZN(new_n19545_));
  AOI21_X1   g16541(.A1(new_n19544_), .A2(new_n11924_), .B(new_n19545_), .ZN(new_n19546_));
  NAND2_X1   g16542(.A1(new_n19543_), .A2(new_n11924_), .ZN(new_n19547_));
  OAI22_X1   g16543(.A1(new_n19547_), .A2(pi0609), .B1(new_n12996_), .B2(new_n19531_), .ZN(new_n19548_));
  NAND2_X1   g16544(.A1(new_n19548_), .A2(new_n11912_), .ZN(new_n19549_));
  OAI22_X1   g16545(.A1(new_n19547_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n19531_), .ZN(new_n19550_));
  NAND2_X1   g16546(.A1(new_n19550_), .A2(pi1155), .ZN(new_n19551_));
  AOI21_X1   g16547(.A1(new_n19549_), .A2(new_n19551_), .B(new_n11870_), .ZN(new_n19552_));
  XOR2_X1    g16548(.A1(new_n19552_), .A2(new_n19546_), .Z(new_n19553_));
  OAI21_X1   g16549(.A1(new_n19532_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n19554_));
  AOI21_X1   g16550(.A1(new_n19553_), .A2(pi0618), .B(new_n19554_), .ZN(new_n19555_));
  NAND2_X1   g16551(.A1(new_n19553_), .A2(pi0618), .ZN(new_n19556_));
  AOI21_X1   g16552(.A1(new_n19532_), .A2(new_n11934_), .B(pi1154), .ZN(new_n19557_));
  NAND2_X1   g16553(.A1(new_n19556_), .A2(new_n19557_), .ZN(new_n19558_));
  NAND2_X1   g16554(.A1(new_n19558_), .A2(new_n19555_), .ZN(new_n19559_));
  MUX2_X1    g16555(.I0(new_n19559_), .I1(new_n19553_), .S(new_n11969_), .Z(new_n19560_));
  NAND2_X1   g16556(.A1(new_n19560_), .A2(new_n11985_), .ZN(new_n19561_));
  NOR3_X1    g16557(.A1(new_n19531_), .A2(pi0619), .A3(pi1159), .ZN(new_n19562_));
  NOR2_X1    g16558(.A1(new_n19562_), .A2(new_n11985_), .ZN(new_n19563_));
  XOR2_X1    g16559(.A1(new_n19561_), .A2(new_n19563_), .Z(new_n19564_));
  OAI21_X1   g16560(.A1(new_n19564_), .A2(new_n11997_), .B(new_n19533_), .ZN(new_n19565_));
  NOR2_X1    g16561(.A1(new_n19531_), .A2(new_n12054_), .ZN(new_n19566_));
  AOI21_X1   g16562(.A1(new_n19565_), .A2(new_n12054_), .B(new_n19566_), .ZN(new_n19567_));
  NAND2_X1   g16563(.A1(new_n19532_), .A2(new_n12091_), .ZN(new_n19568_));
  OAI21_X1   g16564(.A1(new_n19567_), .A2(new_n12091_), .B(new_n19568_), .ZN(new_n19569_));
  AOI21_X1   g16565(.A1(new_n19531_), .A2(pi0644), .B(new_n12099_), .ZN(new_n19570_));
  OAI21_X1   g16566(.A1(new_n19569_), .A2(pi0644), .B(new_n19570_), .ZN(new_n19571_));
  AND2_X2    g16567(.A1(new_n19571_), .A2(new_n12081_), .Z(new_n19572_));
  NOR2_X1    g16568(.A1(new_n19532_), .A2(pi0647), .ZN(new_n19573_));
  NOR2_X1    g16569(.A1(new_n19531_), .A2(new_n13114_), .ZN(new_n19574_));
  NOR2_X1    g16570(.A1(new_n19532_), .A2(new_n12014_), .ZN(new_n19575_));
  NOR2_X1    g16571(.A1(new_n19531_), .A2(new_n11961_), .ZN(new_n19576_));
  OAI21_X1   g16572(.A1(new_n15189_), .A2(new_n19539_), .B(new_n15535_), .ZN(new_n19577_));
  NOR2_X1    g16573(.A1(new_n13395_), .A2(new_n7180_), .ZN(new_n19578_));
  NOR2_X1    g16574(.A1(new_n19578_), .A2(pi0038), .ZN(new_n19579_));
  OAI22_X1   g16575(.A1(new_n19579_), .A2(new_n3232_), .B1(pi0183), .B2(new_n13399_), .ZN(new_n19580_));
  NOR2_X1    g16576(.A1(new_n3232_), .A2(pi0725), .ZN(new_n19581_));
  AOI22_X1   g16577(.A1(new_n19532_), .A2(new_n19581_), .B1(new_n19577_), .B2(new_n19580_), .ZN(new_n19582_));
  NOR3_X1    g16578(.A1(new_n19532_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n19583_));
  NOR4_X1    g16579(.A1(new_n19582_), .A2(new_n12970_), .A3(pi1153), .A4(new_n19531_), .ZN(new_n19584_));
  NOR2_X1    g16580(.A1(new_n19584_), .A2(new_n19583_), .ZN(new_n19585_));
  MUX2_X1    g16581(.I0(new_n19585_), .I1(new_n19582_), .S(new_n11891_), .Z(new_n19586_));
  NOR2_X1    g16582(.A1(new_n19586_), .A2(new_n13024_), .ZN(new_n19587_));
  AOI21_X1   g16583(.A1(new_n13024_), .A2(new_n19531_), .B(new_n19587_), .ZN(new_n19588_));
  AOI21_X1   g16584(.A1(new_n19588_), .A2(new_n11961_), .B(new_n19576_), .ZN(new_n19589_));
  AOI21_X1   g16585(.A1(new_n19589_), .A2(new_n12014_), .B(new_n19575_), .ZN(new_n19590_));
  AOI21_X1   g16586(.A1(new_n19590_), .A2(new_n13114_), .B(new_n19574_), .ZN(new_n19591_));
  INV_X1     g16587(.I(new_n19591_), .ZN(new_n19592_));
  NAND3_X1   g16588(.A1(new_n19531_), .A2(pi0628), .A3(pi1156), .ZN(new_n19593_));
  NOR4_X1    g16589(.A1(new_n19591_), .A2(new_n12031_), .A3(pi1156), .A4(new_n19531_), .ZN(new_n19594_));
  INV_X1     g16590(.I(new_n19594_), .ZN(new_n19595_));
  NAND2_X1   g16591(.A1(new_n19595_), .A2(new_n19593_), .ZN(new_n19596_));
  MUX2_X1    g16592(.I0(new_n19596_), .I1(new_n19592_), .S(new_n11868_), .Z(new_n19597_));
  AOI21_X1   g16593(.A1(new_n19597_), .A2(pi0647), .B(new_n19573_), .ZN(new_n19598_));
  NAND2_X1   g16594(.A1(new_n19598_), .A2(pi1157), .ZN(new_n19599_));
  NOR2_X1    g16595(.A1(new_n19532_), .A2(new_n12061_), .ZN(new_n19600_));
  AOI21_X1   g16596(.A1(new_n19597_), .A2(new_n12061_), .B(new_n19600_), .ZN(new_n19601_));
  NAND2_X1   g16597(.A1(new_n19601_), .A2(new_n12049_), .ZN(new_n19602_));
  NAND2_X1   g16598(.A1(new_n19599_), .A2(new_n19602_), .ZN(new_n19603_));
  NOR2_X1    g16599(.A1(new_n19597_), .A2(pi0787), .ZN(new_n19604_));
  AOI21_X1   g16600(.A1(new_n19603_), .A2(pi0787), .B(new_n19604_), .ZN(new_n19605_));
  AOI21_X1   g16601(.A1(new_n19605_), .A2(pi0644), .B(pi0715), .ZN(new_n19606_));
  NOR2_X1    g16602(.A1(new_n19572_), .A2(new_n19606_), .ZN(new_n19607_));
  NAND3_X1   g16603(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n19608_));
  OR2_X2     g16604(.A1(new_n19569_), .A2(new_n19608_), .Z(new_n19609_));
  NAND2_X1   g16605(.A1(new_n19609_), .A2(pi0715), .ZN(new_n19610_));
  AOI21_X1   g16606(.A1(new_n12082_), .A2(new_n19605_), .B(new_n19610_), .ZN(new_n19611_));
  OAI21_X1   g16607(.A1(new_n19611_), .A2(new_n19607_), .B(pi0790), .ZN(new_n19612_));
  NAND2_X1   g16608(.A1(new_n19560_), .A2(pi0619), .ZN(new_n19613_));
  NAND2_X1   g16609(.A1(new_n19531_), .A2(pi0619), .ZN(new_n19614_));
  NOR3_X1    g16610(.A1(new_n19541_), .A2(new_n15535_), .A3(new_n3231_), .ZN(new_n19624_));
  AOI21_X1   g16611(.A1(pi0183), .A2(new_n3232_), .B(new_n19624_), .ZN(new_n19625_));
  INV_X1     g16612(.I(new_n19584_), .ZN(new_n19626_));
  NAND2_X1   g16613(.A1(new_n19625_), .A2(pi0625), .ZN(new_n19627_));
  NAND2_X1   g16614(.A1(new_n19544_), .A2(pi0625), .ZN(new_n19628_));
  NAND4_X1   g16615(.A1(new_n19628_), .A2(new_n12977_), .A3(new_n19626_), .A4(new_n19627_), .ZN(new_n19629_));
  NAND2_X1   g16616(.A1(new_n19543_), .A2(new_n12970_), .ZN(new_n19630_));
  AND3_X2    g16617(.A1(new_n19627_), .A2(new_n11893_), .A3(new_n19630_), .Z(new_n19631_));
  OAI21_X1   g16618(.A1(new_n19631_), .A2(new_n19583_), .B(new_n13657_), .ZN(new_n19632_));
  AOI21_X1   g16619(.A1(new_n19632_), .A2(new_n19629_), .B(new_n11891_), .ZN(new_n19633_));
  AOI21_X1   g16620(.A1(new_n11891_), .A2(new_n19625_), .B(new_n19633_), .ZN(new_n19634_));
  NOR2_X1    g16621(.A1(new_n19634_), .A2(pi0785), .ZN(new_n19635_));
  INV_X1     g16622(.I(new_n19586_), .ZN(new_n19636_));
  NAND3_X1   g16623(.A1(new_n19636_), .A2(pi0609), .A3(pi1155), .ZN(new_n19637_));
  NAND3_X1   g16624(.A1(new_n19637_), .A2(new_n11923_), .A3(new_n19551_), .ZN(new_n19638_));
  NOR4_X1    g16625(.A1(new_n19634_), .A2(new_n11903_), .A3(pi1155), .A4(new_n19636_), .ZN(new_n19639_));
  NAND2_X1   g16626(.A1(new_n19549_), .A2(pi0660), .ZN(new_n19640_));
  NOR2_X1    g16627(.A1(new_n19639_), .A2(new_n19640_), .ZN(new_n19641_));
  NOR2_X1    g16628(.A1(new_n19641_), .A2(new_n11870_), .ZN(new_n19642_));
  AOI21_X1   g16629(.A1(new_n19642_), .A2(new_n19638_), .B(new_n19635_), .ZN(new_n19643_));
  INV_X1     g16630(.I(new_n19588_), .ZN(new_n19644_));
  NOR4_X1    g16631(.A1(new_n19643_), .A2(new_n11934_), .A3(pi1154), .A4(new_n19644_), .ZN(new_n19645_));
  NAND2_X1   g16632(.A1(new_n19555_), .A2(pi0627), .ZN(new_n19646_));
  NOR3_X1    g16633(.A1(new_n19588_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n19647_));
  NAND2_X1   g16634(.A1(new_n19558_), .A2(new_n11949_), .ZN(new_n19648_));
  OAI22_X1   g16635(.A1(new_n19645_), .A2(new_n19646_), .B1(new_n19647_), .B2(new_n19648_), .ZN(new_n19649_));
  MUX2_X1    g16636(.I0(new_n19649_), .I1(new_n19643_), .S(new_n11969_), .Z(new_n19650_));
  XNOR2_X1   g16637(.A1(new_n19650_), .A2(new_n19589_), .ZN(new_n19651_));
  NOR2_X1    g16638(.A1(new_n19651_), .A2(new_n11967_), .ZN(new_n19652_));
  NAND3_X1   g16639(.A1(new_n19613_), .A2(new_n11869_), .A3(new_n19614_), .ZN(new_n19653_));
  XNOR2_X1   g16640(.A1(new_n19652_), .A2(new_n19650_), .ZN(new_n19654_));
  NAND2_X1   g16641(.A1(new_n19654_), .A2(new_n11869_), .ZN(new_n19655_));
  AOI21_X1   g16642(.A1(new_n19532_), .A2(new_n11967_), .B(pi1159), .ZN(new_n19656_));
  AOI21_X1   g16643(.A1(new_n19613_), .A2(new_n19656_), .B(pi0648), .ZN(new_n19657_));
  INV_X1     g16644(.I(new_n19564_), .ZN(new_n19658_));
  MUX2_X1    g16645(.I0(new_n19658_), .I1(new_n19532_), .S(new_n11994_), .Z(new_n19659_));
  AOI21_X1   g16646(.A1(new_n19564_), .A2(new_n19532_), .B(new_n11994_), .ZN(new_n19660_));
  OAI21_X1   g16647(.A1(new_n19590_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n19661_));
  AOI21_X1   g16648(.A1(new_n19660_), .A2(new_n11990_), .B(new_n19661_), .ZN(new_n19662_));
  OAI21_X1   g16649(.A1(new_n19659_), .A2(new_n17167_), .B(new_n19662_), .ZN(new_n19663_));
  OAI21_X1   g16650(.A1(new_n19650_), .A2(pi0789), .B(new_n11998_), .ZN(new_n19664_));
  NAND3_X1   g16651(.A1(new_n19663_), .A2(new_n17372_), .A3(new_n19664_), .ZN(new_n19665_));
  AOI21_X1   g16652(.A1(new_n19655_), .A2(new_n19657_), .B(new_n19665_), .ZN(new_n19666_));
  NAND2_X1   g16653(.A1(new_n19593_), .A2(pi0629), .ZN(new_n19667_));
  OAI21_X1   g16654(.A1(new_n19594_), .A2(pi0629), .B(new_n19667_), .ZN(new_n19668_));
  NAND2_X1   g16655(.A1(new_n19565_), .A2(new_n15222_), .ZN(new_n19669_));
  NAND2_X1   g16656(.A1(new_n19669_), .A2(new_n19668_), .ZN(new_n19670_));
  AOI22_X1   g16657(.A1(new_n19666_), .A2(new_n19653_), .B1(pi0792), .B2(new_n19670_), .ZN(new_n19671_));
  NAND2_X1   g16658(.A1(new_n19598_), .A2(new_n12060_), .ZN(new_n19672_));
  AOI21_X1   g16659(.A1(new_n19601_), .A2(pi0630), .B(new_n15214_), .ZN(new_n19673_));
  NAND2_X1   g16660(.A1(new_n19673_), .A2(new_n19672_), .ZN(new_n19674_));
  NOR2_X1    g16661(.A1(new_n19567_), .A2(new_n15183_), .ZN(new_n19675_));
  NAND2_X1   g16662(.A1(new_n19572_), .A2(new_n12082_), .ZN(new_n19676_));
  AOI21_X1   g16663(.A1(new_n19609_), .A2(pi0644), .B(pi0790), .ZN(new_n19677_));
  AOI22_X1   g16664(.A1(new_n19676_), .A2(new_n19677_), .B1(new_n19674_), .B2(new_n19675_), .ZN(new_n19678_));
  OAI21_X1   g16665(.A1(new_n19671_), .A2(new_n14725_), .B(new_n19678_), .ZN(new_n19679_));
  AOI21_X1   g16666(.A1(new_n19679_), .A2(new_n19612_), .B(po1038), .ZN(new_n19680_));
  OAI21_X1   g16667(.A1(new_n6845_), .A2(pi0183), .B(new_n13184_), .ZN(new_n19681_));
  OAI21_X1   g16668(.A1(new_n19680_), .A2(new_n19681_), .B(new_n19530_), .ZN(po0340));
  NOR2_X1    g16669(.A1(new_n2925_), .A2(pi0184), .ZN(new_n19683_));
  NOR2_X1    g16670(.A1(new_n11877_), .A2(pi0777), .ZN(new_n19684_));
  NOR2_X1    g16671(.A1(new_n19684_), .A2(new_n19683_), .ZN(new_n19685_));
  AOI21_X1   g16672(.A1(new_n11886_), .A2(new_n16072_), .B(new_n19683_), .ZN(new_n19686_));
  NOR2_X1    g16673(.A1(new_n19686_), .A2(new_n11874_), .ZN(new_n19687_));
  INV_X1     g16674(.I(new_n19687_), .ZN(new_n19688_));
  NAND2_X1   g16675(.A1(new_n19688_), .A2(new_n19685_), .ZN(new_n19689_));
  NAND2_X1   g16676(.A1(new_n19689_), .A2(new_n11891_), .ZN(new_n19690_));
  NOR2_X1    g16677(.A1(new_n19688_), .A2(new_n12970_), .ZN(new_n19691_));
  NOR4_X1    g16678(.A1(new_n19691_), .A2(new_n11893_), .A3(new_n19683_), .A4(new_n19684_), .ZN(new_n19692_));
  NOR3_X1    g16679(.A1(new_n11894_), .A2(pi0625), .A3(pi0737), .ZN(new_n19693_));
  NOR2_X1    g16680(.A1(new_n19683_), .A2(pi1153), .ZN(new_n19694_));
  INV_X1     g16681(.I(new_n19694_), .ZN(new_n19695_));
  NOR2_X1    g16682(.A1(new_n19693_), .A2(new_n19695_), .ZN(new_n19696_));
  INV_X1     g16683(.I(new_n19696_), .ZN(new_n19697_));
  NAND2_X1   g16684(.A1(new_n19697_), .A2(pi0608), .ZN(new_n19698_));
  INV_X1     g16685(.I(new_n19691_), .ZN(new_n19699_));
  AOI21_X1   g16686(.A1(new_n19699_), .A2(new_n19689_), .B(new_n19695_), .ZN(new_n19700_));
  OAI21_X1   g16687(.A1(new_n19693_), .A2(new_n19686_), .B(pi1153), .ZN(new_n19701_));
  NAND2_X1   g16688(.A1(new_n19701_), .A2(new_n13657_), .ZN(new_n19702_));
  OAI22_X1   g16689(.A1(new_n19700_), .A2(new_n19702_), .B1(new_n19692_), .B2(new_n19698_), .ZN(new_n19703_));
  NAND2_X1   g16690(.A1(new_n19703_), .A2(pi0778), .ZN(new_n19704_));
  XOR2_X1    g16691(.A1(new_n19704_), .A2(new_n19690_), .Z(new_n19705_));
  INV_X1     g16692(.I(new_n19705_), .ZN(new_n19706_));
  NAND2_X1   g16693(.A1(new_n19697_), .A2(new_n19701_), .ZN(new_n19707_));
  MUX2_X1    g16694(.I0(new_n19707_), .I1(new_n19686_), .S(new_n11891_), .Z(new_n19708_));
  XNOR2_X1   g16695(.A1(new_n19705_), .A2(new_n19708_), .ZN(new_n19709_));
  NAND2_X1   g16696(.A1(new_n19709_), .A2(pi0609), .ZN(new_n19710_));
  XOR2_X1    g16697(.A1(new_n19710_), .A2(new_n19705_), .Z(new_n19711_));
  NAND2_X1   g16698(.A1(new_n19711_), .A2(new_n11912_), .ZN(new_n19712_));
  NOR2_X1    g16699(.A1(new_n19685_), .A2(new_n11925_), .ZN(new_n19713_));
  INV_X1     g16700(.I(new_n19713_), .ZN(new_n19714_));
  NOR3_X1    g16701(.A1(new_n12997_), .A2(new_n11877_), .A3(pi0777), .ZN(new_n19715_));
  NAND3_X1   g16702(.A1(new_n19714_), .A2(new_n11912_), .A3(new_n19715_), .ZN(new_n19716_));
  NAND3_X1   g16703(.A1(new_n19712_), .A2(new_n11923_), .A3(new_n19716_), .ZN(new_n19717_));
  NOR4_X1    g16704(.A1(new_n19715_), .A2(new_n11923_), .A3(pi1155), .A4(new_n19683_), .ZN(new_n19719_));
  NOR2_X1    g16705(.A1(new_n19719_), .A2(new_n11870_), .ZN(new_n19720_));
  AOI22_X1   g16706(.A1(new_n19717_), .A2(new_n19720_), .B1(new_n11870_), .B2(new_n19706_), .ZN(new_n19721_));
  NOR2_X1    g16707(.A1(new_n19721_), .A2(pi0781), .ZN(new_n19722_));
  NOR4_X1    g16708(.A1(new_n19708_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n19723_));
  NOR3_X1    g16709(.A1(new_n19715_), .A2(pi1155), .A3(new_n19683_), .ZN(new_n19724_));
  NAND2_X1   g16710(.A1(new_n19716_), .A2(new_n19724_), .ZN(new_n19725_));
  MUX2_X1    g16711(.I0(new_n19725_), .I1(new_n19714_), .S(new_n11870_), .Z(new_n19726_));
  INV_X1     g16712(.I(new_n19726_), .ZN(new_n19727_));
  OAI21_X1   g16713(.A1(new_n19727_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n19728_));
  OAI21_X1   g16714(.A1(new_n19727_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n19729_));
  NOR2_X1    g16715(.A1(new_n19708_), .A2(new_n11939_), .ZN(new_n19730_));
  NOR4_X1    g16716(.A1(new_n19721_), .A2(new_n11934_), .A3(pi1154), .A4(new_n19730_), .ZN(new_n19731_));
  NOR2_X1    g16717(.A1(new_n19731_), .A2(new_n19729_), .ZN(new_n19732_));
  OAI22_X1   g16718(.A1(new_n19732_), .A2(pi0627), .B1(new_n19723_), .B2(new_n19728_), .ZN(new_n19733_));
  AOI21_X1   g16719(.A1(new_n19733_), .A2(pi0781), .B(new_n19722_), .ZN(new_n19734_));
  INV_X1     g16720(.I(new_n19730_), .ZN(new_n19735_));
  NOR2_X1    g16721(.A1(new_n19735_), .A2(new_n11962_), .ZN(new_n19736_));
  NOR4_X1    g16722(.A1(new_n19734_), .A2(new_n11967_), .A3(pi1159), .A4(new_n19736_), .ZN(new_n19737_));
  NOR2_X1    g16723(.A1(new_n19727_), .A2(pi0781), .ZN(new_n19738_));
  AOI21_X1   g16724(.A1(new_n11944_), .A2(new_n19726_), .B(new_n19729_), .ZN(new_n19739_));
  NOR2_X1    g16725(.A1(new_n19739_), .A2(new_n11969_), .ZN(new_n19740_));
  XOR2_X1    g16726(.A1(new_n19740_), .A2(new_n19738_), .Z(new_n19741_));
  AOI21_X1   g16727(.A1(new_n19741_), .A2(new_n16479_), .B(pi1159), .ZN(new_n19742_));
  INV_X1     g16728(.I(new_n19742_), .ZN(new_n19743_));
  NOR3_X1    g16729(.A1(new_n19737_), .A2(new_n11966_), .A3(new_n19743_), .ZN(new_n19744_));
  NOR4_X1    g16730(.A1(new_n19735_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n19745_));
  INV_X1     g16731(.I(new_n19741_), .ZN(new_n19746_));
  NOR2_X1    g16732(.A1(new_n19746_), .A2(new_n16482_), .ZN(new_n19747_));
  NOR3_X1    g16733(.A1(new_n19747_), .A2(pi0648), .A3(new_n19745_), .ZN(new_n19748_));
  AOI21_X1   g16734(.A1(new_n19734_), .A2(new_n11998_), .B(pi0789), .ZN(new_n19749_));
  OAI21_X1   g16735(.A1(new_n19744_), .A2(new_n19748_), .B(new_n19749_), .ZN(new_n19750_));
  NAND2_X1   g16736(.A1(new_n19736_), .A2(new_n17450_), .ZN(new_n19751_));
  NOR2_X1    g16737(.A1(new_n19751_), .A2(new_n17153_), .ZN(new_n19752_));
  NOR2_X1    g16738(.A1(new_n14624_), .A2(new_n19683_), .ZN(new_n19753_));
  NOR2_X1    g16739(.A1(new_n19746_), .A2(pi0789), .ZN(new_n19754_));
  NOR2_X1    g16740(.A1(new_n19743_), .A2(new_n19747_), .ZN(new_n19755_));
  NOR2_X1    g16741(.A1(new_n19755_), .A2(new_n11985_), .ZN(new_n19756_));
  XOR2_X1    g16742(.A1(new_n19756_), .A2(new_n19754_), .Z(new_n19757_));
  AOI21_X1   g16743(.A1(new_n19757_), .A2(new_n14624_), .B(new_n19753_), .ZN(new_n19758_));
  AOI22_X1   g16744(.A1(new_n19758_), .A2(new_n12064_), .B1(new_n15080_), .B2(new_n19752_), .ZN(new_n19759_));
  NOR2_X1    g16745(.A1(new_n19759_), .A2(new_n12030_), .ZN(new_n19760_));
  NAND2_X1   g16746(.A1(new_n19758_), .A2(new_n12063_), .ZN(new_n19761_));
  AOI21_X1   g16747(.A1(new_n19752_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n19762_));
  NAND2_X1   g16748(.A1(new_n19761_), .A2(new_n19762_), .ZN(new_n19763_));
  OAI21_X1   g16749(.A1(new_n19760_), .A2(new_n19763_), .B(new_n14726_), .ZN(new_n19764_));
  INV_X1     g16750(.I(new_n19683_), .ZN(new_n19765_));
  MUX2_X1    g16751(.I0(new_n19757_), .I1(new_n19765_), .S(new_n11994_), .Z(new_n19766_));
  INV_X1     g16752(.I(new_n19757_), .ZN(new_n19767_));
  AOI21_X1   g16753(.A1(new_n19767_), .A2(new_n19765_), .B(new_n11994_), .ZN(new_n19768_));
  OAI21_X1   g16754(.A1(new_n19751_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n19769_));
  AOI21_X1   g16755(.A1(new_n19768_), .A2(new_n11990_), .B(new_n19769_), .ZN(new_n19770_));
  OAI21_X1   g16756(.A1(new_n17167_), .A2(new_n19766_), .B(new_n19770_), .ZN(new_n19771_));
  NAND4_X1   g16757(.A1(new_n19750_), .A2(new_n14732_), .A3(new_n19764_), .A4(new_n19771_), .ZN(new_n19772_));
  NAND3_X1   g16758(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n19683_), .ZN(new_n19773_));
  NAND2_X1   g16759(.A1(new_n19752_), .A2(new_n15050_), .ZN(new_n19774_));
  NAND2_X1   g16760(.A1(new_n19774_), .A2(pi0647), .ZN(new_n19775_));
  NAND2_X1   g16761(.A1(new_n19683_), .A2(pi0647), .ZN(new_n19776_));
  NAND3_X1   g16762(.A1(new_n19775_), .A2(new_n12049_), .A3(new_n19776_), .ZN(new_n19777_));
  NAND2_X1   g16763(.A1(new_n19777_), .A2(pi0630), .ZN(new_n19778_));
  NOR2_X1    g16764(.A1(new_n19774_), .A2(new_n12061_), .ZN(new_n19779_));
  AOI21_X1   g16765(.A1(new_n12061_), .A2(new_n19683_), .B(new_n19779_), .ZN(new_n19780_));
  NAND2_X1   g16766(.A1(new_n19780_), .A2(new_n12088_), .ZN(new_n19781_));
  NAND4_X1   g16767(.A1(new_n19781_), .A2(new_n19778_), .A3(pi0787), .A4(new_n19773_), .ZN(new_n19782_));
  AND2_X2    g16768(.A1(new_n19772_), .A2(new_n19782_), .Z(new_n19783_));
  NOR2_X1    g16769(.A1(new_n19783_), .A2(new_n12082_), .ZN(new_n19784_));
  NAND4_X1   g16770(.A1(new_n19775_), .A2(pi0787), .A3(new_n12049_), .A4(new_n19776_), .ZN(new_n19785_));
  OAI21_X1   g16771(.A1(pi0787), .A2(new_n19774_), .B(new_n19785_), .ZN(new_n19786_));
  NOR2_X1    g16772(.A1(new_n19786_), .A2(pi0644), .ZN(new_n19787_));
  OR3_X2     g16773(.A1(new_n19784_), .A2(pi0715), .A3(new_n19787_), .Z(new_n19788_));
  MUX2_X1    g16774(.I0(new_n19758_), .I1(new_n19683_), .S(new_n16841_), .Z(new_n19789_));
  INV_X1     g16775(.I(new_n19789_), .ZN(new_n19790_));
  OAI21_X1   g16776(.A1(new_n19789_), .A2(new_n19683_), .B(new_n12082_), .ZN(new_n19791_));
  AOI21_X1   g16777(.A1(new_n19683_), .A2(new_n19789_), .B(new_n19791_), .ZN(new_n19792_));
  OAI21_X1   g16778(.A1(new_n19792_), .A2(new_n19790_), .B(new_n12099_), .ZN(new_n19793_));
  AOI21_X1   g16779(.A1(new_n19790_), .A2(new_n19792_), .B(new_n19793_), .ZN(new_n19794_));
  AOI21_X1   g16780(.A1(new_n19788_), .A2(new_n19794_), .B(pi1160), .ZN(new_n19795_));
  XOR2_X1    g16781(.A1(new_n19792_), .A2(new_n19683_), .Z(new_n19796_));
  AOI21_X1   g16782(.A1(new_n19786_), .A2(pi0644), .B(new_n13169_), .ZN(new_n19797_));
  OAI21_X1   g16783(.A1(new_n19796_), .A2(new_n12099_), .B(new_n19797_), .ZN(new_n19798_));
  OAI21_X1   g16784(.A1(new_n19784_), .A2(new_n19798_), .B(pi0790), .ZN(new_n19799_));
  NOR2_X1    g16785(.A1(new_n19783_), .A2(new_n14748_), .ZN(new_n19800_));
  OAI21_X1   g16786(.A1(new_n19795_), .A2(new_n19799_), .B(new_n19800_), .ZN(new_n19801_));
  NOR2_X1    g16787(.A1(new_n12965_), .A2(pi0184), .ZN(new_n19802_));
  INV_X1     g16788(.I(new_n19802_), .ZN(new_n19803_));
  NAND2_X1   g16789(.A1(new_n19803_), .A2(new_n11997_), .ZN(new_n19804_));
  AOI21_X1   g16790(.A1(new_n12794_), .A2(new_n8883_), .B(pi0777), .ZN(new_n19805_));
  NAND3_X1   g16791(.A1(new_n13381_), .A2(new_n8883_), .A3(new_n14362_), .ZN(new_n19806_));
  OAI21_X1   g16792(.A1(new_n13381_), .A2(pi0184), .B(new_n12694_), .ZN(new_n19807_));
  NAND3_X1   g16793(.A1(new_n19807_), .A2(new_n19806_), .A3(new_n16049_), .ZN(new_n19808_));
  NOR2_X1    g16794(.A1(new_n19808_), .A2(new_n19805_), .ZN(new_n19809_));
  NOR2_X1    g16795(.A1(new_n12828_), .A2(pi0184), .ZN(new_n19810_));
  OAI21_X1   g16796(.A1(new_n13367_), .A2(pi0777), .B(pi0038), .ZN(new_n19811_));
  OAI22_X1   g16797(.A1(new_n19809_), .A2(pi0038), .B1(new_n19810_), .B2(new_n19811_), .ZN(new_n19812_));
  NOR2_X1    g16798(.A1(new_n19812_), .A2(new_n3232_), .ZN(new_n19813_));
  AOI21_X1   g16799(.A1(new_n8883_), .A2(new_n3232_), .B(new_n19813_), .ZN(new_n19814_));
  INV_X1     g16800(.I(new_n19814_), .ZN(new_n19815_));
  OAI21_X1   g16801(.A1(new_n19803_), .A2(new_n11924_), .B(new_n11870_), .ZN(new_n19816_));
  AOI21_X1   g16802(.A1(new_n19815_), .A2(new_n11924_), .B(new_n19816_), .ZN(new_n19817_));
  NAND2_X1   g16803(.A1(new_n19814_), .A2(new_n11924_), .ZN(new_n19818_));
  OAI22_X1   g16804(.A1(new_n19818_), .A2(pi0609), .B1(new_n12996_), .B2(new_n19802_), .ZN(new_n19819_));
  NAND2_X1   g16805(.A1(new_n19819_), .A2(new_n11912_), .ZN(new_n19820_));
  OAI22_X1   g16806(.A1(new_n19818_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n19802_), .ZN(new_n19821_));
  NAND2_X1   g16807(.A1(new_n19821_), .A2(pi1155), .ZN(new_n19822_));
  AOI21_X1   g16808(.A1(new_n19820_), .A2(new_n19822_), .B(new_n11870_), .ZN(new_n19823_));
  XOR2_X1    g16809(.A1(new_n19823_), .A2(new_n19817_), .Z(new_n19824_));
  OAI21_X1   g16810(.A1(new_n19803_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n19825_));
  AOI21_X1   g16811(.A1(new_n19824_), .A2(pi0618), .B(new_n19825_), .ZN(new_n19826_));
  NAND2_X1   g16812(.A1(new_n19824_), .A2(pi0618), .ZN(new_n19827_));
  AOI21_X1   g16813(.A1(new_n19803_), .A2(new_n11934_), .B(pi1154), .ZN(new_n19828_));
  NAND2_X1   g16814(.A1(new_n19827_), .A2(new_n19828_), .ZN(new_n19829_));
  NAND2_X1   g16815(.A1(new_n19829_), .A2(new_n19826_), .ZN(new_n19830_));
  MUX2_X1    g16816(.I0(new_n19830_), .I1(new_n19824_), .S(new_n11969_), .Z(new_n19831_));
  NAND2_X1   g16817(.A1(new_n19831_), .A2(new_n11985_), .ZN(new_n19832_));
  NOR3_X1    g16818(.A1(new_n19802_), .A2(pi0619), .A3(pi1159), .ZN(new_n19833_));
  NOR2_X1    g16819(.A1(new_n19833_), .A2(new_n11985_), .ZN(new_n19834_));
  XOR2_X1    g16820(.A1(new_n19832_), .A2(new_n19834_), .Z(new_n19835_));
  OAI21_X1   g16821(.A1(new_n19835_), .A2(new_n11997_), .B(new_n19804_), .ZN(new_n19836_));
  NOR2_X1    g16822(.A1(new_n19802_), .A2(new_n12054_), .ZN(new_n19837_));
  AOI21_X1   g16823(.A1(new_n19836_), .A2(new_n12054_), .B(new_n19837_), .ZN(new_n19838_));
  NAND2_X1   g16824(.A1(new_n19803_), .A2(new_n12091_), .ZN(new_n19839_));
  OAI21_X1   g16825(.A1(new_n19838_), .A2(new_n12091_), .B(new_n19839_), .ZN(new_n19840_));
  AOI21_X1   g16826(.A1(new_n19802_), .A2(pi0644), .B(new_n12099_), .ZN(new_n19841_));
  OAI21_X1   g16827(.A1(new_n19840_), .A2(pi0644), .B(new_n19841_), .ZN(new_n19842_));
  AND2_X2    g16828(.A1(new_n19842_), .A2(new_n12081_), .Z(new_n19843_));
  NOR2_X1    g16829(.A1(new_n19803_), .A2(pi0647), .ZN(new_n19844_));
  NOR2_X1    g16830(.A1(new_n19802_), .A2(new_n13114_), .ZN(new_n19845_));
  NOR2_X1    g16831(.A1(new_n19803_), .A2(new_n12014_), .ZN(new_n19846_));
  NOR2_X1    g16832(.A1(new_n19802_), .A2(new_n11961_), .ZN(new_n19847_));
  OAI21_X1   g16833(.A1(new_n15189_), .A2(new_n19810_), .B(new_n16072_), .ZN(new_n19848_));
  NOR2_X1    g16834(.A1(new_n13395_), .A2(new_n8883_), .ZN(new_n19849_));
  NOR2_X1    g16835(.A1(new_n19849_), .A2(pi0038), .ZN(new_n19850_));
  OAI22_X1   g16836(.A1(new_n19850_), .A2(new_n3232_), .B1(pi0184), .B2(new_n13399_), .ZN(new_n19851_));
  NOR2_X1    g16837(.A1(new_n3232_), .A2(pi0737), .ZN(new_n19852_));
  AOI22_X1   g16838(.A1(new_n19803_), .A2(new_n19852_), .B1(new_n19848_), .B2(new_n19851_), .ZN(new_n19853_));
  NOR3_X1    g16839(.A1(new_n19803_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n19854_));
  NOR4_X1    g16840(.A1(new_n19853_), .A2(new_n12970_), .A3(pi1153), .A4(new_n19802_), .ZN(new_n19855_));
  NOR2_X1    g16841(.A1(new_n19855_), .A2(new_n19854_), .ZN(new_n19856_));
  MUX2_X1    g16842(.I0(new_n19856_), .I1(new_n19853_), .S(new_n11891_), .Z(new_n19857_));
  NOR2_X1    g16843(.A1(new_n19857_), .A2(new_n13024_), .ZN(new_n19858_));
  AOI21_X1   g16844(.A1(new_n13024_), .A2(new_n19802_), .B(new_n19858_), .ZN(new_n19859_));
  AOI21_X1   g16845(.A1(new_n19859_), .A2(new_n11961_), .B(new_n19847_), .ZN(new_n19860_));
  AOI21_X1   g16846(.A1(new_n19860_), .A2(new_n12014_), .B(new_n19846_), .ZN(new_n19861_));
  AOI21_X1   g16847(.A1(new_n19861_), .A2(new_n13114_), .B(new_n19845_), .ZN(new_n19862_));
  INV_X1     g16848(.I(new_n19862_), .ZN(new_n19863_));
  NAND3_X1   g16849(.A1(new_n19802_), .A2(pi0628), .A3(pi1156), .ZN(new_n19864_));
  NOR4_X1    g16850(.A1(new_n19862_), .A2(new_n12031_), .A3(pi1156), .A4(new_n19802_), .ZN(new_n19865_));
  INV_X1     g16851(.I(new_n19865_), .ZN(new_n19866_));
  NAND2_X1   g16852(.A1(new_n19866_), .A2(new_n19864_), .ZN(new_n19867_));
  MUX2_X1    g16853(.I0(new_n19867_), .I1(new_n19863_), .S(new_n11868_), .Z(new_n19868_));
  AOI21_X1   g16854(.A1(new_n19868_), .A2(pi0647), .B(new_n19844_), .ZN(new_n19869_));
  NAND2_X1   g16855(.A1(new_n19869_), .A2(pi1157), .ZN(new_n19870_));
  NOR2_X1    g16856(.A1(new_n19803_), .A2(new_n12061_), .ZN(new_n19871_));
  AOI21_X1   g16857(.A1(new_n19868_), .A2(new_n12061_), .B(new_n19871_), .ZN(new_n19872_));
  NAND2_X1   g16858(.A1(new_n19872_), .A2(new_n12049_), .ZN(new_n19873_));
  NAND2_X1   g16859(.A1(new_n19870_), .A2(new_n19873_), .ZN(new_n19874_));
  NOR2_X1    g16860(.A1(new_n19868_), .A2(pi0787), .ZN(new_n19875_));
  AOI21_X1   g16861(.A1(new_n19874_), .A2(pi0787), .B(new_n19875_), .ZN(new_n19876_));
  AOI21_X1   g16862(.A1(new_n19876_), .A2(pi0644), .B(pi0715), .ZN(new_n19877_));
  NOR2_X1    g16863(.A1(new_n19843_), .A2(new_n19877_), .ZN(new_n19878_));
  NAND3_X1   g16864(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n19879_));
  OR2_X2     g16865(.A1(new_n19840_), .A2(new_n19879_), .Z(new_n19880_));
  NAND2_X1   g16866(.A1(new_n19880_), .A2(pi0715), .ZN(new_n19881_));
  AOI21_X1   g16867(.A1(new_n12082_), .A2(new_n19876_), .B(new_n19881_), .ZN(new_n19882_));
  OAI21_X1   g16868(.A1(new_n19882_), .A2(new_n19878_), .B(pi0790), .ZN(new_n19883_));
  NAND2_X1   g16869(.A1(new_n19831_), .A2(pi0619), .ZN(new_n19884_));
  NAND2_X1   g16870(.A1(new_n19802_), .A2(pi0619), .ZN(new_n19885_));
  NOR3_X1    g16871(.A1(new_n19812_), .A2(new_n16072_), .A3(new_n3231_), .ZN(new_n19895_));
  AOI21_X1   g16872(.A1(pi0184), .A2(new_n3232_), .B(new_n19895_), .ZN(new_n19896_));
  INV_X1     g16873(.I(new_n19855_), .ZN(new_n19897_));
  NAND2_X1   g16874(.A1(new_n19896_), .A2(pi0625), .ZN(new_n19898_));
  NAND2_X1   g16875(.A1(new_n19815_), .A2(pi0625), .ZN(new_n19899_));
  NAND4_X1   g16876(.A1(new_n19899_), .A2(new_n12977_), .A3(new_n19897_), .A4(new_n19898_), .ZN(new_n19900_));
  NAND2_X1   g16877(.A1(new_n19814_), .A2(new_n12970_), .ZN(new_n19901_));
  AND3_X2    g16878(.A1(new_n19898_), .A2(new_n11893_), .A3(new_n19901_), .Z(new_n19902_));
  OAI21_X1   g16879(.A1(new_n19902_), .A2(new_n19854_), .B(new_n13657_), .ZN(new_n19903_));
  AOI21_X1   g16880(.A1(new_n19903_), .A2(new_n19900_), .B(new_n11891_), .ZN(new_n19904_));
  AOI21_X1   g16881(.A1(new_n11891_), .A2(new_n19896_), .B(new_n19904_), .ZN(new_n19905_));
  NOR2_X1    g16882(.A1(new_n19905_), .A2(pi0785), .ZN(new_n19906_));
  INV_X1     g16883(.I(new_n19857_), .ZN(new_n19907_));
  NAND3_X1   g16884(.A1(new_n19907_), .A2(pi0609), .A3(pi1155), .ZN(new_n19908_));
  NAND3_X1   g16885(.A1(new_n19908_), .A2(new_n11923_), .A3(new_n19822_), .ZN(new_n19909_));
  NOR4_X1    g16886(.A1(new_n19905_), .A2(new_n11903_), .A3(pi1155), .A4(new_n19907_), .ZN(new_n19910_));
  NAND2_X1   g16887(.A1(new_n19820_), .A2(pi0660), .ZN(new_n19911_));
  NOR2_X1    g16888(.A1(new_n19910_), .A2(new_n19911_), .ZN(new_n19912_));
  NOR2_X1    g16889(.A1(new_n19912_), .A2(new_n11870_), .ZN(new_n19913_));
  AOI21_X1   g16890(.A1(new_n19913_), .A2(new_n19909_), .B(new_n19906_), .ZN(new_n19914_));
  INV_X1     g16891(.I(new_n19859_), .ZN(new_n19915_));
  NOR4_X1    g16892(.A1(new_n19914_), .A2(new_n11934_), .A3(pi1154), .A4(new_n19915_), .ZN(new_n19916_));
  NAND2_X1   g16893(.A1(new_n19826_), .A2(pi0627), .ZN(new_n19917_));
  NOR3_X1    g16894(.A1(new_n19859_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n19918_));
  NAND2_X1   g16895(.A1(new_n19829_), .A2(new_n11949_), .ZN(new_n19919_));
  OAI22_X1   g16896(.A1(new_n19916_), .A2(new_n19917_), .B1(new_n19918_), .B2(new_n19919_), .ZN(new_n19920_));
  MUX2_X1    g16897(.I0(new_n19920_), .I1(new_n19914_), .S(new_n11969_), .Z(new_n19921_));
  XNOR2_X1   g16898(.A1(new_n19921_), .A2(new_n19860_), .ZN(new_n19922_));
  NOR2_X1    g16899(.A1(new_n19922_), .A2(new_n11967_), .ZN(new_n19923_));
  NAND3_X1   g16900(.A1(new_n19884_), .A2(new_n11869_), .A3(new_n19885_), .ZN(new_n19924_));
  XNOR2_X1   g16901(.A1(new_n19923_), .A2(new_n19921_), .ZN(new_n19925_));
  NAND2_X1   g16902(.A1(new_n19925_), .A2(new_n11869_), .ZN(new_n19926_));
  AOI21_X1   g16903(.A1(new_n19803_), .A2(new_n11967_), .B(pi1159), .ZN(new_n19927_));
  AOI21_X1   g16904(.A1(new_n19884_), .A2(new_n19927_), .B(pi0648), .ZN(new_n19928_));
  INV_X1     g16905(.I(new_n19835_), .ZN(new_n19929_));
  MUX2_X1    g16906(.I0(new_n19929_), .I1(new_n19803_), .S(new_n11994_), .Z(new_n19930_));
  AOI21_X1   g16907(.A1(new_n19835_), .A2(new_n19803_), .B(new_n11994_), .ZN(new_n19931_));
  OAI21_X1   g16908(.A1(new_n19861_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n19932_));
  AOI21_X1   g16909(.A1(new_n19931_), .A2(new_n11990_), .B(new_n19932_), .ZN(new_n19933_));
  OAI21_X1   g16910(.A1(new_n19930_), .A2(new_n17167_), .B(new_n19933_), .ZN(new_n19934_));
  OAI21_X1   g16911(.A1(new_n19921_), .A2(pi0789), .B(new_n11998_), .ZN(new_n19935_));
  NAND3_X1   g16912(.A1(new_n19934_), .A2(new_n17372_), .A3(new_n19935_), .ZN(new_n19936_));
  AOI21_X1   g16913(.A1(new_n19926_), .A2(new_n19928_), .B(new_n19936_), .ZN(new_n19937_));
  NAND2_X1   g16914(.A1(new_n19864_), .A2(pi0629), .ZN(new_n19938_));
  OAI21_X1   g16915(.A1(new_n19865_), .A2(pi0629), .B(new_n19938_), .ZN(new_n19939_));
  NAND2_X1   g16916(.A1(new_n19836_), .A2(new_n15222_), .ZN(new_n19940_));
  NAND2_X1   g16917(.A1(new_n19940_), .A2(new_n19939_), .ZN(new_n19941_));
  AOI22_X1   g16918(.A1(new_n19937_), .A2(new_n19924_), .B1(pi0792), .B2(new_n19941_), .ZN(new_n19942_));
  NAND2_X1   g16919(.A1(new_n19869_), .A2(new_n12060_), .ZN(new_n19943_));
  AOI21_X1   g16920(.A1(new_n19872_), .A2(pi0630), .B(new_n15214_), .ZN(new_n19944_));
  NAND2_X1   g16921(.A1(new_n19944_), .A2(new_n19943_), .ZN(new_n19945_));
  NOR2_X1    g16922(.A1(new_n19838_), .A2(new_n15183_), .ZN(new_n19946_));
  NAND2_X1   g16923(.A1(new_n19843_), .A2(new_n12082_), .ZN(new_n19947_));
  AOI21_X1   g16924(.A1(new_n19880_), .A2(pi0644), .B(pi0790), .ZN(new_n19948_));
  AOI22_X1   g16925(.A1(new_n19947_), .A2(new_n19948_), .B1(new_n19945_), .B2(new_n19946_), .ZN(new_n19949_));
  OAI21_X1   g16926(.A1(new_n19942_), .A2(new_n14725_), .B(new_n19949_), .ZN(new_n19950_));
  AOI21_X1   g16927(.A1(new_n19950_), .A2(new_n19883_), .B(po1038), .ZN(new_n19951_));
  OAI21_X1   g16928(.A1(new_n6845_), .A2(pi0184), .B(new_n13184_), .ZN(new_n19952_));
  OAI21_X1   g16929(.A1(new_n19951_), .A2(new_n19952_), .B(new_n19801_), .ZN(po0341));
  NOR2_X1    g16930(.A1(new_n2925_), .A2(pi0185), .ZN(new_n19954_));
  NOR2_X1    g16931(.A1(new_n11877_), .A2(pi0751), .ZN(new_n19955_));
  NOR2_X1    g16932(.A1(new_n19955_), .A2(new_n19954_), .ZN(new_n19956_));
  AOI21_X1   g16933(.A1(new_n11886_), .A2(new_n15564_), .B(new_n19954_), .ZN(new_n19957_));
  NOR2_X1    g16934(.A1(new_n19957_), .A2(new_n11874_), .ZN(new_n19958_));
  INV_X1     g16935(.I(new_n19958_), .ZN(new_n19959_));
  NAND2_X1   g16936(.A1(new_n19959_), .A2(new_n19956_), .ZN(new_n19960_));
  NAND2_X1   g16937(.A1(new_n19960_), .A2(new_n11891_), .ZN(new_n19961_));
  NOR2_X1    g16938(.A1(new_n19959_), .A2(new_n12970_), .ZN(new_n19962_));
  NOR4_X1    g16939(.A1(new_n19962_), .A2(new_n11893_), .A3(new_n19954_), .A4(new_n19955_), .ZN(new_n19963_));
  NOR3_X1    g16940(.A1(new_n11894_), .A2(pi0625), .A3(pi0701), .ZN(new_n19964_));
  NOR2_X1    g16941(.A1(new_n19954_), .A2(pi1153), .ZN(new_n19965_));
  INV_X1     g16942(.I(new_n19965_), .ZN(new_n19966_));
  NOR2_X1    g16943(.A1(new_n19964_), .A2(new_n19966_), .ZN(new_n19967_));
  INV_X1     g16944(.I(new_n19967_), .ZN(new_n19968_));
  NAND2_X1   g16945(.A1(new_n19968_), .A2(pi0608), .ZN(new_n19969_));
  INV_X1     g16946(.I(new_n19962_), .ZN(new_n19970_));
  AOI21_X1   g16947(.A1(new_n19970_), .A2(new_n19960_), .B(new_n19966_), .ZN(new_n19971_));
  OAI21_X1   g16948(.A1(new_n19964_), .A2(new_n19957_), .B(pi1153), .ZN(new_n19972_));
  NAND2_X1   g16949(.A1(new_n19972_), .A2(new_n13657_), .ZN(new_n19973_));
  OAI22_X1   g16950(.A1(new_n19971_), .A2(new_n19973_), .B1(new_n19963_), .B2(new_n19969_), .ZN(new_n19974_));
  NAND2_X1   g16951(.A1(new_n19974_), .A2(pi0778), .ZN(new_n19975_));
  XOR2_X1    g16952(.A1(new_n19975_), .A2(new_n19961_), .Z(new_n19976_));
  INV_X1     g16953(.I(new_n19976_), .ZN(new_n19977_));
  NAND2_X1   g16954(.A1(new_n19968_), .A2(new_n19972_), .ZN(new_n19978_));
  MUX2_X1    g16955(.I0(new_n19978_), .I1(new_n19957_), .S(new_n11891_), .Z(new_n19979_));
  XNOR2_X1   g16956(.A1(new_n19976_), .A2(new_n19979_), .ZN(new_n19980_));
  NAND2_X1   g16957(.A1(new_n19980_), .A2(pi0609), .ZN(new_n19981_));
  XOR2_X1    g16958(.A1(new_n19981_), .A2(new_n19976_), .Z(new_n19982_));
  NAND2_X1   g16959(.A1(new_n19982_), .A2(new_n11912_), .ZN(new_n19983_));
  NOR2_X1    g16960(.A1(new_n19956_), .A2(new_n11925_), .ZN(new_n19984_));
  INV_X1     g16961(.I(new_n19984_), .ZN(new_n19985_));
  NOR3_X1    g16962(.A1(new_n12997_), .A2(new_n11877_), .A3(pi0751), .ZN(new_n19986_));
  NAND3_X1   g16963(.A1(new_n19985_), .A2(new_n11912_), .A3(new_n19986_), .ZN(new_n19987_));
  NAND3_X1   g16964(.A1(new_n19983_), .A2(new_n11923_), .A3(new_n19987_), .ZN(new_n19988_));
  NOR4_X1    g16965(.A1(new_n19986_), .A2(new_n11923_), .A3(pi1155), .A4(new_n19954_), .ZN(new_n19990_));
  NOR2_X1    g16966(.A1(new_n19990_), .A2(new_n11870_), .ZN(new_n19991_));
  AOI22_X1   g16967(.A1(new_n19988_), .A2(new_n19991_), .B1(new_n11870_), .B2(new_n19977_), .ZN(new_n19992_));
  NOR2_X1    g16968(.A1(new_n19992_), .A2(pi0781), .ZN(new_n19993_));
  NOR4_X1    g16969(.A1(new_n19979_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n19994_));
  NOR3_X1    g16970(.A1(new_n19986_), .A2(pi1155), .A3(new_n19954_), .ZN(new_n19995_));
  NAND2_X1   g16971(.A1(new_n19987_), .A2(new_n19995_), .ZN(new_n19996_));
  MUX2_X1    g16972(.I0(new_n19996_), .I1(new_n19985_), .S(new_n11870_), .Z(new_n19997_));
  INV_X1     g16973(.I(new_n19997_), .ZN(new_n19998_));
  OAI21_X1   g16974(.A1(new_n19998_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n19999_));
  OAI21_X1   g16975(.A1(new_n19998_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n20000_));
  NOR2_X1    g16976(.A1(new_n19979_), .A2(new_n11939_), .ZN(new_n20001_));
  NOR4_X1    g16977(.A1(new_n19992_), .A2(new_n11934_), .A3(pi1154), .A4(new_n20001_), .ZN(new_n20002_));
  NOR2_X1    g16978(.A1(new_n20002_), .A2(new_n20000_), .ZN(new_n20003_));
  OAI22_X1   g16979(.A1(new_n20003_), .A2(pi0627), .B1(new_n19994_), .B2(new_n19999_), .ZN(new_n20004_));
  AOI21_X1   g16980(.A1(new_n20004_), .A2(pi0781), .B(new_n19993_), .ZN(new_n20005_));
  INV_X1     g16981(.I(new_n20001_), .ZN(new_n20006_));
  NOR2_X1    g16982(.A1(new_n20006_), .A2(new_n11962_), .ZN(new_n20007_));
  NOR4_X1    g16983(.A1(new_n20005_), .A2(new_n11967_), .A3(pi1159), .A4(new_n20007_), .ZN(new_n20008_));
  NOR2_X1    g16984(.A1(new_n19998_), .A2(pi0781), .ZN(new_n20009_));
  AOI21_X1   g16985(.A1(new_n11944_), .A2(new_n19997_), .B(new_n20000_), .ZN(new_n20010_));
  NOR2_X1    g16986(.A1(new_n20010_), .A2(new_n11969_), .ZN(new_n20011_));
  XOR2_X1    g16987(.A1(new_n20011_), .A2(new_n20009_), .Z(new_n20012_));
  AOI21_X1   g16988(.A1(new_n20012_), .A2(new_n16479_), .B(pi1159), .ZN(new_n20013_));
  INV_X1     g16989(.I(new_n20013_), .ZN(new_n20014_));
  NOR3_X1    g16990(.A1(new_n20008_), .A2(new_n11966_), .A3(new_n20014_), .ZN(new_n20015_));
  NOR4_X1    g16991(.A1(new_n20006_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n20016_));
  INV_X1     g16992(.I(new_n20012_), .ZN(new_n20017_));
  NOR2_X1    g16993(.A1(new_n20017_), .A2(new_n16482_), .ZN(new_n20018_));
  NOR3_X1    g16994(.A1(new_n20018_), .A2(pi0648), .A3(new_n20016_), .ZN(new_n20019_));
  AOI21_X1   g16995(.A1(new_n20005_), .A2(new_n11998_), .B(pi0789), .ZN(new_n20020_));
  OAI21_X1   g16996(.A1(new_n20015_), .A2(new_n20019_), .B(new_n20020_), .ZN(new_n20021_));
  NAND2_X1   g16997(.A1(new_n20007_), .A2(new_n17450_), .ZN(new_n20022_));
  NOR2_X1    g16998(.A1(new_n20022_), .A2(new_n17153_), .ZN(new_n20023_));
  NOR2_X1    g16999(.A1(new_n14624_), .A2(new_n19954_), .ZN(new_n20024_));
  NOR2_X1    g17000(.A1(new_n20017_), .A2(pi0789), .ZN(new_n20025_));
  NOR2_X1    g17001(.A1(new_n20014_), .A2(new_n20018_), .ZN(new_n20026_));
  NOR2_X1    g17002(.A1(new_n20026_), .A2(new_n11985_), .ZN(new_n20027_));
  XOR2_X1    g17003(.A1(new_n20027_), .A2(new_n20025_), .Z(new_n20028_));
  AOI21_X1   g17004(.A1(new_n20028_), .A2(new_n14624_), .B(new_n20024_), .ZN(new_n20029_));
  AOI22_X1   g17005(.A1(new_n20029_), .A2(new_n12064_), .B1(new_n15080_), .B2(new_n20023_), .ZN(new_n20030_));
  NOR2_X1    g17006(.A1(new_n20030_), .A2(new_n12030_), .ZN(new_n20031_));
  NAND2_X1   g17007(.A1(new_n20029_), .A2(new_n12063_), .ZN(new_n20032_));
  AOI21_X1   g17008(.A1(new_n20023_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n20033_));
  NAND2_X1   g17009(.A1(new_n20032_), .A2(new_n20033_), .ZN(new_n20034_));
  OAI21_X1   g17010(.A1(new_n20031_), .A2(new_n20034_), .B(new_n14726_), .ZN(new_n20035_));
  INV_X1     g17011(.I(new_n19954_), .ZN(new_n20036_));
  MUX2_X1    g17012(.I0(new_n20028_), .I1(new_n20036_), .S(new_n11994_), .Z(new_n20037_));
  INV_X1     g17013(.I(new_n20028_), .ZN(new_n20038_));
  AOI21_X1   g17014(.A1(new_n20038_), .A2(new_n20036_), .B(new_n11994_), .ZN(new_n20039_));
  OAI21_X1   g17015(.A1(new_n20022_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n20040_));
  AOI21_X1   g17016(.A1(new_n20039_), .A2(new_n11990_), .B(new_n20040_), .ZN(new_n20041_));
  OAI21_X1   g17017(.A1(new_n17167_), .A2(new_n20037_), .B(new_n20041_), .ZN(new_n20042_));
  NAND4_X1   g17018(.A1(new_n20021_), .A2(new_n14732_), .A3(new_n20035_), .A4(new_n20042_), .ZN(new_n20043_));
  NAND3_X1   g17019(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n19954_), .ZN(new_n20044_));
  NAND2_X1   g17020(.A1(new_n20023_), .A2(new_n15050_), .ZN(new_n20045_));
  NAND2_X1   g17021(.A1(new_n20045_), .A2(pi0647), .ZN(new_n20046_));
  NAND2_X1   g17022(.A1(new_n19954_), .A2(pi0647), .ZN(new_n20047_));
  NAND3_X1   g17023(.A1(new_n20046_), .A2(new_n12049_), .A3(new_n20047_), .ZN(new_n20048_));
  NAND2_X1   g17024(.A1(new_n20048_), .A2(pi0630), .ZN(new_n20049_));
  NOR2_X1    g17025(.A1(new_n20045_), .A2(new_n12061_), .ZN(new_n20050_));
  AOI21_X1   g17026(.A1(new_n12061_), .A2(new_n19954_), .B(new_n20050_), .ZN(new_n20051_));
  NAND2_X1   g17027(.A1(new_n20051_), .A2(new_n12088_), .ZN(new_n20052_));
  NAND4_X1   g17028(.A1(new_n20052_), .A2(new_n20049_), .A3(pi0787), .A4(new_n20044_), .ZN(new_n20053_));
  AND2_X2    g17029(.A1(new_n20043_), .A2(new_n20053_), .Z(new_n20054_));
  NOR2_X1    g17030(.A1(new_n20054_), .A2(new_n12082_), .ZN(new_n20055_));
  NAND4_X1   g17031(.A1(new_n20046_), .A2(pi0787), .A3(new_n12049_), .A4(new_n20047_), .ZN(new_n20056_));
  OAI21_X1   g17032(.A1(pi0787), .A2(new_n20045_), .B(new_n20056_), .ZN(new_n20057_));
  NOR2_X1    g17033(.A1(new_n20057_), .A2(pi0644), .ZN(new_n20058_));
  OR3_X2     g17034(.A1(new_n20055_), .A2(pi0715), .A3(new_n20058_), .Z(new_n20059_));
  MUX2_X1    g17035(.I0(new_n20029_), .I1(new_n19954_), .S(new_n16841_), .Z(new_n20060_));
  INV_X1     g17036(.I(new_n20060_), .ZN(new_n20061_));
  OAI21_X1   g17037(.A1(new_n20060_), .A2(new_n19954_), .B(new_n12082_), .ZN(new_n20062_));
  AOI21_X1   g17038(.A1(new_n19954_), .A2(new_n20060_), .B(new_n20062_), .ZN(new_n20063_));
  OAI21_X1   g17039(.A1(new_n20063_), .A2(new_n20061_), .B(new_n12099_), .ZN(new_n20064_));
  AOI21_X1   g17040(.A1(new_n20061_), .A2(new_n20063_), .B(new_n20064_), .ZN(new_n20065_));
  AOI21_X1   g17041(.A1(new_n20059_), .A2(new_n20065_), .B(pi1160), .ZN(new_n20066_));
  XOR2_X1    g17042(.A1(new_n20063_), .A2(new_n19954_), .Z(new_n20067_));
  AOI21_X1   g17043(.A1(new_n20057_), .A2(pi0644), .B(new_n13169_), .ZN(new_n20068_));
  OAI21_X1   g17044(.A1(new_n20067_), .A2(new_n12099_), .B(new_n20068_), .ZN(new_n20069_));
  OAI21_X1   g17045(.A1(new_n20055_), .A2(new_n20069_), .B(pi0790), .ZN(new_n20070_));
  NOR2_X1    g17046(.A1(new_n20054_), .A2(new_n14748_), .ZN(new_n20071_));
  OAI21_X1   g17047(.A1(new_n20066_), .A2(new_n20070_), .B(new_n20071_), .ZN(new_n20072_));
  NOR2_X1    g17048(.A1(new_n12965_), .A2(pi0185), .ZN(new_n20073_));
  INV_X1     g17049(.I(new_n20073_), .ZN(new_n20074_));
  NAND2_X1   g17050(.A1(new_n20074_), .A2(new_n11997_), .ZN(new_n20075_));
  NAND2_X1   g17051(.A1(new_n12894_), .A2(pi0751), .ZN(new_n20076_));
  NOR2_X1    g17052(.A1(new_n15546_), .A2(pi0185), .ZN(new_n20077_));
  OAI21_X1   g17053(.A1(new_n14361_), .A2(new_n10066_), .B(pi0039), .ZN(new_n20080_));
  AOI21_X1   g17054(.A1(new_n12824_), .A2(new_n20077_), .B(new_n20080_), .ZN(new_n20081_));
  NOR2_X1    g17055(.A1(new_n12828_), .A2(pi0185), .ZN(new_n20082_));
  AOI21_X1   g17056(.A1(new_n12829_), .A2(new_n15546_), .B(pi0038), .ZN(new_n20083_));
  INV_X1     g17057(.I(new_n20083_), .ZN(new_n20084_));
  AOI21_X1   g17058(.A1(new_n20081_), .A2(new_n20076_), .B(new_n20084_), .ZN(new_n20085_));
  NOR2_X1    g17059(.A1(new_n20085_), .A2(new_n3232_), .ZN(new_n20086_));
  AOI21_X1   g17060(.A1(new_n10066_), .A2(new_n3232_), .B(new_n20086_), .ZN(new_n20087_));
  OAI21_X1   g17061(.A1(new_n20087_), .A2(new_n11914_), .B(new_n11870_), .ZN(new_n20088_));
  AOI21_X1   g17062(.A1(new_n11914_), .A2(new_n20073_), .B(new_n20088_), .ZN(new_n20089_));
  NAND2_X1   g17063(.A1(new_n20087_), .A2(new_n11924_), .ZN(new_n20090_));
  OAI22_X1   g17064(.A1(new_n20090_), .A2(pi0609), .B1(new_n12996_), .B2(new_n20073_), .ZN(new_n20091_));
  NAND2_X1   g17065(.A1(new_n20091_), .A2(new_n11912_), .ZN(new_n20092_));
  OAI22_X1   g17066(.A1(new_n20090_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n20073_), .ZN(new_n20093_));
  NAND2_X1   g17067(.A1(new_n20093_), .A2(pi1155), .ZN(new_n20094_));
  AOI21_X1   g17068(.A1(new_n20092_), .A2(new_n20094_), .B(new_n11870_), .ZN(new_n20095_));
  XNOR2_X1   g17069(.A1(new_n20095_), .A2(new_n20089_), .ZN(new_n20096_));
  NOR2_X1    g17070(.A1(new_n20096_), .A2(pi0781), .ZN(new_n20097_));
  NOR3_X1    g17071(.A1(new_n20073_), .A2(pi0618), .A3(pi1154), .ZN(new_n20098_));
  NOR2_X1    g17072(.A1(new_n20098_), .A2(new_n11969_), .ZN(new_n20099_));
  XOR2_X1    g17073(.A1(new_n20097_), .A2(new_n20099_), .Z(new_n20100_));
  NAND2_X1   g17074(.A1(new_n20100_), .A2(new_n11985_), .ZN(new_n20101_));
  NAND3_X1   g17075(.A1(new_n20074_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n20102_));
  NAND2_X1   g17076(.A1(new_n20102_), .A2(pi0789), .ZN(new_n20103_));
  XNOR2_X1   g17077(.A1(new_n20101_), .A2(new_n20103_), .ZN(new_n20104_));
  OAI21_X1   g17078(.A1(new_n20104_), .A2(new_n11997_), .B(new_n20075_), .ZN(new_n20105_));
  NOR2_X1    g17079(.A1(new_n20073_), .A2(new_n12054_), .ZN(new_n20106_));
  AOI21_X1   g17080(.A1(new_n20105_), .A2(new_n12054_), .B(new_n20106_), .ZN(new_n20107_));
  NAND2_X1   g17081(.A1(new_n20074_), .A2(new_n12091_), .ZN(new_n20108_));
  OAI21_X1   g17082(.A1(new_n20107_), .A2(new_n12091_), .B(new_n20108_), .ZN(new_n20109_));
  OR2_X2     g17083(.A1(new_n20109_), .A2(pi0644), .Z(new_n20110_));
  AOI21_X1   g17084(.A1(new_n20073_), .A2(pi0644), .B(new_n12099_), .ZN(new_n20111_));
  AOI21_X1   g17085(.A1(new_n20110_), .A2(new_n20111_), .B(pi1160), .ZN(new_n20112_));
  NOR2_X1    g17086(.A1(new_n20073_), .A2(new_n13114_), .ZN(new_n20113_));
  NOR2_X1    g17087(.A1(new_n20074_), .A2(new_n12014_), .ZN(new_n20114_));
  NOR2_X1    g17088(.A1(new_n20073_), .A2(new_n11961_), .ZN(new_n20115_));
  OAI21_X1   g17089(.A1(new_n15189_), .A2(new_n20082_), .B(new_n15564_), .ZN(new_n20116_));
  NOR2_X1    g17090(.A1(new_n13395_), .A2(new_n10066_), .ZN(new_n20117_));
  NOR2_X1    g17091(.A1(new_n20117_), .A2(pi0038), .ZN(new_n20118_));
  OAI22_X1   g17092(.A1(new_n20118_), .A2(new_n3232_), .B1(pi0185), .B2(new_n13399_), .ZN(new_n20119_));
  NOR2_X1    g17093(.A1(new_n3232_), .A2(pi0701), .ZN(new_n20120_));
  AOI22_X1   g17094(.A1(new_n20074_), .A2(new_n20120_), .B1(new_n20116_), .B2(new_n20119_), .ZN(new_n20121_));
  NOR3_X1    g17095(.A1(new_n20074_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n20122_));
  NOR4_X1    g17096(.A1(new_n20121_), .A2(new_n12970_), .A3(pi1153), .A4(new_n20073_), .ZN(new_n20123_));
  NOR2_X1    g17097(.A1(new_n20123_), .A2(new_n20122_), .ZN(new_n20124_));
  MUX2_X1    g17098(.I0(new_n20124_), .I1(new_n20121_), .S(new_n11891_), .Z(new_n20125_));
  INV_X1     g17099(.I(new_n20125_), .ZN(new_n20126_));
  NOR2_X1    g17100(.A1(new_n20074_), .A2(new_n11938_), .ZN(new_n20127_));
  AOI21_X1   g17101(.A1(new_n20126_), .A2(new_n11938_), .B(new_n20127_), .ZN(new_n20128_));
  AOI21_X1   g17102(.A1(new_n20128_), .A2(new_n11961_), .B(new_n20115_), .ZN(new_n20129_));
  AOI21_X1   g17103(.A1(new_n20129_), .A2(new_n12014_), .B(new_n20114_), .ZN(new_n20130_));
  AOI21_X1   g17104(.A1(new_n20130_), .A2(new_n13114_), .B(new_n20113_), .ZN(new_n20131_));
  NOR3_X1    g17105(.A1(new_n20074_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n20132_));
  NOR4_X1    g17106(.A1(new_n20131_), .A2(new_n12031_), .A3(pi1156), .A4(new_n20073_), .ZN(new_n20133_));
  NOR2_X1    g17107(.A1(new_n20133_), .A2(new_n20132_), .ZN(new_n20134_));
  MUX2_X1    g17108(.I0(new_n20134_), .I1(new_n20131_), .S(new_n11868_), .Z(new_n20135_));
  NOR2_X1    g17109(.A1(new_n20135_), .A2(new_n12061_), .ZN(new_n20136_));
  AOI21_X1   g17110(.A1(new_n12061_), .A2(new_n20073_), .B(new_n20136_), .ZN(new_n20137_));
  NAND2_X1   g17111(.A1(new_n20137_), .A2(pi1157), .ZN(new_n20138_));
  NOR2_X1    g17112(.A1(new_n20135_), .A2(pi0647), .ZN(new_n20139_));
  AOI21_X1   g17113(.A1(pi0647), .A2(new_n20073_), .B(new_n20139_), .ZN(new_n20140_));
  NAND2_X1   g17114(.A1(new_n20140_), .A2(new_n12049_), .ZN(new_n20141_));
  AOI21_X1   g17115(.A1(new_n20141_), .A2(new_n20138_), .B(new_n12048_), .ZN(new_n20142_));
  AOI21_X1   g17116(.A1(new_n12048_), .A2(new_n20135_), .B(new_n20142_), .ZN(new_n20143_));
  NAND2_X1   g17117(.A1(new_n20143_), .A2(pi0644), .ZN(new_n20144_));
  AOI21_X1   g17118(.A1(new_n20144_), .A2(new_n12099_), .B(new_n20112_), .ZN(new_n20145_));
  NAND3_X1   g17119(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n20146_));
  OAI21_X1   g17120(.A1(new_n20109_), .A2(new_n20146_), .B(pi0715), .ZN(new_n20147_));
  AOI21_X1   g17121(.A1(new_n20143_), .A2(new_n12082_), .B(new_n20147_), .ZN(new_n20148_));
  OAI21_X1   g17122(.A1(new_n20145_), .A2(new_n20148_), .B(pi0790), .ZN(new_n20149_));
  NAND2_X1   g17123(.A1(new_n20100_), .A2(pi0619), .ZN(new_n20150_));
  NAND2_X1   g17124(.A1(new_n20073_), .A2(pi0619), .ZN(new_n20151_));
  INV_X1     g17125(.I(new_n20123_), .ZN(new_n20152_));
  INV_X1     g17126(.I(new_n20087_), .ZN(new_n20153_));
  OR3_X2     g17127(.A1(new_n20085_), .A2(new_n15564_), .A3(new_n3231_), .Z(new_n20163_));
  OAI21_X1   g17128(.A1(new_n10066_), .A2(new_n3231_), .B(new_n20163_), .ZN(new_n20164_));
  OAI21_X1   g17129(.A1(new_n20164_), .A2(pi0625), .B(new_n20153_), .ZN(new_n20165_));
  NAND3_X1   g17130(.A1(new_n20164_), .A2(new_n12970_), .A3(new_n20087_), .ZN(new_n20166_));
  NAND4_X1   g17131(.A1(new_n20152_), .A2(new_n12977_), .A3(new_n20165_), .A4(new_n20166_), .ZN(new_n20167_));
  NOR4_X1    g17132(.A1(new_n20164_), .A2(new_n20153_), .A3(new_n12970_), .A4(pi1153), .ZN(new_n20168_));
  OAI21_X1   g17133(.A1(new_n20168_), .A2(new_n20122_), .B(new_n13657_), .ZN(new_n20169_));
  NAND2_X1   g17134(.A1(new_n20167_), .A2(new_n20169_), .ZN(new_n20170_));
  NOR2_X1    g17135(.A1(new_n20164_), .A2(pi0778), .ZN(new_n20171_));
  AOI21_X1   g17136(.A1(new_n20170_), .A2(pi0778), .B(new_n20171_), .ZN(new_n20172_));
  NOR2_X1    g17137(.A1(new_n20172_), .A2(pi0785), .ZN(new_n20173_));
  NAND3_X1   g17138(.A1(new_n20126_), .A2(pi0609), .A3(pi1155), .ZN(new_n20174_));
  NAND3_X1   g17139(.A1(new_n20174_), .A2(new_n11923_), .A3(new_n20094_), .ZN(new_n20175_));
  NAND2_X1   g17140(.A1(new_n20172_), .A2(pi0609), .ZN(new_n20176_));
  NAND3_X1   g17141(.A1(new_n20176_), .A2(new_n13621_), .A3(new_n20125_), .ZN(new_n20177_));
  NAND3_X1   g17142(.A1(new_n20177_), .A2(pi0660), .A3(new_n20092_), .ZN(new_n20178_));
  AND3_X2    g17143(.A1(new_n20178_), .A2(pi0785), .A3(new_n20175_), .Z(new_n20179_));
  NOR2_X1    g17144(.A1(new_n20179_), .A2(new_n20173_), .ZN(new_n20180_));
  NAND2_X1   g17145(.A1(new_n20180_), .A2(new_n11969_), .ZN(new_n20181_));
  NAND2_X1   g17146(.A1(new_n20180_), .A2(pi0618), .ZN(new_n20182_));
  AND2_X2    g17147(.A1(new_n20128_), .A2(new_n14633_), .Z(new_n20183_));
  NOR2_X1    g17148(.A1(new_n20096_), .A2(new_n11934_), .ZN(new_n20184_));
  OAI21_X1   g17149(.A1(new_n20074_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n20185_));
  OR3_X2     g17150(.A1(new_n20184_), .A2(new_n11949_), .A3(new_n20185_), .Z(new_n20186_));
  AOI21_X1   g17151(.A1(new_n20182_), .A2(new_n20183_), .B(new_n20186_), .ZN(new_n20187_));
  NOR3_X1    g17152(.A1(new_n20128_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n20188_));
  OAI21_X1   g17153(.A1(new_n20073_), .A2(pi0618), .B(new_n11950_), .ZN(new_n20189_));
  OAI21_X1   g17154(.A1(new_n20184_), .A2(new_n20189_), .B(new_n11949_), .ZN(new_n20190_));
  NOR2_X1    g17155(.A1(new_n20190_), .A2(new_n20188_), .ZN(new_n20191_));
  OAI21_X1   g17156(.A1(new_n20187_), .A2(new_n20191_), .B(pi0781), .ZN(new_n20192_));
  XOR2_X1    g17157(.A1(new_n20192_), .A2(new_n20181_), .Z(new_n20193_));
  XNOR2_X1   g17158(.A1(new_n20193_), .A2(new_n20129_), .ZN(new_n20194_));
  NOR2_X1    g17159(.A1(new_n20194_), .A2(new_n11967_), .ZN(new_n20195_));
  NAND3_X1   g17160(.A1(new_n20150_), .A2(new_n11869_), .A3(new_n20151_), .ZN(new_n20196_));
  XNOR2_X1   g17161(.A1(new_n20195_), .A2(new_n20193_), .ZN(new_n20197_));
  NAND2_X1   g17162(.A1(new_n20197_), .A2(new_n11869_), .ZN(new_n20198_));
  AOI21_X1   g17163(.A1(new_n20074_), .A2(new_n11967_), .B(pi1159), .ZN(new_n20199_));
  AOI21_X1   g17164(.A1(new_n20150_), .A2(new_n20199_), .B(pi0648), .ZN(new_n20200_));
  OAI21_X1   g17165(.A1(new_n20193_), .A2(pi0789), .B(new_n11998_), .ZN(new_n20201_));
  MUX2_X1    g17166(.I0(new_n20104_), .I1(new_n20073_), .S(new_n11994_), .Z(new_n20202_));
  NAND2_X1   g17167(.A1(new_n20202_), .A2(new_n11988_), .ZN(new_n20203_));
  AOI21_X1   g17168(.A1(new_n20104_), .A2(new_n20074_), .B(new_n11994_), .ZN(new_n20204_));
  OAI21_X1   g17169(.A1(new_n20130_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n20205_));
  AOI21_X1   g17170(.A1(new_n20204_), .A2(new_n11990_), .B(new_n20205_), .ZN(new_n20206_));
  AOI21_X1   g17171(.A1(new_n20203_), .A2(new_n20206_), .B(new_n18842_), .ZN(new_n20207_));
  NAND2_X1   g17172(.A1(new_n20201_), .A2(new_n20207_), .ZN(new_n20208_));
  AOI21_X1   g17173(.A1(new_n20198_), .A2(new_n20200_), .B(new_n20208_), .ZN(new_n20209_));
  NOR2_X1    g17174(.A1(new_n20132_), .A2(new_n12030_), .ZN(new_n20210_));
  NOR2_X1    g17175(.A1(new_n20133_), .A2(pi0629), .ZN(new_n20211_));
  NAND2_X1   g17176(.A1(new_n20105_), .A2(new_n15222_), .ZN(new_n20212_));
  OAI21_X1   g17177(.A1(new_n20210_), .A2(new_n20211_), .B(new_n20212_), .ZN(new_n20213_));
  AOI22_X1   g17178(.A1(new_n20209_), .A2(new_n20196_), .B1(pi0792), .B2(new_n20213_), .ZN(new_n20214_));
  NAND2_X1   g17179(.A1(new_n20137_), .A2(new_n12060_), .ZN(new_n20215_));
  AOI21_X1   g17180(.A1(new_n20140_), .A2(pi0630), .B(new_n15214_), .ZN(new_n20216_));
  NAND2_X1   g17181(.A1(new_n20216_), .A2(new_n20215_), .ZN(new_n20217_));
  NOR2_X1    g17182(.A1(new_n20107_), .A2(new_n15183_), .ZN(new_n20218_));
  OAI21_X1   g17183(.A1(new_n20109_), .A2(new_n20146_), .B(pi0644), .ZN(new_n20219_));
  NAND2_X1   g17184(.A1(new_n20219_), .A2(new_n11867_), .ZN(new_n20220_));
  AOI21_X1   g17185(.A1(new_n20112_), .A2(new_n12082_), .B(new_n20220_), .ZN(new_n20221_));
  AOI21_X1   g17186(.A1(new_n20217_), .A2(new_n20218_), .B(new_n20221_), .ZN(new_n20222_));
  OAI21_X1   g17187(.A1(new_n20214_), .A2(new_n14725_), .B(new_n20222_), .ZN(new_n20223_));
  AOI21_X1   g17188(.A1(new_n20223_), .A2(new_n20149_), .B(po1038), .ZN(new_n20224_));
  OAI21_X1   g17189(.A1(new_n6845_), .A2(pi0185), .B(new_n13184_), .ZN(new_n20225_));
  OAI21_X1   g17190(.A1(new_n20224_), .A2(new_n20225_), .B(new_n20072_), .ZN(po0342));
  NOR2_X1    g17191(.A1(new_n2925_), .A2(pi0186), .ZN(new_n20227_));
  NOR2_X1    g17192(.A1(new_n11877_), .A2(pi0752), .ZN(new_n20228_));
  NOR2_X1    g17193(.A1(new_n20228_), .A2(new_n20227_), .ZN(new_n20229_));
  INV_X1     g17194(.I(new_n20229_), .ZN(new_n20230_));
  AOI21_X1   g17195(.A1(new_n11886_), .A2(pi0703), .B(new_n20227_), .ZN(new_n20231_));
  NOR2_X1    g17196(.A1(new_n20231_), .A2(new_n11874_), .ZN(new_n20232_));
  NOR2_X1    g17197(.A1(new_n20230_), .A2(new_n20232_), .ZN(new_n20233_));
  NOR2_X1    g17198(.A1(new_n20233_), .A2(pi0778), .ZN(new_n20234_));
  NAND2_X1   g17199(.A1(new_n20232_), .A2(pi0625), .ZN(new_n20235_));
  NOR2_X1    g17200(.A1(new_n13201_), .A2(new_n16094_), .ZN(new_n20236_));
  NOR4_X1    g17201(.A1(new_n20228_), .A2(pi0608), .A3(new_n11893_), .A4(new_n20227_), .ZN(new_n20237_));
  OAI21_X1   g17202(.A1(new_n20230_), .A2(new_n20232_), .B(new_n20235_), .ZN(new_n20238_));
  NOR3_X1    g17203(.A1(new_n20227_), .A2(pi0608), .A3(pi1153), .ZN(new_n20239_));
  AOI22_X1   g17204(.A1(new_n20238_), .A2(new_n20239_), .B1(new_n20235_), .B2(new_n20237_), .ZN(new_n20240_));
  NOR2_X1    g17205(.A1(new_n20240_), .A2(new_n11891_), .ZN(new_n20241_));
  XOR2_X1    g17206(.A1(new_n20241_), .A2(new_n20234_), .Z(new_n20242_));
  INV_X1     g17207(.I(new_n20242_), .ZN(new_n20243_));
  NAND2_X1   g17208(.A1(new_n20243_), .A2(new_n11870_), .ZN(new_n20244_));
  AOI21_X1   g17209(.A1(new_n20242_), .A2(new_n11903_), .B(pi1155), .ZN(new_n20245_));
  INV_X1     g17210(.I(new_n20231_), .ZN(new_n20246_));
  XOR2_X1    g17211(.A1(new_n20236_), .A2(pi1153), .Z(new_n20247_));
  NAND2_X1   g17212(.A1(new_n20247_), .A2(new_n20246_), .ZN(new_n20248_));
  OAI21_X1   g17213(.A1(new_n20236_), .A2(new_n20227_), .B(new_n11893_), .ZN(new_n20249_));
  AOI21_X1   g17214(.A1(new_n20248_), .A2(new_n20249_), .B(new_n11891_), .ZN(new_n20250_));
  NOR2_X1    g17215(.A1(new_n20231_), .A2(pi0778), .ZN(new_n20251_));
  OAI21_X1   g17216(.A1(new_n20250_), .A2(new_n20251_), .B(pi0609), .ZN(new_n20252_));
  AOI21_X1   g17217(.A1(new_n20230_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n20253_));
  NOR2_X1    g17218(.A1(new_n20253_), .A2(pi0660), .ZN(new_n20254_));
  OAI21_X1   g17219(.A1(new_n20245_), .A2(new_n20252_), .B(new_n20254_), .ZN(new_n20255_));
  NOR2_X1    g17220(.A1(new_n20250_), .A2(new_n20251_), .ZN(new_n20256_));
  NAND4_X1   g17221(.A1(new_n20243_), .A2(pi0609), .A3(new_n11912_), .A4(new_n20256_), .ZN(new_n20257_));
  NOR2_X1    g17222(.A1(new_n20229_), .A2(new_n11925_), .ZN(new_n20258_));
  AOI21_X1   g17223(.A1(new_n20258_), .A2(new_n11928_), .B(pi1155), .ZN(new_n20259_));
  NOR2_X1    g17224(.A1(new_n20259_), .A2(new_n11923_), .ZN(new_n20260_));
  NAND2_X1   g17225(.A1(new_n20257_), .A2(new_n20260_), .ZN(new_n20261_));
  NAND3_X1   g17226(.A1(new_n20261_), .A2(pi0785), .A3(new_n20255_), .ZN(new_n20262_));
  NAND2_X1   g17227(.A1(new_n20262_), .A2(new_n20244_), .ZN(new_n20263_));
  NOR4_X1    g17228(.A1(new_n20256_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n20265_));
  NOR2_X1    g17229(.A1(new_n20258_), .A2(pi0785), .ZN(new_n20266_));
  OAI21_X1   g17230(.A1(new_n20259_), .A2(new_n20253_), .B(pi0785), .ZN(new_n20267_));
  XNOR2_X1   g17231(.A1(new_n20267_), .A2(new_n20266_), .ZN(new_n20268_));
  INV_X1     g17232(.I(new_n20268_), .ZN(new_n20269_));
  NOR2_X1    g17233(.A1(new_n20269_), .A2(new_n11945_), .ZN(new_n20270_));
  NOR3_X1    g17234(.A1(new_n20265_), .A2(new_n20270_), .A3(pi0627), .ZN(new_n20271_));
  AOI21_X1   g17235(.A1(new_n20268_), .A2(new_n11951_), .B(pi1154), .ZN(new_n20272_));
  NOR2_X1    g17236(.A1(new_n20256_), .A2(new_n11939_), .ZN(new_n20273_));
  INV_X1     g17237(.I(new_n20273_), .ZN(new_n20274_));
  NAND4_X1   g17238(.A1(new_n20263_), .A2(pi0618), .A3(new_n11950_), .A4(new_n20274_), .ZN(new_n20275_));
  NAND2_X1   g17239(.A1(new_n20275_), .A2(new_n20272_), .ZN(new_n20276_));
  AOI21_X1   g17240(.A1(new_n20276_), .A2(new_n11949_), .B(new_n20271_), .ZN(new_n20277_));
  NOR2_X1    g17241(.A1(new_n20277_), .A2(new_n11969_), .ZN(new_n20278_));
  AOI21_X1   g17242(.A1(new_n11969_), .A2(new_n20263_), .B(new_n20278_), .ZN(new_n20279_));
  NOR2_X1    g17243(.A1(new_n20274_), .A2(new_n11962_), .ZN(new_n20280_));
  NOR4_X1    g17244(.A1(new_n20279_), .A2(new_n11967_), .A3(pi1159), .A4(new_n20280_), .ZN(new_n20281_));
  INV_X1     g17245(.I(new_n20270_), .ZN(new_n20282_));
  NAND2_X1   g17246(.A1(new_n20282_), .A2(new_n20272_), .ZN(new_n20283_));
  MUX2_X1    g17247(.I0(new_n20283_), .I1(new_n20268_), .S(new_n11969_), .Z(new_n20284_));
  NAND2_X1   g17248(.A1(new_n20284_), .A2(pi0619), .ZN(new_n20285_));
  INV_X1     g17249(.I(new_n20285_), .ZN(new_n20286_));
  INV_X1     g17250(.I(new_n20227_), .ZN(new_n20287_));
  OAI21_X1   g17251(.A1(new_n20287_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n20288_));
  NOR4_X1    g17252(.A1(new_n20281_), .A2(new_n11966_), .A3(new_n20286_), .A4(new_n20288_), .ZN(new_n20289_));
  NOR4_X1    g17253(.A1(new_n20274_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n20290_));
  OAI21_X1   g17254(.A1(new_n20227_), .A2(pi0619), .B(new_n11869_), .ZN(new_n20291_));
  OAI21_X1   g17255(.A1(new_n20286_), .A2(new_n20291_), .B(new_n11966_), .ZN(new_n20292_));
  NOR2_X1    g17256(.A1(new_n20292_), .A2(new_n20290_), .ZN(new_n20293_));
  AOI21_X1   g17257(.A1(new_n20279_), .A2(new_n11998_), .B(pi0789), .ZN(new_n20294_));
  OAI21_X1   g17258(.A1(new_n20289_), .A2(new_n20293_), .B(new_n20294_), .ZN(new_n20295_));
  NAND2_X1   g17259(.A1(new_n20280_), .A2(new_n17450_), .ZN(new_n20296_));
  NOR2_X1    g17260(.A1(new_n20296_), .A2(new_n17153_), .ZN(new_n20297_));
  INV_X1     g17261(.I(new_n20297_), .ZN(new_n20298_));
  NOR2_X1    g17262(.A1(new_n20298_), .A2(new_n17151_), .ZN(new_n20299_));
  NOR2_X1    g17263(.A1(new_n14624_), .A2(new_n20227_), .ZN(new_n20300_));
  NAND3_X1   g17264(.A1(new_n20287_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n20301_));
  MUX2_X1    g17265(.I0(new_n20301_), .I1(new_n20284_), .S(new_n11985_), .Z(new_n20302_));
  AOI21_X1   g17266(.A1(new_n20302_), .A2(new_n14624_), .B(new_n20300_), .ZN(new_n20303_));
  AND2_X2    g17267(.A1(new_n20303_), .A2(new_n12064_), .Z(new_n20304_));
  OAI21_X1   g17268(.A1(new_n20304_), .A2(new_n20299_), .B(pi0629), .ZN(new_n20305_));
  NAND2_X1   g17269(.A1(new_n20303_), .A2(new_n12063_), .ZN(new_n20306_));
  NAND2_X1   g17270(.A1(new_n20297_), .A2(new_n15084_), .ZN(new_n20307_));
  NAND4_X1   g17271(.A1(new_n20305_), .A2(new_n15085_), .A3(new_n20306_), .A4(new_n20307_), .ZN(new_n20308_));
  MUX2_X1    g17272(.I0(new_n20302_), .I1(new_n20287_), .S(new_n11994_), .Z(new_n20309_));
  NOR2_X1    g17273(.A1(new_n20309_), .A2(new_n17167_), .ZN(new_n20310_));
  OAI21_X1   g17274(.A1(new_n20302_), .A2(new_n20227_), .B(pi0626), .ZN(new_n20311_));
  NOR2_X1    g17275(.A1(new_n20296_), .A2(new_n12020_), .ZN(new_n20312_));
  NOR2_X1    g17276(.A1(new_n20312_), .A2(pi0788), .ZN(new_n20313_));
  OAI21_X1   g17277(.A1(new_n20311_), .A2(new_n17171_), .B(new_n20313_), .ZN(new_n20314_));
  OAI21_X1   g17278(.A1(new_n20310_), .A2(new_n20314_), .B(new_n14732_), .ZN(new_n20315_));
  AOI21_X1   g17279(.A1(new_n20308_), .A2(new_n14726_), .B(new_n20315_), .ZN(new_n20316_));
  NAND3_X1   g17280(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n20227_), .ZN(new_n20317_));
  NOR2_X1    g17281(.A1(new_n20298_), .A2(new_n12068_), .ZN(new_n20318_));
  INV_X1     g17282(.I(new_n20318_), .ZN(new_n20319_));
  NAND2_X1   g17283(.A1(new_n20319_), .A2(pi0647), .ZN(new_n20320_));
  NAND2_X1   g17284(.A1(new_n20227_), .A2(pi0647), .ZN(new_n20321_));
  NAND3_X1   g17285(.A1(new_n20320_), .A2(new_n12049_), .A3(new_n20321_), .ZN(new_n20322_));
  NOR2_X1    g17286(.A1(new_n20287_), .A2(pi0647), .ZN(new_n20323_));
  AOI21_X1   g17287(.A1(new_n20318_), .A2(pi0647), .B(new_n20323_), .ZN(new_n20324_));
  NAND2_X1   g17288(.A1(new_n20324_), .A2(new_n12088_), .ZN(new_n20325_));
  NAND2_X1   g17289(.A1(new_n20325_), .A2(pi0787), .ZN(new_n20326_));
  AOI21_X1   g17290(.A1(pi0630), .A2(new_n20322_), .B(new_n20326_), .ZN(new_n20327_));
  AOI22_X1   g17291(.A1(new_n20295_), .A2(new_n20316_), .B1(new_n20317_), .B2(new_n20327_), .ZN(new_n20328_));
  NOR2_X1    g17292(.A1(new_n20328_), .A2(new_n12082_), .ZN(new_n20329_));
  NAND4_X1   g17293(.A1(new_n20320_), .A2(pi0787), .A3(new_n12049_), .A4(new_n20321_), .ZN(new_n20330_));
  OAI21_X1   g17294(.A1(pi0787), .A2(new_n20319_), .B(new_n20330_), .ZN(new_n20331_));
  NOR2_X1    g17295(.A1(new_n20331_), .A2(pi0644), .ZN(new_n20332_));
  OR3_X2     g17296(.A1(new_n20329_), .A2(pi0715), .A3(new_n20332_), .Z(new_n20333_));
  MUX2_X1    g17297(.I0(new_n20303_), .I1(new_n20227_), .S(new_n16841_), .Z(new_n20334_));
  INV_X1     g17298(.I(new_n20334_), .ZN(new_n20335_));
  OAI21_X1   g17299(.A1(new_n20334_), .A2(new_n20227_), .B(new_n12082_), .ZN(new_n20336_));
  AOI21_X1   g17300(.A1(new_n20227_), .A2(new_n20334_), .B(new_n20336_), .ZN(new_n20337_));
  OAI21_X1   g17301(.A1(new_n20337_), .A2(new_n20335_), .B(new_n12099_), .ZN(new_n20338_));
  AOI21_X1   g17302(.A1(new_n20335_), .A2(new_n20337_), .B(new_n20338_), .ZN(new_n20339_));
  AOI21_X1   g17303(.A1(new_n20333_), .A2(new_n20339_), .B(pi1160), .ZN(new_n20340_));
  XOR2_X1    g17304(.A1(new_n20337_), .A2(new_n20227_), .Z(new_n20341_));
  AOI21_X1   g17305(.A1(new_n20331_), .A2(pi0644), .B(new_n13169_), .ZN(new_n20342_));
  OAI21_X1   g17306(.A1(new_n20341_), .A2(new_n12099_), .B(new_n20342_), .ZN(new_n20343_));
  OAI21_X1   g17307(.A1(new_n20329_), .A2(new_n20343_), .B(pi0790), .ZN(new_n20344_));
  NOR2_X1    g17308(.A1(new_n20328_), .A2(new_n14748_), .ZN(new_n20345_));
  OAI21_X1   g17309(.A1(new_n20340_), .A2(new_n20344_), .B(new_n20345_), .ZN(new_n20346_));
  NOR2_X1    g17310(.A1(new_n3231_), .A2(pi0186), .ZN(new_n20347_));
  INV_X1     g17311(.I(new_n20347_), .ZN(new_n20348_));
  NAND4_X1   g17312(.A1(new_n14351_), .A2(pi0186), .A3(new_n16089_), .A4(new_n14352_), .ZN(new_n20349_));
  NAND3_X1   g17313(.A1(new_n14347_), .A2(new_n20349_), .A3(new_n7109_), .ZN(new_n20350_));
  NAND3_X1   g17314(.A1(new_n14355_), .A2(new_n7109_), .A3(new_n12901_), .ZN(new_n20351_));
  NAND2_X1   g17315(.A1(new_n20351_), .A2(new_n16089_), .ZN(new_n20352_));
  NOR2_X1    g17316(.A1(new_n12694_), .A2(pi0038), .ZN(new_n20353_));
  NOR2_X1    g17317(.A1(new_n20353_), .A2(new_n7109_), .ZN(new_n20354_));
  INV_X1     g17318(.I(new_n14365_), .ZN(new_n20355_));
  NOR3_X1    g17319(.A1(new_n20355_), .A2(pi0186), .A3(pi0752), .ZN(new_n20356_));
  OAI21_X1   g17320(.A1(new_n20356_), .A2(new_n20354_), .B(new_n17798_), .ZN(new_n20357_));
  NAND4_X1   g17321(.A1(new_n20357_), .A2(new_n20352_), .A3(new_n20350_), .A4(new_n16094_), .ZN(new_n20358_));
  NAND2_X1   g17322(.A1(new_n20358_), .A2(new_n3231_), .ZN(new_n20359_));
  XOR2_X1    g17323(.A1(new_n20359_), .A2(new_n20348_), .Z(new_n20360_));
  NAND2_X1   g17324(.A1(new_n20360_), .A2(pi0625), .ZN(new_n20361_));
  NAND4_X1   g17325(.A1(new_n14355_), .A2(new_n7109_), .A3(pi0752), .A4(new_n12901_), .ZN(new_n20362_));
  NAND3_X1   g17326(.A1(new_n20357_), .A2(new_n20362_), .A3(new_n3231_), .ZN(new_n20363_));
  NAND2_X1   g17327(.A1(new_n20363_), .A2(new_n20348_), .ZN(new_n20364_));
  INV_X1     g17328(.I(new_n20364_), .ZN(new_n20365_));
  AOI21_X1   g17329(.A1(new_n20365_), .A2(new_n12970_), .B(pi1153), .ZN(new_n20366_));
  NAND2_X1   g17330(.A1(new_n20361_), .A2(new_n20366_), .ZN(new_n20367_));
  NOR3_X1    g17331(.A1(new_n13399_), .A2(pi0186), .A3(new_n13396_), .ZN(new_n20368_));
  INV_X1     g17332(.I(new_n20368_), .ZN(new_n20369_));
  AOI21_X1   g17333(.A1(new_n13399_), .A2(new_n7109_), .B(new_n13395_), .ZN(new_n20370_));
  NOR2_X1    g17334(.A1(new_n12828_), .A2(pi0186), .ZN(new_n20371_));
  NOR4_X1    g17335(.A1(new_n15189_), .A2(pi0038), .A3(pi0703), .A4(new_n20371_), .ZN(new_n20372_));
  INV_X1     g17336(.I(new_n20372_), .ZN(new_n20373_));
  NOR2_X1    g17337(.A1(new_n20370_), .A2(new_n20373_), .ZN(new_n20374_));
  AOI22_X1   g17338(.A1(new_n20374_), .A2(new_n20369_), .B1(new_n16094_), .B2(new_n20351_), .ZN(new_n20375_));
  NOR3_X1    g17339(.A1(new_n20375_), .A2(new_n3232_), .A3(new_n20348_), .ZN(new_n20376_));
  NOR2_X1    g17340(.A1(new_n20375_), .A2(new_n3232_), .ZN(new_n20377_));
  NOR2_X1    g17341(.A1(new_n20377_), .A2(new_n20347_), .ZN(new_n20378_));
  NOR2_X1    g17342(.A1(new_n20378_), .A2(new_n20376_), .ZN(new_n20379_));
  NAND2_X1   g17343(.A1(new_n20379_), .A2(pi0625), .ZN(new_n20380_));
  NOR2_X1    g17344(.A1(new_n12965_), .A2(pi0186), .ZN(new_n20381_));
  AOI21_X1   g17345(.A1(new_n20381_), .A2(pi0625), .B(pi1153), .ZN(new_n20382_));
  NAND3_X1   g17346(.A1(new_n20380_), .A2(pi0608), .A3(new_n20382_), .ZN(new_n20383_));
  INV_X1     g17347(.I(new_n20383_), .ZN(new_n20384_));
  INV_X1     g17348(.I(new_n20381_), .ZN(new_n20385_));
  AOI21_X1   g17349(.A1(new_n20385_), .A2(new_n12970_), .B(pi1153), .ZN(new_n20386_));
  AOI21_X1   g17350(.A1(new_n20364_), .A2(pi0625), .B(new_n12978_), .ZN(new_n20387_));
  INV_X1     g17351(.I(new_n20387_), .ZN(new_n20388_));
  AOI21_X1   g17352(.A1(new_n20380_), .A2(new_n20386_), .B(new_n20388_), .ZN(new_n20389_));
  AOI22_X1   g17353(.A1(new_n20367_), .A2(new_n20384_), .B1(new_n20361_), .B2(new_n20389_), .ZN(new_n20390_));
  MUX2_X1    g17354(.I0(new_n20390_), .I1(new_n20360_), .S(new_n11891_), .Z(new_n20391_));
  NAND2_X1   g17355(.A1(new_n20391_), .A2(new_n11870_), .ZN(new_n20392_));
  NAND2_X1   g17356(.A1(new_n20379_), .A2(new_n11891_), .ZN(new_n20393_));
  INV_X1     g17357(.I(new_n20393_), .ZN(new_n20394_));
  NAND4_X1   g17358(.A1(new_n20380_), .A2(new_n12970_), .A3(new_n11893_), .A4(new_n20385_), .ZN(new_n20395_));
  NAND3_X1   g17359(.A1(new_n20395_), .A2(pi0778), .A3(new_n20394_), .ZN(new_n20396_));
  INV_X1     g17360(.I(new_n20396_), .ZN(new_n20397_));
  AOI21_X1   g17361(.A1(new_n20395_), .A2(pi0778), .B(new_n20394_), .ZN(new_n20398_));
  OAI21_X1   g17362(.A1(new_n20397_), .A2(new_n20398_), .B(new_n11903_), .ZN(new_n20399_));
  NOR2_X1    g17363(.A1(new_n20381_), .A2(new_n12996_), .ZN(new_n20400_));
  NOR3_X1    g17364(.A1(new_n20364_), .A2(pi0609), .A3(new_n11914_), .ZN(new_n20401_));
  OAI21_X1   g17365(.A1(new_n20401_), .A2(new_n20400_), .B(new_n11912_), .ZN(new_n20402_));
  AOI21_X1   g17366(.A1(new_n20402_), .A2(pi0660), .B(new_n11903_), .ZN(new_n20403_));
  INV_X1     g17367(.I(new_n20403_), .ZN(new_n20404_));
  AOI21_X1   g17368(.A1(new_n20399_), .A2(pi1155), .B(new_n20404_), .ZN(new_n20405_));
  INV_X1     g17369(.I(new_n20361_), .ZN(new_n20406_));
  INV_X1     g17370(.I(new_n20366_), .ZN(new_n20407_));
  AOI21_X1   g17371(.A1(new_n20360_), .A2(pi0625), .B(new_n20407_), .ZN(new_n20408_));
  INV_X1     g17372(.I(new_n20389_), .ZN(new_n20409_));
  OAI22_X1   g17373(.A1(new_n20409_), .A2(new_n20406_), .B1(new_n20383_), .B2(new_n20408_), .ZN(new_n20410_));
  NAND3_X1   g17374(.A1(new_n20410_), .A2(pi0778), .A3(new_n20360_), .ZN(new_n20411_));
  INV_X1     g17375(.I(new_n20360_), .ZN(new_n20412_));
  OAI21_X1   g17376(.A1(new_n20410_), .A2(new_n11891_), .B(new_n20412_), .ZN(new_n20413_));
  NAND3_X1   g17377(.A1(new_n20413_), .A2(new_n20411_), .A3(new_n11903_), .ZN(new_n20414_));
  NAND2_X1   g17378(.A1(new_n20395_), .A2(pi0778), .ZN(new_n20415_));
  NAND2_X1   g17379(.A1(new_n20415_), .A2(new_n20393_), .ZN(new_n20416_));
  NAND2_X1   g17380(.A1(new_n20416_), .A2(new_n20396_), .ZN(new_n20417_));
  NOR2_X1    g17381(.A1(new_n20381_), .A2(new_n11915_), .ZN(new_n20418_));
  NOR3_X1    g17382(.A1(new_n20364_), .A2(new_n11903_), .A3(new_n11914_), .ZN(new_n20419_));
  NOR2_X1    g17383(.A1(new_n11923_), .A2(pi1155), .ZN(new_n20421_));
  INV_X1     g17384(.I(new_n20421_), .ZN(new_n20422_));
  AOI21_X1   g17385(.A1(new_n20417_), .A2(pi0609), .B(new_n20422_), .ZN(new_n20423_));
  AOI22_X1   g17386(.A1(new_n20414_), .A2(new_n20423_), .B1(new_n20405_), .B2(new_n20391_), .ZN(new_n20424_));
  NOR3_X1    g17387(.A1(new_n20424_), .A2(new_n11870_), .A3(new_n20392_), .ZN(new_n20425_));
  INV_X1     g17388(.I(new_n20392_), .ZN(new_n20426_));
  NAND2_X1   g17389(.A1(new_n20413_), .A2(new_n20411_), .ZN(new_n20427_));
  AOI21_X1   g17390(.A1(new_n20416_), .A2(new_n20396_), .B(pi0609), .ZN(new_n20428_));
  OAI21_X1   g17391(.A1(new_n20428_), .A2(new_n11912_), .B(new_n20403_), .ZN(new_n20429_));
  NOR3_X1    g17392(.A1(new_n20390_), .A2(new_n11891_), .A3(new_n20412_), .ZN(new_n20430_));
  AOI21_X1   g17393(.A1(new_n20390_), .A2(pi0778), .B(new_n20360_), .ZN(new_n20431_));
  NOR3_X1    g17394(.A1(new_n20430_), .A2(new_n20431_), .A3(pi0609), .ZN(new_n20432_));
  NOR2_X1    g17395(.A1(new_n20397_), .A2(new_n20398_), .ZN(new_n20433_));
  OAI21_X1   g17396(.A1(new_n20433_), .A2(new_n11903_), .B(new_n20421_), .ZN(new_n20434_));
  OAI22_X1   g17397(.A1(new_n20432_), .A2(new_n20434_), .B1(new_n20427_), .B2(new_n20429_), .ZN(new_n20435_));
  AOI21_X1   g17398(.A1(new_n20435_), .A2(pi0785), .B(new_n20426_), .ZN(new_n20436_));
  NOR3_X1    g17399(.A1(new_n20436_), .A2(new_n20425_), .A3(pi0781), .ZN(new_n20437_));
  INV_X1     g17400(.I(new_n20437_), .ZN(new_n20438_));
  NOR2_X1    g17401(.A1(new_n20436_), .A2(new_n20425_), .ZN(new_n20439_));
  NOR2_X1    g17402(.A1(new_n20385_), .A2(new_n11938_), .ZN(new_n20440_));
  AOI21_X1   g17403(.A1(new_n20417_), .A2(new_n11938_), .B(new_n20440_), .ZN(new_n20441_));
  OAI21_X1   g17404(.A1(new_n20441_), .A2(pi0618), .B(pi1154), .ZN(new_n20442_));
  NOR2_X1    g17405(.A1(new_n20365_), .A2(new_n11914_), .ZN(new_n20443_));
  NOR2_X1    g17406(.A1(new_n20385_), .A2(new_n11924_), .ZN(new_n20444_));
  NOR3_X1    g17407(.A1(new_n20443_), .A2(pi0785), .A3(new_n20444_), .ZN(new_n20445_));
  OAI21_X1   g17408(.A1(new_n20419_), .A2(new_n20418_), .B(pi1155), .ZN(new_n20446_));
  AOI21_X1   g17409(.A1(new_n20402_), .A2(new_n20446_), .B(new_n11870_), .ZN(new_n20447_));
  NAND2_X1   g17410(.A1(new_n20447_), .A2(new_n20445_), .ZN(new_n20448_));
  OR2_X2     g17411(.A1(new_n20447_), .A2(new_n20445_), .Z(new_n20449_));
  NAND3_X1   g17412(.A1(new_n20449_), .A2(pi0618), .A3(new_n20448_), .ZN(new_n20450_));
  NAND2_X1   g17413(.A1(new_n20381_), .A2(pi0618), .ZN(new_n20451_));
  NAND4_X1   g17414(.A1(new_n20450_), .A2(pi0627), .A3(new_n11950_), .A4(new_n20451_), .ZN(new_n20452_));
  AND3_X2    g17415(.A1(new_n20442_), .A2(pi0618), .A3(new_n20452_), .Z(new_n20453_));
  NAND3_X1   g17416(.A1(new_n20435_), .A2(new_n20426_), .A3(pi0785), .ZN(new_n20454_));
  OAI21_X1   g17417(.A1(new_n20424_), .A2(new_n11870_), .B(new_n20392_), .ZN(new_n20455_));
  NAND3_X1   g17418(.A1(new_n20454_), .A2(new_n20455_), .A3(new_n11934_), .ZN(new_n20456_));
  NOR2_X1    g17419(.A1(new_n20441_), .A2(new_n11934_), .ZN(new_n20457_));
  AOI21_X1   g17420(.A1(new_n20385_), .A2(new_n11934_), .B(pi1154), .ZN(new_n20458_));
  AOI21_X1   g17421(.A1(new_n20450_), .A2(new_n20458_), .B(pi0627), .ZN(new_n20459_));
  NOR3_X1    g17422(.A1(new_n20457_), .A2(pi1154), .A3(new_n20459_), .ZN(new_n20460_));
  AOI22_X1   g17423(.A1(new_n20456_), .A2(new_n20460_), .B1(new_n20439_), .B2(new_n20453_), .ZN(new_n20461_));
  NOR3_X1    g17424(.A1(new_n20461_), .A2(new_n11969_), .A3(new_n20438_), .ZN(new_n20462_));
  NAND3_X1   g17425(.A1(new_n20454_), .A2(new_n20453_), .A3(new_n20455_), .ZN(new_n20463_));
  NOR3_X1    g17426(.A1(new_n20436_), .A2(new_n20425_), .A3(pi0618), .ZN(new_n20464_));
  INV_X1     g17427(.I(new_n20460_), .ZN(new_n20465_));
  OAI21_X1   g17428(.A1(new_n20464_), .A2(new_n20465_), .B(new_n20463_), .ZN(new_n20466_));
  AOI21_X1   g17429(.A1(new_n20466_), .A2(pi0781), .B(new_n20437_), .ZN(new_n20467_));
  NOR3_X1    g17430(.A1(new_n20462_), .A2(new_n20467_), .A3(pi0789), .ZN(new_n20468_));
  NAND3_X1   g17431(.A1(new_n20466_), .A2(pi0781), .A3(new_n20437_), .ZN(new_n20469_));
  OAI21_X1   g17432(.A1(new_n20461_), .A2(new_n11969_), .B(new_n20438_), .ZN(new_n20470_));
  AND2_X2    g17433(.A1(new_n20449_), .A2(new_n20448_), .Z(new_n20471_));
  NAND3_X1   g17434(.A1(new_n20385_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n20472_));
  MUX2_X1    g17435(.I0(new_n20472_), .I1(new_n20471_), .S(new_n11969_), .Z(new_n20473_));
  OAI21_X1   g17436(.A1(new_n20385_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n20474_));
  AOI21_X1   g17437(.A1(new_n20473_), .A2(pi0619), .B(new_n20474_), .ZN(new_n20475_));
  NOR2_X1    g17438(.A1(new_n20381_), .A2(new_n11961_), .ZN(new_n20476_));
  AOI21_X1   g17439(.A1(new_n20441_), .A2(new_n11961_), .B(new_n20476_), .ZN(new_n20477_));
  NAND2_X1   g17440(.A1(new_n11869_), .A2(pi0619), .ZN(new_n20478_));
  AOI21_X1   g17441(.A1(new_n20475_), .A2(pi0648), .B(new_n20478_), .ZN(new_n20479_));
  NAND3_X1   g17442(.A1(new_n20470_), .A2(new_n20469_), .A3(new_n20479_), .ZN(new_n20480_));
  NOR3_X1    g17443(.A1(new_n20462_), .A2(new_n20467_), .A3(pi0619), .ZN(new_n20481_));
  NAND2_X1   g17444(.A1(new_n20473_), .A2(pi0619), .ZN(new_n20482_));
  AOI21_X1   g17445(.A1(new_n20385_), .A2(new_n11967_), .B(pi1159), .ZN(new_n20483_));
  NAND2_X1   g17446(.A1(new_n20482_), .A2(new_n20483_), .ZN(new_n20484_));
  NAND2_X1   g17447(.A1(new_n20484_), .A2(new_n11966_), .ZN(new_n20485_));
  NAND2_X1   g17448(.A1(new_n20477_), .A2(pi0619), .ZN(new_n20486_));
  NAND3_X1   g17449(.A1(new_n20485_), .A2(new_n11869_), .A3(new_n20486_), .ZN(new_n20487_));
  OAI21_X1   g17450(.A1(new_n20481_), .A2(new_n20487_), .B(new_n20480_), .ZN(new_n20488_));
  NAND3_X1   g17451(.A1(new_n20488_), .A2(pi0789), .A3(new_n20468_), .ZN(new_n20489_));
  INV_X1     g17452(.I(new_n20468_), .ZN(new_n20490_));
  NOR2_X1    g17453(.A1(new_n20462_), .A2(new_n20467_), .ZN(new_n20491_));
  NAND3_X1   g17454(.A1(new_n20470_), .A2(new_n20469_), .A3(new_n11967_), .ZN(new_n20492_));
  INV_X1     g17455(.I(new_n20487_), .ZN(new_n20493_));
  AOI22_X1   g17456(.A1(new_n20492_), .A2(new_n20493_), .B1(new_n20491_), .B2(new_n20479_), .ZN(new_n20494_));
  OAI21_X1   g17457(.A1(new_n20494_), .A2(new_n11985_), .B(new_n20490_), .ZN(new_n20495_));
  NAND2_X1   g17458(.A1(new_n20495_), .A2(new_n20489_), .ZN(new_n20496_));
  NOR3_X1    g17459(.A1(new_n20494_), .A2(new_n11985_), .A3(new_n20490_), .ZN(new_n20497_));
  AOI21_X1   g17460(.A1(new_n20488_), .A2(pi0789), .B(new_n20468_), .ZN(new_n20498_));
  NAND2_X1   g17461(.A1(new_n20473_), .A2(new_n11985_), .ZN(new_n20499_));
  AOI21_X1   g17462(.A1(new_n20484_), .A2(new_n20475_), .B(new_n11985_), .ZN(new_n20500_));
  XNOR2_X1   g17463(.A1(new_n20500_), .A2(new_n20499_), .ZN(new_n20501_));
  NOR3_X1    g17464(.A1(new_n11994_), .A2(new_n11989_), .A3(pi1158), .ZN(new_n20502_));
  NAND2_X1   g17465(.A1(new_n20501_), .A2(new_n20502_), .ZN(new_n20503_));
  NOR2_X1    g17466(.A1(new_n20385_), .A2(new_n12014_), .ZN(new_n20504_));
  AOI21_X1   g17467(.A1(new_n20477_), .A2(new_n12014_), .B(new_n20504_), .ZN(new_n20505_));
  NOR2_X1    g17468(.A1(new_n11994_), .A2(pi0641), .ZN(new_n20506_));
  NAND2_X1   g17469(.A1(new_n20503_), .A2(new_n20506_), .ZN(new_n20507_));
  INV_X1     g17470(.I(new_n20507_), .ZN(new_n20508_));
  INV_X1     g17471(.I(new_n20501_), .ZN(new_n20509_));
  NOR2_X1    g17472(.A1(new_n20509_), .A2(pi0626), .ZN(new_n20510_));
  OAI21_X1   g17473(.A1(new_n20381_), .A2(new_n11994_), .B(pi0641), .ZN(new_n20511_));
  NOR3_X1    g17474(.A1(new_n11989_), .A2(pi0626), .A3(pi1158), .ZN(new_n20512_));
  OAI21_X1   g17475(.A1(new_n20510_), .A2(new_n20511_), .B(new_n20512_), .ZN(new_n20513_));
  INV_X1     g17476(.I(new_n20513_), .ZN(new_n20514_));
  OAI22_X1   g17477(.A1(new_n20497_), .A2(new_n20498_), .B1(new_n20508_), .B2(new_n20514_), .ZN(new_n20515_));
  NOR3_X1    g17478(.A1(new_n20515_), .A2(new_n11986_), .A3(new_n20496_), .ZN(new_n20516_));
  NOR2_X1    g17479(.A1(new_n20497_), .A2(new_n20498_), .ZN(new_n20517_));
  AOI21_X1   g17480(.A1(new_n20515_), .A2(pi0788), .B(new_n20517_), .ZN(new_n20518_));
  NOR2_X1    g17481(.A1(new_n20516_), .A2(new_n20518_), .ZN(new_n20519_));
  NAND2_X1   g17482(.A1(new_n20385_), .A2(new_n11997_), .ZN(new_n20520_));
  OAI21_X1   g17483(.A1(new_n20509_), .A2(new_n11997_), .B(new_n20520_), .ZN(new_n20521_));
  NOR2_X1    g17484(.A1(new_n20521_), .A2(pi0628), .ZN(new_n20522_));
  NOR2_X1    g17485(.A1(new_n20381_), .A2(new_n13114_), .ZN(new_n20523_));
  AOI21_X1   g17486(.A1(new_n20505_), .A2(new_n13114_), .B(new_n20523_), .ZN(new_n20524_));
  NOR3_X1    g17487(.A1(new_n20385_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n20525_));
  OAI21_X1   g17488(.A1(new_n20525_), .A2(new_n12030_), .B(pi0628), .ZN(new_n20526_));
  INV_X1     g17489(.I(new_n20526_), .ZN(new_n20527_));
  OAI21_X1   g17490(.A1(new_n20522_), .A2(new_n12026_), .B(new_n20527_), .ZN(new_n20528_));
  INV_X1     g17491(.I(new_n20528_), .ZN(new_n20529_));
  NOR2_X1    g17492(.A1(new_n20521_), .A2(new_n12031_), .ZN(new_n20530_));
  NOR2_X1    g17493(.A1(new_n12030_), .A2(pi0628), .ZN(new_n20531_));
  OAI21_X1   g17494(.A1(new_n20530_), .A2(pi1156), .B(new_n20531_), .ZN(new_n20532_));
  INV_X1     g17495(.I(new_n20532_), .ZN(new_n20533_));
  OAI22_X1   g17496(.A1(new_n20516_), .A2(new_n20518_), .B1(new_n20529_), .B2(new_n20533_), .ZN(new_n20534_));
  MUX2_X1    g17497(.I0(new_n20534_), .I1(new_n20519_), .S(new_n11868_), .Z(new_n20535_));
  AOI22_X1   g17498(.A1(new_n20495_), .A2(new_n20489_), .B1(new_n20507_), .B2(new_n20513_), .ZN(new_n20536_));
  NAND3_X1   g17499(.A1(new_n20536_), .A2(pi0788), .A3(new_n20517_), .ZN(new_n20537_));
  OAI21_X1   g17500(.A1(new_n20536_), .A2(new_n11986_), .B(new_n20496_), .ZN(new_n20538_));
  AOI21_X1   g17501(.A1(new_n20538_), .A2(new_n20537_), .B(new_n20528_), .ZN(new_n20539_));
  NAND3_X1   g17502(.A1(new_n20539_), .A2(new_n20519_), .A3(pi0792), .ZN(new_n20540_));
  NAND2_X1   g17503(.A1(new_n20538_), .A2(new_n20537_), .ZN(new_n20541_));
  AOI22_X1   g17504(.A1(new_n20538_), .A2(new_n20537_), .B1(new_n20528_), .B2(new_n20532_), .ZN(new_n20542_));
  OAI21_X1   g17505(.A1(new_n20542_), .A2(new_n11868_), .B(new_n20541_), .ZN(new_n20543_));
  NAND2_X1   g17506(.A1(new_n20543_), .A2(new_n20540_), .ZN(new_n20544_));
  NOR4_X1    g17507(.A1(new_n20524_), .A2(new_n12031_), .A3(pi1156), .A4(new_n20381_), .ZN(new_n20545_));
  NOR2_X1    g17508(.A1(new_n20545_), .A2(new_n20525_), .ZN(new_n20546_));
  MUX2_X1    g17509(.I0(new_n20546_), .I1(new_n20524_), .S(new_n11868_), .Z(new_n20547_));
  NAND2_X1   g17510(.A1(new_n20547_), .A2(pi0647), .ZN(new_n20548_));
  AOI21_X1   g17511(.A1(new_n20381_), .A2(pi0647), .B(pi1157), .ZN(new_n20549_));
  NAND2_X1   g17512(.A1(new_n20548_), .A2(new_n20549_), .ZN(new_n20550_));
  NOR2_X1    g17513(.A1(new_n20381_), .A2(new_n12054_), .ZN(new_n20551_));
  AOI21_X1   g17514(.A1(new_n20521_), .A2(new_n12054_), .B(new_n20551_), .ZN(new_n20552_));
  NOR2_X1    g17515(.A1(new_n12061_), .A2(pi1157), .ZN(new_n20553_));
  OAI21_X1   g17516(.A1(new_n20550_), .A2(new_n12060_), .B(new_n20553_), .ZN(new_n20554_));
  NOR3_X1    g17517(.A1(new_n20534_), .A2(new_n11868_), .A3(new_n20541_), .ZN(new_n20555_));
  AOI21_X1   g17518(.A1(new_n20534_), .A2(pi0792), .B(new_n20519_), .ZN(new_n20556_));
  NOR3_X1    g17519(.A1(new_n20555_), .A2(new_n20556_), .A3(pi0647), .ZN(new_n20557_));
  AOI21_X1   g17520(.A1(new_n20385_), .A2(new_n12061_), .B(pi1157), .ZN(new_n20558_));
  NAND2_X1   g17521(.A1(new_n20548_), .A2(new_n20558_), .ZN(new_n20559_));
  NAND2_X1   g17522(.A1(new_n20559_), .A2(new_n12060_), .ZN(new_n20560_));
  AOI21_X1   g17523(.A1(new_n20552_), .A2(pi0647), .B(pi1157), .ZN(new_n20561_));
  AND2_X2    g17524(.A1(new_n20561_), .A2(new_n20560_), .Z(new_n20562_));
  INV_X1     g17525(.I(new_n20562_), .ZN(new_n20563_));
  OAI22_X1   g17526(.A1(new_n20557_), .A2(new_n20563_), .B1(new_n20544_), .B2(new_n20554_), .ZN(new_n20564_));
  MUX2_X1    g17527(.I0(new_n20564_), .I1(new_n20535_), .S(new_n12048_), .Z(new_n20565_));
  NAND2_X1   g17528(.A1(new_n20547_), .A2(new_n12048_), .ZN(new_n20566_));
  INV_X1     g17529(.I(new_n20559_), .ZN(new_n20567_));
  OAI21_X1   g17530(.A1(new_n20567_), .A2(new_n20550_), .B(pi0787), .ZN(new_n20568_));
  XOR2_X1    g17531(.A1(new_n20568_), .A2(new_n20566_), .Z(new_n20569_));
  NOR2_X1    g17532(.A1(new_n20385_), .A2(new_n12092_), .ZN(new_n20570_));
  AOI21_X1   g17533(.A1(new_n20552_), .A2(new_n12092_), .B(new_n20570_), .ZN(new_n20571_));
  INV_X1     g17534(.I(new_n20571_), .ZN(new_n20572_));
  NOR2_X1    g17535(.A1(pi0644), .A2(pi0715), .ZN(new_n20573_));
  AOI21_X1   g17536(.A1(new_n20572_), .A2(new_n20573_), .B(new_n13169_), .ZN(new_n20574_));
  OAI21_X1   g17537(.A1(new_n20569_), .A2(new_n12082_), .B(new_n20574_), .ZN(new_n20575_));
  AOI21_X1   g17538(.A1(new_n20565_), .A2(new_n12082_), .B(new_n20575_), .ZN(new_n20576_));
  INV_X1     g17539(.I(new_n20554_), .ZN(new_n20577_));
  NAND3_X1   g17540(.A1(new_n20543_), .A2(new_n20540_), .A3(new_n12061_), .ZN(new_n20578_));
  AOI22_X1   g17541(.A1(new_n20578_), .A2(new_n20562_), .B1(new_n20535_), .B2(new_n20577_), .ZN(new_n20579_));
  MUX2_X1    g17542(.I0(new_n20579_), .I1(new_n20544_), .S(new_n12048_), .Z(new_n20580_));
  INV_X1     g17543(.I(new_n20569_), .ZN(new_n20581_));
  NAND3_X1   g17544(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n20582_));
  OAI21_X1   g17545(.A1(new_n20571_), .A2(new_n20582_), .B(new_n13179_), .ZN(new_n20583_));
  NOR2_X1    g17546(.A1(new_n20581_), .A2(new_n20583_), .ZN(new_n20584_));
  OAI21_X1   g17547(.A1(new_n20580_), .A2(new_n12082_), .B(new_n20584_), .ZN(new_n20585_));
  NOR2_X1    g17548(.A1(new_n20576_), .A2(new_n20585_), .ZN(new_n20586_));
  NAND2_X1   g17549(.A1(po1038), .A2(new_n7109_), .ZN(new_n20587_));
  AOI21_X1   g17550(.A1(new_n20587_), .A2(new_n13184_), .B(po1038), .ZN(new_n20588_));
  OAI21_X1   g17551(.A1(new_n20565_), .A2(pi0790), .B(new_n20588_), .ZN(new_n20589_));
  OAI21_X1   g17552(.A1(new_n20586_), .A2(new_n20589_), .B(new_n20346_), .ZN(po0343));
  NOR2_X1    g17553(.A1(new_n2925_), .A2(pi0187), .ZN(new_n20591_));
  NOR2_X1    g17554(.A1(new_n11877_), .A2(pi0770), .ZN(new_n20592_));
  NOR2_X1    g17555(.A1(new_n20592_), .A2(new_n20591_), .ZN(new_n20593_));
  INV_X1     g17556(.I(new_n20593_), .ZN(new_n20594_));
  AOI21_X1   g17557(.A1(new_n11886_), .A2(pi0726), .B(new_n20591_), .ZN(new_n20595_));
  NOR2_X1    g17558(.A1(new_n20595_), .A2(new_n11874_), .ZN(new_n20596_));
  NOR2_X1    g17559(.A1(new_n20594_), .A2(new_n20596_), .ZN(new_n20597_));
  NOR2_X1    g17560(.A1(new_n20597_), .A2(pi0778), .ZN(new_n20598_));
  NAND2_X1   g17561(.A1(new_n20596_), .A2(pi0625), .ZN(new_n20599_));
  NOR2_X1    g17562(.A1(new_n13201_), .A2(new_n15463_), .ZN(new_n20600_));
  NOR4_X1    g17563(.A1(new_n20592_), .A2(pi0608), .A3(new_n11893_), .A4(new_n20591_), .ZN(new_n20601_));
  OAI21_X1   g17564(.A1(new_n20594_), .A2(new_n20596_), .B(new_n20599_), .ZN(new_n20602_));
  NOR3_X1    g17565(.A1(new_n20591_), .A2(pi0608), .A3(pi1153), .ZN(new_n20603_));
  AOI22_X1   g17566(.A1(new_n20602_), .A2(new_n20603_), .B1(new_n20599_), .B2(new_n20601_), .ZN(new_n20604_));
  NOR2_X1    g17567(.A1(new_n20604_), .A2(new_n11891_), .ZN(new_n20605_));
  XOR2_X1    g17568(.A1(new_n20605_), .A2(new_n20598_), .Z(new_n20606_));
  INV_X1     g17569(.I(new_n20606_), .ZN(new_n20607_));
  NAND2_X1   g17570(.A1(new_n20607_), .A2(new_n11870_), .ZN(new_n20608_));
  AOI21_X1   g17571(.A1(new_n20606_), .A2(new_n11903_), .B(pi1155), .ZN(new_n20609_));
  INV_X1     g17572(.I(new_n20595_), .ZN(new_n20610_));
  XOR2_X1    g17573(.A1(new_n20600_), .A2(pi1153), .Z(new_n20611_));
  NAND2_X1   g17574(.A1(new_n20611_), .A2(new_n20610_), .ZN(new_n20612_));
  OAI21_X1   g17575(.A1(new_n20600_), .A2(new_n20591_), .B(new_n11893_), .ZN(new_n20613_));
  AOI21_X1   g17576(.A1(new_n20612_), .A2(new_n20613_), .B(new_n11891_), .ZN(new_n20614_));
  NOR2_X1    g17577(.A1(new_n20595_), .A2(pi0778), .ZN(new_n20615_));
  OAI21_X1   g17578(.A1(new_n20614_), .A2(new_n20615_), .B(pi0609), .ZN(new_n20616_));
  AOI21_X1   g17579(.A1(new_n20594_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n20617_));
  NOR2_X1    g17580(.A1(new_n20617_), .A2(pi0660), .ZN(new_n20618_));
  OAI21_X1   g17581(.A1(new_n20609_), .A2(new_n20616_), .B(new_n20618_), .ZN(new_n20619_));
  NOR2_X1    g17582(.A1(new_n20614_), .A2(new_n20615_), .ZN(new_n20620_));
  NAND4_X1   g17583(.A1(new_n20607_), .A2(pi0609), .A3(new_n11912_), .A4(new_n20620_), .ZN(new_n20621_));
  NOR2_X1    g17584(.A1(new_n20593_), .A2(new_n11925_), .ZN(new_n20622_));
  AOI21_X1   g17585(.A1(new_n20622_), .A2(new_n11928_), .B(pi1155), .ZN(new_n20623_));
  NOR2_X1    g17586(.A1(new_n20623_), .A2(new_n11923_), .ZN(new_n20624_));
  NAND2_X1   g17587(.A1(new_n20621_), .A2(new_n20624_), .ZN(new_n20625_));
  NAND3_X1   g17588(.A1(new_n20625_), .A2(pi0785), .A3(new_n20619_), .ZN(new_n20626_));
  NAND2_X1   g17589(.A1(new_n20626_), .A2(new_n20608_), .ZN(new_n20627_));
  NOR4_X1    g17590(.A1(new_n20620_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n20629_));
  NOR2_X1    g17591(.A1(new_n20622_), .A2(pi0785), .ZN(new_n20630_));
  OAI21_X1   g17592(.A1(new_n20623_), .A2(new_n20617_), .B(pi0785), .ZN(new_n20631_));
  XNOR2_X1   g17593(.A1(new_n20631_), .A2(new_n20630_), .ZN(new_n20632_));
  INV_X1     g17594(.I(new_n20632_), .ZN(new_n20633_));
  NOR2_X1    g17595(.A1(new_n20633_), .A2(new_n11945_), .ZN(new_n20634_));
  NOR3_X1    g17596(.A1(new_n20629_), .A2(new_n20634_), .A3(pi0627), .ZN(new_n20635_));
  AOI21_X1   g17597(.A1(new_n20632_), .A2(new_n11951_), .B(pi1154), .ZN(new_n20636_));
  NOR2_X1    g17598(.A1(new_n20620_), .A2(new_n11939_), .ZN(new_n20637_));
  INV_X1     g17599(.I(new_n20637_), .ZN(new_n20638_));
  NAND4_X1   g17600(.A1(new_n20627_), .A2(pi0618), .A3(new_n11950_), .A4(new_n20638_), .ZN(new_n20639_));
  NAND2_X1   g17601(.A1(new_n20639_), .A2(new_n20636_), .ZN(new_n20640_));
  AOI21_X1   g17602(.A1(new_n20640_), .A2(new_n11949_), .B(new_n20635_), .ZN(new_n20641_));
  NOR2_X1    g17603(.A1(new_n20641_), .A2(new_n11969_), .ZN(new_n20642_));
  AOI21_X1   g17604(.A1(new_n11969_), .A2(new_n20627_), .B(new_n20642_), .ZN(new_n20643_));
  NOR2_X1    g17605(.A1(new_n20638_), .A2(new_n11962_), .ZN(new_n20644_));
  NOR4_X1    g17606(.A1(new_n20643_), .A2(new_n11967_), .A3(pi1159), .A4(new_n20644_), .ZN(new_n20645_));
  INV_X1     g17607(.I(new_n20634_), .ZN(new_n20646_));
  NAND2_X1   g17608(.A1(new_n20646_), .A2(new_n20636_), .ZN(new_n20647_));
  MUX2_X1    g17609(.I0(new_n20647_), .I1(new_n20632_), .S(new_n11969_), .Z(new_n20648_));
  NAND2_X1   g17610(.A1(new_n20648_), .A2(pi0619), .ZN(new_n20649_));
  INV_X1     g17611(.I(new_n20649_), .ZN(new_n20650_));
  INV_X1     g17612(.I(new_n20591_), .ZN(new_n20651_));
  OAI21_X1   g17613(.A1(new_n20651_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n20652_));
  NOR4_X1    g17614(.A1(new_n20645_), .A2(new_n11966_), .A3(new_n20650_), .A4(new_n20652_), .ZN(new_n20653_));
  NOR4_X1    g17615(.A1(new_n20638_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n20654_));
  OAI21_X1   g17616(.A1(new_n20591_), .A2(pi0619), .B(new_n11869_), .ZN(new_n20655_));
  OAI21_X1   g17617(.A1(new_n20650_), .A2(new_n20655_), .B(new_n11966_), .ZN(new_n20656_));
  NOR2_X1    g17618(.A1(new_n20656_), .A2(new_n20654_), .ZN(new_n20657_));
  AOI21_X1   g17619(.A1(new_n20643_), .A2(new_n11998_), .B(pi0789), .ZN(new_n20658_));
  OAI21_X1   g17620(.A1(new_n20653_), .A2(new_n20657_), .B(new_n20658_), .ZN(new_n20659_));
  NAND2_X1   g17621(.A1(new_n20644_), .A2(new_n17450_), .ZN(new_n20660_));
  NOR2_X1    g17622(.A1(new_n20660_), .A2(new_n17153_), .ZN(new_n20661_));
  INV_X1     g17623(.I(new_n20661_), .ZN(new_n20662_));
  NOR2_X1    g17624(.A1(new_n20662_), .A2(new_n17151_), .ZN(new_n20663_));
  NOR2_X1    g17625(.A1(new_n14624_), .A2(new_n20591_), .ZN(new_n20664_));
  NAND3_X1   g17626(.A1(new_n20651_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n20665_));
  MUX2_X1    g17627(.I0(new_n20665_), .I1(new_n20648_), .S(new_n11985_), .Z(new_n20666_));
  AOI21_X1   g17628(.A1(new_n20666_), .A2(new_n14624_), .B(new_n20664_), .ZN(new_n20667_));
  AND2_X2    g17629(.A1(new_n20667_), .A2(new_n12064_), .Z(new_n20668_));
  OAI21_X1   g17630(.A1(new_n20668_), .A2(new_n20663_), .B(pi0629), .ZN(new_n20669_));
  NAND2_X1   g17631(.A1(new_n20667_), .A2(new_n12063_), .ZN(new_n20670_));
  NAND2_X1   g17632(.A1(new_n20661_), .A2(new_n15084_), .ZN(new_n20671_));
  NAND4_X1   g17633(.A1(new_n20669_), .A2(new_n15085_), .A3(new_n20670_), .A4(new_n20671_), .ZN(new_n20672_));
  MUX2_X1    g17634(.I0(new_n20666_), .I1(new_n20651_), .S(new_n11994_), .Z(new_n20673_));
  NOR2_X1    g17635(.A1(new_n20673_), .A2(new_n17167_), .ZN(new_n20674_));
  OAI21_X1   g17636(.A1(new_n20666_), .A2(new_n20591_), .B(pi0626), .ZN(new_n20675_));
  NOR2_X1    g17637(.A1(new_n20660_), .A2(new_n12020_), .ZN(new_n20676_));
  NOR2_X1    g17638(.A1(new_n20676_), .A2(pi0788), .ZN(new_n20677_));
  OAI21_X1   g17639(.A1(new_n20675_), .A2(new_n17171_), .B(new_n20677_), .ZN(new_n20678_));
  OAI21_X1   g17640(.A1(new_n20674_), .A2(new_n20678_), .B(new_n14732_), .ZN(new_n20679_));
  AOI21_X1   g17641(.A1(new_n20672_), .A2(new_n14726_), .B(new_n20679_), .ZN(new_n20680_));
  NAND3_X1   g17642(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n20591_), .ZN(new_n20681_));
  NOR2_X1    g17643(.A1(new_n20662_), .A2(new_n12068_), .ZN(new_n20682_));
  INV_X1     g17644(.I(new_n20682_), .ZN(new_n20683_));
  NAND2_X1   g17645(.A1(new_n20683_), .A2(pi0647), .ZN(new_n20684_));
  NAND2_X1   g17646(.A1(new_n20591_), .A2(pi0647), .ZN(new_n20685_));
  NAND3_X1   g17647(.A1(new_n20684_), .A2(new_n12049_), .A3(new_n20685_), .ZN(new_n20686_));
  NOR2_X1    g17648(.A1(new_n20651_), .A2(pi0647), .ZN(new_n20687_));
  AOI21_X1   g17649(.A1(new_n20682_), .A2(pi0647), .B(new_n20687_), .ZN(new_n20688_));
  NAND2_X1   g17650(.A1(new_n20688_), .A2(new_n12088_), .ZN(new_n20689_));
  NAND2_X1   g17651(.A1(new_n20689_), .A2(pi0787), .ZN(new_n20690_));
  AOI21_X1   g17652(.A1(pi0630), .A2(new_n20686_), .B(new_n20690_), .ZN(new_n20691_));
  AOI22_X1   g17653(.A1(new_n20659_), .A2(new_n20680_), .B1(new_n20681_), .B2(new_n20691_), .ZN(new_n20692_));
  NOR2_X1    g17654(.A1(new_n20692_), .A2(new_n12082_), .ZN(new_n20693_));
  NAND4_X1   g17655(.A1(new_n20684_), .A2(pi0787), .A3(new_n12049_), .A4(new_n20685_), .ZN(new_n20694_));
  OAI21_X1   g17656(.A1(pi0787), .A2(new_n20683_), .B(new_n20694_), .ZN(new_n20695_));
  NOR2_X1    g17657(.A1(new_n20695_), .A2(pi0644), .ZN(new_n20696_));
  OR3_X2     g17658(.A1(new_n20693_), .A2(pi0715), .A3(new_n20696_), .Z(new_n20697_));
  MUX2_X1    g17659(.I0(new_n20667_), .I1(new_n20591_), .S(new_n16841_), .Z(new_n20698_));
  INV_X1     g17660(.I(new_n20698_), .ZN(new_n20699_));
  OAI21_X1   g17661(.A1(new_n20698_), .A2(new_n20591_), .B(new_n12082_), .ZN(new_n20700_));
  AOI21_X1   g17662(.A1(new_n20591_), .A2(new_n20698_), .B(new_n20700_), .ZN(new_n20701_));
  OAI21_X1   g17663(.A1(new_n20701_), .A2(new_n20699_), .B(new_n12099_), .ZN(new_n20702_));
  AOI21_X1   g17664(.A1(new_n20699_), .A2(new_n20701_), .B(new_n20702_), .ZN(new_n20703_));
  AOI21_X1   g17665(.A1(new_n20697_), .A2(new_n20703_), .B(pi1160), .ZN(new_n20704_));
  XOR2_X1    g17666(.A1(new_n20701_), .A2(new_n20591_), .Z(new_n20705_));
  AOI21_X1   g17667(.A1(new_n20695_), .A2(pi0644), .B(new_n13169_), .ZN(new_n20706_));
  OAI21_X1   g17668(.A1(new_n20705_), .A2(new_n12099_), .B(new_n20706_), .ZN(new_n20707_));
  OAI21_X1   g17669(.A1(new_n20693_), .A2(new_n20707_), .B(pi0790), .ZN(new_n20708_));
  NOR2_X1    g17670(.A1(new_n20692_), .A2(new_n14748_), .ZN(new_n20709_));
  OAI21_X1   g17671(.A1(new_n20704_), .A2(new_n20708_), .B(new_n20709_), .ZN(new_n20710_));
  NOR2_X1    g17672(.A1(new_n3231_), .A2(pi0187), .ZN(new_n20711_));
  NOR2_X1    g17673(.A1(pi0187), .A2(pi0726), .ZN(new_n20712_));
  OAI21_X1   g17674(.A1(new_n14363_), .A2(new_n8861_), .B(new_n17798_), .ZN(new_n20713_));
  NAND2_X1   g17675(.A1(new_n12901_), .A2(new_n15427_), .ZN(new_n20714_));
  OAI22_X1   g17676(.A1(new_n14355_), .A2(new_n20714_), .B1(pi0770), .B2(new_n14365_), .ZN(new_n20715_));
  AOI22_X1   g17677(.A1(new_n20715_), .A2(new_n8861_), .B1(new_n15427_), .B2(new_n20713_), .ZN(new_n20716_));
  AOI22_X1   g17678(.A1(new_n20716_), .A2(new_n15463_), .B1(new_n14347_), .B2(new_n20712_), .ZN(new_n20717_));
  NOR2_X1    g17679(.A1(new_n20717_), .A2(new_n3232_), .ZN(new_n20718_));
  XOR2_X1    g17680(.A1(new_n20718_), .A2(new_n20711_), .Z(new_n20719_));
  AOI21_X1   g17681(.A1(new_n20716_), .A2(new_n3231_), .B(new_n20711_), .ZN(new_n20720_));
  OAI21_X1   g17682(.A1(new_n20720_), .A2(pi0625), .B(pi1153), .ZN(new_n20721_));
  INV_X1     g17683(.I(new_n13900_), .ZN(new_n20722_));
  NOR2_X1    g17684(.A1(new_n20722_), .A2(pi1153), .ZN(new_n20723_));
  NAND2_X1   g17685(.A1(new_n8861_), .A2(new_n15463_), .ZN(new_n20724_));
  OAI21_X1   g17686(.A1(new_n12902_), .A2(new_n20724_), .B(new_n3231_), .ZN(new_n20725_));
  NOR3_X1    g17687(.A1(new_n13399_), .A2(pi0187), .A3(new_n13396_), .ZN(new_n20726_));
  AOI21_X1   g17688(.A1(new_n13399_), .A2(new_n8861_), .B(new_n13395_), .ZN(new_n20727_));
  NAND2_X1   g17689(.A1(new_n13368_), .A2(new_n8861_), .ZN(new_n20728_));
  NAND4_X1   g17690(.A1(new_n20728_), .A2(new_n3172_), .A3(new_n15463_), .A4(new_n13403_), .ZN(new_n20729_));
  NOR3_X1    g17691(.A1(new_n20726_), .A2(new_n20727_), .A3(new_n20729_), .ZN(new_n20730_));
  AOI22_X1   g17692(.A1(new_n20730_), .A2(new_n20725_), .B1(pi0187), .B2(new_n3232_), .ZN(new_n20731_));
  INV_X1     g17693(.I(new_n20731_), .ZN(new_n20732_));
  NOR2_X1    g17694(.A1(new_n12965_), .A2(pi0187), .ZN(new_n20733_));
  AOI21_X1   g17695(.A1(new_n20732_), .A2(new_n20723_), .B(new_n12970_), .ZN(new_n20734_));
  NAND2_X1   g17696(.A1(new_n20734_), .A2(new_n20721_), .ZN(new_n20735_));
  NOR2_X1    g17697(.A1(new_n20720_), .A2(new_n12970_), .ZN(new_n20736_));
  NOR2_X1    g17698(.A1(pi0608), .A2(pi0625), .ZN(new_n20738_));
  OAI21_X1   g17699(.A1(new_n20736_), .A2(pi1153), .B(new_n20738_), .ZN(new_n20739_));
  AOI21_X1   g17700(.A1(new_n20735_), .A2(new_n20739_), .B(new_n20719_), .ZN(new_n20740_));
  NAND3_X1   g17701(.A1(new_n20740_), .A2(pi0778), .A3(new_n20719_), .ZN(new_n20741_));
  INV_X1     g17702(.I(new_n20719_), .ZN(new_n20742_));
  OAI21_X1   g17703(.A1(new_n20740_), .A2(new_n11891_), .B(new_n20742_), .ZN(new_n20743_));
  NAND2_X1   g17704(.A1(new_n20743_), .A2(new_n20741_), .ZN(new_n20744_));
  NOR2_X1    g17705(.A1(new_n20744_), .A2(pi0785), .ZN(new_n20745_));
  INV_X1     g17706(.I(new_n20745_), .ZN(new_n20746_));
  INV_X1     g17707(.I(new_n20744_), .ZN(new_n20747_));
  NOR2_X1    g17708(.A1(new_n20731_), .A2(pi0778), .ZN(new_n20748_));
  INV_X1     g17709(.I(new_n20733_), .ZN(new_n20749_));
  MUX2_X1    g17710(.I0(new_n20749_), .I1(new_n20731_), .S(new_n13435_), .Z(new_n20750_));
  NOR2_X1    g17711(.A1(new_n20750_), .A2(new_n11891_), .ZN(new_n20751_));
  NOR2_X1    g17712(.A1(new_n20751_), .A2(new_n20748_), .ZN(new_n20752_));
  INV_X1     g17713(.I(new_n20752_), .ZN(new_n20753_));
  AOI21_X1   g17714(.A1(new_n20753_), .A2(new_n11903_), .B(new_n11912_), .ZN(new_n20754_));
  NOR2_X1    g17715(.A1(new_n20733_), .A2(new_n12996_), .ZN(new_n20755_));
  INV_X1     g17716(.I(new_n20755_), .ZN(new_n20756_));
  NAND3_X1   g17717(.A1(new_n20720_), .A2(new_n11903_), .A3(new_n11924_), .ZN(new_n20757_));
  AOI21_X1   g17718(.A1(new_n20757_), .A2(new_n20756_), .B(pi1155), .ZN(new_n20758_));
  NOR2_X1    g17719(.A1(new_n20758_), .A2(new_n11923_), .ZN(new_n20759_));
  NOR3_X1    g17720(.A1(new_n20754_), .A2(new_n11903_), .A3(new_n20759_), .ZN(new_n20760_));
  NAND3_X1   g17721(.A1(new_n20743_), .A2(new_n20741_), .A3(new_n11903_), .ZN(new_n20761_));
  INV_X1     g17722(.I(new_n20720_), .ZN(new_n20762_));
  NOR2_X1    g17723(.A1(new_n20762_), .A2(new_n11914_), .ZN(new_n20763_));
  AOI22_X1   g17724(.A1(new_n20763_), .A2(pi0609), .B1(new_n13010_), .B2(new_n20749_), .ZN(new_n20764_));
  NOR2_X1    g17725(.A1(new_n11923_), .A2(pi1155), .ZN(new_n20765_));
  OAI21_X1   g17726(.A1(new_n20752_), .A2(new_n11903_), .B(new_n20765_), .ZN(new_n20766_));
  INV_X1     g17727(.I(new_n20766_), .ZN(new_n20767_));
  AOI22_X1   g17728(.A1(new_n20747_), .A2(new_n20760_), .B1(new_n20761_), .B2(new_n20767_), .ZN(new_n20768_));
  NOR3_X1    g17729(.A1(new_n20768_), .A2(new_n11870_), .A3(new_n20746_), .ZN(new_n20769_));
  NAND2_X1   g17730(.A1(new_n20747_), .A2(new_n20760_), .ZN(new_n20770_));
  NAND2_X1   g17731(.A1(new_n20761_), .A2(new_n20767_), .ZN(new_n20771_));
  NAND2_X1   g17732(.A1(new_n20770_), .A2(new_n20771_), .ZN(new_n20772_));
  AOI21_X1   g17733(.A1(new_n20772_), .A2(pi0785), .B(new_n20745_), .ZN(new_n20773_));
  NOR3_X1    g17734(.A1(new_n20773_), .A2(pi0781), .A3(new_n20769_), .ZN(new_n20774_));
  INV_X1     g17735(.I(new_n20774_), .ZN(new_n20775_));
  NOR2_X1    g17736(.A1(new_n20773_), .A2(new_n20769_), .ZN(new_n20776_));
  NOR2_X1    g17737(.A1(new_n20749_), .A2(new_n11938_), .ZN(new_n20777_));
  AOI21_X1   g17738(.A1(new_n20753_), .A2(new_n11938_), .B(new_n20777_), .ZN(new_n20778_));
  INV_X1     g17739(.I(new_n20778_), .ZN(new_n20779_));
  AOI21_X1   g17740(.A1(new_n20779_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n20780_));
  AOI21_X1   g17741(.A1(new_n20733_), .A2(new_n11914_), .B(pi0785), .ZN(new_n20781_));
  OAI21_X1   g17742(.A1(new_n20720_), .A2(new_n11914_), .B(new_n20781_), .ZN(new_n20782_));
  NOR2_X1    g17743(.A1(new_n20764_), .A2(new_n11912_), .ZN(new_n20783_));
  OAI21_X1   g17744(.A1(new_n20783_), .A2(new_n20758_), .B(pi0785), .ZN(new_n20784_));
  NOR2_X1    g17745(.A1(new_n20784_), .A2(new_n20782_), .ZN(new_n20785_));
  AND2_X2    g17746(.A1(new_n20784_), .A2(new_n20782_), .Z(new_n20786_));
  NOR3_X1    g17747(.A1(new_n20786_), .A2(new_n11934_), .A3(new_n20785_), .ZN(new_n20787_));
  NOR2_X1    g17748(.A1(new_n20749_), .A2(new_n11934_), .ZN(new_n20788_));
  NOR4_X1    g17749(.A1(new_n20787_), .A2(new_n11949_), .A3(pi1154), .A4(new_n20788_), .ZN(new_n20789_));
  NOR3_X1    g17750(.A1(new_n20789_), .A2(new_n11934_), .A3(new_n20780_), .ZN(new_n20790_));
  NAND3_X1   g17751(.A1(new_n20772_), .A2(pi0785), .A3(new_n20745_), .ZN(new_n20791_));
  OAI21_X1   g17752(.A1(new_n20768_), .A2(new_n11870_), .B(new_n20746_), .ZN(new_n20792_));
  NAND3_X1   g17753(.A1(new_n20791_), .A2(new_n20792_), .A3(new_n11934_), .ZN(new_n20793_));
  NOR2_X1    g17754(.A1(new_n20733_), .A2(pi0618), .ZN(new_n20794_));
  OR3_X2     g17755(.A1(new_n20787_), .A2(pi1154), .A3(new_n20794_), .Z(new_n20795_));
  AOI21_X1   g17756(.A1(new_n20779_), .A2(pi0618), .B(pi1154), .ZN(new_n20796_));
  INV_X1     g17757(.I(new_n20796_), .ZN(new_n20797_));
  AOI21_X1   g17758(.A1(new_n20795_), .A2(new_n11949_), .B(new_n20797_), .ZN(new_n20798_));
  AOI22_X1   g17759(.A1(new_n20793_), .A2(new_n20798_), .B1(new_n20776_), .B2(new_n20790_), .ZN(new_n20799_));
  NOR3_X1    g17760(.A1(new_n20799_), .A2(new_n11969_), .A3(new_n20775_), .ZN(new_n20800_));
  NAND3_X1   g17761(.A1(new_n20791_), .A2(new_n20790_), .A3(new_n20792_), .ZN(new_n20801_));
  NOR3_X1    g17762(.A1(new_n20773_), .A2(new_n20769_), .A3(pi0618), .ZN(new_n20802_));
  INV_X1     g17763(.I(new_n20798_), .ZN(new_n20803_));
  OAI21_X1   g17764(.A1(new_n20802_), .A2(new_n20803_), .B(new_n20801_), .ZN(new_n20804_));
  AOI21_X1   g17765(.A1(new_n20804_), .A2(pi0781), .B(new_n20774_), .ZN(new_n20805_));
  NOR3_X1    g17766(.A1(new_n20800_), .A2(new_n20805_), .A3(pi0789), .ZN(new_n20806_));
  INV_X1     g17767(.I(new_n20806_), .ZN(new_n20807_));
  NOR2_X1    g17768(.A1(new_n20800_), .A2(new_n20805_), .ZN(new_n20808_));
  NOR2_X1    g17769(.A1(new_n20786_), .A2(new_n20785_), .ZN(new_n20809_));
  NAND3_X1   g17770(.A1(new_n20749_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n20810_));
  MUX2_X1    g17771(.I0(new_n20810_), .I1(new_n20809_), .S(new_n11969_), .Z(new_n20811_));
  NAND2_X1   g17772(.A1(new_n20811_), .A2(pi0619), .ZN(new_n20812_));
  AOI21_X1   g17773(.A1(new_n20733_), .A2(pi0619), .B(pi1159), .ZN(new_n20813_));
  AND3_X2    g17774(.A1(new_n20812_), .A2(pi0648), .A3(new_n20813_), .Z(new_n20814_));
  NOR2_X1    g17775(.A1(new_n20733_), .A2(new_n11961_), .ZN(new_n20815_));
  AOI21_X1   g17776(.A1(new_n20778_), .A2(new_n11961_), .B(new_n20815_), .ZN(new_n20816_));
  NOR3_X1    g17777(.A1(new_n20814_), .A2(new_n11967_), .A3(pi1159), .ZN(new_n20817_));
  NAND3_X1   g17778(.A1(new_n20804_), .A2(new_n20774_), .A3(pi0781), .ZN(new_n20818_));
  OAI21_X1   g17779(.A1(new_n20799_), .A2(new_n11969_), .B(new_n20775_), .ZN(new_n20819_));
  NAND3_X1   g17780(.A1(new_n20819_), .A2(new_n20818_), .A3(new_n11967_), .ZN(new_n20820_));
  AOI21_X1   g17781(.A1(new_n20749_), .A2(new_n11967_), .B(pi1159), .ZN(new_n20821_));
  NAND2_X1   g17782(.A1(new_n20812_), .A2(new_n20821_), .ZN(new_n20822_));
  NAND2_X1   g17783(.A1(new_n20822_), .A2(new_n11966_), .ZN(new_n20823_));
  AOI21_X1   g17784(.A1(new_n20816_), .A2(pi0619), .B(pi1159), .ZN(new_n20824_));
  NAND2_X1   g17785(.A1(new_n20823_), .A2(new_n20824_), .ZN(new_n20825_));
  INV_X1     g17786(.I(new_n20825_), .ZN(new_n20826_));
  AOI22_X1   g17787(.A1(new_n20820_), .A2(new_n20826_), .B1(new_n20808_), .B2(new_n20817_), .ZN(new_n20827_));
  NOR3_X1    g17788(.A1(new_n20827_), .A2(new_n11985_), .A3(new_n20807_), .ZN(new_n20828_));
  NAND3_X1   g17789(.A1(new_n20819_), .A2(new_n20818_), .A3(new_n20817_), .ZN(new_n20829_));
  NOR3_X1    g17790(.A1(new_n20800_), .A2(new_n20805_), .A3(pi0619), .ZN(new_n20830_));
  OAI21_X1   g17791(.A1(new_n20830_), .A2(new_n20825_), .B(new_n20829_), .ZN(new_n20831_));
  AOI21_X1   g17792(.A1(new_n20831_), .A2(pi0789), .B(new_n20806_), .ZN(new_n20832_));
  NOR2_X1    g17793(.A1(new_n20828_), .A2(new_n20832_), .ZN(new_n20833_));
  NAND3_X1   g17794(.A1(new_n20831_), .A2(pi0789), .A3(new_n20806_), .ZN(new_n20834_));
  OAI21_X1   g17795(.A1(new_n20827_), .A2(new_n11985_), .B(new_n20807_), .ZN(new_n20835_));
  NAND2_X1   g17796(.A1(new_n20811_), .A2(new_n11985_), .ZN(new_n20836_));
  NOR3_X1    g17797(.A1(new_n20733_), .A2(pi0619), .A3(pi1159), .ZN(new_n20837_));
  NOR2_X1    g17798(.A1(new_n20837_), .A2(new_n11985_), .ZN(new_n20838_));
  XOR2_X1    g17799(.A1(new_n20836_), .A2(new_n20838_), .Z(new_n20839_));
  INV_X1     g17800(.I(new_n20839_), .ZN(new_n20840_));
  NOR3_X1    g17801(.A1(new_n11994_), .A2(new_n11989_), .A3(pi1158), .ZN(new_n20841_));
  NAND2_X1   g17802(.A1(new_n20840_), .A2(new_n20841_), .ZN(new_n20842_));
  NOR2_X1    g17803(.A1(new_n20749_), .A2(new_n12014_), .ZN(new_n20843_));
  AOI21_X1   g17804(.A1(new_n20816_), .A2(new_n12014_), .B(new_n20843_), .ZN(new_n20844_));
  NOR2_X1    g17805(.A1(new_n11994_), .A2(pi0641), .ZN(new_n20845_));
  NAND2_X1   g17806(.A1(new_n20842_), .A2(new_n20845_), .ZN(new_n20846_));
  NOR2_X1    g17807(.A1(new_n20839_), .A2(pi0626), .ZN(new_n20847_));
  OAI21_X1   g17808(.A1(new_n20733_), .A2(new_n11994_), .B(pi0641), .ZN(new_n20848_));
  NOR3_X1    g17809(.A1(new_n11989_), .A2(pi0626), .A3(pi1158), .ZN(new_n20849_));
  OAI21_X1   g17810(.A1(new_n20847_), .A2(new_n20848_), .B(new_n20849_), .ZN(new_n20850_));
  AOI22_X1   g17811(.A1(new_n20835_), .A2(new_n20834_), .B1(new_n20846_), .B2(new_n20850_), .ZN(new_n20851_));
  NAND3_X1   g17812(.A1(new_n20851_), .A2(pi0788), .A3(new_n20833_), .ZN(new_n20852_));
  NAND2_X1   g17813(.A1(new_n20835_), .A2(new_n20834_), .ZN(new_n20853_));
  OAI21_X1   g17814(.A1(new_n20851_), .A2(new_n11986_), .B(new_n20853_), .ZN(new_n20854_));
  NAND2_X1   g17815(.A1(new_n20854_), .A2(new_n20852_), .ZN(new_n20855_));
  INV_X1     g17816(.I(new_n20846_), .ZN(new_n20856_));
  INV_X1     g17817(.I(new_n20850_), .ZN(new_n20857_));
  OAI22_X1   g17818(.A1(new_n20828_), .A2(new_n20832_), .B1(new_n20856_), .B2(new_n20857_), .ZN(new_n20858_));
  NOR3_X1    g17819(.A1(new_n20858_), .A2(new_n11986_), .A3(new_n20853_), .ZN(new_n20859_));
  AOI21_X1   g17820(.A1(new_n20858_), .A2(pi0788), .B(new_n20833_), .ZN(new_n20860_));
  NOR2_X1    g17821(.A1(new_n20839_), .A2(new_n11997_), .ZN(new_n20861_));
  AOI21_X1   g17822(.A1(new_n11997_), .A2(new_n20749_), .B(new_n20861_), .ZN(new_n20862_));
  INV_X1     g17823(.I(new_n20862_), .ZN(new_n20863_));
  OAI21_X1   g17824(.A1(new_n20863_), .A2(pi0628), .B(pi1156), .ZN(new_n20864_));
  NOR2_X1    g17825(.A1(new_n20733_), .A2(new_n13114_), .ZN(new_n20865_));
  AOI21_X1   g17826(.A1(new_n20844_), .A2(new_n13114_), .B(new_n20865_), .ZN(new_n20866_));
  NOR3_X1    g17827(.A1(new_n20749_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n20867_));
  NOR2_X1    g17828(.A1(new_n20867_), .A2(new_n12030_), .ZN(new_n20868_));
  NOR2_X1    g17829(.A1(new_n20868_), .A2(new_n12031_), .ZN(new_n20869_));
  NAND2_X1   g17830(.A1(new_n20864_), .A2(new_n20869_), .ZN(new_n20870_));
  INV_X1     g17831(.I(new_n20870_), .ZN(new_n20871_));
  NOR2_X1    g17832(.A1(new_n20863_), .A2(new_n12031_), .ZN(new_n20872_));
  NOR2_X1    g17833(.A1(new_n12030_), .A2(pi0628), .ZN(new_n20873_));
  OAI21_X1   g17834(.A1(new_n20872_), .A2(pi1156), .B(new_n20873_), .ZN(new_n20874_));
  INV_X1     g17835(.I(new_n20874_), .ZN(new_n20875_));
  OAI22_X1   g17836(.A1(new_n20859_), .A2(new_n20860_), .B1(new_n20871_), .B2(new_n20875_), .ZN(new_n20876_));
  NOR3_X1    g17837(.A1(new_n20876_), .A2(new_n11868_), .A3(new_n20855_), .ZN(new_n20877_));
  NOR2_X1    g17838(.A1(new_n20859_), .A2(new_n20860_), .ZN(new_n20878_));
  AOI21_X1   g17839(.A1(new_n20876_), .A2(pi0792), .B(new_n20878_), .ZN(new_n20879_));
  NOR2_X1    g17840(.A1(new_n20877_), .A2(new_n20879_), .ZN(new_n20880_));
  AOI22_X1   g17841(.A1(new_n20854_), .A2(new_n20852_), .B1(new_n20870_), .B2(new_n20874_), .ZN(new_n20881_));
  NAND3_X1   g17842(.A1(new_n20881_), .A2(pi0792), .A3(new_n20878_), .ZN(new_n20882_));
  OAI21_X1   g17843(.A1(new_n20881_), .A2(new_n11868_), .B(new_n20855_), .ZN(new_n20883_));
  NAND2_X1   g17844(.A1(new_n20883_), .A2(new_n20882_), .ZN(new_n20884_));
  NOR4_X1    g17845(.A1(new_n20866_), .A2(new_n12031_), .A3(pi1156), .A4(new_n20733_), .ZN(new_n20885_));
  NOR2_X1    g17846(.A1(new_n20885_), .A2(new_n20867_), .ZN(new_n20886_));
  MUX2_X1    g17847(.I0(new_n20886_), .I1(new_n20866_), .S(new_n11868_), .Z(new_n20887_));
  NAND2_X1   g17848(.A1(new_n20887_), .A2(pi0647), .ZN(new_n20888_));
  AOI21_X1   g17849(.A1(new_n20733_), .A2(pi0647), .B(pi1157), .ZN(new_n20889_));
  NAND2_X1   g17850(.A1(new_n20888_), .A2(new_n20889_), .ZN(new_n20890_));
  NOR2_X1    g17851(.A1(new_n20733_), .A2(new_n12054_), .ZN(new_n20891_));
  AOI21_X1   g17852(.A1(new_n20863_), .A2(new_n12054_), .B(new_n20891_), .ZN(new_n20892_));
  NOR2_X1    g17853(.A1(new_n12061_), .A2(pi1157), .ZN(new_n20893_));
  OAI21_X1   g17854(.A1(new_n20890_), .A2(new_n12060_), .B(new_n20893_), .ZN(new_n20894_));
  NOR3_X1    g17855(.A1(new_n20877_), .A2(new_n20879_), .A3(pi0647), .ZN(new_n20895_));
  AOI21_X1   g17856(.A1(new_n20749_), .A2(new_n12061_), .B(pi1157), .ZN(new_n20896_));
  NAND2_X1   g17857(.A1(new_n20888_), .A2(new_n20896_), .ZN(new_n20897_));
  NAND2_X1   g17858(.A1(new_n20897_), .A2(new_n12060_), .ZN(new_n20898_));
  AOI21_X1   g17859(.A1(new_n20892_), .A2(pi0647), .B(pi1157), .ZN(new_n20899_));
  AND2_X2    g17860(.A1(new_n20899_), .A2(new_n20898_), .Z(new_n20900_));
  INV_X1     g17861(.I(new_n20900_), .ZN(new_n20901_));
  OAI22_X1   g17862(.A1(new_n20895_), .A2(new_n20901_), .B1(new_n20884_), .B2(new_n20894_), .ZN(new_n20902_));
  MUX2_X1    g17863(.I0(new_n20902_), .I1(new_n20880_), .S(new_n12048_), .Z(new_n20903_));
  INV_X1     g17864(.I(new_n20887_), .ZN(new_n20904_));
  NOR3_X1    g17865(.A1(new_n20733_), .A2(pi0647), .A3(pi1157), .ZN(new_n20905_));
  MUX2_X1    g17866(.I0(new_n20905_), .I1(new_n20904_), .S(new_n12048_), .Z(new_n20906_));
  NAND2_X1   g17867(.A1(new_n20906_), .A2(pi0644), .ZN(new_n20907_));
  NOR2_X1    g17868(.A1(new_n20749_), .A2(new_n12092_), .ZN(new_n20908_));
  AOI21_X1   g17869(.A1(new_n20892_), .A2(new_n12092_), .B(new_n20908_), .ZN(new_n20909_));
  NAND2_X1   g17870(.A1(new_n12082_), .A2(new_n12099_), .ZN(new_n20910_));
  OR2_X2     g17871(.A1(new_n20909_), .A2(new_n20910_), .Z(new_n20911_));
  NAND3_X1   g17872(.A1(new_n20911_), .A2(new_n20907_), .A3(new_n13168_), .ZN(new_n20912_));
  AOI21_X1   g17873(.A1(new_n20903_), .A2(new_n12082_), .B(new_n20912_), .ZN(new_n20913_));
  INV_X1     g17874(.I(new_n20894_), .ZN(new_n20914_));
  NAND3_X1   g17875(.A1(new_n20883_), .A2(new_n20882_), .A3(new_n12061_), .ZN(new_n20915_));
  AOI22_X1   g17876(.A1(new_n20915_), .A2(new_n20900_), .B1(new_n20880_), .B2(new_n20914_), .ZN(new_n20916_));
  MUX2_X1    g17877(.I0(new_n20916_), .I1(new_n20884_), .S(new_n12048_), .Z(new_n20917_));
  NAND3_X1   g17878(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n20918_));
  OAI21_X1   g17879(.A1(new_n20909_), .A2(new_n20918_), .B(new_n13179_), .ZN(new_n20919_));
  NOR2_X1    g17880(.A1(new_n20919_), .A2(new_n20906_), .ZN(new_n20920_));
  OAI21_X1   g17881(.A1(new_n20917_), .A2(new_n12082_), .B(new_n20920_), .ZN(new_n20921_));
  NOR2_X1    g17882(.A1(new_n20921_), .A2(new_n20913_), .ZN(new_n20922_));
  NAND2_X1   g17883(.A1(po1038), .A2(new_n8861_), .ZN(new_n20923_));
  AOI21_X1   g17884(.A1(new_n20923_), .A2(new_n13184_), .B(po1038), .ZN(new_n20924_));
  OAI21_X1   g17885(.A1(new_n20903_), .A2(pi0790), .B(new_n20924_), .ZN(new_n20925_));
  OAI21_X1   g17886(.A1(new_n20922_), .A2(new_n20925_), .B(new_n20710_), .ZN(po0344));
  NOR2_X1    g17887(.A1(new_n2925_), .A2(pi0188), .ZN(new_n20927_));
  NOR2_X1    g17888(.A1(new_n11877_), .A2(pi0768), .ZN(new_n20928_));
  NOR2_X1    g17889(.A1(new_n20928_), .A2(new_n20927_), .ZN(new_n20929_));
  INV_X1     g17890(.I(new_n20929_), .ZN(new_n20930_));
  AOI21_X1   g17891(.A1(new_n11886_), .A2(pi0705), .B(new_n20927_), .ZN(new_n20931_));
  NOR2_X1    g17892(.A1(new_n20931_), .A2(new_n11874_), .ZN(new_n20932_));
  NOR2_X1    g17893(.A1(new_n20930_), .A2(new_n20932_), .ZN(new_n20933_));
  NOR2_X1    g17894(.A1(new_n20933_), .A2(pi0778), .ZN(new_n20934_));
  NAND2_X1   g17895(.A1(new_n20932_), .A2(pi0625), .ZN(new_n20935_));
  NOR2_X1    g17896(.A1(new_n13201_), .A2(new_n16198_), .ZN(new_n20936_));
  NOR4_X1    g17897(.A1(new_n20928_), .A2(pi0608), .A3(new_n11893_), .A4(new_n20927_), .ZN(new_n20937_));
  OAI21_X1   g17898(.A1(new_n20930_), .A2(new_n20932_), .B(new_n20935_), .ZN(new_n20938_));
  NOR3_X1    g17899(.A1(new_n20927_), .A2(pi0608), .A3(pi1153), .ZN(new_n20939_));
  AOI22_X1   g17900(.A1(new_n20938_), .A2(new_n20939_), .B1(new_n20935_), .B2(new_n20937_), .ZN(new_n20940_));
  NOR2_X1    g17901(.A1(new_n20940_), .A2(new_n11891_), .ZN(new_n20941_));
  XOR2_X1    g17902(.A1(new_n20941_), .A2(new_n20934_), .Z(new_n20942_));
  INV_X1     g17903(.I(new_n20942_), .ZN(new_n20943_));
  NAND2_X1   g17904(.A1(new_n20943_), .A2(new_n11870_), .ZN(new_n20944_));
  AOI21_X1   g17905(.A1(new_n20942_), .A2(new_n11903_), .B(pi1155), .ZN(new_n20945_));
  INV_X1     g17906(.I(new_n20931_), .ZN(new_n20946_));
  XOR2_X1    g17907(.A1(new_n20936_), .A2(pi1153), .Z(new_n20947_));
  NAND2_X1   g17908(.A1(new_n20947_), .A2(new_n20946_), .ZN(new_n20948_));
  OAI21_X1   g17909(.A1(new_n20936_), .A2(new_n20927_), .B(new_n11893_), .ZN(new_n20949_));
  AOI21_X1   g17910(.A1(new_n20948_), .A2(new_n20949_), .B(new_n11891_), .ZN(new_n20950_));
  NOR2_X1    g17911(.A1(new_n20931_), .A2(pi0778), .ZN(new_n20951_));
  OAI21_X1   g17912(.A1(new_n20950_), .A2(new_n20951_), .B(pi0609), .ZN(new_n20952_));
  AOI21_X1   g17913(.A1(new_n20930_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n20953_));
  NOR2_X1    g17914(.A1(new_n20953_), .A2(pi0660), .ZN(new_n20954_));
  OAI21_X1   g17915(.A1(new_n20945_), .A2(new_n20952_), .B(new_n20954_), .ZN(new_n20955_));
  NOR2_X1    g17916(.A1(new_n20950_), .A2(new_n20951_), .ZN(new_n20956_));
  NAND4_X1   g17917(.A1(new_n20943_), .A2(pi0609), .A3(new_n11912_), .A4(new_n20956_), .ZN(new_n20957_));
  NOR2_X1    g17918(.A1(new_n20929_), .A2(new_n11925_), .ZN(new_n20958_));
  AOI21_X1   g17919(.A1(new_n20958_), .A2(new_n11928_), .B(pi1155), .ZN(new_n20959_));
  NOR2_X1    g17920(.A1(new_n20959_), .A2(new_n11923_), .ZN(new_n20960_));
  NAND2_X1   g17921(.A1(new_n20957_), .A2(new_n20960_), .ZN(new_n20961_));
  NAND3_X1   g17922(.A1(new_n20961_), .A2(pi0785), .A3(new_n20955_), .ZN(new_n20962_));
  NAND2_X1   g17923(.A1(new_n20962_), .A2(new_n20944_), .ZN(new_n20963_));
  NOR4_X1    g17924(.A1(new_n20956_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n20965_));
  NOR2_X1    g17925(.A1(new_n20958_), .A2(pi0785), .ZN(new_n20966_));
  OAI21_X1   g17926(.A1(new_n20959_), .A2(new_n20953_), .B(pi0785), .ZN(new_n20967_));
  XNOR2_X1   g17927(.A1(new_n20967_), .A2(new_n20966_), .ZN(new_n20968_));
  INV_X1     g17928(.I(new_n20968_), .ZN(new_n20969_));
  NOR2_X1    g17929(.A1(new_n20969_), .A2(new_n11945_), .ZN(new_n20970_));
  NOR3_X1    g17930(.A1(new_n20965_), .A2(new_n20970_), .A3(pi0627), .ZN(new_n20971_));
  AOI21_X1   g17931(.A1(new_n20968_), .A2(new_n11951_), .B(pi1154), .ZN(new_n20972_));
  NOR2_X1    g17932(.A1(new_n20956_), .A2(new_n11939_), .ZN(new_n20973_));
  INV_X1     g17933(.I(new_n20973_), .ZN(new_n20974_));
  NAND4_X1   g17934(.A1(new_n20963_), .A2(pi0618), .A3(new_n11950_), .A4(new_n20974_), .ZN(new_n20975_));
  NAND2_X1   g17935(.A1(new_n20975_), .A2(new_n20972_), .ZN(new_n20976_));
  AOI21_X1   g17936(.A1(new_n20976_), .A2(new_n11949_), .B(new_n20971_), .ZN(new_n20977_));
  NOR2_X1    g17937(.A1(new_n20977_), .A2(new_n11969_), .ZN(new_n20978_));
  AOI21_X1   g17938(.A1(new_n11969_), .A2(new_n20963_), .B(new_n20978_), .ZN(new_n20979_));
  NOR2_X1    g17939(.A1(new_n20974_), .A2(new_n11962_), .ZN(new_n20980_));
  NOR4_X1    g17940(.A1(new_n20979_), .A2(new_n11967_), .A3(pi1159), .A4(new_n20980_), .ZN(new_n20981_));
  INV_X1     g17941(.I(new_n20970_), .ZN(new_n20982_));
  NAND2_X1   g17942(.A1(new_n20982_), .A2(new_n20972_), .ZN(new_n20983_));
  MUX2_X1    g17943(.I0(new_n20983_), .I1(new_n20968_), .S(new_n11969_), .Z(new_n20984_));
  NAND2_X1   g17944(.A1(new_n20984_), .A2(pi0619), .ZN(new_n20985_));
  INV_X1     g17945(.I(new_n20985_), .ZN(new_n20986_));
  INV_X1     g17946(.I(new_n20927_), .ZN(new_n20987_));
  OAI21_X1   g17947(.A1(new_n20987_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n20988_));
  NOR4_X1    g17948(.A1(new_n20981_), .A2(new_n11966_), .A3(new_n20986_), .A4(new_n20988_), .ZN(new_n20989_));
  NOR4_X1    g17949(.A1(new_n20974_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n20990_));
  OAI21_X1   g17950(.A1(new_n20927_), .A2(pi0619), .B(new_n11869_), .ZN(new_n20991_));
  OAI21_X1   g17951(.A1(new_n20986_), .A2(new_n20991_), .B(new_n11966_), .ZN(new_n20992_));
  NOR2_X1    g17952(.A1(new_n20992_), .A2(new_n20990_), .ZN(new_n20993_));
  AOI21_X1   g17953(.A1(new_n20979_), .A2(new_n11998_), .B(pi0789), .ZN(new_n20994_));
  OAI21_X1   g17954(.A1(new_n20989_), .A2(new_n20993_), .B(new_n20994_), .ZN(new_n20995_));
  NAND2_X1   g17955(.A1(new_n20980_), .A2(new_n17450_), .ZN(new_n20996_));
  NOR2_X1    g17956(.A1(new_n20996_), .A2(new_n17153_), .ZN(new_n20997_));
  INV_X1     g17957(.I(new_n20997_), .ZN(new_n20998_));
  NOR2_X1    g17958(.A1(new_n20998_), .A2(new_n17151_), .ZN(new_n20999_));
  NOR2_X1    g17959(.A1(new_n14624_), .A2(new_n20927_), .ZN(new_n21000_));
  NAND3_X1   g17960(.A1(new_n20987_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n21001_));
  MUX2_X1    g17961(.I0(new_n21001_), .I1(new_n20984_), .S(new_n11985_), .Z(new_n21002_));
  AOI21_X1   g17962(.A1(new_n21002_), .A2(new_n14624_), .B(new_n21000_), .ZN(new_n21003_));
  AND2_X2    g17963(.A1(new_n21003_), .A2(new_n12064_), .Z(new_n21004_));
  OAI21_X1   g17964(.A1(new_n21004_), .A2(new_n20999_), .B(pi0629), .ZN(new_n21005_));
  NAND2_X1   g17965(.A1(new_n21003_), .A2(new_n12063_), .ZN(new_n21006_));
  NAND2_X1   g17966(.A1(new_n20997_), .A2(new_n15084_), .ZN(new_n21007_));
  NAND4_X1   g17967(.A1(new_n21005_), .A2(new_n15085_), .A3(new_n21006_), .A4(new_n21007_), .ZN(new_n21008_));
  MUX2_X1    g17968(.I0(new_n21002_), .I1(new_n20987_), .S(new_n11994_), .Z(new_n21009_));
  NOR2_X1    g17969(.A1(new_n21009_), .A2(new_n17167_), .ZN(new_n21010_));
  OAI21_X1   g17970(.A1(new_n21002_), .A2(new_n20927_), .B(pi0626), .ZN(new_n21011_));
  NOR2_X1    g17971(.A1(new_n20996_), .A2(new_n12020_), .ZN(new_n21012_));
  NOR2_X1    g17972(.A1(new_n21012_), .A2(pi0788), .ZN(new_n21013_));
  OAI21_X1   g17973(.A1(new_n21011_), .A2(new_n17171_), .B(new_n21013_), .ZN(new_n21014_));
  OAI21_X1   g17974(.A1(new_n21010_), .A2(new_n21014_), .B(new_n14732_), .ZN(new_n21015_));
  AOI21_X1   g17975(.A1(new_n21008_), .A2(new_n14726_), .B(new_n21015_), .ZN(new_n21016_));
  NAND3_X1   g17976(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n20927_), .ZN(new_n21017_));
  NOR2_X1    g17977(.A1(new_n20998_), .A2(new_n12068_), .ZN(new_n21018_));
  INV_X1     g17978(.I(new_n21018_), .ZN(new_n21019_));
  NAND2_X1   g17979(.A1(new_n21019_), .A2(pi0647), .ZN(new_n21020_));
  NAND2_X1   g17980(.A1(new_n20927_), .A2(pi0647), .ZN(new_n21021_));
  NAND3_X1   g17981(.A1(new_n21020_), .A2(new_n12049_), .A3(new_n21021_), .ZN(new_n21022_));
  NOR2_X1    g17982(.A1(new_n20987_), .A2(pi0647), .ZN(new_n21023_));
  AOI21_X1   g17983(.A1(new_n21018_), .A2(pi0647), .B(new_n21023_), .ZN(new_n21024_));
  NAND2_X1   g17984(.A1(new_n21024_), .A2(new_n12088_), .ZN(new_n21025_));
  NAND2_X1   g17985(.A1(new_n21025_), .A2(pi0787), .ZN(new_n21026_));
  AOI21_X1   g17986(.A1(pi0630), .A2(new_n21022_), .B(new_n21026_), .ZN(new_n21027_));
  AOI22_X1   g17987(.A1(new_n20995_), .A2(new_n21016_), .B1(new_n21017_), .B2(new_n21027_), .ZN(new_n21028_));
  NOR2_X1    g17988(.A1(new_n21028_), .A2(new_n12082_), .ZN(new_n21029_));
  NAND4_X1   g17989(.A1(new_n21020_), .A2(pi0787), .A3(new_n12049_), .A4(new_n21021_), .ZN(new_n21030_));
  OAI21_X1   g17990(.A1(pi0787), .A2(new_n21019_), .B(new_n21030_), .ZN(new_n21031_));
  NOR2_X1    g17991(.A1(new_n21031_), .A2(pi0644), .ZN(new_n21032_));
  OR3_X2     g17992(.A1(new_n21029_), .A2(pi0715), .A3(new_n21032_), .Z(new_n21033_));
  MUX2_X1    g17993(.I0(new_n21003_), .I1(new_n20927_), .S(new_n16841_), .Z(new_n21034_));
  INV_X1     g17994(.I(new_n21034_), .ZN(new_n21035_));
  OAI21_X1   g17995(.A1(new_n21034_), .A2(new_n20927_), .B(new_n12082_), .ZN(new_n21036_));
  AOI21_X1   g17996(.A1(new_n20927_), .A2(new_n21034_), .B(new_n21036_), .ZN(new_n21037_));
  OAI21_X1   g17997(.A1(new_n21037_), .A2(new_n21035_), .B(new_n12099_), .ZN(new_n21038_));
  AOI21_X1   g17998(.A1(new_n21035_), .A2(new_n21037_), .B(new_n21038_), .ZN(new_n21039_));
  AOI21_X1   g17999(.A1(new_n21033_), .A2(new_n21039_), .B(pi1160), .ZN(new_n21040_));
  XOR2_X1    g18000(.A1(new_n21037_), .A2(new_n20927_), .Z(new_n21041_));
  AOI21_X1   g18001(.A1(new_n21031_), .A2(pi0644), .B(new_n13169_), .ZN(new_n21042_));
  OAI21_X1   g18002(.A1(new_n21041_), .A2(new_n12099_), .B(new_n21042_), .ZN(new_n21043_));
  OAI21_X1   g18003(.A1(new_n21029_), .A2(new_n21043_), .B(pi0790), .ZN(new_n21044_));
  NOR2_X1    g18004(.A1(new_n21028_), .A2(new_n14748_), .ZN(new_n21045_));
  OAI21_X1   g18005(.A1(new_n21040_), .A2(new_n21044_), .B(new_n21045_), .ZN(new_n21046_));
  NOR2_X1    g18006(.A1(new_n3231_), .A2(pi0188), .ZN(new_n21047_));
  INV_X1     g18007(.I(new_n21047_), .ZN(new_n21048_));
  NOR2_X1    g18008(.A1(pi0188), .A2(pi0705), .ZN(new_n21049_));
  NAND2_X1   g18009(.A1(new_n20353_), .A2(pi0188), .ZN(new_n21050_));
  AOI21_X1   g18010(.A1(new_n21050_), .A2(new_n17798_), .B(pi0768), .ZN(new_n21051_));
  OAI21_X1   g18011(.A1(pi0768), .A2(new_n14365_), .B(new_n16211_), .ZN(new_n21052_));
  AOI21_X1   g18012(.A1(new_n21052_), .A2(new_n7356_), .B(new_n21051_), .ZN(new_n21053_));
  AOI22_X1   g18013(.A1(new_n21053_), .A2(new_n16198_), .B1(new_n14347_), .B2(new_n21049_), .ZN(new_n21054_));
  NOR2_X1    g18014(.A1(new_n21054_), .A2(new_n3232_), .ZN(new_n21055_));
  XOR2_X1    g18015(.A1(new_n21055_), .A2(new_n21048_), .Z(new_n21056_));
  AOI21_X1   g18016(.A1(new_n21053_), .A2(new_n3231_), .B(new_n21047_), .ZN(new_n21057_));
  INV_X1     g18017(.I(new_n21057_), .ZN(new_n21058_));
  AOI21_X1   g18018(.A1(new_n21058_), .A2(new_n12970_), .B(new_n11893_), .ZN(new_n21059_));
  NAND2_X1   g18019(.A1(new_n7356_), .A2(new_n16198_), .ZN(new_n21060_));
  OAI21_X1   g18020(.A1(new_n12902_), .A2(new_n21060_), .B(new_n3231_), .ZN(new_n21061_));
  NOR3_X1    g18021(.A1(new_n13399_), .A2(pi0188), .A3(new_n13396_), .ZN(new_n21062_));
  AOI21_X1   g18022(.A1(new_n13399_), .A2(new_n7356_), .B(new_n13395_), .ZN(new_n21063_));
  NAND2_X1   g18023(.A1(new_n13368_), .A2(new_n7356_), .ZN(new_n21064_));
  NAND4_X1   g18024(.A1(new_n21064_), .A2(new_n3172_), .A3(new_n16198_), .A4(new_n13403_), .ZN(new_n21065_));
  NOR3_X1    g18025(.A1(new_n21062_), .A2(new_n21063_), .A3(new_n21065_), .ZN(new_n21066_));
  AOI22_X1   g18026(.A1(new_n21066_), .A2(new_n21061_), .B1(pi0188), .B2(new_n3232_), .ZN(new_n21067_));
  INV_X1     g18027(.I(new_n21067_), .ZN(new_n21068_));
  NOR2_X1    g18028(.A1(new_n12965_), .A2(pi0188), .ZN(new_n21069_));
  AOI21_X1   g18029(.A1(new_n21068_), .A2(new_n20723_), .B(new_n12970_), .ZN(new_n21070_));
  INV_X1     g18030(.I(new_n21070_), .ZN(new_n21071_));
  OR2_X2     g18031(.A1(new_n21059_), .A2(new_n21071_), .Z(new_n21072_));
  NOR2_X1    g18032(.A1(new_n21057_), .A2(new_n12970_), .ZN(new_n21073_));
  NOR2_X1    g18033(.A1(pi0608), .A2(pi0625), .ZN(new_n21075_));
  OAI21_X1   g18034(.A1(new_n21073_), .A2(pi1153), .B(new_n21075_), .ZN(new_n21076_));
  NAND4_X1   g18035(.A1(new_n21072_), .A2(new_n21056_), .A3(pi0778), .A4(new_n21076_), .ZN(new_n21077_));
  NOR2_X1    g18036(.A1(new_n21077_), .A2(new_n21056_), .ZN(new_n21078_));
  XOR2_X1    g18037(.A1(new_n21055_), .A2(new_n21047_), .Z(new_n21079_));
  NOR2_X1    g18038(.A1(new_n21059_), .A2(new_n21071_), .ZN(new_n21080_));
  INV_X1     g18039(.I(new_n21076_), .ZN(new_n21081_));
  NOR4_X1    g18040(.A1(new_n21079_), .A2(new_n11891_), .A3(new_n21080_), .A4(new_n21081_), .ZN(new_n21082_));
  NOR2_X1    g18041(.A1(new_n21082_), .A2(new_n21079_), .ZN(new_n21083_));
  NOR2_X1    g18042(.A1(new_n21078_), .A2(new_n21083_), .ZN(new_n21084_));
  NAND2_X1   g18043(.A1(new_n21084_), .A2(new_n11870_), .ZN(new_n21085_));
  NOR2_X1    g18044(.A1(new_n21067_), .A2(pi0778), .ZN(new_n21086_));
  INV_X1     g18045(.I(new_n21069_), .ZN(new_n21087_));
  MUX2_X1    g18046(.I0(new_n21087_), .I1(new_n21067_), .S(new_n13435_), .Z(new_n21088_));
  NOR2_X1    g18047(.A1(new_n21088_), .A2(new_n11891_), .ZN(new_n21089_));
  NOR2_X1    g18048(.A1(new_n21089_), .A2(new_n21086_), .ZN(new_n21090_));
  INV_X1     g18049(.I(new_n21090_), .ZN(new_n21091_));
  NAND2_X1   g18050(.A1(new_n21091_), .A2(new_n11903_), .ZN(new_n21092_));
  NAND2_X1   g18051(.A1(new_n21092_), .A2(pi1155), .ZN(new_n21093_));
  NOR2_X1    g18052(.A1(new_n21069_), .A2(new_n12996_), .ZN(new_n21094_));
  INV_X1     g18053(.I(new_n21094_), .ZN(new_n21095_));
  NAND3_X1   g18054(.A1(new_n21057_), .A2(new_n11903_), .A3(new_n11924_), .ZN(new_n21096_));
  AOI21_X1   g18055(.A1(new_n21096_), .A2(new_n21095_), .B(pi1155), .ZN(new_n21097_));
  OR2_X2     g18056(.A1(new_n21097_), .A2(new_n11923_), .Z(new_n21098_));
  NAND3_X1   g18057(.A1(new_n21093_), .A2(pi0609), .A3(new_n21098_), .ZN(new_n21099_));
  INV_X1     g18058(.I(new_n21099_), .ZN(new_n21100_));
  NOR2_X1    g18059(.A1(new_n21072_), .A2(new_n21079_), .ZN(new_n21101_));
  NAND3_X1   g18060(.A1(new_n21101_), .A2(pi0778), .A3(new_n21079_), .ZN(new_n21102_));
  NAND2_X1   g18061(.A1(new_n21077_), .A2(new_n21056_), .ZN(new_n21103_));
  NAND3_X1   g18062(.A1(new_n21103_), .A2(new_n21102_), .A3(new_n11903_), .ZN(new_n21104_));
  NOR2_X1    g18063(.A1(new_n21058_), .A2(new_n11914_), .ZN(new_n21105_));
  NOR2_X1    g18064(.A1(new_n21069_), .A2(new_n11915_), .ZN(new_n21106_));
  AOI21_X1   g18065(.A1(new_n21105_), .A2(pi0609), .B(new_n21106_), .ZN(new_n21107_));
  NOR2_X1    g18066(.A1(new_n11923_), .A2(pi1155), .ZN(new_n21108_));
  OAI21_X1   g18067(.A1(new_n21090_), .A2(new_n11903_), .B(new_n21108_), .ZN(new_n21109_));
  INV_X1     g18068(.I(new_n21109_), .ZN(new_n21110_));
  AOI22_X1   g18069(.A1(new_n21104_), .A2(new_n21110_), .B1(new_n21084_), .B2(new_n21100_), .ZN(new_n21111_));
  NOR3_X1    g18070(.A1(new_n21111_), .A2(new_n11870_), .A3(new_n21085_), .ZN(new_n21112_));
  NAND2_X1   g18071(.A1(new_n21103_), .A2(new_n21102_), .ZN(new_n21113_));
  NOR2_X1    g18072(.A1(new_n21113_), .A2(pi0785), .ZN(new_n21114_));
  NOR3_X1    g18073(.A1(new_n21078_), .A2(new_n21083_), .A3(pi0609), .ZN(new_n21115_));
  OAI22_X1   g18074(.A1(new_n21115_), .A2(new_n21109_), .B1(new_n21113_), .B2(new_n21099_), .ZN(new_n21116_));
  AOI21_X1   g18075(.A1(new_n21116_), .A2(pi0785), .B(new_n21114_), .ZN(new_n21117_));
  NOR2_X1    g18076(.A1(new_n21112_), .A2(new_n21117_), .ZN(new_n21118_));
  NAND2_X1   g18077(.A1(new_n21118_), .A2(new_n11969_), .ZN(new_n21119_));
  INV_X1     g18078(.I(new_n21119_), .ZN(new_n21120_));
  NAND3_X1   g18079(.A1(new_n21116_), .A2(pi0785), .A3(new_n21114_), .ZN(new_n21121_));
  OAI21_X1   g18080(.A1(new_n21111_), .A2(new_n11870_), .B(new_n21085_), .ZN(new_n21122_));
  NOR2_X1    g18081(.A1(new_n21087_), .A2(new_n11938_), .ZN(new_n21123_));
  AOI21_X1   g18082(.A1(new_n21091_), .A2(new_n11938_), .B(new_n21123_), .ZN(new_n21124_));
  INV_X1     g18083(.I(new_n21124_), .ZN(new_n21125_));
  AOI21_X1   g18084(.A1(new_n21125_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n21126_));
  AOI21_X1   g18085(.A1(new_n21069_), .A2(new_n11914_), .B(pi0785), .ZN(new_n21127_));
  OAI21_X1   g18086(.A1(new_n21057_), .A2(new_n11914_), .B(new_n21127_), .ZN(new_n21128_));
  NOR2_X1    g18087(.A1(new_n21107_), .A2(new_n11912_), .ZN(new_n21129_));
  OAI21_X1   g18088(.A1(new_n21129_), .A2(new_n21097_), .B(pi0785), .ZN(new_n21130_));
  NOR2_X1    g18089(.A1(new_n21130_), .A2(new_n21128_), .ZN(new_n21131_));
  AND2_X2    g18090(.A1(new_n21130_), .A2(new_n21128_), .Z(new_n21132_));
  NOR3_X1    g18091(.A1(new_n21132_), .A2(new_n11934_), .A3(new_n21131_), .ZN(new_n21133_));
  OAI21_X1   g18092(.A1(new_n21087_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n21134_));
  NOR3_X1    g18093(.A1(new_n21133_), .A2(new_n11949_), .A3(new_n21134_), .ZN(new_n21135_));
  NOR3_X1    g18094(.A1(new_n21135_), .A2(new_n11934_), .A3(new_n21126_), .ZN(new_n21136_));
  NAND3_X1   g18095(.A1(new_n21136_), .A2(new_n21122_), .A3(new_n21121_), .ZN(new_n21137_));
  NOR3_X1    g18096(.A1(new_n21112_), .A2(new_n21117_), .A3(pi0618), .ZN(new_n21138_));
  NOR2_X1    g18097(.A1(new_n21069_), .A2(pi0618), .ZN(new_n21139_));
  OR3_X2     g18098(.A1(new_n21133_), .A2(pi1154), .A3(new_n21139_), .Z(new_n21140_));
  AOI21_X1   g18099(.A1(new_n21125_), .A2(pi0618), .B(pi1154), .ZN(new_n21141_));
  INV_X1     g18100(.I(new_n21141_), .ZN(new_n21142_));
  AOI21_X1   g18101(.A1(new_n21140_), .A2(new_n11949_), .B(new_n21142_), .ZN(new_n21143_));
  INV_X1     g18102(.I(new_n21143_), .ZN(new_n21144_));
  OAI21_X1   g18103(.A1(new_n21144_), .A2(new_n21138_), .B(new_n21137_), .ZN(new_n21145_));
  NAND3_X1   g18104(.A1(new_n21145_), .A2(new_n21120_), .A3(pi0781), .ZN(new_n21146_));
  NAND3_X1   g18105(.A1(new_n21122_), .A2(new_n21121_), .A3(new_n11934_), .ZN(new_n21147_));
  AOI22_X1   g18106(.A1(new_n21147_), .A2(new_n21143_), .B1(new_n21118_), .B2(new_n21136_), .ZN(new_n21148_));
  OAI21_X1   g18107(.A1(new_n21148_), .A2(new_n11969_), .B(new_n21119_), .ZN(new_n21149_));
  NAND2_X1   g18108(.A1(new_n21146_), .A2(new_n21149_), .ZN(new_n21150_));
  NOR2_X1    g18109(.A1(new_n21150_), .A2(pi0789), .ZN(new_n21151_));
  NOR2_X1    g18110(.A1(new_n21132_), .A2(new_n21131_), .ZN(new_n21152_));
  NAND3_X1   g18111(.A1(new_n21087_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n21153_));
  MUX2_X1    g18112(.I0(new_n21153_), .I1(new_n21152_), .S(new_n11969_), .Z(new_n21154_));
  AND2_X2    g18113(.A1(new_n21154_), .A2(pi0619), .Z(new_n21155_));
  OAI21_X1   g18114(.A1(new_n21087_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n21156_));
  NOR3_X1    g18115(.A1(new_n21155_), .A2(new_n11966_), .A3(new_n21156_), .ZN(new_n21157_));
  NOR2_X1    g18116(.A1(new_n21069_), .A2(new_n11961_), .ZN(new_n21158_));
  AOI21_X1   g18117(.A1(new_n21124_), .A2(new_n11961_), .B(new_n21158_), .ZN(new_n21159_));
  NOR3_X1    g18118(.A1(new_n21157_), .A2(new_n11967_), .A3(pi1159), .ZN(new_n21160_));
  NAND3_X1   g18119(.A1(new_n21146_), .A2(new_n21149_), .A3(new_n21160_), .ZN(new_n21161_));
  NOR3_X1    g18120(.A1(new_n21148_), .A2(new_n11969_), .A3(new_n21119_), .ZN(new_n21162_));
  AOI21_X1   g18121(.A1(new_n21145_), .A2(pi0781), .B(new_n21120_), .ZN(new_n21163_));
  NOR3_X1    g18122(.A1(new_n21163_), .A2(new_n21162_), .A3(pi0619), .ZN(new_n21164_));
  NOR2_X1    g18123(.A1(new_n21069_), .A2(pi0619), .ZN(new_n21165_));
  OR3_X2     g18124(.A1(new_n21155_), .A2(pi1159), .A3(new_n21165_), .Z(new_n21166_));
  AOI21_X1   g18125(.A1(new_n21159_), .A2(pi0619), .B(pi1159), .ZN(new_n21167_));
  INV_X1     g18126(.I(new_n21167_), .ZN(new_n21168_));
  AOI21_X1   g18127(.A1(new_n21166_), .A2(new_n11966_), .B(new_n21168_), .ZN(new_n21169_));
  INV_X1     g18128(.I(new_n21169_), .ZN(new_n21170_));
  OAI21_X1   g18129(.A1(new_n21164_), .A2(new_n21170_), .B(new_n21161_), .ZN(new_n21171_));
  NAND3_X1   g18130(.A1(new_n21171_), .A2(pi0789), .A3(new_n21151_), .ZN(new_n21172_));
  MUX2_X1    g18131(.I0(new_n21145_), .I1(new_n21118_), .S(new_n11969_), .Z(new_n21173_));
  NAND2_X1   g18132(.A1(new_n21173_), .A2(new_n11985_), .ZN(new_n21174_));
  NAND3_X1   g18133(.A1(new_n21146_), .A2(new_n21149_), .A3(new_n11967_), .ZN(new_n21175_));
  AOI22_X1   g18134(.A1(new_n21175_), .A2(new_n21169_), .B1(new_n21173_), .B2(new_n21160_), .ZN(new_n21176_));
  OAI21_X1   g18135(.A1(new_n21176_), .A2(new_n11985_), .B(new_n21174_), .ZN(new_n21177_));
  NAND2_X1   g18136(.A1(new_n21177_), .A2(new_n21172_), .ZN(new_n21178_));
  NOR3_X1    g18137(.A1(new_n21176_), .A2(new_n11985_), .A3(new_n21174_), .ZN(new_n21179_));
  AOI21_X1   g18138(.A1(new_n21171_), .A2(pi0789), .B(new_n21151_), .ZN(new_n21180_));
  NAND2_X1   g18139(.A1(new_n21154_), .A2(new_n11985_), .ZN(new_n21181_));
  NOR3_X1    g18140(.A1(new_n21069_), .A2(pi0619), .A3(pi1159), .ZN(new_n21182_));
  NOR2_X1    g18141(.A1(new_n21182_), .A2(new_n11985_), .ZN(new_n21183_));
  XNOR2_X1   g18142(.A1(new_n21181_), .A2(new_n21183_), .ZN(new_n21184_));
  NOR3_X1    g18143(.A1(new_n11994_), .A2(new_n11989_), .A3(pi1158), .ZN(new_n21185_));
  NAND2_X1   g18144(.A1(new_n21184_), .A2(new_n21185_), .ZN(new_n21186_));
  NOR2_X1    g18145(.A1(new_n21087_), .A2(new_n12014_), .ZN(new_n21187_));
  AOI21_X1   g18146(.A1(new_n21159_), .A2(new_n12014_), .B(new_n21187_), .ZN(new_n21188_));
  NOR2_X1    g18147(.A1(new_n11994_), .A2(pi0641), .ZN(new_n21189_));
  NAND2_X1   g18148(.A1(new_n21186_), .A2(new_n21189_), .ZN(new_n21190_));
  INV_X1     g18149(.I(new_n21190_), .ZN(new_n21191_));
  AND2_X2    g18150(.A1(new_n21184_), .A2(new_n11994_), .Z(new_n21192_));
  OAI21_X1   g18151(.A1(new_n21069_), .A2(new_n11994_), .B(pi0641), .ZN(new_n21193_));
  NOR3_X1    g18152(.A1(new_n11989_), .A2(pi0626), .A3(pi1158), .ZN(new_n21194_));
  OAI21_X1   g18153(.A1(new_n21192_), .A2(new_n21193_), .B(new_n21194_), .ZN(new_n21195_));
  INV_X1     g18154(.I(new_n21195_), .ZN(new_n21196_));
  OAI22_X1   g18155(.A1(new_n21180_), .A2(new_n21179_), .B1(new_n21191_), .B2(new_n21196_), .ZN(new_n21197_));
  NOR3_X1    g18156(.A1(new_n21197_), .A2(new_n11986_), .A3(new_n21178_), .ZN(new_n21198_));
  NOR2_X1    g18157(.A1(new_n21180_), .A2(new_n21179_), .ZN(new_n21199_));
  AOI21_X1   g18158(.A1(new_n21197_), .A2(pi0788), .B(new_n21199_), .ZN(new_n21200_));
  NOR2_X1    g18159(.A1(new_n21198_), .A2(new_n21200_), .ZN(new_n21201_));
  NOR2_X1    g18160(.A1(new_n21069_), .A2(new_n14624_), .ZN(new_n21202_));
  AOI21_X1   g18161(.A1(new_n21184_), .A2(new_n14624_), .B(new_n21202_), .ZN(new_n21203_));
  INV_X1     g18162(.I(new_n21203_), .ZN(new_n21204_));
  NOR2_X1    g18163(.A1(new_n21204_), .A2(pi0628), .ZN(new_n21205_));
  NOR2_X1    g18164(.A1(new_n21069_), .A2(new_n13114_), .ZN(new_n21206_));
  AOI21_X1   g18165(.A1(new_n21188_), .A2(new_n13114_), .B(new_n21206_), .ZN(new_n21207_));
  NOR3_X1    g18166(.A1(new_n21087_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n21208_));
  NOR2_X1    g18167(.A1(new_n21208_), .A2(new_n12030_), .ZN(new_n21209_));
  NOR2_X1    g18168(.A1(new_n21209_), .A2(new_n12031_), .ZN(new_n21210_));
  OAI21_X1   g18169(.A1(new_n21205_), .A2(new_n12026_), .B(new_n21210_), .ZN(new_n21211_));
  INV_X1     g18170(.I(new_n21211_), .ZN(new_n21212_));
  NOR2_X1    g18171(.A1(new_n21204_), .A2(new_n12031_), .ZN(new_n21213_));
  NOR2_X1    g18172(.A1(new_n12030_), .A2(pi0628), .ZN(new_n21214_));
  OAI21_X1   g18173(.A1(new_n21213_), .A2(pi1156), .B(new_n21214_), .ZN(new_n21215_));
  INV_X1     g18174(.I(new_n21215_), .ZN(new_n21216_));
  OAI22_X1   g18175(.A1(new_n21198_), .A2(new_n21200_), .B1(new_n21212_), .B2(new_n21216_), .ZN(new_n21217_));
  MUX2_X1    g18176(.I0(new_n21217_), .I1(new_n21201_), .S(new_n11868_), .Z(new_n21218_));
  AOI22_X1   g18177(.A1(new_n21177_), .A2(new_n21172_), .B1(new_n21190_), .B2(new_n21195_), .ZN(new_n21219_));
  NAND3_X1   g18178(.A1(new_n21219_), .A2(pi0788), .A3(new_n21199_), .ZN(new_n21220_));
  OAI21_X1   g18179(.A1(new_n21219_), .A2(new_n11986_), .B(new_n21178_), .ZN(new_n21221_));
  AOI22_X1   g18180(.A1(new_n21221_), .A2(new_n21220_), .B1(new_n21211_), .B2(new_n21215_), .ZN(new_n21222_));
  NAND3_X1   g18181(.A1(new_n21222_), .A2(pi0792), .A3(new_n21201_), .ZN(new_n21223_));
  NAND2_X1   g18182(.A1(new_n21221_), .A2(new_n21220_), .ZN(new_n21224_));
  OAI21_X1   g18183(.A1(new_n21222_), .A2(new_n11868_), .B(new_n21224_), .ZN(new_n21225_));
  NAND2_X1   g18184(.A1(new_n21225_), .A2(new_n21223_), .ZN(new_n21226_));
  NOR4_X1    g18185(.A1(new_n21207_), .A2(new_n12031_), .A3(pi1156), .A4(new_n21069_), .ZN(new_n21227_));
  NOR2_X1    g18186(.A1(new_n21227_), .A2(new_n21208_), .ZN(new_n21228_));
  MUX2_X1    g18187(.I0(new_n21228_), .I1(new_n21207_), .S(new_n11868_), .Z(new_n21229_));
  NAND2_X1   g18188(.A1(new_n21229_), .A2(pi0647), .ZN(new_n21230_));
  AOI21_X1   g18189(.A1(new_n21069_), .A2(pi0647), .B(pi1157), .ZN(new_n21231_));
  NAND2_X1   g18190(.A1(new_n21230_), .A2(new_n21231_), .ZN(new_n21232_));
  NOR2_X1    g18191(.A1(new_n21069_), .A2(new_n12054_), .ZN(new_n21233_));
  AOI21_X1   g18192(.A1(new_n21204_), .A2(new_n12054_), .B(new_n21233_), .ZN(new_n21234_));
  NOR2_X1    g18193(.A1(new_n12061_), .A2(pi1157), .ZN(new_n21235_));
  OAI21_X1   g18194(.A1(new_n21232_), .A2(new_n12060_), .B(new_n21235_), .ZN(new_n21236_));
  NOR3_X1    g18195(.A1(new_n21217_), .A2(new_n11868_), .A3(new_n21224_), .ZN(new_n21237_));
  AOI21_X1   g18196(.A1(new_n21217_), .A2(pi0792), .B(new_n21201_), .ZN(new_n21238_));
  NOR3_X1    g18197(.A1(new_n21237_), .A2(new_n21238_), .A3(pi0647), .ZN(new_n21239_));
  AOI21_X1   g18198(.A1(new_n21087_), .A2(new_n12061_), .B(pi1157), .ZN(new_n21240_));
  NAND2_X1   g18199(.A1(new_n21230_), .A2(new_n21240_), .ZN(new_n21241_));
  NAND2_X1   g18200(.A1(new_n21241_), .A2(new_n12060_), .ZN(new_n21242_));
  AOI21_X1   g18201(.A1(new_n21234_), .A2(pi0647), .B(pi1157), .ZN(new_n21243_));
  AND2_X2    g18202(.A1(new_n21243_), .A2(new_n21242_), .Z(new_n21244_));
  INV_X1     g18203(.I(new_n21244_), .ZN(new_n21245_));
  OAI22_X1   g18204(.A1(new_n21239_), .A2(new_n21245_), .B1(new_n21226_), .B2(new_n21236_), .ZN(new_n21246_));
  MUX2_X1    g18205(.I0(new_n21246_), .I1(new_n21218_), .S(new_n12048_), .Z(new_n21247_));
  INV_X1     g18206(.I(new_n21229_), .ZN(new_n21248_));
  NOR3_X1    g18207(.A1(new_n21069_), .A2(pi0647), .A3(pi1157), .ZN(new_n21249_));
  MUX2_X1    g18208(.I0(new_n21249_), .I1(new_n21248_), .S(new_n12048_), .Z(new_n21250_));
  NAND2_X1   g18209(.A1(new_n21250_), .A2(pi0644), .ZN(new_n21251_));
  NOR2_X1    g18210(.A1(new_n21087_), .A2(new_n12092_), .ZN(new_n21252_));
  AOI21_X1   g18211(.A1(new_n21234_), .A2(new_n12092_), .B(new_n21252_), .ZN(new_n21253_));
  NAND2_X1   g18212(.A1(new_n12082_), .A2(new_n12099_), .ZN(new_n21254_));
  OR2_X2     g18213(.A1(new_n21253_), .A2(new_n21254_), .Z(new_n21255_));
  NAND3_X1   g18214(.A1(new_n21255_), .A2(new_n21251_), .A3(new_n13168_), .ZN(new_n21256_));
  AOI21_X1   g18215(.A1(new_n21247_), .A2(new_n12082_), .B(new_n21256_), .ZN(new_n21257_));
  INV_X1     g18216(.I(new_n21236_), .ZN(new_n21258_));
  NAND3_X1   g18217(.A1(new_n21225_), .A2(new_n21223_), .A3(new_n12061_), .ZN(new_n21259_));
  AOI22_X1   g18218(.A1(new_n21259_), .A2(new_n21244_), .B1(new_n21218_), .B2(new_n21258_), .ZN(new_n21260_));
  MUX2_X1    g18219(.I0(new_n21260_), .I1(new_n21226_), .S(new_n12048_), .Z(new_n21261_));
  NAND3_X1   g18220(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n21262_));
  OAI21_X1   g18221(.A1(new_n21253_), .A2(new_n21262_), .B(new_n13179_), .ZN(new_n21263_));
  NOR2_X1    g18222(.A1(new_n21263_), .A2(new_n21250_), .ZN(new_n21264_));
  OAI21_X1   g18223(.A1(new_n21261_), .A2(new_n12082_), .B(new_n21264_), .ZN(new_n21265_));
  NOR2_X1    g18224(.A1(new_n21257_), .A2(new_n21265_), .ZN(new_n21266_));
  NAND2_X1   g18225(.A1(po1038), .A2(new_n7356_), .ZN(new_n21267_));
  AOI21_X1   g18226(.A1(new_n21267_), .A2(new_n13184_), .B(po1038), .ZN(new_n21268_));
  OAI21_X1   g18227(.A1(new_n21247_), .A2(pi0790), .B(new_n21268_), .ZN(new_n21269_));
  OAI21_X1   g18228(.A1(new_n21266_), .A2(new_n21269_), .B(new_n21046_), .ZN(po0345));
  NOR2_X1    g18229(.A1(new_n2925_), .A2(new_n8872_), .ZN(new_n21271_));
  NOR2_X1    g18230(.A1(new_n11894_), .A2(new_n16128_), .ZN(new_n21272_));
  NOR2_X1    g18231(.A1(new_n21272_), .A2(new_n21271_), .ZN(new_n21273_));
  INV_X1     g18232(.I(new_n21273_), .ZN(new_n21274_));
  INV_X1     g18233(.I(new_n21272_), .ZN(new_n21275_));
  NOR3_X1    g18234(.A1(new_n21275_), .A2(new_n13659_), .A3(new_n21271_), .ZN(new_n21276_));
  INV_X1     g18235(.I(new_n21271_), .ZN(new_n21277_));
  NOR3_X1    g18236(.A1(new_n21272_), .A2(new_n12970_), .A3(new_n21277_), .ZN(new_n21278_));
  AOI21_X1   g18237(.A1(new_n21275_), .A2(new_n21277_), .B(pi0625), .ZN(new_n21279_));
  NOR3_X1    g18238(.A1(new_n21279_), .A2(pi1153), .A3(new_n21278_), .ZN(new_n21280_));
  INV_X1     g18239(.I(new_n21280_), .ZN(new_n21281_));
  NOR2_X1    g18240(.A1(new_n21281_), .A2(new_n21276_), .ZN(new_n21282_));
  MUX2_X1    g18241(.I0(new_n21282_), .I1(new_n21274_), .S(new_n11891_), .Z(new_n21283_));
  NOR2_X1    g18242(.A1(new_n21283_), .A2(new_n13717_), .ZN(new_n21284_));
  INV_X1     g18243(.I(new_n21284_), .ZN(new_n21285_));
  NOR2_X1    g18244(.A1(new_n21285_), .A2(new_n12066_), .ZN(new_n21286_));
  AOI21_X1   g18245(.A1(new_n21286_), .A2(new_n13748_), .B(new_n21271_), .ZN(new_n21287_));
  INV_X1     g18246(.I(new_n21287_), .ZN(new_n21288_));
  NOR2_X1    g18247(.A1(new_n11877_), .A2(new_n16129_), .ZN(new_n21289_));
  INV_X1     g18248(.I(new_n21289_), .ZN(new_n21290_));
  NOR2_X1    g18249(.A1(new_n21290_), .A2(new_n14627_), .ZN(new_n21291_));
  INV_X1     g18250(.I(new_n21291_), .ZN(new_n21292_));
  NOR2_X1    g18251(.A1(new_n21292_), .A2(new_n14644_), .ZN(new_n21293_));
  INV_X1     g18252(.I(new_n21293_), .ZN(new_n21294_));
  NOR2_X1    g18253(.A1(new_n21294_), .A2(new_n11997_), .ZN(new_n21295_));
  AOI21_X1   g18254(.A1(new_n21295_), .A2(new_n16762_), .B(new_n12061_), .ZN(new_n21296_));
  OAI21_X1   g18255(.A1(new_n21286_), .A2(pi0630), .B(new_n21296_), .ZN(new_n21297_));
  OAI22_X1   g18256(.A1(new_n21286_), .A2(new_n12060_), .B1(new_n16765_), .B2(new_n21295_), .ZN(new_n21298_));
  NAND2_X1   g18257(.A1(new_n21298_), .A2(new_n12049_), .ZN(new_n21299_));
  NAND2_X1   g18258(.A1(new_n21299_), .A2(new_n21297_), .ZN(new_n21300_));
  NOR2_X1    g18259(.A1(new_n21271_), .A2(new_n12048_), .ZN(new_n21301_));
  NOR4_X1    g18260(.A1(new_n21285_), .A2(new_n12031_), .A3(pi0629), .A4(pi1156), .ZN(new_n21302_));
  INV_X1     g18261(.I(new_n21295_), .ZN(new_n21303_));
  OAI21_X1   g18262(.A1(new_n21303_), .A2(pi0629), .B(pi0628), .ZN(new_n21304_));
  NAND2_X1   g18263(.A1(new_n21285_), .A2(pi0629), .ZN(new_n21305_));
  AOI21_X1   g18264(.A1(new_n21305_), .A2(new_n21304_), .B(pi1156), .ZN(new_n21306_));
  NOR2_X1    g18265(.A1(new_n21271_), .A2(new_n11868_), .ZN(new_n21307_));
  OAI21_X1   g18266(.A1(new_n21306_), .A2(new_n21302_), .B(new_n21307_), .ZN(new_n21308_));
  INV_X1     g18267(.I(new_n21283_), .ZN(new_n21309_));
  AOI21_X1   g18268(.A1(new_n21309_), .A2(new_n11938_), .B(new_n21271_), .ZN(new_n21310_));
  INV_X1     g18269(.I(new_n21310_), .ZN(new_n21311_));
  NAND2_X1   g18270(.A1(new_n12118_), .A2(pi0727), .ZN(new_n21312_));
  AND3_X2    g18271(.A1(new_n21312_), .A2(new_n21277_), .A3(new_n21290_), .Z(new_n21313_));
  NOR2_X1    g18272(.A1(new_n13649_), .A2(new_n16128_), .ZN(new_n21314_));
  NAND3_X1   g18273(.A1(new_n21290_), .A2(pi1153), .A3(new_n21277_), .ZN(new_n21315_));
  OAI21_X1   g18274(.A1(new_n21314_), .A2(new_n21315_), .B(pi0608), .ZN(new_n21316_));
  INV_X1     g18275(.I(new_n21313_), .ZN(new_n21317_));
  NOR2_X1    g18276(.A1(new_n21317_), .A2(new_n21314_), .ZN(new_n21318_));
  OAI21_X1   g18277(.A1(new_n21276_), .A2(pi0608), .B(new_n11893_), .ZN(new_n21319_));
  OAI22_X1   g18278(.A1(new_n21281_), .A2(new_n21316_), .B1(new_n21318_), .B2(new_n21319_), .ZN(new_n21320_));
  MUX2_X1    g18279(.I0(new_n21320_), .I1(new_n21313_), .S(new_n11891_), .Z(new_n21321_));
  NOR3_X1    g18280(.A1(new_n21283_), .A2(new_n11903_), .A3(new_n11912_), .ZN(new_n21322_));
  NOR4_X1    g18281(.A1(new_n21290_), .A2(pi1155), .A3(new_n13010_), .A4(new_n21271_), .ZN(new_n21323_));
  NOR3_X1    g18282(.A1(new_n21322_), .A2(pi0660), .A3(new_n21323_), .ZN(new_n21324_));
  NOR4_X1    g18283(.A1(new_n21321_), .A2(new_n11903_), .A3(pi1155), .A4(new_n21309_), .ZN(new_n21325_));
  NOR2_X1    g18284(.A1(new_n21271_), .A2(new_n14671_), .ZN(new_n21326_));
  OAI21_X1   g18285(.A1(new_n21290_), .A2(new_n12997_), .B(new_n21326_), .ZN(new_n21327_));
  OAI21_X1   g18286(.A1(new_n21325_), .A2(new_n21327_), .B(pi0785), .ZN(new_n21328_));
  OAI22_X1   g18287(.A1(new_n21328_), .A2(new_n21324_), .B1(pi0785), .B2(new_n21321_), .ZN(new_n21329_));
  XOR2_X1    g18288(.A1(new_n21329_), .A2(new_n21311_), .Z(new_n21330_));
  NOR2_X1    g18289(.A1(new_n21330_), .A2(new_n11934_), .ZN(new_n21331_));
  XOR2_X1    g18290(.A1(new_n21331_), .A2(new_n21311_), .Z(new_n21332_));
  NOR2_X1    g18291(.A1(new_n21332_), .A2(new_n11950_), .ZN(new_n21333_));
  NOR2_X1    g18292(.A1(new_n21271_), .A2(pi1154), .ZN(new_n21334_));
  OAI21_X1   g18293(.A1(new_n21292_), .A2(new_n14686_), .B(new_n21334_), .ZN(new_n21335_));
  OAI21_X1   g18294(.A1(new_n21333_), .A2(new_n21335_), .B(new_n11949_), .ZN(new_n21336_));
  XOR2_X1    g18295(.A1(new_n21331_), .A2(new_n21329_), .Z(new_n21337_));
  NAND2_X1   g18296(.A1(new_n21337_), .A2(new_n11950_), .ZN(new_n21338_));
  NOR4_X1    g18297(.A1(new_n11914_), .A2(new_n11934_), .A3(pi1154), .A4(new_n21271_), .ZN(new_n21339_));
  AOI21_X1   g18298(.A1(new_n21291_), .A2(new_n21339_), .B(pi0627), .ZN(new_n21340_));
  AOI21_X1   g18299(.A1(new_n21338_), .A2(new_n21340_), .B(new_n11969_), .ZN(new_n21341_));
  OAI21_X1   g18300(.A1(new_n21329_), .A2(pi0781), .B(new_n16811_), .ZN(new_n21342_));
  AOI21_X1   g18301(.A1(new_n21336_), .A2(new_n21341_), .B(new_n21342_), .ZN(new_n21343_));
  NOR2_X1    g18302(.A1(new_n21283_), .A2(new_n13716_), .ZN(new_n21344_));
  AOI21_X1   g18303(.A1(new_n21291_), .A2(new_n14697_), .B(pi0648), .ZN(new_n21345_));
  OAI21_X1   g18304(.A1(new_n21292_), .A2(new_n16816_), .B(pi0648), .ZN(new_n21346_));
  NAND2_X1   g18305(.A1(new_n21346_), .A2(new_n12012_), .ZN(new_n21347_));
  NOR4_X1    g18306(.A1(new_n14640_), .A2(new_n16809_), .A3(new_n21271_), .A4(pi0789), .ZN(new_n21348_));
  OAI21_X1   g18307(.A1(new_n21347_), .A2(new_n21345_), .B(new_n21348_), .ZN(new_n21349_));
  NOR2_X1    g18308(.A1(new_n21344_), .A2(new_n21349_), .ZN(new_n21350_));
  AOI21_X1   g18309(.A1(new_n21344_), .A2(new_n12014_), .B(new_n21271_), .ZN(new_n21351_));
  OAI21_X1   g18310(.A1(new_n21294_), .A2(pi0626), .B(new_n21277_), .ZN(new_n21352_));
  NAND2_X1   g18311(.A1(new_n21352_), .A2(new_n11987_), .ZN(new_n21353_));
  NAND4_X1   g18312(.A1(new_n21351_), .A2(new_n11989_), .A3(new_n16822_), .A4(new_n21353_), .ZN(new_n21354_));
  NAND2_X1   g18313(.A1(new_n21351_), .A2(new_n16827_), .ZN(new_n21355_));
  OAI21_X1   g18314(.A1(new_n21294_), .A2(new_n11994_), .B(new_n21277_), .ZN(new_n21356_));
  NAND2_X1   g18315(.A1(new_n21356_), .A2(pi1158), .ZN(new_n21357_));
  NAND4_X1   g18316(.A1(new_n21354_), .A2(new_n11989_), .A3(new_n21355_), .A4(new_n21357_), .ZN(new_n21358_));
  AOI21_X1   g18317(.A1(new_n21358_), .A2(new_n11986_), .B(new_n16832_), .ZN(new_n21359_));
  OAI21_X1   g18318(.A1(new_n21343_), .A2(new_n21350_), .B(new_n21359_), .ZN(new_n21360_));
  NAND2_X1   g18319(.A1(new_n21360_), .A2(new_n21308_), .ZN(new_n21361_));
  AOI22_X1   g18320(.A1(new_n21361_), .A2(new_n14726_), .B1(new_n21300_), .B2(new_n21301_), .ZN(new_n21362_));
  NOR3_X1    g18321(.A1(new_n21362_), .A2(pi0644), .A3(new_n21288_), .ZN(new_n21363_));
  AOI21_X1   g18322(.A1(new_n21362_), .A2(new_n12082_), .B(new_n21287_), .ZN(new_n21364_));
  NOR4_X1    g18323(.A1(new_n21303_), .A2(new_n14740_), .A3(new_n16841_), .A4(new_n21271_), .ZN(new_n21365_));
  NOR4_X1    g18324(.A1(new_n21363_), .A2(new_n21364_), .A3(new_n13169_), .A4(new_n21365_), .ZN(new_n21366_));
  NOR3_X1    g18325(.A1(new_n21303_), .A2(new_n12082_), .A3(new_n16841_), .ZN(new_n21367_));
  NOR3_X1    g18326(.A1(new_n21367_), .A2(pi0715), .A3(new_n21271_), .ZN(new_n21368_));
  OAI21_X1   g18327(.A1(new_n21368_), .A2(pi1160), .B(pi0790), .ZN(new_n21369_));
  AND2_X2    g18328(.A1(new_n21362_), .A2(new_n14747_), .Z(new_n21370_));
  OAI21_X1   g18329(.A1(new_n21366_), .A2(new_n21369_), .B(new_n21370_), .ZN(new_n21371_));
  NOR2_X1    g18330(.A1(new_n11875_), .A2(new_n16129_), .ZN(new_n21372_));
  INV_X1     g18331(.I(new_n21372_), .ZN(new_n21373_));
  NOR3_X1    g18332(.A1(new_n13368_), .A2(pi0189), .A3(new_n21373_), .ZN(new_n21374_));
  AOI21_X1   g18333(.A1(new_n12828_), .A2(new_n21373_), .B(new_n8872_), .ZN(new_n21375_));
  OAI21_X1   g18334(.A1(new_n21374_), .A2(new_n21375_), .B(pi0038), .ZN(new_n21376_));
  NAND2_X1   g18335(.A1(new_n8872_), .A2(pi0772), .ZN(new_n21377_));
  NAND2_X1   g18336(.A1(new_n12793_), .A2(new_n16129_), .ZN(new_n21378_));
  AOI21_X1   g18337(.A1(new_n12823_), .A2(pi0772), .B(new_n3154_), .ZN(new_n21379_));
  OAI21_X1   g18338(.A1(pi0772), .A2(new_n12852_), .B(new_n13346_), .ZN(new_n21380_));
  NAND3_X1   g18339(.A1(new_n12664_), .A2(new_n16129_), .A3(new_n12852_), .ZN(new_n21381_));
  NAND3_X1   g18340(.A1(new_n21380_), .A2(new_n21381_), .A3(new_n3154_), .ZN(new_n21382_));
  AOI21_X1   g18341(.A1(new_n21378_), .A2(new_n21379_), .B(new_n21382_), .ZN(new_n21383_));
  OAI22_X1   g18342(.A1(new_n21383_), .A2(new_n8872_), .B1(new_n12694_), .B2(new_n21377_), .ZN(new_n21384_));
  NAND2_X1   g18343(.A1(new_n21384_), .A2(new_n3172_), .ZN(new_n21385_));
  NAND2_X1   g18344(.A1(new_n21385_), .A2(new_n21376_), .ZN(new_n21386_));
  NAND2_X1   g18345(.A1(new_n12277_), .A2(new_n8872_), .ZN(new_n21387_));
  NOR4_X1    g18346(.A1(new_n12349_), .A2(pi0039), .A3(pi0189), .A4(pi0772), .ZN(new_n21388_));
  NAND2_X1   g18347(.A1(pi0189), .A2(pi0772), .ZN(new_n21389_));
  AOI21_X1   g18348(.A1(new_n21387_), .A2(new_n21388_), .B(new_n21389_), .ZN(new_n21390_));
  NAND2_X1   g18349(.A1(new_n21390_), .A2(new_n13332_), .ZN(new_n21391_));
  AOI21_X1   g18350(.A1(new_n13362_), .A2(pi0189), .B(pi0772), .ZN(new_n21392_));
  OAI21_X1   g18351(.A1(pi0189), .A2(new_n13360_), .B(new_n21392_), .ZN(new_n21393_));
  NOR4_X1    g18352(.A1(new_n12668_), .A2(new_n8872_), .A3(pi0772), .A4(new_n13347_), .ZN(new_n21394_));
  NOR2_X1    g18353(.A1(new_n21394_), .A2(pi0039), .ZN(new_n21395_));
  NAND3_X1   g18354(.A1(new_n21376_), .A2(pi0727), .A3(new_n14352_), .ZN(new_n21396_));
  NAND2_X1   g18355(.A1(new_n21396_), .A2(new_n14778_), .ZN(new_n21397_));
  AOI21_X1   g18356(.A1(new_n21393_), .A2(new_n21395_), .B(new_n21397_), .ZN(new_n21398_));
  AOI21_X1   g18357(.A1(new_n21398_), .A2(new_n21391_), .B(pi0727), .ZN(new_n21399_));
  AOI22_X1   g18358(.A1(new_n21386_), .A2(new_n21399_), .B1(pi0189), .B2(new_n3232_), .ZN(new_n21400_));
  INV_X1     g18359(.I(new_n21400_), .ZN(new_n21401_));
  NOR2_X1    g18360(.A1(new_n3231_), .A2(pi0189), .ZN(new_n21402_));
  AOI21_X1   g18361(.A1(new_n21386_), .A2(new_n3231_), .B(new_n21402_), .ZN(new_n21403_));
  AOI21_X1   g18362(.A1(new_n21403_), .A2(new_n12970_), .B(pi1153), .ZN(new_n21404_));
  OAI21_X1   g18363(.A1(new_n12970_), .A2(new_n21401_), .B(new_n21404_), .ZN(new_n21405_));
  NAND3_X1   g18364(.A1(new_n14382_), .A2(new_n8872_), .A3(new_n13395_), .ZN(new_n21406_));
  OAI21_X1   g18365(.A1(pi0189), .A2(new_n13395_), .B(new_n13399_), .ZN(new_n21407_));
  NOR3_X1    g18366(.A1(new_n3232_), .A2(pi0038), .A3(new_n16128_), .ZN(new_n21410_));
  AND3_X2    g18367(.A1(new_n21406_), .A2(new_n21407_), .A3(new_n21410_), .Z(new_n21411_));
  AOI22_X1   g18368(.A1(new_n14396_), .A2(pi0189), .B1(pi0727), .B2(new_n3231_), .ZN(new_n21412_));
  NOR2_X1    g18369(.A1(new_n21411_), .A2(new_n21412_), .ZN(new_n21413_));
  INV_X1     g18370(.I(new_n21413_), .ZN(new_n21414_));
  NAND2_X1   g18371(.A1(new_n14396_), .A2(pi0189), .ZN(new_n21415_));
  NAND2_X1   g18372(.A1(new_n21415_), .A2(pi0625), .ZN(new_n21416_));
  NAND2_X1   g18373(.A1(new_n21416_), .A2(new_n11893_), .ZN(new_n21417_));
  AOI21_X1   g18374(.A1(new_n21414_), .A2(new_n12970_), .B(new_n21417_), .ZN(new_n21418_));
  NOR2_X1    g18375(.A1(new_n21418_), .A2(new_n13657_), .ZN(new_n21419_));
  NAND2_X1   g18376(.A1(new_n21413_), .A2(pi0625), .ZN(new_n21420_));
  AOI21_X1   g18377(.A1(new_n21420_), .A2(new_n21416_), .B(new_n11893_), .ZN(new_n21421_));
  INV_X1     g18378(.I(new_n21421_), .ZN(new_n21422_));
  OAI21_X1   g18379(.A1(new_n21403_), .A2(new_n12970_), .B(new_n12977_), .ZN(new_n21423_));
  AOI21_X1   g18380(.A1(pi0625), .A2(new_n21400_), .B(new_n21423_), .ZN(new_n21424_));
  AOI22_X1   g18381(.A1(new_n21422_), .A2(new_n21424_), .B1(new_n21419_), .B2(new_n21405_), .ZN(new_n21425_));
  MUX2_X1    g18382(.I0(new_n21425_), .I1(new_n21400_), .S(new_n11891_), .Z(new_n21426_));
  INV_X1     g18383(.I(new_n21426_), .ZN(new_n21427_));
  NOR2_X1    g18384(.A1(new_n21427_), .A2(pi0785), .ZN(new_n21428_));
  INV_X1     g18385(.I(new_n21428_), .ZN(new_n21429_));
  NOR2_X1    g18386(.A1(new_n21421_), .A2(new_n21418_), .ZN(new_n21430_));
  MUX2_X1    g18387(.I0(new_n21430_), .I1(new_n21414_), .S(new_n11891_), .Z(new_n21431_));
  OAI21_X1   g18388(.A1(new_n21431_), .A2(pi0609), .B(pi1155), .ZN(new_n21432_));
  NOR2_X1    g18389(.A1(new_n21415_), .A2(new_n11924_), .ZN(new_n21433_));
  AOI21_X1   g18390(.A1(new_n21403_), .A2(new_n11924_), .B(new_n21433_), .ZN(new_n21434_));
  INV_X1     g18391(.I(new_n21434_), .ZN(new_n21435_));
  NOR3_X1    g18392(.A1(new_n21435_), .A2(new_n11903_), .A3(new_n21415_), .ZN(new_n21436_));
  AOI21_X1   g18393(.A1(pi0609), .A2(new_n21415_), .B(new_n21434_), .ZN(new_n21437_));
  OAI21_X1   g18394(.A1(new_n21436_), .A2(new_n21437_), .B(new_n11912_), .ZN(new_n21438_));
  NAND2_X1   g18395(.A1(new_n21438_), .A2(pi0660), .ZN(new_n21439_));
  AND3_X2    g18396(.A1(new_n21426_), .A2(pi0609), .A3(new_n21439_), .Z(new_n21440_));
  NOR2_X1    g18397(.A1(new_n12965_), .A2(new_n8872_), .ZN(new_n21441_));
  NOR3_X1    g18398(.A1(new_n21434_), .A2(new_n11903_), .A3(new_n21441_), .ZN(new_n21442_));
  AOI21_X1   g18399(.A1(new_n21434_), .A2(pi0609), .B(new_n21415_), .ZN(new_n21443_));
  NOR2_X1    g18400(.A1(new_n11923_), .A2(pi1155), .ZN(new_n21444_));
  OAI21_X1   g18401(.A1(new_n21431_), .A2(new_n11903_), .B(new_n21444_), .ZN(new_n21445_));
  AOI21_X1   g18402(.A1(new_n21426_), .A2(new_n11903_), .B(new_n21445_), .ZN(new_n21446_));
  AOI21_X1   g18403(.A1(new_n21440_), .A2(new_n21432_), .B(new_n21446_), .ZN(new_n21447_));
  NOR3_X1    g18404(.A1(new_n21447_), .A2(new_n11870_), .A3(new_n21429_), .ZN(new_n21448_));
  NAND4_X1   g18405(.A1(new_n21426_), .A2(pi0609), .A3(new_n21432_), .A4(new_n21439_), .ZN(new_n21449_));
  NOR2_X1    g18406(.A1(new_n21427_), .A2(pi0609), .ZN(new_n21450_));
  OAI21_X1   g18407(.A1(new_n21450_), .A2(new_n21445_), .B(new_n21449_), .ZN(new_n21451_));
  AOI21_X1   g18408(.A1(new_n21451_), .A2(pi0785), .B(new_n21428_), .ZN(new_n21452_));
  NOR2_X1    g18409(.A1(new_n21448_), .A2(new_n21452_), .ZN(new_n21453_));
  NAND2_X1   g18410(.A1(new_n21453_), .A2(new_n11969_), .ZN(new_n21454_));
  OAI21_X1   g18411(.A1(new_n21442_), .A2(new_n21443_), .B(pi1155), .ZN(new_n21455_));
  NAND2_X1   g18412(.A1(new_n21438_), .A2(new_n21455_), .ZN(new_n21456_));
  MUX2_X1    g18413(.I0(new_n21456_), .I1(new_n21435_), .S(new_n11870_), .Z(new_n21457_));
  NAND3_X1   g18414(.A1(new_n21457_), .A2(new_n11934_), .A3(new_n21441_), .ZN(new_n21458_));
  OAI21_X1   g18415(.A1(new_n21457_), .A2(pi0618), .B(new_n21415_), .ZN(new_n21459_));
  NAND3_X1   g18416(.A1(new_n21459_), .A2(new_n21458_), .A3(new_n11950_), .ZN(new_n21460_));
  NOR2_X1    g18417(.A1(new_n21460_), .A2(new_n11949_), .ZN(new_n21461_));
  INV_X1     g18418(.I(new_n21461_), .ZN(new_n21462_));
  NOR2_X1    g18419(.A1(new_n21415_), .A2(new_n11938_), .ZN(new_n21463_));
  AOI21_X1   g18420(.A1(new_n21431_), .A2(new_n11938_), .B(new_n21463_), .ZN(new_n21464_));
  NOR4_X1    g18421(.A1(new_n21448_), .A2(new_n21452_), .A3(new_n11934_), .A4(pi1154), .ZN(new_n21465_));
  NAND3_X1   g18422(.A1(new_n21451_), .A2(pi0785), .A3(new_n21428_), .ZN(new_n21466_));
  OAI21_X1   g18423(.A1(new_n21447_), .A2(new_n11870_), .B(new_n21429_), .ZN(new_n21467_));
  NAND3_X1   g18424(.A1(new_n21467_), .A2(new_n21466_), .A3(new_n11934_), .ZN(new_n21468_));
  AOI21_X1   g18425(.A1(new_n21464_), .A2(pi0618), .B(new_n14687_), .ZN(new_n21469_));
  AOI22_X1   g18426(.A1(new_n21465_), .A2(new_n21462_), .B1(new_n21468_), .B2(new_n21469_), .ZN(new_n21470_));
  NOR3_X1    g18427(.A1(new_n21470_), .A2(new_n11969_), .A3(new_n21454_), .ZN(new_n21471_));
  INV_X1     g18428(.I(new_n21454_), .ZN(new_n21472_));
  NAND4_X1   g18429(.A1(new_n21467_), .A2(new_n21466_), .A3(pi0618), .A4(new_n11950_), .ZN(new_n21473_));
  NOR3_X1    g18430(.A1(new_n21448_), .A2(new_n21452_), .A3(pi0618), .ZN(new_n21474_));
  INV_X1     g18431(.I(new_n21469_), .ZN(new_n21475_));
  OAI22_X1   g18432(.A1(new_n21461_), .A2(new_n21473_), .B1(new_n21474_), .B2(new_n21475_), .ZN(new_n21476_));
  AOI21_X1   g18433(.A1(new_n21476_), .A2(pi0781), .B(new_n21472_), .ZN(new_n21477_));
  NOR3_X1    g18434(.A1(new_n21477_), .A2(new_n21471_), .A3(pi0789), .ZN(new_n21478_));
  INV_X1     g18435(.I(new_n21457_), .ZN(new_n21479_));
  MUX2_X1    g18436(.I0(new_n21460_), .I1(new_n21479_), .S(new_n11969_), .Z(new_n21480_));
  NOR3_X1    g18437(.A1(new_n21480_), .A2(pi0619), .A3(new_n21415_), .ZN(new_n21481_));
  AOI21_X1   g18438(.A1(new_n21480_), .A2(new_n11967_), .B(new_n21441_), .ZN(new_n21482_));
  NOR3_X1    g18439(.A1(new_n21481_), .A2(new_n21482_), .A3(pi1159), .ZN(new_n21483_));
  NAND2_X1   g18440(.A1(new_n21483_), .A2(pi0648), .ZN(new_n21484_));
  INV_X1     g18441(.I(new_n21484_), .ZN(new_n21485_));
  NAND3_X1   g18442(.A1(new_n21476_), .A2(new_n21472_), .A3(pi0781), .ZN(new_n21486_));
  OAI21_X1   g18443(.A1(new_n21470_), .A2(new_n11969_), .B(new_n21454_), .ZN(new_n21487_));
  NOR2_X1    g18444(.A1(new_n21441_), .A2(new_n11961_), .ZN(new_n21488_));
  AOI21_X1   g18445(.A1(new_n21464_), .A2(new_n11961_), .B(new_n21488_), .ZN(new_n21489_));
  NAND4_X1   g18446(.A1(new_n21486_), .A2(new_n21487_), .A3(pi0619), .A4(new_n11869_), .ZN(new_n21490_));
  NOR3_X1    g18447(.A1(new_n21477_), .A2(new_n21471_), .A3(pi0619), .ZN(new_n21491_));
  INV_X1     g18448(.I(new_n21489_), .ZN(new_n21492_));
  AOI21_X1   g18449(.A1(new_n21492_), .A2(pi0619), .B(new_n14904_), .ZN(new_n21493_));
  INV_X1     g18450(.I(new_n21493_), .ZN(new_n21494_));
  OAI22_X1   g18451(.A1(new_n21491_), .A2(new_n21494_), .B1(new_n21490_), .B2(new_n21485_), .ZN(new_n21495_));
  NAND3_X1   g18452(.A1(new_n21495_), .A2(pi0789), .A3(new_n21478_), .ZN(new_n21496_));
  INV_X1     g18453(.I(new_n21478_), .ZN(new_n21497_));
  NOR4_X1    g18454(.A1(new_n21477_), .A2(new_n21471_), .A3(new_n11967_), .A4(pi1159), .ZN(new_n21498_));
  NAND3_X1   g18455(.A1(new_n21486_), .A2(new_n21487_), .A3(new_n11967_), .ZN(new_n21499_));
  AOI22_X1   g18456(.A1(new_n21498_), .A2(new_n21484_), .B1(new_n21499_), .B2(new_n21493_), .ZN(new_n21500_));
  OAI21_X1   g18457(.A1(new_n21500_), .A2(new_n11985_), .B(new_n21497_), .ZN(new_n21501_));
  NAND2_X1   g18458(.A1(new_n21496_), .A2(new_n21501_), .ZN(new_n21502_));
  NOR3_X1    g18459(.A1(new_n21500_), .A2(new_n11985_), .A3(new_n21497_), .ZN(new_n21503_));
  AOI21_X1   g18460(.A1(new_n21495_), .A2(pi0789), .B(new_n21478_), .ZN(new_n21504_));
  INV_X1     g18461(.I(new_n21480_), .ZN(new_n21505_));
  MUX2_X1    g18462(.I0(new_n21483_), .I1(new_n21505_), .S(new_n11985_), .Z(new_n21506_));
  INV_X1     g18463(.I(new_n21506_), .ZN(new_n21507_));
  NOR3_X1    g18464(.A1(new_n11994_), .A2(new_n11989_), .A3(pi1158), .ZN(new_n21508_));
  NOR2_X1    g18465(.A1(new_n21415_), .A2(new_n12014_), .ZN(new_n21509_));
  AOI21_X1   g18466(.A1(new_n21489_), .A2(new_n12014_), .B(new_n21509_), .ZN(new_n21510_));
  NOR2_X1    g18467(.A1(new_n11994_), .A2(pi0641), .ZN(new_n21511_));
  INV_X1     g18468(.I(new_n21511_), .ZN(new_n21512_));
  AOI21_X1   g18469(.A1(new_n21507_), .A2(new_n21508_), .B(new_n21512_), .ZN(new_n21513_));
  INV_X1     g18470(.I(new_n21483_), .ZN(new_n21514_));
  NOR2_X1    g18471(.A1(new_n21505_), .A2(pi0789), .ZN(new_n21515_));
  NAND3_X1   g18472(.A1(new_n21514_), .A2(pi0789), .A3(new_n21515_), .ZN(new_n21516_));
  INV_X1     g18473(.I(new_n21515_), .ZN(new_n21517_));
  OAI21_X1   g18474(.A1(new_n21483_), .A2(new_n11985_), .B(new_n21517_), .ZN(new_n21518_));
  NAND3_X1   g18475(.A1(new_n21516_), .A2(new_n11994_), .A3(new_n21518_), .ZN(new_n21519_));
  AOI21_X1   g18476(.A1(new_n21441_), .A2(pi0626), .B(new_n11989_), .ZN(new_n21520_));
  NOR3_X1    g18477(.A1(new_n11989_), .A2(pi0626), .A3(pi1158), .ZN(new_n21521_));
  INV_X1     g18478(.I(new_n21521_), .ZN(new_n21522_));
  AOI21_X1   g18479(.A1(new_n21519_), .A2(new_n21520_), .B(new_n21522_), .ZN(new_n21523_));
  OAI22_X1   g18480(.A1(new_n21504_), .A2(new_n21503_), .B1(new_n21513_), .B2(new_n21523_), .ZN(new_n21524_));
  NOR3_X1    g18481(.A1(new_n21524_), .A2(new_n11986_), .A3(new_n21502_), .ZN(new_n21525_));
  NOR2_X1    g18482(.A1(new_n21504_), .A2(new_n21503_), .ZN(new_n21526_));
  AOI21_X1   g18483(.A1(new_n21524_), .A2(pi0788), .B(new_n21526_), .ZN(new_n21527_));
  NOR2_X1    g18484(.A1(new_n21525_), .A2(new_n21527_), .ZN(new_n21528_));
  NAND2_X1   g18485(.A1(new_n21506_), .A2(new_n14624_), .ZN(new_n21529_));
  NAND2_X1   g18486(.A1(new_n21415_), .A2(new_n11997_), .ZN(new_n21530_));
  AOI21_X1   g18487(.A1(new_n21529_), .A2(new_n21530_), .B(pi0628), .ZN(new_n21531_));
  NOR2_X1    g18488(.A1(new_n21441_), .A2(new_n13114_), .ZN(new_n21532_));
  AOI21_X1   g18489(.A1(new_n21510_), .A2(new_n13114_), .B(new_n21532_), .ZN(new_n21533_));
  INV_X1     g18490(.I(new_n21533_), .ZN(new_n21534_));
  NAND3_X1   g18491(.A1(new_n21534_), .A2(new_n12031_), .A3(new_n21441_), .ZN(new_n21535_));
  OAI21_X1   g18492(.A1(new_n21534_), .A2(pi0628), .B(new_n21415_), .ZN(new_n21536_));
  NAND3_X1   g18493(.A1(new_n21536_), .A2(new_n21535_), .A3(new_n12026_), .ZN(new_n21537_));
  INV_X1     g18494(.I(new_n21537_), .ZN(new_n21538_));
  AOI21_X1   g18495(.A1(new_n21538_), .A2(pi0629), .B(new_n12031_), .ZN(new_n21539_));
  OAI21_X1   g18496(.A1(new_n21531_), .A2(new_n12026_), .B(new_n21539_), .ZN(new_n21540_));
  INV_X1     g18497(.I(new_n21540_), .ZN(new_n21541_));
  AND2_X2    g18498(.A1(new_n21529_), .A2(new_n21530_), .Z(new_n21542_));
  NOR3_X1    g18499(.A1(new_n12030_), .A2(new_n12026_), .A3(pi0628), .ZN(new_n21543_));
  OAI22_X1   g18500(.A1(new_n21525_), .A2(new_n21527_), .B1(new_n21541_), .B2(new_n21543_), .ZN(new_n21544_));
  MUX2_X1    g18501(.I0(new_n21544_), .I1(new_n21528_), .S(new_n11868_), .Z(new_n21545_));
  INV_X1     g18502(.I(new_n21545_), .ZN(new_n21546_));
  NAND2_X1   g18503(.A1(new_n21415_), .A2(new_n12053_), .ZN(new_n21547_));
  OAI21_X1   g18504(.A1(new_n21542_), .A2(new_n12053_), .B(new_n21547_), .ZN(new_n21548_));
  AOI21_X1   g18505(.A1(new_n21548_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n21549_));
  MUX2_X1    g18506(.I0(new_n21538_), .I1(new_n21534_), .S(new_n11868_), .Z(new_n21550_));
  NAND3_X1   g18507(.A1(new_n21550_), .A2(new_n12061_), .A3(new_n21441_), .ZN(new_n21551_));
  OAI21_X1   g18508(.A1(new_n21550_), .A2(pi0647), .B(new_n21415_), .ZN(new_n21552_));
  NAND3_X1   g18509(.A1(new_n21552_), .A2(new_n21551_), .A3(new_n12049_), .ZN(new_n21553_));
  NOR2_X1    g18510(.A1(new_n21553_), .A2(new_n12060_), .ZN(new_n21554_));
  NOR3_X1    g18511(.A1(new_n21549_), .A2(new_n12061_), .A3(new_n21554_), .ZN(new_n21555_));
  INV_X1     g18512(.I(new_n21513_), .ZN(new_n21556_));
  OAI21_X1   g18513(.A1(new_n21506_), .A2(pi0626), .B(new_n21520_), .ZN(new_n21557_));
  NAND2_X1   g18514(.A1(new_n21557_), .A2(new_n21521_), .ZN(new_n21558_));
  AOI22_X1   g18515(.A1(new_n21496_), .A2(new_n21501_), .B1(new_n21556_), .B2(new_n21558_), .ZN(new_n21559_));
  NAND3_X1   g18516(.A1(new_n21559_), .A2(pi0788), .A3(new_n21526_), .ZN(new_n21560_));
  OAI21_X1   g18517(.A1(new_n21559_), .A2(new_n11986_), .B(new_n21502_), .ZN(new_n21561_));
  AOI21_X1   g18518(.A1(new_n21561_), .A2(new_n21560_), .B(new_n21540_), .ZN(new_n21562_));
  NAND3_X1   g18519(.A1(new_n21562_), .A2(new_n21528_), .A3(pi0792), .ZN(new_n21563_));
  NAND2_X1   g18520(.A1(new_n21561_), .A2(new_n21560_), .ZN(new_n21564_));
  INV_X1     g18521(.I(new_n21543_), .ZN(new_n21565_));
  AOI22_X1   g18522(.A1(new_n21561_), .A2(new_n21560_), .B1(new_n21540_), .B2(new_n21565_), .ZN(new_n21566_));
  OAI21_X1   g18523(.A1(new_n21566_), .A2(new_n11868_), .B(new_n21564_), .ZN(new_n21567_));
  NAND3_X1   g18524(.A1(new_n21567_), .A2(new_n21563_), .A3(new_n12061_), .ZN(new_n21568_));
  AOI21_X1   g18525(.A1(new_n21548_), .A2(pi0647), .B(new_n13743_), .ZN(new_n21569_));
  AOI22_X1   g18526(.A1(new_n21568_), .A2(new_n21569_), .B1(new_n21545_), .B2(new_n21555_), .ZN(new_n21570_));
  MUX2_X1    g18527(.I0(new_n21570_), .I1(new_n21546_), .S(new_n12048_), .Z(new_n21571_));
  NOR2_X1    g18528(.A1(new_n21548_), .A2(new_n12091_), .ZN(new_n21572_));
  AOI21_X1   g18529(.A1(new_n12091_), .A2(new_n21441_), .B(new_n21572_), .ZN(new_n21573_));
  NAND2_X1   g18530(.A1(new_n21573_), .A2(new_n12082_), .ZN(new_n21574_));
  AOI21_X1   g18531(.A1(new_n21415_), .A2(pi0644), .B(new_n12099_), .ZN(new_n21575_));
  NOR2_X1    g18532(.A1(new_n21550_), .A2(pi0787), .ZN(new_n21576_));
  NAND2_X1   g18533(.A1(new_n21553_), .A2(pi0787), .ZN(new_n21577_));
  XNOR2_X1   g18534(.A1(new_n21577_), .A2(new_n21576_), .ZN(new_n21578_));
  OAI21_X1   g18535(.A1(new_n21578_), .A2(new_n12082_), .B(new_n13168_), .ZN(new_n21579_));
  AOI21_X1   g18536(.A1(new_n21574_), .A2(new_n21575_), .B(new_n21579_), .ZN(new_n21580_));
  OAI21_X1   g18537(.A1(new_n21571_), .A2(pi0644), .B(new_n21580_), .ZN(new_n21581_));
  NAND2_X1   g18538(.A1(new_n21545_), .A2(new_n12048_), .ZN(new_n21582_));
  OR3_X2     g18539(.A1(new_n21570_), .A2(new_n12048_), .A3(new_n21582_), .Z(new_n21583_));
  OAI21_X1   g18540(.A1(new_n21570_), .A2(new_n12048_), .B(new_n21582_), .ZN(new_n21584_));
  NOR3_X1    g18541(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n21585_));
  NAND2_X1   g18542(.A1(new_n21573_), .A2(new_n21585_), .ZN(new_n21586_));
  NOR2_X1    g18543(.A1(new_n12082_), .A2(pi0715), .ZN(new_n21587_));
  NAND4_X1   g18544(.A1(new_n21583_), .A2(new_n21584_), .A3(new_n21586_), .A4(new_n21587_), .ZN(new_n21588_));
  OAI21_X1   g18545(.A1(new_n21571_), .A2(new_n5223_), .B(new_n11867_), .ZN(new_n21589_));
  AOI21_X1   g18546(.A1(new_n21581_), .A2(new_n21588_), .B(new_n21589_), .ZN(new_n21590_));
  NAND2_X1   g18547(.A1(pi0057), .A2(pi0189), .ZN(new_n21591_));
  AOI21_X1   g18548(.A1(new_n21591_), .A2(new_n13184_), .B(pi0057), .ZN(new_n21592_));
  OAI21_X1   g18549(.A1(new_n5224_), .A2(pi0189), .B(new_n21592_), .ZN(new_n21593_));
  OAI21_X1   g18550(.A1(new_n21590_), .A2(new_n21593_), .B(new_n21371_), .ZN(po0346));
  NOR2_X1    g18551(.A1(new_n2925_), .A2(pi0190), .ZN(new_n21595_));
  NOR2_X1    g18552(.A1(new_n11877_), .A2(new_n16222_), .ZN(new_n21596_));
  NOR2_X1    g18553(.A1(new_n21596_), .A2(new_n21595_), .ZN(new_n21597_));
  AOI21_X1   g18554(.A1(new_n11886_), .A2(pi0699), .B(new_n21595_), .ZN(new_n21598_));
  NOR2_X1    g18555(.A1(new_n21598_), .A2(new_n11874_), .ZN(new_n21599_));
  INV_X1     g18556(.I(new_n21599_), .ZN(new_n21600_));
  NAND2_X1   g18557(.A1(new_n21600_), .A2(new_n21597_), .ZN(new_n21601_));
  NAND2_X1   g18558(.A1(new_n21601_), .A2(new_n11891_), .ZN(new_n21602_));
  NOR2_X1    g18559(.A1(new_n21600_), .A2(new_n12970_), .ZN(new_n21603_));
  NOR4_X1    g18560(.A1(new_n21603_), .A2(new_n11893_), .A3(new_n21595_), .A4(new_n21596_), .ZN(new_n21604_));
  NOR2_X1    g18561(.A1(new_n13201_), .A2(new_n16255_), .ZN(new_n21605_));
  NOR2_X1    g18562(.A1(new_n21595_), .A2(pi1153), .ZN(new_n21606_));
  INV_X1     g18563(.I(new_n21606_), .ZN(new_n21607_));
  NOR2_X1    g18564(.A1(new_n21605_), .A2(new_n21607_), .ZN(new_n21608_));
  INV_X1     g18565(.I(new_n21608_), .ZN(new_n21609_));
  NAND2_X1   g18566(.A1(new_n21609_), .A2(pi0608), .ZN(new_n21610_));
  INV_X1     g18567(.I(new_n21603_), .ZN(new_n21611_));
  AOI21_X1   g18568(.A1(new_n21611_), .A2(new_n21601_), .B(new_n21607_), .ZN(new_n21612_));
  OAI21_X1   g18569(.A1(new_n21605_), .A2(new_n21598_), .B(pi1153), .ZN(new_n21613_));
  NAND2_X1   g18570(.A1(new_n21613_), .A2(new_n13657_), .ZN(new_n21614_));
  OAI22_X1   g18571(.A1(new_n21610_), .A2(new_n21604_), .B1(new_n21612_), .B2(new_n21614_), .ZN(new_n21615_));
  NAND2_X1   g18572(.A1(new_n21615_), .A2(pi0778), .ZN(new_n21616_));
  XOR2_X1    g18573(.A1(new_n21616_), .A2(new_n21602_), .Z(new_n21617_));
  INV_X1     g18574(.I(new_n21617_), .ZN(new_n21618_));
  NAND2_X1   g18575(.A1(new_n21609_), .A2(new_n21613_), .ZN(new_n21619_));
  MUX2_X1    g18576(.I0(new_n21619_), .I1(new_n21598_), .S(new_n11891_), .Z(new_n21620_));
  XNOR2_X1   g18577(.A1(new_n21617_), .A2(new_n21620_), .ZN(new_n21621_));
  NAND2_X1   g18578(.A1(new_n21621_), .A2(pi0609), .ZN(new_n21622_));
  XOR2_X1    g18579(.A1(new_n21622_), .A2(new_n21618_), .Z(new_n21623_));
  INV_X1     g18580(.I(new_n21596_), .ZN(new_n21624_));
  NOR2_X1    g18581(.A1(new_n21597_), .A2(new_n11925_), .ZN(new_n21625_));
  NOR4_X1    g18582(.A1(new_n21625_), .A2(pi1155), .A3(new_n12997_), .A4(new_n21624_), .ZN(new_n21626_));
  NOR2_X1    g18583(.A1(new_n21626_), .A2(pi0660), .ZN(new_n21627_));
  OAI21_X1   g18584(.A1(new_n21623_), .A2(pi1155), .B(new_n21627_), .ZN(new_n21628_));
  NOR2_X1    g18585(.A1(new_n21624_), .A2(new_n12997_), .ZN(new_n21629_));
  NOR4_X1    g18586(.A1(new_n21629_), .A2(new_n11923_), .A3(pi1155), .A4(new_n21595_), .ZN(new_n21631_));
  NOR2_X1    g18587(.A1(new_n21631_), .A2(new_n11870_), .ZN(new_n21632_));
  AOI22_X1   g18588(.A1(new_n21628_), .A2(new_n21632_), .B1(new_n11870_), .B2(new_n21618_), .ZN(new_n21633_));
  NOR2_X1    g18589(.A1(new_n21633_), .A2(pi0781), .ZN(new_n21634_));
  NOR4_X1    g18590(.A1(new_n21620_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n21635_));
  NOR2_X1    g18591(.A1(new_n21625_), .A2(pi0785), .ZN(new_n21636_));
  NOR4_X1    g18592(.A1(new_n21626_), .A2(pi1155), .A3(new_n21595_), .A4(new_n21629_), .ZN(new_n21637_));
  NOR2_X1    g18593(.A1(new_n21637_), .A2(new_n11870_), .ZN(new_n21638_));
  XOR2_X1    g18594(.A1(new_n21638_), .A2(new_n21636_), .Z(new_n21639_));
  INV_X1     g18595(.I(new_n21639_), .ZN(new_n21640_));
  OAI21_X1   g18596(.A1(new_n21640_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n21641_));
  OAI21_X1   g18597(.A1(new_n21640_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n21642_));
  NOR2_X1    g18598(.A1(new_n21620_), .A2(new_n11939_), .ZN(new_n21643_));
  NOR4_X1    g18599(.A1(new_n21633_), .A2(new_n11934_), .A3(pi1154), .A4(new_n21643_), .ZN(new_n21644_));
  NOR2_X1    g18600(.A1(new_n21644_), .A2(new_n21642_), .ZN(new_n21645_));
  OAI22_X1   g18601(.A1(new_n21645_), .A2(pi0627), .B1(new_n21635_), .B2(new_n21641_), .ZN(new_n21646_));
  AOI21_X1   g18602(.A1(new_n21646_), .A2(pi0781), .B(new_n21634_), .ZN(new_n21647_));
  INV_X1     g18603(.I(new_n21643_), .ZN(new_n21648_));
  NOR2_X1    g18604(.A1(new_n21648_), .A2(new_n11962_), .ZN(new_n21649_));
  NOR4_X1    g18605(.A1(new_n21647_), .A2(new_n11967_), .A3(pi1159), .A4(new_n21649_), .ZN(new_n21650_));
  NOR2_X1    g18606(.A1(new_n21640_), .A2(pi0781), .ZN(new_n21651_));
  AOI21_X1   g18607(.A1(new_n11944_), .A2(new_n21639_), .B(new_n21642_), .ZN(new_n21652_));
  NOR2_X1    g18608(.A1(new_n21652_), .A2(new_n11969_), .ZN(new_n21653_));
  XOR2_X1    g18609(.A1(new_n21653_), .A2(new_n21651_), .Z(new_n21654_));
  AOI21_X1   g18610(.A1(new_n21654_), .A2(new_n16479_), .B(pi1159), .ZN(new_n21655_));
  INV_X1     g18611(.I(new_n21655_), .ZN(new_n21656_));
  NOR3_X1    g18612(.A1(new_n21650_), .A2(new_n11966_), .A3(new_n21656_), .ZN(new_n21657_));
  NOR4_X1    g18613(.A1(new_n21648_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n21658_));
  INV_X1     g18614(.I(new_n21654_), .ZN(new_n21659_));
  NOR2_X1    g18615(.A1(new_n21659_), .A2(new_n16482_), .ZN(new_n21660_));
  NOR3_X1    g18616(.A1(new_n21660_), .A2(pi0648), .A3(new_n21658_), .ZN(new_n21661_));
  AOI21_X1   g18617(.A1(new_n21647_), .A2(new_n11998_), .B(pi0789), .ZN(new_n21662_));
  OAI21_X1   g18618(.A1(new_n21657_), .A2(new_n21661_), .B(new_n21662_), .ZN(new_n21663_));
  NOR3_X1    g18619(.A1(new_n21648_), .A2(new_n11962_), .A3(new_n12015_), .ZN(new_n21664_));
  NAND2_X1   g18620(.A1(new_n21664_), .A2(new_n17154_), .ZN(new_n21665_));
  NOR2_X1    g18621(.A1(new_n14624_), .A2(new_n21595_), .ZN(new_n21666_));
  OAI21_X1   g18622(.A1(new_n16482_), .A2(new_n21659_), .B(new_n21655_), .ZN(new_n21667_));
  MUX2_X1    g18623(.I0(new_n21667_), .I1(new_n21654_), .S(new_n11985_), .Z(new_n21668_));
  AOI21_X1   g18624(.A1(new_n21668_), .A2(new_n14624_), .B(new_n21666_), .ZN(new_n21669_));
  INV_X1     g18625(.I(new_n21669_), .ZN(new_n21670_));
  OAI22_X1   g18626(.A1(new_n21670_), .A2(new_n17150_), .B1(new_n17151_), .B2(new_n21665_), .ZN(new_n21671_));
  NAND2_X1   g18627(.A1(new_n21671_), .A2(pi0629), .ZN(new_n21672_));
  OAI21_X1   g18628(.A1(new_n21665_), .A2(new_n17163_), .B(new_n15085_), .ZN(new_n21673_));
  AOI21_X1   g18629(.A1(new_n21669_), .A2(new_n12063_), .B(new_n21673_), .ZN(new_n21674_));
  NAND2_X1   g18630(.A1(new_n21672_), .A2(new_n21674_), .ZN(new_n21675_));
  INV_X1     g18631(.I(new_n21595_), .ZN(new_n21676_));
  MUX2_X1    g18632(.I0(new_n21668_), .I1(new_n21676_), .S(new_n11994_), .Z(new_n21677_));
  NOR2_X1    g18633(.A1(new_n21677_), .A2(new_n17167_), .ZN(new_n21678_));
  OAI21_X1   g18634(.A1(new_n21668_), .A2(new_n21595_), .B(pi0626), .ZN(new_n21679_));
  AOI21_X1   g18635(.A1(new_n21664_), .A2(new_n17173_), .B(pi0788), .ZN(new_n21680_));
  OAI21_X1   g18636(.A1(new_n21679_), .A2(new_n17171_), .B(new_n21680_), .ZN(new_n21681_));
  OAI21_X1   g18637(.A1(new_n21678_), .A2(new_n21681_), .B(new_n14732_), .ZN(new_n21682_));
  AOI21_X1   g18638(.A1(new_n21675_), .A2(new_n14726_), .B(new_n21682_), .ZN(new_n21683_));
  NAND3_X1   g18639(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n21595_), .ZN(new_n21684_));
  NOR2_X1    g18640(.A1(new_n21665_), .A2(new_n12068_), .ZN(new_n21685_));
  AOI21_X1   g18641(.A1(new_n21595_), .A2(pi0647), .B(pi1157), .ZN(new_n21686_));
  OAI21_X1   g18642(.A1(new_n21685_), .A2(new_n12061_), .B(new_n21686_), .ZN(new_n21687_));
  NOR2_X1    g18643(.A1(new_n21676_), .A2(pi0647), .ZN(new_n21688_));
  AOI21_X1   g18644(.A1(new_n21685_), .A2(pi0647), .B(new_n21688_), .ZN(new_n21689_));
  NAND2_X1   g18645(.A1(new_n21689_), .A2(new_n12088_), .ZN(new_n21690_));
  NAND2_X1   g18646(.A1(new_n21690_), .A2(pi0787), .ZN(new_n21691_));
  AOI21_X1   g18647(.A1(pi0630), .A2(new_n21687_), .B(new_n21691_), .ZN(new_n21692_));
  AOI22_X1   g18648(.A1(new_n21663_), .A2(new_n21683_), .B1(new_n21684_), .B2(new_n21692_), .ZN(new_n21693_));
  OR2_X2     g18649(.A1(new_n21693_), .A2(new_n12082_), .Z(new_n21694_));
  MUX2_X1    g18650(.I0(new_n21670_), .I1(new_n21676_), .S(new_n16841_), .Z(new_n21695_));
  MUX2_X1    g18651(.I0(new_n21695_), .I1(new_n21676_), .S(pi0644), .Z(new_n21696_));
  NAND2_X1   g18652(.A1(new_n21689_), .A2(pi1157), .ZN(new_n21697_));
  NOR2_X1    g18653(.A1(new_n21687_), .A2(new_n12048_), .ZN(new_n21698_));
  AOI22_X1   g18654(.A1(new_n21698_), .A2(new_n21697_), .B1(new_n12048_), .B2(new_n21685_), .ZN(new_n21699_));
  OAI21_X1   g18655(.A1(new_n21699_), .A2(new_n12082_), .B(new_n13168_), .ZN(new_n21700_));
  AOI21_X1   g18656(.A1(new_n21696_), .A2(pi0715), .B(new_n21700_), .ZN(new_n21701_));
  AOI21_X1   g18657(.A1(new_n21699_), .A2(new_n12082_), .B(pi0715), .ZN(new_n21702_));
  NAND2_X1   g18658(.A1(new_n21694_), .A2(new_n21702_), .ZN(new_n21703_));
  NAND3_X1   g18659(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n21704_));
  NOR2_X1    g18660(.A1(new_n21695_), .A2(new_n21704_), .ZN(new_n21705_));
  AOI22_X1   g18661(.A1(new_n21703_), .A2(new_n21705_), .B1(new_n21694_), .B2(new_n21701_), .ZN(new_n21706_));
  AOI21_X1   g18662(.A1(new_n21693_), .A2(new_n11867_), .B(new_n13184_), .ZN(new_n21707_));
  OAI21_X1   g18663(.A1(new_n21706_), .A2(new_n11867_), .B(new_n21707_), .ZN(new_n21708_));
  NOR2_X1    g18664(.A1(new_n12965_), .A2(pi0190), .ZN(new_n21709_));
  INV_X1     g18665(.I(new_n21709_), .ZN(new_n21710_));
  NAND2_X1   g18666(.A1(new_n21710_), .A2(new_n11997_), .ZN(new_n21711_));
  NOR2_X1    g18667(.A1(new_n16222_), .A2(pi0190), .ZN(new_n21712_));
  OAI21_X1   g18668(.A1(new_n14361_), .A2(new_n10096_), .B(pi0039), .ZN(new_n21713_));
  AOI21_X1   g18669(.A1(new_n13381_), .A2(new_n21712_), .B(new_n21713_), .ZN(new_n21714_));
  OAI21_X1   g18670(.A1(pi0763), .A2(new_n12793_), .B(new_n21714_), .ZN(new_n21715_));
  NOR2_X1    g18671(.A1(new_n12828_), .A2(pi0190), .ZN(new_n21716_));
  AOI21_X1   g18672(.A1(new_n12829_), .A2(pi0763), .B(pi0038), .ZN(new_n21717_));
  AOI21_X1   g18673(.A1(new_n21715_), .A2(new_n21717_), .B(new_n3232_), .ZN(new_n21718_));
  AOI21_X1   g18674(.A1(new_n10096_), .A2(new_n3232_), .B(new_n21718_), .ZN(new_n21719_));
  OAI21_X1   g18675(.A1(new_n21719_), .A2(new_n11914_), .B(new_n11870_), .ZN(new_n21720_));
  AOI21_X1   g18676(.A1(new_n11914_), .A2(new_n21709_), .B(new_n21720_), .ZN(new_n21721_));
  NAND2_X1   g18677(.A1(new_n21719_), .A2(new_n11924_), .ZN(new_n21722_));
  OAI22_X1   g18678(.A1(new_n21722_), .A2(pi0609), .B1(new_n12996_), .B2(new_n21709_), .ZN(new_n21723_));
  NAND2_X1   g18679(.A1(new_n21723_), .A2(new_n11912_), .ZN(new_n21724_));
  OAI22_X1   g18680(.A1(new_n21722_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n21709_), .ZN(new_n21725_));
  NAND2_X1   g18681(.A1(new_n21725_), .A2(pi1155), .ZN(new_n21726_));
  NAND2_X1   g18682(.A1(new_n21724_), .A2(new_n21726_), .ZN(new_n21727_));
  NAND2_X1   g18683(.A1(new_n21727_), .A2(pi0785), .ZN(new_n21728_));
  XNOR2_X1   g18684(.A1(new_n21728_), .A2(new_n21721_), .ZN(new_n21729_));
  OAI21_X1   g18685(.A1(new_n21710_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n21730_));
  AOI21_X1   g18686(.A1(new_n21729_), .A2(pi0618), .B(new_n21730_), .ZN(new_n21731_));
  INV_X1     g18687(.I(new_n21729_), .ZN(new_n21732_));
  AOI21_X1   g18688(.A1(new_n21710_), .A2(new_n11934_), .B(pi1154), .ZN(new_n21733_));
  OAI21_X1   g18689(.A1(new_n21732_), .A2(new_n11934_), .B(new_n21733_), .ZN(new_n21734_));
  NAND2_X1   g18690(.A1(new_n21734_), .A2(new_n21731_), .ZN(new_n21735_));
  MUX2_X1    g18691(.I0(new_n21735_), .I1(new_n21729_), .S(new_n11969_), .Z(new_n21736_));
  NAND2_X1   g18692(.A1(new_n21736_), .A2(new_n11985_), .ZN(new_n21737_));
  NOR3_X1    g18693(.A1(new_n21709_), .A2(pi0619), .A3(pi1159), .ZN(new_n21738_));
  NOR2_X1    g18694(.A1(new_n21738_), .A2(new_n11985_), .ZN(new_n21739_));
  XOR2_X1    g18695(.A1(new_n21737_), .A2(new_n21739_), .Z(new_n21740_));
  OAI21_X1   g18696(.A1(new_n21740_), .A2(new_n11997_), .B(new_n21711_), .ZN(new_n21741_));
  NOR2_X1    g18697(.A1(new_n21709_), .A2(new_n12054_), .ZN(new_n21742_));
  AOI21_X1   g18698(.A1(new_n21741_), .A2(new_n12054_), .B(new_n21742_), .ZN(new_n21743_));
  INV_X1     g18699(.I(new_n21743_), .ZN(new_n21744_));
  NOR2_X1    g18700(.A1(new_n21709_), .A2(new_n12092_), .ZN(new_n21745_));
  AOI21_X1   g18701(.A1(new_n21744_), .A2(new_n12092_), .B(new_n21745_), .ZN(new_n21746_));
  NAND2_X1   g18702(.A1(new_n21746_), .A2(new_n12082_), .ZN(new_n21747_));
  AOI21_X1   g18703(.A1(new_n21709_), .A2(pi0644), .B(new_n12099_), .ZN(new_n21748_));
  AOI21_X1   g18704(.A1(new_n21747_), .A2(new_n21748_), .B(pi1160), .ZN(new_n21749_));
  NOR2_X1    g18705(.A1(new_n21709_), .A2(new_n13114_), .ZN(new_n21750_));
  NOR2_X1    g18706(.A1(new_n21710_), .A2(new_n12014_), .ZN(new_n21751_));
  NOR2_X1    g18707(.A1(new_n21709_), .A2(new_n11961_), .ZN(new_n21752_));
  NAND2_X1   g18708(.A1(new_n10096_), .A2(new_n16255_), .ZN(new_n21753_));
  OAI21_X1   g18709(.A1(new_n12902_), .A2(new_n21753_), .B(new_n3231_), .ZN(new_n21754_));
  NOR3_X1    g18710(.A1(new_n13399_), .A2(pi0190), .A3(new_n13396_), .ZN(new_n21755_));
  AOI21_X1   g18711(.A1(new_n13399_), .A2(new_n10096_), .B(new_n13395_), .ZN(new_n21756_));
  NAND3_X1   g18712(.A1(new_n13403_), .A2(new_n3172_), .A3(new_n16255_), .ZN(new_n21757_));
  NOR4_X1    g18713(.A1(new_n21755_), .A2(new_n21756_), .A3(new_n21716_), .A4(new_n21757_), .ZN(new_n21758_));
  AOI22_X1   g18714(.A1(new_n21758_), .A2(new_n21754_), .B1(pi0190), .B2(new_n3232_), .ZN(new_n21759_));
  NAND2_X1   g18715(.A1(new_n21759_), .A2(new_n11891_), .ZN(new_n21760_));
  AOI21_X1   g18716(.A1(new_n21759_), .A2(new_n12970_), .B(new_n21710_), .ZN(new_n21761_));
  NOR3_X1    g18717(.A1(new_n21759_), .A2(pi0625), .A3(new_n21709_), .ZN(new_n21762_));
  NOR3_X1    g18718(.A1(new_n21762_), .A2(new_n21761_), .A3(pi1153), .ZN(new_n21763_));
  NAND4_X1   g18719(.A1(new_n21759_), .A2(pi0625), .A3(new_n11893_), .A4(new_n21710_), .ZN(new_n21764_));
  NAND2_X1   g18720(.A1(new_n21763_), .A2(new_n21764_), .ZN(new_n21765_));
  NAND2_X1   g18721(.A1(new_n21765_), .A2(pi0778), .ZN(new_n21766_));
  XOR2_X1    g18722(.A1(new_n21766_), .A2(new_n21760_), .Z(new_n21767_));
  NOR2_X1    g18723(.A1(new_n21767_), .A2(new_n13024_), .ZN(new_n21768_));
  AOI21_X1   g18724(.A1(new_n13024_), .A2(new_n21709_), .B(new_n21768_), .ZN(new_n21769_));
  AOI21_X1   g18725(.A1(new_n21769_), .A2(new_n11961_), .B(new_n21752_), .ZN(new_n21770_));
  AOI21_X1   g18726(.A1(new_n21770_), .A2(new_n12014_), .B(new_n21751_), .ZN(new_n21771_));
  AOI21_X1   g18727(.A1(new_n21771_), .A2(new_n13114_), .B(new_n21750_), .ZN(new_n21772_));
  NOR2_X1    g18728(.A1(new_n21772_), .A2(pi0628), .ZN(new_n21773_));
  AOI21_X1   g18729(.A1(pi0628), .A2(new_n21710_), .B(new_n21773_), .ZN(new_n21774_));
  NOR2_X1    g18730(.A1(new_n21774_), .A2(pi1156), .ZN(new_n21775_));
  NOR2_X1    g18731(.A1(new_n21772_), .A2(new_n12031_), .ZN(new_n21776_));
  AOI21_X1   g18732(.A1(new_n12031_), .A2(new_n21710_), .B(new_n21776_), .ZN(new_n21777_));
  NOR2_X1    g18733(.A1(new_n21777_), .A2(new_n12026_), .ZN(new_n21778_));
  OAI21_X1   g18734(.A1(new_n21775_), .A2(new_n21778_), .B(pi0792), .ZN(new_n21779_));
  OAI21_X1   g18735(.A1(pi0792), .A2(new_n21772_), .B(new_n21779_), .ZN(new_n21780_));
  NOR2_X1    g18736(.A1(new_n21709_), .A2(new_n12061_), .ZN(new_n21781_));
  AOI21_X1   g18737(.A1(new_n21780_), .A2(new_n12061_), .B(new_n21781_), .ZN(new_n21782_));
  NOR2_X1    g18738(.A1(new_n21782_), .A2(pi1157), .ZN(new_n21783_));
  NOR2_X1    g18739(.A1(new_n21709_), .A2(pi0647), .ZN(new_n21784_));
  AOI21_X1   g18740(.A1(new_n21780_), .A2(pi0647), .B(new_n21784_), .ZN(new_n21785_));
  NOR2_X1    g18741(.A1(new_n21785_), .A2(new_n12049_), .ZN(new_n21786_));
  NOR2_X1    g18742(.A1(new_n21783_), .A2(new_n21786_), .ZN(new_n21787_));
  NOR2_X1    g18743(.A1(new_n21787_), .A2(new_n12048_), .ZN(new_n21788_));
  AOI21_X1   g18744(.A1(new_n12048_), .A2(new_n21780_), .B(new_n21788_), .ZN(new_n21789_));
  NAND2_X1   g18745(.A1(new_n21789_), .A2(pi0644), .ZN(new_n21790_));
  AOI21_X1   g18746(.A1(new_n21790_), .A2(new_n12099_), .B(new_n21749_), .ZN(new_n21791_));
  NOR3_X1    g18747(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n21792_));
  NAND2_X1   g18748(.A1(new_n21746_), .A2(new_n21792_), .ZN(new_n21793_));
  NAND2_X1   g18749(.A1(new_n21793_), .A2(pi0715), .ZN(new_n21794_));
  AOI21_X1   g18750(.A1(new_n21789_), .A2(new_n12082_), .B(new_n21794_), .ZN(new_n21795_));
  OAI21_X1   g18751(.A1(new_n21791_), .A2(new_n21795_), .B(pi0790), .ZN(new_n21796_));
  NAND2_X1   g18752(.A1(new_n21749_), .A2(new_n12082_), .ZN(new_n21797_));
  AOI21_X1   g18753(.A1(new_n21793_), .A2(pi0644), .B(pi0790), .ZN(new_n21798_));
  NAND2_X1   g18754(.A1(new_n21797_), .A2(new_n21798_), .ZN(new_n21799_));
  NAND2_X1   g18755(.A1(new_n21785_), .A2(new_n12060_), .ZN(new_n21800_));
  AOI21_X1   g18756(.A1(new_n21782_), .A2(pi0630), .B(new_n12090_), .ZN(new_n21801_));
  NAND2_X1   g18757(.A1(new_n21744_), .A2(new_n15078_), .ZN(new_n21802_));
  AOI21_X1   g18758(.A1(new_n21801_), .A2(new_n21800_), .B(new_n21802_), .ZN(new_n21803_));
  AND2_X2    g18759(.A1(new_n21777_), .A2(new_n12030_), .Z(new_n21804_));
  NAND2_X1   g18760(.A1(new_n21774_), .A2(pi0629), .ZN(new_n21805_));
  NAND2_X1   g18761(.A1(new_n21805_), .A2(new_n17299_), .ZN(new_n21806_));
  OR2_X2     g18762(.A1(new_n21806_), .A2(new_n21804_), .Z(new_n21807_));
  NAND3_X1   g18763(.A1(new_n21807_), .A2(new_n17304_), .A3(new_n21741_), .ZN(new_n21808_));
  NAND2_X1   g18764(.A1(new_n21736_), .A2(pi0619), .ZN(new_n21809_));
  NAND2_X1   g18765(.A1(new_n21709_), .A2(pi0619), .ZN(new_n21810_));
  INV_X1     g18766(.I(new_n21719_), .ZN(new_n21811_));
  NAND2_X1   g18767(.A1(new_n17309_), .A2(new_n16222_), .ZN(new_n21812_));
  AOI21_X1   g18768(.A1(new_n12122_), .A2(new_n21812_), .B(pi0039), .ZN(new_n21813_));
  AOI21_X1   g18769(.A1(new_n13644_), .A2(new_n21624_), .B(new_n10096_), .ZN(new_n21814_));
  AOI21_X1   g18770(.A1(new_n21814_), .A2(new_n5156_), .B(new_n3172_), .ZN(new_n21815_));
  OAI21_X1   g18771(.A1(new_n21813_), .A2(pi0190), .B(new_n21815_), .ZN(new_n21816_));
  NOR2_X1    g18772(.A1(new_n13333_), .A2(new_n10096_), .ZN(new_n21817_));
  OAI21_X1   g18773(.A1(new_n12515_), .A2(new_n10096_), .B(new_n16222_), .ZN(new_n21818_));
  NOR3_X1    g18774(.A1(new_n12645_), .A2(new_n10096_), .A3(new_n13347_), .ZN(new_n21819_));
  AOI21_X1   g18775(.A1(new_n12645_), .A2(pi0190), .B(new_n12665_), .ZN(new_n21820_));
  OAI21_X1   g18776(.A1(new_n21819_), .A2(new_n21820_), .B(pi0763), .ZN(new_n21821_));
  NAND2_X1   g18777(.A1(new_n13360_), .A2(pi0190), .ZN(new_n21822_));
  NAND2_X1   g18778(.A1(new_n13362_), .A2(pi0190), .ZN(new_n21823_));
  NAND4_X1   g18779(.A1(new_n21821_), .A2(new_n16242_), .A3(new_n21822_), .A4(new_n21823_), .ZN(new_n21824_));
  AOI21_X1   g18780(.A1(new_n21824_), .A2(new_n3172_), .B(pi0039), .ZN(new_n21825_));
  OAI21_X1   g18781(.A1(new_n21817_), .A2(new_n21818_), .B(new_n21825_), .ZN(new_n21826_));
  NAND2_X1   g18782(.A1(new_n3232_), .A2(new_n16255_), .ZN(new_n21827_));
  AOI21_X1   g18783(.A1(new_n21826_), .A2(new_n21816_), .B(new_n21827_), .ZN(new_n21828_));
  NAND2_X1   g18784(.A1(new_n21715_), .A2(new_n21717_), .ZN(new_n21829_));
  NAND2_X1   g18785(.A1(new_n21829_), .A2(new_n16255_), .ZN(new_n21830_));
  OAI22_X1   g18786(.A1(new_n21828_), .A2(new_n21830_), .B1(new_n10096_), .B2(new_n3231_), .ZN(new_n21831_));
  OAI21_X1   g18787(.A1(new_n21831_), .A2(pi0625), .B(new_n21811_), .ZN(new_n21832_));
  NAND3_X1   g18788(.A1(new_n21831_), .A2(new_n12970_), .A3(new_n21719_), .ZN(new_n21833_));
  NAND4_X1   g18789(.A1(new_n21832_), .A2(new_n21833_), .A3(new_n12977_), .A4(new_n21764_), .ZN(new_n21834_));
  INV_X1     g18790(.I(new_n21763_), .ZN(new_n21835_));
  NOR4_X1    g18791(.A1(new_n21831_), .A2(new_n12970_), .A3(pi1153), .A4(new_n21811_), .ZN(new_n21836_));
  OAI21_X1   g18792(.A1(new_n21836_), .A2(new_n21835_), .B(new_n13657_), .ZN(new_n21837_));
  NAND2_X1   g18793(.A1(new_n21834_), .A2(new_n21837_), .ZN(new_n21838_));
  NOR2_X1    g18794(.A1(new_n21831_), .A2(pi0778), .ZN(new_n21839_));
  AOI21_X1   g18795(.A1(new_n21838_), .A2(pi0778), .B(new_n21839_), .ZN(new_n21840_));
  NOR2_X1    g18796(.A1(new_n21840_), .A2(pi0785), .ZN(new_n21841_));
  INV_X1     g18797(.I(new_n21767_), .ZN(new_n21842_));
  NAND3_X1   g18798(.A1(new_n21842_), .A2(pi0609), .A3(pi1155), .ZN(new_n21843_));
  NAND3_X1   g18799(.A1(new_n21843_), .A2(new_n11923_), .A3(new_n21726_), .ZN(new_n21844_));
  NOR4_X1    g18800(.A1(new_n21840_), .A2(new_n11903_), .A3(new_n21842_), .A4(pi1155), .ZN(new_n21845_));
  NAND2_X1   g18801(.A1(new_n21724_), .A2(pi0660), .ZN(new_n21846_));
  NOR2_X1    g18802(.A1(new_n21845_), .A2(new_n21846_), .ZN(new_n21847_));
  NOR2_X1    g18803(.A1(new_n21847_), .A2(new_n11870_), .ZN(new_n21848_));
  AOI21_X1   g18804(.A1(new_n21848_), .A2(new_n21844_), .B(new_n21841_), .ZN(new_n21849_));
  INV_X1     g18805(.I(new_n21769_), .ZN(new_n21850_));
  NOR4_X1    g18806(.A1(new_n21849_), .A2(new_n11934_), .A3(pi1154), .A4(new_n21850_), .ZN(new_n21851_));
  NAND2_X1   g18807(.A1(new_n21731_), .A2(pi0627), .ZN(new_n21852_));
  NOR3_X1    g18808(.A1(new_n21769_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n21853_));
  NAND2_X1   g18809(.A1(new_n21734_), .A2(new_n11949_), .ZN(new_n21854_));
  OAI22_X1   g18810(.A1(new_n21851_), .A2(new_n21852_), .B1(new_n21853_), .B2(new_n21854_), .ZN(new_n21855_));
  MUX2_X1    g18811(.I0(new_n21855_), .I1(new_n21849_), .S(new_n11969_), .Z(new_n21856_));
  XNOR2_X1   g18812(.A1(new_n21856_), .A2(new_n21770_), .ZN(new_n21857_));
  NOR2_X1    g18813(.A1(new_n21857_), .A2(new_n11967_), .ZN(new_n21858_));
  NAND3_X1   g18814(.A1(new_n21809_), .A2(new_n11869_), .A3(new_n21810_), .ZN(new_n21859_));
  XOR2_X1    g18815(.A1(new_n21858_), .A2(new_n21856_), .Z(new_n21860_));
  AOI21_X1   g18816(.A1(new_n21710_), .A2(new_n11967_), .B(pi1159), .ZN(new_n21861_));
  AOI21_X1   g18817(.A1(new_n21809_), .A2(new_n21861_), .B(pi0648), .ZN(new_n21862_));
  OAI21_X1   g18818(.A1(new_n21860_), .A2(pi1159), .B(new_n21862_), .ZN(new_n21863_));
  OR2_X2     g18819(.A1(new_n21856_), .A2(pi0789), .Z(new_n21864_));
  NAND3_X1   g18820(.A1(new_n21740_), .A2(pi0626), .A3(new_n21710_), .ZN(new_n21865_));
  OAI21_X1   g18821(.A1(new_n21740_), .A2(new_n11994_), .B(new_n21709_), .ZN(new_n21866_));
  AOI21_X1   g18822(.A1(new_n21866_), .A2(new_n21865_), .B(new_n17167_), .ZN(new_n21867_));
  AOI21_X1   g18823(.A1(new_n21740_), .A2(new_n21710_), .B(new_n11994_), .ZN(new_n21868_));
  NAND2_X1   g18824(.A1(new_n21868_), .A2(new_n11990_), .ZN(new_n21869_));
  NOR2_X1    g18825(.A1(new_n21771_), .A2(new_n12020_), .ZN(new_n21870_));
  NOR2_X1    g18826(.A1(new_n21870_), .A2(pi0788), .ZN(new_n21871_));
  NAND2_X1   g18827(.A1(new_n21869_), .A2(new_n21871_), .ZN(new_n21872_));
  OAI21_X1   g18828(.A1(new_n21872_), .A2(new_n21867_), .B(new_n17372_), .ZN(new_n21873_));
  AOI21_X1   g18829(.A1(new_n11998_), .A2(new_n21864_), .B(new_n21873_), .ZN(new_n21874_));
  NAND3_X1   g18830(.A1(new_n21863_), .A2(new_n21859_), .A3(new_n21874_), .ZN(new_n21875_));
  AOI21_X1   g18831(.A1(new_n21875_), .A2(new_n21808_), .B(new_n14725_), .ZN(new_n21876_));
  OAI21_X1   g18832(.A1(new_n21876_), .A2(new_n21803_), .B(new_n21799_), .ZN(new_n21877_));
  AOI21_X1   g18833(.A1(new_n21796_), .A2(new_n21877_), .B(po1038), .ZN(new_n21878_));
  OAI21_X1   g18834(.A1(new_n6845_), .A2(pi0190), .B(new_n13184_), .ZN(new_n21879_));
  OAI21_X1   g18835(.A1(new_n21878_), .A2(new_n21879_), .B(new_n21708_), .ZN(po0347));
  NOR2_X1    g18836(.A1(new_n2925_), .A2(pi0191), .ZN(new_n21881_));
  NOR2_X1    g18837(.A1(new_n11877_), .A2(new_n16270_), .ZN(new_n21882_));
  NOR2_X1    g18838(.A1(new_n21882_), .A2(new_n21881_), .ZN(new_n21883_));
  AOI21_X1   g18839(.A1(new_n11886_), .A2(pi0729), .B(new_n21881_), .ZN(new_n21884_));
  NOR2_X1    g18840(.A1(new_n21884_), .A2(new_n11874_), .ZN(new_n21885_));
  INV_X1     g18841(.I(new_n21885_), .ZN(new_n21886_));
  NAND2_X1   g18842(.A1(new_n21886_), .A2(new_n21883_), .ZN(new_n21887_));
  NAND2_X1   g18843(.A1(new_n21887_), .A2(new_n11891_), .ZN(new_n21888_));
  NOR2_X1    g18844(.A1(new_n21886_), .A2(new_n12970_), .ZN(new_n21889_));
  NOR4_X1    g18845(.A1(new_n21889_), .A2(new_n11893_), .A3(new_n21881_), .A4(new_n21882_), .ZN(new_n21890_));
  NOR2_X1    g18846(.A1(new_n13201_), .A2(new_n16303_), .ZN(new_n21891_));
  NOR2_X1    g18847(.A1(new_n21881_), .A2(pi1153), .ZN(new_n21892_));
  INV_X1     g18848(.I(new_n21892_), .ZN(new_n21893_));
  NOR2_X1    g18849(.A1(new_n21891_), .A2(new_n21893_), .ZN(new_n21894_));
  INV_X1     g18850(.I(new_n21894_), .ZN(new_n21895_));
  NAND2_X1   g18851(.A1(new_n21895_), .A2(pi0608), .ZN(new_n21896_));
  INV_X1     g18852(.I(new_n21889_), .ZN(new_n21897_));
  AOI21_X1   g18853(.A1(new_n21897_), .A2(new_n21887_), .B(new_n21893_), .ZN(new_n21898_));
  OAI21_X1   g18854(.A1(new_n21891_), .A2(new_n21884_), .B(pi1153), .ZN(new_n21899_));
  NAND2_X1   g18855(.A1(new_n21899_), .A2(new_n13657_), .ZN(new_n21900_));
  OAI22_X1   g18856(.A1(new_n21896_), .A2(new_n21890_), .B1(new_n21898_), .B2(new_n21900_), .ZN(new_n21901_));
  NAND2_X1   g18857(.A1(new_n21901_), .A2(pi0778), .ZN(new_n21902_));
  XOR2_X1    g18858(.A1(new_n21902_), .A2(new_n21888_), .Z(new_n21903_));
  INV_X1     g18859(.I(new_n21903_), .ZN(new_n21904_));
  NAND2_X1   g18860(.A1(new_n21895_), .A2(new_n21899_), .ZN(new_n21905_));
  MUX2_X1    g18861(.I0(new_n21905_), .I1(new_n21884_), .S(new_n11891_), .Z(new_n21906_));
  XNOR2_X1   g18862(.A1(new_n21903_), .A2(new_n21906_), .ZN(new_n21907_));
  NAND2_X1   g18863(.A1(new_n21907_), .A2(pi0609), .ZN(new_n21908_));
  XOR2_X1    g18864(.A1(new_n21908_), .A2(new_n21904_), .Z(new_n21909_));
  INV_X1     g18865(.I(new_n21882_), .ZN(new_n21910_));
  NOR2_X1    g18866(.A1(new_n21883_), .A2(new_n11925_), .ZN(new_n21911_));
  NOR4_X1    g18867(.A1(new_n21911_), .A2(pi1155), .A3(new_n12997_), .A4(new_n21910_), .ZN(new_n21912_));
  NOR2_X1    g18868(.A1(new_n21912_), .A2(pi0660), .ZN(new_n21913_));
  OAI21_X1   g18869(.A1(new_n21909_), .A2(pi1155), .B(new_n21913_), .ZN(new_n21914_));
  NOR2_X1    g18870(.A1(new_n21910_), .A2(new_n12997_), .ZN(new_n21915_));
  NOR4_X1    g18871(.A1(new_n21915_), .A2(new_n11923_), .A3(pi1155), .A4(new_n21881_), .ZN(new_n21917_));
  NOR2_X1    g18872(.A1(new_n21917_), .A2(new_n11870_), .ZN(new_n21918_));
  AOI22_X1   g18873(.A1(new_n21914_), .A2(new_n21918_), .B1(new_n11870_), .B2(new_n21904_), .ZN(new_n21919_));
  NOR2_X1    g18874(.A1(new_n21919_), .A2(pi0781), .ZN(new_n21920_));
  NOR4_X1    g18875(.A1(new_n21906_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n21921_));
  NOR2_X1    g18876(.A1(new_n21911_), .A2(pi0785), .ZN(new_n21922_));
  NOR4_X1    g18877(.A1(new_n21912_), .A2(pi1155), .A3(new_n21881_), .A4(new_n21915_), .ZN(new_n21923_));
  NOR2_X1    g18878(.A1(new_n21923_), .A2(new_n11870_), .ZN(new_n21924_));
  XOR2_X1    g18879(.A1(new_n21924_), .A2(new_n21922_), .Z(new_n21925_));
  INV_X1     g18880(.I(new_n21925_), .ZN(new_n21926_));
  OAI21_X1   g18881(.A1(new_n21926_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n21927_));
  OAI21_X1   g18882(.A1(new_n21926_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n21928_));
  NOR2_X1    g18883(.A1(new_n21906_), .A2(new_n11939_), .ZN(new_n21929_));
  NOR4_X1    g18884(.A1(new_n21919_), .A2(new_n11934_), .A3(pi1154), .A4(new_n21929_), .ZN(new_n21930_));
  NOR2_X1    g18885(.A1(new_n21930_), .A2(new_n21928_), .ZN(new_n21931_));
  OAI22_X1   g18886(.A1(new_n21931_), .A2(pi0627), .B1(new_n21921_), .B2(new_n21927_), .ZN(new_n21932_));
  AOI21_X1   g18887(.A1(new_n21932_), .A2(pi0781), .B(new_n21920_), .ZN(new_n21933_));
  INV_X1     g18888(.I(new_n21929_), .ZN(new_n21934_));
  NOR2_X1    g18889(.A1(new_n21934_), .A2(new_n11962_), .ZN(new_n21935_));
  NOR4_X1    g18890(.A1(new_n21933_), .A2(new_n11967_), .A3(pi1159), .A4(new_n21935_), .ZN(new_n21936_));
  NOR2_X1    g18891(.A1(new_n21926_), .A2(pi0781), .ZN(new_n21937_));
  AOI21_X1   g18892(.A1(new_n11944_), .A2(new_n21925_), .B(new_n21928_), .ZN(new_n21938_));
  NOR2_X1    g18893(.A1(new_n21938_), .A2(new_n11969_), .ZN(new_n21939_));
  XOR2_X1    g18894(.A1(new_n21939_), .A2(new_n21937_), .Z(new_n21940_));
  AOI21_X1   g18895(.A1(new_n21940_), .A2(new_n16479_), .B(pi1159), .ZN(new_n21941_));
  INV_X1     g18896(.I(new_n21941_), .ZN(new_n21942_));
  NOR3_X1    g18897(.A1(new_n21936_), .A2(new_n11966_), .A3(new_n21942_), .ZN(new_n21943_));
  NOR4_X1    g18898(.A1(new_n21934_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n21944_));
  INV_X1     g18899(.I(new_n21940_), .ZN(new_n21945_));
  NOR2_X1    g18900(.A1(new_n21945_), .A2(new_n16482_), .ZN(new_n21946_));
  NOR3_X1    g18901(.A1(new_n21946_), .A2(pi0648), .A3(new_n21944_), .ZN(new_n21947_));
  AOI21_X1   g18902(.A1(new_n21933_), .A2(new_n11998_), .B(pi0789), .ZN(new_n21948_));
  OAI21_X1   g18903(.A1(new_n21943_), .A2(new_n21947_), .B(new_n21948_), .ZN(new_n21949_));
  NOR3_X1    g18904(.A1(new_n21934_), .A2(new_n11962_), .A3(new_n12015_), .ZN(new_n21950_));
  NAND2_X1   g18905(.A1(new_n21950_), .A2(new_n17154_), .ZN(new_n21951_));
  NOR2_X1    g18906(.A1(new_n14624_), .A2(new_n21881_), .ZN(new_n21952_));
  OAI21_X1   g18907(.A1(new_n16482_), .A2(new_n21945_), .B(new_n21941_), .ZN(new_n21953_));
  MUX2_X1    g18908(.I0(new_n21953_), .I1(new_n21940_), .S(new_n11985_), .Z(new_n21954_));
  AOI21_X1   g18909(.A1(new_n21954_), .A2(new_n14624_), .B(new_n21952_), .ZN(new_n21955_));
  INV_X1     g18910(.I(new_n21955_), .ZN(new_n21956_));
  OAI22_X1   g18911(.A1(new_n21956_), .A2(new_n17150_), .B1(new_n17151_), .B2(new_n21951_), .ZN(new_n21957_));
  NAND2_X1   g18912(.A1(new_n21957_), .A2(pi0629), .ZN(new_n21958_));
  OAI21_X1   g18913(.A1(new_n21951_), .A2(new_n17163_), .B(new_n15085_), .ZN(new_n21959_));
  AOI21_X1   g18914(.A1(new_n21955_), .A2(new_n12063_), .B(new_n21959_), .ZN(new_n21960_));
  NAND2_X1   g18915(.A1(new_n21958_), .A2(new_n21960_), .ZN(new_n21961_));
  INV_X1     g18916(.I(new_n21881_), .ZN(new_n21962_));
  MUX2_X1    g18917(.I0(new_n21954_), .I1(new_n21962_), .S(new_n11994_), .Z(new_n21963_));
  NOR2_X1    g18918(.A1(new_n21963_), .A2(new_n17167_), .ZN(new_n21964_));
  OAI21_X1   g18919(.A1(new_n21954_), .A2(new_n21881_), .B(pi0626), .ZN(new_n21965_));
  AOI21_X1   g18920(.A1(new_n21950_), .A2(new_n17173_), .B(pi0788), .ZN(new_n21966_));
  OAI21_X1   g18921(.A1(new_n21965_), .A2(new_n17171_), .B(new_n21966_), .ZN(new_n21967_));
  OAI21_X1   g18922(.A1(new_n21964_), .A2(new_n21967_), .B(new_n14732_), .ZN(new_n21968_));
  AOI21_X1   g18923(.A1(new_n21961_), .A2(new_n14726_), .B(new_n21968_), .ZN(new_n21969_));
  NAND3_X1   g18924(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n21881_), .ZN(new_n21970_));
  NOR2_X1    g18925(.A1(new_n21951_), .A2(new_n12068_), .ZN(new_n21971_));
  AOI21_X1   g18926(.A1(new_n21881_), .A2(pi0647), .B(pi1157), .ZN(new_n21972_));
  OAI21_X1   g18927(.A1(new_n21971_), .A2(new_n12061_), .B(new_n21972_), .ZN(new_n21973_));
  NOR2_X1    g18928(.A1(new_n21962_), .A2(pi0647), .ZN(new_n21974_));
  AOI21_X1   g18929(.A1(new_n21971_), .A2(pi0647), .B(new_n21974_), .ZN(new_n21975_));
  NAND2_X1   g18930(.A1(new_n21975_), .A2(new_n12088_), .ZN(new_n21976_));
  NAND2_X1   g18931(.A1(new_n21976_), .A2(pi0787), .ZN(new_n21977_));
  AOI21_X1   g18932(.A1(pi0630), .A2(new_n21973_), .B(new_n21977_), .ZN(new_n21978_));
  AOI22_X1   g18933(.A1(new_n21949_), .A2(new_n21969_), .B1(new_n21970_), .B2(new_n21978_), .ZN(new_n21979_));
  OR2_X2     g18934(.A1(new_n21979_), .A2(new_n12082_), .Z(new_n21980_));
  MUX2_X1    g18935(.I0(new_n21956_), .I1(new_n21962_), .S(new_n16841_), .Z(new_n21981_));
  MUX2_X1    g18936(.I0(new_n21981_), .I1(new_n21962_), .S(pi0644), .Z(new_n21982_));
  NAND2_X1   g18937(.A1(new_n21975_), .A2(pi1157), .ZN(new_n21983_));
  NOR2_X1    g18938(.A1(new_n21973_), .A2(new_n12048_), .ZN(new_n21984_));
  AOI22_X1   g18939(.A1(new_n21984_), .A2(new_n21983_), .B1(new_n12048_), .B2(new_n21971_), .ZN(new_n21985_));
  OAI21_X1   g18940(.A1(new_n21985_), .A2(new_n12082_), .B(new_n13168_), .ZN(new_n21986_));
  AOI21_X1   g18941(.A1(new_n21982_), .A2(pi0715), .B(new_n21986_), .ZN(new_n21987_));
  AOI21_X1   g18942(.A1(new_n21985_), .A2(new_n12082_), .B(pi0715), .ZN(new_n21988_));
  NAND2_X1   g18943(.A1(new_n21980_), .A2(new_n21988_), .ZN(new_n21989_));
  NAND3_X1   g18944(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n21990_));
  NOR2_X1    g18945(.A1(new_n21981_), .A2(new_n21990_), .ZN(new_n21991_));
  AOI22_X1   g18946(.A1(new_n21989_), .A2(new_n21991_), .B1(new_n21980_), .B2(new_n21987_), .ZN(new_n21992_));
  AOI21_X1   g18947(.A1(new_n21979_), .A2(new_n11867_), .B(new_n13184_), .ZN(new_n21993_));
  OAI21_X1   g18948(.A1(new_n21992_), .A2(new_n11867_), .B(new_n21993_), .ZN(new_n21994_));
  NOR2_X1    g18949(.A1(new_n12965_), .A2(pi0191), .ZN(new_n21995_));
  INV_X1     g18950(.I(new_n21995_), .ZN(new_n21996_));
  NAND2_X1   g18951(.A1(new_n21996_), .A2(new_n11997_), .ZN(new_n21997_));
  NOR2_X1    g18952(.A1(new_n16270_), .A2(pi0191), .ZN(new_n21998_));
  OAI21_X1   g18953(.A1(new_n14361_), .A2(new_n11361_), .B(pi0039), .ZN(new_n21999_));
  AOI21_X1   g18954(.A1(new_n13381_), .A2(new_n21998_), .B(new_n21999_), .ZN(new_n22000_));
  OAI21_X1   g18955(.A1(pi0746), .A2(new_n12793_), .B(new_n22000_), .ZN(new_n22001_));
  NOR2_X1    g18956(.A1(new_n12828_), .A2(pi0191), .ZN(new_n22002_));
  AOI21_X1   g18957(.A1(new_n12829_), .A2(pi0746), .B(pi0038), .ZN(new_n22003_));
  AOI21_X1   g18958(.A1(new_n22001_), .A2(new_n22003_), .B(new_n3232_), .ZN(new_n22004_));
  AOI21_X1   g18959(.A1(new_n11361_), .A2(new_n3232_), .B(new_n22004_), .ZN(new_n22005_));
  OAI21_X1   g18960(.A1(new_n22005_), .A2(new_n11914_), .B(new_n11870_), .ZN(new_n22006_));
  AOI21_X1   g18961(.A1(new_n11914_), .A2(new_n21995_), .B(new_n22006_), .ZN(new_n22007_));
  NAND2_X1   g18962(.A1(new_n22005_), .A2(new_n11924_), .ZN(new_n22008_));
  OAI22_X1   g18963(.A1(new_n22008_), .A2(pi0609), .B1(new_n12996_), .B2(new_n21995_), .ZN(new_n22009_));
  NAND2_X1   g18964(.A1(new_n22009_), .A2(new_n11912_), .ZN(new_n22010_));
  OAI22_X1   g18965(.A1(new_n22008_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n21995_), .ZN(new_n22011_));
  NAND2_X1   g18966(.A1(new_n22011_), .A2(pi1155), .ZN(new_n22012_));
  NAND2_X1   g18967(.A1(new_n22010_), .A2(new_n22012_), .ZN(new_n22013_));
  NAND2_X1   g18968(.A1(new_n22013_), .A2(pi0785), .ZN(new_n22014_));
  XNOR2_X1   g18969(.A1(new_n22014_), .A2(new_n22007_), .ZN(new_n22015_));
  OAI21_X1   g18970(.A1(new_n21996_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n22016_));
  AOI21_X1   g18971(.A1(new_n22015_), .A2(pi0618), .B(new_n22016_), .ZN(new_n22017_));
  INV_X1     g18972(.I(new_n22015_), .ZN(new_n22018_));
  AOI21_X1   g18973(.A1(new_n21996_), .A2(new_n11934_), .B(pi1154), .ZN(new_n22019_));
  OAI21_X1   g18974(.A1(new_n22018_), .A2(new_n11934_), .B(new_n22019_), .ZN(new_n22020_));
  NAND2_X1   g18975(.A1(new_n22020_), .A2(new_n22017_), .ZN(new_n22021_));
  MUX2_X1    g18976(.I0(new_n22021_), .I1(new_n22015_), .S(new_n11969_), .Z(new_n22022_));
  NAND2_X1   g18977(.A1(new_n22022_), .A2(new_n11985_), .ZN(new_n22023_));
  NOR3_X1    g18978(.A1(new_n21995_), .A2(pi0619), .A3(pi1159), .ZN(new_n22024_));
  NOR2_X1    g18979(.A1(new_n22024_), .A2(new_n11985_), .ZN(new_n22025_));
  XOR2_X1    g18980(.A1(new_n22023_), .A2(new_n22025_), .Z(new_n22026_));
  OAI21_X1   g18981(.A1(new_n22026_), .A2(new_n11997_), .B(new_n21997_), .ZN(new_n22027_));
  NOR2_X1    g18982(.A1(new_n21995_), .A2(new_n12054_), .ZN(new_n22028_));
  AOI21_X1   g18983(.A1(new_n22027_), .A2(new_n12054_), .B(new_n22028_), .ZN(new_n22029_));
  INV_X1     g18984(.I(new_n22029_), .ZN(new_n22030_));
  NOR2_X1    g18985(.A1(new_n21995_), .A2(new_n12092_), .ZN(new_n22031_));
  AOI21_X1   g18986(.A1(new_n22030_), .A2(new_n12092_), .B(new_n22031_), .ZN(new_n22032_));
  NAND2_X1   g18987(.A1(new_n22032_), .A2(new_n12082_), .ZN(new_n22033_));
  AOI21_X1   g18988(.A1(new_n21995_), .A2(pi0644), .B(new_n12099_), .ZN(new_n22034_));
  AOI21_X1   g18989(.A1(new_n22033_), .A2(new_n22034_), .B(pi1160), .ZN(new_n22035_));
  NOR2_X1    g18990(.A1(new_n21995_), .A2(new_n13114_), .ZN(new_n22036_));
  NOR2_X1    g18991(.A1(new_n21996_), .A2(new_n12014_), .ZN(new_n22037_));
  NOR2_X1    g18992(.A1(new_n21995_), .A2(new_n11961_), .ZN(new_n22038_));
  NAND2_X1   g18993(.A1(new_n11361_), .A2(new_n16303_), .ZN(new_n22039_));
  OAI21_X1   g18994(.A1(new_n12902_), .A2(new_n22039_), .B(new_n3231_), .ZN(new_n22040_));
  NOR3_X1    g18995(.A1(new_n13399_), .A2(pi0191), .A3(new_n13396_), .ZN(new_n22041_));
  AOI21_X1   g18996(.A1(new_n13399_), .A2(new_n11361_), .B(new_n13395_), .ZN(new_n22042_));
  NAND3_X1   g18997(.A1(new_n13403_), .A2(new_n3172_), .A3(new_n16303_), .ZN(new_n22043_));
  NOR4_X1    g18998(.A1(new_n22041_), .A2(new_n22042_), .A3(new_n22002_), .A4(new_n22043_), .ZN(new_n22044_));
  AOI22_X1   g18999(.A1(new_n22044_), .A2(new_n22040_), .B1(pi0191), .B2(new_n3232_), .ZN(new_n22045_));
  NAND2_X1   g19000(.A1(new_n22045_), .A2(new_n11891_), .ZN(new_n22046_));
  AOI21_X1   g19001(.A1(new_n22045_), .A2(new_n12970_), .B(new_n21996_), .ZN(new_n22047_));
  NOR3_X1    g19002(.A1(new_n22045_), .A2(pi0625), .A3(new_n21995_), .ZN(new_n22048_));
  NOR3_X1    g19003(.A1(new_n22048_), .A2(new_n22047_), .A3(pi1153), .ZN(new_n22049_));
  NAND4_X1   g19004(.A1(new_n22045_), .A2(pi0625), .A3(new_n11893_), .A4(new_n21996_), .ZN(new_n22050_));
  NAND2_X1   g19005(.A1(new_n22049_), .A2(new_n22050_), .ZN(new_n22051_));
  NAND2_X1   g19006(.A1(new_n22051_), .A2(pi0778), .ZN(new_n22052_));
  XOR2_X1    g19007(.A1(new_n22052_), .A2(new_n22046_), .Z(new_n22053_));
  NOR2_X1    g19008(.A1(new_n22053_), .A2(new_n13024_), .ZN(new_n22054_));
  AOI21_X1   g19009(.A1(new_n13024_), .A2(new_n21995_), .B(new_n22054_), .ZN(new_n22055_));
  AOI21_X1   g19010(.A1(new_n22055_), .A2(new_n11961_), .B(new_n22038_), .ZN(new_n22056_));
  AOI21_X1   g19011(.A1(new_n22056_), .A2(new_n12014_), .B(new_n22037_), .ZN(new_n22057_));
  AOI21_X1   g19012(.A1(new_n22057_), .A2(new_n13114_), .B(new_n22036_), .ZN(new_n22058_));
  NOR2_X1    g19013(.A1(new_n22058_), .A2(pi0628), .ZN(new_n22059_));
  AOI21_X1   g19014(.A1(pi0628), .A2(new_n21996_), .B(new_n22059_), .ZN(new_n22060_));
  NOR2_X1    g19015(.A1(new_n22060_), .A2(pi1156), .ZN(new_n22061_));
  NOR2_X1    g19016(.A1(new_n22058_), .A2(new_n12031_), .ZN(new_n22062_));
  AOI21_X1   g19017(.A1(new_n12031_), .A2(new_n21996_), .B(new_n22062_), .ZN(new_n22063_));
  NOR2_X1    g19018(.A1(new_n22063_), .A2(new_n12026_), .ZN(new_n22064_));
  OAI21_X1   g19019(.A1(new_n22061_), .A2(new_n22064_), .B(pi0792), .ZN(new_n22065_));
  OAI21_X1   g19020(.A1(pi0792), .A2(new_n22058_), .B(new_n22065_), .ZN(new_n22066_));
  NOR2_X1    g19021(.A1(new_n21995_), .A2(new_n12061_), .ZN(new_n22067_));
  AOI21_X1   g19022(.A1(new_n22066_), .A2(new_n12061_), .B(new_n22067_), .ZN(new_n22068_));
  NOR2_X1    g19023(.A1(new_n22068_), .A2(pi1157), .ZN(new_n22069_));
  NOR2_X1    g19024(.A1(new_n21995_), .A2(pi0647), .ZN(new_n22070_));
  AOI21_X1   g19025(.A1(new_n22066_), .A2(pi0647), .B(new_n22070_), .ZN(new_n22071_));
  NOR2_X1    g19026(.A1(new_n22071_), .A2(new_n12049_), .ZN(new_n22072_));
  NOR2_X1    g19027(.A1(new_n22069_), .A2(new_n22072_), .ZN(new_n22073_));
  NOR2_X1    g19028(.A1(new_n22073_), .A2(new_n12048_), .ZN(new_n22074_));
  AOI21_X1   g19029(.A1(new_n12048_), .A2(new_n22066_), .B(new_n22074_), .ZN(new_n22075_));
  NAND2_X1   g19030(.A1(new_n22075_), .A2(pi0644), .ZN(new_n22076_));
  AOI21_X1   g19031(.A1(new_n22076_), .A2(new_n12099_), .B(new_n22035_), .ZN(new_n22077_));
  NOR3_X1    g19032(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n22078_));
  NAND2_X1   g19033(.A1(new_n22032_), .A2(new_n22078_), .ZN(new_n22079_));
  NAND2_X1   g19034(.A1(new_n22079_), .A2(pi0715), .ZN(new_n22080_));
  AOI21_X1   g19035(.A1(new_n22075_), .A2(new_n12082_), .B(new_n22080_), .ZN(new_n22081_));
  OAI21_X1   g19036(.A1(new_n22077_), .A2(new_n22081_), .B(pi0790), .ZN(new_n22082_));
  NAND2_X1   g19037(.A1(new_n22035_), .A2(new_n12082_), .ZN(new_n22083_));
  AOI21_X1   g19038(.A1(new_n22079_), .A2(pi0644), .B(pi0790), .ZN(new_n22084_));
  NAND2_X1   g19039(.A1(new_n22083_), .A2(new_n22084_), .ZN(new_n22085_));
  NAND2_X1   g19040(.A1(new_n22071_), .A2(new_n12060_), .ZN(new_n22086_));
  AOI21_X1   g19041(.A1(new_n22068_), .A2(pi0630), .B(new_n12090_), .ZN(new_n22087_));
  NAND2_X1   g19042(.A1(new_n22030_), .A2(new_n15078_), .ZN(new_n22088_));
  AOI21_X1   g19043(.A1(new_n22087_), .A2(new_n22086_), .B(new_n22088_), .ZN(new_n22089_));
  AND2_X2    g19044(.A1(new_n22063_), .A2(new_n12030_), .Z(new_n22090_));
  NAND2_X1   g19045(.A1(new_n22060_), .A2(pi0629), .ZN(new_n22091_));
  NAND2_X1   g19046(.A1(new_n22091_), .A2(new_n17299_), .ZN(new_n22092_));
  OR2_X2     g19047(.A1(new_n22092_), .A2(new_n22090_), .Z(new_n22093_));
  NAND3_X1   g19048(.A1(new_n22093_), .A2(new_n17304_), .A3(new_n22027_), .ZN(new_n22094_));
  NAND2_X1   g19049(.A1(new_n22022_), .A2(pi0619), .ZN(new_n22095_));
  NAND2_X1   g19050(.A1(new_n21995_), .A2(pi0619), .ZN(new_n22096_));
  INV_X1     g19051(.I(new_n22005_), .ZN(new_n22097_));
  NAND2_X1   g19052(.A1(new_n17309_), .A2(new_n16270_), .ZN(new_n22098_));
  AOI21_X1   g19053(.A1(new_n12122_), .A2(new_n22098_), .B(pi0039), .ZN(new_n22099_));
  AOI21_X1   g19054(.A1(new_n13644_), .A2(new_n21910_), .B(new_n11361_), .ZN(new_n22100_));
  AOI21_X1   g19055(.A1(new_n22100_), .A2(new_n5156_), .B(new_n3172_), .ZN(new_n22101_));
  OAI21_X1   g19056(.A1(new_n22099_), .A2(pi0191), .B(new_n22101_), .ZN(new_n22102_));
  NOR2_X1    g19057(.A1(new_n13333_), .A2(new_n11361_), .ZN(new_n22103_));
  OAI21_X1   g19058(.A1(new_n12515_), .A2(new_n11361_), .B(new_n16270_), .ZN(new_n22104_));
  NOR3_X1    g19059(.A1(new_n12645_), .A2(new_n11361_), .A3(new_n13347_), .ZN(new_n22105_));
  AOI21_X1   g19060(.A1(new_n12645_), .A2(pi0191), .B(new_n12665_), .ZN(new_n22106_));
  OAI21_X1   g19061(.A1(new_n22105_), .A2(new_n22106_), .B(pi0746), .ZN(new_n22107_));
  NAND2_X1   g19062(.A1(new_n13360_), .A2(pi0191), .ZN(new_n22108_));
  NAND2_X1   g19063(.A1(new_n13362_), .A2(pi0191), .ZN(new_n22109_));
  NAND4_X1   g19064(.A1(new_n22107_), .A2(new_n16290_), .A3(new_n22108_), .A4(new_n22109_), .ZN(new_n22110_));
  AOI21_X1   g19065(.A1(new_n22110_), .A2(new_n3172_), .B(pi0039), .ZN(new_n22111_));
  OAI21_X1   g19066(.A1(new_n22103_), .A2(new_n22104_), .B(new_n22111_), .ZN(new_n22112_));
  NAND2_X1   g19067(.A1(new_n3232_), .A2(new_n16303_), .ZN(new_n22113_));
  AOI21_X1   g19068(.A1(new_n22112_), .A2(new_n22102_), .B(new_n22113_), .ZN(new_n22114_));
  NAND2_X1   g19069(.A1(new_n22001_), .A2(new_n22003_), .ZN(new_n22115_));
  NAND2_X1   g19070(.A1(new_n22115_), .A2(new_n16303_), .ZN(new_n22116_));
  OAI22_X1   g19071(.A1(new_n22114_), .A2(new_n22116_), .B1(new_n11361_), .B2(new_n3231_), .ZN(new_n22117_));
  OAI21_X1   g19072(.A1(new_n22117_), .A2(pi0625), .B(new_n22097_), .ZN(new_n22118_));
  NAND3_X1   g19073(.A1(new_n22117_), .A2(new_n12970_), .A3(new_n22005_), .ZN(new_n22119_));
  NAND4_X1   g19074(.A1(new_n22118_), .A2(new_n22119_), .A3(new_n12977_), .A4(new_n22050_), .ZN(new_n22120_));
  INV_X1     g19075(.I(new_n22049_), .ZN(new_n22121_));
  NOR4_X1    g19076(.A1(new_n22117_), .A2(new_n12970_), .A3(pi1153), .A4(new_n22097_), .ZN(new_n22122_));
  OAI21_X1   g19077(.A1(new_n22122_), .A2(new_n22121_), .B(new_n13657_), .ZN(new_n22123_));
  NAND2_X1   g19078(.A1(new_n22120_), .A2(new_n22123_), .ZN(new_n22124_));
  NOR2_X1    g19079(.A1(new_n22117_), .A2(pi0778), .ZN(new_n22125_));
  AOI21_X1   g19080(.A1(new_n22124_), .A2(pi0778), .B(new_n22125_), .ZN(new_n22126_));
  NOR2_X1    g19081(.A1(new_n22126_), .A2(pi0785), .ZN(new_n22127_));
  INV_X1     g19082(.I(new_n22053_), .ZN(new_n22128_));
  NAND3_X1   g19083(.A1(new_n22128_), .A2(pi0609), .A3(pi1155), .ZN(new_n22129_));
  NAND3_X1   g19084(.A1(new_n22129_), .A2(new_n11923_), .A3(new_n22012_), .ZN(new_n22130_));
  NOR4_X1    g19085(.A1(new_n22126_), .A2(new_n11903_), .A3(new_n22128_), .A4(pi1155), .ZN(new_n22131_));
  NAND2_X1   g19086(.A1(new_n22010_), .A2(pi0660), .ZN(new_n22132_));
  NOR2_X1    g19087(.A1(new_n22131_), .A2(new_n22132_), .ZN(new_n22133_));
  NOR2_X1    g19088(.A1(new_n22133_), .A2(new_n11870_), .ZN(new_n22134_));
  AOI21_X1   g19089(.A1(new_n22134_), .A2(new_n22130_), .B(new_n22127_), .ZN(new_n22135_));
  INV_X1     g19090(.I(new_n22055_), .ZN(new_n22136_));
  NOR4_X1    g19091(.A1(new_n22135_), .A2(new_n11934_), .A3(pi1154), .A4(new_n22136_), .ZN(new_n22137_));
  NAND2_X1   g19092(.A1(new_n22017_), .A2(pi0627), .ZN(new_n22138_));
  NOR3_X1    g19093(.A1(new_n22055_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n22139_));
  NAND2_X1   g19094(.A1(new_n22020_), .A2(new_n11949_), .ZN(new_n22140_));
  OAI22_X1   g19095(.A1(new_n22137_), .A2(new_n22138_), .B1(new_n22139_), .B2(new_n22140_), .ZN(new_n22141_));
  MUX2_X1    g19096(.I0(new_n22141_), .I1(new_n22135_), .S(new_n11969_), .Z(new_n22142_));
  XNOR2_X1   g19097(.A1(new_n22142_), .A2(new_n22056_), .ZN(new_n22143_));
  NOR2_X1    g19098(.A1(new_n22143_), .A2(new_n11967_), .ZN(new_n22144_));
  NAND3_X1   g19099(.A1(new_n22095_), .A2(new_n11869_), .A3(new_n22096_), .ZN(new_n22145_));
  XOR2_X1    g19100(.A1(new_n22144_), .A2(new_n22142_), .Z(new_n22146_));
  AOI21_X1   g19101(.A1(new_n21996_), .A2(new_n11967_), .B(pi1159), .ZN(new_n22147_));
  AOI21_X1   g19102(.A1(new_n22095_), .A2(new_n22147_), .B(pi0648), .ZN(new_n22148_));
  OAI21_X1   g19103(.A1(new_n22146_), .A2(pi1159), .B(new_n22148_), .ZN(new_n22149_));
  OR2_X2     g19104(.A1(new_n22142_), .A2(pi0789), .Z(new_n22150_));
  NAND3_X1   g19105(.A1(new_n22026_), .A2(pi0626), .A3(new_n21996_), .ZN(new_n22151_));
  OAI21_X1   g19106(.A1(new_n22026_), .A2(new_n11994_), .B(new_n21995_), .ZN(new_n22152_));
  AOI21_X1   g19107(.A1(new_n22152_), .A2(new_n22151_), .B(new_n17167_), .ZN(new_n22153_));
  AOI21_X1   g19108(.A1(new_n22026_), .A2(new_n21996_), .B(new_n11994_), .ZN(new_n22154_));
  NAND2_X1   g19109(.A1(new_n22154_), .A2(new_n11990_), .ZN(new_n22155_));
  NOR2_X1    g19110(.A1(new_n22057_), .A2(new_n12020_), .ZN(new_n22156_));
  NOR2_X1    g19111(.A1(new_n22156_), .A2(pi0788), .ZN(new_n22157_));
  NAND2_X1   g19112(.A1(new_n22155_), .A2(new_n22157_), .ZN(new_n22158_));
  OAI21_X1   g19113(.A1(new_n22158_), .A2(new_n22153_), .B(new_n17372_), .ZN(new_n22159_));
  AOI21_X1   g19114(.A1(new_n11998_), .A2(new_n22150_), .B(new_n22159_), .ZN(new_n22160_));
  NAND3_X1   g19115(.A1(new_n22149_), .A2(new_n22145_), .A3(new_n22160_), .ZN(new_n22161_));
  AOI21_X1   g19116(.A1(new_n22161_), .A2(new_n22094_), .B(new_n14725_), .ZN(new_n22162_));
  OAI21_X1   g19117(.A1(new_n22162_), .A2(new_n22089_), .B(new_n22085_), .ZN(new_n22163_));
  AOI21_X1   g19118(.A1(new_n22082_), .A2(new_n22163_), .B(po1038), .ZN(new_n22164_));
  OAI21_X1   g19119(.A1(new_n6845_), .A2(pi0191), .B(new_n13184_), .ZN(new_n22165_));
  OAI21_X1   g19120(.A1(new_n22164_), .A2(new_n22165_), .B(new_n21994_), .ZN(po0348));
  NOR2_X1    g19121(.A1(new_n2925_), .A2(pi0192), .ZN(new_n22167_));
  NOR2_X1    g19122(.A1(new_n11877_), .A2(new_n16368_), .ZN(new_n22168_));
  NOR2_X1    g19123(.A1(new_n22168_), .A2(new_n22167_), .ZN(new_n22169_));
  AOI21_X1   g19124(.A1(new_n11886_), .A2(pi0691), .B(new_n22167_), .ZN(new_n22170_));
  NOR2_X1    g19125(.A1(new_n22170_), .A2(new_n11874_), .ZN(new_n22171_));
  INV_X1     g19126(.I(new_n22171_), .ZN(new_n22172_));
  NAND2_X1   g19127(.A1(new_n22172_), .A2(new_n22169_), .ZN(new_n22173_));
  NAND2_X1   g19128(.A1(new_n22173_), .A2(new_n11891_), .ZN(new_n22174_));
  NOR2_X1    g19129(.A1(new_n22172_), .A2(new_n12970_), .ZN(new_n22175_));
  NOR4_X1    g19130(.A1(new_n22175_), .A2(new_n11893_), .A3(new_n22167_), .A4(new_n22168_), .ZN(new_n22176_));
  NOR2_X1    g19131(.A1(new_n13201_), .A2(new_n16401_), .ZN(new_n22177_));
  NOR2_X1    g19132(.A1(new_n22167_), .A2(pi1153), .ZN(new_n22178_));
  INV_X1     g19133(.I(new_n22178_), .ZN(new_n22179_));
  NOR2_X1    g19134(.A1(new_n22177_), .A2(new_n22179_), .ZN(new_n22180_));
  INV_X1     g19135(.I(new_n22180_), .ZN(new_n22181_));
  NAND2_X1   g19136(.A1(new_n22181_), .A2(pi0608), .ZN(new_n22182_));
  INV_X1     g19137(.I(new_n22175_), .ZN(new_n22183_));
  AOI21_X1   g19138(.A1(new_n22183_), .A2(new_n22173_), .B(new_n22179_), .ZN(new_n22184_));
  OAI21_X1   g19139(.A1(new_n22177_), .A2(new_n22170_), .B(pi1153), .ZN(new_n22185_));
  NAND2_X1   g19140(.A1(new_n22185_), .A2(new_n13657_), .ZN(new_n22186_));
  OAI22_X1   g19141(.A1(new_n22182_), .A2(new_n22176_), .B1(new_n22184_), .B2(new_n22186_), .ZN(new_n22187_));
  NAND2_X1   g19142(.A1(new_n22187_), .A2(pi0778), .ZN(new_n22188_));
  XOR2_X1    g19143(.A1(new_n22188_), .A2(new_n22174_), .Z(new_n22189_));
  INV_X1     g19144(.I(new_n22189_), .ZN(new_n22190_));
  NAND2_X1   g19145(.A1(new_n22181_), .A2(new_n22185_), .ZN(new_n22191_));
  MUX2_X1    g19146(.I0(new_n22191_), .I1(new_n22170_), .S(new_n11891_), .Z(new_n22192_));
  XNOR2_X1   g19147(.A1(new_n22189_), .A2(new_n22192_), .ZN(new_n22193_));
  NAND2_X1   g19148(.A1(new_n22193_), .A2(pi0609), .ZN(new_n22194_));
  XOR2_X1    g19149(.A1(new_n22194_), .A2(new_n22190_), .Z(new_n22195_));
  INV_X1     g19150(.I(new_n22168_), .ZN(new_n22196_));
  NOR2_X1    g19151(.A1(new_n22169_), .A2(new_n11925_), .ZN(new_n22197_));
  NOR4_X1    g19152(.A1(new_n22197_), .A2(pi1155), .A3(new_n12997_), .A4(new_n22196_), .ZN(new_n22198_));
  NOR2_X1    g19153(.A1(new_n22198_), .A2(pi0660), .ZN(new_n22199_));
  OAI21_X1   g19154(.A1(new_n22195_), .A2(pi1155), .B(new_n22199_), .ZN(new_n22200_));
  NOR2_X1    g19155(.A1(new_n22196_), .A2(new_n12997_), .ZN(new_n22201_));
  NOR4_X1    g19156(.A1(new_n22201_), .A2(new_n11923_), .A3(pi1155), .A4(new_n22167_), .ZN(new_n22203_));
  NOR2_X1    g19157(.A1(new_n22203_), .A2(new_n11870_), .ZN(new_n22204_));
  AOI22_X1   g19158(.A1(new_n22200_), .A2(new_n22204_), .B1(new_n11870_), .B2(new_n22190_), .ZN(new_n22205_));
  NOR2_X1    g19159(.A1(new_n22205_), .A2(pi0781), .ZN(new_n22206_));
  NOR4_X1    g19160(.A1(new_n22192_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n22207_));
  NOR2_X1    g19161(.A1(new_n22197_), .A2(pi0785), .ZN(new_n22208_));
  NOR4_X1    g19162(.A1(new_n22198_), .A2(pi1155), .A3(new_n22167_), .A4(new_n22201_), .ZN(new_n22209_));
  NOR2_X1    g19163(.A1(new_n22209_), .A2(new_n11870_), .ZN(new_n22210_));
  XOR2_X1    g19164(.A1(new_n22210_), .A2(new_n22208_), .Z(new_n22211_));
  INV_X1     g19165(.I(new_n22211_), .ZN(new_n22212_));
  OAI21_X1   g19166(.A1(new_n22212_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n22213_));
  OAI21_X1   g19167(.A1(new_n22212_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n22214_));
  NOR2_X1    g19168(.A1(new_n22192_), .A2(new_n11939_), .ZN(new_n22215_));
  NOR4_X1    g19169(.A1(new_n22205_), .A2(new_n11934_), .A3(pi1154), .A4(new_n22215_), .ZN(new_n22216_));
  NOR2_X1    g19170(.A1(new_n22216_), .A2(new_n22214_), .ZN(new_n22217_));
  OAI22_X1   g19171(.A1(new_n22217_), .A2(pi0627), .B1(new_n22207_), .B2(new_n22213_), .ZN(new_n22218_));
  AOI21_X1   g19172(.A1(new_n22218_), .A2(pi0781), .B(new_n22206_), .ZN(new_n22219_));
  INV_X1     g19173(.I(new_n22215_), .ZN(new_n22220_));
  NOR2_X1    g19174(.A1(new_n22220_), .A2(new_n11962_), .ZN(new_n22221_));
  NOR4_X1    g19175(.A1(new_n22219_), .A2(new_n11967_), .A3(pi1159), .A4(new_n22221_), .ZN(new_n22222_));
  NOR2_X1    g19176(.A1(new_n22212_), .A2(pi0781), .ZN(new_n22223_));
  AOI21_X1   g19177(.A1(new_n11944_), .A2(new_n22211_), .B(new_n22214_), .ZN(new_n22224_));
  NOR2_X1    g19178(.A1(new_n22224_), .A2(new_n11969_), .ZN(new_n22225_));
  XOR2_X1    g19179(.A1(new_n22225_), .A2(new_n22223_), .Z(new_n22226_));
  AOI21_X1   g19180(.A1(new_n22226_), .A2(new_n16479_), .B(pi1159), .ZN(new_n22227_));
  INV_X1     g19181(.I(new_n22227_), .ZN(new_n22228_));
  NOR3_X1    g19182(.A1(new_n22222_), .A2(new_n11966_), .A3(new_n22228_), .ZN(new_n22229_));
  NOR4_X1    g19183(.A1(new_n22220_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n22230_));
  INV_X1     g19184(.I(new_n22226_), .ZN(new_n22231_));
  NOR2_X1    g19185(.A1(new_n22231_), .A2(new_n16482_), .ZN(new_n22232_));
  NOR3_X1    g19186(.A1(new_n22232_), .A2(pi0648), .A3(new_n22230_), .ZN(new_n22233_));
  AOI21_X1   g19187(.A1(new_n22219_), .A2(new_n11998_), .B(pi0789), .ZN(new_n22234_));
  OAI21_X1   g19188(.A1(new_n22229_), .A2(new_n22233_), .B(new_n22234_), .ZN(new_n22235_));
  NOR3_X1    g19189(.A1(new_n22220_), .A2(new_n11962_), .A3(new_n12015_), .ZN(new_n22236_));
  NAND2_X1   g19190(.A1(new_n22236_), .A2(new_n17154_), .ZN(new_n22237_));
  NOR2_X1    g19191(.A1(new_n14624_), .A2(new_n22167_), .ZN(new_n22238_));
  OAI21_X1   g19192(.A1(new_n16482_), .A2(new_n22231_), .B(new_n22227_), .ZN(new_n22239_));
  MUX2_X1    g19193(.I0(new_n22239_), .I1(new_n22226_), .S(new_n11985_), .Z(new_n22240_));
  AOI21_X1   g19194(.A1(new_n22240_), .A2(new_n14624_), .B(new_n22238_), .ZN(new_n22241_));
  INV_X1     g19195(.I(new_n22241_), .ZN(new_n22242_));
  OAI22_X1   g19196(.A1(new_n22242_), .A2(new_n17150_), .B1(new_n17151_), .B2(new_n22237_), .ZN(new_n22243_));
  NAND2_X1   g19197(.A1(new_n22243_), .A2(pi0629), .ZN(new_n22244_));
  OAI21_X1   g19198(.A1(new_n22237_), .A2(new_n17163_), .B(new_n15085_), .ZN(new_n22245_));
  AOI21_X1   g19199(.A1(new_n22241_), .A2(new_n12063_), .B(new_n22245_), .ZN(new_n22246_));
  NAND2_X1   g19200(.A1(new_n22244_), .A2(new_n22246_), .ZN(new_n22247_));
  INV_X1     g19201(.I(new_n22167_), .ZN(new_n22248_));
  MUX2_X1    g19202(.I0(new_n22240_), .I1(new_n22248_), .S(new_n11994_), .Z(new_n22249_));
  NOR2_X1    g19203(.A1(new_n22249_), .A2(new_n17167_), .ZN(new_n22250_));
  OAI21_X1   g19204(.A1(new_n22240_), .A2(new_n22167_), .B(pi0626), .ZN(new_n22251_));
  AOI21_X1   g19205(.A1(new_n22236_), .A2(new_n17173_), .B(pi0788), .ZN(new_n22252_));
  OAI21_X1   g19206(.A1(new_n22251_), .A2(new_n17171_), .B(new_n22252_), .ZN(new_n22253_));
  OAI21_X1   g19207(.A1(new_n22250_), .A2(new_n22253_), .B(new_n14732_), .ZN(new_n22254_));
  AOI21_X1   g19208(.A1(new_n22247_), .A2(new_n14726_), .B(new_n22254_), .ZN(new_n22255_));
  NAND3_X1   g19209(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n22167_), .ZN(new_n22256_));
  NOR2_X1    g19210(.A1(new_n22237_), .A2(new_n12068_), .ZN(new_n22257_));
  AOI21_X1   g19211(.A1(new_n22167_), .A2(pi0647), .B(pi1157), .ZN(new_n22258_));
  OAI21_X1   g19212(.A1(new_n22257_), .A2(new_n12061_), .B(new_n22258_), .ZN(new_n22259_));
  NOR2_X1    g19213(.A1(new_n22248_), .A2(pi0647), .ZN(new_n22260_));
  AOI21_X1   g19214(.A1(new_n22257_), .A2(pi0647), .B(new_n22260_), .ZN(new_n22261_));
  NAND2_X1   g19215(.A1(new_n22261_), .A2(new_n12088_), .ZN(new_n22262_));
  NAND2_X1   g19216(.A1(new_n22262_), .A2(pi0787), .ZN(new_n22263_));
  AOI21_X1   g19217(.A1(pi0630), .A2(new_n22259_), .B(new_n22263_), .ZN(new_n22264_));
  AOI22_X1   g19218(.A1(new_n22235_), .A2(new_n22255_), .B1(new_n22256_), .B2(new_n22264_), .ZN(new_n22265_));
  OR2_X2     g19219(.A1(new_n22265_), .A2(new_n12082_), .Z(new_n22266_));
  MUX2_X1    g19220(.I0(new_n22242_), .I1(new_n22248_), .S(new_n16841_), .Z(new_n22267_));
  MUX2_X1    g19221(.I0(new_n22267_), .I1(new_n22248_), .S(pi0644), .Z(new_n22268_));
  NAND2_X1   g19222(.A1(new_n22261_), .A2(pi1157), .ZN(new_n22269_));
  NOR2_X1    g19223(.A1(new_n22259_), .A2(new_n12048_), .ZN(new_n22270_));
  AOI22_X1   g19224(.A1(new_n22270_), .A2(new_n22269_), .B1(new_n12048_), .B2(new_n22257_), .ZN(new_n22271_));
  OAI21_X1   g19225(.A1(new_n22271_), .A2(new_n12082_), .B(new_n13168_), .ZN(new_n22272_));
  AOI21_X1   g19226(.A1(new_n22268_), .A2(pi0715), .B(new_n22272_), .ZN(new_n22273_));
  AOI21_X1   g19227(.A1(new_n22271_), .A2(new_n12082_), .B(pi0715), .ZN(new_n22274_));
  NAND2_X1   g19228(.A1(new_n22266_), .A2(new_n22274_), .ZN(new_n22275_));
  NAND3_X1   g19229(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n22276_));
  NOR2_X1    g19230(.A1(new_n22267_), .A2(new_n22276_), .ZN(new_n22277_));
  AOI22_X1   g19231(.A1(new_n22275_), .A2(new_n22277_), .B1(new_n22266_), .B2(new_n22273_), .ZN(new_n22278_));
  AOI21_X1   g19232(.A1(new_n22265_), .A2(new_n11867_), .B(new_n13184_), .ZN(new_n22279_));
  OAI21_X1   g19233(.A1(new_n22278_), .A2(new_n11867_), .B(new_n22279_), .ZN(new_n22280_));
  NOR2_X1    g19234(.A1(new_n12965_), .A2(pi0192), .ZN(new_n22281_));
  INV_X1     g19235(.I(new_n22281_), .ZN(new_n22282_));
  NAND2_X1   g19236(.A1(new_n22282_), .A2(new_n11997_), .ZN(new_n22283_));
  NOR2_X1    g19237(.A1(new_n16368_), .A2(pi0192), .ZN(new_n22284_));
  OAI21_X1   g19238(.A1(new_n14361_), .A2(new_n11572_), .B(pi0039), .ZN(new_n22285_));
  AOI21_X1   g19239(.A1(new_n13381_), .A2(new_n22284_), .B(new_n22285_), .ZN(new_n22286_));
  OAI21_X1   g19240(.A1(pi0764), .A2(new_n12793_), .B(new_n22286_), .ZN(new_n22287_));
  NOR2_X1    g19241(.A1(new_n12828_), .A2(pi0192), .ZN(new_n22288_));
  AOI21_X1   g19242(.A1(new_n12829_), .A2(pi0764), .B(pi0038), .ZN(new_n22289_));
  AOI21_X1   g19243(.A1(new_n22287_), .A2(new_n22289_), .B(new_n3232_), .ZN(new_n22290_));
  AOI21_X1   g19244(.A1(new_n11572_), .A2(new_n3232_), .B(new_n22290_), .ZN(new_n22291_));
  OAI21_X1   g19245(.A1(new_n22291_), .A2(new_n11914_), .B(new_n11870_), .ZN(new_n22292_));
  AOI21_X1   g19246(.A1(new_n11914_), .A2(new_n22281_), .B(new_n22292_), .ZN(new_n22293_));
  NAND2_X1   g19247(.A1(new_n22291_), .A2(new_n11924_), .ZN(new_n22294_));
  OAI22_X1   g19248(.A1(new_n22294_), .A2(pi0609), .B1(new_n12996_), .B2(new_n22281_), .ZN(new_n22295_));
  NAND2_X1   g19249(.A1(new_n22295_), .A2(new_n11912_), .ZN(new_n22296_));
  OAI22_X1   g19250(.A1(new_n22294_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n22281_), .ZN(new_n22297_));
  NAND2_X1   g19251(.A1(new_n22297_), .A2(pi1155), .ZN(new_n22298_));
  NAND2_X1   g19252(.A1(new_n22296_), .A2(new_n22298_), .ZN(new_n22299_));
  NAND2_X1   g19253(.A1(new_n22299_), .A2(pi0785), .ZN(new_n22300_));
  XNOR2_X1   g19254(.A1(new_n22300_), .A2(new_n22293_), .ZN(new_n22301_));
  OAI21_X1   g19255(.A1(new_n22282_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n22302_));
  AOI21_X1   g19256(.A1(new_n22301_), .A2(pi0618), .B(new_n22302_), .ZN(new_n22303_));
  INV_X1     g19257(.I(new_n22301_), .ZN(new_n22304_));
  AOI21_X1   g19258(.A1(new_n22282_), .A2(new_n11934_), .B(pi1154), .ZN(new_n22305_));
  OAI21_X1   g19259(.A1(new_n22304_), .A2(new_n11934_), .B(new_n22305_), .ZN(new_n22306_));
  NAND2_X1   g19260(.A1(new_n22306_), .A2(new_n22303_), .ZN(new_n22307_));
  MUX2_X1    g19261(.I0(new_n22307_), .I1(new_n22301_), .S(new_n11969_), .Z(new_n22308_));
  NAND2_X1   g19262(.A1(new_n22308_), .A2(new_n11985_), .ZN(new_n22309_));
  NOR3_X1    g19263(.A1(new_n22281_), .A2(pi0619), .A3(pi1159), .ZN(new_n22310_));
  NOR2_X1    g19264(.A1(new_n22310_), .A2(new_n11985_), .ZN(new_n22311_));
  XOR2_X1    g19265(.A1(new_n22309_), .A2(new_n22311_), .Z(new_n22312_));
  OAI21_X1   g19266(.A1(new_n22312_), .A2(new_n11997_), .B(new_n22283_), .ZN(new_n22313_));
  NOR2_X1    g19267(.A1(new_n22281_), .A2(new_n12054_), .ZN(new_n22314_));
  AOI21_X1   g19268(.A1(new_n22313_), .A2(new_n12054_), .B(new_n22314_), .ZN(new_n22315_));
  INV_X1     g19269(.I(new_n22315_), .ZN(new_n22316_));
  NOR2_X1    g19270(.A1(new_n22281_), .A2(new_n12092_), .ZN(new_n22317_));
  AOI21_X1   g19271(.A1(new_n22316_), .A2(new_n12092_), .B(new_n22317_), .ZN(new_n22318_));
  NAND2_X1   g19272(.A1(new_n22318_), .A2(new_n12082_), .ZN(new_n22319_));
  AOI21_X1   g19273(.A1(new_n22281_), .A2(pi0644), .B(new_n12099_), .ZN(new_n22320_));
  AOI21_X1   g19274(.A1(new_n22319_), .A2(new_n22320_), .B(pi1160), .ZN(new_n22321_));
  NOR2_X1    g19275(.A1(new_n22281_), .A2(new_n13114_), .ZN(new_n22322_));
  NOR2_X1    g19276(.A1(new_n22282_), .A2(new_n12014_), .ZN(new_n22323_));
  NOR2_X1    g19277(.A1(new_n22281_), .A2(new_n11961_), .ZN(new_n22324_));
  NAND2_X1   g19278(.A1(new_n11572_), .A2(new_n16401_), .ZN(new_n22325_));
  OAI21_X1   g19279(.A1(new_n12902_), .A2(new_n22325_), .B(new_n3231_), .ZN(new_n22326_));
  NOR3_X1    g19280(.A1(new_n13399_), .A2(pi0192), .A3(new_n13396_), .ZN(new_n22327_));
  AOI21_X1   g19281(.A1(new_n13399_), .A2(new_n11572_), .B(new_n13395_), .ZN(new_n22328_));
  NAND3_X1   g19282(.A1(new_n13403_), .A2(new_n3172_), .A3(new_n16401_), .ZN(new_n22329_));
  NOR4_X1    g19283(.A1(new_n22327_), .A2(new_n22328_), .A3(new_n22288_), .A4(new_n22329_), .ZN(new_n22330_));
  AOI22_X1   g19284(.A1(new_n22330_), .A2(new_n22326_), .B1(pi0192), .B2(new_n3232_), .ZN(new_n22331_));
  NAND2_X1   g19285(.A1(new_n22331_), .A2(new_n11891_), .ZN(new_n22332_));
  AOI21_X1   g19286(.A1(new_n22331_), .A2(new_n12970_), .B(new_n22282_), .ZN(new_n22333_));
  NOR3_X1    g19287(.A1(new_n22331_), .A2(pi0625), .A3(new_n22281_), .ZN(new_n22334_));
  NOR3_X1    g19288(.A1(new_n22334_), .A2(new_n22333_), .A3(pi1153), .ZN(new_n22335_));
  NAND4_X1   g19289(.A1(new_n22331_), .A2(pi0625), .A3(new_n11893_), .A4(new_n22282_), .ZN(new_n22336_));
  NAND2_X1   g19290(.A1(new_n22335_), .A2(new_n22336_), .ZN(new_n22337_));
  NAND2_X1   g19291(.A1(new_n22337_), .A2(pi0778), .ZN(new_n22338_));
  XOR2_X1    g19292(.A1(new_n22338_), .A2(new_n22332_), .Z(new_n22339_));
  NOR2_X1    g19293(.A1(new_n22339_), .A2(new_n13024_), .ZN(new_n22340_));
  AOI21_X1   g19294(.A1(new_n13024_), .A2(new_n22281_), .B(new_n22340_), .ZN(new_n22341_));
  AOI21_X1   g19295(.A1(new_n22341_), .A2(new_n11961_), .B(new_n22324_), .ZN(new_n22342_));
  AOI21_X1   g19296(.A1(new_n22342_), .A2(new_n12014_), .B(new_n22323_), .ZN(new_n22343_));
  AOI21_X1   g19297(.A1(new_n22343_), .A2(new_n13114_), .B(new_n22322_), .ZN(new_n22344_));
  NOR2_X1    g19298(.A1(new_n22344_), .A2(pi0628), .ZN(new_n22345_));
  AOI21_X1   g19299(.A1(pi0628), .A2(new_n22282_), .B(new_n22345_), .ZN(new_n22346_));
  NOR2_X1    g19300(.A1(new_n22346_), .A2(pi1156), .ZN(new_n22347_));
  NOR2_X1    g19301(.A1(new_n22344_), .A2(new_n12031_), .ZN(new_n22348_));
  AOI21_X1   g19302(.A1(new_n12031_), .A2(new_n22282_), .B(new_n22348_), .ZN(new_n22349_));
  NOR2_X1    g19303(.A1(new_n22349_), .A2(new_n12026_), .ZN(new_n22350_));
  OAI21_X1   g19304(.A1(new_n22347_), .A2(new_n22350_), .B(pi0792), .ZN(new_n22351_));
  OAI21_X1   g19305(.A1(pi0792), .A2(new_n22344_), .B(new_n22351_), .ZN(new_n22352_));
  NOR2_X1    g19306(.A1(new_n22281_), .A2(new_n12061_), .ZN(new_n22353_));
  AOI21_X1   g19307(.A1(new_n22352_), .A2(new_n12061_), .B(new_n22353_), .ZN(new_n22354_));
  NOR2_X1    g19308(.A1(new_n22354_), .A2(pi1157), .ZN(new_n22355_));
  NOR2_X1    g19309(.A1(new_n22281_), .A2(pi0647), .ZN(new_n22356_));
  AOI21_X1   g19310(.A1(new_n22352_), .A2(pi0647), .B(new_n22356_), .ZN(new_n22357_));
  NOR2_X1    g19311(.A1(new_n22357_), .A2(new_n12049_), .ZN(new_n22358_));
  NOR2_X1    g19312(.A1(new_n22355_), .A2(new_n22358_), .ZN(new_n22359_));
  NOR2_X1    g19313(.A1(new_n22359_), .A2(new_n12048_), .ZN(new_n22360_));
  AOI21_X1   g19314(.A1(new_n12048_), .A2(new_n22352_), .B(new_n22360_), .ZN(new_n22361_));
  NAND2_X1   g19315(.A1(new_n22361_), .A2(pi0644), .ZN(new_n22362_));
  AOI21_X1   g19316(.A1(new_n22362_), .A2(new_n12099_), .B(new_n22321_), .ZN(new_n22363_));
  NOR3_X1    g19317(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n22364_));
  NAND2_X1   g19318(.A1(new_n22318_), .A2(new_n22364_), .ZN(new_n22365_));
  NAND2_X1   g19319(.A1(new_n22365_), .A2(pi0715), .ZN(new_n22366_));
  AOI21_X1   g19320(.A1(new_n22361_), .A2(new_n12082_), .B(new_n22366_), .ZN(new_n22367_));
  OAI21_X1   g19321(.A1(new_n22363_), .A2(new_n22367_), .B(pi0790), .ZN(new_n22368_));
  NAND2_X1   g19322(.A1(new_n22321_), .A2(new_n12082_), .ZN(new_n22369_));
  AOI21_X1   g19323(.A1(new_n22365_), .A2(pi0644), .B(pi0790), .ZN(new_n22370_));
  NAND2_X1   g19324(.A1(new_n22369_), .A2(new_n22370_), .ZN(new_n22371_));
  NAND2_X1   g19325(.A1(new_n22357_), .A2(new_n12060_), .ZN(new_n22372_));
  AOI21_X1   g19326(.A1(new_n22354_), .A2(pi0630), .B(new_n12090_), .ZN(new_n22373_));
  NAND2_X1   g19327(.A1(new_n22316_), .A2(new_n15078_), .ZN(new_n22374_));
  AOI21_X1   g19328(.A1(new_n22373_), .A2(new_n22372_), .B(new_n22374_), .ZN(new_n22375_));
  AND2_X2    g19329(.A1(new_n22349_), .A2(new_n12030_), .Z(new_n22376_));
  NAND2_X1   g19330(.A1(new_n22346_), .A2(pi0629), .ZN(new_n22377_));
  NAND2_X1   g19331(.A1(new_n22377_), .A2(new_n17299_), .ZN(new_n22378_));
  OR2_X2     g19332(.A1(new_n22378_), .A2(new_n22376_), .Z(new_n22379_));
  NAND3_X1   g19333(.A1(new_n22379_), .A2(new_n17304_), .A3(new_n22313_), .ZN(new_n22380_));
  NAND2_X1   g19334(.A1(new_n22308_), .A2(pi0619), .ZN(new_n22381_));
  NAND2_X1   g19335(.A1(new_n22281_), .A2(pi0619), .ZN(new_n22382_));
  INV_X1     g19336(.I(new_n22291_), .ZN(new_n22383_));
  NAND2_X1   g19337(.A1(new_n17309_), .A2(new_n16368_), .ZN(new_n22384_));
  AOI21_X1   g19338(.A1(new_n12122_), .A2(new_n22384_), .B(pi0039), .ZN(new_n22385_));
  AOI21_X1   g19339(.A1(new_n13644_), .A2(new_n22196_), .B(new_n11572_), .ZN(new_n22386_));
  AOI21_X1   g19340(.A1(new_n22386_), .A2(new_n5156_), .B(new_n3172_), .ZN(new_n22387_));
  OAI21_X1   g19341(.A1(new_n22385_), .A2(pi0192), .B(new_n22387_), .ZN(new_n22388_));
  NOR2_X1    g19342(.A1(new_n13333_), .A2(new_n11572_), .ZN(new_n22389_));
  OAI21_X1   g19343(.A1(new_n12515_), .A2(new_n11572_), .B(new_n16368_), .ZN(new_n22390_));
  NOR3_X1    g19344(.A1(new_n12645_), .A2(new_n11572_), .A3(new_n13347_), .ZN(new_n22391_));
  AOI21_X1   g19345(.A1(new_n12645_), .A2(pi0192), .B(new_n12665_), .ZN(new_n22392_));
  OAI21_X1   g19346(.A1(new_n22391_), .A2(new_n22392_), .B(pi0764), .ZN(new_n22393_));
  NAND2_X1   g19347(.A1(new_n13360_), .A2(pi0192), .ZN(new_n22394_));
  NAND2_X1   g19348(.A1(new_n13362_), .A2(pi0192), .ZN(new_n22395_));
  NAND4_X1   g19349(.A1(new_n22393_), .A2(new_n16388_), .A3(new_n22394_), .A4(new_n22395_), .ZN(new_n22396_));
  AOI21_X1   g19350(.A1(new_n22396_), .A2(new_n3172_), .B(pi0039), .ZN(new_n22397_));
  OAI21_X1   g19351(.A1(new_n22389_), .A2(new_n22390_), .B(new_n22397_), .ZN(new_n22398_));
  NAND2_X1   g19352(.A1(new_n3232_), .A2(new_n16401_), .ZN(new_n22399_));
  AOI21_X1   g19353(.A1(new_n22398_), .A2(new_n22388_), .B(new_n22399_), .ZN(new_n22400_));
  NAND2_X1   g19354(.A1(new_n22287_), .A2(new_n22289_), .ZN(new_n22401_));
  NAND2_X1   g19355(.A1(new_n22401_), .A2(new_n16401_), .ZN(new_n22402_));
  OAI22_X1   g19356(.A1(new_n22400_), .A2(new_n22402_), .B1(new_n11572_), .B2(new_n3231_), .ZN(new_n22403_));
  OAI21_X1   g19357(.A1(new_n22403_), .A2(pi0625), .B(new_n22383_), .ZN(new_n22404_));
  NAND3_X1   g19358(.A1(new_n22403_), .A2(new_n12970_), .A3(new_n22291_), .ZN(new_n22405_));
  NAND4_X1   g19359(.A1(new_n22404_), .A2(new_n22405_), .A3(new_n12977_), .A4(new_n22336_), .ZN(new_n22406_));
  INV_X1     g19360(.I(new_n22335_), .ZN(new_n22407_));
  NOR4_X1    g19361(.A1(new_n22403_), .A2(new_n12970_), .A3(pi1153), .A4(new_n22383_), .ZN(new_n22408_));
  OAI21_X1   g19362(.A1(new_n22408_), .A2(new_n22407_), .B(new_n13657_), .ZN(new_n22409_));
  NAND2_X1   g19363(.A1(new_n22406_), .A2(new_n22409_), .ZN(new_n22410_));
  NOR2_X1    g19364(.A1(new_n22403_), .A2(pi0778), .ZN(new_n22411_));
  AOI21_X1   g19365(.A1(new_n22410_), .A2(pi0778), .B(new_n22411_), .ZN(new_n22412_));
  NOR2_X1    g19366(.A1(new_n22412_), .A2(pi0785), .ZN(new_n22413_));
  INV_X1     g19367(.I(new_n22339_), .ZN(new_n22414_));
  NAND3_X1   g19368(.A1(new_n22414_), .A2(pi0609), .A3(pi1155), .ZN(new_n22415_));
  NAND3_X1   g19369(.A1(new_n22415_), .A2(new_n11923_), .A3(new_n22298_), .ZN(new_n22416_));
  NOR4_X1    g19370(.A1(new_n22412_), .A2(new_n11903_), .A3(new_n22414_), .A4(pi1155), .ZN(new_n22417_));
  NAND2_X1   g19371(.A1(new_n22296_), .A2(pi0660), .ZN(new_n22418_));
  NOR2_X1    g19372(.A1(new_n22417_), .A2(new_n22418_), .ZN(new_n22419_));
  NOR2_X1    g19373(.A1(new_n22419_), .A2(new_n11870_), .ZN(new_n22420_));
  AOI21_X1   g19374(.A1(new_n22420_), .A2(new_n22416_), .B(new_n22413_), .ZN(new_n22421_));
  INV_X1     g19375(.I(new_n22341_), .ZN(new_n22422_));
  NOR4_X1    g19376(.A1(new_n22421_), .A2(new_n11934_), .A3(pi1154), .A4(new_n22422_), .ZN(new_n22423_));
  NAND2_X1   g19377(.A1(new_n22303_), .A2(pi0627), .ZN(new_n22424_));
  NOR3_X1    g19378(.A1(new_n22341_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n22425_));
  NAND2_X1   g19379(.A1(new_n22306_), .A2(new_n11949_), .ZN(new_n22426_));
  OAI22_X1   g19380(.A1(new_n22423_), .A2(new_n22424_), .B1(new_n22425_), .B2(new_n22426_), .ZN(new_n22427_));
  MUX2_X1    g19381(.I0(new_n22427_), .I1(new_n22421_), .S(new_n11969_), .Z(new_n22428_));
  XNOR2_X1   g19382(.A1(new_n22428_), .A2(new_n22342_), .ZN(new_n22429_));
  NOR2_X1    g19383(.A1(new_n22429_), .A2(new_n11967_), .ZN(new_n22430_));
  NAND3_X1   g19384(.A1(new_n22381_), .A2(new_n11869_), .A3(new_n22382_), .ZN(new_n22431_));
  XOR2_X1    g19385(.A1(new_n22430_), .A2(new_n22428_), .Z(new_n22432_));
  AOI21_X1   g19386(.A1(new_n22282_), .A2(new_n11967_), .B(pi1159), .ZN(new_n22433_));
  AOI21_X1   g19387(.A1(new_n22381_), .A2(new_n22433_), .B(pi0648), .ZN(new_n22434_));
  OAI21_X1   g19388(.A1(new_n22432_), .A2(pi1159), .B(new_n22434_), .ZN(new_n22435_));
  OR2_X2     g19389(.A1(new_n22428_), .A2(pi0789), .Z(new_n22436_));
  NAND3_X1   g19390(.A1(new_n22312_), .A2(pi0626), .A3(new_n22282_), .ZN(new_n22437_));
  OAI21_X1   g19391(.A1(new_n22312_), .A2(new_n11994_), .B(new_n22281_), .ZN(new_n22438_));
  AOI21_X1   g19392(.A1(new_n22438_), .A2(new_n22437_), .B(new_n17167_), .ZN(new_n22439_));
  AOI21_X1   g19393(.A1(new_n22312_), .A2(new_n22282_), .B(new_n11994_), .ZN(new_n22440_));
  NAND2_X1   g19394(.A1(new_n22440_), .A2(new_n11990_), .ZN(new_n22441_));
  NOR2_X1    g19395(.A1(new_n22343_), .A2(new_n12020_), .ZN(new_n22442_));
  NOR2_X1    g19396(.A1(new_n22442_), .A2(pi0788), .ZN(new_n22443_));
  NAND2_X1   g19397(.A1(new_n22441_), .A2(new_n22443_), .ZN(new_n22444_));
  OAI21_X1   g19398(.A1(new_n22444_), .A2(new_n22439_), .B(new_n17372_), .ZN(new_n22445_));
  AOI21_X1   g19399(.A1(new_n11998_), .A2(new_n22436_), .B(new_n22445_), .ZN(new_n22446_));
  NAND3_X1   g19400(.A1(new_n22435_), .A2(new_n22431_), .A3(new_n22446_), .ZN(new_n22447_));
  AOI21_X1   g19401(.A1(new_n22447_), .A2(new_n22380_), .B(new_n14725_), .ZN(new_n22448_));
  OAI21_X1   g19402(.A1(new_n22448_), .A2(new_n22375_), .B(new_n22371_), .ZN(new_n22449_));
  AOI21_X1   g19403(.A1(new_n22368_), .A2(new_n22449_), .B(po1038), .ZN(new_n22450_));
  OAI21_X1   g19404(.A1(new_n6845_), .A2(pi0192), .B(new_n13184_), .ZN(new_n22451_));
  OAI21_X1   g19405(.A1(new_n22450_), .A2(new_n22451_), .B(new_n22280_), .ZN(po0349));
  NOR2_X1    g19406(.A1(new_n2925_), .A2(pi0193), .ZN(new_n22453_));
  NOR2_X1    g19407(.A1(new_n11877_), .A2(new_n16415_), .ZN(new_n22454_));
  NOR2_X1    g19408(.A1(new_n22454_), .A2(new_n22453_), .ZN(new_n22455_));
  AOI21_X1   g19409(.A1(new_n11886_), .A2(pi0690), .B(new_n22453_), .ZN(new_n22456_));
  NOR2_X1    g19410(.A1(new_n22456_), .A2(new_n11874_), .ZN(new_n22457_));
  INV_X1     g19411(.I(new_n22457_), .ZN(new_n22458_));
  NAND2_X1   g19412(.A1(new_n22458_), .A2(new_n22455_), .ZN(new_n22459_));
  NAND2_X1   g19413(.A1(new_n22459_), .A2(new_n11891_), .ZN(new_n22460_));
  NOR2_X1    g19414(.A1(new_n22458_), .A2(new_n12970_), .ZN(new_n22461_));
  NOR4_X1    g19415(.A1(new_n22461_), .A2(new_n11893_), .A3(new_n22453_), .A4(new_n22454_), .ZN(new_n22462_));
  NOR2_X1    g19416(.A1(new_n13201_), .A2(new_n16448_), .ZN(new_n22463_));
  NOR2_X1    g19417(.A1(new_n22453_), .A2(pi1153), .ZN(new_n22464_));
  INV_X1     g19418(.I(new_n22464_), .ZN(new_n22465_));
  NOR2_X1    g19419(.A1(new_n22463_), .A2(new_n22465_), .ZN(new_n22466_));
  INV_X1     g19420(.I(new_n22466_), .ZN(new_n22467_));
  NAND2_X1   g19421(.A1(new_n22467_), .A2(pi0608), .ZN(new_n22468_));
  INV_X1     g19422(.I(new_n22461_), .ZN(new_n22469_));
  AOI21_X1   g19423(.A1(new_n22469_), .A2(new_n22459_), .B(new_n22465_), .ZN(new_n22470_));
  OAI21_X1   g19424(.A1(new_n22463_), .A2(new_n22456_), .B(pi1153), .ZN(new_n22471_));
  NAND2_X1   g19425(.A1(new_n22471_), .A2(new_n13657_), .ZN(new_n22472_));
  OAI22_X1   g19426(.A1(new_n22468_), .A2(new_n22462_), .B1(new_n22470_), .B2(new_n22472_), .ZN(new_n22473_));
  NAND2_X1   g19427(.A1(new_n22473_), .A2(pi0778), .ZN(new_n22474_));
  XOR2_X1    g19428(.A1(new_n22474_), .A2(new_n22460_), .Z(new_n22475_));
  INV_X1     g19429(.I(new_n22475_), .ZN(new_n22476_));
  NAND2_X1   g19430(.A1(new_n22467_), .A2(new_n22471_), .ZN(new_n22477_));
  MUX2_X1    g19431(.I0(new_n22477_), .I1(new_n22456_), .S(new_n11891_), .Z(new_n22478_));
  XNOR2_X1   g19432(.A1(new_n22475_), .A2(new_n22478_), .ZN(new_n22479_));
  NAND2_X1   g19433(.A1(new_n22479_), .A2(pi0609), .ZN(new_n22480_));
  XOR2_X1    g19434(.A1(new_n22480_), .A2(new_n22476_), .Z(new_n22481_));
  INV_X1     g19435(.I(new_n22454_), .ZN(new_n22482_));
  NOR2_X1    g19436(.A1(new_n22455_), .A2(new_n11925_), .ZN(new_n22483_));
  NOR4_X1    g19437(.A1(new_n22483_), .A2(pi1155), .A3(new_n12997_), .A4(new_n22482_), .ZN(new_n22484_));
  NOR2_X1    g19438(.A1(new_n22484_), .A2(pi0660), .ZN(new_n22485_));
  OAI21_X1   g19439(.A1(new_n22481_), .A2(pi1155), .B(new_n22485_), .ZN(new_n22486_));
  NOR2_X1    g19440(.A1(new_n22482_), .A2(new_n12997_), .ZN(new_n22487_));
  NOR4_X1    g19441(.A1(new_n22487_), .A2(new_n11923_), .A3(pi1155), .A4(new_n22453_), .ZN(new_n22489_));
  NOR2_X1    g19442(.A1(new_n22489_), .A2(new_n11870_), .ZN(new_n22490_));
  AOI22_X1   g19443(.A1(new_n22486_), .A2(new_n22490_), .B1(new_n11870_), .B2(new_n22476_), .ZN(new_n22491_));
  NOR2_X1    g19444(.A1(new_n22491_), .A2(pi0781), .ZN(new_n22492_));
  NOR4_X1    g19445(.A1(new_n22478_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n22493_));
  NOR2_X1    g19446(.A1(new_n22483_), .A2(pi0785), .ZN(new_n22494_));
  NOR4_X1    g19447(.A1(new_n22484_), .A2(pi1155), .A3(new_n22453_), .A4(new_n22487_), .ZN(new_n22495_));
  NOR2_X1    g19448(.A1(new_n22495_), .A2(new_n11870_), .ZN(new_n22496_));
  XOR2_X1    g19449(.A1(new_n22496_), .A2(new_n22494_), .Z(new_n22497_));
  INV_X1     g19450(.I(new_n22497_), .ZN(new_n22498_));
  OAI21_X1   g19451(.A1(new_n22498_), .A2(new_n11945_), .B(new_n11949_), .ZN(new_n22499_));
  OAI21_X1   g19452(.A1(new_n22498_), .A2(new_n11952_), .B(new_n11950_), .ZN(new_n22500_));
  NOR2_X1    g19453(.A1(new_n22478_), .A2(new_n11939_), .ZN(new_n22501_));
  NOR4_X1    g19454(.A1(new_n22491_), .A2(new_n11934_), .A3(pi1154), .A4(new_n22501_), .ZN(new_n22502_));
  NOR2_X1    g19455(.A1(new_n22502_), .A2(new_n22500_), .ZN(new_n22503_));
  OAI22_X1   g19456(.A1(new_n22503_), .A2(pi0627), .B1(new_n22493_), .B2(new_n22499_), .ZN(new_n22504_));
  AOI21_X1   g19457(.A1(new_n22504_), .A2(pi0781), .B(new_n22492_), .ZN(new_n22505_));
  INV_X1     g19458(.I(new_n22501_), .ZN(new_n22506_));
  NOR2_X1    g19459(.A1(new_n22506_), .A2(new_n11962_), .ZN(new_n22507_));
  NOR4_X1    g19460(.A1(new_n22505_), .A2(new_n11967_), .A3(pi1159), .A4(new_n22507_), .ZN(new_n22508_));
  NOR2_X1    g19461(.A1(new_n22498_), .A2(pi0781), .ZN(new_n22509_));
  AOI21_X1   g19462(.A1(new_n11944_), .A2(new_n22497_), .B(new_n22500_), .ZN(new_n22510_));
  NOR2_X1    g19463(.A1(new_n22510_), .A2(new_n11969_), .ZN(new_n22511_));
  XOR2_X1    g19464(.A1(new_n22511_), .A2(new_n22509_), .Z(new_n22512_));
  AOI21_X1   g19465(.A1(new_n22512_), .A2(new_n16479_), .B(pi1159), .ZN(new_n22513_));
  INV_X1     g19466(.I(new_n22513_), .ZN(new_n22514_));
  NOR3_X1    g19467(.A1(new_n22508_), .A2(new_n11966_), .A3(new_n22514_), .ZN(new_n22515_));
  NOR4_X1    g19468(.A1(new_n22506_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n22516_));
  INV_X1     g19469(.I(new_n22512_), .ZN(new_n22517_));
  NOR2_X1    g19470(.A1(new_n22517_), .A2(new_n16482_), .ZN(new_n22518_));
  NOR3_X1    g19471(.A1(new_n22518_), .A2(pi0648), .A3(new_n22516_), .ZN(new_n22519_));
  AOI21_X1   g19472(.A1(new_n22505_), .A2(new_n11998_), .B(pi0789), .ZN(new_n22520_));
  OAI21_X1   g19473(.A1(new_n22515_), .A2(new_n22519_), .B(new_n22520_), .ZN(new_n22521_));
  NAND2_X1   g19474(.A1(new_n22507_), .A2(new_n17450_), .ZN(new_n22522_));
  NOR2_X1    g19475(.A1(new_n22522_), .A2(new_n17153_), .ZN(new_n22523_));
  NOR2_X1    g19476(.A1(new_n14624_), .A2(new_n22453_), .ZN(new_n22524_));
  NOR2_X1    g19477(.A1(new_n22517_), .A2(pi0789), .ZN(new_n22525_));
  NOR2_X1    g19478(.A1(new_n22514_), .A2(new_n22518_), .ZN(new_n22526_));
  NOR2_X1    g19479(.A1(new_n22526_), .A2(new_n11985_), .ZN(new_n22527_));
  XOR2_X1    g19480(.A1(new_n22527_), .A2(new_n22525_), .Z(new_n22528_));
  AOI21_X1   g19481(.A1(new_n22528_), .A2(new_n14624_), .B(new_n22524_), .ZN(new_n22529_));
  AOI22_X1   g19482(.A1(new_n22529_), .A2(new_n12064_), .B1(new_n15080_), .B2(new_n22523_), .ZN(new_n22530_));
  NOR2_X1    g19483(.A1(new_n22530_), .A2(new_n12030_), .ZN(new_n22531_));
  NAND2_X1   g19484(.A1(new_n22529_), .A2(new_n12063_), .ZN(new_n22532_));
  AOI21_X1   g19485(.A1(new_n22523_), .A2(new_n15084_), .B(new_n15086_), .ZN(new_n22533_));
  NAND2_X1   g19486(.A1(new_n22532_), .A2(new_n22533_), .ZN(new_n22534_));
  OAI21_X1   g19487(.A1(new_n22531_), .A2(new_n22534_), .B(new_n14726_), .ZN(new_n22535_));
  INV_X1     g19488(.I(new_n22453_), .ZN(new_n22536_));
  MUX2_X1    g19489(.I0(new_n22528_), .I1(new_n22536_), .S(new_n11994_), .Z(new_n22537_));
  INV_X1     g19490(.I(new_n22528_), .ZN(new_n22538_));
  AOI21_X1   g19491(.A1(new_n22538_), .A2(new_n22536_), .B(new_n11994_), .ZN(new_n22539_));
  OAI21_X1   g19492(.A1(new_n22522_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n22540_));
  AOI21_X1   g19493(.A1(new_n22539_), .A2(new_n11990_), .B(new_n22540_), .ZN(new_n22541_));
  OAI21_X1   g19494(.A1(new_n17167_), .A2(new_n22537_), .B(new_n22541_), .ZN(new_n22542_));
  NAND4_X1   g19495(.A1(new_n22521_), .A2(new_n22535_), .A3(new_n22542_), .A4(new_n14732_), .ZN(new_n22543_));
  NAND3_X1   g19496(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n22453_), .ZN(new_n22544_));
  NAND2_X1   g19497(.A1(new_n22523_), .A2(new_n15050_), .ZN(new_n22545_));
  NAND2_X1   g19498(.A1(new_n22545_), .A2(pi0647), .ZN(new_n22546_));
  NAND2_X1   g19499(.A1(new_n22453_), .A2(pi0647), .ZN(new_n22547_));
  NAND3_X1   g19500(.A1(new_n22546_), .A2(new_n12049_), .A3(new_n22547_), .ZN(new_n22548_));
  NAND2_X1   g19501(.A1(new_n22548_), .A2(pi0630), .ZN(new_n22549_));
  NOR2_X1    g19502(.A1(new_n22545_), .A2(new_n12061_), .ZN(new_n22550_));
  AOI21_X1   g19503(.A1(new_n12061_), .A2(new_n22453_), .B(new_n22550_), .ZN(new_n22551_));
  NAND2_X1   g19504(.A1(new_n22551_), .A2(new_n12088_), .ZN(new_n22552_));
  NAND4_X1   g19505(.A1(new_n22552_), .A2(new_n22549_), .A3(pi0787), .A4(new_n22544_), .ZN(new_n22553_));
  AND2_X2    g19506(.A1(new_n22543_), .A2(new_n22553_), .Z(new_n22554_));
  NOR2_X1    g19507(.A1(new_n22554_), .A2(new_n12082_), .ZN(new_n22555_));
  NAND4_X1   g19508(.A1(new_n22546_), .A2(pi0787), .A3(new_n12049_), .A4(new_n22547_), .ZN(new_n22556_));
  OAI21_X1   g19509(.A1(pi0787), .A2(new_n22545_), .B(new_n22556_), .ZN(new_n22557_));
  NOR2_X1    g19510(.A1(new_n22557_), .A2(pi0644), .ZN(new_n22558_));
  OR3_X2     g19511(.A1(new_n22555_), .A2(pi0715), .A3(new_n22558_), .Z(new_n22559_));
  MUX2_X1    g19512(.I0(new_n22529_), .I1(new_n22453_), .S(new_n16841_), .Z(new_n22560_));
  INV_X1     g19513(.I(new_n22560_), .ZN(new_n22561_));
  OAI21_X1   g19514(.A1(new_n22560_), .A2(new_n22453_), .B(new_n12082_), .ZN(new_n22562_));
  AOI21_X1   g19515(.A1(new_n22453_), .A2(new_n22560_), .B(new_n22562_), .ZN(new_n22563_));
  OAI21_X1   g19516(.A1(new_n22563_), .A2(new_n22561_), .B(new_n12099_), .ZN(new_n22564_));
  AOI21_X1   g19517(.A1(new_n22561_), .A2(new_n22563_), .B(new_n22564_), .ZN(new_n22565_));
  AOI21_X1   g19518(.A1(new_n22559_), .A2(new_n22565_), .B(pi1160), .ZN(new_n22566_));
  XOR2_X1    g19519(.A1(new_n22563_), .A2(new_n22453_), .Z(new_n22567_));
  AOI21_X1   g19520(.A1(new_n22557_), .A2(pi0644), .B(new_n13169_), .ZN(new_n22568_));
  OAI21_X1   g19521(.A1(new_n22567_), .A2(new_n12099_), .B(new_n22568_), .ZN(new_n22569_));
  OAI21_X1   g19522(.A1(new_n22569_), .A2(new_n22555_), .B(pi0790), .ZN(new_n22570_));
  NOR2_X1    g19523(.A1(new_n22554_), .A2(new_n14748_), .ZN(new_n22571_));
  OAI21_X1   g19524(.A1(new_n22566_), .A2(new_n22570_), .B(new_n22571_), .ZN(new_n22572_));
  NOR2_X1    g19525(.A1(new_n12965_), .A2(pi0193), .ZN(new_n22573_));
  INV_X1     g19526(.I(new_n22573_), .ZN(new_n22574_));
  NAND2_X1   g19527(.A1(new_n22574_), .A2(new_n11997_), .ZN(new_n22575_));
  NOR3_X1    g19528(.A1(new_n15144_), .A2(pi0193), .A3(pi0739), .ZN(new_n22576_));
  INV_X1     g19529(.I(new_n22576_), .ZN(new_n22577_));
  MUX2_X1    g19530(.I0(new_n13381_), .I1(new_n14362_), .S(new_n7179_), .Z(new_n22578_));
  AOI21_X1   g19531(.A1(new_n22578_), .A2(new_n16415_), .B(pi0038), .ZN(new_n22579_));
  NOR2_X1    g19532(.A1(new_n12828_), .A2(pi0193), .ZN(new_n22580_));
  NOR2_X1    g19533(.A1(new_n13367_), .A2(new_n16415_), .ZN(new_n22581_));
  NOR3_X1    g19534(.A1(new_n22581_), .A2(new_n3172_), .A3(new_n22580_), .ZN(new_n22582_));
  AOI21_X1   g19535(.A1(new_n22579_), .A2(new_n22577_), .B(new_n22582_), .ZN(new_n22583_));
  NOR2_X1    g19536(.A1(new_n3231_), .A2(pi0193), .ZN(new_n22584_));
  AOI21_X1   g19537(.A1(new_n22583_), .A2(new_n3231_), .B(new_n22584_), .ZN(new_n22585_));
  NOR2_X1    g19538(.A1(new_n22585_), .A2(new_n11914_), .ZN(new_n22586_));
  OAI21_X1   g19539(.A1(new_n22574_), .A2(new_n11924_), .B(new_n11870_), .ZN(new_n22587_));
  NOR2_X1    g19540(.A1(new_n22586_), .A2(new_n22587_), .ZN(new_n22588_));
  NAND2_X1   g19541(.A1(new_n22585_), .A2(new_n11924_), .ZN(new_n22589_));
  OAI22_X1   g19542(.A1(new_n22589_), .A2(pi0609), .B1(new_n12996_), .B2(new_n22573_), .ZN(new_n22590_));
  NAND2_X1   g19543(.A1(new_n22590_), .A2(new_n11912_), .ZN(new_n22591_));
  OAI22_X1   g19544(.A1(new_n22589_), .A2(new_n11903_), .B1(new_n11915_), .B2(new_n22573_), .ZN(new_n22592_));
  NAND2_X1   g19545(.A1(new_n22592_), .A2(pi1155), .ZN(new_n22593_));
  AOI21_X1   g19546(.A1(new_n22591_), .A2(new_n22593_), .B(new_n11870_), .ZN(new_n22594_));
  XOR2_X1    g19547(.A1(new_n22594_), .A2(new_n22588_), .Z(new_n22595_));
  NAND3_X1   g19548(.A1(new_n22574_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n22596_));
  MUX2_X1    g19549(.I0(new_n22596_), .I1(new_n22595_), .S(new_n11969_), .Z(new_n22597_));
  NOR3_X1    g19550(.A1(new_n22573_), .A2(pi0619), .A3(pi1159), .ZN(new_n22598_));
  INV_X1     g19551(.I(new_n22598_), .ZN(new_n22599_));
  MUX2_X1    g19552(.I0(new_n22599_), .I1(new_n22597_), .S(new_n11985_), .Z(new_n22600_));
  NAND2_X1   g19553(.A1(new_n22600_), .A2(new_n14624_), .ZN(new_n22601_));
  AOI21_X1   g19554(.A1(new_n22601_), .A2(new_n22575_), .B(new_n12053_), .ZN(new_n22602_));
  NOR2_X1    g19555(.A1(new_n22573_), .A2(new_n12054_), .ZN(new_n22603_));
  OAI21_X1   g19556(.A1(new_n22602_), .A2(new_n22603_), .B(new_n12092_), .ZN(new_n22604_));
  NAND2_X1   g19557(.A1(new_n22574_), .A2(new_n12091_), .ZN(new_n22605_));
  NAND3_X1   g19558(.A1(new_n22604_), .A2(new_n12082_), .A3(new_n22605_), .ZN(new_n22606_));
  AOI21_X1   g19559(.A1(new_n22573_), .A2(pi0644), .B(new_n12099_), .ZN(new_n22607_));
  NAND2_X1   g19560(.A1(new_n22606_), .A2(new_n22607_), .ZN(new_n22608_));
  NOR2_X1    g19561(.A1(new_n22573_), .A2(new_n13114_), .ZN(new_n22609_));
  NOR2_X1    g19562(.A1(new_n22574_), .A2(new_n12014_), .ZN(new_n22610_));
  NOR2_X1    g19563(.A1(new_n22573_), .A2(new_n11961_), .ZN(new_n22611_));
  NOR2_X1    g19564(.A1(new_n13395_), .A2(new_n7179_), .ZN(new_n22612_));
  NOR2_X1    g19565(.A1(new_n22612_), .A2(pi0038), .ZN(new_n22613_));
  OAI22_X1   g19566(.A1(new_n22613_), .A2(new_n3232_), .B1(pi0193), .B2(new_n13399_), .ZN(new_n22614_));
  NOR3_X1    g19567(.A1(new_n15189_), .A2(pi0690), .A3(new_n22580_), .ZN(new_n22615_));
  NOR2_X1    g19568(.A1(new_n3232_), .A2(new_n16448_), .ZN(new_n22616_));
  AOI22_X1   g19569(.A1(new_n22574_), .A2(new_n22616_), .B1(new_n22614_), .B2(new_n22615_), .ZN(new_n22617_));
  NOR3_X1    g19570(.A1(new_n22574_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n22618_));
  NOR4_X1    g19571(.A1(new_n22617_), .A2(new_n12970_), .A3(pi1153), .A4(new_n22573_), .ZN(new_n22619_));
  NOR2_X1    g19572(.A1(new_n22619_), .A2(new_n22618_), .ZN(new_n22620_));
  MUX2_X1    g19573(.I0(new_n22620_), .I1(new_n22617_), .S(new_n11891_), .Z(new_n22621_));
  NOR2_X1    g19574(.A1(new_n22621_), .A2(new_n13024_), .ZN(new_n22622_));
  AOI21_X1   g19575(.A1(new_n13024_), .A2(new_n22573_), .B(new_n22622_), .ZN(new_n22623_));
  AOI21_X1   g19576(.A1(new_n22623_), .A2(new_n11961_), .B(new_n22611_), .ZN(new_n22624_));
  AOI21_X1   g19577(.A1(new_n22624_), .A2(new_n12014_), .B(new_n22610_), .ZN(new_n22625_));
  AOI21_X1   g19578(.A1(new_n22625_), .A2(new_n13114_), .B(new_n22609_), .ZN(new_n22626_));
  NOR3_X1    g19579(.A1(new_n22574_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n22627_));
  NOR4_X1    g19580(.A1(new_n22626_), .A2(new_n12031_), .A3(pi1156), .A4(new_n22573_), .ZN(new_n22628_));
  NOR2_X1    g19581(.A1(new_n22628_), .A2(new_n22627_), .ZN(new_n22629_));
  MUX2_X1    g19582(.I0(new_n22629_), .I1(new_n22626_), .S(new_n11868_), .Z(new_n22630_));
  NOR2_X1    g19583(.A1(new_n22630_), .A2(new_n12061_), .ZN(new_n22631_));
  AOI21_X1   g19584(.A1(new_n12061_), .A2(new_n22573_), .B(new_n22631_), .ZN(new_n22632_));
  NAND2_X1   g19585(.A1(new_n22632_), .A2(pi1157), .ZN(new_n22633_));
  NOR2_X1    g19586(.A1(new_n22630_), .A2(pi0647), .ZN(new_n22634_));
  AOI21_X1   g19587(.A1(pi0647), .A2(new_n22573_), .B(new_n22634_), .ZN(new_n22635_));
  NAND2_X1   g19588(.A1(new_n22635_), .A2(new_n12049_), .ZN(new_n22636_));
  AOI21_X1   g19589(.A1(new_n22636_), .A2(new_n22633_), .B(new_n12048_), .ZN(new_n22637_));
  AOI21_X1   g19590(.A1(new_n12048_), .A2(new_n22630_), .B(new_n22637_), .ZN(new_n22638_));
  NAND2_X1   g19591(.A1(new_n22638_), .A2(pi0644), .ZN(new_n22639_));
  AOI22_X1   g19592(.A1(new_n22639_), .A2(new_n12099_), .B1(new_n12081_), .B2(new_n22608_), .ZN(new_n22640_));
  NOR3_X1    g19593(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n22641_));
  NAND3_X1   g19594(.A1(new_n22604_), .A2(new_n22605_), .A3(new_n22641_), .ZN(new_n22642_));
  NAND2_X1   g19595(.A1(new_n22642_), .A2(pi0715), .ZN(new_n22643_));
  AOI21_X1   g19596(.A1(new_n22638_), .A2(new_n12082_), .B(new_n22643_), .ZN(new_n22644_));
  OAI21_X1   g19597(.A1(new_n22640_), .A2(new_n22644_), .B(pi0790), .ZN(new_n22645_));
  NAND2_X1   g19598(.A1(new_n22597_), .A2(pi0619), .ZN(new_n22646_));
  NAND2_X1   g19599(.A1(new_n22573_), .A2(pi0619), .ZN(new_n22647_));
  NAND2_X1   g19600(.A1(new_n17309_), .A2(new_n16415_), .ZN(new_n22648_));
  AOI21_X1   g19601(.A1(new_n12122_), .A2(new_n22648_), .B(pi0039), .ZN(new_n22649_));
  OR2_X2     g19602(.A1(new_n22649_), .A2(pi0193), .Z(new_n22650_));
  AOI21_X1   g19603(.A1(new_n13644_), .A2(new_n22482_), .B(new_n7179_), .ZN(new_n22651_));
  AOI21_X1   g19604(.A1(new_n22651_), .A2(new_n5156_), .B(new_n3172_), .ZN(new_n22652_));
  AOI21_X1   g19605(.A1(new_n13337_), .A2(pi0193), .B(pi0739), .ZN(new_n22653_));
  OAI21_X1   g19606(.A1(new_n13333_), .A2(new_n7179_), .B(new_n22653_), .ZN(new_n22654_));
  NOR3_X1    g19607(.A1(new_n12633_), .A2(new_n7179_), .A3(new_n12616_), .ZN(new_n22655_));
  AOI21_X1   g19608(.A1(new_n12633_), .A2(pi0193), .B(new_n13362_), .ZN(new_n22656_));
  OAI21_X1   g19609(.A1(new_n22655_), .A2(new_n22656_), .B(new_n16415_), .ZN(new_n22657_));
  INV_X1     g19610(.I(new_n22657_), .ZN(new_n22658_));
  OAI21_X1   g19611(.A1(new_n12668_), .A2(new_n7179_), .B(new_n16415_), .ZN(new_n22659_));
  AOI21_X1   g19612(.A1(new_n7179_), .A2(new_n12665_), .B(new_n22659_), .ZN(new_n22660_));
  NOR4_X1    g19613(.A1(new_n22658_), .A2(pi0038), .A3(pi0039), .A4(new_n22660_), .ZN(new_n22661_));
  AOI22_X1   g19614(.A1(new_n22661_), .A2(new_n22654_), .B1(new_n22650_), .B2(new_n22652_), .ZN(new_n22662_));
  NOR4_X1    g19615(.A1(new_n22662_), .A2(pi0690), .A3(new_n3231_), .A4(new_n22583_), .ZN(new_n22663_));
  AOI21_X1   g19616(.A1(pi0193), .A2(new_n3232_), .B(new_n22663_), .ZN(new_n22664_));
  NAND2_X1   g19617(.A1(new_n22664_), .A2(pi0625), .ZN(new_n22665_));
  OAI21_X1   g19618(.A1(new_n22585_), .A2(new_n12970_), .B(new_n12977_), .ZN(new_n22666_));
  NOR2_X1    g19619(.A1(new_n22619_), .A2(new_n22666_), .ZN(new_n22667_));
  INV_X1     g19620(.I(new_n22618_), .ZN(new_n22668_));
  AOI21_X1   g19621(.A1(new_n22585_), .A2(new_n12970_), .B(pi1153), .ZN(new_n22669_));
  NAND2_X1   g19622(.A1(new_n22665_), .A2(new_n22669_), .ZN(new_n22670_));
  NAND2_X1   g19623(.A1(new_n22670_), .A2(new_n22668_), .ZN(new_n22671_));
  AOI22_X1   g19624(.A1(new_n22671_), .A2(new_n13657_), .B1(new_n22665_), .B2(new_n22667_), .ZN(new_n22672_));
  NOR2_X1    g19625(.A1(new_n22672_), .A2(new_n11891_), .ZN(new_n22673_));
  AOI21_X1   g19626(.A1(new_n11891_), .A2(new_n22664_), .B(new_n22673_), .ZN(new_n22674_));
  NOR2_X1    g19627(.A1(new_n22674_), .A2(pi0785), .ZN(new_n22675_));
  INV_X1     g19628(.I(new_n22621_), .ZN(new_n22676_));
  NAND3_X1   g19629(.A1(new_n22676_), .A2(pi0609), .A3(pi1155), .ZN(new_n22677_));
  NAND3_X1   g19630(.A1(new_n22677_), .A2(new_n11923_), .A3(new_n22593_), .ZN(new_n22678_));
  NOR4_X1    g19631(.A1(new_n22674_), .A2(new_n11903_), .A3(pi1155), .A4(new_n22676_), .ZN(new_n22679_));
  NAND2_X1   g19632(.A1(new_n22591_), .A2(pi0660), .ZN(new_n22680_));
  NOR2_X1    g19633(.A1(new_n22679_), .A2(new_n22680_), .ZN(new_n22681_));
  NOR2_X1    g19634(.A1(new_n22681_), .A2(new_n11870_), .ZN(new_n22682_));
  AOI21_X1   g19635(.A1(new_n22682_), .A2(new_n22678_), .B(new_n22675_), .ZN(new_n22683_));
  INV_X1     g19636(.I(new_n22623_), .ZN(new_n22684_));
  NOR4_X1    g19637(.A1(new_n22683_), .A2(new_n11934_), .A3(pi1154), .A4(new_n22684_), .ZN(new_n22685_));
  NAND2_X1   g19638(.A1(new_n22595_), .A2(pi0618), .ZN(new_n22686_));
  NAND2_X1   g19639(.A1(new_n22573_), .A2(pi0618), .ZN(new_n22687_));
  NAND4_X1   g19640(.A1(new_n22686_), .A2(pi0627), .A3(new_n11950_), .A4(new_n22687_), .ZN(new_n22688_));
  NOR3_X1    g19641(.A1(new_n22623_), .A2(new_n11934_), .A3(new_n11950_), .ZN(new_n22689_));
  AOI21_X1   g19642(.A1(new_n22574_), .A2(new_n11934_), .B(pi1154), .ZN(new_n22690_));
  NAND2_X1   g19643(.A1(new_n22686_), .A2(new_n22690_), .ZN(new_n22691_));
  NAND2_X1   g19644(.A1(new_n22691_), .A2(new_n11949_), .ZN(new_n22692_));
  OAI22_X1   g19645(.A1(new_n22685_), .A2(new_n22688_), .B1(new_n22689_), .B2(new_n22692_), .ZN(new_n22693_));
  MUX2_X1    g19646(.I0(new_n22693_), .I1(new_n22683_), .S(new_n11969_), .Z(new_n22694_));
  XNOR2_X1   g19647(.A1(new_n22694_), .A2(new_n22624_), .ZN(new_n22695_));
  NOR2_X1    g19648(.A1(new_n22695_), .A2(new_n11967_), .ZN(new_n22696_));
  NAND3_X1   g19649(.A1(new_n22646_), .A2(new_n11869_), .A3(new_n22647_), .ZN(new_n22697_));
  XNOR2_X1   g19650(.A1(new_n22696_), .A2(new_n22694_), .ZN(new_n22698_));
  NAND2_X1   g19651(.A1(new_n22698_), .A2(new_n11869_), .ZN(new_n22699_));
  AOI21_X1   g19652(.A1(new_n22574_), .A2(new_n11967_), .B(pi1159), .ZN(new_n22700_));
  AOI21_X1   g19653(.A1(new_n22646_), .A2(new_n22700_), .B(pi0648), .ZN(new_n22701_));
  NOR3_X1    g19654(.A1(new_n22600_), .A2(new_n11994_), .A3(new_n22573_), .ZN(new_n22702_));
  AOI21_X1   g19655(.A1(new_n22600_), .A2(pi0626), .B(new_n22574_), .ZN(new_n22703_));
  OAI21_X1   g19656(.A1(new_n22702_), .A2(new_n22703_), .B(new_n11988_), .ZN(new_n22704_));
  NAND2_X1   g19657(.A1(new_n22600_), .A2(pi0626), .ZN(new_n22705_));
  OAI21_X1   g19658(.A1(new_n11994_), .A2(new_n22574_), .B(new_n22705_), .ZN(new_n22706_));
  OAI21_X1   g19659(.A1(new_n22625_), .A2(new_n12020_), .B(new_n11986_), .ZN(new_n22707_));
  AOI21_X1   g19660(.A1(new_n22706_), .A2(new_n11990_), .B(new_n22707_), .ZN(new_n22708_));
  NAND2_X1   g19661(.A1(new_n22708_), .A2(new_n22704_), .ZN(new_n22709_));
  OAI21_X1   g19662(.A1(new_n22694_), .A2(pi0789), .B(new_n11998_), .ZN(new_n22710_));
  NAND3_X1   g19663(.A1(new_n22710_), .A2(new_n17372_), .A3(new_n22709_), .ZN(new_n22711_));
  AOI21_X1   g19664(.A1(new_n22699_), .A2(new_n22701_), .B(new_n22711_), .ZN(new_n22712_));
  OR2_X2     g19665(.A1(new_n22627_), .A2(new_n12030_), .Z(new_n22713_));
  OAI21_X1   g19666(.A1(new_n22628_), .A2(pi0629), .B(new_n22713_), .ZN(new_n22714_));
  NAND2_X1   g19667(.A1(new_n22601_), .A2(new_n22575_), .ZN(new_n22715_));
  NAND2_X1   g19668(.A1(new_n22715_), .A2(new_n15222_), .ZN(new_n22716_));
  NAND2_X1   g19669(.A1(new_n22716_), .A2(new_n22714_), .ZN(new_n22717_));
  AOI22_X1   g19670(.A1(new_n22712_), .A2(new_n22697_), .B1(pi0792), .B2(new_n22717_), .ZN(new_n22718_));
  NAND2_X1   g19671(.A1(new_n22632_), .A2(new_n12060_), .ZN(new_n22719_));
  AOI21_X1   g19672(.A1(new_n22635_), .A2(pi0630), .B(new_n15214_), .ZN(new_n22720_));
  NAND2_X1   g19673(.A1(new_n22720_), .A2(new_n22719_), .ZN(new_n22721_));
  NOR2_X1    g19674(.A1(new_n22602_), .A2(new_n22603_), .ZN(new_n22722_));
  NOR2_X1    g19675(.A1(new_n22722_), .A2(new_n15183_), .ZN(new_n22723_));
  NAND3_X1   g19676(.A1(new_n22608_), .A2(new_n12082_), .A3(new_n12081_), .ZN(new_n22724_));
  AOI21_X1   g19677(.A1(new_n22642_), .A2(pi0644), .B(pi0790), .ZN(new_n22725_));
  AOI22_X1   g19678(.A1(new_n22721_), .A2(new_n22723_), .B1(new_n22724_), .B2(new_n22725_), .ZN(new_n22726_));
  OAI21_X1   g19679(.A1(new_n22718_), .A2(new_n14725_), .B(new_n22726_), .ZN(new_n22727_));
  AOI21_X1   g19680(.A1(new_n22727_), .A2(new_n22645_), .B(po1038), .ZN(new_n22728_));
  OAI21_X1   g19681(.A1(new_n6845_), .A2(pi0193), .B(new_n13184_), .ZN(new_n22729_));
  OAI21_X1   g19682(.A1(new_n22728_), .A2(new_n22729_), .B(new_n22572_), .ZN(po0350));
  NOR2_X1    g19683(.A1(new_n2925_), .A2(pi0194), .ZN(new_n22731_));
  NOR2_X1    g19684(.A1(new_n11877_), .A2(new_n16315_), .ZN(new_n22732_));
  NOR2_X1    g19685(.A1(new_n22732_), .A2(new_n22731_), .ZN(new_n22733_));
  INV_X1     g19686(.I(new_n22733_), .ZN(new_n22734_));
  AOI21_X1   g19687(.A1(new_n11886_), .A2(pi0730), .B(new_n22731_), .ZN(new_n22735_));
  NOR2_X1    g19688(.A1(new_n22735_), .A2(new_n11874_), .ZN(new_n22736_));
  NOR2_X1    g19689(.A1(new_n22734_), .A2(new_n22736_), .ZN(new_n22737_));
  NOR2_X1    g19690(.A1(new_n22737_), .A2(pi0778), .ZN(new_n22738_));
  NAND2_X1   g19691(.A1(new_n22736_), .A2(pi0625), .ZN(new_n22739_));
  NOR2_X1    g19692(.A1(new_n13201_), .A2(new_n16318_), .ZN(new_n22740_));
  NOR4_X1    g19693(.A1(new_n22732_), .A2(pi0608), .A3(new_n11893_), .A4(new_n22731_), .ZN(new_n22741_));
  OAI21_X1   g19694(.A1(new_n22734_), .A2(new_n22736_), .B(new_n22739_), .ZN(new_n22742_));
  NOR3_X1    g19695(.A1(new_n22731_), .A2(pi0608), .A3(pi1153), .ZN(new_n22743_));
  AOI22_X1   g19696(.A1(new_n22742_), .A2(new_n22743_), .B1(new_n22739_), .B2(new_n22741_), .ZN(new_n22744_));
  NOR2_X1    g19697(.A1(new_n22744_), .A2(new_n11891_), .ZN(new_n22745_));
  XOR2_X1    g19698(.A1(new_n22745_), .A2(new_n22738_), .Z(new_n22746_));
  INV_X1     g19699(.I(new_n22746_), .ZN(new_n22747_));
  NAND2_X1   g19700(.A1(new_n22747_), .A2(new_n11870_), .ZN(new_n22748_));
  AOI21_X1   g19701(.A1(new_n22746_), .A2(new_n11903_), .B(pi1155), .ZN(new_n22749_));
  INV_X1     g19702(.I(new_n22735_), .ZN(new_n22750_));
  XOR2_X1    g19703(.A1(new_n22740_), .A2(pi1153), .Z(new_n22751_));
  NAND2_X1   g19704(.A1(new_n22751_), .A2(new_n22750_), .ZN(new_n22752_));
  OAI21_X1   g19705(.A1(new_n22740_), .A2(new_n22731_), .B(new_n11893_), .ZN(new_n22753_));
  AOI21_X1   g19706(.A1(new_n22752_), .A2(new_n22753_), .B(new_n11891_), .ZN(new_n22754_));
  NOR2_X1    g19707(.A1(new_n22735_), .A2(pi0778), .ZN(new_n22755_));
  OAI21_X1   g19708(.A1(new_n22754_), .A2(new_n22755_), .B(pi0609), .ZN(new_n22756_));
  AOI21_X1   g19709(.A1(new_n22734_), .A2(new_n11917_), .B(new_n11912_), .ZN(new_n22757_));
  NOR2_X1    g19710(.A1(new_n22757_), .A2(pi0660), .ZN(new_n22758_));
  OAI21_X1   g19711(.A1(new_n22749_), .A2(new_n22756_), .B(new_n22758_), .ZN(new_n22759_));
  NOR2_X1    g19712(.A1(new_n22754_), .A2(new_n22755_), .ZN(new_n22760_));
  NAND4_X1   g19713(.A1(new_n22747_), .A2(pi0609), .A3(new_n11912_), .A4(new_n22760_), .ZN(new_n22761_));
  NOR2_X1    g19714(.A1(new_n22733_), .A2(new_n11925_), .ZN(new_n22762_));
  AOI21_X1   g19715(.A1(new_n22762_), .A2(new_n11928_), .B(pi1155), .ZN(new_n22763_));
  NOR2_X1    g19716(.A1(new_n22763_), .A2(new_n11923_), .ZN(new_n22764_));
  NAND2_X1   g19717(.A1(new_n22761_), .A2(new_n22764_), .ZN(new_n22765_));
  NAND3_X1   g19718(.A1(new_n22765_), .A2(pi0785), .A3(new_n22759_), .ZN(new_n22766_));
  NAND2_X1   g19719(.A1(new_n22766_), .A2(new_n22748_), .ZN(new_n22767_));
  NOR4_X1    g19720(.A1(new_n22760_), .A2(new_n11934_), .A3(new_n11950_), .A4(new_n11939_), .ZN(new_n22769_));
  NOR2_X1    g19721(.A1(new_n22762_), .A2(pi0785), .ZN(new_n22770_));
  OAI21_X1   g19722(.A1(new_n22763_), .A2(new_n22757_), .B(pi0785), .ZN(new_n22771_));
  XNOR2_X1   g19723(.A1(new_n22771_), .A2(new_n22770_), .ZN(new_n22772_));
  INV_X1     g19724(.I(new_n22772_), .ZN(new_n22773_));
  NOR2_X1    g19725(.A1(new_n22773_), .A2(new_n11945_), .ZN(new_n22774_));
  NOR3_X1    g19726(.A1(new_n22769_), .A2(new_n22774_), .A3(pi0627), .ZN(new_n22775_));
  AOI21_X1   g19727(.A1(new_n22772_), .A2(new_n11951_), .B(pi1154), .ZN(new_n22776_));
  NOR2_X1    g19728(.A1(new_n22760_), .A2(new_n11939_), .ZN(new_n22777_));
  INV_X1     g19729(.I(new_n22777_), .ZN(new_n22778_));
  NAND4_X1   g19730(.A1(new_n22767_), .A2(pi0618), .A3(new_n11950_), .A4(new_n22778_), .ZN(new_n22779_));
  NAND2_X1   g19731(.A1(new_n22779_), .A2(new_n22776_), .ZN(new_n22780_));
  AOI21_X1   g19732(.A1(new_n22780_), .A2(new_n11949_), .B(new_n22775_), .ZN(new_n22781_));
  NOR2_X1    g19733(.A1(new_n22781_), .A2(new_n11969_), .ZN(new_n22782_));
  AOI21_X1   g19734(.A1(new_n11969_), .A2(new_n22767_), .B(new_n22782_), .ZN(new_n22783_));
  NOR2_X1    g19735(.A1(new_n22778_), .A2(new_n11962_), .ZN(new_n22784_));
  NOR4_X1    g19736(.A1(new_n22783_), .A2(new_n11967_), .A3(pi1159), .A4(new_n22784_), .ZN(new_n22785_));
  INV_X1     g19737(.I(new_n22774_), .ZN(new_n22786_));
  NAND2_X1   g19738(.A1(new_n22786_), .A2(new_n22776_), .ZN(new_n22787_));
  MUX2_X1    g19739(.I0(new_n22787_), .I1(new_n22772_), .S(new_n11969_), .Z(new_n22788_));
  NAND2_X1   g19740(.A1(new_n22788_), .A2(pi0619), .ZN(new_n22789_));
  INV_X1     g19741(.I(new_n22789_), .ZN(new_n22790_));
  INV_X1     g19742(.I(new_n22731_), .ZN(new_n22791_));
  OAI21_X1   g19743(.A1(new_n22791_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n22792_));
  NOR4_X1    g19744(.A1(new_n22785_), .A2(new_n11966_), .A3(new_n22790_), .A4(new_n22792_), .ZN(new_n22793_));
  NOR4_X1    g19745(.A1(new_n22778_), .A2(new_n11967_), .A3(new_n11869_), .A4(new_n11962_), .ZN(new_n22794_));
  OAI21_X1   g19746(.A1(new_n22731_), .A2(pi0619), .B(new_n11869_), .ZN(new_n22795_));
  OAI21_X1   g19747(.A1(new_n22790_), .A2(new_n22795_), .B(new_n11966_), .ZN(new_n22796_));
  NOR2_X1    g19748(.A1(new_n22796_), .A2(new_n22794_), .ZN(new_n22797_));
  AOI21_X1   g19749(.A1(new_n22783_), .A2(new_n11998_), .B(pi0789), .ZN(new_n22798_));
  OAI21_X1   g19750(.A1(new_n22793_), .A2(new_n22797_), .B(new_n22798_), .ZN(new_n22799_));
  NAND2_X1   g19751(.A1(new_n22784_), .A2(new_n17450_), .ZN(new_n22800_));
  NOR2_X1    g19752(.A1(new_n22800_), .A2(new_n17153_), .ZN(new_n22801_));
  INV_X1     g19753(.I(new_n22801_), .ZN(new_n22802_));
  NOR2_X1    g19754(.A1(new_n22802_), .A2(new_n17151_), .ZN(new_n22803_));
  NOR2_X1    g19755(.A1(new_n14624_), .A2(new_n22731_), .ZN(new_n22804_));
  NAND3_X1   g19756(.A1(new_n22791_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n22805_));
  MUX2_X1    g19757(.I0(new_n22805_), .I1(new_n22788_), .S(new_n11985_), .Z(new_n22806_));
  AOI21_X1   g19758(.A1(new_n22806_), .A2(new_n14624_), .B(new_n22804_), .ZN(new_n22807_));
  AND2_X2    g19759(.A1(new_n22807_), .A2(new_n12064_), .Z(new_n22808_));
  OAI21_X1   g19760(.A1(new_n22808_), .A2(new_n22803_), .B(pi0629), .ZN(new_n22809_));
  NAND2_X1   g19761(.A1(new_n22807_), .A2(new_n12063_), .ZN(new_n22810_));
  NAND2_X1   g19762(.A1(new_n22801_), .A2(new_n15084_), .ZN(new_n22811_));
  NAND4_X1   g19763(.A1(new_n22809_), .A2(new_n15085_), .A3(new_n22810_), .A4(new_n22811_), .ZN(new_n22812_));
  MUX2_X1    g19764(.I0(new_n22806_), .I1(new_n22791_), .S(new_n11994_), .Z(new_n22813_));
  NOR2_X1    g19765(.A1(new_n22813_), .A2(new_n17167_), .ZN(new_n22814_));
  OAI21_X1   g19766(.A1(new_n22806_), .A2(new_n22731_), .B(pi0626), .ZN(new_n22815_));
  NOR2_X1    g19767(.A1(new_n22800_), .A2(new_n12020_), .ZN(new_n22816_));
  NOR2_X1    g19768(.A1(new_n22816_), .A2(pi0788), .ZN(new_n22817_));
  OAI21_X1   g19769(.A1(new_n22815_), .A2(new_n17171_), .B(new_n22817_), .ZN(new_n22818_));
  OAI21_X1   g19770(.A1(new_n22814_), .A2(new_n22818_), .B(new_n14732_), .ZN(new_n22819_));
  AOI21_X1   g19771(.A1(new_n22812_), .A2(new_n14726_), .B(new_n22819_), .ZN(new_n22820_));
  NAND3_X1   g19772(.A1(new_n15077_), .A2(new_n12053_), .A3(new_n22731_), .ZN(new_n22821_));
  NOR2_X1    g19773(.A1(new_n22802_), .A2(new_n12068_), .ZN(new_n22822_));
  INV_X1     g19774(.I(new_n22822_), .ZN(new_n22823_));
  NAND2_X1   g19775(.A1(new_n22823_), .A2(pi0647), .ZN(new_n22824_));
  NAND2_X1   g19776(.A1(new_n22731_), .A2(pi0647), .ZN(new_n22825_));
  NAND3_X1   g19777(.A1(new_n22824_), .A2(new_n12049_), .A3(new_n22825_), .ZN(new_n22826_));
  NOR2_X1    g19778(.A1(new_n22791_), .A2(pi0647), .ZN(new_n22827_));
  AOI21_X1   g19779(.A1(new_n22822_), .A2(pi0647), .B(new_n22827_), .ZN(new_n22828_));
  NAND2_X1   g19780(.A1(new_n22828_), .A2(new_n12088_), .ZN(new_n22829_));
  NAND2_X1   g19781(.A1(new_n22829_), .A2(pi0787), .ZN(new_n22830_));
  AOI21_X1   g19782(.A1(pi0630), .A2(new_n22826_), .B(new_n22830_), .ZN(new_n22831_));
  AOI22_X1   g19783(.A1(new_n22799_), .A2(new_n22820_), .B1(new_n22821_), .B2(new_n22831_), .ZN(new_n22832_));
  NOR2_X1    g19784(.A1(new_n22832_), .A2(new_n12082_), .ZN(new_n22833_));
  NAND4_X1   g19785(.A1(new_n22824_), .A2(pi0787), .A3(new_n12049_), .A4(new_n22825_), .ZN(new_n22834_));
  OAI21_X1   g19786(.A1(pi0787), .A2(new_n22823_), .B(new_n22834_), .ZN(new_n22835_));
  NOR2_X1    g19787(.A1(new_n22835_), .A2(pi0644), .ZN(new_n22836_));
  OR3_X2     g19788(.A1(new_n22833_), .A2(pi0715), .A3(new_n22836_), .Z(new_n22837_));
  MUX2_X1    g19789(.I0(new_n22807_), .I1(new_n22731_), .S(new_n16841_), .Z(new_n22838_));
  INV_X1     g19790(.I(new_n22838_), .ZN(new_n22839_));
  OAI21_X1   g19791(.A1(new_n22838_), .A2(new_n22731_), .B(new_n12082_), .ZN(new_n22840_));
  AOI21_X1   g19792(.A1(new_n22731_), .A2(new_n22838_), .B(new_n22840_), .ZN(new_n22841_));
  OAI21_X1   g19793(.A1(new_n22841_), .A2(new_n22839_), .B(new_n12099_), .ZN(new_n22842_));
  AOI21_X1   g19794(.A1(new_n22839_), .A2(new_n22841_), .B(new_n22842_), .ZN(new_n22843_));
  AOI21_X1   g19795(.A1(new_n22837_), .A2(new_n22843_), .B(pi1160), .ZN(new_n22844_));
  XOR2_X1    g19796(.A1(new_n22841_), .A2(new_n22731_), .Z(new_n22845_));
  AOI21_X1   g19797(.A1(new_n22835_), .A2(pi0644), .B(new_n13169_), .ZN(new_n22846_));
  OAI21_X1   g19798(.A1(new_n22845_), .A2(new_n12099_), .B(new_n22846_), .ZN(new_n22847_));
  OAI21_X1   g19799(.A1(new_n22833_), .A2(new_n22847_), .B(pi0790), .ZN(new_n22848_));
  NOR2_X1    g19800(.A1(new_n22832_), .A2(new_n14748_), .ZN(new_n22849_));
  OAI21_X1   g19801(.A1(new_n22844_), .A2(new_n22848_), .B(new_n22849_), .ZN(new_n22850_));
  AOI21_X1   g19802(.A1(new_n17788_), .A2(new_n3172_), .B(new_n14340_), .ZN(new_n22851_));
  NOR2_X1    g19803(.A1(pi0194), .A2(pi0748), .ZN(new_n22852_));
  INV_X1     g19804(.I(new_n22852_), .ZN(new_n22853_));
  NOR2_X1    g19805(.A1(new_n12900_), .A2(pi0194), .ZN(new_n22854_));
  INV_X1     g19806(.I(new_n22854_), .ZN(new_n22855_));
  NOR3_X1    g19807(.A1(new_n16210_), .A2(pi0748), .A3(new_n22855_), .ZN(new_n22856_));
  NAND2_X1   g19808(.A1(new_n17506_), .A2(pi0194), .ZN(new_n22857_));
  NAND2_X1   g19809(.A1(new_n20355_), .A2(new_n11628_), .ZN(new_n22858_));
  NAND3_X1   g19810(.A1(new_n22858_), .A2(pi0748), .A3(new_n22857_), .ZN(new_n22859_));
  NAND2_X1   g19811(.A1(new_n22859_), .A2(new_n16318_), .ZN(new_n22860_));
  OAI22_X1   g19812(.A1(new_n22860_), .A2(new_n22856_), .B1(new_n22851_), .B2(new_n22853_), .ZN(new_n22861_));
  MUX2_X1    g19813(.I0(new_n22861_), .I1(new_n11628_), .S(new_n3232_), .Z(new_n22862_));
  INV_X1     g19814(.I(new_n22862_), .ZN(new_n22863_));
  NAND2_X1   g19815(.A1(new_n22862_), .A2(pi0625), .ZN(new_n22864_));
  NOR2_X1    g19816(.A1(new_n3231_), .A2(pi0194), .ZN(new_n22865_));
  INV_X1     g19817(.I(new_n22865_), .ZN(new_n22866_));
  NOR2_X1    g19818(.A1(new_n16210_), .A2(new_n22855_), .ZN(new_n22867_));
  NOR2_X1    g19819(.A1(new_n22867_), .A2(pi0748), .ZN(new_n22868_));
  AOI21_X1   g19820(.A1(new_n22858_), .A2(new_n22857_), .B(new_n16315_), .ZN(new_n22869_));
  NOR2_X1    g19821(.A1(new_n22868_), .A2(new_n22869_), .ZN(new_n22870_));
  OAI21_X1   g19822(.A1(new_n22870_), .A2(new_n3232_), .B(new_n22866_), .ZN(new_n22871_));
  INV_X1     g19823(.I(new_n22871_), .ZN(new_n22872_));
  AOI21_X1   g19824(.A1(new_n22872_), .A2(new_n12970_), .B(pi1153), .ZN(new_n22873_));
  NAND2_X1   g19825(.A1(new_n22864_), .A2(new_n22873_), .ZN(new_n22874_));
  NAND3_X1   g19826(.A1(new_n22867_), .A2(new_n16318_), .A3(new_n3231_), .ZN(new_n22875_));
  OAI21_X1   g19827(.A1(new_n11628_), .A2(new_n17547_), .B(new_n22875_), .ZN(new_n22876_));
  NOR2_X1    g19828(.A1(new_n22876_), .A2(new_n12970_), .ZN(new_n22877_));
  NOR2_X1    g19829(.A1(new_n12965_), .A2(pi0194), .ZN(new_n22878_));
  NAND2_X1   g19830(.A1(new_n22878_), .A2(pi0625), .ZN(new_n22879_));
  INV_X1     g19831(.I(new_n22879_), .ZN(new_n22880_));
  NOR4_X1    g19832(.A1(new_n22877_), .A2(new_n13657_), .A3(pi1153), .A4(new_n22880_), .ZN(new_n22881_));
  OAI21_X1   g19833(.A1(new_n22878_), .A2(pi0625), .B(new_n11893_), .ZN(new_n22882_));
  OAI21_X1   g19834(.A1(new_n22877_), .A2(new_n22882_), .B(new_n12977_), .ZN(new_n22883_));
  AOI21_X1   g19835(.A1(pi0625), .A2(new_n22871_), .B(new_n22883_), .ZN(new_n22884_));
  AOI22_X1   g19836(.A1(new_n22874_), .A2(new_n22881_), .B1(new_n22864_), .B2(new_n22884_), .ZN(new_n22885_));
  NOR3_X1    g19837(.A1(new_n22885_), .A2(new_n11891_), .A3(new_n22863_), .ZN(new_n22886_));
  AOI21_X1   g19838(.A1(new_n22885_), .A2(pi0778), .B(new_n22862_), .ZN(new_n22887_));
  NOR2_X1    g19839(.A1(new_n22886_), .A2(new_n22887_), .ZN(new_n22888_));
  NAND2_X1   g19840(.A1(new_n22888_), .A2(new_n11870_), .ZN(new_n22889_));
  NOR2_X1    g19841(.A1(new_n22876_), .A2(pi0778), .ZN(new_n22890_));
  NOR4_X1    g19842(.A1(new_n22877_), .A2(pi0625), .A3(pi1153), .A4(new_n22878_), .ZN(new_n22891_));
  NOR2_X1    g19843(.A1(new_n22891_), .A2(new_n11891_), .ZN(new_n22892_));
  XNOR2_X1   g19844(.A1(new_n22892_), .A2(new_n22890_), .ZN(new_n22893_));
  AOI21_X1   g19845(.A1(new_n22893_), .A2(new_n11903_), .B(new_n11912_), .ZN(new_n22894_));
  INV_X1     g19846(.I(new_n22878_), .ZN(new_n22895_));
  NOR2_X1    g19847(.A1(new_n22871_), .A2(new_n11914_), .ZN(new_n22896_));
  AOI22_X1   g19848(.A1(new_n22896_), .A2(new_n11903_), .B1(new_n12997_), .B2(new_n22895_), .ZN(new_n22897_));
  NOR2_X1    g19849(.A1(new_n22897_), .A2(pi1155), .ZN(new_n22898_));
  OAI21_X1   g19850(.A1(new_n22898_), .A2(new_n11923_), .B(pi0609), .ZN(new_n22899_));
  NOR2_X1    g19851(.A1(new_n22894_), .A2(new_n22899_), .ZN(new_n22900_));
  NOR3_X1    g19852(.A1(new_n22886_), .A2(new_n22887_), .A3(pi0609), .ZN(new_n22901_));
  NAND2_X1   g19853(.A1(new_n22893_), .A2(pi0609), .ZN(new_n22902_));
  NOR3_X1    g19854(.A1(new_n22871_), .A2(new_n11903_), .A3(new_n11914_), .ZN(new_n22903_));
  NOR2_X1    g19855(.A1(new_n11923_), .A2(pi1155), .ZN(new_n22904_));
  NAND2_X1   g19856(.A1(new_n22902_), .A2(new_n22904_), .ZN(new_n22905_));
  NOR2_X1    g19857(.A1(new_n22901_), .A2(new_n22905_), .ZN(new_n22906_));
  AOI21_X1   g19858(.A1(new_n22888_), .A2(new_n22900_), .B(new_n22906_), .ZN(new_n22907_));
  NOR3_X1    g19859(.A1(new_n22907_), .A2(new_n11870_), .A3(new_n22889_), .ZN(new_n22908_));
  INV_X1     g19860(.I(new_n22889_), .ZN(new_n22909_));
  INV_X1     g19861(.I(new_n22888_), .ZN(new_n22910_));
  INV_X1     g19862(.I(new_n22900_), .ZN(new_n22911_));
  OAI22_X1   g19863(.A1(new_n22911_), .A2(new_n22910_), .B1(new_n22901_), .B2(new_n22905_), .ZN(new_n22912_));
  AOI21_X1   g19864(.A1(new_n22912_), .A2(pi0785), .B(new_n22909_), .ZN(new_n22913_));
  NOR2_X1    g19865(.A1(new_n22908_), .A2(new_n22913_), .ZN(new_n22914_));
  NAND3_X1   g19866(.A1(new_n22912_), .A2(pi0785), .A3(new_n22909_), .ZN(new_n22915_));
  OAI21_X1   g19867(.A1(new_n22907_), .A2(new_n11870_), .B(new_n22889_), .ZN(new_n22916_));
  OAI21_X1   g19868(.A1(new_n22895_), .A2(new_n11924_), .B(new_n11870_), .ZN(new_n22917_));
  AOI21_X1   g19869(.A1(new_n22871_), .A2(new_n11924_), .B(new_n22917_), .ZN(new_n22918_));
  AOI21_X1   g19870(.A1(new_n13010_), .A2(new_n22895_), .B(new_n22903_), .ZN(new_n22919_));
  NOR2_X1    g19871(.A1(new_n22919_), .A2(new_n11912_), .ZN(new_n22920_));
  OAI21_X1   g19872(.A1(new_n22920_), .A2(new_n22898_), .B(pi0785), .ZN(new_n22921_));
  XOR2_X1    g19873(.A1(new_n22921_), .A2(new_n22918_), .Z(new_n22922_));
  NOR2_X1    g19874(.A1(new_n22922_), .A2(new_n11934_), .ZN(new_n22923_));
  NOR2_X1    g19875(.A1(new_n22895_), .A2(new_n11934_), .ZN(new_n22924_));
  NOR4_X1    g19876(.A1(new_n22923_), .A2(new_n11949_), .A3(pi1154), .A4(new_n22924_), .ZN(new_n22925_));
  NOR2_X1    g19877(.A1(new_n22895_), .A2(new_n11938_), .ZN(new_n22926_));
  AOI21_X1   g19878(.A1(new_n22893_), .A2(new_n11938_), .B(new_n22926_), .ZN(new_n22927_));
  NOR3_X1    g19879(.A1(new_n22925_), .A2(new_n11934_), .A3(pi1154), .ZN(new_n22928_));
  NAND3_X1   g19880(.A1(new_n22916_), .A2(new_n22915_), .A3(new_n22928_), .ZN(new_n22929_));
  NOR3_X1    g19881(.A1(new_n22908_), .A2(pi0618), .A3(new_n22913_), .ZN(new_n22930_));
  AOI21_X1   g19882(.A1(new_n22895_), .A2(new_n11934_), .B(pi1154), .ZN(new_n22931_));
  OAI21_X1   g19883(.A1(new_n22922_), .A2(new_n11934_), .B(new_n22931_), .ZN(new_n22932_));
  OAI21_X1   g19884(.A1(new_n22927_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n22933_));
  AOI21_X1   g19885(.A1(new_n22932_), .A2(new_n11949_), .B(new_n22933_), .ZN(new_n22934_));
  INV_X1     g19886(.I(new_n22934_), .ZN(new_n22935_));
  OAI21_X1   g19887(.A1(new_n22930_), .A2(new_n22935_), .B(new_n22929_), .ZN(new_n22936_));
  MUX2_X1    g19888(.I0(new_n22936_), .I1(new_n22914_), .S(new_n11969_), .Z(new_n22937_));
  NAND2_X1   g19889(.A1(new_n22937_), .A2(new_n11985_), .ZN(new_n22938_));
  INV_X1     g19890(.I(new_n22938_), .ZN(new_n22939_));
  NOR3_X1    g19891(.A1(new_n22908_), .A2(pi0781), .A3(new_n22913_), .ZN(new_n22940_));
  NAND3_X1   g19892(.A1(new_n22936_), .A2(new_n22940_), .A3(pi0781), .ZN(new_n22941_));
  INV_X1     g19893(.I(new_n22940_), .ZN(new_n22942_));
  NAND3_X1   g19894(.A1(new_n22916_), .A2(new_n22915_), .A3(new_n11934_), .ZN(new_n22943_));
  AOI22_X1   g19895(.A1(new_n22943_), .A2(new_n22934_), .B1(new_n22914_), .B2(new_n22928_), .ZN(new_n22944_));
  OAI21_X1   g19896(.A1(new_n22944_), .A2(new_n11969_), .B(new_n22942_), .ZN(new_n22945_));
  INV_X1     g19897(.I(new_n22922_), .ZN(new_n22946_));
  NOR3_X1    g19898(.A1(new_n22878_), .A2(pi0618), .A3(pi1154), .ZN(new_n22947_));
  INV_X1     g19899(.I(new_n22947_), .ZN(new_n22948_));
  MUX2_X1    g19900(.I0(new_n22948_), .I1(new_n22946_), .S(new_n11969_), .Z(new_n22949_));
  OAI21_X1   g19901(.A1(new_n22895_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n22950_));
  AOI21_X1   g19902(.A1(new_n22949_), .A2(pi0619), .B(new_n22950_), .ZN(new_n22951_));
  NOR2_X1    g19903(.A1(new_n22878_), .A2(new_n11961_), .ZN(new_n22952_));
  AOI21_X1   g19904(.A1(new_n22927_), .A2(new_n11961_), .B(new_n22952_), .ZN(new_n22953_));
  NAND2_X1   g19905(.A1(new_n11869_), .A2(pi0619), .ZN(new_n22954_));
  AOI21_X1   g19906(.A1(new_n22951_), .A2(pi0648), .B(new_n22954_), .ZN(new_n22955_));
  NAND3_X1   g19907(.A1(new_n22945_), .A2(new_n22941_), .A3(new_n22955_), .ZN(new_n22956_));
  NOR3_X1    g19908(.A1(new_n22944_), .A2(new_n11969_), .A3(new_n22942_), .ZN(new_n22957_));
  AOI21_X1   g19909(.A1(new_n22936_), .A2(pi0781), .B(new_n22940_), .ZN(new_n22958_));
  NOR3_X1    g19910(.A1(new_n22957_), .A2(new_n22958_), .A3(pi0619), .ZN(new_n22959_));
  NAND2_X1   g19911(.A1(new_n22949_), .A2(pi0619), .ZN(new_n22960_));
  AOI21_X1   g19912(.A1(new_n22895_), .A2(new_n11967_), .B(pi1159), .ZN(new_n22961_));
  NAND2_X1   g19913(.A1(new_n22960_), .A2(new_n22961_), .ZN(new_n22962_));
  NAND2_X1   g19914(.A1(new_n22962_), .A2(new_n11966_), .ZN(new_n22963_));
  AOI21_X1   g19915(.A1(new_n22953_), .A2(pi0619), .B(pi1159), .ZN(new_n22964_));
  NAND2_X1   g19916(.A1(new_n22963_), .A2(new_n22964_), .ZN(new_n22965_));
  OAI21_X1   g19917(.A1(new_n22959_), .A2(new_n22965_), .B(new_n22956_), .ZN(new_n22966_));
  NAND3_X1   g19918(.A1(new_n22966_), .A2(new_n22939_), .A3(pi0789), .ZN(new_n22967_));
  NAND3_X1   g19919(.A1(new_n22945_), .A2(new_n22941_), .A3(new_n11967_), .ZN(new_n22968_));
  INV_X1     g19920(.I(new_n22965_), .ZN(new_n22969_));
  AOI22_X1   g19921(.A1(new_n22968_), .A2(new_n22969_), .B1(new_n22937_), .B2(new_n22955_), .ZN(new_n22970_));
  OAI21_X1   g19922(.A1(new_n22970_), .A2(new_n11985_), .B(new_n22938_), .ZN(new_n22971_));
  NAND2_X1   g19923(.A1(new_n22971_), .A2(new_n22967_), .ZN(new_n22972_));
  NOR3_X1    g19924(.A1(new_n22970_), .A2(new_n11985_), .A3(new_n22938_), .ZN(new_n22973_));
  AOI21_X1   g19925(.A1(new_n22966_), .A2(pi0789), .B(new_n22939_), .ZN(new_n22974_));
  NOR3_X1    g19926(.A1(new_n22878_), .A2(pi0619), .A3(pi1159), .ZN(new_n22975_));
  INV_X1     g19927(.I(new_n22975_), .ZN(new_n22976_));
  MUX2_X1    g19928(.I0(new_n22976_), .I1(new_n22949_), .S(new_n11985_), .Z(new_n22977_));
  NOR3_X1    g19929(.A1(new_n11994_), .A2(new_n11989_), .A3(pi1158), .ZN(new_n22978_));
  NAND2_X1   g19930(.A1(new_n22977_), .A2(new_n22978_), .ZN(new_n22979_));
  NOR2_X1    g19931(.A1(new_n22895_), .A2(new_n12014_), .ZN(new_n22980_));
  AOI21_X1   g19932(.A1(new_n22953_), .A2(new_n12014_), .B(new_n22980_), .ZN(new_n22981_));
  NOR2_X1    g19933(.A1(new_n11994_), .A2(pi0641), .ZN(new_n22982_));
  NAND2_X1   g19934(.A1(new_n22979_), .A2(new_n22982_), .ZN(new_n22983_));
  INV_X1     g19935(.I(new_n22983_), .ZN(new_n22984_));
  NAND2_X1   g19936(.A1(new_n22977_), .A2(new_n11994_), .ZN(new_n22985_));
  AOI21_X1   g19937(.A1(new_n22895_), .A2(pi0626), .B(new_n11989_), .ZN(new_n22986_));
  NAND2_X1   g19938(.A1(new_n22985_), .A2(new_n22986_), .ZN(new_n22987_));
  NOR3_X1    g19939(.A1(new_n11989_), .A2(pi0626), .A3(pi1158), .ZN(new_n22988_));
  NAND2_X1   g19940(.A1(new_n22987_), .A2(new_n22988_), .ZN(new_n22989_));
  INV_X1     g19941(.I(new_n22989_), .ZN(new_n22990_));
  OAI22_X1   g19942(.A1(new_n22974_), .A2(new_n22973_), .B1(new_n22984_), .B2(new_n22990_), .ZN(new_n22991_));
  NOR3_X1    g19943(.A1(new_n22991_), .A2(new_n11986_), .A3(new_n22972_), .ZN(new_n22992_));
  NOR2_X1    g19944(.A1(new_n22974_), .A2(new_n22973_), .ZN(new_n22993_));
  AOI21_X1   g19945(.A1(new_n22991_), .A2(pi0788), .B(new_n22993_), .ZN(new_n22994_));
  NOR2_X1    g19946(.A1(new_n22992_), .A2(new_n22994_), .ZN(new_n22995_));
  NOR2_X1    g19947(.A1(new_n22878_), .A2(new_n14624_), .ZN(new_n22996_));
  AOI21_X1   g19948(.A1(new_n22977_), .A2(new_n14624_), .B(new_n22996_), .ZN(new_n22997_));
  NAND2_X1   g19949(.A1(new_n22997_), .A2(new_n12031_), .ZN(new_n22998_));
  NAND2_X1   g19950(.A1(new_n22998_), .A2(pi1156), .ZN(new_n22999_));
  NOR2_X1    g19951(.A1(new_n22878_), .A2(new_n13114_), .ZN(new_n23000_));
  AOI21_X1   g19952(.A1(new_n22981_), .A2(new_n13114_), .B(new_n23000_), .ZN(new_n23001_));
  NOR3_X1    g19953(.A1(new_n22895_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n23002_));
  NOR2_X1    g19954(.A1(new_n23002_), .A2(new_n12030_), .ZN(new_n23003_));
  NOR2_X1    g19955(.A1(new_n23003_), .A2(new_n12031_), .ZN(new_n23004_));
  NAND2_X1   g19956(.A1(new_n22999_), .A2(new_n23004_), .ZN(new_n23005_));
  INV_X1     g19957(.I(new_n23005_), .ZN(new_n23006_));
  NAND2_X1   g19958(.A1(new_n22997_), .A2(pi0628), .ZN(new_n23007_));
  INV_X1     g19959(.I(new_n23007_), .ZN(new_n23008_));
  NOR2_X1    g19960(.A1(new_n12030_), .A2(pi0628), .ZN(new_n23009_));
  OAI21_X1   g19961(.A1(new_n23008_), .A2(pi1156), .B(new_n23009_), .ZN(new_n23010_));
  INV_X1     g19962(.I(new_n23010_), .ZN(new_n23011_));
  OAI22_X1   g19963(.A1(new_n22992_), .A2(new_n22994_), .B1(new_n23006_), .B2(new_n23011_), .ZN(new_n23012_));
  MUX2_X1    g19964(.I0(new_n23012_), .I1(new_n22995_), .S(new_n11868_), .Z(new_n23013_));
  AOI22_X1   g19965(.A1(new_n22971_), .A2(new_n22967_), .B1(new_n22983_), .B2(new_n22989_), .ZN(new_n23014_));
  NAND3_X1   g19966(.A1(new_n23014_), .A2(pi0788), .A3(new_n22993_), .ZN(new_n23015_));
  OAI21_X1   g19967(.A1(new_n23014_), .A2(new_n11986_), .B(new_n22972_), .ZN(new_n23016_));
  AOI21_X1   g19968(.A1(new_n23016_), .A2(new_n23015_), .B(new_n23005_), .ZN(new_n23017_));
  NAND3_X1   g19969(.A1(new_n23017_), .A2(new_n22995_), .A3(pi0792), .ZN(new_n23018_));
  NAND2_X1   g19970(.A1(new_n23016_), .A2(new_n23015_), .ZN(new_n23019_));
  AOI22_X1   g19971(.A1(new_n23016_), .A2(new_n23015_), .B1(new_n23005_), .B2(new_n23010_), .ZN(new_n23020_));
  OAI21_X1   g19972(.A1(new_n23020_), .A2(new_n11868_), .B(new_n23019_), .ZN(new_n23021_));
  NAND2_X1   g19973(.A1(new_n23021_), .A2(new_n23018_), .ZN(new_n23022_));
  NOR2_X1    g19974(.A1(new_n22997_), .A2(new_n12053_), .ZN(new_n23023_));
  AOI21_X1   g19975(.A1(new_n12053_), .A2(new_n22895_), .B(new_n23023_), .ZN(new_n23024_));
  AOI21_X1   g19976(.A1(new_n23024_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n23025_));
  NOR4_X1    g19977(.A1(new_n23001_), .A2(new_n12031_), .A3(pi1156), .A4(new_n22878_), .ZN(new_n23026_));
  NOR2_X1    g19978(.A1(new_n23026_), .A2(new_n23002_), .ZN(new_n23027_));
  MUX2_X1    g19979(.I0(new_n23027_), .I1(new_n23001_), .S(new_n11868_), .Z(new_n23028_));
  NAND2_X1   g19980(.A1(new_n23028_), .A2(pi0647), .ZN(new_n23029_));
  NAND2_X1   g19981(.A1(new_n22878_), .A2(pi0647), .ZN(new_n23030_));
  NAND4_X1   g19982(.A1(new_n23029_), .A2(pi0630), .A3(new_n12049_), .A4(new_n23030_), .ZN(new_n23031_));
  INV_X1     g19983(.I(new_n23031_), .ZN(new_n23032_));
  NOR3_X1    g19984(.A1(new_n23032_), .A2(new_n12061_), .A3(new_n23025_), .ZN(new_n23033_));
  INV_X1     g19985(.I(new_n23033_), .ZN(new_n23034_));
  NOR3_X1    g19986(.A1(new_n23012_), .A2(new_n11868_), .A3(new_n23019_), .ZN(new_n23035_));
  AOI21_X1   g19987(.A1(new_n23012_), .A2(pi0792), .B(new_n22995_), .ZN(new_n23036_));
  NOR3_X1    g19988(.A1(new_n23035_), .A2(new_n23036_), .A3(pi0647), .ZN(new_n23037_));
  NAND2_X1   g19989(.A1(new_n23024_), .A2(pi0647), .ZN(new_n23038_));
  AOI21_X1   g19990(.A1(new_n22895_), .A2(new_n12061_), .B(pi1157), .ZN(new_n23039_));
  NAND2_X1   g19991(.A1(new_n23029_), .A2(new_n23039_), .ZN(new_n23040_));
  NAND2_X1   g19992(.A1(new_n23040_), .A2(new_n12060_), .ZN(new_n23041_));
  NAND3_X1   g19993(.A1(new_n23041_), .A2(new_n12049_), .A3(new_n23038_), .ZN(new_n23042_));
  OAI22_X1   g19994(.A1(new_n23037_), .A2(new_n23042_), .B1(new_n23022_), .B2(new_n23034_), .ZN(new_n23043_));
  MUX2_X1    g19995(.I0(new_n23043_), .I1(new_n23013_), .S(new_n12048_), .Z(new_n23044_));
  INV_X1     g19996(.I(new_n23028_), .ZN(new_n23045_));
  NOR3_X1    g19997(.A1(new_n22878_), .A2(pi0647), .A3(pi1157), .ZN(new_n23046_));
  MUX2_X1    g19998(.I0(new_n23046_), .I1(new_n23045_), .S(new_n12048_), .Z(new_n23047_));
  NAND2_X1   g19999(.A1(new_n23047_), .A2(pi0644), .ZN(new_n23048_));
  NOR2_X1    g20000(.A1(new_n22895_), .A2(new_n12092_), .ZN(new_n23049_));
  AOI21_X1   g20001(.A1(new_n23024_), .A2(new_n12092_), .B(new_n23049_), .ZN(new_n23050_));
  NAND2_X1   g20002(.A1(new_n12082_), .A2(new_n12099_), .ZN(new_n23051_));
  OR2_X2     g20003(.A1(new_n23050_), .A2(new_n23051_), .Z(new_n23052_));
  NAND3_X1   g20004(.A1(new_n23052_), .A2(new_n13168_), .A3(new_n23048_), .ZN(new_n23053_));
  AOI21_X1   g20005(.A1(new_n23044_), .A2(new_n12082_), .B(new_n23053_), .ZN(new_n23054_));
  NAND3_X1   g20006(.A1(new_n23021_), .A2(new_n23018_), .A3(new_n12061_), .ZN(new_n23055_));
  INV_X1     g20007(.I(new_n23042_), .ZN(new_n23056_));
  AOI22_X1   g20008(.A1(new_n23055_), .A2(new_n23056_), .B1(new_n23013_), .B2(new_n23033_), .ZN(new_n23057_));
  MUX2_X1    g20009(.I0(new_n23057_), .I1(new_n23022_), .S(new_n12048_), .Z(new_n23058_));
  NAND3_X1   g20010(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n23059_));
  OAI21_X1   g20011(.A1(new_n23050_), .A2(new_n23059_), .B(new_n13179_), .ZN(new_n23060_));
  NOR2_X1    g20012(.A1(new_n23060_), .A2(new_n23047_), .ZN(new_n23061_));
  OAI21_X1   g20013(.A1(new_n23058_), .A2(new_n12082_), .B(new_n23061_), .ZN(new_n23062_));
  NOR2_X1    g20014(.A1(new_n23054_), .A2(new_n23062_), .ZN(new_n23063_));
  NAND2_X1   g20015(.A1(po1038), .A2(new_n11628_), .ZN(new_n23064_));
  AOI21_X1   g20016(.A1(new_n23064_), .A2(new_n13184_), .B(po1038), .ZN(new_n23065_));
  OAI21_X1   g20017(.A1(new_n23044_), .A2(pi0790), .B(new_n23065_), .ZN(new_n23066_));
  OAI21_X1   g20018(.A1(new_n23063_), .A2(new_n23066_), .B(new_n22850_), .ZN(po0351));
  INV_X1     g20019(.I(new_n11844_), .ZN(new_n23068_));
  NAND4_X1   g20020(.A1(new_n7519_), .A2(new_n11572_), .A3(new_n5987_), .A4(new_n2587_), .ZN(new_n23070_));
  NAND4_X1   g20021(.A1(new_n11762_), .A2(pi0192), .A3(new_n11771_), .A4(new_n23070_), .ZN(new_n23071_));
  INV_X1     g20022(.I(new_n3319_), .ZN(new_n23072_));
  NAND2_X1   g20023(.A1(new_n11785_), .A2(pi0192), .ZN(new_n23073_));
  NOR2_X1    g20024(.A1(new_n11832_), .A2(pi0171), .ZN(new_n23074_));
  OAI21_X1   g20025(.A1(new_n11787_), .A2(new_n23074_), .B(new_n7170_), .ZN(new_n23075_));
  AOI21_X1   g20026(.A1(new_n11780_), .A2(new_n11572_), .B(new_n11837_), .ZN(new_n23076_));
  NAND3_X1   g20027(.A1(new_n23073_), .A2(new_n23075_), .A3(new_n23076_), .ZN(new_n23077_));
  AOI21_X1   g20028(.A1(new_n23077_), .A2(new_n11782_), .B(new_n23072_), .ZN(new_n23078_));
  AOI21_X1   g20029(.A1(new_n23071_), .A2(new_n23078_), .B(pi0087), .ZN(new_n23079_));
  OAI21_X1   g20030(.A1(new_n23079_), .A2(new_n11757_), .B(new_n3203_), .ZN(new_n23080_));
  AOI21_X1   g20031(.A1(new_n23080_), .A2(new_n11795_), .B(new_n23068_), .ZN(new_n23081_));
  NOR2_X1    g20032(.A1(new_n11818_), .A2(pi0138), .ZN(new_n23082_));
  INV_X1     g20033(.I(new_n23082_), .ZN(new_n23083_));
  NOR2_X1    g20034(.A1(new_n23083_), .A2(pi0196), .ZN(new_n23084_));
  NAND2_X1   g20035(.A1(new_n7681_), .A2(pi0195), .ZN(new_n23085_));
  OAI21_X1   g20036(.A1(new_n23085_), .A2(new_n23084_), .B(new_n2533_), .ZN(new_n23086_));
  NOR3_X1    g20037(.A1(new_n5143_), .A2(new_n3842_), .A3(new_n2587_), .ZN(new_n23087_));
  NOR2_X1    g20038(.A1(new_n11807_), .A2(new_n11572_), .ZN(new_n23088_));
  OAI21_X1   g20039(.A1(new_n11853_), .A2(new_n11572_), .B(new_n2587_), .ZN(new_n23089_));
  OAI22_X1   g20040(.A1(new_n23089_), .A2(new_n23088_), .B1(new_n8688_), .B2(new_n23087_), .ZN(new_n23090_));
  AOI21_X1   g20041(.A1(new_n5987_), .A2(new_n8691_), .B(new_n23090_), .ZN(new_n23091_));
  NAND3_X1   g20042(.A1(new_n23090_), .A2(new_n5987_), .A3(new_n8690_), .ZN(new_n23092_));
  OAI21_X1   g20043(.A1(new_n11802_), .A2(new_n11574_), .B(new_n3154_), .ZN(new_n23093_));
  NOR4_X1    g20044(.A1(new_n23083_), .A2(pi0195), .A3(pi0196), .A4(new_n7855_), .ZN(new_n23094_));
  AOI21_X1   g20045(.A1(new_n23093_), .A2(new_n23094_), .B(new_n3154_), .ZN(new_n23095_));
  NAND2_X1   g20046(.A1(new_n23092_), .A2(new_n23095_), .ZN(new_n23096_));
  OAI22_X1   g20047(.A1(new_n23081_), .A2(new_n23086_), .B1(new_n23091_), .B2(new_n23096_), .ZN(po0352));
  INV_X1     g20048(.I(new_n11756_), .ZN(new_n23098_));
  INV_X1     g20049(.I(new_n11797_), .ZN(new_n23099_));
  NOR2_X1    g20050(.A1(new_n11832_), .A2(pi0170), .ZN(new_n23100_));
  OAI21_X1   g20051(.A1(new_n11787_), .A2(new_n23100_), .B(new_n7170_), .ZN(new_n23101_));
  AOI21_X1   g20052(.A1(new_n23101_), .A2(new_n7597_), .B(new_n11779_), .ZN(new_n23102_));
  OAI21_X1   g20053(.A1(new_n23102_), .A2(new_n5987_), .B(new_n11782_), .ZN(new_n23103_));
  INV_X1     g20054(.I(new_n23103_), .ZN(new_n23104_));
  NOR2_X1    g20055(.A1(new_n11785_), .A2(new_n7178_), .ZN(new_n23105_));
  NOR2_X1    g20056(.A1(new_n11628_), .A2(pi0038), .ZN(new_n23106_));
  INV_X1     g20057(.I(new_n23106_), .ZN(new_n23107_));
  AOI21_X1   g20058(.A1(new_n23104_), .A2(new_n23105_), .B(new_n23107_), .ZN(new_n23108_));
  AND2_X2    g20059(.A1(new_n11761_), .A2(new_n23108_), .Z(new_n23109_));
  MUX2_X1    g20060(.I0(new_n7453_), .I1(new_n7406_), .S(new_n11630_), .Z(new_n23110_));
  NOR2_X1    g20061(.A1(pi0038), .A2(pi0194), .ZN(new_n23111_));
  OAI21_X1   g20062(.A1(new_n23104_), .A2(pi0039), .B(new_n23111_), .ZN(new_n23112_));
  AOI21_X1   g20063(.A1(new_n23112_), .A2(new_n11768_), .B(new_n11465_), .ZN(new_n23113_));
  NAND2_X1   g20064(.A1(new_n23110_), .A2(new_n23113_), .ZN(new_n23114_));
  NOR2_X1    g20065(.A1(new_n23108_), .A2(new_n23112_), .ZN(new_n23115_));
  OAI22_X1   g20066(.A1(new_n23109_), .A2(new_n23114_), .B1(new_n11770_), .B2(new_n23115_), .ZN(new_n23116_));
  AOI21_X1   g20067(.A1(new_n23116_), .A2(new_n3205_), .B(new_n11757_), .ZN(new_n23117_));
  OAI21_X1   g20068(.A1(new_n23117_), .A2(new_n23099_), .B(new_n3227_), .ZN(new_n23118_));
  NAND2_X1   g20069(.A1(new_n23118_), .A2(new_n23098_), .ZN(new_n23119_));
  AOI21_X1   g20070(.A1(new_n23119_), .A2(new_n2533_), .B(new_n7682_), .ZN(new_n23120_));
  NAND2_X1   g20071(.A1(new_n7171_), .A2(new_n3984_), .ZN(new_n23121_));
  NOR2_X1    g20072(.A1(new_n11806_), .A2(new_n10180_), .ZN(new_n23122_));
  AOI22_X1   g20073(.A1(new_n23122_), .A2(new_n23121_), .B1(new_n9702_), .B2(new_n11806_), .ZN(new_n23123_));
  MUX2_X1    g20074(.I0(new_n23123_), .I1(new_n8691_), .S(new_n5987_), .Z(new_n23124_));
  AOI21_X1   g20075(.A1(new_n11853_), .A2(new_n2587_), .B(new_n3154_), .ZN(new_n23125_));
  OAI21_X1   g20076(.A1(new_n23124_), .A2(new_n2587_), .B(new_n23125_), .ZN(new_n23126_));
  NAND2_X1   g20077(.A1(new_n11802_), .A2(new_n11631_), .ZN(new_n23127_));
  AOI21_X1   g20078(.A1(new_n23127_), .A2(new_n3154_), .B(pi0038), .ZN(new_n23128_));
  AOI21_X1   g20079(.A1(new_n23126_), .A2(new_n23128_), .B(new_n11628_), .ZN(new_n23129_));
  OAI21_X1   g20080(.A1(new_n11801_), .A2(new_n11663_), .B(new_n3154_), .ZN(new_n23130_));
  NAND2_X1   g20081(.A1(new_n23130_), .A2(new_n23106_), .ZN(new_n23131_));
  AOI21_X1   g20082(.A1(new_n23124_), .A2(pi0039), .B(new_n23131_), .ZN(new_n23132_));
  OAI21_X1   g20083(.A1(new_n23129_), .A2(new_n23132_), .B(new_n7832_), .ZN(new_n23133_));
  AOI21_X1   g20084(.A1(new_n23133_), .A2(new_n11820_), .B(new_n23082_), .ZN(new_n23134_));
  OAI21_X1   g20085(.A1(new_n23120_), .A2(new_n11820_), .B(new_n23134_), .ZN(new_n23135_));
  INV_X1     g20086(.I(new_n23120_), .ZN(new_n23136_));
  NOR2_X1    g20087(.A1(new_n11819_), .A2(pi0196), .ZN(new_n23137_));
  MUX2_X1    g20088(.I0(new_n23133_), .I1(new_n23136_), .S(new_n23137_), .Z(new_n23138_));
  OAI21_X1   g20089(.A1(new_n23138_), .A2(new_n23083_), .B(new_n23135_), .ZN(po0353));
  NOR2_X1    g20090(.A1(new_n15399_), .A2(new_n5339_), .ZN(new_n23140_));
  NAND2_X1   g20091(.A1(new_n15376_), .A2(new_n5339_), .ZN(new_n23141_));
  NAND3_X1   g20092(.A1(new_n15378_), .A2(new_n15145_), .A3(new_n23141_), .ZN(new_n23142_));
  NAND4_X1   g20093(.A1(new_n23142_), .A2(pi0197), .A3(new_n15145_), .A4(new_n6593_), .ZN(new_n23143_));
  NOR2_X1    g20094(.A1(new_n15367_), .A2(new_n23143_), .ZN(new_n23144_));
  OAI21_X1   g20095(.A1(new_n5339_), .A2(new_n15419_), .B(new_n23144_), .ZN(new_n23145_));
  OAI21_X1   g20096(.A1(new_n12852_), .A2(pi0197), .B(new_n3154_), .ZN(new_n23146_));
  NOR2_X1    g20097(.A1(new_n5473_), .A2(pi0767), .ZN(new_n23147_));
  NAND3_X1   g20098(.A1(new_n23146_), .A2(new_n12852_), .A3(new_n23147_), .ZN(new_n23148_));
  OAI22_X1   g20099(.A1(new_n23145_), .A2(new_n23140_), .B1(new_n15373_), .B2(new_n23148_), .ZN(new_n23149_));
  NAND2_X1   g20100(.A1(new_n13368_), .A2(new_n5339_), .ZN(new_n23150_));
  NOR4_X1    g20101(.A1(new_n15523_), .A2(pi0039), .A3(new_n15145_), .A4(new_n5473_), .ZN(new_n23151_));
  NOR2_X1    g20102(.A1(new_n23151_), .A2(new_n3172_), .ZN(new_n23152_));
  AOI22_X1   g20103(.A1(new_n23149_), .A2(new_n3172_), .B1(new_n23150_), .B2(new_n23152_), .ZN(new_n23153_));
  AOI21_X1   g20104(.A1(new_n15487_), .A2(new_n15489_), .B(new_n5339_), .ZN(new_n23154_));
  NAND2_X1   g20105(.A1(new_n23154_), .A2(pi0299), .ZN(new_n23155_));
  NOR2_X1    g20106(.A1(pi0039), .A2(pi0767), .ZN(new_n23156_));
  OAI21_X1   g20107(.A1(new_n12894_), .A2(pi0197), .B(new_n23156_), .ZN(new_n23157_));
  NAND2_X1   g20108(.A1(new_n15451_), .A2(new_n23141_), .ZN(new_n23158_));
  NAND4_X1   g20109(.A1(new_n23155_), .A2(new_n15145_), .A3(new_n23157_), .A4(new_n23158_), .ZN(new_n23159_));
  AOI21_X1   g20110(.A1(new_n12899_), .A2(pi0197), .B(pi0038), .ZN(new_n23161_));
  NAND3_X1   g20111(.A1(new_n23159_), .A2(new_n23148_), .A3(new_n23161_), .ZN(new_n23162_));
  AOI21_X1   g20112(.A1(new_n23162_), .A2(pi0698), .B(new_n7833_), .ZN(new_n23163_));
  OAI21_X1   g20113(.A1(new_n23153_), .A2(pi0698), .B(new_n23163_), .ZN(new_n23164_));
  AOI21_X1   g20114(.A1(new_n7833_), .A2(new_n5339_), .B(pi0832), .ZN(new_n23165_));
  AOI21_X1   g20115(.A1(new_n15051_), .A2(new_n15351_), .B(new_n23147_), .ZN(new_n23166_));
  MUX2_X1    g20116(.I0(new_n23166_), .I1(pi0197), .S(new_n2926_), .Z(new_n23167_));
  AOI22_X1   g20117(.A1(new_n23164_), .A2(new_n23165_), .B1(pi0832), .B2(new_n23167_), .ZN(po0354));
  OAI21_X1   g20118(.A1(new_n12852_), .A2(new_n2545_), .B(new_n13972_), .ZN(new_n23169_));
  NAND2_X1   g20119(.A1(new_n23169_), .A2(pi0198), .ZN(new_n23170_));
  NOR2_X1    g20120(.A1(new_n12132_), .A2(new_n2601_), .ZN(new_n23171_));
  INV_X1     g20121(.I(new_n23171_), .ZN(new_n23172_));
  NAND2_X1   g20122(.A1(new_n23172_), .A2(new_n2614_), .ZN(new_n23173_));
  OAI21_X1   g20123(.A1(new_n12809_), .A2(new_n2601_), .B(new_n5141_), .ZN(new_n23174_));
  NOR2_X1    g20124(.A1(new_n12495_), .A2(new_n2601_), .ZN(new_n23175_));
  NAND2_X1   g20125(.A1(new_n23175_), .A2(po1101), .ZN(new_n23176_));
  OAI21_X1   g20126(.A1(po1101), .A2(new_n23172_), .B(new_n23176_), .ZN(new_n23177_));
  AOI21_X1   g20127(.A1(new_n23177_), .A2(new_n5141_), .B(new_n2614_), .ZN(new_n23178_));
  AOI22_X1   g20128(.A1(new_n23178_), .A2(new_n23174_), .B1(new_n2604_), .B2(new_n23173_), .ZN(new_n23179_));
  OAI21_X1   g20129(.A1(new_n12809_), .A2(new_n2601_), .B(new_n5094_), .ZN(new_n23180_));
  AOI21_X1   g20130(.A1(new_n23177_), .A2(new_n5094_), .B(new_n3284_), .ZN(new_n23181_));
  NOR2_X1    g20131(.A1(new_n12473_), .A2(new_n2601_), .ZN(new_n23182_));
  INV_X1     g20132(.I(new_n23182_), .ZN(new_n23183_));
  AOI21_X1   g20133(.A1(new_n5107_), .A2(new_n23172_), .B(new_n23183_), .ZN(new_n23184_));
  OAI21_X1   g20134(.A1(new_n12464_), .A2(new_n12262_), .B(new_n5106_), .ZN(new_n23185_));
  NOR2_X1    g20135(.A1(new_n23185_), .A2(new_n2601_), .ZN(new_n23186_));
  AOI21_X1   g20136(.A1(new_n23186_), .A2(new_n6445_), .B(new_n23184_), .ZN(new_n23187_));
  NAND2_X1   g20137(.A1(new_n23172_), .A2(new_n3284_), .ZN(new_n23188_));
  AOI21_X1   g20138(.A1(new_n23188_), .A2(new_n2566_), .B(pi0299), .ZN(new_n23189_));
  OAI21_X1   g20139(.A1(new_n23187_), .A2(new_n2566_), .B(new_n23189_), .ZN(new_n23190_));
  AOI21_X1   g20140(.A1(new_n23181_), .A2(new_n23180_), .B(new_n23190_), .ZN(new_n23191_));
  AOI21_X1   g20141(.A1(new_n23186_), .A2(new_n6460_), .B(new_n23184_), .ZN(new_n23192_));
  NOR3_X1    g20142(.A1(new_n3232_), .A2(pi0299), .A3(new_n8533_), .ZN(new_n23193_));
  OAI21_X1   g20143(.A1(new_n23192_), .A2(new_n2604_), .B(new_n23193_), .ZN(new_n23194_));
  OR3_X2     g20144(.A1(new_n23179_), .A2(new_n23191_), .A3(new_n23194_), .Z(new_n23195_));
  NAND2_X1   g20145(.A1(new_n23170_), .A2(new_n23195_), .ZN(new_n23196_));
  NAND2_X1   g20146(.A1(new_n23196_), .A2(new_n12053_), .ZN(new_n23197_));
  INV_X1     g20147(.I(new_n23196_), .ZN(new_n23198_));
  NAND2_X1   g20148(.A1(new_n23198_), .A2(new_n11997_), .ZN(new_n23199_));
  NOR2_X1    g20149(.A1(new_n3231_), .A2(pi0198), .ZN(new_n23200_));
  INV_X1     g20150(.I(new_n23200_), .ZN(new_n23201_));
  INV_X1     g20151(.I(pi0633), .ZN(new_n23202_));
  NOR2_X1    g20152(.A1(new_n11875_), .A2(new_n23202_), .ZN(new_n23203_));
  MUX2_X1    g20153(.I0(pi0198), .I1(new_n23203_), .S(new_n12109_), .Z(new_n23204_));
  INV_X1     g20154(.I(new_n23204_), .ZN(new_n23205_));
  MUX2_X1    g20155(.I0(new_n23205_), .I1(pi0198), .S(pi0039), .Z(new_n23206_));
  NOR2_X1    g20156(.A1(new_n23206_), .A2(new_n3172_), .ZN(new_n23207_));
  NOR2_X1    g20157(.A1(new_n12590_), .A2(new_n2601_), .ZN(new_n23208_));
  INV_X1     g20158(.I(new_n23208_), .ZN(new_n23209_));
  NOR2_X1    g20159(.A1(new_n12613_), .A2(pi0198), .ZN(new_n23210_));
  AOI21_X1   g20160(.A1(pi0198), .A2(new_n12627_), .B(new_n23210_), .ZN(new_n23211_));
  NAND2_X1   g20161(.A1(new_n23202_), .A2(pi0603), .ZN(new_n23212_));
  MUX2_X1    g20162(.I0(new_n23211_), .I1(new_n23209_), .S(new_n23212_), .Z(new_n23213_));
  NAND2_X1   g20163(.A1(new_n13849_), .A2(new_n5101_), .ZN(new_n23214_));
  INV_X1     g20164(.I(new_n12565_), .ZN(new_n23215_));
  NOR2_X1    g20165(.A1(new_n23215_), .A2(new_n2601_), .ZN(new_n23216_));
  INV_X1     g20166(.I(new_n23216_), .ZN(new_n23217_));
  NOR2_X1    g20167(.A1(new_n12603_), .A2(new_n12582_), .ZN(new_n23218_));
  NAND2_X1   g20168(.A1(new_n23218_), .A2(pi0198), .ZN(new_n23219_));
  AOI21_X1   g20169(.A1(new_n23219_), .A2(new_n13343_), .B(new_n23202_), .ZN(new_n23220_));
  OAI21_X1   g20170(.A1(new_n13343_), .A2(new_n23219_), .B(new_n23220_), .ZN(new_n23221_));
  NAND2_X1   g20171(.A1(new_n23221_), .A2(new_n23217_), .ZN(new_n23222_));
  NAND2_X1   g20172(.A1(new_n23222_), .A2(new_n23214_), .ZN(new_n23223_));
  AOI21_X1   g20173(.A1(new_n2587_), .A2(new_n23223_), .B(new_n23213_), .ZN(new_n23224_));
  INV_X1     g20174(.I(new_n23223_), .ZN(new_n23225_));
  NAND3_X1   g20175(.A1(new_n23225_), .A2(new_n23213_), .A3(new_n2587_), .ZN(new_n23226_));
  INV_X1     g20176(.I(new_n23226_), .ZN(new_n23227_));
  NOR2_X1    g20177(.A1(new_n11873_), .A2(new_n23202_), .ZN(new_n23228_));
  NOR3_X1    g20178(.A1(new_n23228_), .A2(new_n2601_), .A3(new_n12132_), .ZN(new_n23229_));
  INV_X1     g20179(.I(new_n23228_), .ZN(new_n23230_));
  AOI21_X1   g20180(.A1(new_n2601_), .A2(new_n12133_), .B(new_n23230_), .ZN(new_n23231_));
  NOR2_X1    g20181(.A1(new_n23231_), .A2(new_n23229_), .ZN(new_n23232_));
  INV_X1     g20182(.I(new_n23232_), .ZN(new_n23233_));
  NOR2_X1    g20183(.A1(new_n23171_), .A2(pi0603), .ZN(new_n23234_));
  AOI21_X1   g20184(.A1(new_n23233_), .A2(pi0603), .B(new_n23234_), .ZN(new_n23235_));
  NAND2_X1   g20185(.A1(new_n23235_), .A2(new_n12168_), .ZN(new_n23236_));
  NOR2_X1    g20186(.A1(new_n23172_), .A2(pi0603), .ZN(new_n23237_));
  NOR3_X1    g20187(.A1(new_n12262_), .A2(new_n12133_), .A3(new_n23230_), .ZN(new_n23238_));
  AOI21_X1   g20188(.A1(new_n5108_), .A2(new_n23232_), .B(new_n23238_), .ZN(new_n23239_));
  AOI21_X1   g20189(.A1(new_n23183_), .A2(new_n23239_), .B(new_n5101_), .ZN(new_n23240_));
  OAI21_X1   g20190(.A1(new_n23240_), .A2(new_n23237_), .B(new_n12187_), .ZN(new_n23241_));
  XOR2_X1    g20191(.A1(new_n23241_), .A2(new_n23236_), .Z(new_n23242_));
  NOR2_X1    g20192(.A1(new_n23240_), .A2(new_n23182_), .ZN(new_n23243_));
  MUX2_X1    g20193(.I0(new_n23243_), .I1(new_n23242_), .S(new_n5217_), .Z(new_n23244_));
  INV_X1     g20194(.I(new_n23244_), .ZN(new_n23245_));
  AND3_X2    g20195(.A1(new_n12250_), .A2(pi0633), .A3(new_n12251_), .Z(new_n23246_));
  NOR2_X1    g20196(.A1(new_n23246_), .A2(new_n23186_), .ZN(new_n23247_));
  NOR2_X1    g20197(.A1(new_n12242_), .A2(new_n2601_), .ZN(new_n23248_));
  NOR2_X1    g20198(.A1(new_n23238_), .A2(new_n23248_), .ZN(new_n23249_));
  NOR2_X1    g20199(.A1(new_n23249_), .A2(new_n12797_), .ZN(new_n23250_));
  MUX2_X1    g20200(.I0(new_n23250_), .I1(new_n23247_), .S(new_n5217_), .Z(new_n23251_));
  AOI21_X1   g20201(.A1(new_n23251_), .A2(new_n6460_), .B(pi0223), .ZN(new_n23252_));
  OAI21_X1   g20202(.A1(new_n23245_), .A2(new_n6460_), .B(new_n23252_), .ZN(new_n23253_));
  NOR2_X1    g20203(.A1(new_n12156_), .A2(new_n2601_), .ZN(new_n23254_));
  AOI21_X1   g20204(.A1(pi0633), .A2(new_n12170_), .B(new_n23254_), .ZN(new_n23255_));
  NOR4_X1    g20205(.A1(new_n23255_), .A2(pi0603), .A3(new_n5109_), .A4(new_n23233_), .ZN(new_n23256_));
  AOI21_X1   g20206(.A1(new_n23232_), .A2(new_n5105_), .B(new_n5101_), .ZN(new_n23257_));
  NOR4_X1    g20207(.A1(new_n23233_), .A2(new_n5101_), .A3(pi0642), .A4(new_n5104_), .ZN(new_n23258_));
  OAI21_X1   g20208(.A1(new_n23234_), .A2(new_n23257_), .B(new_n23258_), .ZN(new_n23259_));
  INV_X1     g20209(.I(new_n23259_), .ZN(new_n23260_));
  OAI21_X1   g20210(.A1(new_n23256_), .A2(pi0642), .B(new_n23260_), .ZN(new_n23261_));
  NAND2_X1   g20211(.A1(new_n23261_), .A2(new_n5217_), .ZN(new_n23262_));
  AOI21_X1   g20212(.A1(new_n5101_), .A2(new_n23175_), .B(new_n23256_), .ZN(new_n23263_));
  NOR2_X1    g20213(.A1(new_n23263_), .A2(new_n5217_), .ZN(new_n23264_));
  XOR2_X1    g20214(.A1(new_n23264_), .A2(new_n23262_), .Z(new_n23265_));
  NAND3_X1   g20215(.A1(new_n12158_), .A2(pi0198), .A3(new_n5101_), .ZN(new_n23266_));
  NOR2_X1    g20216(.A1(pi0332), .A2(pi0468), .ZN(new_n23267_));
  NAND2_X1   g20217(.A1(new_n23255_), .A2(new_n23267_), .ZN(new_n23268_));
  NOR2_X1    g20218(.A1(new_n23255_), .A2(new_n5101_), .ZN(new_n23269_));
  AOI22_X1   g20219(.A1(new_n12187_), .A2(new_n23269_), .B1(new_n23268_), .B2(new_n23266_), .ZN(new_n23270_));
  NOR2_X1    g20220(.A1(new_n23269_), .A2(new_n23254_), .ZN(new_n23271_));
  MUX2_X1    g20221(.I0(new_n23271_), .I1(new_n23270_), .S(new_n5217_), .Z(new_n23272_));
  OAI21_X1   g20222(.A1(new_n23272_), .A2(new_n5141_), .B(new_n23265_), .ZN(new_n23273_));
  INV_X1     g20223(.I(new_n23265_), .ZN(new_n23274_));
  NAND3_X1   g20224(.A1(new_n23274_), .A2(new_n6460_), .A3(new_n23272_), .ZN(new_n23275_));
  NOR2_X1    g20225(.A1(new_n2614_), .A2(pi0223), .ZN(new_n23276_));
  NAND3_X1   g20226(.A1(new_n23275_), .A2(new_n23273_), .A3(new_n23276_), .ZN(new_n23277_));
  AOI21_X1   g20227(.A1(new_n23277_), .A2(new_n23253_), .B(pi0299), .ZN(new_n23278_));
  AOI21_X1   g20228(.A1(new_n23251_), .A2(new_n6445_), .B(pi0215), .ZN(new_n23279_));
  OAI21_X1   g20229(.A1(new_n23245_), .A2(new_n6445_), .B(new_n23279_), .ZN(new_n23280_));
  OAI21_X1   g20230(.A1(new_n23272_), .A2(new_n5094_), .B(new_n23265_), .ZN(new_n23281_));
  NAND3_X1   g20231(.A1(new_n23274_), .A2(new_n6445_), .A3(new_n23272_), .ZN(new_n23282_));
  NOR2_X1    g20232(.A1(new_n3284_), .A2(pi0215), .ZN(new_n23283_));
  NAND4_X1   g20233(.A1(new_n23282_), .A2(new_n23280_), .A3(new_n23281_), .A4(new_n23283_), .ZN(new_n23284_));
  NAND2_X1   g20234(.A1(new_n23284_), .A2(new_n13820_), .ZN(new_n23285_));
  NOR2_X1    g20235(.A1(new_n23278_), .A2(new_n23285_), .ZN(new_n23286_));
  NOR4_X1    g20236(.A1(new_n23286_), .A2(pi0039), .A3(new_n23224_), .A4(new_n23227_), .ZN(new_n23287_));
  NOR2_X1    g20237(.A1(new_n23287_), .A2(pi0038), .ZN(new_n23288_));
  OAI21_X1   g20238(.A1(new_n23288_), .A2(new_n23207_), .B(new_n3231_), .ZN(new_n23289_));
  XOR2_X1    g20239(.A1(new_n23289_), .A2(new_n23201_), .Z(new_n23290_));
  AOI21_X1   g20240(.A1(new_n23196_), .A2(new_n11914_), .B(pi0785), .ZN(new_n23291_));
  OAI21_X1   g20241(.A1(new_n23290_), .A2(new_n11914_), .B(new_n23291_), .ZN(new_n23292_));
  OAI21_X1   g20242(.A1(new_n23290_), .A2(new_n12996_), .B(new_n23196_), .ZN(new_n23293_));
  NAND3_X1   g20243(.A1(new_n23290_), .A2(new_n12997_), .A3(new_n23198_), .ZN(new_n23294_));
  NAND3_X1   g20244(.A1(new_n23293_), .A2(new_n23294_), .A3(new_n11912_), .ZN(new_n23295_));
  INV_X1     g20245(.I(new_n23290_), .ZN(new_n23296_));
  OAI21_X1   g20246(.A1(new_n13010_), .A2(new_n23198_), .B(new_n23296_), .ZN(new_n23297_));
  NAND3_X1   g20247(.A1(new_n23290_), .A2(new_n11915_), .A3(new_n23198_), .ZN(new_n23298_));
  NAND3_X1   g20248(.A1(new_n23297_), .A2(pi1155), .A3(new_n23298_), .ZN(new_n23299_));
  AOI21_X1   g20249(.A1(new_n23299_), .A2(new_n23295_), .B(new_n11870_), .ZN(new_n23300_));
  XNOR2_X1   g20250(.A1(new_n23300_), .A2(new_n23292_), .ZN(new_n23301_));
  NOR3_X1    g20251(.A1(new_n23196_), .A2(pi0618), .A3(pi1154), .ZN(new_n23302_));
  INV_X1     g20252(.I(new_n23302_), .ZN(new_n23303_));
  MUX2_X1    g20253(.I0(new_n23303_), .I1(new_n23301_), .S(new_n11969_), .Z(new_n23304_));
  INV_X1     g20254(.I(new_n23304_), .ZN(new_n23305_));
  NOR3_X1    g20255(.A1(new_n23196_), .A2(pi0619), .A3(pi1159), .ZN(new_n23306_));
  MUX2_X1    g20256(.I0(new_n23306_), .I1(new_n23305_), .S(new_n11985_), .Z(new_n23307_));
  OAI21_X1   g20257(.A1(new_n23307_), .A2(new_n11997_), .B(new_n23199_), .ZN(new_n23308_));
  OAI21_X1   g20258(.A1(new_n23308_), .A2(new_n12053_), .B(new_n23197_), .ZN(new_n23309_));
  NOR2_X1    g20259(.A1(new_n23309_), .A2(new_n15077_), .ZN(new_n23310_));
  INV_X1     g20260(.I(new_n23310_), .ZN(new_n23311_));
  NOR2_X1    g20261(.A1(new_n23198_), .A2(new_n11961_), .ZN(new_n23312_));
  NOR2_X1    g20262(.A1(new_n23196_), .A2(new_n11938_), .ZN(new_n23313_));
  NAND2_X1   g20263(.A1(new_n11884_), .A2(pi0634), .ZN(new_n23314_));
  MUX2_X1    g20264(.I0(new_n2601_), .I1(new_n23314_), .S(new_n12109_), .Z(new_n23315_));
  MUX2_X1    g20265(.I0(new_n23315_), .I1(pi0198), .S(pi0039), .Z(new_n23316_));
  NOR2_X1    g20266(.A1(new_n23316_), .A2(new_n3172_), .ZN(new_n23317_));
  INV_X1     g20267(.I(pi0634), .ZN(new_n23318_));
  NOR2_X1    g20268(.A1(new_n12655_), .A2(new_n2601_), .ZN(new_n23319_));
  AOI21_X1   g20269(.A1(new_n2601_), .A2(new_n12630_), .B(new_n23319_), .ZN(new_n23320_));
  NOR3_X1    g20270(.A1(new_n23320_), .A2(new_n23318_), .A3(new_n5095_), .ZN(new_n23321_));
  NOR2_X1    g20271(.A1(new_n23318_), .A2(new_n5095_), .ZN(new_n23322_));
  OAI21_X1   g20272(.A1(new_n23208_), .A2(new_n23322_), .B(pi0299), .ZN(new_n23323_));
  OAI21_X1   g20273(.A1(new_n12638_), .A2(pi0198), .B(new_n23322_), .ZN(new_n23324_));
  NOR3_X1    g20274(.A1(new_n12564_), .A2(new_n2601_), .A3(new_n11882_), .ZN(new_n23325_));
  AOI21_X1   g20275(.A1(new_n23325_), .A2(new_n23324_), .B(new_n23216_), .ZN(new_n23326_));
  AOI21_X1   g20276(.A1(new_n23326_), .A2(new_n2587_), .B(pi0039), .ZN(new_n23327_));
  OAI21_X1   g20277(.A1(new_n23321_), .A2(new_n23323_), .B(new_n23327_), .ZN(new_n23328_));
  INV_X1     g20278(.I(new_n12161_), .ZN(new_n23329_));
  AOI21_X1   g20279(.A1(pi0634), .A2(new_n23329_), .B(new_n23254_), .ZN(new_n23330_));
  INV_X1     g20280(.I(new_n23330_), .ZN(new_n23331_));
  NOR2_X1    g20281(.A1(new_n12160_), .A2(new_n23318_), .ZN(new_n23332_));
  NOR2_X1    g20282(.A1(new_n23332_), .A2(new_n23171_), .ZN(new_n23333_));
  NOR2_X1    g20283(.A1(new_n23333_), .A2(new_n5108_), .ZN(new_n23334_));
  AOI21_X1   g20284(.A1(new_n23331_), .A2(new_n5108_), .B(new_n23334_), .ZN(new_n23335_));
  INV_X1     g20285(.I(new_n23335_), .ZN(new_n23336_));
  MUX2_X1    g20286(.I0(new_n23331_), .I1(new_n23336_), .S(new_n5427_), .Z(new_n23337_));
  OAI22_X1   g20287(.A1(new_n12424_), .A2(new_n2601_), .B1(new_n23331_), .B2(new_n5100_), .ZN(new_n23338_));
  AOI21_X1   g20288(.A1(new_n23337_), .A2(new_n12130_), .B(new_n23338_), .ZN(new_n23339_));
  NAND2_X1   g20289(.A1(new_n12242_), .A2(new_n23332_), .ZN(new_n23340_));
  XOR2_X1    g20290(.A1(new_n23248_), .A2(new_n23340_), .Z(new_n23341_));
  INV_X1     g20291(.I(new_n23341_), .ZN(new_n23342_));
  AOI21_X1   g20292(.A1(new_n23341_), .A2(new_n5108_), .B(new_n23334_), .ZN(new_n23343_));
  MUX2_X1    g20293(.I0(new_n23342_), .I1(new_n23343_), .S(new_n5427_), .Z(new_n23344_));
  NOR2_X1    g20294(.A1(new_n23344_), .A2(new_n12222_), .ZN(new_n23345_));
  NAND2_X1   g20295(.A1(new_n23186_), .A2(new_n5095_), .ZN(new_n23346_));
  OAI21_X1   g20296(.A1(new_n5100_), .A2(new_n23341_), .B(new_n23346_), .ZN(new_n23347_));
  NOR2_X1    g20297(.A1(new_n23345_), .A2(new_n23347_), .ZN(new_n23348_));
  NOR2_X1    g20298(.A1(new_n23346_), .A2(new_n23183_), .ZN(new_n23349_));
  INV_X1     g20299(.I(new_n23333_), .ZN(new_n23350_));
  NOR2_X1    g20300(.A1(new_n23350_), .A2(new_n5109_), .ZN(new_n23351_));
  INV_X1     g20301(.I(new_n23351_), .ZN(new_n23352_));
  OAI21_X1   g20302(.A1(new_n23341_), .A2(new_n5108_), .B(new_n23352_), .ZN(new_n23353_));
  NOR2_X1    g20303(.A1(new_n23353_), .A2(new_n5427_), .ZN(new_n23354_));
  OAI21_X1   g20304(.A1(new_n23333_), .A2(new_n5106_), .B(new_n12222_), .ZN(new_n23355_));
  OAI22_X1   g20305(.A1(new_n23354_), .A2(new_n23355_), .B1(new_n5217_), .B2(new_n23353_), .ZN(new_n23356_));
  NOR2_X1    g20306(.A1(new_n23356_), .A2(new_n23349_), .ZN(new_n23357_));
  NAND4_X1   g20307(.A1(new_n23348_), .A2(new_n2566_), .A3(new_n5094_), .A4(new_n23357_), .ZN(new_n23358_));
  AOI21_X1   g20308(.A1(new_n23330_), .A2(new_n5109_), .B(new_n23351_), .ZN(new_n23359_));
  AOI21_X1   g20309(.A1(new_n23359_), .A2(new_n5106_), .B(new_n23355_), .ZN(new_n23360_));
  NOR2_X1    g20310(.A1(new_n23175_), .A2(new_n5427_), .ZN(new_n23361_));
  OAI21_X1   g20311(.A1(new_n5106_), .A2(new_n23171_), .B(new_n5095_), .ZN(new_n23362_));
  OAI22_X1   g20312(.A1(new_n23359_), .A2(new_n5100_), .B1(new_n23361_), .B2(new_n23362_), .ZN(new_n23363_));
  NOR2_X1    g20313(.A1(new_n23363_), .A2(new_n23360_), .ZN(new_n23364_));
  NAND2_X1   g20314(.A1(new_n23364_), .A2(new_n5094_), .ZN(new_n23365_));
  AOI21_X1   g20315(.A1(new_n23332_), .A2(pi0680), .B(new_n23171_), .ZN(new_n23366_));
  NOR3_X1    g20316(.A1(new_n3284_), .A2(new_n2566_), .A3(pi0299), .ZN(new_n23367_));
  NAND3_X1   g20317(.A1(new_n23358_), .A2(new_n23365_), .A3(new_n23367_), .ZN(new_n23368_));
  AOI21_X1   g20318(.A1(new_n6445_), .A2(new_n23339_), .B(new_n23368_), .ZN(new_n23369_));
  NAND2_X1   g20319(.A1(new_n23339_), .A2(new_n6460_), .ZN(new_n23370_));
  AOI21_X1   g20320(.A1(new_n23364_), .A2(new_n5141_), .B(new_n2614_), .ZN(new_n23371_));
  NAND4_X1   g20321(.A1(new_n23348_), .A2(new_n2604_), .A3(new_n5141_), .A4(new_n23357_), .ZN(new_n23372_));
  NOR2_X1    g20322(.A1(new_n23366_), .A2(new_n3155_), .ZN(new_n23373_));
  NOR2_X1    g20323(.A1(new_n23373_), .A2(new_n3294_), .ZN(new_n23374_));
  NAND2_X1   g20324(.A1(new_n23372_), .A2(new_n23374_), .ZN(new_n23375_));
  AOI21_X1   g20325(.A1(new_n23370_), .A2(new_n23371_), .B(new_n23375_), .ZN(new_n23376_));
  OAI21_X1   g20326(.A1(new_n23376_), .A2(new_n23369_), .B(pi0039), .ZN(new_n23377_));
  AOI21_X1   g20327(.A1(new_n23377_), .A2(new_n23328_), .B(pi0038), .ZN(new_n23378_));
  OAI21_X1   g20328(.A1(new_n23378_), .A2(new_n23317_), .B(new_n3231_), .ZN(new_n23379_));
  XOR2_X1    g20329(.A1(new_n23379_), .A2(new_n23201_), .Z(new_n23380_));
  NAND3_X1   g20330(.A1(new_n23198_), .A2(new_n12970_), .A3(new_n11893_), .ZN(new_n23381_));
  MUX2_X1    g20331(.I0(new_n23381_), .I1(new_n23380_), .S(new_n11891_), .Z(new_n23382_));
  AOI21_X1   g20332(.A1(new_n23382_), .A2(new_n11938_), .B(new_n23313_), .ZN(new_n23383_));
  AOI21_X1   g20333(.A1(new_n23383_), .A2(new_n11961_), .B(new_n23312_), .ZN(new_n23384_));
  INV_X1     g20334(.I(new_n23384_), .ZN(new_n23385_));
  MUX2_X1    g20335(.I0(new_n23198_), .I1(new_n23385_), .S(new_n13713_), .Z(new_n23386_));
  NOR2_X1    g20336(.A1(new_n23386_), .A2(new_n12031_), .ZN(new_n23387_));
  AOI21_X1   g20337(.A1(new_n12031_), .A2(new_n23198_), .B(new_n23387_), .ZN(new_n23388_));
  NOR2_X1    g20338(.A1(new_n23388_), .A2(new_n12026_), .ZN(new_n23389_));
  NOR3_X1    g20339(.A1(new_n23198_), .A2(new_n12031_), .A3(new_n12026_), .ZN(new_n23390_));
  NOR3_X1    g20340(.A1(new_n23389_), .A2(new_n11868_), .A3(new_n23390_), .ZN(new_n23391_));
  AOI21_X1   g20341(.A1(new_n11868_), .A2(new_n23386_), .B(new_n23391_), .ZN(new_n23392_));
  INV_X1     g20342(.I(new_n23392_), .ZN(new_n23393_));
  NOR2_X1    g20343(.A1(new_n23393_), .A2(new_n12061_), .ZN(new_n23394_));
  NOR2_X1    g20344(.A1(new_n23198_), .A2(new_n12061_), .ZN(new_n23395_));
  NOR3_X1    g20345(.A1(new_n23394_), .A2(pi1157), .A3(new_n23395_), .ZN(new_n23396_));
  INV_X1     g20346(.I(new_n23396_), .ZN(new_n23397_));
  NOR2_X1    g20347(.A1(new_n23198_), .A2(pi0647), .ZN(new_n23398_));
  AOI21_X1   g20348(.A1(new_n23393_), .A2(pi0647), .B(new_n23398_), .ZN(new_n23399_));
  AOI22_X1   g20349(.A1(new_n23397_), .A2(pi0630), .B1(new_n12088_), .B2(new_n23399_), .ZN(new_n23400_));
  AOI21_X1   g20350(.A1(new_n23311_), .A2(new_n23400_), .B(new_n12048_), .ZN(new_n23401_));
  INV_X1     g20351(.I(new_n12050_), .ZN(new_n23402_));
  INV_X1     g20352(.I(new_n23390_), .ZN(new_n23403_));
  OAI22_X1   g20353(.A1(new_n23388_), .A2(new_n23402_), .B1(new_n12030_), .B2(new_n23403_), .ZN(new_n23404_));
  AOI21_X1   g20354(.A1(new_n23308_), .A2(new_n15222_), .B(new_n23404_), .ZN(new_n23405_));
  NAND2_X1   g20355(.A1(new_n23405_), .A2(pi0792), .ZN(new_n23406_));
  NOR2_X1    g20356(.A1(new_n23305_), .A2(new_n11967_), .ZN(new_n23407_));
  OAI21_X1   g20357(.A1(new_n23198_), .A2(new_n11967_), .B(new_n11869_), .ZN(new_n23408_));
  OR3_X2     g20358(.A1(new_n23407_), .A2(new_n11966_), .A3(new_n23408_), .Z(new_n23409_));
  NAND2_X1   g20359(.A1(new_n23359_), .A2(new_n5101_), .ZN(new_n23410_));
  NOR4_X1    g20360(.A1(new_n23233_), .A2(new_n23318_), .A3(pi0665), .A4(new_n12292_), .ZN(new_n23411_));
  NOR3_X1    g20361(.A1(new_n23411_), .A2(pi0603), .A3(new_n5109_), .ZN(new_n23412_));
  OAI21_X1   g20362(.A1(new_n23318_), .A2(new_n12485_), .B(new_n23255_), .ZN(new_n23413_));
  AOI21_X1   g20363(.A1(new_n23413_), .A2(new_n23412_), .B(new_n12461_), .ZN(new_n23414_));
  AOI21_X1   g20364(.A1(new_n23413_), .A2(new_n23412_), .B(new_n12384_), .ZN(new_n23415_));
  NOR2_X1    g20365(.A1(new_n23411_), .A2(new_n5101_), .ZN(new_n23416_));
  INV_X1     g20366(.I(new_n23416_), .ZN(new_n23417_));
  NOR2_X1    g20367(.A1(new_n23417_), .A2(new_n12384_), .ZN(new_n23418_));
  NOR2_X1    g20368(.A1(new_n23333_), .A2(pi0603), .ZN(new_n23419_));
  NOR4_X1    g20369(.A1(new_n23415_), .A2(new_n5105_), .A3(new_n23418_), .A4(new_n23419_), .ZN(new_n23420_));
  INV_X1     g20370(.I(new_n23420_), .ZN(new_n23421_));
  NOR2_X1    g20371(.A1(new_n23416_), .A2(new_n23419_), .ZN(new_n23422_));
  INV_X1     g20372(.I(new_n23422_), .ZN(new_n23423_));
  AOI21_X1   g20373(.A1(new_n23423_), .A2(new_n5105_), .B(new_n12129_), .ZN(new_n23424_));
  AOI22_X1   g20374(.A1(new_n23421_), .A2(new_n23424_), .B1(new_n23414_), .B2(new_n23410_), .ZN(new_n23425_));
  MUX2_X1    g20375(.I0(new_n23425_), .I1(new_n23261_), .S(new_n5095_), .Z(new_n23426_));
  NOR4_X1    g20376(.A1(new_n23232_), .A2(pi0603), .A3(new_n5108_), .A4(new_n12187_), .ZN(new_n23429_));
  AOI21_X1   g20377(.A1(new_n23416_), .A2(new_n12168_), .B(new_n23429_), .ZN(new_n23430_));
  NOR2_X1    g20378(.A1(new_n23430_), .A2(new_n5108_), .ZN(new_n23431_));
  OR3_X2     g20379(.A1(new_n23426_), .A2(new_n3285_), .A3(new_n6445_), .Z(new_n23438_));
  NOR3_X1    g20380(.A1(new_n12212_), .A2(new_n2601_), .A3(pi0665), .ZN(new_n23439_));
  NOR2_X1    g20381(.A1(pi0198), .A2(pi0665), .ZN(new_n23440_));
  INV_X1     g20382(.I(new_n23440_), .ZN(new_n23441_));
  NOR2_X1    g20383(.A1(new_n12290_), .A2(new_n23441_), .ZN(new_n23442_));
  NOR3_X1    g20384(.A1(new_n23442_), .A2(new_n23248_), .A3(new_n23439_), .ZN(new_n23443_));
  AND3_X2    g20385(.A1(new_n23443_), .A2(new_n23318_), .A3(new_n23248_), .Z(new_n23444_));
  INV_X1     g20386(.I(new_n23248_), .ZN(new_n23445_));
  AOI21_X1   g20387(.A1(new_n23318_), .A2(new_n23445_), .B(new_n23443_), .ZN(new_n23446_));
  NOR3_X1    g20388(.A1(new_n23444_), .A2(new_n23238_), .A3(new_n23446_), .ZN(new_n23447_));
  NAND3_X1   g20389(.A1(new_n23429_), .A2(pi0603), .A3(new_n12187_), .ZN(new_n23448_));
  NAND2_X1   g20390(.A1(new_n23447_), .A2(new_n23448_), .ZN(new_n23449_));
  NOR2_X1    g20391(.A1(new_n23343_), .A2(pi0603), .ZN(new_n23450_));
  NOR2_X1    g20392(.A1(new_n23450_), .A2(new_n23431_), .ZN(new_n23451_));
  AOI21_X1   g20393(.A1(new_n23451_), .A2(new_n23449_), .B(new_n12222_), .ZN(new_n23452_));
  OAI21_X1   g20394(.A1(new_n23342_), .A2(pi0603), .B(new_n5217_), .ZN(new_n23453_));
  AOI21_X1   g20395(.A1(new_n23447_), .A2(pi0603), .B(new_n23453_), .ZN(new_n23454_));
  NOR3_X1    g20396(.A1(new_n23246_), .A2(pi0680), .A3(new_n23186_), .ZN(new_n23455_));
  OAI21_X1   g20397(.A1(new_n23452_), .A2(new_n23454_), .B(new_n23455_), .ZN(new_n23456_));
  NAND2_X1   g20398(.A1(new_n23456_), .A2(new_n6445_), .ZN(new_n23457_));
  NAND2_X1   g20399(.A1(new_n23447_), .A2(new_n23412_), .ZN(new_n23458_));
  INV_X1     g20400(.I(new_n23458_), .ZN(new_n23459_));
  AOI21_X1   g20401(.A1(new_n23423_), .A2(new_n12130_), .B(new_n12187_), .ZN(new_n23460_));
  OAI21_X1   g20402(.A1(new_n23459_), .A2(new_n23419_), .B(new_n23460_), .ZN(new_n23461_));
  NOR2_X1    g20403(.A1(new_n23353_), .A2(pi0603), .ZN(new_n23462_));
  OR3_X2     g20404(.A1(new_n23459_), .A2(new_n5100_), .A3(new_n23462_), .Z(new_n23463_));
  OR2_X2     g20405(.A1(new_n23242_), .A2(pi0680), .Z(new_n23464_));
  AND3_X2    g20406(.A1(new_n23464_), .A2(new_n23461_), .A3(new_n23463_), .Z(new_n23465_));
  AOI21_X1   g20407(.A1(new_n23465_), .A2(new_n5094_), .B(pi0215), .ZN(new_n23466_));
  INV_X1     g20408(.I(new_n23235_), .ZN(new_n23467_));
  NOR2_X1    g20409(.A1(new_n12159_), .A2(new_n23171_), .ZN(new_n23468_));
  NOR4_X1    g20410(.A1(new_n23467_), .A2(new_n23318_), .A3(new_n12114_), .A4(new_n23468_), .ZN(new_n23469_));
  NAND2_X1   g20411(.A1(new_n23469_), .A2(new_n3284_), .ZN(new_n23470_));
  NAND2_X1   g20412(.A1(new_n23470_), .A2(new_n2566_), .ZN(new_n23471_));
  AOI21_X1   g20413(.A1(new_n23466_), .A2(new_n23457_), .B(new_n23471_), .ZN(new_n23472_));
  AOI21_X1   g20414(.A1(new_n23438_), .A2(new_n23472_), .B(new_n15651_), .ZN(new_n23473_));
  NOR3_X1    g20415(.A1(new_n23426_), .A2(new_n3155_), .A3(new_n6460_), .ZN(new_n23474_));
  NAND2_X1   g20416(.A1(new_n23456_), .A2(new_n6460_), .ZN(new_n23475_));
  NAND2_X1   g20417(.A1(new_n23465_), .A2(new_n5141_), .ZN(new_n23476_));
  NAND3_X1   g20418(.A1(new_n23476_), .A2(new_n2604_), .A3(new_n23475_), .ZN(new_n23477_));
  NAND2_X1   g20419(.A1(new_n23469_), .A2(new_n2614_), .ZN(new_n23478_));
  NAND3_X1   g20420(.A1(new_n23477_), .A2(new_n2604_), .A3(new_n23478_), .ZN(new_n23479_));
  OAI21_X1   g20421(.A1(new_n23479_), .A2(new_n23474_), .B(new_n2587_), .ZN(new_n23480_));
  NOR2_X1    g20422(.A1(new_n23473_), .A2(new_n23480_), .ZN(new_n23481_));
  NOR3_X1    g20423(.A1(new_n23318_), .A2(new_n5095_), .A3(pi0299), .ZN(new_n23482_));
  MUX2_X1    g20424(.I0(new_n12641_), .I1(pi0665), .S(new_n2601_), .Z(new_n23483_));
  NOR2_X1    g20425(.A1(new_n23211_), .A2(pi0633), .ZN(new_n23484_));
  INV_X1     g20426(.I(new_n12613_), .ZN(new_n23485_));
  NAND2_X1   g20427(.A1(new_n23485_), .A2(new_n12655_), .ZN(new_n23486_));
  NAND2_X1   g20428(.A1(new_n2601_), .A2(new_n23202_), .ZN(new_n23487_));
  AOI21_X1   g20429(.A1(new_n12658_), .A2(new_n23441_), .B(new_n23487_), .ZN(new_n23488_));
  AOI22_X1   g20430(.A1(new_n23484_), .A2(new_n23483_), .B1(new_n23486_), .B2(new_n23488_), .ZN(new_n23489_));
  MUX2_X1    g20431(.I0(new_n23489_), .I1(new_n23320_), .S(new_n5101_), .Z(new_n23490_));
  NOR2_X1    g20432(.A1(new_n12564_), .A2(new_n11882_), .ZN(new_n23491_));
  NOR3_X1    g20433(.A1(new_n12605_), .A2(new_n23491_), .A3(new_n2601_), .ZN(new_n23492_));
  INV_X1     g20434(.I(new_n23492_), .ZN(new_n23493_));
  AOI21_X1   g20435(.A1(new_n23217_), .A2(new_n23318_), .B(new_n23493_), .ZN(new_n23494_));
  NOR3_X1    g20436(.A1(new_n23217_), .A2(pi0634), .A3(new_n23492_), .ZN(new_n23495_));
  NOR3_X1    g20437(.A1(new_n23495_), .A2(new_n23494_), .A3(pi0633), .ZN(new_n23496_));
  OAI21_X1   g20438(.A1(new_n23326_), .A2(pi0603), .B(pi0680), .ZN(new_n23497_));
  NOR4_X1    g20439(.A1(new_n2601_), .A2(pi0633), .A3(pi0634), .A4(pi0665), .ZN(new_n23498_));
  NOR2_X1    g20440(.A1(new_n23498_), .A2(pi0603), .ZN(new_n23499_));
  NAND4_X1   g20441(.A1(new_n23497_), .A2(new_n13342_), .A3(new_n23221_), .A4(new_n23499_), .ZN(new_n23500_));
  AOI21_X1   g20442(.A1(new_n23225_), .A2(new_n5095_), .B(new_n6594_), .ZN(new_n23501_));
  OAI21_X1   g20443(.A1(new_n23496_), .A2(new_n23500_), .B(new_n23501_), .ZN(new_n23502_));
  AOI21_X1   g20444(.A1(new_n23490_), .A2(new_n23482_), .B(new_n23502_), .ZN(new_n23503_));
  OAI21_X1   g20445(.A1(new_n23503_), .A2(new_n23481_), .B(new_n3172_), .ZN(new_n23507_));
  NAND2_X1   g20446(.A1(new_n23507_), .A2(new_n3231_), .ZN(new_n23508_));
  XOR2_X1    g20447(.A1(new_n23508_), .A2(new_n23201_), .Z(new_n23509_));
  NAND2_X1   g20448(.A1(new_n23380_), .A2(pi0625), .ZN(new_n23510_));
  AOI21_X1   g20449(.A1(new_n23198_), .A2(new_n12970_), .B(pi1153), .ZN(new_n23511_));
  NAND2_X1   g20450(.A1(new_n23510_), .A2(new_n23511_), .ZN(new_n23512_));
  NAND2_X1   g20451(.A1(new_n23296_), .A2(pi0625), .ZN(new_n23513_));
  INV_X1     g20452(.I(new_n23509_), .ZN(new_n23514_));
  NOR2_X1    g20453(.A1(new_n23514_), .A2(new_n12970_), .ZN(new_n23515_));
  INV_X1     g20454(.I(new_n23515_), .ZN(new_n23516_));
  NAND4_X1   g20455(.A1(new_n23516_), .A2(new_n12977_), .A3(new_n23513_), .A4(new_n23512_), .ZN(new_n23517_));
  AOI21_X1   g20456(.A1(new_n23196_), .A2(pi0625), .B(pi1153), .ZN(new_n23518_));
  NAND2_X1   g20457(.A1(new_n23510_), .A2(new_n23518_), .ZN(new_n23519_));
  NOR2_X1    g20458(.A1(new_n23296_), .A2(pi0625), .ZN(new_n23520_));
  NOR3_X1    g20459(.A1(new_n23520_), .A2(pi1153), .A3(new_n23515_), .ZN(new_n23521_));
  OAI21_X1   g20460(.A1(new_n23521_), .A2(new_n23519_), .B(new_n13657_), .ZN(new_n23522_));
  AOI21_X1   g20461(.A1(new_n23522_), .A2(new_n23517_), .B(new_n11891_), .ZN(new_n23523_));
  AOI21_X1   g20462(.A1(new_n11891_), .A2(new_n23509_), .B(new_n23523_), .ZN(new_n23524_));
  NAND2_X1   g20463(.A1(new_n23524_), .A2(new_n11870_), .ZN(new_n23525_));
  NOR2_X1    g20464(.A1(new_n11903_), .A2(pi1155), .ZN(new_n23526_));
  NAND2_X1   g20465(.A1(new_n23524_), .A2(new_n23526_), .ZN(new_n23527_));
  AOI21_X1   g20466(.A1(pi0660), .A2(new_n23295_), .B(new_n23527_), .ZN(new_n23528_));
  NAND2_X1   g20467(.A1(new_n23299_), .A2(new_n11923_), .ZN(new_n23529_));
  NOR2_X1    g20468(.A1(new_n23382_), .A2(new_n11903_), .ZN(new_n23530_));
  NOR2_X1    g20469(.A1(new_n23530_), .A2(pi1155), .ZN(new_n23531_));
  NAND2_X1   g20470(.A1(new_n23529_), .A2(new_n23531_), .ZN(new_n23532_));
  AOI21_X1   g20471(.A1(new_n23524_), .A2(new_n11903_), .B(new_n23532_), .ZN(new_n23533_));
  OAI21_X1   g20472(.A1(new_n23528_), .A2(new_n23533_), .B(pi0785), .ZN(new_n23534_));
  XOR2_X1    g20473(.A1(new_n23534_), .A2(new_n23525_), .Z(new_n23535_));
  INV_X1     g20474(.I(new_n23535_), .ZN(new_n23536_));
  NOR2_X1    g20475(.A1(new_n23536_), .A2(pi0781), .ZN(new_n23537_));
  INV_X1     g20476(.I(new_n23537_), .ZN(new_n23538_));
  NAND2_X1   g20477(.A1(new_n23301_), .A2(pi0618), .ZN(new_n23539_));
  NAND2_X1   g20478(.A1(new_n23196_), .A2(pi0618), .ZN(new_n23540_));
  NAND4_X1   g20479(.A1(new_n23539_), .A2(pi0627), .A3(new_n11950_), .A4(new_n23540_), .ZN(new_n23541_));
  NOR2_X1    g20480(.A1(new_n11934_), .A2(pi1154), .ZN(new_n23542_));
  AND2_X2    g20481(.A1(new_n23535_), .A2(new_n23542_), .Z(new_n23543_));
  NAND2_X1   g20482(.A1(new_n23535_), .A2(new_n11934_), .ZN(new_n23544_));
  AOI21_X1   g20483(.A1(new_n23198_), .A2(new_n11934_), .B(pi1154), .ZN(new_n23545_));
  NAND2_X1   g20484(.A1(new_n23539_), .A2(new_n23545_), .ZN(new_n23546_));
  NAND2_X1   g20485(.A1(new_n23546_), .A2(new_n11949_), .ZN(new_n23547_));
  AOI21_X1   g20486(.A1(new_n23383_), .A2(pi0618), .B(pi1154), .ZN(new_n23548_));
  NAND2_X1   g20487(.A1(new_n23547_), .A2(new_n23548_), .ZN(new_n23549_));
  INV_X1     g20488(.I(new_n23549_), .ZN(new_n23550_));
  AOI22_X1   g20489(.A1(new_n23543_), .A2(new_n23541_), .B1(new_n23544_), .B2(new_n23550_), .ZN(new_n23551_));
  NOR3_X1    g20490(.A1(new_n23551_), .A2(new_n11969_), .A3(new_n23538_), .ZN(new_n23552_));
  OAI21_X1   g20491(.A1(new_n23551_), .A2(new_n11969_), .B(new_n23538_), .ZN(new_n23553_));
  INV_X1     g20492(.I(new_n23553_), .ZN(new_n23554_));
  NOR2_X1    g20493(.A1(new_n23554_), .A2(new_n23552_), .ZN(new_n23555_));
  NOR2_X1    g20494(.A1(new_n11967_), .A2(pi1159), .ZN(new_n23556_));
  AND2_X2    g20495(.A1(new_n23555_), .A2(new_n23556_), .Z(new_n23557_));
  NAND2_X1   g20496(.A1(new_n23555_), .A2(new_n11967_), .ZN(new_n23558_));
  AOI21_X1   g20497(.A1(new_n23198_), .A2(new_n11967_), .B(pi1159), .ZN(new_n23559_));
  OAI21_X1   g20498(.A1(new_n23305_), .A2(new_n11967_), .B(new_n23559_), .ZN(new_n23560_));
  AOI21_X1   g20499(.A1(new_n23385_), .A2(pi0619), .B(pi1159), .ZN(new_n23561_));
  INV_X1     g20500(.I(new_n23561_), .ZN(new_n23562_));
  AOI21_X1   g20501(.A1(new_n23560_), .A2(new_n11966_), .B(new_n23562_), .ZN(new_n23563_));
  AOI22_X1   g20502(.A1(new_n23557_), .A2(new_n23409_), .B1(new_n23558_), .B2(new_n23563_), .ZN(new_n23564_));
  INV_X1     g20503(.I(new_n23555_), .ZN(new_n23565_));
  OAI21_X1   g20504(.A1(new_n23565_), .A2(new_n11999_), .B(new_n11985_), .ZN(new_n23566_));
  INV_X1     g20505(.I(new_n23307_), .ZN(new_n23567_));
  MUX2_X1    g20506(.I0(new_n23567_), .I1(new_n23198_), .S(new_n11994_), .Z(new_n23568_));
  NOR2_X1    g20507(.A1(new_n23568_), .A2(new_n17167_), .ZN(new_n23569_));
  OAI21_X1   g20508(.A1(new_n23567_), .A2(new_n23196_), .B(pi0626), .ZN(new_n23570_));
  OAI21_X1   g20509(.A1(new_n23384_), .A2(new_n23196_), .B(new_n12013_), .ZN(new_n23571_));
  OAI22_X1   g20510(.A1(new_n23570_), .A2(new_n17171_), .B1(new_n12020_), .B2(new_n23571_), .ZN(new_n23572_));
  NOR2_X1    g20511(.A1(new_n23569_), .A2(new_n23572_), .ZN(new_n23573_));
  OAI22_X1   g20512(.A1(new_n23564_), .A2(new_n23566_), .B1(new_n11986_), .B2(new_n23573_), .ZN(new_n23574_));
  OAI21_X1   g20513(.A1(new_n23405_), .A2(new_n14732_), .B(new_n14726_), .ZN(new_n23575_));
  AOI21_X1   g20514(.A1(new_n23574_), .A2(new_n23406_), .B(new_n23575_), .ZN(new_n23576_));
  OR2_X2     g20515(.A1(new_n23576_), .A2(new_n23401_), .Z(new_n23577_));
  NAND2_X1   g20516(.A1(new_n23198_), .A2(new_n12091_), .ZN(new_n23578_));
  OAI21_X1   g20517(.A1(new_n23309_), .A2(new_n12091_), .B(new_n23578_), .ZN(new_n23579_));
  MUX2_X1    g20518(.I0(new_n23579_), .I1(new_n23198_), .S(pi0644), .Z(new_n23580_));
  AOI21_X1   g20519(.A1(new_n23580_), .A2(pi0715), .B(pi1160), .ZN(new_n23581_));
  NAND2_X1   g20520(.A1(new_n12082_), .A2(pi0715), .ZN(new_n23584_));
  NOR4_X1    g20521(.A1(new_n23576_), .A2(new_n23401_), .A3(new_n23581_), .A4(new_n23584_), .ZN(new_n23585_));
  NOR4_X1    g20522(.A1(new_n23309_), .A2(pi0644), .A3(new_n12091_), .A4(new_n23198_), .ZN(new_n23586_));
  AOI21_X1   g20523(.A1(new_n12082_), .A2(new_n23198_), .B(new_n23579_), .ZN(new_n23587_));
  NOR4_X1    g20524(.A1(new_n23587_), .A2(pi0715), .A3(new_n12081_), .A4(new_n23586_), .ZN(new_n23588_));
  NOR2_X1    g20525(.A1(new_n12082_), .A2(pi0715), .ZN(new_n23589_));
  INV_X1     g20526(.I(new_n23589_), .ZN(new_n23590_));
  NOR4_X1    g20527(.A1(new_n23576_), .A2(new_n23401_), .A3(new_n23588_), .A4(new_n23590_), .ZN(new_n23591_));
  NOR2_X1    g20528(.A1(new_n23585_), .A2(new_n23591_), .ZN(new_n23592_));
  AOI21_X1   g20529(.A1(new_n23592_), .A2(pi0790), .B(new_n23577_), .ZN(new_n23593_));
  NAND3_X1   g20530(.A1(new_n23577_), .A2(pi0790), .A3(new_n23585_), .ZN(new_n23594_));
  NAND2_X1   g20531(.A1(new_n23594_), .A2(new_n6845_), .ZN(new_n23595_));
  OAI22_X1   g20532(.A1(new_n23595_), .A2(new_n23593_), .B1(new_n2601_), .B2(new_n6845_), .ZN(po0355));
  NAND2_X1   g20533(.A1(po1038), .A2(pi0199), .ZN(new_n23597_));
  INV_X1     g20534(.I(pi0637), .ZN(new_n23598_));
  MUX2_X1    g20535(.I0(new_n12391_), .I1(new_n12363_), .S(new_n6445_), .Z(new_n23599_));
  NOR2_X1    g20536(.A1(new_n23599_), .A2(new_n2566_), .ZN(new_n23600_));
  OAI21_X1   g20537(.A1(new_n5094_), .A2(new_n12430_), .B(new_n12423_), .ZN(new_n23601_));
  NAND3_X1   g20538(.A1(new_n23601_), .A2(new_n3285_), .A3(new_n13328_), .ZN(new_n23602_));
  AOI21_X1   g20539(.A1(new_n23602_), .A2(new_n13327_), .B(new_n23600_), .ZN(new_n23603_));
  NOR3_X1    g20540(.A1(new_n12438_), .A2(new_n6460_), .A3(new_n12391_), .ZN(new_n23604_));
  OAI21_X1   g20541(.A1(new_n23604_), .A2(new_n12394_), .B(pi0223), .ZN(new_n23605_));
  INV_X1     g20542(.I(new_n12436_), .ZN(new_n23606_));
  AOI21_X1   g20543(.A1(new_n23605_), .A2(new_n23606_), .B(new_n15651_), .ZN(new_n23607_));
  OAI21_X1   g20544(.A1(new_n23603_), .A2(new_n2587_), .B(new_n23607_), .ZN(new_n23608_));
  AOI21_X1   g20545(.A1(new_n23608_), .A2(new_n14342_), .B(pi0038), .ZN(new_n23609_));
  NAND2_X1   g20546(.A1(new_n23609_), .A2(pi0199), .ZN(new_n23610_));
  OAI21_X1   g20547(.A1(new_n14351_), .A2(new_n17581_), .B(new_n3231_), .ZN(new_n23611_));
  NAND2_X1   g20548(.A1(new_n23611_), .A2(new_n8094_), .ZN(new_n23612_));
  NOR2_X1    g20549(.A1(new_n14340_), .A2(pi0617), .ZN(new_n23613_));
  NAND3_X1   g20550(.A1(new_n23612_), .A2(new_n23610_), .A3(new_n23613_), .ZN(new_n23614_));
  INV_X1     g20551(.I(pi0617), .ZN(new_n23615_));
  NOR3_X1    g20552(.A1(new_n12121_), .A2(new_n3172_), .A3(new_n3154_), .ZN(new_n23616_));
  NOR2_X1    g20553(.A1(new_n12121_), .A2(new_n3154_), .ZN(new_n23617_));
  NOR3_X1    g20554(.A1(new_n12657_), .A2(new_n12664_), .A3(new_n12122_), .ZN(new_n23618_));
  AOI21_X1   g20555(.A1(new_n12602_), .A2(new_n13346_), .B(new_n12121_), .ZN(new_n23619_));
  NOR3_X1    g20556(.A1(new_n23619_), .A2(new_n23618_), .A3(pi0039), .ZN(new_n23620_));
  NOR3_X1    g20557(.A1(new_n23620_), .A2(pi0038), .A3(new_n23617_), .ZN(new_n23621_));
  OAI21_X1   g20558(.A1(new_n12343_), .A2(new_n12348_), .B(pi0039), .ZN(new_n23622_));
  NOR4_X1    g20559(.A1(new_n23621_), .A2(new_n8094_), .A3(new_n23616_), .A4(new_n23622_), .ZN(new_n23623_));
  OAI21_X1   g20560(.A1(new_n23623_), .A2(new_n23615_), .B(new_n3231_), .ZN(new_n23624_));
  NAND3_X1   g20561(.A1(new_n23614_), .A2(pi0199), .A3(new_n23624_), .ZN(new_n23625_));
  NOR2_X1    g20562(.A1(new_n23625_), .A2(new_n23598_), .ZN(new_n23626_));
  AOI21_X1   g20563(.A1(new_n12694_), .A2(new_n8094_), .B(pi0038), .ZN(new_n23627_));
  NAND2_X1   g20564(.A1(new_n13381_), .A2(pi0199), .ZN(new_n23628_));
  NAND2_X1   g20565(.A1(new_n14359_), .A2(new_n8094_), .ZN(new_n23629_));
  AOI21_X1   g20566(.A1(new_n23629_), .A2(new_n14364_), .B(new_n3232_), .ZN(new_n23630_));
  OAI21_X1   g20567(.A1(new_n23628_), .A2(new_n23627_), .B(new_n23630_), .ZN(new_n23631_));
  NAND4_X1   g20568(.A1(new_n23631_), .A2(new_n8094_), .A3(new_n23615_), .A4(new_n3231_), .ZN(new_n23632_));
  NAND2_X1   g20569(.A1(new_n14396_), .A2(pi0199), .ZN(new_n23633_));
  NAND2_X1   g20570(.A1(new_n23633_), .A2(new_n23615_), .ZN(new_n23634_));
  NAND2_X1   g20571(.A1(new_n23634_), .A2(new_n23632_), .ZN(new_n23635_));
  AOI21_X1   g20572(.A1(new_n23598_), .A2(new_n23635_), .B(new_n23626_), .ZN(new_n23636_));
  AOI21_X1   g20573(.A1(new_n23635_), .A2(pi0625), .B(pi1153), .ZN(new_n23637_));
  NAND3_X1   g20574(.A1(new_n13356_), .A2(new_n13359_), .A3(new_n3154_), .ZN(new_n23638_));
  NAND3_X1   g20575(.A1(new_n13336_), .A2(new_n13335_), .A3(pi0039), .ZN(new_n23639_));
  NAND3_X1   g20576(.A1(new_n23638_), .A2(new_n23639_), .A3(new_n3172_), .ZN(new_n23640_));
  AOI21_X1   g20577(.A1(new_n23640_), .A2(new_n14352_), .B(new_n3232_), .ZN(new_n23641_));
  OAI21_X1   g20578(.A1(new_n23641_), .A2(pi0199), .B(new_n23613_), .ZN(new_n23642_));
  AOI21_X1   g20579(.A1(pi0199), .A2(new_n23609_), .B(new_n23642_), .ZN(new_n23643_));
  NAND2_X1   g20580(.A1(new_n23624_), .A2(pi0199), .ZN(new_n23644_));
  NOR2_X1    g20581(.A1(new_n23643_), .A2(new_n23644_), .ZN(new_n23645_));
  AND2_X2    g20582(.A1(new_n23634_), .A2(new_n23632_), .Z(new_n23646_));
  NAND3_X1   g20583(.A1(new_n23646_), .A2(new_n23645_), .A3(new_n23598_), .ZN(new_n23647_));
  AOI21_X1   g20584(.A1(new_n23598_), .A2(new_n23635_), .B(new_n23645_), .ZN(new_n23648_));
  NOR2_X1    g20585(.A1(new_n23648_), .A2(pi0625), .ZN(new_n23649_));
  AOI21_X1   g20586(.A1(new_n23649_), .A2(new_n23647_), .B(new_n23637_), .ZN(new_n23650_));
  MUX2_X1    g20587(.I0(new_n23635_), .I1(new_n23625_), .S(new_n23598_), .Z(new_n23651_));
  AOI21_X1   g20588(.A1(new_n23635_), .A2(new_n12970_), .B(new_n11893_), .ZN(new_n23652_));
  NOR2_X1    g20589(.A1(new_n12965_), .A2(new_n8094_), .ZN(new_n23653_));
  NOR3_X1    g20590(.A1(new_n13368_), .A2(pi0199), .A3(new_n11885_), .ZN(new_n23654_));
  AOI21_X1   g20591(.A1(new_n12828_), .A2(new_n11885_), .B(new_n8094_), .ZN(new_n23655_));
  OAI21_X1   g20592(.A1(new_n23654_), .A2(new_n23655_), .B(pi0038), .ZN(new_n23656_));
  OAI21_X1   g20593(.A1(new_n12937_), .A2(new_n12954_), .B(pi0199), .ZN(new_n23657_));
  NOR2_X1    g20594(.A1(new_n23657_), .A2(new_n3154_), .ZN(new_n23658_));
  NAND3_X1   g20595(.A1(new_n12643_), .A2(new_n12602_), .A3(new_n8094_), .ZN(new_n23659_));
  OAI21_X1   g20596(.A1(new_n12643_), .A2(pi0199), .B(new_n12657_), .ZN(new_n23660_));
  NAND3_X1   g20597(.A1(new_n23660_), .A2(new_n23659_), .A3(new_n2544_), .ZN(new_n23661_));
  OAI21_X1   g20598(.A1(new_n23658_), .A2(new_n23661_), .B(new_n23656_), .ZN(new_n23662_));
  NOR4_X1    g20599(.A1(new_n23662_), .A2(pi0199), .A3(pi0637), .A4(new_n3232_), .ZN(new_n23663_));
  NOR2_X1    g20600(.A1(new_n23653_), .A2(pi0637), .ZN(new_n23664_));
  NOR2_X1    g20601(.A1(new_n23664_), .A2(new_n23663_), .ZN(new_n23665_));
  NOR4_X1    g20602(.A1(new_n23665_), .A2(pi0625), .A3(pi1153), .A4(new_n23653_), .ZN(new_n23666_));
  NOR4_X1    g20603(.A1(new_n23651_), .A2(new_n20722_), .A3(new_n23652_), .A4(new_n23666_), .ZN(new_n23667_));
  OAI21_X1   g20604(.A1(new_n23653_), .A2(pi0625), .B(pi1153), .ZN(new_n23668_));
  NOR2_X1    g20605(.A1(new_n23665_), .A2(new_n12970_), .ZN(new_n23669_));
  AOI21_X1   g20606(.A1(new_n23669_), .A2(new_n23668_), .B(pi0608), .ZN(new_n23670_));
  INV_X1     g20607(.I(new_n23670_), .ZN(new_n23671_));
  NOR3_X1    g20608(.A1(new_n23650_), .A2(new_n23667_), .A3(new_n23671_), .ZN(new_n23672_));
  MUX2_X1    g20609(.I0(new_n23672_), .I1(new_n23636_), .S(new_n11891_), .Z(new_n23673_));
  NAND2_X1   g20610(.A1(new_n23673_), .A2(new_n11870_), .ZN(new_n23674_));
  AOI21_X1   g20611(.A1(new_n23668_), .A2(new_n23669_), .B(new_n23666_), .ZN(new_n23675_));
  NOR3_X1    g20612(.A1(new_n23675_), .A2(new_n11891_), .A3(new_n23665_), .ZN(new_n23676_));
  INV_X1     g20613(.I(new_n23665_), .ZN(new_n23677_));
  AOI21_X1   g20614(.A1(new_n23675_), .A2(pi0778), .B(new_n23677_), .ZN(new_n23678_));
  OAI21_X1   g20615(.A1(new_n23676_), .A2(new_n23678_), .B(new_n11903_), .ZN(new_n23679_));
  NAND3_X1   g20616(.A1(new_n23634_), .A2(new_n11924_), .A3(new_n23632_), .ZN(new_n23680_));
  NAND2_X1   g20617(.A1(new_n23653_), .A2(new_n11914_), .ZN(new_n23681_));
  NAND2_X1   g20618(.A1(new_n23680_), .A2(new_n23681_), .ZN(new_n23682_));
  NOR3_X1    g20619(.A1(new_n23682_), .A2(new_n11903_), .A3(new_n23633_), .ZN(new_n23683_));
  AOI22_X1   g20620(.A1(new_n23680_), .A2(new_n23681_), .B1(pi0609), .B2(new_n23633_), .ZN(new_n23684_));
  OAI21_X1   g20621(.A1(new_n23683_), .A2(new_n23684_), .B(new_n11912_), .ZN(new_n23685_));
  NAND2_X1   g20622(.A1(new_n23685_), .A2(pi0660), .ZN(new_n23686_));
  NAND2_X1   g20623(.A1(new_n23686_), .A2(pi0609), .ZN(new_n23687_));
  AOI21_X1   g20624(.A1(pi1155), .A2(new_n23679_), .B(new_n23687_), .ZN(new_n23688_));
  INV_X1     g20625(.I(new_n23637_), .ZN(new_n23689_));
  OAI21_X1   g20626(.A1(new_n23646_), .A2(pi0637), .B(new_n23625_), .ZN(new_n23690_));
  NAND3_X1   g20627(.A1(new_n23690_), .A2(new_n23647_), .A3(new_n12970_), .ZN(new_n23691_));
  NAND2_X1   g20628(.A1(new_n23691_), .A2(new_n23689_), .ZN(new_n23692_));
  INV_X1     g20629(.I(new_n23651_), .ZN(new_n23693_));
  NOR3_X1    g20630(.A1(new_n23666_), .A2(new_n20722_), .A3(new_n23652_), .ZN(new_n23694_));
  NAND2_X1   g20631(.A1(new_n23693_), .A2(new_n23694_), .ZN(new_n23695_));
  NAND3_X1   g20632(.A1(new_n23692_), .A2(new_n23695_), .A3(new_n23670_), .ZN(new_n23696_));
  NAND3_X1   g20633(.A1(new_n23696_), .A2(pi0778), .A3(new_n23636_), .ZN(new_n23697_));
  INV_X1     g20634(.I(new_n23636_), .ZN(new_n23698_));
  OAI21_X1   g20635(.A1(new_n23696_), .A2(new_n11891_), .B(new_n23698_), .ZN(new_n23699_));
  NAND3_X1   g20636(.A1(new_n23699_), .A2(new_n23697_), .A3(new_n11903_), .ZN(new_n23700_));
  NOR2_X1    g20637(.A1(new_n23676_), .A2(new_n23678_), .ZN(new_n23701_));
  NOR2_X1    g20638(.A1(new_n11923_), .A2(pi1155), .ZN(new_n23704_));
  OAI21_X1   g20639(.A1(new_n23701_), .A2(new_n11903_), .B(new_n23704_), .ZN(new_n23705_));
  INV_X1     g20640(.I(new_n23705_), .ZN(new_n23706_));
  AOI22_X1   g20641(.A1(new_n23700_), .A2(new_n23706_), .B1(new_n23673_), .B2(new_n23688_), .ZN(new_n23707_));
  NOR3_X1    g20642(.A1(new_n23707_), .A2(new_n11870_), .A3(new_n23674_), .ZN(new_n23708_));
  NAND2_X1   g20643(.A1(new_n23699_), .A2(new_n23697_), .ZN(new_n23709_));
  NOR2_X1    g20644(.A1(new_n23709_), .A2(pi0785), .ZN(new_n23710_));
  INV_X1     g20645(.I(new_n23688_), .ZN(new_n23711_));
  NOR3_X1    g20646(.A1(new_n23672_), .A2(new_n11891_), .A3(new_n23698_), .ZN(new_n23712_));
  AOI21_X1   g20647(.A1(new_n23672_), .A2(pi0778), .B(new_n23636_), .ZN(new_n23713_));
  NOR3_X1    g20648(.A1(new_n23712_), .A2(new_n23713_), .A3(pi0609), .ZN(new_n23714_));
  OAI22_X1   g20649(.A1(new_n23714_), .A2(new_n23705_), .B1(new_n23711_), .B2(new_n23709_), .ZN(new_n23715_));
  AOI21_X1   g20650(.A1(new_n23715_), .A2(pi0785), .B(new_n23710_), .ZN(new_n23716_));
  NOR3_X1    g20651(.A1(new_n23716_), .A2(new_n23708_), .A3(pi0781), .ZN(new_n23717_));
  INV_X1     g20652(.I(new_n23717_), .ZN(new_n23718_));
  NAND3_X1   g20653(.A1(new_n23682_), .A2(pi0609), .A3(new_n23633_), .ZN(new_n23719_));
  OAI21_X1   g20654(.A1(new_n23682_), .A2(new_n11903_), .B(new_n23653_), .ZN(new_n23720_));
  AND2_X2    g20655(.A1(new_n23720_), .A2(new_n23719_), .Z(new_n23721_));
  OAI21_X1   g20656(.A1(new_n23721_), .A2(new_n11912_), .B(new_n23685_), .ZN(new_n23722_));
  MUX2_X1    g20657(.I0(new_n23722_), .I1(new_n23682_), .S(new_n11870_), .Z(new_n23723_));
  NAND3_X1   g20658(.A1(new_n23723_), .A2(new_n11934_), .A3(new_n23653_), .ZN(new_n23724_));
  OAI21_X1   g20659(.A1(new_n23723_), .A2(pi0618), .B(new_n23633_), .ZN(new_n23725_));
  NAND4_X1   g20660(.A1(new_n23725_), .A2(new_n23724_), .A3(pi0627), .A4(new_n11950_), .ZN(new_n23726_));
  NOR2_X1    g20661(.A1(new_n23633_), .A2(new_n11938_), .ZN(new_n23727_));
  AOI21_X1   g20662(.A1(new_n23701_), .A2(new_n11938_), .B(new_n23727_), .ZN(new_n23728_));
  NOR4_X1    g20663(.A1(new_n23716_), .A2(new_n23708_), .A3(new_n11934_), .A4(pi1154), .ZN(new_n23729_));
  NAND3_X1   g20664(.A1(new_n23715_), .A2(pi0785), .A3(new_n23710_), .ZN(new_n23730_));
  OAI21_X1   g20665(.A1(new_n23707_), .A2(new_n11870_), .B(new_n23674_), .ZN(new_n23731_));
  NAND3_X1   g20666(.A1(new_n23730_), .A2(new_n23731_), .A3(new_n11934_), .ZN(new_n23732_));
  AOI21_X1   g20667(.A1(new_n23728_), .A2(pi0618), .B(new_n14687_), .ZN(new_n23733_));
  AOI22_X1   g20668(.A1(new_n23729_), .A2(new_n23726_), .B1(new_n23732_), .B2(new_n23733_), .ZN(new_n23734_));
  NOR3_X1    g20669(.A1(new_n23734_), .A2(new_n11969_), .A3(new_n23718_), .ZN(new_n23735_));
  NOR2_X1    g20670(.A1(new_n11934_), .A2(pi1154), .ZN(new_n23736_));
  NAND4_X1   g20671(.A1(new_n23730_), .A2(new_n23731_), .A3(new_n23726_), .A4(new_n23736_), .ZN(new_n23737_));
  NOR3_X1    g20672(.A1(new_n23716_), .A2(new_n23708_), .A3(pi0618), .ZN(new_n23738_));
  INV_X1     g20673(.I(new_n23733_), .ZN(new_n23739_));
  OAI21_X1   g20674(.A1(new_n23738_), .A2(new_n23739_), .B(new_n23737_), .ZN(new_n23740_));
  AOI21_X1   g20675(.A1(new_n23740_), .A2(pi0781), .B(new_n23717_), .ZN(new_n23741_));
  NOR2_X1    g20676(.A1(new_n23735_), .A2(new_n23741_), .ZN(new_n23742_));
  INV_X1     g20677(.I(new_n23682_), .ZN(new_n23743_));
  INV_X1     g20678(.I(new_n23685_), .ZN(new_n23744_));
  AOI21_X1   g20679(.A1(new_n23720_), .A2(new_n23719_), .B(new_n11912_), .ZN(new_n23745_));
  NOR2_X1    g20680(.A1(new_n23744_), .A2(new_n23745_), .ZN(new_n23746_));
  MUX2_X1    g20681(.I0(new_n23746_), .I1(new_n23743_), .S(new_n11870_), .Z(new_n23747_));
  NOR3_X1    g20682(.A1(new_n23747_), .A2(pi0618), .A3(new_n23633_), .ZN(new_n23748_));
  AOI21_X1   g20683(.A1(new_n23747_), .A2(new_n11934_), .B(new_n23653_), .ZN(new_n23749_));
  NOR3_X1    g20684(.A1(new_n23748_), .A2(new_n23749_), .A3(pi1154), .ZN(new_n23750_));
  MUX2_X1    g20685(.I0(new_n23750_), .I1(new_n23723_), .S(new_n11969_), .Z(new_n23751_));
  NAND3_X1   g20686(.A1(new_n23751_), .A2(new_n11967_), .A3(new_n23653_), .ZN(new_n23752_));
  OAI21_X1   g20687(.A1(new_n23751_), .A2(pi0619), .B(new_n23633_), .ZN(new_n23753_));
  NAND3_X1   g20688(.A1(new_n23753_), .A2(new_n23752_), .A3(new_n11869_), .ZN(new_n23754_));
  NOR2_X1    g20689(.A1(new_n23754_), .A2(new_n11966_), .ZN(new_n23755_));
  NAND3_X1   g20690(.A1(new_n23740_), .A2(pi0781), .A3(new_n23717_), .ZN(new_n23756_));
  OAI21_X1   g20691(.A1(new_n23734_), .A2(new_n11969_), .B(new_n23718_), .ZN(new_n23757_));
  NOR2_X1    g20692(.A1(new_n23653_), .A2(new_n11961_), .ZN(new_n23758_));
  AOI21_X1   g20693(.A1(new_n23728_), .A2(new_n11961_), .B(new_n23758_), .ZN(new_n23759_));
  NOR2_X1    g20694(.A1(new_n11967_), .A2(pi1159), .ZN(new_n23760_));
  NAND3_X1   g20695(.A1(new_n23757_), .A2(new_n23756_), .A3(new_n23760_), .ZN(new_n23761_));
  NOR3_X1    g20696(.A1(new_n23735_), .A2(new_n23741_), .A3(pi0619), .ZN(new_n23762_));
  INV_X1     g20697(.I(new_n23759_), .ZN(new_n23763_));
  AOI21_X1   g20698(.A1(new_n23763_), .A2(pi0619), .B(new_n14904_), .ZN(new_n23764_));
  INV_X1     g20699(.I(new_n23764_), .ZN(new_n23765_));
  OAI22_X1   g20700(.A1(new_n23762_), .A2(new_n23765_), .B1(new_n23761_), .B2(new_n23755_), .ZN(new_n23766_));
  MUX2_X1    g20701(.I0(new_n23766_), .I1(new_n23742_), .S(new_n11985_), .Z(new_n23767_));
  NOR3_X1    g20702(.A1(new_n23735_), .A2(new_n23741_), .A3(pi0789), .ZN(new_n23768_));
  NAND3_X1   g20703(.A1(new_n23766_), .A2(pi0789), .A3(new_n23768_), .ZN(new_n23769_));
  INV_X1     g20704(.I(new_n23768_), .ZN(new_n23770_));
  NAND3_X1   g20705(.A1(new_n23725_), .A2(new_n23724_), .A3(new_n11950_), .ZN(new_n23771_));
  MUX2_X1    g20706(.I0(new_n23771_), .I1(new_n23747_), .S(new_n11969_), .Z(new_n23772_));
  NOR3_X1    g20707(.A1(new_n23772_), .A2(pi0619), .A3(new_n23633_), .ZN(new_n23773_));
  AOI21_X1   g20708(.A1(new_n23772_), .A2(new_n11967_), .B(new_n23653_), .ZN(new_n23774_));
  NOR3_X1    g20709(.A1(new_n23773_), .A2(new_n23774_), .A3(pi1159), .ZN(new_n23775_));
  NAND2_X1   g20710(.A1(new_n23775_), .A2(pi0648), .ZN(new_n23776_));
  NOR4_X1    g20711(.A1(new_n23735_), .A2(new_n23741_), .A3(new_n11967_), .A4(pi1159), .ZN(new_n23777_));
  NAND3_X1   g20712(.A1(new_n23757_), .A2(new_n23756_), .A3(new_n11967_), .ZN(new_n23778_));
  AOI22_X1   g20713(.A1(new_n23777_), .A2(new_n23776_), .B1(new_n23778_), .B2(new_n23764_), .ZN(new_n23779_));
  OAI21_X1   g20714(.A1(new_n23779_), .A2(new_n11985_), .B(new_n23770_), .ZN(new_n23780_));
  MUX2_X1    g20715(.I0(new_n23754_), .I1(new_n23772_), .S(new_n11985_), .Z(new_n23781_));
  NOR3_X1    g20716(.A1(new_n11994_), .A2(new_n11989_), .A3(pi1158), .ZN(new_n23782_));
  NOR2_X1    g20717(.A1(new_n23633_), .A2(new_n12014_), .ZN(new_n23783_));
  AOI21_X1   g20718(.A1(new_n23759_), .A2(new_n12014_), .B(new_n23783_), .ZN(new_n23784_));
  NOR2_X1    g20719(.A1(new_n11994_), .A2(pi0641), .ZN(new_n23785_));
  INV_X1     g20720(.I(new_n23785_), .ZN(new_n23786_));
  AOI21_X1   g20721(.A1(new_n23781_), .A2(new_n23782_), .B(new_n23786_), .ZN(new_n23787_));
  INV_X1     g20722(.I(new_n23787_), .ZN(new_n23788_));
  AOI21_X1   g20723(.A1(new_n23780_), .A2(new_n23769_), .B(new_n23788_), .ZN(new_n23789_));
  NAND2_X1   g20724(.A1(new_n23781_), .A2(new_n11994_), .ZN(new_n23790_));
  AOI21_X1   g20725(.A1(new_n23653_), .A2(pi0626), .B(new_n11989_), .ZN(new_n23791_));
  NOR3_X1    g20726(.A1(new_n11989_), .A2(pi0626), .A3(pi1158), .ZN(new_n23792_));
  INV_X1     g20727(.I(new_n23792_), .ZN(new_n23793_));
  AOI21_X1   g20728(.A1(new_n23790_), .A2(new_n23791_), .B(new_n23793_), .ZN(new_n23794_));
  NAND3_X1   g20729(.A1(new_n23789_), .A2(pi0788), .A3(new_n23767_), .ZN(new_n23795_));
  NAND2_X1   g20730(.A1(new_n23780_), .A2(new_n23769_), .ZN(new_n23796_));
  MUX2_X1    g20731(.I0(new_n23775_), .I1(new_n23751_), .S(new_n11985_), .Z(new_n23797_));
  NOR2_X1    g20732(.A1(new_n23797_), .A2(pi0626), .ZN(new_n23798_));
  INV_X1     g20733(.I(new_n23791_), .ZN(new_n23799_));
  OAI21_X1   g20734(.A1(new_n23798_), .A2(new_n23799_), .B(new_n23792_), .ZN(new_n23800_));
  AOI22_X1   g20735(.A1(new_n23780_), .A2(new_n23769_), .B1(new_n23788_), .B2(new_n23800_), .ZN(new_n23801_));
  OAI21_X1   g20736(.A1(new_n23801_), .A2(new_n11986_), .B(new_n23796_), .ZN(new_n23802_));
  NAND2_X1   g20737(.A1(new_n23802_), .A2(new_n23795_), .ZN(new_n23803_));
  NOR3_X1    g20738(.A1(new_n23779_), .A2(new_n11985_), .A3(new_n23770_), .ZN(new_n23804_));
  AOI21_X1   g20739(.A1(new_n23766_), .A2(pi0789), .B(new_n23768_), .ZN(new_n23805_));
  OAI22_X1   g20740(.A1(new_n23804_), .A2(new_n23805_), .B1(new_n23794_), .B2(new_n23787_), .ZN(new_n23806_));
  NOR3_X1    g20741(.A1(new_n23806_), .A2(new_n11986_), .A3(new_n23796_), .ZN(new_n23807_));
  AOI21_X1   g20742(.A1(new_n23806_), .A2(pi0788), .B(new_n23767_), .ZN(new_n23808_));
  NOR2_X1    g20743(.A1(new_n23653_), .A2(new_n14624_), .ZN(new_n23809_));
  AOI21_X1   g20744(.A1(new_n23797_), .A2(new_n14624_), .B(new_n23809_), .ZN(new_n23810_));
  OR2_X2     g20745(.A1(new_n23810_), .A2(pi0628), .Z(new_n23811_));
  NAND2_X1   g20746(.A1(new_n23784_), .A2(new_n13114_), .ZN(new_n23812_));
  OAI21_X1   g20747(.A1(new_n13114_), .A2(new_n23653_), .B(new_n23812_), .ZN(new_n23813_));
  NAND3_X1   g20748(.A1(new_n23813_), .A2(new_n12031_), .A3(new_n23653_), .ZN(new_n23814_));
  OAI21_X1   g20749(.A1(new_n23813_), .A2(pi0628), .B(new_n23633_), .ZN(new_n23815_));
  AND3_X2    g20750(.A1(new_n23815_), .A2(new_n23814_), .A3(new_n12026_), .Z(new_n23816_));
  AOI21_X1   g20751(.A1(new_n23816_), .A2(pi0629), .B(new_n12031_), .ZN(new_n23817_));
  INV_X1     g20752(.I(new_n23817_), .ZN(new_n23818_));
  AOI21_X1   g20753(.A1(new_n23811_), .A2(pi1156), .B(new_n23818_), .ZN(new_n23819_));
  OAI21_X1   g20754(.A1(new_n23807_), .A2(new_n23808_), .B(new_n23819_), .ZN(new_n23820_));
  NOR3_X1    g20755(.A1(new_n12030_), .A2(new_n12026_), .A3(pi0628), .ZN(new_n23821_));
  NOR3_X1    g20756(.A1(new_n23820_), .A2(new_n11868_), .A3(new_n23803_), .ZN(new_n23822_));
  NOR2_X1    g20757(.A1(new_n23807_), .A2(new_n23808_), .ZN(new_n23823_));
  OAI22_X1   g20758(.A1(new_n23807_), .A2(new_n23808_), .B1(new_n23819_), .B2(new_n23821_), .ZN(new_n23824_));
  AOI21_X1   g20759(.A1(new_n23824_), .A2(pi0792), .B(new_n23823_), .ZN(new_n23825_));
  NOR3_X1    g20760(.A1(new_n23825_), .A2(new_n23822_), .A3(pi0787), .ZN(new_n23826_));
  NAND2_X1   g20761(.A1(new_n23811_), .A2(pi1156), .ZN(new_n23827_));
  NAND2_X1   g20762(.A1(new_n23827_), .A2(new_n23817_), .ZN(new_n23828_));
  AOI21_X1   g20763(.A1(new_n23802_), .A2(new_n23795_), .B(new_n23828_), .ZN(new_n23829_));
  NAND3_X1   g20764(.A1(new_n23823_), .A2(new_n23829_), .A3(pi0792), .ZN(new_n23830_));
  INV_X1     g20765(.I(new_n23821_), .ZN(new_n23831_));
  AOI22_X1   g20766(.A1(new_n23802_), .A2(new_n23795_), .B1(new_n23828_), .B2(new_n23831_), .ZN(new_n23832_));
  OAI21_X1   g20767(.A1(new_n23832_), .A2(new_n11868_), .B(new_n23803_), .ZN(new_n23833_));
  NAND2_X1   g20768(.A1(new_n23633_), .A2(new_n12053_), .ZN(new_n23834_));
  OAI21_X1   g20769(.A1(new_n23810_), .A2(new_n12053_), .B(new_n23834_), .ZN(new_n23835_));
  AOI21_X1   g20770(.A1(new_n23835_), .A2(new_n12061_), .B(new_n12049_), .ZN(new_n23836_));
  MUX2_X1    g20771(.I0(new_n23816_), .I1(new_n23813_), .S(new_n11868_), .Z(new_n23837_));
  NAND3_X1   g20772(.A1(new_n23837_), .A2(new_n12061_), .A3(new_n23653_), .ZN(new_n23838_));
  OAI21_X1   g20773(.A1(new_n23837_), .A2(pi0647), .B(new_n23633_), .ZN(new_n23839_));
  NAND3_X1   g20774(.A1(new_n23839_), .A2(new_n23838_), .A3(new_n12049_), .ZN(new_n23840_));
  OAI21_X1   g20775(.A1(new_n23840_), .A2(new_n12060_), .B(pi0647), .ZN(new_n23841_));
  NOR2_X1    g20776(.A1(new_n23841_), .A2(new_n23836_), .ZN(new_n23842_));
  NAND3_X1   g20777(.A1(new_n23833_), .A2(new_n23830_), .A3(new_n23842_), .ZN(new_n23843_));
  NOR3_X1    g20778(.A1(new_n23825_), .A2(new_n23822_), .A3(pi0647), .ZN(new_n23844_));
  AOI21_X1   g20779(.A1(new_n23835_), .A2(pi0647), .B(new_n13743_), .ZN(new_n23845_));
  INV_X1     g20780(.I(new_n23845_), .ZN(new_n23846_));
  OAI21_X1   g20781(.A1(new_n23844_), .A2(new_n23846_), .B(new_n23843_), .ZN(new_n23847_));
  NAND3_X1   g20782(.A1(new_n23847_), .A2(pi0787), .A3(new_n23826_), .ZN(new_n23848_));
  INV_X1     g20783(.I(new_n23826_), .ZN(new_n23849_));
  NOR2_X1    g20784(.A1(new_n23825_), .A2(new_n23822_), .ZN(new_n23850_));
  NAND3_X1   g20785(.A1(new_n23833_), .A2(new_n23830_), .A3(new_n12061_), .ZN(new_n23851_));
  AOI22_X1   g20786(.A1(new_n23851_), .A2(new_n23845_), .B1(new_n23850_), .B2(new_n23842_), .ZN(new_n23852_));
  OAI21_X1   g20787(.A1(new_n23852_), .A2(new_n12048_), .B(new_n23849_), .ZN(new_n23853_));
  NAND2_X1   g20788(.A1(new_n23853_), .A2(new_n23848_), .ZN(new_n23854_));
  NOR2_X1    g20789(.A1(new_n23854_), .A2(pi0790), .ZN(new_n23855_));
  NOR3_X1    g20790(.A1(new_n23852_), .A2(new_n12048_), .A3(new_n23849_), .ZN(new_n23856_));
  AOI21_X1   g20791(.A1(new_n23847_), .A2(pi0787), .B(new_n23826_), .ZN(new_n23857_));
  NOR3_X1    g20792(.A1(new_n23856_), .A2(new_n23857_), .A3(pi0644), .ZN(new_n23858_));
  NOR2_X1    g20793(.A1(new_n23633_), .A2(new_n12092_), .ZN(new_n23859_));
  NOR2_X1    g20794(.A1(new_n23835_), .A2(new_n12091_), .ZN(new_n23860_));
  NOR3_X1    g20795(.A1(new_n23860_), .A2(pi0644), .A3(new_n23859_), .ZN(new_n23861_));
  OAI21_X1   g20796(.A1(new_n23653_), .A2(new_n12082_), .B(pi0715), .ZN(new_n23862_));
  NOR2_X1    g20797(.A1(new_n23837_), .A2(pi0787), .ZN(new_n23863_));
  NAND2_X1   g20798(.A1(new_n23840_), .A2(pi0787), .ZN(new_n23864_));
  XOR2_X1    g20799(.A1(new_n23864_), .A2(new_n23863_), .Z(new_n23865_));
  AOI21_X1   g20800(.A1(new_n23865_), .A2(pi0644), .B(new_n13169_), .ZN(new_n23866_));
  OAI21_X1   g20801(.A1(new_n23861_), .A2(new_n23862_), .B(new_n23866_), .ZN(new_n23867_));
  NOR2_X1    g20802(.A1(new_n23860_), .A2(new_n23859_), .ZN(new_n23868_));
  NOR3_X1    g20803(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n23869_));
  NOR2_X1    g20804(.A1(new_n12082_), .A2(pi0715), .ZN(new_n23871_));
  INV_X1     g20805(.I(new_n23871_), .ZN(new_n23872_));
  AOI21_X1   g20806(.A1(new_n23868_), .A2(new_n23869_), .B(new_n23872_), .ZN(new_n23873_));
  INV_X1     g20807(.I(new_n23873_), .ZN(new_n23874_));
  OAI22_X1   g20808(.A1(new_n23858_), .A2(new_n23867_), .B1(new_n23854_), .B2(new_n23874_), .ZN(new_n23875_));
  AOI21_X1   g20809(.A1(new_n23875_), .A2(pi0790), .B(new_n23855_), .ZN(new_n23876_));
  INV_X1     g20810(.I(new_n23855_), .ZN(new_n23877_));
  MUX2_X1    g20811(.I0(new_n23847_), .I1(new_n23850_), .S(new_n12048_), .Z(new_n23878_));
  AOI21_X1   g20812(.A1(new_n23878_), .A2(new_n12082_), .B(new_n23867_), .ZN(new_n23879_));
  NOR3_X1    g20813(.A1(new_n23856_), .A2(new_n23857_), .A3(new_n23874_), .ZN(new_n23880_));
  OAI21_X1   g20814(.A1(new_n23879_), .A2(new_n23880_), .B(pi0790), .ZN(new_n23881_));
  OAI21_X1   g20815(.A1(new_n23881_), .A2(new_n23877_), .B(new_n6845_), .ZN(new_n23882_));
  OAI21_X1   g20816(.A1(new_n23882_), .A2(new_n23876_), .B(new_n23597_), .ZN(po0356));
  NOR2_X1    g20817(.A1(new_n12965_), .A2(new_n8098_), .ZN(new_n23884_));
  NOR2_X1    g20818(.A1(new_n23884_), .A2(new_n13114_), .ZN(new_n23885_));
  INV_X1     g20819(.I(new_n23884_), .ZN(new_n23886_));
  NOR2_X1    g20820(.A1(new_n23886_), .A2(new_n12014_), .ZN(new_n23887_));
  NAND2_X1   g20821(.A1(new_n23884_), .A2(new_n13024_), .ZN(new_n23888_));
  NOR3_X1    g20822(.A1(new_n13368_), .A2(pi0200), .A3(new_n11885_), .ZN(new_n23889_));
  AOI21_X1   g20823(.A1(new_n12828_), .A2(new_n11885_), .B(new_n8098_), .ZN(new_n23890_));
  OAI21_X1   g20824(.A1(new_n23889_), .A2(new_n23890_), .B(pi0038), .ZN(new_n23891_));
  NOR4_X1    g20825(.A1(new_n12936_), .A2(new_n8098_), .A3(pi0299), .A4(new_n12952_), .ZN(new_n23892_));
  NAND2_X1   g20826(.A1(new_n12930_), .A2(pi0200), .ZN(new_n23893_));
  AOI21_X1   g20827(.A1(new_n12950_), .A2(pi0200), .B(pi0299), .ZN(new_n23894_));
  NAND2_X1   g20828(.A1(new_n23893_), .A2(new_n23894_), .ZN(new_n23895_));
  OAI21_X1   g20829(.A1(new_n23895_), .A2(new_n23892_), .B(pi0039), .ZN(new_n23896_));
  NOR2_X1    g20830(.A1(new_n3154_), .A2(new_n8098_), .ZN(new_n23897_));
  AOI21_X1   g20831(.A1(new_n12602_), .A2(new_n23897_), .B(pi0038), .ZN(new_n23898_));
  NAND2_X1   g20832(.A1(new_n23896_), .A2(new_n23898_), .ZN(new_n23899_));
  AOI21_X1   g20833(.A1(new_n23899_), .A2(new_n23891_), .B(new_n3232_), .ZN(new_n23900_));
  INV_X1     g20834(.I(pi0643), .ZN(new_n23901_));
  NAND3_X1   g20835(.A1(new_n3231_), .A2(new_n8098_), .A3(new_n23901_), .ZN(new_n23902_));
  OAI22_X1   g20836(.A1(new_n23884_), .A2(pi0643), .B1(new_n23900_), .B2(new_n23902_), .ZN(new_n23903_));
  INV_X1     g20837(.I(new_n23903_), .ZN(new_n23904_));
  XOR2_X1    g20838(.A1(new_n23903_), .A2(new_n23886_), .Z(new_n23905_));
  NAND2_X1   g20839(.A1(new_n23905_), .A2(pi0625), .ZN(new_n23906_));
  NOR2_X1    g20840(.A1(new_n23906_), .A2(new_n23904_), .ZN(new_n23907_));
  AOI21_X1   g20841(.A1(pi0625), .A2(new_n23886_), .B(new_n23903_), .ZN(new_n23908_));
  OAI21_X1   g20842(.A1(new_n23908_), .A2(new_n23907_), .B(new_n11893_), .ZN(new_n23909_));
  XOR2_X1    g20843(.A1(new_n23906_), .A2(new_n23884_), .Z(new_n23910_));
  OAI21_X1   g20844(.A1(new_n23910_), .A2(new_n11893_), .B(new_n23909_), .ZN(new_n23911_));
  MUX2_X1    g20845(.I0(new_n23911_), .I1(new_n23904_), .S(new_n11891_), .Z(new_n23912_));
  OAI21_X1   g20846(.A1(new_n23912_), .A2(new_n13024_), .B(new_n23888_), .ZN(new_n23913_));
  NOR2_X1    g20847(.A1(new_n23913_), .A2(new_n13714_), .ZN(new_n23914_));
  AOI21_X1   g20848(.A1(new_n13714_), .A2(new_n23886_), .B(new_n23914_), .ZN(new_n23915_));
  AOI21_X1   g20849(.A1(new_n23915_), .A2(new_n12014_), .B(new_n23887_), .ZN(new_n23916_));
  AOI21_X1   g20850(.A1(new_n23916_), .A2(new_n13114_), .B(new_n23885_), .ZN(new_n23917_));
  NOR3_X1    g20851(.A1(new_n23917_), .A2(pi0628), .A3(new_n23886_), .ZN(new_n23918_));
  AOI21_X1   g20852(.A1(new_n23917_), .A2(new_n12031_), .B(new_n23884_), .ZN(new_n23919_));
  NOR3_X1    g20853(.A1(new_n23918_), .A2(new_n23919_), .A3(pi1156), .ZN(new_n23920_));
  INV_X1     g20854(.I(new_n23920_), .ZN(new_n23921_));
  MUX2_X1    g20855(.I0(new_n23921_), .I1(new_n23917_), .S(new_n11868_), .Z(new_n23922_));
  NOR2_X1    g20856(.A1(new_n23922_), .A2(new_n12061_), .ZN(new_n23923_));
  OAI21_X1   g20857(.A1(new_n23884_), .A2(pi0647), .B(pi1157), .ZN(new_n23924_));
  NOR2_X1    g20858(.A1(new_n23923_), .A2(new_n23924_), .ZN(new_n23925_));
  NAND2_X1   g20859(.A1(new_n23925_), .A2(new_n12060_), .ZN(new_n23926_));
  NOR3_X1    g20860(.A1(new_n23922_), .A2(pi0647), .A3(new_n23886_), .ZN(new_n23927_));
  AOI21_X1   g20861(.A1(new_n23922_), .A2(new_n12061_), .B(new_n23884_), .ZN(new_n23928_));
  NOR3_X1    g20862(.A1(new_n23927_), .A2(new_n23928_), .A3(pi1157), .ZN(new_n23929_));
  NOR2_X1    g20863(.A1(new_n23929_), .A2(new_n12060_), .ZN(new_n23930_));
  NAND2_X1   g20864(.A1(new_n23930_), .A2(new_n23926_), .ZN(new_n23931_));
  NAND2_X1   g20865(.A1(new_n23925_), .A2(new_n12060_), .ZN(new_n23932_));
  OAI21_X1   g20866(.A1(new_n14362_), .A2(pi0200), .B(new_n3172_), .ZN(new_n23933_));
  NAND3_X1   g20867(.A1(new_n23933_), .A2(pi0200), .A3(new_n13381_), .ZN(new_n23934_));
  NAND2_X1   g20868(.A1(new_n14359_), .A2(new_n8098_), .ZN(new_n23935_));
  AOI21_X1   g20869(.A1(new_n23935_), .A2(new_n14364_), .B(new_n3232_), .ZN(new_n23936_));
  INV_X1     g20870(.I(pi0606), .ZN(new_n23937_));
  NAND3_X1   g20871(.A1(new_n3231_), .A2(new_n8098_), .A3(new_n23937_), .ZN(new_n23938_));
  AOI21_X1   g20872(.A1(new_n23934_), .A2(new_n23936_), .B(new_n23938_), .ZN(new_n23939_));
  NOR2_X1    g20873(.A1(new_n23884_), .A2(pi0606), .ZN(new_n23940_));
  NOR2_X1    g20874(.A1(new_n23940_), .A2(new_n23939_), .ZN(new_n23941_));
  NOR2_X1    g20875(.A1(new_n23886_), .A2(new_n11924_), .ZN(new_n23942_));
  AOI21_X1   g20876(.A1(new_n23941_), .A2(new_n11924_), .B(new_n23942_), .ZN(new_n23943_));
  NAND3_X1   g20877(.A1(new_n23943_), .A2(pi0609), .A3(new_n23884_), .ZN(new_n23944_));
  INV_X1     g20878(.I(new_n23943_), .ZN(new_n23945_));
  OAI21_X1   g20879(.A1(new_n11903_), .A2(new_n23884_), .B(new_n23945_), .ZN(new_n23946_));
  AOI21_X1   g20880(.A1(new_n23946_), .A2(new_n23944_), .B(pi1155), .ZN(new_n23947_));
  MUX2_X1    g20881(.I0(new_n23943_), .I1(new_n23886_), .S(new_n11903_), .Z(new_n23948_));
  NOR2_X1    g20882(.A1(new_n23948_), .A2(new_n11912_), .ZN(new_n23949_));
  NOR2_X1    g20883(.A1(new_n23947_), .A2(new_n23949_), .ZN(new_n23950_));
  MUX2_X1    g20884(.I0(new_n23950_), .I1(new_n23943_), .S(new_n11870_), .Z(new_n23951_));
  NOR2_X1    g20885(.A1(new_n23951_), .A2(pi0781), .ZN(new_n23952_));
  INV_X1     g20886(.I(new_n23951_), .ZN(new_n23953_));
  MUX2_X1    g20887(.I0(new_n23953_), .I1(new_n23886_), .S(new_n15166_), .Z(new_n23954_));
  AOI21_X1   g20888(.A1(new_n23954_), .A2(pi0781), .B(new_n23952_), .ZN(new_n23955_));
  NAND2_X1   g20889(.A1(new_n23955_), .A2(new_n11985_), .ZN(new_n23956_));
  NOR3_X1    g20890(.A1(new_n23955_), .A2(pi0619), .A3(new_n23886_), .ZN(new_n23957_));
  AOI21_X1   g20891(.A1(new_n23955_), .A2(new_n11967_), .B(new_n23884_), .ZN(new_n23958_));
  NOR3_X1    g20892(.A1(new_n23957_), .A2(new_n23958_), .A3(pi1159), .ZN(new_n23959_));
  NOR2_X1    g20893(.A1(new_n23959_), .A2(new_n11985_), .ZN(new_n23960_));
  XNOR2_X1   g20894(.A1(new_n23960_), .A2(new_n23956_), .ZN(new_n23961_));
  INV_X1     g20895(.I(new_n23961_), .ZN(new_n23962_));
  NOR2_X1    g20896(.A1(new_n23884_), .A2(new_n14624_), .ZN(new_n23963_));
  AOI21_X1   g20897(.A1(new_n23962_), .A2(new_n14624_), .B(new_n23963_), .ZN(new_n23964_));
  NOR2_X1    g20898(.A1(new_n23884_), .A2(new_n12054_), .ZN(new_n23965_));
  INV_X1     g20899(.I(new_n23965_), .ZN(new_n23966_));
  OAI21_X1   g20900(.A1(new_n23964_), .A2(new_n12053_), .B(new_n23966_), .ZN(new_n23967_));
  OAI21_X1   g20901(.A1(new_n23967_), .A2(new_n15077_), .B(new_n12048_), .ZN(new_n23968_));
  AOI21_X1   g20902(.A1(new_n23931_), .A2(new_n23932_), .B(new_n23968_), .ZN(new_n23969_));
  NAND2_X1   g20903(.A1(new_n23964_), .A2(new_n15222_), .ZN(new_n23970_));
  AOI21_X1   g20904(.A1(new_n23921_), .A2(pi0629), .B(pi0792), .ZN(new_n23971_));
  NAND2_X1   g20905(.A1(new_n23970_), .A2(new_n23971_), .ZN(new_n23972_));
  MUX2_X1    g20906(.I0(new_n23961_), .I1(new_n23884_), .S(pi0626), .Z(new_n23973_));
  NOR2_X1    g20907(.A1(new_n23973_), .A2(new_n17171_), .ZN(new_n23974_));
  NOR4_X1    g20908(.A1(new_n23961_), .A2(new_n11994_), .A3(new_n11988_), .A4(new_n23884_), .ZN(new_n23975_));
  NOR2_X1    g20909(.A1(new_n23916_), .A2(new_n17173_), .ZN(new_n23976_));
  OR3_X2     g20910(.A1(new_n23975_), .A2(new_n11986_), .A3(new_n23976_), .Z(new_n23977_));
  OAI21_X1   g20911(.A1(new_n23977_), .A2(new_n23974_), .B(new_n14732_), .ZN(new_n23978_));
  NAND2_X1   g20912(.A1(new_n13657_), .A2(new_n11893_), .ZN(new_n23979_));
  INV_X1     g20913(.I(new_n23941_), .ZN(new_n23980_));
  NOR2_X1    g20914(.A1(new_n17790_), .A2(new_n17791_), .ZN(new_n23981_));
  AOI21_X1   g20915(.A1(new_n23981_), .A2(new_n8098_), .B(pi0038), .ZN(new_n23982_));
  OAI21_X1   g20916(.A1(new_n8098_), .A2(new_n17789_), .B(new_n23982_), .ZN(new_n23983_));
  AOI21_X1   g20917(.A1(new_n12114_), .A2(new_n15189_), .B(new_n23891_), .ZN(new_n23984_));
  NOR2_X1    g20918(.A1(new_n23984_), .A2(pi0606), .ZN(new_n23985_));
  NAND2_X1   g20919(.A1(new_n23983_), .A2(new_n23985_), .ZN(new_n23986_));
  AOI22_X1   g20920(.A1(new_n12277_), .A2(pi0039), .B1(pi0038), .B2(new_n17783_), .ZN(new_n23987_));
  NAND2_X1   g20921(.A1(new_n17777_), .A2(pi0200), .ZN(new_n23988_));
  AOI21_X1   g20922(.A1(new_n17780_), .A2(new_n8098_), .B(pi0038), .ZN(new_n23989_));
  NAND3_X1   g20923(.A1(new_n17784_), .A2(pi0038), .A3(pi0200), .ZN(new_n23990_));
  NAND3_X1   g20924(.A1(new_n23990_), .A2(pi0606), .A3(new_n3231_), .ZN(new_n23991_));
  AOI21_X1   g20925(.A1(new_n23988_), .A2(new_n23989_), .B(new_n23991_), .ZN(new_n23992_));
  NOR2_X1    g20926(.A1(new_n3231_), .A2(new_n8098_), .ZN(new_n23993_));
  OAI22_X1   g20927(.A1(new_n23992_), .A2(new_n23993_), .B1(pi0200), .B2(new_n23987_), .ZN(new_n23994_));
  NAND4_X1   g20928(.A1(new_n23986_), .A2(pi0643), .A3(new_n3232_), .A4(new_n23994_), .ZN(new_n23995_));
  OAI21_X1   g20929(.A1(pi0643), .A2(new_n23941_), .B(new_n23995_), .ZN(new_n23996_));
  MUX2_X1    g20930(.I0(new_n23996_), .I1(new_n23980_), .S(pi0625), .Z(new_n23997_));
  OAI22_X1   g20931(.A1(new_n23909_), .A2(pi0608), .B1(new_n23979_), .B2(new_n23997_), .ZN(new_n23998_));
  NOR2_X1    g20932(.A1(new_n23996_), .A2(pi0778), .ZN(new_n23999_));
  AOI21_X1   g20933(.A1(new_n23998_), .A2(pi0778), .B(new_n23999_), .ZN(new_n24000_));
  NOR4_X1    g20934(.A1(new_n23912_), .A2(new_n11903_), .A3(pi1155), .A4(new_n24000_), .ZN(new_n24001_));
  OR2_X2     g20935(.A1(new_n23947_), .A2(new_n11923_), .Z(new_n24002_));
  AND3_X2    g20936(.A1(new_n23912_), .A2(pi0609), .A3(pi1155), .Z(new_n24003_));
  OAI21_X1   g20937(.A1(new_n23948_), .A2(new_n11912_), .B(new_n11923_), .ZN(new_n24004_));
  OAI22_X1   g20938(.A1(new_n24003_), .A2(new_n24004_), .B1(new_n24001_), .B2(new_n24002_), .ZN(new_n24005_));
  MUX2_X1    g20939(.I0(new_n24005_), .I1(new_n24000_), .S(new_n11870_), .Z(new_n24006_));
  NAND2_X1   g20940(.A1(new_n24006_), .A2(new_n11969_), .ZN(new_n24007_));
  OAI21_X1   g20941(.A1(new_n23913_), .A2(pi0618), .B(pi1154), .ZN(new_n24008_));
  NOR3_X1    g20942(.A1(new_n11950_), .A2(pi0618), .A3(pi0627), .ZN(new_n24009_));
  NAND2_X1   g20943(.A1(new_n23953_), .A2(new_n24009_), .ZN(new_n24010_));
  NAND4_X1   g20944(.A1(new_n24006_), .A2(pi0618), .A3(new_n24008_), .A4(new_n24010_), .ZN(new_n24011_));
  AND2_X2    g20945(.A1(new_n24006_), .A2(new_n11934_), .Z(new_n24012_));
  NOR2_X1    g20946(.A1(new_n11934_), .A2(pi1154), .ZN(new_n24013_));
  NAND2_X1   g20947(.A1(new_n23953_), .A2(new_n24013_), .ZN(new_n24014_));
  AND3_X2    g20948(.A1(new_n24014_), .A2(new_n11949_), .A3(new_n11950_), .Z(new_n24015_));
  OAI21_X1   g20949(.A1(new_n11934_), .A2(new_n23913_), .B(new_n24015_), .ZN(new_n24016_));
  OAI21_X1   g20950(.A1(new_n24012_), .A2(new_n24016_), .B(new_n24011_), .ZN(new_n24017_));
  NAND2_X1   g20951(.A1(new_n24017_), .A2(pi0781), .ZN(new_n24018_));
  XOR2_X1    g20952(.A1(new_n24018_), .A2(new_n24007_), .Z(new_n24019_));
  OR3_X2     g20953(.A1(new_n23915_), .A2(new_n11967_), .A3(new_n11869_), .Z(new_n24020_));
  NAND2_X1   g20954(.A1(new_n24020_), .A2(new_n11966_), .ZN(new_n24021_));
  INV_X1     g20955(.I(new_n24019_), .ZN(new_n24022_));
  NAND4_X1   g20956(.A1(new_n24022_), .A2(pi0619), .A3(new_n11869_), .A4(new_n23915_), .ZN(new_n24023_));
  NAND2_X1   g20957(.A1(new_n24023_), .A2(new_n23959_), .ZN(new_n24024_));
  NAND2_X1   g20958(.A1(new_n24022_), .A2(new_n11985_), .ZN(new_n24025_));
  AOI21_X1   g20959(.A1(new_n24025_), .A2(new_n11998_), .B(new_n17371_), .ZN(new_n24026_));
  NAND4_X1   g20960(.A1(new_n24024_), .A2(new_n24026_), .A3(new_n23978_), .A4(new_n24021_), .ZN(new_n24027_));
  AOI21_X1   g20961(.A1(new_n24027_), .A2(new_n23972_), .B(new_n14725_), .ZN(new_n24028_));
  NOR2_X1    g20962(.A1(new_n24028_), .A2(new_n23969_), .ZN(new_n24029_));
  NOR2_X1    g20963(.A1(new_n23922_), .A2(pi0787), .ZN(new_n24030_));
  NOR2_X1    g20964(.A1(new_n23925_), .A2(new_n12048_), .ZN(new_n24031_));
  AND2_X2    g20965(.A1(new_n24031_), .A2(new_n23929_), .Z(new_n24032_));
  OAI21_X1   g20966(.A1(new_n24032_), .A2(new_n24030_), .B(new_n12082_), .ZN(new_n24033_));
  NOR2_X1    g20967(.A1(new_n23884_), .A2(new_n12092_), .ZN(new_n24034_));
  AOI21_X1   g20968(.A1(new_n23967_), .A2(new_n12092_), .B(new_n24034_), .ZN(new_n24035_));
  NAND3_X1   g20969(.A1(new_n12081_), .A2(pi0644), .A3(pi0715), .ZN(new_n24036_));
  OAI21_X1   g20970(.A1(new_n24035_), .A2(new_n24036_), .B(pi0644), .ZN(new_n24037_));
  AOI21_X1   g20971(.A1(new_n24033_), .A2(pi0715), .B(new_n24037_), .ZN(new_n24038_));
  OAI21_X1   g20972(.A1(new_n24032_), .A2(new_n24030_), .B(pi0644), .ZN(new_n24039_));
  NAND2_X1   g20973(.A1(new_n12082_), .A2(new_n12099_), .ZN(new_n24040_));
  NOR2_X1    g20974(.A1(pi0644), .A2(pi1160), .ZN(new_n24041_));
  OAI21_X1   g20975(.A1(new_n24035_), .A2(new_n24040_), .B(new_n24041_), .ZN(new_n24042_));
  AOI21_X1   g20976(.A1(new_n24039_), .A2(new_n12099_), .B(new_n24042_), .ZN(new_n24043_));
  NOR4_X1    g20977(.A1(new_n24038_), .A2(new_n24043_), .A3(new_n24029_), .A4(new_n11867_), .ZN(new_n24044_));
  XOR2_X1    g20978(.A1(new_n24044_), .A2(new_n24029_), .Z(new_n24045_));
  NAND2_X1   g20979(.A1(po1038), .A2(pi0200), .ZN(new_n24046_));
  OAI21_X1   g20980(.A1(new_n24045_), .A2(po1038), .B(new_n24046_), .ZN(po0357));
  INV_X1     g20981(.I(pi0201), .ZN(new_n24048_));
  NAND2_X1   g20982(.A1(new_n2891_), .A2(new_n8589_), .ZN(new_n24049_));
  NOR3_X1    g20983(.A1(new_n3227_), .A2(new_n3202_), .A3(new_n2563_), .ZN(new_n24058_));
  NOR2_X1    g20984(.A1(new_n3234_), .A2(new_n5429_), .ZN(new_n24059_));
  AOI21_X1   g20985(.A1(new_n24059_), .A2(new_n2490_), .B(pi0332), .ZN(new_n24060_));
  NOR4_X1    g20986(.A1(new_n24060_), .A2(new_n3227_), .A3(new_n2533_), .A4(new_n24058_), .ZN(new_n24061_));
  INV_X1     g20987(.I(new_n24060_), .ZN(new_n24062_));
  NAND4_X1   g20988(.A1(new_n24062_), .A2(new_n5205_), .A3(new_n2563_), .A4(new_n5222_), .ZN(new_n24063_));
  NOR2_X1    g20989(.A1(new_n3503_), .A2(pi0332), .ZN(new_n24064_));
  NOR4_X1    g20990(.A1(new_n24064_), .A2(new_n5055_), .A3(new_n2563_), .A4(new_n3405_), .ZN(new_n24065_));
  NAND2_X1   g20991(.A1(new_n24063_), .A2(new_n24065_), .ZN(new_n24066_));
  NOR2_X1    g20992(.A1(new_n24066_), .A2(new_n24061_), .ZN(new_n24067_));
  INV_X1     g20993(.I(new_n24067_), .ZN(new_n24068_));
  INV_X1     g20994(.I(pi0233), .ZN(new_n24069_));
  INV_X1     g20995(.I(pi0237), .ZN(new_n24070_));
  NOR2_X1    g20996(.A1(new_n24069_), .A2(new_n24070_), .ZN(new_n24071_));
  NAND3_X1   g20997(.A1(new_n24068_), .A2(new_n24048_), .A3(new_n24071_), .ZN(new_n24072_));
  INV_X1     g20998(.I(new_n24071_), .ZN(new_n24073_));
  NAND2_X1   g20999(.A1(pi0096), .A2(pi0210), .ZN(new_n24074_));
  NOR4_X1    g21000(.A1(new_n5432_), .A2(new_n11749_), .A3(new_n2659_), .A4(new_n2601_), .ZN(new_n24075_));
  OAI21_X1   g21001(.A1(new_n5429_), .A2(new_n24074_), .B(new_n24075_), .ZN(new_n24076_));
  NOR2_X1    g21002(.A1(new_n24076_), .A2(new_n24073_), .ZN(new_n24077_));
  NAND2_X1   g21003(.A1(new_n24077_), .A2(pi0201), .ZN(new_n24078_));
  NAND2_X1   g21004(.A1(new_n24072_), .A2(new_n24078_), .ZN(po0358));
  NOR2_X1    g21005(.A1(new_n24070_), .A2(pi0233), .ZN(new_n24080_));
  NAND2_X1   g21006(.A1(new_n24068_), .A2(new_n24080_), .ZN(new_n24081_));
  INV_X1     g21007(.I(new_n24080_), .ZN(new_n24082_));
  NOR2_X1    g21008(.A1(new_n24076_), .A2(new_n24082_), .ZN(new_n24083_));
  NAND2_X1   g21009(.A1(new_n24083_), .A2(pi0202), .ZN(new_n24084_));
  OAI21_X1   g21010(.A1(new_n24081_), .A2(pi0202), .B(new_n24084_), .ZN(po0359));
  NOR2_X1    g21011(.A1(pi0233), .A2(pi0237), .ZN(new_n24086_));
  INV_X1     g21012(.I(new_n24086_), .ZN(new_n24087_));
  NOR2_X1    g21013(.A1(new_n24067_), .A2(new_n24087_), .ZN(new_n24088_));
  NOR2_X1    g21014(.A1(new_n24076_), .A2(new_n24087_), .ZN(new_n24089_));
  NAND2_X1   g21015(.A1(new_n24089_), .A2(pi0203), .ZN(new_n24090_));
  OAI21_X1   g21016(.A1(new_n24088_), .A2(pi0203), .B(new_n24090_), .ZN(po0360));
  NAND2_X1   g21017(.A1(new_n2587_), .A2(new_n5394_), .ZN(new_n24092_));
  AOI21_X1   g21018(.A1(new_n15305_), .A2(pi0299), .B(pi0468), .ZN(new_n24093_));
  AOI22_X1   g21019(.A1(new_n5100_), .A2(pi0468), .B1(new_n24092_), .B2(new_n24093_), .ZN(new_n24094_));
  OAI21_X1   g21020(.A1(new_n24049_), .A2(new_n24094_), .B(new_n2563_), .ZN(new_n24095_));
  NAND2_X1   g21021(.A1(new_n24095_), .A2(new_n5918_), .ZN(new_n24096_));
  NAND2_X1   g21022(.A1(new_n5217_), .A2(pi0468), .ZN(new_n24097_));
  NAND2_X1   g21023(.A1(new_n9909_), .A2(new_n5394_), .ZN(new_n24098_));
  NAND4_X1   g21024(.A1(new_n5220_), .A2(pi0299), .A3(new_n24097_), .A4(new_n24098_), .ZN(new_n24099_));
  OAI21_X1   g21025(.A1(new_n24099_), .A2(new_n2490_), .B(new_n2563_), .ZN(new_n24100_));
  AOI21_X1   g21026(.A1(new_n24100_), .A2(new_n11280_), .B(pi0074), .ZN(new_n24101_));
  NOR3_X1    g21027(.A1(new_n5219_), .A2(new_n2491_), .A3(new_n3234_), .ZN(new_n24102_));
  NOR2_X1    g21028(.A1(new_n24102_), .A2(pi0332), .ZN(new_n24103_));
  NOR2_X1    g21029(.A1(new_n24103_), .A2(new_n3227_), .ZN(new_n24104_));
  NOR3_X1    g21030(.A1(new_n11279_), .A2(pi0074), .A3(pi0332), .ZN(new_n24105_));
  OAI22_X1   g21031(.A1(new_n24104_), .A2(new_n3503_), .B1(pi0055), .B2(new_n24105_), .ZN(new_n24106_));
  AOI21_X1   g21032(.A1(new_n24096_), .A2(new_n24101_), .B(new_n24106_), .ZN(new_n24107_));
  NAND4_X1   g21033(.A1(new_n24102_), .A2(new_n5205_), .A3(new_n2563_), .A4(new_n5222_), .ZN(new_n24108_));
  NAND2_X1   g21034(.A1(new_n24108_), .A2(new_n24065_), .ZN(new_n24109_));
  NOR2_X1    g21035(.A1(new_n24107_), .A2(new_n24109_), .ZN(new_n24110_));
  INV_X1     g21036(.I(new_n24110_), .ZN(new_n24111_));
  NAND2_X1   g21037(.A1(new_n24111_), .A2(new_n24071_), .ZN(new_n24112_));
  NOR4_X1    g21038(.A1(new_n5227_), .A2(new_n2659_), .A3(new_n2601_), .A4(new_n11749_), .ZN(new_n24113_));
  OAI21_X1   g21039(.A1(new_n5219_), .A2(new_n24074_), .B(new_n24113_), .ZN(new_n24114_));
  NOR2_X1    g21040(.A1(new_n24114_), .A2(new_n24073_), .ZN(new_n24115_));
  NAND2_X1   g21041(.A1(new_n24115_), .A2(pi0204), .ZN(new_n24116_));
  OAI21_X1   g21042(.A1(new_n24112_), .A2(pi0204), .B(new_n24116_), .ZN(po0361));
  NAND2_X1   g21043(.A1(new_n24111_), .A2(new_n24080_), .ZN(new_n24118_));
  NOR2_X1    g21044(.A1(new_n24114_), .A2(new_n24082_), .ZN(new_n24119_));
  NAND2_X1   g21045(.A1(new_n24119_), .A2(pi0205), .ZN(new_n24120_));
  OAI21_X1   g21046(.A1(new_n24118_), .A2(pi0205), .B(new_n24120_), .ZN(po0362));
  NOR2_X1    g21047(.A1(new_n24069_), .A2(pi0237), .ZN(new_n24122_));
  NAND2_X1   g21048(.A1(new_n24111_), .A2(new_n24122_), .ZN(new_n24123_));
  INV_X1     g21049(.I(new_n24122_), .ZN(new_n24124_));
  NOR2_X1    g21050(.A1(new_n24114_), .A2(new_n24124_), .ZN(new_n24125_));
  NAND2_X1   g21051(.A1(new_n24125_), .A2(pi0206), .ZN(new_n24126_));
  OAI21_X1   g21052(.A1(new_n24123_), .A2(pi0206), .B(new_n24126_), .ZN(po0363));
  NOR2_X1    g21053(.A1(new_n12965_), .A2(new_n14624_), .ZN(new_n24128_));
  NOR2_X1    g21054(.A1(new_n20355_), .A2(new_n3232_), .ZN(new_n24129_));
  AOI21_X1   g21055(.A1(new_n24129_), .A2(new_n11924_), .B(pi0785), .ZN(new_n24130_));
  OAI21_X1   g21056(.A1(new_n11924_), .A2(new_n14396_), .B(new_n24130_), .ZN(new_n24131_));
  NOR2_X1    g21057(.A1(new_n24129_), .A2(new_n11914_), .ZN(new_n24132_));
  AOI22_X1   g21058(.A1(new_n24132_), .A2(new_n11903_), .B1(new_n14396_), .B2(new_n12997_), .ZN(new_n24133_));
  NOR2_X1    g21059(.A1(new_n24133_), .A2(pi1155), .ZN(new_n24134_));
  AOI21_X1   g21060(.A1(new_n24132_), .A2(pi0609), .B(pi1155), .ZN(new_n24135_));
  OAI21_X1   g21061(.A1(new_n11915_), .A2(new_n12965_), .B(new_n24135_), .ZN(new_n24136_));
  AOI21_X1   g21062(.A1(new_n24136_), .A2(new_n24134_), .B(new_n11870_), .ZN(new_n24137_));
  XNOR2_X1   g21063(.A1(new_n24137_), .A2(new_n24131_), .ZN(new_n24138_));
  NAND2_X1   g21064(.A1(new_n24138_), .A2(pi0618), .ZN(new_n24139_));
  AOI21_X1   g21065(.A1(new_n14396_), .A2(new_n11934_), .B(pi1154), .ZN(new_n24140_));
  NAND2_X1   g21066(.A1(new_n24139_), .A2(new_n24140_), .ZN(new_n24141_));
  OAI21_X1   g21067(.A1(new_n14396_), .A2(new_n11934_), .B(new_n11950_), .ZN(new_n24142_));
  AOI21_X1   g21068(.A1(new_n24138_), .A2(pi0618), .B(new_n24142_), .ZN(new_n24143_));
  NAND2_X1   g21069(.A1(new_n24141_), .A2(new_n24143_), .ZN(new_n24144_));
  MUX2_X1    g21070(.I0(new_n24144_), .I1(new_n24138_), .S(new_n11969_), .Z(new_n24145_));
  NAND2_X1   g21071(.A1(new_n24145_), .A2(new_n11985_), .ZN(new_n24146_));
  NAND2_X1   g21072(.A1(new_n24145_), .A2(pi0619), .ZN(new_n24147_));
  AOI21_X1   g21073(.A1(new_n14396_), .A2(new_n11967_), .B(pi1159), .ZN(new_n24148_));
  NAND2_X1   g21074(.A1(new_n24147_), .A2(new_n24148_), .ZN(new_n24149_));
  INV_X1     g21075(.I(new_n24149_), .ZN(new_n24150_));
  AOI21_X1   g21076(.A1(new_n12965_), .A2(pi0619), .B(pi1159), .ZN(new_n24151_));
  NAND2_X1   g21077(.A1(new_n24147_), .A2(new_n24151_), .ZN(new_n24152_));
  OAI21_X1   g21078(.A1(new_n24150_), .A2(new_n24152_), .B(pi0789), .ZN(new_n24153_));
  XOR2_X1    g21079(.A1(new_n24153_), .A2(new_n24146_), .Z(new_n24154_));
  AOI21_X1   g21080(.A1(new_n24154_), .A2(new_n14624_), .B(new_n24128_), .ZN(new_n24155_));
  NOR2_X1    g21081(.A1(new_n12965_), .A2(new_n12054_), .ZN(new_n24156_));
  INV_X1     g21082(.I(new_n24156_), .ZN(new_n24157_));
  OAI21_X1   g21083(.A1(new_n24155_), .A2(new_n12053_), .B(new_n24157_), .ZN(new_n24158_));
  NAND3_X1   g21084(.A1(new_n17506_), .A2(new_n3231_), .A3(new_n11924_), .ZN(new_n24159_));
  NOR2_X1    g21085(.A1(new_n24159_), .A2(new_n14627_), .ZN(new_n24160_));
  INV_X1     g21086(.I(new_n24160_), .ZN(new_n24161_));
  NOR2_X1    g21087(.A1(new_n24161_), .A2(new_n14636_), .ZN(new_n24162_));
  NOR2_X1    g21088(.A1(new_n24162_), .A2(new_n14642_), .ZN(new_n24163_));
  INV_X1     g21089(.I(new_n24163_), .ZN(new_n24164_));
  NOR2_X1    g21090(.A1(new_n24164_), .A2(new_n11997_), .ZN(new_n24165_));
  INV_X1     g21091(.I(new_n24165_), .ZN(new_n24166_));
  NOR2_X1    g21092(.A1(new_n24166_), .A2(new_n12053_), .ZN(new_n24167_));
  INV_X1     g21093(.I(new_n24167_), .ZN(new_n24168_));
  AOI21_X1   g21094(.A1(new_n24158_), .A2(new_n24168_), .B(new_n8087_), .ZN(new_n24169_));
  NAND2_X1   g21095(.A1(new_n24169_), .A2(pi0623), .ZN(new_n24170_));
  NOR2_X1    g21096(.A1(new_n12965_), .A2(pi0207), .ZN(new_n24171_));
  INV_X1     g21097(.I(new_n24171_), .ZN(new_n24172_));
  OAI21_X1   g21098(.A1(pi0623), .A2(new_n24172_), .B(new_n24170_), .ZN(new_n24173_));
  INV_X1     g21099(.I(pi0710), .ZN(new_n24174_));
  NOR2_X1    g21100(.A1(new_n14396_), .A2(new_n12067_), .ZN(new_n24175_));
  NOR2_X1    g21101(.A1(new_n12965_), .A2(new_n13114_), .ZN(new_n24176_));
  NOR2_X1    g21102(.A1(new_n14396_), .A2(new_n12014_), .ZN(new_n24177_));
  NOR2_X1    g21103(.A1(new_n12965_), .A2(new_n11961_), .ZN(new_n24178_));
  NAND3_X1   g21104(.A1(new_n12970_), .A2(new_n11893_), .A3(pi0778), .ZN(new_n24179_));
  NOR2_X1    g21105(.A1(new_n13024_), .A2(new_n24179_), .ZN(new_n24180_));
  AOI21_X1   g21106(.A1(new_n12965_), .A2(new_n13024_), .B(new_n24180_), .ZN(new_n24181_));
  INV_X1     g21107(.I(new_n24181_), .ZN(new_n24182_));
  NOR2_X1    g21108(.A1(new_n24182_), .A2(new_n13714_), .ZN(new_n24183_));
  NOR2_X1    g21109(.A1(new_n24183_), .A2(new_n24178_), .ZN(new_n24184_));
  AOI21_X1   g21110(.A1(new_n24184_), .A2(new_n12014_), .B(new_n24177_), .ZN(new_n24185_));
  AOI21_X1   g21111(.A1(new_n24185_), .A2(new_n13114_), .B(new_n24176_), .ZN(new_n24186_));
  INV_X1     g21112(.I(new_n24186_), .ZN(new_n24187_));
  NOR2_X1    g21113(.A1(new_n24187_), .A2(new_n12066_), .ZN(new_n24188_));
  NOR2_X1    g21114(.A1(new_n24188_), .A2(new_n24175_), .ZN(new_n24189_));
  INV_X1     g21115(.I(new_n17547_), .ZN(new_n24190_));
  NOR2_X1    g21116(.A1(new_n24190_), .A2(new_n13636_), .ZN(new_n24191_));
  INV_X1     g21117(.I(new_n24191_), .ZN(new_n24192_));
  NOR2_X1    g21118(.A1(new_n24192_), .A2(new_n13717_), .ZN(new_n24193_));
  INV_X1     g21119(.I(new_n24193_), .ZN(new_n24194_));
  NOR2_X1    g21120(.A1(new_n24194_), .A2(new_n12066_), .ZN(new_n24195_));
  INV_X1     g21121(.I(new_n24195_), .ZN(new_n24196_));
  NOR2_X1    g21122(.A1(new_n24196_), .A2(new_n8087_), .ZN(new_n24197_));
  AOI21_X1   g21123(.A1(new_n24189_), .A2(new_n8087_), .B(new_n24197_), .ZN(new_n24198_));
  NOR2_X1    g21124(.A1(new_n24198_), .A2(new_n24174_), .ZN(new_n24199_));
  AOI21_X1   g21125(.A1(new_n24174_), .A2(new_n24171_), .B(new_n24199_), .ZN(new_n24200_));
  NAND2_X1   g21126(.A1(new_n24200_), .A2(pi0647), .ZN(new_n24201_));
  AOI21_X1   g21127(.A1(new_n24172_), .A2(new_n12061_), .B(pi1157), .ZN(new_n24202_));
  AOI21_X1   g21128(.A1(new_n24201_), .A2(new_n24202_), .B(pi0630), .ZN(new_n24203_));
  AOI21_X1   g21129(.A1(new_n24171_), .A2(pi0647), .B(pi1157), .ZN(new_n24204_));
  AND3_X2    g21130(.A1(new_n24201_), .A2(pi0630), .A3(new_n24204_), .Z(new_n24205_));
  NOR4_X1    g21131(.A1(new_n24173_), .A2(new_n15183_), .A3(new_n24203_), .A4(new_n24205_), .ZN(new_n24206_));
  INV_X1     g21132(.I(new_n12051_), .ZN(new_n24207_));
  MUX2_X1    g21133(.I0(new_n24186_), .I1(new_n12965_), .S(pi0628), .Z(new_n24208_));
  NOR2_X1    g21134(.A1(new_n24208_), .A2(new_n24207_), .ZN(new_n24209_));
  INV_X1     g21135(.I(new_n24209_), .ZN(new_n24210_));
  NOR3_X1    g21136(.A1(new_n12031_), .A2(new_n12026_), .A3(pi0792), .ZN(new_n24211_));
  NAND2_X1   g21137(.A1(new_n24210_), .A2(new_n24211_), .ZN(new_n24212_));
  NAND3_X1   g21138(.A1(new_n14346_), .A2(new_n3231_), .A3(new_n14341_), .ZN(new_n24213_));
  NAND4_X1   g21139(.A1(new_n24213_), .A2(new_n14396_), .A3(pi0625), .A4(new_n11893_), .ZN(new_n24214_));
  OAI21_X1   g21140(.A1(new_n14396_), .A2(new_n12970_), .B(new_n11893_), .ZN(new_n24215_));
  NOR2_X1    g21141(.A1(new_n24215_), .A2(new_n13657_), .ZN(new_n24216_));
  NOR3_X1    g21142(.A1(new_n23609_), .A2(new_n3232_), .A3(new_n14340_), .ZN(new_n24217_));
  OAI21_X1   g21143(.A1(new_n24217_), .A2(pi0625), .B(new_n12965_), .ZN(new_n24218_));
  NOR3_X1    g21144(.A1(new_n24213_), .A2(new_n12965_), .A3(pi0625), .ZN(new_n24219_));
  OAI21_X1   g21145(.A1(new_n12965_), .A2(new_n13659_), .B(new_n12977_), .ZN(new_n24220_));
  NOR2_X1    g21146(.A1(new_n24219_), .A2(new_n24220_), .ZN(new_n24221_));
  AOI22_X1   g21147(.A1(new_n24221_), .A2(new_n24218_), .B1(new_n24216_), .B2(new_n24214_), .ZN(new_n24222_));
  MUX2_X1    g21148(.I0(new_n24222_), .I1(new_n24213_), .S(new_n11891_), .Z(new_n24223_));
  NOR2_X1    g21149(.A1(new_n24179_), .A2(pi0609), .ZN(new_n24224_));
  INV_X1     g21150(.I(new_n24224_), .ZN(new_n24225_));
  OAI21_X1   g21151(.A1(new_n24223_), .A2(new_n11903_), .B(new_n24225_), .ZN(new_n24226_));
  MUX2_X1    g21152(.I0(new_n24226_), .I1(new_n12965_), .S(new_n11912_), .Z(new_n24227_));
  NOR3_X1    g21153(.A1(new_n24222_), .A2(new_n11891_), .A3(new_n24217_), .ZN(new_n24228_));
  AOI21_X1   g21154(.A1(new_n24222_), .A2(pi0778), .B(new_n24213_), .ZN(new_n24229_));
  OAI21_X1   g21155(.A1(new_n24228_), .A2(new_n24229_), .B(new_n11903_), .ZN(new_n24230_));
  NOR2_X1    g21156(.A1(new_n24179_), .A2(new_n11903_), .ZN(new_n24231_));
  INV_X1     g21157(.I(new_n24231_), .ZN(new_n24232_));
  NAND4_X1   g21158(.A1(new_n24230_), .A2(pi1155), .A3(new_n12965_), .A4(new_n24232_), .ZN(new_n24233_));
  AOI21_X1   g21159(.A1(new_n12965_), .A2(pi0625), .B(pi1153), .ZN(new_n24234_));
  NAND3_X1   g21160(.A1(new_n24214_), .A2(new_n24234_), .A3(pi0608), .ZN(new_n24235_));
  NAND4_X1   g21161(.A1(new_n22851_), .A2(new_n15823_), .A3(new_n12970_), .A4(new_n3231_), .ZN(new_n24236_));
  AOI21_X1   g21162(.A1(new_n14396_), .A2(new_n13434_), .B(new_n12978_), .ZN(new_n24237_));
  NAND3_X1   g21163(.A1(new_n24218_), .A2(new_n24237_), .A3(new_n24236_), .ZN(new_n24238_));
  NAND2_X1   g21164(.A1(new_n24235_), .A2(new_n24238_), .ZN(new_n24239_));
  NAND3_X1   g21165(.A1(new_n24239_), .A2(pi0778), .A3(new_n24213_), .ZN(new_n24240_));
  OAI21_X1   g21166(.A1(new_n24239_), .A2(new_n11891_), .B(new_n24217_), .ZN(new_n24241_));
  AOI21_X1   g21167(.A1(new_n24241_), .A2(new_n24240_), .B(pi0609), .ZN(new_n24242_));
  OAI22_X1   g21168(.A1(new_n24242_), .A2(new_n24231_), .B1(new_n11912_), .B2(new_n12965_), .ZN(new_n24243_));
  AOI21_X1   g21169(.A1(new_n24233_), .A2(new_n24243_), .B(pi0660), .ZN(new_n24244_));
  AOI21_X1   g21170(.A1(new_n24227_), .A2(pi0660), .B(new_n24244_), .ZN(new_n24245_));
  MUX2_X1    g21171(.I0(new_n24245_), .I1(new_n24223_), .S(new_n11870_), .Z(new_n24246_));
  NOR2_X1    g21172(.A1(new_n24181_), .A2(pi0618), .ZN(new_n24247_));
  AOI21_X1   g21173(.A1(new_n24246_), .A2(pi0618), .B(new_n24247_), .ZN(new_n24248_));
  MUX2_X1    g21174(.I0(new_n24248_), .I1(new_n14396_), .S(new_n11950_), .Z(new_n24249_));
  NOR2_X1    g21175(.A1(new_n24181_), .A2(new_n11934_), .ZN(new_n24250_));
  MUX2_X1    g21176(.I0(new_n24239_), .I1(new_n24217_), .S(new_n11891_), .Z(new_n24251_));
  NOR3_X1    g21177(.A1(new_n24245_), .A2(new_n11870_), .A3(new_n24251_), .ZN(new_n24252_));
  AOI21_X1   g21178(.A1(new_n24245_), .A2(pi0785), .B(new_n24223_), .ZN(new_n24253_));
  NOR3_X1    g21179(.A1(new_n24252_), .A2(new_n24253_), .A3(pi0618), .ZN(new_n24254_));
  NOR4_X1    g21180(.A1(new_n24254_), .A2(new_n11950_), .A3(new_n14396_), .A4(new_n24250_), .ZN(new_n24255_));
  INV_X1     g21181(.I(new_n24250_), .ZN(new_n24256_));
  AOI21_X1   g21182(.A1(new_n24251_), .A2(pi0609), .B(new_n24224_), .ZN(new_n24257_));
  NOR3_X1    g21183(.A1(new_n24257_), .A2(new_n11912_), .A3(new_n12965_), .ZN(new_n24258_));
  AOI21_X1   g21184(.A1(new_n24257_), .A2(pi1155), .B(new_n14396_), .ZN(new_n24259_));
  OAI21_X1   g21185(.A1(new_n24258_), .A2(new_n24259_), .B(pi0660), .ZN(new_n24260_));
  NOR4_X1    g21186(.A1(new_n24242_), .A2(new_n11912_), .A3(new_n14396_), .A4(new_n24231_), .ZN(new_n24261_));
  AOI22_X1   g21187(.A1(new_n24230_), .A2(new_n24232_), .B1(pi1155), .B2(new_n14396_), .ZN(new_n24262_));
  OAI21_X1   g21188(.A1(new_n24262_), .A2(new_n24261_), .B(new_n11923_), .ZN(new_n24263_));
  NAND2_X1   g21189(.A1(new_n24260_), .A2(new_n24263_), .ZN(new_n24264_));
  NAND3_X1   g21190(.A1(new_n24264_), .A2(pi0785), .A3(new_n24223_), .ZN(new_n24265_));
  OAI21_X1   g21191(.A1(new_n24264_), .A2(new_n11870_), .B(new_n24251_), .ZN(new_n24266_));
  NAND3_X1   g21192(.A1(new_n24266_), .A2(new_n24265_), .A3(new_n11934_), .ZN(new_n24267_));
  AOI22_X1   g21193(.A1(new_n24267_), .A2(new_n24256_), .B1(pi1154), .B2(new_n14396_), .ZN(new_n24268_));
  OAI21_X1   g21194(.A1(new_n24255_), .A2(new_n24268_), .B(new_n11949_), .ZN(new_n24269_));
  OAI21_X1   g21195(.A1(new_n11949_), .A2(new_n24249_), .B(new_n24269_), .ZN(new_n24270_));
  MUX2_X1    g21196(.I0(new_n24270_), .I1(new_n24246_), .S(new_n11969_), .Z(new_n24271_));
  INV_X1     g21197(.I(new_n24184_), .ZN(new_n24272_));
  NOR2_X1    g21198(.A1(new_n24272_), .A2(pi0619), .ZN(new_n24273_));
  AOI21_X1   g21199(.A1(new_n24271_), .A2(pi0619), .B(new_n24273_), .ZN(new_n24274_));
  MUX2_X1    g21200(.I0(new_n24274_), .I1(new_n14396_), .S(new_n11869_), .Z(new_n24275_));
  NOR2_X1    g21201(.A1(new_n24272_), .A2(new_n11967_), .ZN(new_n24276_));
  MUX2_X1    g21202(.I0(new_n24264_), .I1(new_n24251_), .S(new_n11870_), .Z(new_n24277_));
  NOR2_X1    g21203(.A1(new_n24277_), .A2(pi0781), .ZN(new_n24278_));
  INV_X1     g21204(.I(new_n24278_), .ZN(new_n24279_));
  INV_X1     g21205(.I(new_n24247_), .ZN(new_n24280_));
  OAI21_X1   g21206(.A1(new_n24277_), .A2(new_n11934_), .B(new_n24280_), .ZN(new_n24281_));
  MUX2_X1    g21207(.I0(new_n24281_), .I1(new_n12965_), .S(new_n11950_), .Z(new_n24282_));
  NAND4_X1   g21208(.A1(new_n24267_), .A2(pi1154), .A3(new_n12965_), .A4(new_n24256_), .ZN(new_n24283_));
  OAI22_X1   g21209(.A1(new_n24254_), .A2(new_n24250_), .B1(new_n11950_), .B2(new_n12965_), .ZN(new_n24284_));
  AOI21_X1   g21210(.A1(new_n24284_), .A2(new_n24283_), .B(pi0627), .ZN(new_n24285_));
  AOI21_X1   g21211(.A1(pi0627), .A2(new_n24282_), .B(new_n24285_), .ZN(new_n24286_));
  NOR3_X1    g21212(.A1(new_n24286_), .A2(new_n11969_), .A3(new_n24279_), .ZN(new_n24287_));
  AOI21_X1   g21213(.A1(new_n24270_), .A2(pi0781), .B(new_n24278_), .ZN(new_n24288_));
  NOR3_X1    g21214(.A1(new_n24287_), .A2(new_n24288_), .A3(pi0619), .ZN(new_n24289_));
  NOR4_X1    g21215(.A1(new_n24289_), .A2(new_n11869_), .A3(new_n14396_), .A4(new_n24276_), .ZN(new_n24290_));
  INV_X1     g21216(.I(new_n24276_), .ZN(new_n24291_));
  NAND3_X1   g21217(.A1(new_n24270_), .A2(pi0781), .A3(new_n24278_), .ZN(new_n24292_));
  OAI21_X1   g21218(.A1(new_n24286_), .A2(new_n11969_), .B(new_n24279_), .ZN(new_n24293_));
  NAND3_X1   g21219(.A1(new_n24293_), .A2(new_n24292_), .A3(new_n11967_), .ZN(new_n24294_));
  AOI22_X1   g21220(.A1(new_n24294_), .A2(new_n24291_), .B1(pi1159), .B2(new_n14396_), .ZN(new_n24295_));
  OAI21_X1   g21221(.A1(new_n24290_), .A2(new_n24295_), .B(new_n11966_), .ZN(new_n24296_));
  OAI21_X1   g21222(.A1(new_n11966_), .A2(new_n24275_), .B(new_n24296_), .ZN(new_n24297_));
  MUX2_X1    g21223(.I0(new_n24297_), .I1(new_n24271_), .S(new_n11985_), .Z(new_n24298_));
  NOR2_X1    g21224(.A1(new_n24185_), .A2(pi0626), .ZN(new_n24299_));
  NOR2_X1    g21225(.A1(new_n12965_), .A2(pi0641), .ZN(new_n24300_));
  INV_X1     g21226(.I(new_n24300_), .ZN(new_n24301_));
  AOI21_X1   g21227(.A1(new_n24301_), .A2(pi1158), .B(new_n11994_), .ZN(new_n24302_));
  OAI21_X1   g21228(.A1(new_n24299_), .A2(new_n11989_), .B(new_n24302_), .ZN(new_n24303_));
  INV_X1     g21229(.I(new_n24303_), .ZN(new_n24304_));
  MUX2_X1    g21230(.I0(new_n24286_), .I1(new_n24277_), .S(new_n11969_), .Z(new_n24305_));
  NOR2_X1    g21231(.A1(new_n24305_), .A2(pi0789), .ZN(new_n24306_));
  NAND3_X1   g21232(.A1(new_n24297_), .A2(pi0789), .A3(new_n24306_), .ZN(new_n24307_));
  INV_X1     g21233(.I(new_n24306_), .ZN(new_n24308_));
  INV_X1     g21234(.I(new_n24273_), .ZN(new_n24309_));
  OAI21_X1   g21235(.A1(new_n24305_), .A2(new_n11967_), .B(new_n24309_), .ZN(new_n24310_));
  MUX2_X1    g21236(.I0(new_n24310_), .I1(new_n12965_), .S(new_n11869_), .Z(new_n24311_));
  NAND4_X1   g21237(.A1(new_n24294_), .A2(pi1159), .A3(new_n12965_), .A4(new_n24291_), .ZN(new_n24312_));
  OAI22_X1   g21238(.A1(new_n24289_), .A2(new_n24276_), .B1(new_n11869_), .B2(new_n12965_), .ZN(new_n24313_));
  AOI21_X1   g21239(.A1(new_n24313_), .A2(new_n24312_), .B(pi0648), .ZN(new_n24314_));
  AOI21_X1   g21240(.A1(pi0648), .A2(new_n24311_), .B(new_n24314_), .ZN(new_n24315_));
  OAI21_X1   g21241(.A1(new_n24315_), .A2(new_n11985_), .B(new_n24308_), .ZN(new_n24316_));
  NAND3_X1   g21242(.A1(new_n24307_), .A2(new_n24316_), .A3(new_n11994_), .ZN(new_n24317_));
  NOR2_X1    g21243(.A1(new_n11987_), .A2(pi0641), .ZN(new_n24318_));
  OAI21_X1   g21244(.A1(new_n24185_), .A2(new_n11994_), .B(new_n24318_), .ZN(new_n24319_));
  INV_X1     g21245(.I(new_n24319_), .ZN(new_n24320_));
  AOI22_X1   g21246(.A1(new_n24317_), .A2(new_n24320_), .B1(new_n24298_), .B2(new_n24304_), .ZN(new_n24321_));
  NOR2_X1    g21247(.A1(new_n14732_), .A2(new_n11986_), .ZN(new_n24322_));
  INV_X1     g21248(.I(new_n24322_), .ZN(new_n24323_));
  OAI21_X1   g21249(.A1(new_n24321_), .A2(new_n24323_), .B(new_n24212_), .ZN(new_n24324_));
  INV_X1     g21250(.I(pi0623), .ZN(new_n24325_));
  NOR2_X1    g21251(.A1(new_n12054_), .A2(new_n14727_), .ZN(new_n24326_));
  NOR2_X1    g21252(.A1(new_n24192_), .A2(new_n13716_), .ZN(new_n24327_));
  NOR2_X1    g21253(.A1(new_n14642_), .A2(new_n16809_), .ZN(new_n24328_));
  OAI21_X1   g21254(.A1(new_n24190_), .A2(pi0625), .B(new_n11893_), .ZN(new_n24329_));
  NAND2_X1   g21255(.A1(new_n24329_), .A2(pi0608), .ZN(new_n24330_));
  NOR2_X1    g21256(.A1(new_n23611_), .A2(new_n13659_), .ZN(new_n24331_));
  OAI21_X1   g21257(.A1(new_n24190_), .A2(new_n13659_), .B(new_n13657_), .ZN(new_n24332_));
  OAI21_X1   g21258(.A1(new_n23611_), .A2(pi0625), .B(new_n11893_), .ZN(new_n24333_));
  AOI22_X1   g21259(.A1(new_n24330_), .A2(new_n24331_), .B1(new_n24332_), .B2(new_n24333_), .ZN(new_n24334_));
  MUX2_X1    g21260(.I0(new_n24334_), .I1(new_n23611_), .S(new_n11891_), .Z(new_n24335_));
  AOI21_X1   g21261(.A1(pi0660), .A2(pi1155), .B(new_n11903_), .ZN(new_n24336_));
  NOR2_X1    g21262(.A1(pi0660), .A2(pi1155), .ZN(new_n24337_));
  OAI21_X1   g21263(.A1(new_n24192_), .A2(pi0609), .B(new_n24337_), .ZN(new_n24338_));
  NAND2_X1   g21264(.A1(new_n24335_), .A2(new_n11903_), .ZN(new_n24339_));
  AOI22_X1   g21265(.A1(new_n24339_), .A2(new_n24338_), .B1(new_n24335_), .B2(new_n24336_), .ZN(new_n24340_));
  NAND2_X1   g21266(.A1(new_n24335_), .A2(new_n11870_), .ZN(new_n24341_));
  OAI21_X1   g21267(.A1(new_n24340_), .A2(new_n11870_), .B(new_n24341_), .ZN(new_n24342_));
  NOR2_X1    g21268(.A1(new_n24192_), .A2(new_n13024_), .ZN(new_n24343_));
  NOR2_X1    g21269(.A1(new_n11949_), .A2(new_n11950_), .ZN(new_n24344_));
  OAI21_X1   g21270(.A1(new_n24343_), .A2(pi0618), .B(new_n24344_), .ZN(new_n24345_));
  NAND3_X1   g21271(.A1(new_n24345_), .A2(pi0618), .A3(new_n11969_), .ZN(new_n24346_));
  NOR4_X1    g21272(.A1(new_n24343_), .A2(pi0618), .A3(pi0627), .A4(pi1154), .ZN(new_n24347_));
  NAND3_X1   g21273(.A1(new_n24342_), .A2(new_n24346_), .A3(new_n24347_), .ZN(new_n24348_));
  AOI21_X1   g21274(.A1(new_n24342_), .A2(new_n11969_), .B(new_n16810_), .ZN(new_n24349_));
  AOI22_X1   g21275(.A1(new_n24349_), .A2(new_n24348_), .B1(new_n24327_), .B2(new_n24328_), .ZN(new_n24350_));
  OAI21_X1   g21276(.A1(new_n24350_), .A2(pi0788), .B(new_n14732_), .ZN(new_n24351_));
  NOR3_X1    g21277(.A1(new_n11989_), .A2(pi0626), .A3(pi1158), .ZN(new_n24352_));
  NOR3_X1    g21278(.A1(new_n24192_), .A2(new_n12013_), .A3(new_n13716_), .ZN(new_n24353_));
  NAND3_X1   g21279(.A1(new_n13095_), .A2(pi0626), .A3(new_n11986_), .ZN(new_n24354_));
  NOR3_X1    g21280(.A1(new_n24350_), .A2(new_n24352_), .A3(new_n24354_), .ZN(new_n24355_));
  AOI22_X1   g21281(.A1(new_n24355_), .A2(new_n24351_), .B1(new_n24193_), .B2(new_n24326_), .ZN(new_n24356_));
  NOR2_X1    g21282(.A1(new_n24325_), .A2(pi0207), .ZN(new_n24357_));
  INV_X1     g21283(.I(new_n17304_), .ZN(new_n24358_));
  AOI21_X1   g21284(.A1(new_n12965_), .A2(new_n12031_), .B(pi0629), .ZN(new_n24359_));
  OAI21_X1   g21285(.A1(new_n24187_), .A2(new_n12031_), .B(new_n24359_), .ZN(new_n24360_));
  AND2_X2    g21286(.A1(new_n24360_), .A2(new_n12026_), .Z(new_n24361_));
  NOR4_X1    g21287(.A1(new_n24155_), .A2(new_n24358_), .A3(new_n24209_), .A4(new_n24361_), .ZN(new_n24362_));
  NOR2_X1    g21288(.A1(new_n24184_), .A2(pi0619), .ZN(new_n24363_));
  NOR4_X1    g21289(.A1(new_n23621_), .A2(new_n3232_), .A3(new_n23616_), .A4(new_n23622_), .ZN(new_n24364_));
  INV_X1     g21290(.I(new_n24364_), .ZN(new_n24365_));
  NOR2_X1    g21291(.A1(new_n12965_), .A2(new_n13659_), .ZN(new_n24366_));
  INV_X1     g21292(.I(new_n24129_), .ZN(new_n24367_));
  AOI21_X1   g21293(.A1(new_n24365_), .A2(new_n12970_), .B(new_n24367_), .ZN(new_n24368_));
  NOR3_X1    g21294(.A1(new_n24365_), .A2(pi0625), .A3(new_n24129_), .ZN(new_n24369_));
  NOR4_X1    g21295(.A1(new_n24369_), .A2(new_n24368_), .A3(new_n12978_), .A4(new_n24366_), .ZN(new_n24370_));
  NAND2_X1   g21296(.A1(new_n24364_), .A2(pi0625), .ZN(new_n24371_));
  NAND2_X1   g21297(.A1(new_n24367_), .A2(new_n13434_), .ZN(new_n24372_));
  INV_X1     g21298(.I(new_n24372_), .ZN(new_n24373_));
  AOI21_X1   g21299(.A1(new_n24373_), .A2(new_n24371_), .B(new_n13657_), .ZN(new_n24374_));
  AOI21_X1   g21300(.A1(new_n24234_), .A2(new_n24374_), .B(new_n24370_), .ZN(new_n24375_));
  MUX2_X1    g21301(.I0(new_n24375_), .I1(new_n24365_), .S(new_n11891_), .Z(new_n24376_));
  NAND2_X1   g21302(.A1(new_n24376_), .A2(pi0609), .ZN(new_n24377_));
  NAND2_X1   g21303(.A1(new_n24179_), .A2(new_n11903_), .ZN(new_n24378_));
  NAND3_X1   g21304(.A1(new_n24377_), .A2(new_n11912_), .A3(new_n24378_), .ZN(new_n24379_));
  NAND3_X1   g21305(.A1(new_n24379_), .A2(pi0660), .A3(new_n24134_), .ZN(new_n24380_));
  AND3_X2    g21306(.A1(new_n24136_), .A2(new_n24232_), .A3(new_n24337_), .Z(new_n24381_));
  AOI21_X1   g21307(.A1(new_n24377_), .A2(new_n24381_), .B(new_n11870_), .ZN(new_n24382_));
  NAND2_X1   g21308(.A1(new_n24380_), .A2(new_n24382_), .ZN(new_n24383_));
  NAND2_X1   g21309(.A1(new_n24376_), .A2(new_n11870_), .ZN(new_n24384_));
  NAND2_X1   g21310(.A1(new_n24383_), .A2(new_n24384_), .ZN(new_n24385_));
  INV_X1     g21311(.I(new_n24385_), .ZN(new_n24386_));
  NAND3_X1   g21312(.A1(new_n24182_), .A2(pi0618), .A3(pi1154), .ZN(new_n24387_));
  NAND3_X1   g21313(.A1(new_n24141_), .A2(new_n11949_), .A3(new_n24387_), .ZN(new_n24388_));
  NAND4_X1   g21314(.A1(new_n24385_), .A2(pi0618), .A3(new_n11950_), .A4(new_n24181_), .ZN(new_n24389_));
  NAND2_X1   g21315(.A1(new_n24389_), .A2(new_n24143_), .ZN(new_n24390_));
  NAND2_X1   g21316(.A1(new_n24390_), .A2(new_n11949_), .ZN(new_n24391_));
  NAND2_X1   g21317(.A1(new_n24391_), .A2(new_n24388_), .ZN(new_n24392_));
  MUX2_X1    g21318(.I0(new_n24392_), .I1(new_n24385_), .S(new_n11969_), .Z(new_n24393_));
  AOI21_X1   g21319(.A1(new_n24393_), .A2(pi0619), .B(new_n24363_), .ZN(new_n24394_));
  OAI21_X1   g21320(.A1(new_n24152_), .A2(new_n11966_), .B(pi1159), .ZN(new_n24395_));
  NOR2_X1    g21321(.A1(new_n24386_), .A2(pi0781), .ZN(new_n24396_));
  AOI21_X1   g21322(.A1(new_n24392_), .A2(pi0781), .B(new_n24396_), .ZN(new_n24397_));
  MUX2_X1    g21323(.I0(new_n24397_), .I1(new_n24184_), .S(pi0619), .Z(new_n24398_));
  NOR2_X1    g21324(.A1(new_n24150_), .A2(pi0648), .ZN(new_n24399_));
  NOR4_X1    g21325(.A1(new_n24398_), .A2(pi0789), .A3(pi1159), .A4(new_n24399_), .ZN(new_n24400_));
  OAI21_X1   g21326(.A1(new_n24394_), .A2(new_n24395_), .B(new_n24400_), .ZN(new_n24401_));
  NOR2_X1    g21327(.A1(new_n24397_), .A2(pi0789), .ZN(new_n24402_));
  XNOR2_X1   g21328(.A1(pi0626), .A2(pi0641), .ZN(new_n24403_));
  NOR2_X1    g21329(.A1(new_n12003_), .A2(new_n24403_), .ZN(new_n24404_));
  INV_X1     g21330(.I(new_n24404_), .ZN(new_n24405_));
  NAND2_X1   g21331(.A1(new_n24301_), .A2(new_n11993_), .ZN(new_n24406_));
  AOI21_X1   g21332(.A1(new_n14396_), .A2(pi0641), .B(new_n16827_), .ZN(new_n24407_));
  XOR2_X1    g21333(.A1(new_n24406_), .A2(new_n24407_), .Z(new_n24408_));
  NOR2_X1    g21334(.A1(new_n24408_), .A2(new_n24185_), .ZN(new_n24409_));
  INV_X1     g21335(.I(new_n24409_), .ZN(new_n24410_));
  NOR2_X1    g21336(.A1(new_n24408_), .A2(new_n11989_), .ZN(new_n24411_));
  XOR2_X1    g21337(.A1(new_n24411_), .A2(new_n24406_), .Z(new_n24412_));
  AOI21_X1   g21338(.A1(new_n24412_), .A2(new_n24410_), .B(pi0788), .ZN(new_n24413_));
  OAI21_X1   g21339(.A1(new_n24154_), .A2(new_n24405_), .B(new_n24413_), .ZN(new_n24414_));
  NAND3_X1   g21340(.A1(new_n24414_), .A2(new_n11998_), .A3(new_n14732_), .ZN(new_n24415_));
  NOR2_X1    g21341(.A1(new_n24415_), .A2(new_n24402_), .ZN(new_n24416_));
  AOI21_X1   g21342(.A1(new_n24401_), .A2(new_n24416_), .B(new_n24362_), .ZN(new_n24417_));
  INV_X1     g21343(.I(new_n24417_), .ZN(new_n24418_));
  NAND2_X1   g21344(.A1(new_n24173_), .A2(new_n24174_), .ZN(new_n24419_));
  AOI21_X1   g21345(.A1(new_n24194_), .A2(new_n12026_), .B(new_n15220_), .ZN(new_n24420_));
  INV_X1     g21346(.I(new_n24420_), .ZN(new_n24421_));
  NAND4_X1   g21347(.A1(new_n24193_), .A2(new_n12031_), .A3(new_n12030_), .A4(new_n12026_), .ZN(new_n24422_));
  XOR2_X1    g21348(.A1(new_n24420_), .A2(new_n24422_), .Z(new_n24423_));
  NOR2_X1    g21349(.A1(new_n24423_), .A2(new_n12026_), .ZN(new_n24424_));
  NOR2_X1    g21350(.A1(new_n24424_), .A2(new_n24421_), .ZN(new_n24425_));
  NAND2_X1   g21351(.A1(new_n24424_), .A2(new_n24421_), .ZN(new_n24426_));
  INV_X1     g21352(.I(new_n24426_), .ZN(new_n24427_));
  NOR2_X1    g21353(.A1(new_n24423_), .A2(new_n24166_), .ZN(new_n24428_));
  NOR4_X1    g21354(.A1(new_n24427_), .A2(new_n11868_), .A3(new_n24425_), .A4(new_n24428_), .ZN(new_n24429_));
  NOR2_X1    g21355(.A1(new_n11934_), .A2(new_n11950_), .ZN(new_n24430_));
  NAND2_X1   g21356(.A1(new_n24160_), .A2(new_n24430_), .ZN(new_n24431_));
  INV_X1     g21357(.I(new_n24343_), .ZN(new_n24432_));
  NAND2_X1   g21358(.A1(new_n24432_), .A2(pi0618), .ZN(new_n24433_));
  AOI22_X1   g21359(.A1(new_n24433_), .A2(new_n11950_), .B1(new_n11949_), .B2(new_n24431_), .ZN(new_n24434_));
  NAND3_X1   g21360(.A1(new_n24191_), .A2(new_n11903_), .A3(pi1155), .ZN(new_n24435_));
  AOI21_X1   g21361(.A1(new_n11903_), .A2(new_n11912_), .B(pi0660), .ZN(new_n24436_));
  AND2_X2    g21362(.A1(new_n24159_), .A2(new_n24436_), .Z(new_n24437_));
  NAND3_X1   g21363(.A1(new_n24191_), .A2(pi0609), .A3(new_n11912_), .ZN(new_n24438_));
  NAND2_X1   g21364(.A1(pi0609), .A2(pi1155), .ZN(new_n24439_));
  OAI21_X1   g21365(.A1(new_n24159_), .A2(new_n24439_), .B(new_n11923_), .ZN(new_n24440_));
  AOI22_X1   g21366(.A1(new_n24438_), .A2(new_n24440_), .B1(new_n24435_), .B2(new_n24437_), .ZN(new_n24441_));
  NAND2_X1   g21367(.A1(new_n24441_), .A2(pi0785), .ZN(new_n24442_));
  MUX2_X1    g21368(.I0(new_n24442_), .I1(new_n24432_), .S(new_n11934_), .Z(new_n24443_));
  NOR2_X1    g21369(.A1(new_n24443_), .A2(new_n11950_), .ZN(new_n24444_));
  NOR2_X1    g21370(.A1(pi0618), .A2(pi1154), .ZN(new_n24445_));
  NOR4_X1    g21371(.A1(new_n24444_), .A2(pi0627), .A3(new_n24160_), .A4(new_n24445_), .ZN(new_n24446_));
  OAI21_X1   g21372(.A1(new_n24446_), .A2(new_n24434_), .B(pi0781), .ZN(new_n24447_));
  NOR4_X1    g21373(.A1(new_n24162_), .A2(pi0789), .A3(new_n11869_), .A4(new_n16807_), .ZN(new_n24448_));
  NOR2_X1    g21374(.A1(pi0619), .A2(pi0648), .ZN(new_n24449_));
  NAND4_X1   g21375(.A1(new_n24327_), .A2(new_n11869_), .A3(new_n24449_), .A4(new_n24162_), .ZN(new_n24450_));
  NOR2_X1    g21376(.A1(new_n24450_), .A2(new_n24448_), .ZN(new_n24451_));
  INV_X1     g21377(.I(new_n24451_), .ZN(new_n24452_));
  INV_X1     g21378(.I(new_n24442_), .ZN(new_n24453_));
  AOI21_X1   g21379(.A1(new_n12012_), .A2(new_n16809_), .B(new_n24452_), .ZN(new_n24454_));
  AOI21_X1   g21380(.A1(new_n11934_), .A2(new_n11949_), .B(new_n11969_), .ZN(new_n24455_));
  NOR3_X1    g21381(.A1(new_n24454_), .A2(new_n24453_), .A3(new_n24455_), .ZN(new_n24456_));
  AOI22_X1   g21382(.A1(new_n24447_), .A2(new_n24456_), .B1(pi0789), .B2(new_n24452_), .ZN(new_n24457_));
  NOR4_X1    g21383(.A1(new_n24163_), .A2(pi0626), .A3(new_n11989_), .A4(pi1158), .ZN(new_n24458_));
  NOR2_X1    g21384(.A1(new_n24353_), .A2(pi0626), .ZN(new_n24459_));
  NAND4_X1   g21385(.A1(new_n24457_), .A2(pi0626), .A3(pi0641), .A4(new_n24459_), .ZN(new_n24460_));
  NOR4_X1    g21386(.A1(new_n24164_), .A2(new_n11994_), .A3(pi0641), .A4(pi1158), .ZN(new_n24461_));
  AOI22_X1   g21387(.A1(new_n24460_), .A2(new_n24461_), .B1(new_n24457_), .B2(new_n24458_), .ZN(new_n24462_));
  OR2_X2     g21388(.A1(new_n24462_), .A2(new_n11986_), .Z(new_n24463_));
  AOI21_X1   g21389(.A1(new_n24457_), .A2(new_n11986_), .B(new_n14731_), .ZN(new_n24464_));
  AOI21_X1   g21390(.A1(new_n24463_), .A2(new_n24464_), .B(new_n24429_), .ZN(new_n24465_));
  INV_X1     g21391(.I(new_n24465_), .ZN(new_n24466_));
  NOR2_X1    g21392(.A1(new_n24325_), .A2(pi0710), .ZN(new_n24467_));
  OAI21_X1   g21393(.A1(new_n24466_), .A2(new_n8087_), .B(new_n24467_), .ZN(new_n24468_));
  AOI21_X1   g21394(.A1(new_n24419_), .A2(new_n14726_), .B(new_n24468_), .ZN(new_n24469_));
  OAI21_X1   g21395(.A1(pi0207), .A2(new_n24418_), .B(new_n24469_), .ZN(new_n24470_));
  AOI21_X1   g21396(.A1(new_n24324_), .A2(new_n24357_), .B(new_n24470_), .ZN(new_n24471_));
  NOR2_X1    g21397(.A1(new_n24471_), .A2(new_n24206_), .ZN(new_n24472_));
  NAND3_X1   g21398(.A1(new_n24172_), .A2(new_n12061_), .A3(new_n12049_), .ZN(new_n24473_));
  MUX2_X1    g21399(.I0(new_n24473_), .I1(new_n24200_), .S(new_n12048_), .Z(new_n24474_));
  INV_X1     g21400(.I(new_n24474_), .ZN(new_n24475_));
  AOI21_X1   g21401(.A1(new_n24475_), .A2(pi0644), .B(pi0715), .ZN(new_n24476_));
  NAND2_X1   g21402(.A1(new_n24173_), .A2(new_n12092_), .ZN(new_n24477_));
  OAI21_X1   g21403(.A1(new_n12092_), .A2(new_n24172_), .B(new_n24477_), .ZN(new_n24478_));
  NOR2_X1    g21404(.A1(pi0644), .A2(pi0715), .ZN(new_n24479_));
  NAND2_X1   g21405(.A1(new_n24478_), .A2(new_n24479_), .ZN(new_n24480_));
  NAND2_X1   g21406(.A1(new_n24480_), .A2(new_n24041_), .ZN(new_n24481_));
  NOR2_X1    g21407(.A1(new_n24481_), .A2(new_n24476_), .ZN(new_n24482_));
  AOI21_X1   g21408(.A1(new_n24475_), .A2(new_n12082_), .B(new_n12099_), .ZN(new_n24483_));
  NOR3_X1    g21409(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n24484_));
  NAND2_X1   g21410(.A1(new_n24478_), .A2(new_n24484_), .ZN(new_n24485_));
  NAND2_X1   g21411(.A1(new_n24485_), .A2(pi0644), .ZN(new_n24486_));
  NOR2_X1    g21412(.A1(new_n24486_), .A2(new_n24483_), .ZN(new_n24487_));
  NOR3_X1    g21413(.A1(new_n24472_), .A2(new_n24482_), .A3(new_n24487_), .ZN(new_n24488_));
  AOI21_X1   g21414(.A1(new_n24488_), .A2(pi0790), .B(new_n24472_), .ZN(new_n24489_));
  NAND3_X1   g21415(.A1(new_n24488_), .A2(pi0790), .A3(new_n24472_), .ZN(new_n24490_));
  NAND2_X1   g21416(.A1(new_n24490_), .A2(new_n6845_), .ZN(new_n24491_));
  OAI22_X1   g21417(.A1(new_n24491_), .A2(new_n24489_), .B1(pi0207), .B2(new_n6845_), .ZN(po0364));
  AOI21_X1   g21418(.A1(new_n24158_), .A2(new_n24168_), .B(new_n8088_), .ZN(new_n24493_));
  NAND2_X1   g21419(.A1(new_n24493_), .A2(pi0607), .ZN(new_n24494_));
  NOR2_X1    g21420(.A1(new_n12965_), .A2(pi0208), .ZN(new_n24495_));
  INV_X1     g21421(.I(new_n24495_), .ZN(new_n24496_));
  OAI21_X1   g21422(.A1(pi0607), .A2(new_n24496_), .B(new_n24494_), .ZN(new_n24497_));
  INV_X1     g21423(.I(pi0638), .ZN(new_n24498_));
  NOR2_X1    g21424(.A1(new_n24196_), .A2(new_n8088_), .ZN(new_n24499_));
  AOI21_X1   g21425(.A1(new_n24189_), .A2(new_n8088_), .B(new_n24499_), .ZN(new_n24500_));
  NOR2_X1    g21426(.A1(new_n24500_), .A2(new_n24498_), .ZN(new_n24501_));
  AOI21_X1   g21427(.A1(new_n24498_), .A2(new_n24495_), .B(new_n24501_), .ZN(new_n24502_));
  NAND2_X1   g21428(.A1(new_n24502_), .A2(pi0647), .ZN(new_n24503_));
  AOI21_X1   g21429(.A1(new_n24496_), .A2(new_n12061_), .B(pi1157), .ZN(new_n24504_));
  AOI21_X1   g21430(.A1(new_n24503_), .A2(new_n24504_), .B(pi0630), .ZN(new_n24505_));
  AOI21_X1   g21431(.A1(new_n24495_), .A2(pi0647), .B(pi1157), .ZN(new_n24506_));
  AND3_X2    g21432(.A1(new_n24503_), .A2(pi0630), .A3(new_n24506_), .Z(new_n24507_));
  NOR4_X1    g21433(.A1(new_n24497_), .A2(new_n15183_), .A3(new_n24505_), .A4(new_n24507_), .ZN(new_n24508_));
  INV_X1     g21434(.I(pi0607), .ZN(new_n24509_));
  NOR2_X1    g21435(.A1(new_n24509_), .A2(pi0208), .ZN(new_n24510_));
  NAND2_X1   g21436(.A1(new_n24497_), .A2(new_n24498_), .ZN(new_n24511_));
  NOR2_X1    g21437(.A1(new_n24509_), .A2(pi0638), .ZN(new_n24512_));
  OAI21_X1   g21438(.A1(new_n24466_), .A2(new_n8088_), .B(new_n24512_), .ZN(new_n24513_));
  AOI21_X1   g21439(.A1(new_n24511_), .A2(new_n14726_), .B(new_n24513_), .ZN(new_n24514_));
  OAI21_X1   g21440(.A1(pi0208), .A2(new_n24418_), .B(new_n24514_), .ZN(new_n24515_));
  AOI21_X1   g21441(.A1(new_n24324_), .A2(new_n24510_), .B(new_n24515_), .ZN(new_n24516_));
  NOR2_X1    g21442(.A1(new_n24516_), .A2(new_n24508_), .ZN(new_n24517_));
  NAND3_X1   g21443(.A1(new_n24496_), .A2(new_n12061_), .A3(new_n12049_), .ZN(new_n24518_));
  MUX2_X1    g21444(.I0(new_n24518_), .I1(new_n24502_), .S(new_n12048_), .Z(new_n24519_));
  INV_X1     g21445(.I(new_n24519_), .ZN(new_n24520_));
  AOI21_X1   g21446(.A1(new_n24520_), .A2(pi0644), .B(pi0715), .ZN(new_n24521_));
  NAND2_X1   g21447(.A1(new_n24497_), .A2(new_n12092_), .ZN(new_n24522_));
  OAI21_X1   g21448(.A1(new_n12092_), .A2(new_n24496_), .B(new_n24522_), .ZN(new_n24523_));
  NOR2_X1    g21449(.A1(pi0644), .A2(pi0715), .ZN(new_n24524_));
  NAND2_X1   g21450(.A1(new_n24523_), .A2(new_n24524_), .ZN(new_n24525_));
  NAND2_X1   g21451(.A1(new_n24525_), .A2(new_n24041_), .ZN(new_n24526_));
  NOR2_X1    g21452(.A1(new_n24526_), .A2(new_n24521_), .ZN(new_n24527_));
  AOI21_X1   g21453(.A1(new_n24520_), .A2(new_n12082_), .B(new_n12099_), .ZN(new_n24528_));
  NOR3_X1    g21454(.A1(new_n12082_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n24529_));
  NAND2_X1   g21455(.A1(new_n24523_), .A2(new_n24529_), .ZN(new_n24530_));
  NAND2_X1   g21456(.A1(new_n24530_), .A2(pi0644), .ZN(new_n24531_));
  NOR2_X1    g21457(.A1(new_n24531_), .A2(new_n24528_), .ZN(new_n24532_));
  NOR3_X1    g21458(.A1(new_n24517_), .A2(new_n24527_), .A3(new_n24532_), .ZN(new_n24533_));
  AOI21_X1   g21459(.A1(new_n24533_), .A2(pi0790), .B(new_n24517_), .ZN(new_n24534_));
  NAND3_X1   g21460(.A1(new_n24533_), .A2(pi0790), .A3(new_n24517_), .ZN(new_n24535_));
  NAND2_X1   g21461(.A1(new_n24535_), .A2(new_n6845_), .ZN(new_n24536_));
  OAI22_X1   g21462(.A1(new_n24536_), .A2(new_n24534_), .B1(pi0208), .B2(new_n6845_), .ZN(po0365));
  NOR4_X1    g21463(.A1(new_n24465_), .A2(new_n12061_), .A3(pi1157), .A4(new_n24167_), .ZN(new_n24538_));
  OAI21_X1   g21464(.A1(new_n24196_), .A2(pi0647), .B(new_n12049_), .ZN(new_n24539_));
  NAND2_X1   g21465(.A1(new_n24539_), .A2(pi0630), .ZN(new_n24540_));
  NOR3_X1    g21466(.A1(new_n24168_), .A2(new_n12061_), .A3(new_n12049_), .ZN(new_n24541_));
  AOI21_X1   g21467(.A1(new_n24195_), .A2(new_n13736_), .B(pi0630), .ZN(new_n24542_));
  OAI22_X1   g21468(.A1(new_n24538_), .A2(new_n24540_), .B1(new_n24541_), .B2(new_n24542_), .ZN(new_n24543_));
  MUX2_X1    g21469(.I0(new_n24543_), .I1(new_n24465_), .S(new_n12048_), .Z(new_n24544_));
  NOR2_X1    g21470(.A1(new_n24166_), .A2(new_n16841_), .ZN(new_n24545_));
  NAND3_X1   g21471(.A1(new_n24545_), .A2(new_n12081_), .A3(new_n12095_), .ZN(new_n24546_));
  INV_X1     g21472(.I(new_n13748_), .ZN(new_n24547_));
  NOR2_X1    g21473(.A1(new_n24196_), .A2(new_n24547_), .ZN(new_n24548_));
  NAND3_X1   g21474(.A1(new_n24546_), .A2(pi0644), .A3(new_n12099_), .ZN(new_n24549_));
  NOR4_X1    g21475(.A1(new_n24548_), .A2(pi0644), .A3(pi0715), .A4(pi1160), .ZN(new_n24550_));
  NAND3_X1   g21476(.A1(new_n24545_), .A2(new_n12082_), .A3(pi0715), .ZN(new_n24551_));
  NAND2_X1   g21477(.A1(new_n24551_), .A2(new_n24550_), .ZN(new_n24552_));
  AOI21_X1   g21478(.A1(new_n24549_), .A2(new_n24552_), .B(new_n24544_), .ZN(new_n24553_));
  NOR2_X1    g21479(.A1(new_n6845_), .A2(new_n11867_), .ZN(new_n24554_));
  NAND2_X1   g21480(.A1(new_n24553_), .A2(new_n24554_), .ZN(new_n24555_));
  INV_X1     g21481(.I(pi0622), .ZN(new_n24556_));
  INV_X1     g21482(.I(pi0639), .ZN(new_n24557_));
  XOR2_X1    g21483(.A1(pi0647), .A2(pi1157), .Z(new_n24558_));
  NOR2_X1    g21484(.A1(new_n12092_), .A2(new_n24558_), .ZN(new_n24559_));
  AOI22_X1   g21485(.A1(new_n24356_), .A2(new_n14726_), .B1(new_n24195_), .B2(new_n24559_), .ZN(new_n24560_));
  NAND2_X1   g21486(.A1(new_n24560_), .A2(new_n24550_), .ZN(new_n24561_));
  NOR2_X1    g21487(.A1(new_n24548_), .A2(pi0644), .ZN(new_n24562_));
  AND2_X2    g21488(.A1(new_n24560_), .A2(pi0644), .Z(new_n24563_));
  NOR4_X1    g21489(.A1(new_n24563_), .A2(new_n12099_), .A3(new_n12081_), .A4(new_n24562_), .ZN(new_n24564_));
  INV_X1     g21490(.I(new_n24564_), .ZN(new_n24565_));
  OAI21_X1   g21491(.A1(new_n24560_), .A2(po1038), .B(new_n11867_), .ZN(new_n24566_));
  AOI21_X1   g21492(.A1(new_n24565_), .A2(new_n24561_), .B(new_n24566_), .ZN(new_n24567_));
  NOR2_X1    g21493(.A1(new_n12082_), .A2(pi1160), .ZN(new_n24568_));
  NOR2_X1    g21494(.A1(new_n12081_), .A2(pi0644), .ZN(new_n24569_));
  OAI21_X1   g21495(.A1(new_n24568_), .A2(new_n24569_), .B(pi0790), .ZN(new_n24570_));
  NAND3_X1   g21496(.A1(new_n24545_), .A2(new_n6845_), .A3(new_n24570_), .ZN(new_n24571_));
  NOR3_X1    g21497(.A1(new_n24556_), .A2(new_n24557_), .A3(pi0209), .ZN(new_n24573_));
  NAND2_X1   g21498(.A1(new_n24555_), .A2(new_n24573_), .ZN(new_n24574_));
  NAND3_X1   g21499(.A1(new_n24189_), .A2(new_n12061_), .A3(new_n12965_), .ZN(new_n24575_));
  INV_X1     g21500(.I(new_n24189_), .ZN(new_n24576_));
  OAI21_X1   g21501(.A1(pi0647), .A2(new_n12965_), .B(new_n24576_), .ZN(new_n24577_));
  NAND3_X1   g21502(.A1(new_n24577_), .A2(new_n12060_), .A3(new_n24575_), .ZN(new_n24578_));
  AOI21_X1   g21503(.A1(new_n12061_), .A2(new_n14396_), .B(new_n24578_), .ZN(new_n24579_));
  AOI21_X1   g21504(.A1(new_n12965_), .A2(pi0647), .B(new_n13743_), .ZN(new_n24580_));
  OAI21_X1   g21505(.A1(new_n24189_), .A2(pi0647), .B(new_n24580_), .ZN(new_n24581_));
  INV_X1     g21506(.I(new_n24581_), .ZN(new_n24582_));
  NAND3_X1   g21507(.A1(new_n12048_), .A2(pi0647), .A3(pi1157), .ZN(new_n24583_));
  NOR3_X1    g21508(.A1(new_n24579_), .A2(new_n24582_), .A3(new_n24583_), .ZN(new_n24584_));
  MUX2_X1    g21509(.I0(new_n24315_), .I1(new_n24305_), .S(new_n11985_), .Z(new_n24585_));
  NOR2_X1    g21510(.A1(new_n24585_), .A2(new_n24303_), .ZN(new_n24586_));
  AOI21_X1   g21511(.A1(new_n24298_), .A2(new_n11994_), .B(new_n24319_), .ZN(new_n24587_));
  OAI21_X1   g21512(.A1(new_n24587_), .A2(new_n24586_), .B(new_n24322_), .ZN(new_n24588_));
  AOI21_X1   g21513(.A1(new_n24588_), .A2(new_n24212_), .B(new_n14725_), .ZN(new_n24589_));
  NOR2_X1    g21514(.A1(new_n14396_), .A2(new_n13748_), .ZN(new_n24590_));
  AOI21_X1   g21515(.A1(new_n24576_), .A2(new_n13748_), .B(new_n24590_), .ZN(new_n24591_));
  AOI21_X1   g21516(.A1(new_n24591_), .A2(new_n12082_), .B(new_n12099_), .ZN(new_n24592_));
  OAI21_X1   g21517(.A1(new_n14396_), .A2(pi0715), .B(pi1160), .ZN(new_n24593_));
  NAND2_X1   g21518(.A1(new_n24593_), .A2(pi0644), .ZN(new_n24594_));
  NOR4_X1    g21519(.A1(new_n24589_), .A2(new_n24584_), .A3(new_n24592_), .A4(new_n24594_), .ZN(new_n24595_));
  AOI21_X1   g21520(.A1(new_n24324_), .A2(new_n14726_), .B(new_n24584_), .ZN(new_n24596_));
  NAND2_X1   g21521(.A1(new_n24591_), .A2(pi0644), .ZN(new_n24597_));
  NAND2_X1   g21522(.A1(new_n24597_), .A2(new_n12099_), .ZN(new_n24598_));
  AOI21_X1   g21523(.A1(new_n12965_), .A2(pi0715), .B(pi1160), .ZN(new_n24599_));
  NOR2_X1    g21524(.A1(new_n24598_), .A2(new_n24599_), .ZN(new_n24600_));
  INV_X1     g21525(.I(new_n24600_), .ZN(new_n24601_));
  AOI21_X1   g21526(.A1(new_n24596_), .A2(new_n12082_), .B(new_n24601_), .ZN(new_n24602_));
  NOR2_X1    g21527(.A1(new_n6845_), .A2(new_n11867_), .ZN(new_n24603_));
  OAI21_X1   g21528(.A1(new_n24602_), .A2(new_n24595_), .B(new_n24603_), .ZN(new_n24604_));
  NAND2_X1   g21529(.A1(new_n12902_), .A2(new_n7832_), .ZN(new_n24605_));
  AOI21_X1   g21530(.A1(new_n24557_), .A2(new_n24605_), .B(new_n24604_), .ZN(new_n24606_));
  NOR2_X1    g21531(.A1(new_n24592_), .A2(new_n24594_), .ZN(new_n24607_));
  NAND2_X1   g21532(.A1(new_n24596_), .A2(new_n24607_), .ZN(new_n24608_));
  INV_X1     g21533(.I(new_n24212_), .ZN(new_n24609_));
  NOR3_X1    g21534(.A1(new_n24315_), .A2(new_n11985_), .A3(new_n24308_), .ZN(new_n24610_));
  AOI21_X1   g21535(.A1(new_n24297_), .A2(pi0789), .B(new_n24306_), .ZN(new_n24611_));
  NOR3_X1    g21536(.A1(new_n24611_), .A2(new_n24610_), .A3(pi0626), .ZN(new_n24612_));
  OAI22_X1   g21537(.A1(new_n24612_), .A2(new_n24319_), .B1(new_n24585_), .B2(new_n24303_), .ZN(new_n24613_));
  AOI21_X1   g21538(.A1(new_n24613_), .A2(new_n24322_), .B(new_n24609_), .ZN(new_n24614_));
  INV_X1     g21539(.I(new_n24584_), .ZN(new_n24615_));
  OAI21_X1   g21540(.A1(new_n24614_), .A2(new_n14725_), .B(new_n24615_), .ZN(new_n24616_));
  OAI21_X1   g21541(.A1(new_n24616_), .A2(pi0644), .B(new_n24600_), .ZN(new_n24617_));
  INV_X1     g21542(.I(new_n24603_), .ZN(new_n24618_));
  AOI21_X1   g21543(.A1(new_n24617_), .A2(new_n24608_), .B(new_n24618_), .ZN(new_n24619_));
  NOR3_X1    g21544(.A1(new_n24619_), .A2(pi0639), .A3(new_n24605_), .ZN(new_n24620_));
  NAND2_X1   g21545(.A1(new_n24578_), .A2(pi1157), .ZN(new_n24621_));
  AOI21_X1   g21546(.A1(new_n24158_), .A2(new_n15076_), .B(new_n24582_), .ZN(new_n24622_));
  NAND2_X1   g21547(.A1(new_n24622_), .A2(new_n24621_), .ZN(new_n24623_));
  AOI22_X1   g21548(.A1(new_n24417_), .A2(new_n14726_), .B1(pi0787), .B2(new_n24623_), .ZN(new_n24624_));
  NOR2_X1    g21549(.A1(new_n14396_), .A2(pi0644), .ZN(new_n24625_));
  OR2_X2     g21550(.A1(new_n24158_), .A2(new_n12091_), .Z(new_n24626_));
  OAI21_X1   g21551(.A1(new_n12092_), .A2(new_n14396_), .B(new_n24626_), .ZN(new_n24627_));
  AOI21_X1   g21552(.A1(new_n24627_), .A2(pi0644), .B(new_n24625_), .ZN(new_n24628_));
  OAI21_X1   g21553(.A1(new_n24628_), .A2(pi0715), .B(pi1160), .ZN(new_n24629_));
  NOR2_X1    g21554(.A1(new_n12082_), .A2(pi0715), .ZN(new_n24630_));
  NAND2_X1   g21555(.A1(new_n24629_), .A2(new_n24630_), .ZN(new_n24631_));
  NOR2_X1    g21556(.A1(new_n24624_), .A2(pi0644), .ZN(new_n24632_));
  NOR2_X1    g21557(.A1(new_n14396_), .A2(new_n12082_), .ZN(new_n24633_));
  AOI21_X1   g21558(.A1(new_n24627_), .A2(new_n12082_), .B(new_n24633_), .ZN(new_n24634_));
  NAND3_X1   g21559(.A1(new_n24597_), .A2(new_n12099_), .A3(pi1160), .ZN(new_n24635_));
  OAI22_X1   g21560(.A1(new_n24631_), .A2(new_n24624_), .B1(new_n24632_), .B2(new_n24635_), .ZN(new_n24636_));
  NOR2_X1    g21561(.A1(new_n6845_), .A2(new_n11867_), .ZN(new_n24637_));
  AOI21_X1   g21562(.A1(new_n24636_), .A2(new_n24637_), .B(new_n24557_), .ZN(new_n24638_));
  INV_X1     g21563(.I(new_n24627_), .ZN(new_n24639_));
  NAND4_X1   g21564(.A1(new_n24628_), .A2(new_n24634_), .A3(new_n11867_), .A4(pi1160), .ZN(new_n24640_));
  NAND2_X1   g21565(.A1(new_n24640_), .A2(new_n6845_), .ZN(new_n24641_));
  NAND3_X1   g21566(.A1(new_n24641_), .A2(new_n11867_), .A3(new_n24639_), .ZN(new_n24642_));
  AND2_X2    g21567(.A1(new_n24642_), .A2(new_n24557_), .Z(new_n24643_));
  OAI21_X1   g21568(.A1(new_n24643_), .A2(new_n24638_), .B(new_n24556_), .ZN(new_n24644_));
  NOR3_X1    g21569(.A1(new_n24606_), .A2(new_n24620_), .A3(new_n24644_), .ZN(new_n24645_));
  OAI21_X1   g21570(.A1(new_n24645_), .A2(pi0209), .B(new_n24574_), .ZN(po0366));
  NAND3_X1   g21571(.A1(new_n5473_), .A2(pi0634), .A3(pi0907), .ZN(new_n24647_));
  NAND2_X1   g21572(.A1(pi0633), .A2(pi0947), .ZN(new_n24648_));
  XNOR2_X1   g21573(.A1(new_n24647_), .A2(new_n24648_), .ZN(new_n24649_));
  NOR4_X1    g21574(.A1(new_n13368_), .A2(pi0038), .A3(pi0210), .A4(new_n24649_), .ZN(new_n24650_));
  OAI21_X1   g21575(.A1(new_n12809_), .A2(new_n2631_), .B(new_n5091_), .ZN(new_n24651_));
  OAI21_X1   g21576(.A1(po1101), .A2(new_n12132_), .B(new_n2631_), .ZN(new_n24652_));
  AOI21_X1   g21577(.A1(new_n12231_), .A2(po1101), .B(new_n24652_), .ZN(new_n24653_));
  AOI21_X1   g21578(.A1(new_n24653_), .A2(new_n5090_), .B(pi0907), .ZN(new_n24654_));
  NOR2_X1    g21579(.A1(new_n12156_), .A2(pi0210), .ZN(new_n24655_));
  AOI21_X1   g21580(.A1(new_n23202_), .A2(new_n12156_), .B(new_n24655_), .ZN(new_n24656_));
  INV_X1     g21581(.I(new_n24656_), .ZN(new_n24657_));
  NOR2_X1    g21582(.A1(new_n12132_), .A2(pi0210), .ZN(new_n24658_));
  AOI21_X1   g21583(.A1(new_n23202_), .A2(new_n12132_), .B(new_n24658_), .ZN(new_n24659_));
  INV_X1     g21584(.I(new_n24659_), .ZN(new_n24660_));
  NOR3_X1    g21585(.A1(new_n6446_), .A2(pi0947), .A3(new_n24660_), .ZN(new_n24661_));
  INV_X1     g21586(.I(new_n24661_), .ZN(new_n24662_));
  NOR2_X1    g21587(.A1(new_n24657_), .A2(new_n24662_), .ZN(new_n24663_));
  AOI21_X1   g21588(.A1(new_n23318_), .A2(new_n12156_), .B(new_n24655_), .ZN(new_n24664_));
  AOI21_X1   g21589(.A1(new_n23318_), .A2(new_n12132_), .B(new_n24658_), .ZN(new_n24665_));
  INV_X1     g21590(.I(new_n24665_), .ZN(new_n24666_));
  NOR3_X1    g21591(.A1(new_n6446_), .A2(pi0907), .A3(new_n24666_), .ZN(new_n24667_));
  AOI21_X1   g21592(.A1(new_n24664_), .A2(new_n24667_), .B(pi0947), .ZN(new_n24668_));
  OAI21_X1   g21593(.A1(new_n24663_), .A2(new_n3284_), .B(new_n24668_), .ZN(new_n24669_));
  AOI21_X1   g21594(.A1(new_n24651_), .A2(new_n24654_), .B(new_n24669_), .ZN(new_n24670_));
  NOR2_X1    g21595(.A1(new_n12242_), .A2(pi0210), .ZN(new_n24671_));
  INV_X1     g21596(.I(new_n24671_), .ZN(new_n24672_));
  OAI21_X1   g21597(.A1(pi0633), .A2(new_n12262_), .B(new_n24672_), .ZN(new_n24673_));
  NOR2_X1    g21598(.A1(new_n24673_), .A2(new_n24662_), .ZN(new_n24674_));
  AOI21_X1   g21599(.A1(new_n23318_), .A2(new_n12242_), .B(new_n24671_), .ZN(new_n24675_));
  NAND2_X1   g21600(.A1(new_n24675_), .A2(new_n24667_), .ZN(new_n24676_));
  AOI21_X1   g21601(.A1(new_n12725_), .A2(po1101), .B(new_n24652_), .ZN(new_n24677_));
  NOR3_X1    g21602(.A1(new_n6446_), .A2(new_n2926_), .A3(new_n12680_), .ZN(new_n24678_));
  NOR3_X1    g21603(.A1(new_n24678_), .A2(new_n12242_), .A3(new_n2631_), .ZN(new_n24679_));
  NAND3_X1   g21604(.A1(new_n24677_), .A2(pi0907), .A3(new_n5090_), .ZN(new_n24680_));
  AOI21_X1   g21605(.A1(new_n24680_), .A2(new_n24676_), .B(pi0947), .ZN(new_n24681_));
  INV_X1     g21606(.I(new_n4905_), .ZN(new_n24682_));
  INV_X1     g21607(.I(new_n24658_), .ZN(new_n24683_));
  OAI21_X1   g21608(.A1(new_n24649_), .A2(new_n12133_), .B(new_n24683_), .ZN(new_n24684_));
  AOI21_X1   g21609(.A1(new_n24684_), .A2(new_n3284_), .B(new_n24682_), .ZN(new_n24685_));
  OAI21_X1   g21610(.A1(new_n24681_), .A2(new_n24674_), .B(new_n24685_), .ZN(new_n24686_));
  AOI21_X1   g21611(.A1(new_n5107_), .A2(new_n24660_), .B(new_n5473_), .ZN(new_n24690_));
  NOR2_X1    g21612(.A1(new_n24660_), .A2(new_n5109_), .ZN(new_n24691_));
  NOR3_X1    g21613(.A1(new_n24690_), .A2(new_n5107_), .A3(new_n24691_), .ZN(new_n24692_));
  NAND3_X1   g21614(.A1(new_n24684_), .A2(pi0223), .A3(new_n2614_), .ZN(new_n24701_));
  INV_X1     g21615(.I(new_n24675_), .ZN(new_n24702_));
  NAND3_X1   g21616(.A1(new_n24702_), .A2(new_n5143_), .A3(new_n24665_), .ZN(new_n24703_));
  OAI21_X1   g21617(.A1(new_n24702_), .A2(new_n6548_), .B(new_n24666_), .ZN(new_n24704_));
  AOI21_X1   g21618(.A1(new_n24704_), .A2(new_n24703_), .B(new_n15305_), .ZN(new_n24705_));
  NAND2_X1   g21619(.A1(new_n24677_), .A2(new_n15305_), .ZN(new_n24706_));
  OAI21_X1   g21620(.A1(new_n24673_), .A2(new_n5108_), .B(new_n24692_), .ZN(new_n24707_));
  NAND3_X1   g21621(.A1(new_n24707_), .A2(new_n5473_), .A3(new_n24706_), .ZN(new_n24708_));
  INV_X1     g21622(.I(new_n24676_), .ZN(new_n24709_));
  OAI21_X1   g21623(.A1(new_n24709_), .A2(new_n24679_), .B(new_n5473_), .ZN(new_n24710_));
  NOR2_X1    g21624(.A1(new_n24674_), .A2(new_n5141_), .ZN(new_n24711_));
  NAND2_X1   g21625(.A1(new_n6460_), .A2(new_n2604_), .ZN(new_n24712_));
  AOI21_X1   g21626(.A1(new_n24710_), .A2(new_n24711_), .B(new_n24712_), .ZN(new_n24713_));
  OAI21_X1   g21627(.A1(new_n24705_), .A2(new_n24708_), .B(new_n24713_), .ZN(new_n24714_));
  NAND3_X1   g21628(.A1(new_n24714_), .A2(new_n2587_), .A3(new_n24701_), .ZN(new_n24715_));
  OAI21_X1   g21629(.A1(new_n24670_), .A2(new_n24686_), .B(new_n24715_), .ZN(new_n24716_));
  INV_X1     g21630(.I(new_n24649_), .ZN(new_n24717_));
  NAND3_X1   g21631(.A1(new_n12646_), .A2(pi0210), .A3(new_n24717_), .ZN(new_n24718_));
  OAI21_X1   g21632(.A1(new_n12584_), .A2(pi0210), .B(new_n24649_), .ZN(new_n24719_));
  NOR2_X1    g21633(.A1(pi0039), .A2(pi0299), .ZN(new_n24722_));
  NAND3_X1   g21634(.A1(new_n24718_), .A2(new_n24719_), .A3(new_n24722_), .ZN(new_n24723_));
  AOI21_X1   g21635(.A1(new_n24723_), .A2(new_n3172_), .B(pi0039), .ZN(new_n24724_));
  AOI21_X1   g21636(.A1(new_n24724_), .A2(new_n24716_), .B(new_n24650_), .ZN(new_n24725_));
  MUX2_X1    g21637(.I0(new_n24725_), .I1(pi0210), .S(new_n7833_), .Z(po0367));
  NOR2_X1    g21638(.A1(new_n15444_), .A2(new_n3232_), .ZN(new_n24727_));
  INV_X1     g21639(.I(new_n24727_), .ZN(new_n24728_));
  AOI21_X1   g21640(.A1(new_n23937_), .A2(new_n14396_), .B(new_n24728_), .ZN(new_n24729_));
  NAND3_X1   g21641(.A1(new_n24728_), .A2(new_n23937_), .A3(new_n12965_), .ZN(new_n24730_));
  NOR3_X1    g21642(.A1(new_n3231_), .A2(new_n23937_), .A3(pi0643), .ZN(new_n24731_));
  NOR4_X1    g21643(.A1(new_n24731_), .A2(new_n8077_), .A3(pi0643), .A4(po1038), .ZN(new_n24732_));
  NAND2_X1   g21644(.A1(new_n24730_), .A2(new_n24732_), .ZN(new_n24733_));
  NAND2_X1   g21645(.A1(new_n15804_), .A2(new_n3231_), .ZN(new_n24734_));
  NOR2_X1    g21646(.A1(new_n15802_), .A2(new_n3232_), .ZN(new_n24735_));
  OAI21_X1   g21647(.A1(new_n24735_), .A2(new_n24734_), .B(pi0606), .ZN(new_n24736_));
  NOR2_X1    g21648(.A1(new_n24736_), .A2(new_n23901_), .ZN(new_n24737_));
  NAND2_X1   g21649(.A1(new_n23901_), .A2(pi0606), .ZN(new_n24738_));
  NOR2_X1    g21650(.A1(new_n15461_), .A2(new_n3232_), .ZN(new_n24739_));
  INV_X1     g21651(.I(new_n24739_), .ZN(new_n24740_));
  OAI21_X1   g21652(.A1(new_n24740_), .A2(new_n24738_), .B(new_n6845_), .ZN(new_n24741_));
  NOR2_X1    g21653(.A1(new_n24737_), .A2(new_n24741_), .ZN(new_n24742_));
  OAI22_X1   g21654(.A1(new_n24733_), .A2(new_n24729_), .B1(pi0211), .B2(new_n24742_), .ZN(po0368));
  AOI21_X1   g21655(.A1(new_n24509_), .A2(new_n14396_), .B(new_n24728_), .ZN(new_n24744_));
  NOR3_X1    g21656(.A1(new_n24727_), .A2(pi0607), .A3(new_n14396_), .ZN(new_n24745_));
  NOR3_X1    g21657(.A1(new_n3231_), .A2(new_n24509_), .A3(pi0638), .ZN(new_n24746_));
  NAND2_X1   g21658(.A1(new_n6845_), .A2(new_n24498_), .ZN(new_n24747_));
  NOR4_X1    g21659(.A1(new_n24744_), .A2(new_n24745_), .A3(new_n24746_), .A4(new_n24747_), .ZN(new_n24748_));
  OAI21_X1   g21660(.A1(new_n24735_), .A2(new_n24734_), .B(pi0607), .ZN(new_n24749_));
  AOI21_X1   g21661(.A1(new_n24739_), .A2(new_n24512_), .B(po1038), .ZN(new_n24750_));
  OAI21_X1   g21662(.A1(new_n24749_), .A2(new_n24498_), .B(new_n24750_), .ZN(new_n24751_));
  MUX2_X1    g21663(.I0(new_n24751_), .I1(new_n24748_), .S(new_n8076_), .Z(po0369));
  INV_X1     g21664(.I(pi0213), .ZN(new_n24753_));
  NAND2_X1   g21665(.A1(new_n15796_), .A2(new_n3231_), .ZN(new_n24754_));
  INV_X1     g21666(.I(new_n24754_), .ZN(new_n24755_));
  NOR4_X1    g21667(.A1(new_n24755_), .A2(pi0622), .A3(new_n24557_), .A4(new_n24727_), .ZN(new_n24756_));
  AOI21_X1   g21668(.A1(new_n15823_), .A2(new_n24557_), .B(new_n3232_), .ZN(new_n24757_));
  NOR4_X1    g21669(.A1(new_n24756_), .A2(pi0622), .A3(po1038), .A4(new_n24757_), .ZN(new_n24758_));
  OAI21_X1   g21670(.A1(new_n24735_), .A2(new_n24734_), .B(pi0622), .ZN(new_n24759_));
  NOR2_X1    g21671(.A1(new_n24556_), .A2(pi0639), .ZN(new_n24760_));
  AOI21_X1   g21672(.A1(new_n24739_), .A2(new_n24760_), .B(po1038), .ZN(new_n24761_));
  OAI21_X1   g21673(.A1(new_n24759_), .A2(new_n24557_), .B(new_n24761_), .ZN(new_n24762_));
  MUX2_X1    g21674(.I0(new_n24762_), .I1(new_n24758_), .S(new_n24753_), .Z(po0370));
  AOI21_X1   g21675(.A1(new_n24325_), .A2(new_n14396_), .B(new_n24728_), .ZN(new_n24764_));
  NOR3_X1    g21676(.A1(new_n24727_), .A2(pi0623), .A3(new_n14396_), .ZN(new_n24765_));
  NOR3_X1    g21677(.A1(new_n3231_), .A2(new_n24325_), .A3(pi0710), .ZN(new_n24766_));
  NAND2_X1   g21678(.A1(new_n6845_), .A2(new_n24174_), .ZN(new_n24767_));
  NOR4_X1    g21679(.A1(new_n24764_), .A2(new_n24765_), .A3(new_n24766_), .A4(new_n24767_), .ZN(new_n24768_));
  OAI21_X1   g21680(.A1(new_n24735_), .A2(new_n24734_), .B(pi0623), .ZN(new_n24769_));
  AOI21_X1   g21681(.A1(new_n24739_), .A2(new_n24467_), .B(po1038), .ZN(new_n24770_));
  OAI21_X1   g21682(.A1(new_n24769_), .A2(new_n24174_), .B(new_n24770_), .ZN(new_n24771_));
  MUX2_X1    g21683(.I0(new_n24771_), .I1(new_n24768_), .S(new_n8078_), .Z(po0371));
  NOR2_X1    g21684(.A1(new_n12731_), .A2(new_n15305_), .ZN(new_n24773_));
  NOR2_X1    g21685(.A1(new_n24773_), .A2(pi0947), .ZN(new_n24774_));
  AOI21_X1   g21686(.A1(new_n12384_), .A2(pi0947), .B(new_n24774_), .ZN(new_n24775_));
  NOR4_X1    g21687(.A1(new_n13368_), .A2(pi0038), .A3(pi0215), .A4(new_n24775_), .ZN(new_n24776_));
  NAND2_X1   g21688(.A1(new_n15579_), .A2(new_n5473_), .ZN(new_n24777_));
  INV_X1     g21689(.I(new_n24773_), .ZN(new_n24778_));
  NOR2_X1    g21690(.A1(new_n12242_), .A2(new_n5097_), .ZN(new_n24779_));
  INV_X1     g21691(.I(new_n24779_), .ZN(new_n24780_));
  NOR2_X1    g21692(.A1(new_n24780_), .A2(new_n12128_), .ZN(new_n24781_));
  NOR2_X1    g21693(.A1(new_n24781_), .A2(pi0642), .ZN(new_n24782_));
  NOR2_X1    g21694(.A1(new_n24782_), .A2(new_n5100_), .ZN(new_n24783_));
  NAND2_X1   g21695(.A1(new_n12911_), .A2(new_n24783_), .ZN(new_n24784_));
  INV_X1     g21696(.I(new_n24784_), .ZN(new_n24785_));
  MUX2_X1    g21697(.I0(new_n24785_), .I1(new_n24778_), .S(new_n5473_), .Z(new_n24786_));
  AOI21_X1   g21698(.A1(new_n24777_), .A2(new_n24786_), .B(new_n2587_), .ZN(new_n24787_));
  NOR2_X1    g21699(.A1(new_n24775_), .A2(new_n2614_), .ZN(new_n24788_));
  AOI21_X1   g21700(.A1(new_n24788_), .A2(new_n12132_), .B(pi0223), .ZN(new_n24789_));
  NOR2_X1    g21701(.A1(new_n12198_), .A2(pi0642), .ZN(new_n24790_));
  INV_X1     g21702(.I(new_n24790_), .ZN(new_n24791_));
  NOR2_X1    g21703(.A1(new_n12445_), .A2(new_n12400_), .ZN(new_n24792_));
  NOR2_X1    g21704(.A1(new_n24792_), .A2(new_n12168_), .ZN(new_n24793_));
  NOR2_X1    g21705(.A1(new_n12133_), .A2(new_n5104_), .ZN(new_n24794_));
  INV_X1     g21706(.I(new_n24794_), .ZN(new_n24795_));
  OAI21_X1   g21707(.A1(pi0642), .A2(new_n24795_), .B(new_n5217_), .ZN(new_n24796_));
  NAND2_X1   g21708(.A1(new_n5217_), .A2(new_n12384_), .ZN(new_n24797_));
  OAI22_X1   g21709(.A1(new_n24793_), .A2(new_n24796_), .B1(new_n12231_), .B2(new_n24797_), .ZN(new_n24798_));
  OAI21_X1   g21710(.A1(new_n24791_), .A2(new_n24798_), .B(new_n5141_), .ZN(new_n24799_));
  OAI21_X1   g21711(.A1(new_n24799_), .A2(new_n5473_), .B(new_n3155_), .ZN(new_n24800_));
  AOI21_X1   g21712(.A1(new_n15654_), .A2(new_n24774_), .B(new_n24800_), .ZN(new_n24801_));
  NAND2_X1   g21713(.A1(new_n24784_), .A2(new_n5141_), .ZN(new_n24802_));
  MUX2_X1    g21714(.I0(new_n12473_), .I1(new_n12372_), .S(new_n5217_), .Z(new_n24803_));
  NAND3_X1   g21715(.A1(new_n24803_), .A2(new_n12384_), .A3(new_n5141_), .ZN(new_n24804_));
  AOI21_X1   g21716(.A1(new_n24802_), .A2(new_n24804_), .B(new_n5473_), .ZN(new_n24805_));
  NOR2_X1    g21717(.A1(new_n15390_), .A2(new_n24805_), .ZN(new_n24806_));
  OAI21_X1   g21718(.A1(new_n24778_), .A2(pi0947), .B(pi0223), .ZN(new_n24807_));
  OAI22_X1   g21719(.A1(new_n24801_), .A2(new_n24789_), .B1(new_n24806_), .B2(new_n24807_), .ZN(new_n24808_));
  AOI21_X1   g21720(.A1(new_n24808_), .A2(new_n2587_), .B(new_n24787_), .ZN(new_n24809_));
  NOR2_X1    g21721(.A1(new_n12372_), .A2(new_n6460_), .ZN(new_n24810_));
  OAI21_X1   g21722(.A1(new_n24810_), .A2(new_n24778_), .B(new_n5473_), .ZN(new_n24811_));
  AOI21_X1   g21723(.A1(pi0947), .A2(new_n12464_), .B(new_n12362_), .ZN(new_n24812_));
  NAND2_X1   g21724(.A1(new_n24812_), .A2(new_n6460_), .ZN(new_n24813_));
  INV_X1     g21725(.I(new_n24813_), .ZN(new_n24814_));
  NOR3_X1    g21726(.A1(new_n12461_), .A2(new_n12384_), .A3(new_n12713_), .ZN(new_n24815_));
  NOR2_X1    g21727(.A1(new_n12712_), .A2(new_n12384_), .ZN(new_n24816_));
  NOR4_X1    g21728(.A1(new_n12732_), .A2(pi0947), .A3(new_n24815_), .A4(new_n24816_), .ZN(new_n24817_));
  NOR2_X1    g21729(.A1(new_n24814_), .A2(new_n24817_), .ZN(new_n24818_));
  AOI21_X1   g21730(.A1(new_n24818_), .A2(new_n24811_), .B(new_n2604_), .ZN(new_n24819_));
  NAND3_X1   g21731(.A1(new_n6460_), .A2(new_n5473_), .A3(new_n24773_), .ZN(new_n24822_));
  OAI21_X1   g21732(.A1(new_n12453_), .A2(new_n24822_), .B(new_n3155_), .ZN(new_n24823_));
  NAND2_X1   g21733(.A1(new_n12196_), .A2(new_n24773_), .ZN(new_n24824_));
  AOI21_X1   g21734(.A1(new_n12157_), .A2(new_n5217_), .B(new_n12197_), .ZN(new_n24825_));
  NOR3_X1    g21735(.A1(new_n24825_), .A2(new_n12384_), .A3(new_n12461_), .ZN(new_n24826_));
  NOR3_X1    g21736(.A1(new_n12158_), .A2(new_n12384_), .A3(new_n12129_), .ZN(new_n24827_));
  NOR2_X1    g21737(.A1(new_n24826_), .A2(new_n24827_), .ZN(new_n24828_));
  MUX2_X1    g21738(.I0(new_n24828_), .I1(new_n24824_), .S(new_n5473_), .Z(new_n24829_));
  AND2_X2    g21739(.A1(new_n24829_), .A2(new_n6460_), .Z(new_n24830_));
  NAND3_X1   g21740(.A1(new_n24775_), .A2(new_n2614_), .A3(new_n12132_), .ZN(new_n24831_));
  AOI22_X1   g21741(.A1(new_n24830_), .A2(new_n24823_), .B1(new_n2604_), .B2(new_n24831_), .ZN(new_n24832_));
  OAI21_X1   g21742(.A1(new_n24832_), .A2(new_n24819_), .B(new_n2587_), .ZN(new_n24833_));
  AOI21_X1   g21743(.A1(new_n24775_), .A2(new_n12770_), .B(new_n2587_), .ZN(new_n24834_));
  OAI21_X1   g21744(.A1(new_n24829_), .A2(new_n3284_), .B(new_n24834_), .ZN(new_n24835_));
  NAND2_X1   g21745(.A1(new_n24833_), .A2(new_n24835_), .ZN(new_n24836_));
  AOI21_X1   g21746(.A1(new_n24836_), .A2(new_n2566_), .B(new_n3154_), .ZN(new_n24837_));
  OAI21_X1   g21747(.A1(new_n24809_), .A2(new_n2566_), .B(new_n24837_), .ZN(new_n24838_));
  XOR2_X1    g21748(.A1(new_n24775_), .A2(pi0215), .Z(new_n24839_));
  NAND2_X1   g21749(.A1(new_n12646_), .A2(new_n24839_), .ZN(new_n24840_));
  AOI21_X1   g21750(.A1(new_n24840_), .A2(new_n24775_), .B(new_n6594_), .ZN(new_n24841_));
  NOR2_X1    g21751(.A1(new_n24840_), .A2(new_n24775_), .ZN(new_n24842_));
  NOR3_X1    g21752(.A1(new_n12652_), .A2(new_n24682_), .A3(new_n24775_), .ZN(new_n24843_));
  NOR2_X1    g21753(.A1(new_n24842_), .A2(new_n24843_), .ZN(new_n24844_));
  AOI21_X1   g21754(.A1(new_n24844_), .A2(new_n24841_), .B(pi0038), .ZN(new_n24845_));
  AOI21_X1   g21755(.A1(new_n24838_), .A2(new_n24845_), .B(new_n24776_), .ZN(new_n24846_));
  MUX2_X1    g21756(.I0(new_n24846_), .I1(pi0215), .S(new_n7833_), .Z(po0372));
  INV_X1     g21757(.I(pi0662), .ZN(new_n24848_));
  NOR2_X1    g21758(.A1(new_n15372_), .A2(new_n24848_), .ZN(new_n24849_));
  NOR2_X1    g21759(.A1(new_n12443_), .A2(new_n5473_), .ZN(new_n24850_));
  NOR2_X1    g21760(.A1(new_n24849_), .A2(new_n24850_), .ZN(new_n24851_));
  INV_X1     g21761(.I(new_n24851_), .ZN(new_n24852_));
  NOR3_X1    g21762(.A1(new_n13368_), .A2(new_n3267_), .A3(new_n24852_), .ZN(new_n24853_));
  INV_X1     g21763(.I(new_n15390_), .ZN(new_n24854_));
  NOR3_X1    g21764(.A1(new_n12249_), .A2(new_n5427_), .A3(new_n12242_), .ZN(new_n24855_));
  AOI21_X1   g21765(.A1(new_n5106_), .A2(new_n12242_), .B(new_n12464_), .ZN(new_n24856_));
  OAI22_X1   g21766(.A1(new_n24856_), .A2(new_n24855_), .B1(new_n12443_), .B2(pi0616), .ZN(new_n24857_));
  NAND2_X1   g21767(.A1(new_n24857_), .A2(new_n5100_), .ZN(new_n24858_));
  AOI21_X1   g21768(.A1(new_n12262_), .A2(new_n5100_), .B(pi0614), .ZN(new_n24859_));
  AND2_X2    g21769(.A1(new_n24858_), .A2(new_n24859_), .Z(new_n24860_));
  INV_X1     g21770(.I(new_n24860_), .ZN(new_n24861_));
  NOR2_X1    g21771(.A1(new_n12360_), .A2(new_n12166_), .ZN(new_n24862_));
  NAND2_X1   g21772(.A1(new_n12132_), .A2(pi0616), .ZN(new_n24863_));
  NAND4_X1   g21773(.A1(new_n12725_), .A2(new_n12443_), .A3(new_n5217_), .A4(new_n24863_), .ZN(new_n24864_));
  NOR2_X1    g21774(.A1(new_n24862_), .A2(new_n24864_), .ZN(new_n24865_));
  NOR3_X1    g21775(.A1(new_n24861_), .A2(new_n5141_), .A3(new_n24865_), .ZN(new_n24866_));
  AOI21_X1   g21776(.A1(new_n6460_), .A2(new_n24865_), .B(new_n24860_), .ZN(new_n24867_));
  OAI21_X1   g21777(.A1(new_n24866_), .A2(new_n24867_), .B(new_n5473_), .ZN(new_n24868_));
  INV_X1     g21778(.I(new_n24849_), .ZN(new_n24869_));
  NAND3_X1   g21779(.A1(new_n24869_), .A2(new_n2562_), .A3(pi0223), .ZN(new_n24870_));
  AOI21_X1   g21780(.A1(new_n24854_), .A2(new_n24868_), .B(new_n24870_), .ZN(new_n24871_));
  NOR2_X1    g21781(.A1(new_n24848_), .A2(new_n15305_), .ZN(new_n24872_));
  NAND3_X1   g21782(.A1(new_n12879_), .A2(new_n5473_), .A3(new_n24872_), .ZN(new_n24873_));
  NAND2_X1   g21783(.A1(new_n12863_), .A2(pi0947), .ZN(new_n24874_));
  AOI21_X1   g21784(.A1(new_n24873_), .A2(new_n24874_), .B(new_n6460_), .ZN(new_n24875_));
  NOR2_X1    g21785(.A1(new_n12776_), .A2(pi0947), .ZN(new_n24876_));
  AOI21_X1   g21786(.A1(new_n12809_), .A2(new_n12443_), .B(new_n5473_), .ZN(new_n24877_));
  OR3_X2     g21787(.A1(new_n24877_), .A2(new_n5141_), .A3(new_n24849_), .Z(new_n24878_));
  OAI21_X1   g21788(.A1(new_n24878_), .A2(new_n24876_), .B(new_n3155_), .ZN(new_n24879_));
  NOR2_X1    g21789(.A1(new_n24852_), .A2(new_n2614_), .ZN(new_n24880_));
  AOI21_X1   g21790(.A1(new_n24880_), .A2(new_n12132_), .B(pi0223), .ZN(new_n24881_));
  NAND2_X1   g21791(.A1(new_n24879_), .A2(new_n24881_), .ZN(new_n24882_));
  NOR3_X1    g21792(.A1(new_n24871_), .A2(new_n24875_), .A3(new_n24882_), .ZN(new_n24883_));
  NAND2_X1   g21793(.A1(new_n12412_), .A2(new_n24849_), .ZN(new_n24884_));
  AOI21_X1   g21794(.A1(new_n12757_), .A2(pi0947), .B(new_n6460_), .ZN(new_n24885_));
  INV_X1     g21795(.I(new_n24825_), .ZN(new_n24886_));
  NAND2_X1   g21796(.A1(new_n24886_), .A2(new_n24850_), .ZN(new_n24887_));
  OAI21_X1   g21797(.A1(new_n12326_), .A2(new_n24869_), .B(new_n24887_), .ZN(new_n24888_));
  OAI21_X1   g21798(.A1(new_n24888_), .A2(new_n5141_), .B(new_n3155_), .ZN(new_n24889_));
  AOI21_X1   g21799(.A1(new_n24884_), .A2(new_n24885_), .B(new_n24889_), .ZN(new_n24890_));
  NAND3_X1   g21800(.A1(new_n24852_), .A2(new_n2614_), .A3(new_n12132_), .ZN(new_n24891_));
  NAND2_X1   g21801(.A1(new_n24891_), .A2(new_n2604_), .ZN(new_n24892_));
  NAND2_X1   g21802(.A1(new_n2562_), .A2(new_n2587_), .ZN(new_n24893_));
  INV_X1     g21803(.I(new_n24810_), .ZN(new_n24894_));
  NAND2_X1   g21804(.A1(new_n24894_), .A2(new_n24872_), .ZN(new_n24895_));
  NAND4_X1   g21805(.A1(new_n12716_), .A2(new_n5473_), .A3(new_n12753_), .A4(new_n12755_), .ZN(new_n24896_));
  NAND4_X1   g21806(.A1(new_n24813_), .A2(new_n24895_), .A3(new_n5473_), .A4(new_n24896_), .ZN(new_n24897_));
  AOI21_X1   g21807(.A1(new_n24897_), .A2(pi0223), .B(new_n24893_), .ZN(new_n24898_));
  OAI21_X1   g21808(.A1(new_n24890_), .A2(new_n24892_), .B(new_n24898_), .ZN(new_n24899_));
  OAI21_X1   g21809(.A1(new_n24883_), .A2(new_n24899_), .B(pi0039), .ZN(new_n24900_));
  NAND2_X1   g21810(.A1(new_n15436_), .A2(new_n5473_), .ZN(new_n24901_));
  AOI22_X1   g21811(.A1(new_n24888_), .A2(new_n4135_), .B1(new_n12770_), .B2(new_n24852_), .ZN(new_n24902_));
  NOR4_X1    g21812(.A1(new_n24902_), .A2(new_n2562_), .A3(new_n24849_), .A4(new_n24877_), .ZN(new_n24903_));
  NOR3_X1    g21813(.A1(new_n24896_), .A2(new_n5473_), .A3(new_n12464_), .ZN(new_n24905_));
  OAI21_X1   g21814(.A1(new_n24905_), .A2(pi0216), .B(pi0215), .ZN(new_n24906_));
  OAI21_X1   g21815(.A1(new_n12584_), .A2(pi0216), .B(new_n24852_), .ZN(new_n24907_));
  NAND3_X1   g21816(.A1(new_n12646_), .A2(pi0216), .A3(new_n24851_), .ZN(new_n24908_));
  NAND4_X1   g21817(.A1(new_n12590_), .A2(new_n2562_), .A3(new_n2587_), .A4(new_n24851_), .ZN(new_n24909_));
  NAND4_X1   g21818(.A1(new_n24908_), .A2(new_n24909_), .A3(new_n24907_), .A4(new_n6593_), .ZN(new_n24910_));
  NOR4_X1    g21819(.A1(new_n24849_), .A2(pi0216), .A3(new_n5473_), .A4(new_n24682_), .ZN(new_n24911_));
  NAND2_X1   g21820(.A1(new_n24861_), .A2(new_n24911_), .ZN(new_n24912_));
  AOI21_X1   g21821(.A1(new_n24910_), .A2(new_n3172_), .B(new_n24912_), .ZN(new_n24913_));
  NAND3_X1   g21822(.A1(new_n24913_), .A2(new_n24777_), .A3(new_n24906_), .ZN(new_n24914_));
  AOI21_X1   g21823(.A1(new_n24901_), .A2(new_n24903_), .B(new_n24914_), .ZN(new_n24915_));
  AOI21_X1   g21824(.A1(new_n24915_), .A2(new_n24900_), .B(new_n24853_), .ZN(new_n24916_));
  MUX2_X1    g21825(.I0(new_n24916_), .I1(pi0216), .S(new_n7833_), .Z(po0373));
  NOR2_X1    g21826(.A1(new_n24619_), .A2(pi0695), .ZN(new_n24918_));
  INV_X1     g21827(.I(pi0612), .ZN(new_n24919_));
  INV_X1     g21828(.I(pi0695), .ZN(new_n24920_));
  NAND3_X1   g21829(.A1(new_n24567_), .A2(new_n9637_), .A3(new_n24920_), .ZN(new_n24921_));
  NAND2_X1   g21830(.A1(new_n24605_), .A2(pi0695), .ZN(new_n24922_));
  NAND4_X1   g21831(.A1(new_n24921_), .A2(new_n9637_), .A3(new_n24919_), .A4(new_n24922_), .ZN(new_n24923_));
  NAND2_X1   g21832(.A1(new_n24636_), .A2(new_n24637_), .ZN(new_n24924_));
  MUX2_X1    g21833(.I0(new_n24642_), .I1(new_n24924_), .S(new_n24920_), .Z(new_n24925_));
  NOR2_X1    g21834(.A1(new_n24925_), .A2(pi0217), .ZN(new_n24926_));
  AND4_X2    g21835(.A1(new_n9637_), .A2(new_n24555_), .A3(pi0695), .A4(new_n24571_), .Z(new_n24927_));
  NOR2_X1    g21836(.A1(new_n24926_), .A2(new_n24927_), .ZN(new_n24928_));
  OAI22_X1   g21837(.A1(new_n24928_), .A2(pi0612), .B1(new_n24918_), .B2(new_n24923_), .ZN(po0374));
  NOR2_X1    g21838(.A1(new_n24110_), .A2(new_n24087_), .ZN(new_n24930_));
  NOR2_X1    g21839(.A1(new_n24114_), .A2(new_n24087_), .ZN(new_n24931_));
  NAND2_X1   g21840(.A1(new_n24931_), .A2(pi0218), .ZN(new_n24932_));
  OAI21_X1   g21841(.A1(new_n24930_), .A2(pi0218), .B(new_n24932_), .ZN(po0375));
  AOI21_X1   g21842(.A1(new_n23615_), .A2(new_n14396_), .B(new_n24728_), .ZN(new_n24934_));
  NAND3_X1   g21843(.A1(new_n24728_), .A2(new_n23615_), .A3(new_n12965_), .ZN(new_n24935_));
  NOR3_X1    g21844(.A1(new_n3231_), .A2(new_n23615_), .A3(pi0637), .ZN(new_n24936_));
  NOR4_X1    g21845(.A1(new_n24936_), .A2(new_n8247_), .A3(pi0637), .A4(po1038), .ZN(new_n24937_));
  NAND2_X1   g21846(.A1(new_n24935_), .A2(new_n24937_), .ZN(new_n24938_));
  OAI21_X1   g21847(.A1(new_n24735_), .A2(new_n24734_), .B(pi0617), .ZN(new_n24939_));
  NOR2_X1    g21848(.A1(new_n24939_), .A2(new_n23598_), .ZN(new_n24940_));
  NAND2_X1   g21849(.A1(new_n23598_), .A2(pi0617), .ZN(new_n24941_));
  OAI21_X1   g21850(.A1(new_n24740_), .A2(new_n24941_), .B(new_n6845_), .ZN(new_n24942_));
  NOR2_X1    g21851(.A1(new_n24940_), .A2(new_n24942_), .ZN(new_n24943_));
  OAI22_X1   g21852(.A1(new_n24938_), .A2(new_n24934_), .B1(pi0219), .B2(new_n24943_), .ZN(po0376));
  INV_X1     g21853(.I(pi0220), .ZN(new_n24945_));
  NAND3_X1   g21854(.A1(new_n24068_), .A2(new_n24945_), .A3(new_n24122_), .ZN(new_n24946_));
  NOR2_X1    g21855(.A1(new_n24076_), .A2(new_n24124_), .ZN(new_n24947_));
  NAND2_X1   g21856(.A1(new_n24947_), .A2(pi0220), .ZN(new_n24948_));
  NAND2_X1   g21857(.A1(new_n24946_), .A2(new_n24948_), .ZN(po0377));
  INV_X1     g21858(.I(pi0661), .ZN(new_n24950_));
  NOR2_X1    g21859(.A1(new_n15372_), .A2(new_n24950_), .ZN(new_n24951_));
  NOR2_X1    g21860(.A1(new_n12166_), .A2(new_n5473_), .ZN(new_n24952_));
  NOR2_X1    g21861(.A1(new_n24951_), .A2(new_n24952_), .ZN(new_n24953_));
  INV_X1     g21862(.I(new_n24953_), .ZN(new_n24954_));
  NOR4_X1    g21863(.A1(new_n13368_), .A2(pi0038), .A3(pi0221), .A4(new_n24954_), .ZN(new_n24955_));
  NOR2_X1    g21864(.A1(new_n12156_), .A2(new_n5109_), .ZN(new_n24956_));
  AOI21_X1   g21865(.A1(new_n12452_), .A2(new_n12443_), .B(new_n12721_), .ZN(new_n24957_));
  AOI21_X1   g21866(.A1(new_n24957_), .A2(new_n5109_), .B(new_n24956_), .ZN(new_n24958_));
  NOR3_X1    g21867(.A1(new_n12461_), .A2(pi0616), .A3(pi0947), .ZN(new_n24959_));
  OAI21_X1   g21868(.A1(new_n24790_), .A2(new_n24826_), .B(new_n24959_), .ZN(new_n24960_));
  AOI21_X1   g21869(.A1(new_n24958_), .A2(new_n12718_), .B(new_n24960_), .ZN(new_n24961_));
  INV_X1     g21870(.I(new_n24961_), .ZN(new_n24962_));
  NOR2_X1    g21871(.A1(new_n24950_), .A2(new_n15305_), .ZN(new_n24963_));
  OAI21_X1   g21872(.A1(new_n15436_), .A2(new_n24963_), .B(new_n5473_), .ZN(new_n24964_));
  AOI22_X1   g21873(.A1(new_n24886_), .A2(new_n24952_), .B1(new_n12196_), .B2(new_n24951_), .ZN(new_n24965_));
  NAND3_X1   g21874(.A1(new_n12132_), .A2(pi0216), .A3(new_n2550_), .ZN(new_n24966_));
  OAI21_X1   g21875(.A1(new_n24965_), .A2(new_n24966_), .B(new_n2530_), .ZN(new_n24967_));
  AOI21_X1   g21876(.A1(new_n24964_), .A2(new_n24962_), .B(new_n24967_), .ZN(new_n24968_));
  NOR2_X1    g21877(.A1(new_n12733_), .A2(new_n5473_), .ZN(new_n24969_));
  NOR2_X1    g21878(.A1(new_n24969_), .A2(new_n24951_), .ZN(new_n24970_));
  OAI21_X1   g21879(.A1(new_n24812_), .A2(new_n24970_), .B(new_n2550_), .ZN(new_n24971_));
  NAND2_X1   g21880(.A1(new_n24971_), .A2(pi0215), .ZN(new_n24972_));
  NOR2_X1    g21881(.A1(new_n12360_), .A2(pi0614), .ZN(new_n24973_));
  NOR2_X1    g21882(.A1(new_n24973_), .A2(new_n12249_), .ZN(new_n24974_));
  NOR2_X1    g21883(.A1(new_n24974_), .A2(new_n5100_), .ZN(new_n24975_));
  INV_X1     g21884(.I(new_n24975_), .ZN(new_n24976_));
  NOR2_X1    g21885(.A1(new_n24781_), .A2(pi0616), .ZN(new_n24977_));
  AOI21_X1   g21886(.A1(new_n24976_), .A2(new_n24977_), .B(new_n5473_), .ZN(new_n24978_));
  NOR4_X1    g21887(.A1(new_n24978_), .A2(new_n2550_), .A3(pi0299), .A4(new_n24951_), .ZN(new_n24979_));
  NAND3_X1   g21888(.A1(new_n24777_), .A2(new_n24972_), .A3(new_n24979_), .ZN(new_n24980_));
  NAND3_X1   g21889(.A1(new_n24954_), .A2(new_n2614_), .A3(new_n12132_), .ZN(new_n24981_));
  NAND2_X1   g21890(.A1(new_n12872_), .A2(new_n12754_), .ZN(new_n24982_));
  NAND4_X1   g21891(.A1(new_n12871_), .A2(pi0616), .A3(new_n12129_), .A4(new_n24982_), .ZN(new_n24983_));
  NOR4_X1    g21892(.A1(new_n12759_), .A2(new_n5473_), .A3(new_n5141_), .A4(new_n24983_), .ZN(new_n24984_));
  NOR2_X1    g21893(.A1(new_n24951_), .A2(new_n5141_), .ZN(new_n24985_));
  OAI21_X1   g21894(.A1(new_n24961_), .A2(new_n24876_), .B(new_n24985_), .ZN(new_n24986_));
  OAI21_X1   g21895(.A1(new_n24984_), .A2(new_n24986_), .B(new_n2614_), .ZN(new_n24987_));
  AOI22_X1   g21896(.A1(new_n24987_), .A2(new_n12505_), .B1(new_n2604_), .B2(new_n24981_), .ZN(new_n24988_));
  NAND2_X1   g21897(.A1(new_n12722_), .A2(new_n12727_), .ZN(new_n24989_));
  INV_X1     g21898(.I(new_n12786_), .ZN(new_n24990_));
  MUX2_X1    g21899(.I0(new_n24990_), .I1(new_n24989_), .S(new_n5473_), .Z(new_n24991_));
  AOI21_X1   g21900(.A1(new_n12784_), .A2(new_n5473_), .B(new_n24978_), .ZN(new_n24992_));
  OAI21_X1   g21901(.A1(new_n15372_), .A2(new_n24950_), .B(pi0223), .ZN(new_n24993_));
  NOR4_X1    g21902(.A1(new_n24991_), .A2(new_n5141_), .A3(new_n24992_), .A4(new_n24993_), .ZN(new_n24994_));
  NOR2_X1    g21903(.A1(new_n24988_), .A2(new_n24994_), .ZN(new_n24995_));
  AOI21_X1   g21904(.A1(new_n24894_), .A2(new_n24951_), .B(new_n24969_), .ZN(new_n24996_));
  OAI21_X1   g21905(.A1(new_n24814_), .A2(new_n24996_), .B(pi0223), .ZN(new_n24997_));
  NAND2_X1   g21906(.A1(new_n24997_), .A2(new_n2550_), .ZN(new_n24998_));
  NOR4_X1    g21907(.A1(new_n5141_), .A2(new_n24950_), .A3(new_n15305_), .A4(pi0947), .ZN(new_n25000_));
  NAND2_X1   g21908(.A1(new_n12412_), .A2(new_n25000_), .ZN(new_n25001_));
  NAND2_X1   g21909(.A1(new_n24965_), .A2(new_n6460_), .ZN(new_n25002_));
  NOR2_X1    g21910(.A1(new_n2614_), .A2(new_n2604_), .ZN(new_n25003_));
  NAND4_X1   g21911(.A1(new_n24998_), .A2(new_n25001_), .A3(new_n25002_), .A4(new_n25003_), .ZN(new_n25004_));
  NAND3_X1   g21912(.A1(new_n25004_), .A2(new_n2550_), .A3(new_n2587_), .ZN(new_n25005_));
  OAI22_X1   g21913(.A1(new_n24995_), .A2(new_n25005_), .B1(new_n24968_), .B2(new_n24980_), .ZN(new_n25006_));
  OAI21_X1   g21914(.A1(new_n12584_), .A2(pi0221), .B(new_n24954_), .ZN(new_n25007_));
  NAND3_X1   g21915(.A1(new_n12646_), .A2(pi0221), .A3(new_n24953_), .ZN(new_n25008_));
  NAND4_X1   g21916(.A1(new_n12590_), .A2(new_n2550_), .A3(new_n2587_), .A4(new_n24953_), .ZN(new_n25009_));
  NAND4_X1   g21917(.A1(new_n25008_), .A2(new_n25009_), .A3(new_n25007_), .A4(new_n6593_), .ZN(new_n25010_));
  AOI21_X1   g21918(.A1(new_n25010_), .A2(new_n3172_), .B(pi0039), .ZN(new_n25011_));
  AOI21_X1   g21919(.A1(new_n25006_), .A2(new_n25011_), .B(new_n24955_), .ZN(new_n25012_));
  MUX2_X1    g21920(.I0(new_n25012_), .I1(pi0221), .S(new_n7833_), .Z(po0378));
  AOI21_X1   g21921(.A1(new_n15392_), .A2(pi0223), .B(new_n10309_), .ZN(new_n25014_));
  OAI21_X1   g21922(.A1(new_n15654_), .A2(new_n2604_), .B(new_n25014_), .ZN(new_n25015_));
  NOR2_X1    g21923(.A1(new_n13384_), .A2(pi0038), .ZN(new_n25016_));
  OAI21_X1   g21924(.A1(new_n25015_), .A2(new_n12885_), .B(new_n25016_), .ZN(new_n25017_));
  NAND2_X1   g21925(.A1(new_n25017_), .A2(new_n13972_), .ZN(new_n25018_));
  INV_X1     g21926(.I(new_n25018_), .ZN(new_n25019_));
  NOR2_X1    g21927(.A1(new_n25019_), .A2(new_n2588_), .ZN(new_n25020_));
  NOR2_X1    g21928(.A1(new_n25020_), .A2(new_n12054_), .ZN(new_n25021_));
  INV_X1     g21929(.I(new_n25020_), .ZN(new_n25022_));
  NOR2_X1    g21930(.A1(new_n25022_), .A2(new_n14624_), .ZN(new_n25023_));
  NAND2_X1   g21931(.A1(new_n3232_), .A2(pi0222), .ZN(new_n25024_));
  NAND2_X1   g21932(.A1(new_n12735_), .A2(new_n12723_), .ZN(new_n25025_));
  AOI21_X1   g21933(.A1(pi0616), .A2(new_n12287_), .B(new_n25025_), .ZN(new_n25026_));
  NOR2_X1    g21934(.A1(new_n11875_), .A2(new_n12166_), .ZN(new_n25027_));
  NOR2_X1    g21935(.A1(new_n5096_), .A2(new_n12127_), .ZN(new_n25028_));
  NAND2_X1   g21936(.A1(new_n25026_), .A2(new_n25028_), .ZN(new_n25029_));
  OAI21_X1   g21937(.A1(new_n12127_), .A2(new_n25026_), .B(new_n25029_), .ZN(new_n25030_));
  OR2_X2     g21938(.A1(new_n25030_), .A2(new_n6460_), .Z(new_n25031_));
  NOR2_X1    g21939(.A1(new_n12362_), .A2(new_n5096_), .ZN(new_n25032_));
  NOR2_X1    g21940(.A1(new_n12307_), .A2(new_n12166_), .ZN(new_n25033_));
  NOR2_X1    g21941(.A1(new_n24779_), .A2(new_n25033_), .ZN(new_n25034_));
  NOR3_X1    g21942(.A1(new_n25032_), .A2(new_n12127_), .A3(new_n25034_), .ZN(new_n25035_));
  OAI21_X1   g21943(.A1(new_n12166_), .A2(new_n12307_), .B(new_n12362_), .ZN(new_n25036_));
  AOI21_X1   g21944(.A1(new_n12128_), .A2(new_n25036_), .B(new_n25035_), .ZN(new_n25037_));
  NOR3_X1    g21945(.A1(new_n25037_), .A2(pi0222), .A3(new_n6460_), .ZN(new_n25038_));
  NOR2_X1    g21946(.A1(new_n12209_), .A2(new_n12166_), .ZN(new_n25039_));
  INV_X1     g21947(.I(new_n25039_), .ZN(new_n25040_));
  NAND2_X1   g21948(.A1(new_n12243_), .A2(new_n5100_), .ZN(new_n25041_));
  INV_X1     g21949(.I(new_n25041_), .ZN(new_n25042_));
  NOR2_X1    g21950(.A1(new_n25042_), .A2(new_n25040_), .ZN(new_n25043_));
  NAND4_X1   g21951(.A1(new_n25043_), .A2(new_n2588_), .A3(new_n2604_), .A4(new_n12686_), .ZN(new_n25044_));
  AOI21_X1   g21952(.A1(new_n25038_), .A2(new_n25031_), .B(new_n25044_), .ZN(new_n25045_));
  INV_X1     g21953(.I(new_n12489_), .ZN(new_n25046_));
  NAND2_X1   g21954(.A1(new_n24958_), .A2(new_n12166_), .ZN(new_n25047_));
  OAI21_X1   g21955(.A1(new_n12166_), .A2(new_n25046_), .B(new_n25047_), .ZN(new_n25048_));
  INV_X1     g21956(.I(new_n25048_), .ZN(new_n25049_));
  INV_X1     g21957(.I(new_n25027_), .ZN(new_n25050_));
  OAI21_X1   g21958(.A1(new_n12170_), .A2(new_n25050_), .B(new_n12182_), .ZN(new_n25051_));
  MUX2_X1    g21959(.I0(new_n25048_), .I1(new_n25051_), .S(new_n5097_), .Z(new_n25052_));
  OAI21_X1   g21960(.A1(new_n25052_), .A2(new_n25049_), .B(new_n12128_), .ZN(new_n25053_));
  INV_X1     g21961(.I(new_n24957_), .ZN(new_n25054_));
  NOR2_X1    g21962(.A1(new_n12287_), .A2(new_n12166_), .ZN(new_n25055_));
  AOI21_X1   g21963(.A1(new_n25054_), .A2(new_n12166_), .B(new_n25055_), .ZN(new_n25056_));
  NAND2_X1   g21964(.A1(new_n5097_), .A2(new_n12128_), .ZN(new_n25057_));
  NOR2_X1    g21965(.A1(new_n25056_), .A2(new_n25057_), .ZN(new_n25058_));
  AOI21_X1   g21966(.A1(new_n12128_), .A2(new_n25056_), .B(new_n25058_), .ZN(new_n25059_));
  NOR4_X1    g21967(.A1(new_n25053_), .A2(pi0222), .A3(new_n6460_), .A4(new_n25059_), .ZN(new_n25060_));
  MUX2_X1    g21968(.I0(new_n12208_), .I1(new_n12206_), .S(new_n5100_), .Z(new_n25061_));
  NAND2_X1   g21969(.A1(new_n25061_), .A2(pi0616), .ZN(new_n25062_));
  NAND2_X1   g21970(.A1(new_n12157_), .A2(new_n11874_), .ZN(new_n25063_));
  NOR2_X1    g21971(.A1(new_n25063_), .A2(new_n12166_), .ZN(new_n25064_));
  NOR4_X1    g21972(.A1(new_n12426_), .A2(new_n12166_), .A3(new_n5097_), .A4(new_n12127_), .ZN(new_n25065_));
  INV_X1     g21973(.I(new_n25065_), .ZN(new_n25066_));
  OAI21_X1   g21974(.A1(new_n25064_), .A2(new_n12127_), .B(new_n25066_), .ZN(new_n25067_));
  NAND4_X1   g21975(.A1(new_n25062_), .A2(new_n2595_), .A3(new_n5141_), .A4(new_n25067_), .ZN(new_n25068_));
  AND2_X2    g21976(.A1(new_n25068_), .A2(new_n2588_), .Z(new_n25069_));
  NAND2_X1   g21977(.A1(new_n25040_), .A2(new_n2595_), .ZN(new_n25070_));
  OAI21_X1   g21978(.A1(new_n25069_), .A2(new_n25070_), .B(new_n2604_), .ZN(new_n25071_));
  NOR2_X1    g21979(.A1(new_n25060_), .A2(new_n25071_), .ZN(new_n25072_));
  OAI21_X1   g21980(.A1(new_n25072_), .A2(new_n25045_), .B(new_n2587_), .ZN(new_n25073_));
  NOR4_X1    g21981(.A1(new_n25053_), .A2(pi0222), .A3(new_n6445_), .A4(new_n25059_), .ZN(new_n25074_));
  MUX2_X1    g21982(.I0(new_n25067_), .I1(new_n25062_), .S(new_n5094_), .Z(new_n25075_));
  OAI21_X1   g21983(.A1(new_n25075_), .A2(pi0222), .B(new_n3285_), .ZN(new_n25076_));
  AOI21_X1   g21984(.A1(new_n12133_), .A2(pi0222), .B(new_n3285_), .ZN(new_n25077_));
  AOI21_X1   g21985(.A1(new_n25040_), .A2(new_n25077_), .B(pi0215), .ZN(new_n25078_));
  OAI21_X1   g21986(.A1(new_n25074_), .A2(new_n25076_), .B(new_n25078_), .ZN(new_n25079_));
  INV_X1     g21987(.I(new_n25037_), .ZN(new_n25080_));
  NAND4_X1   g21988(.A1(new_n25080_), .A2(new_n2588_), .A3(new_n25030_), .A4(new_n5094_), .ZN(new_n25081_));
  INV_X1     g21989(.I(new_n25043_), .ZN(new_n25082_));
  OAI21_X1   g21990(.A1(new_n25082_), .A2(pi0222), .B(new_n12676_), .ZN(new_n25083_));
  AOI21_X1   g21991(.A1(new_n25081_), .A2(new_n25083_), .B(new_n24682_), .ZN(new_n25084_));
  AOI21_X1   g21992(.A1(new_n25079_), .A2(new_n25084_), .B(new_n3154_), .ZN(new_n25085_));
  NAND2_X1   g21993(.A1(new_n25085_), .A2(new_n25073_), .ZN(new_n25086_));
  AOI21_X1   g21994(.A1(new_n13368_), .A2(pi0222), .B(new_n3172_), .ZN(new_n25087_));
  NOR4_X1    g21995(.A1(new_n25087_), .A2(new_n12166_), .A3(new_n3231_), .A4(new_n13367_), .ZN(new_n25088_));
  AOI21_X1   g21996(.A1(new_n12667_), .A2(new_n12166_), .B(pi0039), .ZN(new_n25089_));
  OAI21_X1   g21997(.A1(pi0222), .A2(new_n12667_), .B(new_n25089_), .ZN(new_n25090_));
  NAND3_X1   g21998(.A1(new_n25090_), .A2(pi0222), .A3(new_n13346_), .ZN(new_n25091_));
  AOI21_X1   g21999(.A1(new_n25091_), .A2(new_n3172_), .B(new_n25088_), .ZN(new_n25092_));
  NAND2_X1   g22000(.A1(new_n25086_), .A2(new_n25092_), .ZN(new_n25093_));
  NAND2_X1   g22001(.A1(new_n25093_), .A2(new_n25024_), .ZN(new_n25094_));
  NOR2_X1    g22002(.A1(new_n25020_), .A2(new_n11924_), .ZN(new_n25095_));
  AOI21_X1   g22003(.A1(new_n25094_), .A2(new_n11924_), .B(new_n25095_), .ZN(new_n25096_));
  NAND2_X1   g22004(.A1(new_n25096_), .A2(new_n11870_), .ZN(new_n25097_));
  NOR3_X1    g22005(.A1(new_n25096_), .A2(pi0609), .A3(new_n25022_), .ZN(new_n25098_));
  AOI21_X1   g22006(.A1(new_n25096_), .A2(new_n11903_), .B(new_n25020_), .ZN(new_n25099_));
  NOR3_X1    g22007(.A1(new_n25098_), .A2(new_n25099_), .A3(pi1155), .ZN(new_n25100_));
  NOR2_X1    g22008(.A1(new_n25100_), .A2(new_n11870_), .ZN(new_n25101_));
  XOR2_X1    g22009(.A1(new_n25101_), .A2(new_n25097_), .Z(new_n25102_));
  NAND3_X1   g22010(.A1(new_n25102_), .A2(new_n11934_), .A3(new_n25020_), .ZN(new_n25103_));
  OAI21_X1   g22011(.A1(new_n25102_), .A2(pi0618), .B(new_n25022_), .ZN(new_n25104_));
  AND3_X2    g22012(.A1(new_n25104_), .A2(new_n25103_), .A3(new_n11950_), .Z(new_n25105_));
  MUX2_X1    g22013(.I0(new_n25105_), .I1(new_n25102_), .S(new_n11969_), .Z(new_n25106_));
  NOR2_X1    g22014(.A1(new_n25106_), .A2(pi0789), .ZN(new_n25107_));
  NAND3_X1   g22015(.A1(new_n25106_), .A2(new_n11967_), .A3(new_n25020_), .ZN(new_n25108_));
  OAI21_X1   g22016(.A1(new_n25106_), .A2(pi0619), .B(new_n25022_), .ZN(new_n25109_));
  NAND3_X1   g22017(.A1(new_n25109_), .A2(new_n25108_), .A3(new_n11869_), .ZN(new_n25110_));
  NAND2_X1   g22018(.A1(new_n25110_), .A2(pi0789), .ZN(new_n25111_));
  XNOR2_X1   g22019(.A1(new_n25111_), .A2(new_n25107_), .ZN(new_n25112_));
  AOI21_X1   g22020(.A1(new_n25112_), .A2(new_n14624_), .B(new_n25023_), .ZN(new_n25113_));
  AOI21_X1   g22021(.A1(new_n25113_), .A2(new_n12054_), .B(new_n25021_), .ZN(new_n25114_));
  NOR2_X1    g22022(.A1(new_n25020_), .A2(new_n12067_), .ZN(new_n25115_));
  NOR2_X1    g22023(.A1(new_n12731_), .A2(pi0661), .ZN(new_n25116_));
  NAND2_X1   g22024(.A1(new_n12453_), .A2(new_n25116_), .ZN(new_n25117_));
  AOI21_X1   g22025(.A1(new_n12453_), .A2(new_n5095_), .B(new_n12921_), .ZN(new_n25118_));
  NOR2_X1    g22026(.A1(new_n25118_), .A2(new_n24950_), .ZN(new_n25119_));
  XOR2_X1    g22027(.A1(new_n25119_), .A2(new_n25117_), .Z(new_n25120_));
  AOI21_X1   g22028(.A1(new_n12412_), .A2(new_n5096_), .B(new_n12231_), .ZN(new_n25121_));
  NOR3_X1    g22029(.A1(new_n12412_), .A2(new_n5097_), .A3(new_n12495_), .ZN(new_n25122_));
  NOR3_X1    g22030(.A1(new_n25122_), .A2(new_n25121_), .A3(new_n12128_), .ZN(new_n25123_));
  NOR2_X1    g22031(.A1(new_n25120_), .A2(new_n25123_), .ZN(new_n25124_));
  NOR2_X1    g22032(.A1(new_n25124_), .A2(new_n6460_), .ZN(new_n25125_));
  NAND2_X1   g22033(.A1(new_n12776_), .A2(new_n24950_), .ZN(new_n25126_));
  NOR2_X1    g22034(.A1(new_n12322_), .A2(new_n5095_), .ZN(new_n25127_));
  AOI21_X1   g22035(.A1(new_n5095_), .A2(new_n12196_), .B(new_n25127_), .ZN(new_n25128_));
  OAI21_X1   g22036(.A1(new_n24950_), .A2(new_n25128_), .B(new_n25126_), .ZN(new_n25129_));
  OAI21_X1   g22037(.A1(new_n25129_), .A2(new_n5141_), .B(new_n2588_), .ZN(new_n25130_));
  NAND2_X1   g22038(.A1(new_n12913_), .A2(pi0661), .ZN(new_n25131_));
  AOI21_X1   g22039(.A1(new_n12911_), .A2(new_n25116_), .B(new_n25131_), .ZN(new_n25132_));
  NOR3_X1    g22040(.A1(new_n12362_), .A2(pi0661), .A3(new_n12731_), .ZN(new_n25133_));
  OAI22_X1   g22041(.A1(new_n25132_), .A2(new_n25133_), .B1(new_n12128_), .B2(new_n12782_), .ZN(new_n25134_));
  OAI21_X1   g22042(.A1(new_n12382_), .A2(new_n12907_), .B(new_n12374_), .ZN(new_n25135_));
  NOR2_X1    g22043(.A1(new_n25135_), .A2(new_n24950_), .ZN(new_n25136_));
  AOI21_X1   g22044(.A1(new_n24990_), .A2(new_n24950_), .B(new_n25136_), .ZN(new_n25137_));
  NAND4_X1   g22045(.A1(new_n25134_), .A2(new_n2588_), .A3(new_n5141_), .A4(new_n25137_), .ZN(new_n25138_));
  AND3_X2    g22046(.A1(new_n12939_), .A2(pi0661), .A3(new_n2597_), .Z(new_n25139_));
  NOR2_X1    g22047(.A1(new_n24950_), .A2(new_n5095_), .ZN(new_n25140_));
  AOI21_X1   g22048(.A1(new_n12944_), .A2(new_n25140_), .B(new_n6460_), .ZN(new_n25141_));
  NOR2_X1    g22049(.A1(new_n12326_), .A2(new_n11885_), .ZN(new_n25142_));
  INV_X1     g22050(.I(new_n25142_), .ZN(new_n25143_));
  NOR2_X1    g22051(.A1(new_n25143_), .A2(new_n24950_), .ZN(new_n25144_));
  NOR3_X1    g22052(.A1(new_n11885_), .A2(new_n24950_), .A3(new_n12133_), .ZN(new_n25145_));
  AOI21_X1   g22053(.A1(new_n25145_), .A2(new_n2588_), .B(pi0224), .ZN(new_n25146_));
  OAI21_X1   g22054(.A1(new_n25144_), .A2(new_n5141_), .B(new_n25146_), .ZN(new_n25147_));
  OAI21_X1   g22055(.A1(new_n25147_), .A2(new_n25141_), .B(new_n2604_), .ZN(new_n25148_));
  AOI21_X1   g22056(.A1(new_n25138_), .A2(new_n25139_), .B(new_n25148_), .ZN(new_n25149_));
  OAI21_X1   g22057(.A1(new_n25125_), .A2(new_n25130_), .B(new_n25149_), .ZN(new_n25150_));
  INV_X1     g22058(.I(new_n25077_), .ZN(new_n25151_));
  NAND2_X1   g22059(.A1(new_n25151_), .A2(new_n25145_), .ZN(new_n25152_));
  NAND2_X1   g22060(.A1(new_n25152_), .A2(new_n2566_), .ZN(new_n25153_));
  NOR2_X1    g22061(.A1(new_n25124_), .A2(new_n6445_), .ZN(new_n25154_));
  OAI21_X1   g22062(.A1(new_n25129_), .A2(new_n5094_), .B(new_n2588_), .ZN(new_n25155_));
  INV_X1     g22063(.I(new_n12944_), .ZN(new_n25156_));
  INV_X1     g22064(.I(new_n25140_), .ZN(new_n25157_));
  OAI21_X1   g22065(.A1(new_n25156_), .A2(new_n25157_), .B(new_n5094_), .ZN(new_n25158_));
  NOR2_X1    g22066(.A1(new_n25144_), .A2(new_n5094_), .ZN(new_n25159_));
  NOR2_X1    g22067(.A1(new_n25159_), .A2(pi0222), .ZN(new_n25160_));
  AOI21_X1   g22068(.A1(new_n25160_), .A2(new_n25158_), .B(new_n3284_), .ZN(new_n25161_));
  OAI21_X1   g22069(.A1(new_n25154_), .A2(new_n25155_), .B(new_n25161_), .ZN(new_n25162_));
  AND3_X2    g22070(.A1(new_n25137_), .A2(new_n2588_), .A3(new_n5094_), .Z(new_n25163_));
  NAND3_X1   g22071(.A1(new_n12951_), .A2(new_n2588_), .A3(pi0661), .ZN(new_n25164_));
  NAND2_X1   g22072(.A1(new_n25164_), .A2(pi0215), .ZN(new_n25165_));
  AOI21_X1   g22073(.A1(new_n25163_), .A2(new_n25134_), .B(new_n25165_), .ZN(new_n25166_));
  AOI21_X1   g22074(.A1(new_n25162_), .A2(new_n25153_), .B(new_n25166_), .ZN(new_n25167_));
  MUX2_X1    g22075(.I0(new_n25167_), .I1(new_n25150_), .S(new_n2587_), .Z(new_n25168_));
  MUX2_X1    g22076(.I0(new_n25157_), .I1(new_n2588_), .S(new_n12624_), .Z(new_n25169_));
  OAI21_X1   g22077(.A1(new_n12648_), .A2(new_n2588_), .B(new_n2587_), .ZN(new_n25170_));
  MUX2_X1    g22078(.I0(new_n25157_), .I1(new_n2588_), .S(new_n12630_), .Z(new_n25171_));
  OAI21_X1   g22079(.A1(new_n12655_), .A2(new_n2588_), .B(pi0299), .ZN(new_n25172_));
  OAI22_X1   g22080(.A1(new_n25169_), .A2(new_n25170_), .B1(new_n25171_), .B2(new_n25172_), .ZN(new_n25173_));
  AOI21_X1   g22081(.A1(new_n25173_), .A2(new_n3154_), .B(pi0038), .ZN(new_n25174_));
  OAI21_X1   g22082(.A1(new_n25168_), .A2(new_n3154_), .B(new_n25174_), .ZN(new_n25175_));
  NOR4_X1    g22083(.A1(new_n25087_), .A2(new_n24950_), .A3(new_n3231_), .A4(new_n17545_), .ZN(new_n25176_));
  AOI22_X1   g22084(.A1(new_n25175_), .A2(new_n25176_), .B1(pi0222), .B2(new_n3232_), .ZN(new_n25177_));
  NAND2_X1   g22085(.A1(new_n25177_), .A2(new_n11891_), .ZN(new_n25178_));
  NOR3_X1    g22086(.A1(new_n25177_), .A2(pi0625), .A3(new_n25022_), .ZN(new_n25179_));
  AOI21_X1   g22087(.A1(new_n25177_), .A2(new_n12970_), .B(new_n25020_), .ZN(new_n25180_));
  NOR3_X1    g22088(.A1(new_n25179_), .A2(new_n25180_), .A3(pi1153), .ZN(new_n25181_));
  NOR2_X1    g22089(.A1(new_n25181_), .A2(new_n11891_), .ZN(new_n25182_));
  XNOR2_X1   g22090(.A1(new_n25182_), .A2(new_n25178_), .ZN(new_n25183_));
  INV_X1     g22091(.I(new_n25183_), .ZN(new_n25184_));
  NOR2_X1    g22092(.A1(new_n25020_), .A2(new_n11938_), .ZN(new_n25185_));
  AOI21_X1   g22093(.A1(new_n25184_), .A2(new_n11938_), .B(new_n25185_), .ZN(new_n25186_));
  NOR2_X1    g22094(.A1(new_n25186_), .A2(new_n13714_), .ZN(new_n25187_));
  AOI21_X1   g22095(.A1(new_n13714_), .A2(new_n25022_), .B(new_n25187_), .ZN(new_n25188_));
  MUX2_X1    g22096(.I0(new_n25188_), .I1(new_n25020_), .S(new_n13713_), .Z(new_n25189_));
  AOI21_X1   g22097(.A1(new_n25189_), .A2(new_n12067_), .B(new_n25115_), .ZN(new_n25190_));
  MUX2_X1    g22098(.I0(new_n25190_), .I1(new_n25020_), .S(pi0647), .Z(new_n25191_));
  AOI21_X1   g22099(.A1(new_n25191_), .A2(new_n12049_), .B(new_n12060_), .ZN(new_n25192_));
  MUX2_X1    g22100(.I0(new_n25190_), .I1(new_n25020_), .S(new_n12061_), .Z(new_n25193_));
  AOI21_X1   g22101(.A1(new_n25193_), .A2(pi1157), .B(pi0630), .ZN(new_n25194_));
  OAI21_X1   g22102(.A1(new_n25192_), .A2(new_n25194_), .B(new_n12048_), .ZN(new_n25195_));
  AOI21_X1   g22103(.A1(new_n25114_), .A2(new_n15076_), .B(new_n25195_), .ZN(new_n25196_));
  OAI21_X1   g22104(.A1(new_n25020_), .A2(new_n12031_), .B(new_n12051_), .ZN(new_n25197_));
  AOI21_X1   g22105(.A1(new_n25189_), .A2(new_n12031_), .B(new_n25197_), .ZN(new_n25198_));
  INV_X1     g22106(.I(new_n25189_), .ZN(new_n25199_));
  NAND2_X1   g22107(.A1(new_n23402_), .A2(pi0628), .ZN(new_n25200_));
  OAI21_X1   g22108(.A1(new_n25199_), .A2(new_n25200_), .B(new_n17304_), .ZN(new_n25201_));
  OR3_X2     g22109(.A1(new_n25113_), .A2(new_n25198_), .A3(new_n25201_), .Z(new_n25202_));
  INV_X1     g22110(.I(new_n25188_), .ZN(new_n25203_));
  NOR3_X1    g22111(.A1(new_n25203_), .A2(new_n12013_), .A3(new_n25022_), .ZN(new_n25204_));
  AOI21_X1   g22112(.A1(new_n12014_), .A2(new_n25022_), .B(new_n25188_), .ZN(new_n25205_));
  OAI21_X1   g22113(.A1(new_n25204_), .A2(new_n25205_), .B(new_n12020_), .ZN(new_n25206_));
  AND3_X2    g22114(.A1(new_n25112_), .A2(new_n11994_), .A3(new_n25020_), .Z(new_n25207_));
  AOI21_X1   g22115(.A1(new_n11994_), .A2(new_n25022_), .B(new_n25112_), .ZN(new_n25208_));
  NOR2_X1    g22116(.A1(new_n25207_), .A2(new_n25208_), .ZN(new_n25209_));
  OAI21_X1   g22117(.A1(new_n25209_), .A2(new_n11990_), .B(new_n25206_), .ZN(new_n25210_));
  OAI21_X1   g22118(.A1(new_n25210_), .A2(new_n11998_), .B(new_n14732_), .ZN(new_n25211_));
  NAND2_X1   g22119(.A1(new_n25210_), .A2(pi0788), .ZN(new_n25212_));
  NOR2_X1    g22120(.A1(new_n3231_), .A2(pi0222), .ZN(new_n25213_));
  NOR2_X1    g22121(.A1(pi0661), .A2(pi0680), .ZN(new_n25214_));
  AOI21_X1   g22122(.A1(new_n12318_), .A2(new_n5108_), .B(new_n12303_), .ZN(new_n25215_));
  NOR2_X1    g22123(.A1(new_n25215_), .A2(new_n5101_), .ZN(new_n25216_));
  OAI21_X1   g22124(.A1(new_n12156_), .A2(new_n5101_), .B(new_n12417_), .ZN(new_n25217_));
  NOR2_X1    g22125(.A1(new_n25216_), .A2(new_n25217_), .ZN(new_n25218_));
  NAND2_X1   g22126(.A1(new_n25063_), .A2(new_n25215_), .ZN(new_n25219_));
  MUX2_X1    g22127(.I0(new_n25219_), .I1(new_n25218_), .S(pi0642), .Z(new_n25220_));
  NOR2_X1    g22128(.A1(new_n25220_), .A2(new_n5104_), .ZN(new_n25221_));
  INV_X1     g22129(.I(new_n25221_), .ZN(new_n25222_));
  NOR2_X1    g22130(.A1(new_n25215_), .A2(new_n12320_), .ZN(new_n25223_));
  NOR4_X1    g22131(.A1(new_n25219_), .A2(new_n12443_), .A3(pi0616), .A4(pi0680), .ZN(new_n25224_));
  NAND2_X1   g22132(.A1(new_n25222_), .A2(new_n25224_), .ZN(new_n25225_));
  NAND2_X1   g22133(.A1(new_n25225_), .A2(new_n25214_), .ZN(new_n25226_));
  AOI21_X1   g22134(.A1(new_n25226_), .A2(new_n25116_), .B(new_n25049_), .ZN(new_n25227_));
  AOI21_X1   g22135(.A1(new_n12128_), .A2(new_n25052_), .B(new_n25227_), .ZN(new_n25228_));
  NOR2_X1    g22136(.A1(new_n12448_), .A2(pi0616), .ZN(new_n25229_));
  NOR2_X1    g22137(.A1(new_n12331_), .A2(new_n12166_), .ZN(new_n25230_));
  NOR2_X1    g22138(.A1(new_n25230_), .A2(new_n5095_), .ZN(new_n25231_));
  AND3_X2    g22139(.A1(new_n25229_), .A2(new_n12387_), .A3(new_n25231_), .Z(new_n25232_));
  OAI21_X1   g22140(.A1(new_n25056_), .A2(pi0680), .B(pi0661), .ZN(new_n25233_));
  NOR2_X1    g22141(.A1(new_n25056_), .A2(new_n25116_), .ZN(new_n25234_));
  NOR2_X1    g22142(.A1(new_n25058_), .A2(new_n25234_), .ZN(new_n25235_));
  OAI21_X1   g22143(.A1(new_n25232_), .A2(new_n25233_), .B(new_n25235_), .ZN(new_n25236_));
  OAI21_X1   g22144(.A1(new_n25228_), .A2(new_n25236_), .B(new_n5094_), .ZN(new_n25237_));
  NOR4_X1    g22145(.A1(new_n12207_), .A2(new_n12166_), .A3(new_n5097_), .A4(new_n12127_), .ZN(new_n25238_));
  INV_X1     g22146(.I(new_n12226_), .ZN(new_n25239_));
  NAND2_X1   g22147(.A1(new_n12496_), .A2(pi0680), .ZN(new_n25240_));
  OAI21_X1   g22148(.A1(new_n25040_), .A2(pi0680), .B(pi0661), .ZN(new_n25241_));
  NAND4_X1   g22149(.A1(new_n25240_), .A2(pi0616), .A3(new_n25239_), .A4(new_n25241_), .ZN(new_n25242_));
  OAI21_X1   g22150(.A1(new_n25040_), .A2(new_n25116_), .B(new_n25242_), .ZN(new_n25243_));
  NOR2_X1    g22151(.A1(new_n25243_), .A2(new_n25238_), .ZN(new_n25244_));
  NOR2_X1    g22152(.A1(new_n25244_), .A2(new_n6445_), .ZN(new_n25245_));
  INV_X1     g22153(.I(new_n25064_), .ZN(new_n25246_));
  NOR3_X1    g22154(.A1(new_n25246_), .A2(pi0661), .A3(pi0680), .ZN(new_n25247_));
  NOR2_X1    g22155(.A1(new_n25246_), .A2(new_n25116_), .ZN(new_n25248_));
  NOR4_X1    g22156(.A1(new_n25247_), .A2(new_n25248_), .A3(new_n6445_), .A4(new_n25065_), .ZN(new_n25249_));
  NOR3_X1    g22157(.A1(new_n25245_), .A2(pi0222), .A3(new_n25249_), .ZN(new_n25250_));
  OAI21_X1   g22158(.A1(new_n25237_), .A2(new_n2588_), .B(new_n25250_), .ZN(new_n25251_));
  NOR2_X1    g22159(.A1(new_n25239_), .A2(new_n12166_), .ZN(new_n25252_));
  AOI21_X1   g22160(.A1(new_n12166_), .A2(new_n12477_), .B(new_n25252_), .ZN(new_n25253_));
  AOI21_X1   g22161(.A1(new_n25050_), .A2(new_n25157_), .B(new_n25253_), .ZN(new_n25254_));
  OAI21_X1   g22162(.A1(new_n25254_), .A2(new_n25151_), .B(new_n2566_), .ZN(new_n25255_));
  AOI21_X1   g22163(.A1(new_n25251_), .A2(new_n3285_), .B(new_n25255_), .ZN(new_n25256_));
  NOR3_X1    g22164(.A1(new_n25236_), .A2(pi0222), .A3(new_n6460_), .ZN(new_n25257_));
  NOR3_X1    g22165(.A1(new_n25247_), .A2(new_n25248_), .A3(new_n25065_), .ZN(new_n25258_));
  NAND4_X1   g22166(.A1(new_n25244_), .A2(new_n2595_), .A3(new_n5141_), .A4(new_n25258_), .ZN(new_n25259_));
  AND2_X2    g22167(.A1(new_n25253_), .A2(new_n25140_), .Z(new_n25260_));
  OAI21_X1   g22168(.A1(new_n25039_), .A2(new_n25140_), .B(new_n2588_), .ZN(new_n25261_));
  OAI21_X1   g22169(.A1(new_n25260_), .A2(new_n25261_), .B(new_n3300_), .ZN(new_n25262_));
  NAND2_X1   g22170(.A1(new_n25259_), .A2(new_n25262_), .ZN(new_n25263_));
  NAND2_X1   g22171(.A1(new_n25263_), .A2(new_n2604_), .ZN(new_n25264_));
  AOI21_X1   g22172(.A1(new_n25228_), .A2(new_n25257_), .B(new_n25264_), .ZN(new_n25265_));
  NOR2_X1    g22173(.A1(new_n25036_), .A2(new_n25116_), .ZN(new_n25266_));
  AOI21_X1   g22174(.A1(new_n12302_), .A2(new_n12304_), .B(new_n12320_), .ZN(new_n25267_));
  INV_X1     g22175(.I(new_n25267_), .ZN(new_n25268_));
  NAND2_X1   g22176(.A1(new_n24950_), .A2(new_n5095_), .ZN(new_n25270_));
  NOR2_X1    g22177(.A1(new_n25036_), .A2(new_n25270_), .ZN(new_n25271_));
  NOR3_X1    g22178(.A1(new_n25266_), .A2(new_n25271_), .A3(new_n25035_), .ZN(new_n25272_));
  NAND2_X1   g22179(.A1(new_n12389_), .A2(new_n25231_), .ZN(new_n25273_));
  AOI21_X1   g22180(.A1(new_n25026_), .A2(new_n5095_), .B(new_n24950_), .ZN(new_n25274_));
  OAI21_X1   g22181(.A1(pi0661), .A2(new_n12731_), .B(new_n25026_), .ZN(new_n25275_));
  NAND2_X1   g22182(.A1(new_n25275_), .A2(new_n25029_), .ZN(new_n25276_));
  AOI21_X1   g22183(.A1(new_n25273_), .A2(new_n25274_), .B(new_n25276_), .ZN(new_n25277_));
  XOR2_X1    g22184(.A1(new_n25277_), .A2(new_n25272_), .Z(new_n25278_));
  NAND2_X1   g22185(.A1(new_n25278_), .A2(new_n5141_), .ZN(new_n25279_));
  XOR2_X1    g22186(.A1(new_n25279_), .A2(new_n25272_), .Z(new_n25280_));
  NAND2_X1   g22187(.A1(new_n25280_), .A2(pi0222), .ZN(new_n25281_));
  INV_X1     g22188(.I(new_n12475_), .ZN(new_n25282_));
  AOI21_X1   g22189(.A1(new_n25282_), .A2(new_n25157_), .B(new_n25043_), .ZN(new_n25283_));
  INV_X1     g22190(.I(new_n25283_), .ZN(new_n25284_));
  NOR2_X1    g22191(.A1(new_n12250_), .A2(new_n12258_), .ZN(new_n25285_));
  AOI21_X1   g22192(.A1(new_n25285_), .A2(pi0616), .B(new_n5095_), .ZN(new_n25286_));
  NAND2_X1   g22193(.A1(new_n12470_), .A2(new_n25286_), .ZN(new_n25287_));
  INV_X1     g22194(.I(new_n12250_), .ZN(new_n25288_));
  NOR4_X1    g22195(.A1(new_n25288_), .A2(new_n12166_), .A3(pi0661), .A4(pi0680), .ZN(new_n25289_));
  NOR2_X1    g22196(.A1(new_n12262_), .A2(new_n25040_), .ZN(new_n25290_));
  NOR2_X1    g22197(.A1(new_n25288_), .A2(new_n12166_), .ZN(new_n25291_));
  OAI22_X1   g22198(.A1(new_n25291_), .A2(pi0661), .B1(new_n5217_), .B2(new_n25290_), .ZN(new_n25292_));
  AOI21_X1   g22199(.A1(new_n25287_), .A2(new_n25289_), .B(new_n25292_), .ZN(new_n25293_));
  NAND3_X1   g22200(.A1(new_n25293_), .A2(new_n6460_), .A3(new_n25284_), .ZN(new_n25294_));
  OAI21_X1   g22201(.A1(new_n25293_), .A2(new_n5141_), .B(new_n25283_), .ZN(new_n25295_));
  AND3_X2    g22202(.A1(new_n25295_), .A2(new_n25294_), .A3(new_n2588_), .Z(new_n25296_));
  AOI21_X1   g22203(.A1(new_n25281_), .A2(new_n25296_), .B(pi0223), .ZN(new_n25297_));
  OAI21_X1   g22204(.A1(new_n25297_), .A2(pi0299), .B(new_n3154_), .ZN(new_n25298_));
  NAND2_X1   g22205(.A1(new_n25278_), .A2(new_n5094_), .ZN(new_n25299_));
  XOR2_X1    g22206(.A1(new_n25299_), .A2(new_n25272_), .Z(new_n25300_));
  NAND2_X1   g22207(.A1(new_n25300_), .A2(pi0222), .ZN(new_n25301_));
  NAND3_X1   g22208(.A1(new_n25293_), .A2(new_n6445_), .A3(new_n25284_), .ZN(new_n25302_));
  OAI21_X1   g22209(.A1(new_n25293_), .A2(new_n5094_), .B(new_n25283_), .ZN(new_n25303_));
  AND3_X2    g22210(.A1(new_n25303_), .A2(new_n25302_), .A3(new_n2588_), .Z(new_n25304_));
  AOI21_X1   g22211(.A1(new_n25301_), .A2(new_n25304_), .B(new_n24682_), .ZN(new_n25305_));
  OAI21_X1   g22212(.A1(new_n25298_), .A2(new_n25265_), .B(new_n25305_), .ZN(new_n25306_));
  OAI21_X1   g22213(.A1(new_n13830_), .A2(new_n12166_), .B(new_n2588_), .ZN(new_n25307_));
  NAND3_X1   g22214(.A1(new_n13829_), .A2(pi0661), .A3(new_n25307_), .ZN(new_n25308_));
  NAND2_X1   g22215(.A1(new_n12627_), .A2(pi0665), .ZN(new_n25309_));
  MUX2_X1    g22216(.I0(new_n25309_), .I1(new_n12655_), .S(new_n5101_), .Z(new_n25310_));
  OAI21_X1   g22217(.A1(pi0616), .A2(new_n13830_), .B(new_n25310_), .ZN(new_n25311_));
  NAND4_X1   g22218(.A1(new_n25311_), .A2(new_n2588_), .A3(new_n13358_), .A4(new_n25157_), .ZN(new_n25312_));
  NAND3_X1   g22219(.A1(new_n25312_), .A2(pi0299), .A3(new_n25308_), .ZN(new_n25313_));
  NAND2_X1   g22220(.A1(new_n12619_), .A2(pi0665), .ZN(new_n25314_));
  MUX2_X1    g22221(.I0(new_n25314_), .I1(new_n12648_), .S(new_n5101_), .Z(new_n25315_));
  OAI21_X1   g22222(.A1(pi0616), .A2(new_n13858_), .B(new_n25315_), .ZN(new_n25316_));
  NAND4_X1   g22223(.A1(new_n25316_), .A2(new_n2588_), .A3(new_n13355_), .A4(new_n25157_), .ZN(new_n25317_));
  NAND2_X1   g22224(.A1(new_n12610_), .A2(pi0616), .ZN(new_n25318_));
  AOI21_X1   g22225(.A1(new_n25318_), .A2(new_n2588_), .B(new_n24950_), .ZN(new_n25319_));
  AOI21_X1   g22226(.A1(new_n13844_), .A2(new_n25319_), .B(pi0299), .ZN(new_n25320_));
  AOI21_X1   g22227(.A1(new_n25317_), .A2(new_n25320_), .B(pi0039), .ZN(new_n25321_));
  AOI21_X1   g22228(.A1(new_n25313_), .A2(new_n25321_), .B(pi0038), .ZN(new_n25326_));
  OAI21_X1   g22229(.A1(new_n25306_), .A2(new_n25256_), .B(new_n25326_), .ZN(new_n25327_));
  NAND2_X1   g22230(.A1(new_n25327_), .A2(new_n3231_), .ZN(new_n25328_));
  XOR2_X1    g22231(.A1(new_n25328_), .A2(new_n25213_), .Z(new_n25329_));
  OAI21_X1   g22232(.A1(new_n25329_), .A2(pi0625), .B(new_n25094_), .ZN(new_n25330_));
  INV_X1     g22233(.I(new_n25094_), .ZN(new_n25331_));
  NAND3_X1   g22234(.A1(new_n25329_), .A2(new_n12970_), .A3(new_n25331_), .ZN(new_n25332_));
  NAND3_X1   g22235(.A1(new_n25330_), .A2(new_n25332_), .A3(new_n12977_), .ZN(new_n25333_));
  NAND2_X1   g22236(.A1(new_n25329_), .A2(pi0625), .ZN(new_n25334_));
  NAND3_X1   g22237(.A1(new_n25334_), .A2(new_n13434_), .A3(new_n25331_), .ZN(new_n25335_));
  NAND2_X1   g22238(.A1(new_n25335_), .A2(new_n25181_), .ZN(new_n25336_));
  NAND2_X1   g22239(.A1(new_n25336_), .A2(new_n13657_), .ZN(new_n25337_));
  NAND2_X1   g22240(.A1(new_n25337_), .A2(new_n25333_), .ZN(new_n25338_));
  NOR2_X1    g22241(.A1(new_n25329_), .A2(pi0778), .ZN(new_n25339_));
  AOI21_X1   g22242(.A1(new_n25338_), .A2(pi0778), .B(new_n25339_), .ZN(new_n25340_));
  NOR4_X1    g22243(.A1(new_n25340_), .A2(new_n11903_), .A3(pi1155), .A4(new_n25184_), .ZN(new_n25341_));
  NAND2_X1   g22244(.A1(new_n25100_), .A2(pi0660), .ZN(new_n25342_));
  NOR3_X1    g22245(.A1(new_n25183_), .A2(new_n11903_), .A3(new_n11912_), .ZN(new_n25343_));
  OAI22_X1   g22246(.A1(new_n25341_), .A2(new_n25342_), .B1(pi0660), .B2(new_n25343_), .ZN(new_n25344_));
  MUX2_X1    g22247(.I0(new_n25344_), .I1(new_n25340_), .S(new_n11870_), .Z(new_n25345_));
  OAI21_X1   g22248(.A1(new_n25186_), .A2(pi0618), .B(pi1154), .ZN(new_n25346_));
  NAND2_X1   g22249(.A1(new_n25105_), .A2(pi0627), .ZN(new_n25347_));
  NAND4_X1   g22250(.A1(new_n25345_), .A2(pi0618), .A3(new_n25346_), .A4(new_n25347_), .ZN(new_n25348_));
  AND2_X2    g22251(.A1(new_n25345_), .A2(new_n11934_), .Z(new_n25349_));
  OAI21_X1   g22252(.A1(new_n25186_), .A2(new_n11934_), .B(new_n11960_), .ZN(new_n25350_));
  OAI21_X1   g22253(.A1(new_n25349_), .A2(new_n25350_), .B(new_n25348_), .ZN(new_n25351_));
  MUX2_X1    g22254(.I0(new_n25351_), .I1(new_n25345_), .S(new_n11969_), .Z(new_n25352_));
  NOR3_X1    g22255(.A1(new_n25188_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n25353_));
  NOR2_X1    g22256(.A1(new_n25353_), .A2(pi0648), .ZN(new_n25354_));
  NOR4_X1    g22257(.A1(new_n25352_), .A2(new_n11967_), .A3(pi1159), .A4(new_n25203_), .ZN(new_n25355_));
  NOR2_X1    g22258(.A1(new_n25355_), .A2(new_n25110_), .ZN(new_n25356_));
  NOR2_X1    g22259(.A1(new_n25352_), .A2(pi0789), .ZN(new_n25357_));
  NOR4_X1    g22260(.A1(new_n25356_), .A2(new_n17371_), .A3(new_n25354_), .A4(new_n25357_), .ZN(new_n25358_));
  NAND3_X1   g22261(.A1(new_n25358_), .A2(new_n25211_), .A3(new_n25212_), .ZN(new_n25359_));
  AOI21_X1   g22262(.A1(new_n25359_), .A2(new_n25202_), .B(new_n14725_), .ZN(new_n25360_));
  NOR2_X1    g22263(.A1(new_n25360_), .A2(new_n25196_), .ZN(new_n25361_));
  NAND2_X1   g22264(.A1(new_n25114_), .A2(new_n12092_), .ZN(new_n25362_));
  AOI21_X1   g22265(.A1(new_n25020_), .A2(new_n12091_), .B(new_n12082_), .ZN(new_n25363_));
  NAND2_X1   g22266(.A1(new_n25362_), .A2(new_n25363_), .ZN(new_n25364_));
  OAI21_X1   g22267(.A1(new_n12082_), .A2(new_n25022_), .B(new_n25364_), .ZN(new_n25365_));
  AOI21_X1   g22268(.A1(new_n25365_), .A2(pi0715), .B(pi1160), .ZN(new_n25366_));
  NAND2_X1   g22269(.A1(new_n25191_), .A2(new_n12049_), .ZN(new_n25367_));
  NAND2_X1   g22270(.A1(new_n25193_), .A2(pi1157), .ZN(new_n25368_));
  NAND2_X1   g22271(.A1(new_n25367_), .A2(new_n25368_), .ZN(new_n25369_));
  MUX2_X1    g22272(.I0(new_n25369_), .I1(new_n25190_), .S(new_n12048_), .Z(new_n25370_));
  NOR4_X1    g22273(.A1(new_n25361_), .A2(pi0644), .A3(new_n12099_), .A4(new_n25366_), .ZN(new_n25372_));
  AOI21_X1   g22274(.A1(new_n25370_), .A2(new_n12082_), .B(new_n12099_), .ZN(new_n25373_));
  AOI21_X1   g22275(.A1(new_n25022_), .A2(new_n12082_), .B(pi0715), .ZN(new_n25374_));
  AOI21_X1   g22276(.A1(new_n25364_), .A2(new_n25374_), .B(new_n12081_), .ZN(new_n25375_));
  NOR4_X1    g22277(.A1(new_n25361_), .A2(new_n12082_), .A3(new_n25373_), .A4(new_n25375_), .ZN(new_n25376_));
  NOR2_X1    g22278(.A1(new_n25372_), .A2(new_n25376_), .ZN(new_n25377_));
  MUX2_X1    g22279(.I0(new_n25377_), .I1(new_n25361_), .S(new_n11867_), .Z(new_n25378_));
  NAND2_X1   g22280(.A1(po1038), .A2(pi0222), .ZN(new_n25379_));
  OAI21_X1   g22281(.A1(new_n25378_), .A2(po1038), .B(new_n25379_), .ZN(po0379));
  AOI21_X1   g22282(.A1(new_n15389_), .A2(new_n2587_), .B(new_n3154_), .ZN(new_n25381_));
  NAND2_X1   g22283(.A1(new_n12780_), .A2(new_n25381_), .ZN(new_n25382_));
  NOR4_X1    g22284(.A1(new_n13384_), .A2(pi0223), .A3(new_n10843_), .A4(new_n13972_), .ZN(new_n25383_));
  NAND2_X1   g22285(.A1(new_n25383_), .A2(new_n25382_), .ZN(new_n25384_));
  INV_X1     g22286(.I(new_n25384_), .ZN(new_n25385_));
  NOR2_X1    g22287(.A1(new_n25385_), .A2(new_n12054_), .ZN(new_n25386_));
  NOR2_X1    g22288(.A1(new_n25384_), .A2(new_n14624_), .ZN(new_n25387_));
  NOR2_X1    g22289(.A1(new_n25384_), .A2(new_n11924_), .ZN(new_n25388_));
  NOR2_X1    g22290(.A1(new_n3231_), .A2(pi0223), .ZN(new_n25389_));
  INV_X1     g22291(.I(new_n25389_), .ZN(new_n25390_));
  AOI21_X1   g22292(.A1(pi0039), .A2(pi0223), .B(new_n3172_), .ZN(new_n25391_));
  INV_X1     g22293(.I(new_n25391_), .ZN(new_n25392_));
  OAI21_X1   g22294(.A1(new_n12109_), .A2(pi0223), .B(new_n3154_), .ZN(new_n25393_));
  NOR2_X1    g22295(.A1(new_n11875_), .A2(new_n12384_), .ZN(new_n25394_));
  NOR2_X1    g22296(.A1(new_n12110_), .A2(new_n25394_), .ZN(new_n25395_));
  NOR2_X1    g22297(.A1(new_n25395_), .A2(new_n25393_), .ZN(new_n25396_));
  AOI21_X1   g22298(.A1(new_n12133_), .A2(pi0223), .B(new_n3285_), .ZN(new_n25397_));
  NOR2_X1    g22299(.A1(new_n12209_), .A2(new_n12384_), .ZN(new_n25398_));
  INV_X1     g22300(.I(new_n25398_), .ZN(new_n25399_));
  NOR2_X1    g22301(.A1(new_n25399_), .A2(new_n25397_), .ZN(new_n25400_));
  NOR2_X1    g22302(.A1(new_n24795_), .A2(new_n25394_), .ZN(new_n25401_));
  INV_X1     g22303(.I(new_n24792_), .ZN(new_n25402_));
  AOI21_X1   g22304(.A1(new_n25402_), .A2(new_n12287_), .B(new_n12384_), .ZN(new_n25403_));
  AOI21_X1   g22305(.A1(new_n25403_), .A2(new_n5104_), .B(new_n25401_), .ZN(new_n25404_));
  NAND2_X1   g22306(.A1(new_n25404_), .A2(pi0681), .ZN(new_n25405_));
  INV_X1     g22307(.I(new_n25404_), .ZN(new_n25406_));
  AOI21_X1   g22308(.A1(pi0642), .A2(new_n12217_), .B(new_n12231_), .ZN(new_n25407_));
  MUX2_X1    g22309(.I0(new_n25407_), .I1(new_n25406_), .S(new_n5099_), .Z(new_n25408_));
  OAI21_X1   g22310(.A1(new_n25408_), .A2(pi0681), .B(new_n5094_), .ZN(new_n25409_));
  INV_X1     g22311(.I(new_n25409_), .ZN(new_n25410_));
  NOR2_X1    g22312(.A1(new_n12326_), .A2(pi0642), .ZN(new_n25411_));
  AOI21_X1   g22313(.A1(pi0642), .A2(new_n12489_), .B(new_n25411_), .ZN(new_n25412_));
  INV_X1     g22314(.I(new_n25412_), .ZN(new_n25413_));
  NOR4_X1    g22315(.A1(new_n12191_), .A2(pi0681), .A3(new_n5098_), .A4(new_n25394_), .ZN(new_n25414_));
  AOI21_X1   g22316(.A1(new_n25413_), .A2(new_n25414_), .B(new_n5094_), .ZN(new_n25415_));
  NOR2_X1    g22317(.A1(new_n25413_), .A2(new_n12731_), .ZN(new_n25416_));
  OAI21_X1   g22318(.A1(new_n25415_), .A2(new_n25416_), .B(pi0223), .ZN(new_n25417_));
  AOI21_X1   g22319(.A1(new_n25410_), .A2(new_n25405_), .B(new_n25417_), .ZN(new_n25418_));
  NOR3_X1    g22320(.A1(new_n5099_), .A2(new_n12384_), .A3(pi0681), .ZN(new_n25419_));
  INV_X1     g22321(.I(new_n25419_), .ZN(new_n25420_));
  NOR2_X1    g22322(.A1(new_n12207_), .A2(new_n25420_), .ZN(new_n25421_));
  AOI21_X1   g22323(.A1(new_n12731_), .A2(new_n25398_), .B(new_n25421_), .ZN(new_n25422_));
  OR2_X2     g22324(.A1(new_n25422_), .A2(new_n15315_), .Z(new_n25423_));
  INV_X1     g22325(.I(new_n25394_), .ZN(new_n25424_));
  NAND2_X1   g22326(.A1(new_n12157_), .A2(new_n5099_), .ZN(new_n25425_));
  NAND3_X1   g22327(.A1(new_n12425_), .A2(pi0642), .A3(new_n5098_), .ZN(new_n25426_));
  NAND4_X1   g22328(.A1(new_n25425_), .A2(new_n12731_), .A3(new_n25424_), .A4(new_n25426_), .ZN(new_n25427_));
  INV_X1     g22329(.I(new_n25427_), .ZN(new_n25428_));
  AOI21_X1   g22330(.A1(new_n12157_), .A2(new_n25394_), .B(new_n12731_), .ZN(new_n25429_));
  NOR2_X1    g22331(.A1(new_n25428_), .A2(new_n25429_), .ZN(new_n25430_));
  NAND2_X1   g22332(.A1(new_n25430_), .A2(new_n5473_), .ZN(new_n25431_));
  NOR2_X1    g22333(.A1(new_n25430_), .A2(new_n15315_), .ZN(new_n25432_));
  NAND2_X1   g22334(.A1(new_n2604_), .A2(new_n5473_), .ZN(new_n25433_));
  NOR3_X1    g22335(.A1(new_n25432_), .A2(new_n3284_), .A3(new_n25433_), .ZN(new_n25434_));
  NAND3_X1   g22336(.A1(new_n25423_), .A2(new_n25431_), .A3(new_n25434_), .ZN(new_n25435_));
  OAI22_X1   g22337(.A1(new_n25418_), .A2(new_n25435_), .B1(pi0215), .B2(new_n25400_), .ZN(new_n25436_));
  NOR2_X1    g22338(.A1(new_n12310_), .A2(new_n12384_), .ZN(new_n25437_));
  AOI21_X1   g22339(.A1(new_n12362_), .A2(new_n12384_), .B(new_n25437_), .ZN(new_n25438_));
  AOI21_X1   g22340(.A1(pi0642), .A2(new_n12308_), .B(new_n12262_), .ZN(new_n25439_));
  NOR2_X1    g22341(.A1(new_n25439_), .A2(new_n5098_), .ZN(new_n25440_));
  OAI22_X1   g22342(.A1(new_n25438_), .A2(new_n5098_), .B1(pi0681), .B2(new_n25440_), .ZN(new_n25441_));
  NAND2_X1   g22343(.A1(new_n25441_), .A2(new_n6445_), .ZN(new_n25442_));
  NOR4_X1    g22344(.A1(new_n12725_), .A2(new_n5099_), .A3(new_n12110_), .A4(new_n25394_), .ZN(new_n25443_));
  OAI21_X1   g22345(.A1(new_n12384_), .A2(new_n12286_), .B(new_n25026_), .ZN(new_n25444_));
  OAI21_X1   g22346(.A1(new_n24795_), .A2(new_n25394_), .B(new_n25444_), .ZN(new_n25445_));
  OAI21_X1   g22347(.A1(new_n12731_), .A2(new_n5098_), .B(new_n25445_), .ZN(new_n25446_));
  OAI21_X1   g22348(.A1(new_n12731_), .A2(new_n25443_), .B(new_n25446_), .ZN(new_n25447_));
  AOI21_X1   g22349(.A1(new_n25447_), .A2(new_n5094_), .B(pi0223), .ZN(new_n25448_));
  OAI21_X1   g22350(.A1(new_n25439_), .A2(new_n5098_), .B(new_n12731_), .ZN(new_n25449_));
  NOR2_X1    g22351(.A1(new_n12375_), .A2(new_n25420_), .ZN(new_n25450_));
  AOI21_X1   g22352(.A1(new_n12249_), .A2(new_n25449_), .B(new_n25450_), .ZN(new_n25451_));
  NOR4_X1    g22353(.A1(new_n25451_), .A2(new_n12384_), .A3(pi0681), .A4(new_n25288_), .ZN(new_n25452_));
  NOR2_X1    g22354(.A1(new_n25452_), .A2(new_n5473_), .ZN(new_n25453_));
  NAND2_X1   g22355(.A1(new_n25452_), .A2(new_n15315_), .ZN(new_n25454_));
  NOR2_X1    g22356(.A1(new_n25450_), .A2(new_n6445_), .ZN(new_n25455_));
  AOI21_X1   g22357(.A1(new_n25455_), .A2(new_n25398_), .B(new_n25433_), .ZN(new_n25456_));
  NAND2_X1   g22358(.A1(new_n25454_), .A2(new_n25456_), .ZN(new_n25457_));
  OAI21_X1   g22359(.A1(new_n25457_), .A2(new_n25453_), .B(new_n4905_), .ZN(new_n25458_));
  AOI21_X1   g22360(.A1(new_n25448_), .A2(new_n25442_), .B(new_n25458_), .ZN(new_n25459_));
  NAND2_X1   g22361(.A1(new_n25441_), .A2(new_n6460_), .ZN(new_n25460_));
  NAND2_X1   g22362(.A1(new_n25447_), .A2(new_n5141_), .ZN(new_n25461_));
  NAND3_X1   g22363(.A1(new_n25461_), .A2(new_n25460_), .A3(new_n2604_), .ZN(new_n25462_));
  NOR2_X1    g22364(.A1(new_n25422_), .A2(new_n6460_), .ZN(new_n25463_));
  OAI21_X1   g22365(.A1(new_n25430_), .A2(new_n6460_), .B(new_n3155_), .ZN(new_n25464_));
  AOI21_X1   g22366(.A1(new_n25398_), .A2(new_n3155_), .B(pi0223), .ZN(new_n25465_));
  OAI21_X1   g22367(.A1(new_n25463_), .A2(new_n25464_), .B(new_n25465_), .ZN(new_n25466_));
  NAND3_X1   g22368(.A1(new_n25462_), .A2(new_n2587_), .A3(new_n25466_), .ZN(new_n25467_));
  AOI21_X1   g22369(.A1(new_n25436_), .A2(new_n25459_), .B(new_n25467_), .ZN(new_n25468_));
  NAND2_X1   g22370(.A1(new_n12613_), .A2(new_n5102_), .ZN(new_n25469_));
  AND2_X2    g22371(.A1(new_n13837_), .A2(new_n25469_), .Z(new_n25470_));
  NOR3_X1    g22372(.A1(new_n13830_), .A2(new_n12384_), .A3(new_n3294_), .ZN(new_n25471_));
  NOR3_X1    g22373(.A1(new_n25470_), .A2(pi0223), .A3(new_n25471_), .ZN(new_n25472_));
  NAND2_X1   g22374(.A1(new_n2604_), .A2(pi0642), .ZN(new_n25473_));
  OAI21_X1   g22375(.A1(new_n13858_), .A2(new_n25473_), .B(new_n2587_), .ZN(new_n25474_));
  OAI21_X1   g22376(.A1(new_n13858_), .A2(pi0642), .B(pi0223), .ZN(new_n25475_));
  OAI21_X1   g22377(.A1(new_n13859_), .A2(new_n25475_), .B(new_n25474_), .ZN(new_n25476_));
  NAND2_X1   g22378(.A1(new_n25476_), .A2(new_n3154_), .ZN(new_n25477_));
  OAI21_X1   g22379(.A1(new_n25477_), .A2(new_n25472_), .B(new_n3172_), .ZN(new_n25478_));
  NAND2_X1   g22380(.A1(new_n25478_), .A2(new_n3154_), .ZN(new_n25479_));
  OAI22_X1   g22381(.A1(new_n25479_), .A2(new_n25468_), .B1(new_n25392_), .B2(new_n25396_), .ZN(new_n25480_));
  NAND2_X1   g22382(.A1(new_n25480_), .A2(new_n3231_), .ZN(new_n25481_));
  XOR2_X1    g22383(.A1(new_n25481_), .A2(new_n25390_), .Z(new_n25482_));
  AOI21_X1   g22384(.A1(new_n25482_), .A2(new_n11924_), .B(new_n25388_), .ZN(new_n25483_));
  MUX2_X1    g22385(.I0(new_n25483_), .I1(new_n25384_), .S(pi0609), .Z(new_n25484_));
  NOR2_X1    g22386(.A1(new_n25484_), .A2(pi1155), .ZN(new_n25485_));
  MUX2_X1    g22387(.I0(new_n25483_), .I1(new_n25384_), .S(new_n11903_), .Z(new_n25486_));
  NOR2_X1    g22388(.A1(new_n25486_), .A2(new_n11912_), .ZN(new_n25487_));
  NOR2_X1    g22389(.A1(new_n25485_), .A2(new_n25487_), .ZN(new_n25488_));
  MUX2_X1    g22390(.I0(new_n25488_), .I1(new_n25483_), .S(new_n11870_), .Z(new_n25489_));
  NAND2_X1   g22391(.A1(new_n25489_), .A2(new_n11969_), .ZN(new_n25490_));
  NOR3_X1    g22392(.A1(new_n25489_), .A2(pi0618), .A3(new_n25384_), .ZN(new_n25491_));
  AOI21_X1   g22393(.A1(new_n25489_), .A2(new_n11934_), .B(new_n25385_), .ZN(new_n25492_));
  NOR3_X1    g22394(.A1(new_n25491_), .A2(new_n25492_), .A3(pi1154), .ZN(new_n25493_));
  NOR2_X1    g22395(.A1(new_n25493_), .A2(new_n11969_), .ZN(new_n25494_));
  XOR2_X1    g22396(.A1(new_n25494_), .A2(new_n25490_), .Z(new_n25495_));
  INV_X1     g22397(.I(new_n25495_), .ZN(new_n25496_));
  NAND3_X1   g22398(.A1(new_n25495_), .A2(new_n11967_), .A3(new_n25385_), .ZN(new_n25497_));
  OAI21_X1   g22399(.A1(new_n25495_), .A2(pi0619), .B(new_n25384_), .ZN(new_n25498_));
  NAND3_X1   g22400(.A1(new_n25498_), .A2(new_n25497_), .A3(new_n11869_), .ZN(new_n25499_));
  MUX2_X1    g22401(.I0(new_n25499_), .I1(new_n25496_), .S(new_n11985_), .Z(new_n25500_));
  AOI21_X1   g22402(.A1(new_n25500_), .A2(new_n14624_), .B(new_n25387_), .ZN(new_n25501_));
  AOI21_X1   g22403(.A1(new_n25501_), .A2(new_n12054_), .B(new_n25386_), .ZN(new_n25502_));
  NOR2_X1    g22404(.A1(new_n25385_), .A2(new_n12067_), .ZN(new_n25503_));
  NOR2_X1    g22405(.A1(new_n25385_), .A2(new_n11961_), .ZN(new_n25504_));
  NOR2_X1    g22406(.A1(new_n25384_), .A2(new_n11938_), .ZN(new_n25505_));
  NAND2_X1   g22407(.A1(new_n13402_), .A2(pi0681), .ZN(new_n25506_));
  AOI21_X1   g22408(.A1(new_n13368_), .A2(pi0223), .B(new_n3172_), .ZN(new_n25507_));
  NOR2_X1    g22409(.A1(new_n5095_), .A2(new_n12731_), .ZN(new_n25508_));
  NAND3_X1   g22410(.A1(new_n12641_), .A2(new_n2604_), .A3(new_n25508_), .ZN(new_n25509_));
  OAI21_X1   g22411(.A1(new_n12630_), .A2(new_n25508_), .B(pi0223), .ZN(new_n25510_));
  OAI21_X1   g22412(.A1(new_n12655_), .A2(new_n2604_), .B(pi0299), .ZN(new_n25511_));
  AOI21_X1   g22413(.A1(new_n25509_), .A2(new_n25510_), .B(new_n25511_), .ZN(new_n25512_));
  INV_X1     g22414(.I(new_n25508_), .ZN(new_n25513_));
  MUX2_X1    g22415(.I0(new_n25513_), .I1(new_n2604_), .S(new_n12624_), .Z(new_n25514_));
  OAI21_X1   g22416(.A1(new_n12648_), .A2(new_n2604_), .B(new_n2587_), .ZN(new_n25515_));
  OAI21_X1   g22417(.A1(new_n25514_), .A2(new_n25515_), .B(new_n3154_), .ZN(new_n25516_));
  INV_X1     g22418(.I(new_n25397_), .ZN(new_n25517_));
  NAND3_X1   g22419(.A1(new_n12871_), .A2(new_n12731_), .A3(new_n12873_), .ZN(new_n25518_));
  OR2_X2     g22420(.A1(new_n25118_), .A2(new_n12731_), .Z(new_n25519_));
  NOR3_X1    g22421(.A1(new_n12774_), .A2(pi0681), .A3(new_n12760_), .ZN(new_n25520_));
  NOR2_X1    g22422(.A1(new_n12731_), .A2(pi0223), .ZN(new_n25521_));
  NAND2_X1   g22423(.A1(new_n25128_), .A2(new_n25521_), .ZN(new_n25522_));
  OAI21_X1   g22424(.A1(new_n25522_), .A2(new_n25520_), .B(new_n6445_), .ZN(new_n25523_));
  AOI21_X1   g22425(.A1(new_n25519_), .A2(new_n25518_), .B(new_n25523_), .ZN(new_n25524_));
  NAND2_X1   g22426(.A1(new_n12944_), .A2(new_n25508_), .ZN(new_n25525_));
  INV_X1     g22427(.I(new_n25525_), .ZN(new_n25526_));
  NOR2_X1    g22428(.A1(new_n25526_), .A2(new_n6445_), .ZN(new_n25527_));
  NOR2_X1    g22429(.A1(new_n25143_), .A2(new_n12731_), .ZN(new_n25528_));
  OAI21_X1   g22430(.A1(new_n25528_), .A2(new_n5094_), .B(new_n2604_), .ZN(new_n25529_));
  OAI21_X1   g22431(.A1(new_n25529_), .A2(new_n25527_), .B(new_n3285_), .ZN(new_n25530_));
  NOR3_X1    g22432(.A1(new_n11885_), .A2(new_n12731_), .A3(new_n12133_), .ZN(new_n25531_));
  OAI22_X1   g22433(.A1(new_n25524_), .A2(new_n25530_), .B1(new_n25517_), .B2(new_n25531_), .ZN(new_n25532_));
  NAND3_X1   g22434(.A1(new_n12362_), .A2(pi0661), .A3(pi0681), .ZN(new_n25533_));
  NAND2_X1   g22435(.A1(new_n12913_), .A2(pi0681), .ZN(new_n25534_));
  NAND2_X1   g22436(.A1(new_n25534_), .A2(new_n25533_), .ZN(new_n25535_));
  MUX2_X1    g22437(.I0(new_n25135_), .I1(new_n12728_), .S(new_n12731_), .Z(new_n25536_));
  AOI21_X1   g22438(.A1(new_n12951_), .A2(new_n25521_), .B(new_n2566_), .ZN(new_n25537_));
  NOR4_X1    g22439(.A1(new_n25536_), .A2(new_n3294_), .A3(new_n6445_), .A4(new_n25537_), .ZN(new_n25538_));
  NAND2_X1   g22440(.A1(new_n25538_), .A2(new_n25535_), .ZN(new_n25539_));
  AOI21_X1   g22441(.A1(new_n25532_), .A2(new_n2566_), .B(new_n25539_), .ZN(new_n25540_));
  OAI21_X1   g22442(.A1(new_n25535_), .A2(new_n25536_), .B(new_n5141_), .ZN(new_n25541_));
  NOR2_X1    g22443(.A1(new_n25541_), .A2(new_n2604_), .ZN(new_n25542_));
  OAI21_X1   g22444(.A1(new_n5141_), .A2(new_n25528_), .B(new_n25526_), .ZN(new_n25543_));
  NAND3_X1   g22445(.A1(new_n25528_), .A2(new_n6460_), .A3(new_n25525_), .ZN(new_n25544_));
  NAND2_X1   g22446(.A1(new_n2588_), .A2(new_n2595_), .ZN(new_n25545_));
  AND3_X2    g22447(.A1(new_n25543_), .A2(new_n25544_), .A3(new_n25545_), .Z(new_n25546_));
  OAI21_X1   g22448(.A1(new_n25546_), .A2(pi0223), .B(new_n2587_), .ZN(new_n25547_));
  OAI21_X1   g22449(.A1(new_n25547_), .A2(new_n25542_), .B(pi0039), .ZN(new_n25548_));
  OAI22_X1   g22450(.A1(new_n25540_), .A2(new_n25548_), .B1(new_n25512_), .B2(new_n25516_), .ZN(new_n25549_));
  AOI22_X1   g22451(.A1(new_n25549_), .A2(new_n3172_), .B1(new_n25506_), .B2(new_n25507_), .ZN(new_n25550_));
  MUX2_X1    g22452(.I0(new_n25550_), .I1(pi0223), .S(new_n3232_), .Z(new_n25551_));
  NOR2_X1    g22453(.A1(new_n25551_), .A2(pi0778), .ZN(new_n25552_));
  NAND3_X1   g22454(.A1(new_n25551_), .A2(new_n12970_), .A3(new_n25385_), .ZN(new_n25553_));
  OAI21_X1   g22455(.A1(new_n25551_), .A2(pi0625), .B(new_n25384_), .ZN(new_n25554_));
  NAND3_X1   g22456(.A1(new_n25554_), .A2(new_n25553_), .A3(new_n11893_), .ZN(new_n25555_));
  NAND2_X1   g22457(.A1(new_n25555_), .A2(pi0778), .ZN(new_n25556_));
  XNOR2_X1   g22458(.A1(new_n25556_), .A2(new_n25552_), .ZN(new_n25557_));
  AOI21_X1   g22459(.A1(new_n25557_), .A2(new_n11938_), .B(new_n25505_), .ZN(new_n25558_));
  AOI21_X1   g22460(.A1(new_n25558_), .A2(new_n11961_), .B(new_n25504_), .ZN(new_n25559_));
  NAND2_X1   g22461(.A1(new_n25559_), .A2(new_n12032_), .ZN(new_n25560_));
  NAND2_X1   g22462(.A1(new_n25385_), .A2(new_n13713_), .ZN(new_n25561_));
  XOR2_X1    g22463(.A1(new_n25560_), .A2(new_n25561_), .Z(new_n25562_));
  AOI21_X1   g22464(.A1(new_n25562_), .A2(new_n12067_), .B(new_n25503_), .ZN(new_n25563_));
  INV_X1     g22465(.I(new_n25563_), .ZN(new_n25564_));
  MUX2_X1    g22466(.I0(new_n25564_), .I1(new_n25384_), .S(pi0647), .Z(new_n25565_));
  NOR2_X1    g22467(.A1(new_n25565_), .A2(pi1157), .ZN(new_n25566_));
  NOR2_X1    g22468(.A1(new_n25566_), .A2(new_n12060_), .ZN(new_n25567_));
  MUX2_X1    g22469(.I0(new_n25564_), .I1(new_n25384_), .S(new_n12061_), .Z(new_n25568_));
  NOR2_X1    g22470(.A1(new_n25568_), .A2(new_n12049_), .ZN(new_n25569_));
  NOR2_X1    g22471(.A1(new_n25569_), .A2(pi0630), .ZN(new_n25570_));
  OAI21_X1   g22472(.A1(new_n25567_), .A2(new_n25570_), .B(new_n12048_), .ZN(new_n25571_));
  AOI21_X1   g22473(.A1(new_n25502_), .A2(new_n15076_), .B(new_n25571_), .ZN(new_n25572_));
  MUX2_X1    g22474(.I0(new_n25500_), .I1(new_n25385_), .S(pi0626), .Z(new_n25573_));
  NOR2_X1    g22475(.A1(new_n25573_), .A2(new_n17171_), .ZN(new_n25574_));
  AND2_X2    g22476(.A1(new_n25500_), .A2(pi0626), .Z(new_n25575_));
  NOR2_X1    g22477(.A1(new_n11988_), .A2(new_n11994_), .ZN(new_n25576_));
  NAND2_X1   g22478(.A1(new_n25384_), .A2(new_n25576_), .ZN(new_n25577_));
  MUX2_X1    g22479(.I0(new_n25559_), .I1(new_n25385_), .S(new_n12013_), .Z(new_n25578_));
  OAI22_X1   g22480(.A1(new_n25575_), .A2(new_n25577_), .B1(new_n12020_), .B2(new_n25578_), .ZN(new_n25579_));
  OAI21_X1   g22481(.A1(new_n25579_), .A2(new_n25574_), .B(pi0788), .ZN(new_n25580_));
  INV_X1     g22482(.I(new_n25562_), .ZN(new_n25581_));
  NAND2_X1   g22483(.A1(new_n23402_), .A2(pi0628), .ZN(new_n25582_));
  NOR2_X1    g22484(.A1(new_n25581_), .A2(pi0628), .ZN(new_n25583_));
  OAI21_X1   g22485(.A1(new_n25385_), .A2(new_n12031_), .B(new_n12051_), .ZN(new_n25584_));
  OAI22_X1   g22486(.A1(new_n25583_), .A2(new_n25584_), .B1(new_n25581_), .B2(new_n25582_), .ZN(new_n25585_));
  OAI21_X1   g22487(.A1(new_n25501_), .A2(new_n17303_), .B(new_n25585_), .ZN(new_n25586_));
  INV_X1     g22488(.I(new_n25482_), .ZN(new_n25587_));
  NAND2_X1   g22489(.A1(new_n12109_), .A2(new_n12225_), .ZN(new_n25588_));
  NAND2_X1   g22490(.A1(new_n12112_), .A2(new_n12384_), .ZN(new_n25589_));
  NAND2_X1   g22491(.A1(new_n25588_), .A2(new_n25589_), .ZN(new_n25590_));
  MUX2_X1    g22492(.I0(new_n25590_), .I1(new_n25424_), .S(new_n25513_), .Z(new_n25591_));
  INV_X1     g22493(.I(new_n25591_), .ZN(new_n25592_));
  MUX2_X1    g22494(.I0(new_n12320_), .I1(new_n12112_), .S(pi0642), .Z(new_n25593_));
  NOR2_X1    g22495(.A1(new_n12109_), .A2(new_n25593_), .ZN(new_n25594_));
  OR4_X2     g22496(.A1(pi0223), .A2(new_n25395_), .A3(new_n25513_), .A4(new_n25594_), .Z(new_n25595_));
  NAND4_X1   g22497(.A1(new_n25592_), .A2(new_n25392_), .A3(new_n25393_), .A4(new_n25595_), .ZN(new_n25596_));
  OAI21_X1   g22498(.A1(new_n12164_), .A2(new_n12384_), .B(pi0680), .ZN(new_n25597_));
  NOR2_X1    g22499(.A1(new_n5104_), .A2(pi0642), .ZN(new_n25598_));
  NAND3_X1   g22500(.A1(new_n12489_), .A2(new_n12162_), .A3(new_n25598_), .ZN(new_n25599_));
  NOR2_X1    g22501(.A1(new_n12487_), .A2(new_n12187_), .ZN(new_n25600_));
  NAND3_X1   g22502(.A1(new_n25600_), .A2(new_n25597_), .A3(new_n25599_), .ZN(new_n25601_));
  OR2_X2     g22503(.A1(new_n25429_), .A2(new_n25508_), .Z(new_n25602_));
  AOI21_X1   g22504(.A1(new_n25601_), .A2(new_n25602_), .B(new_n25428_), .ZN(new_n25603_));
  NAND2_X1   g22505(.A1(new_n25399_), .A2(new_n5095_), .ZN(new_n25604_));
  NOR2_X1    g22506(.A1(new_n12331_), .A2(new_n12384_), .ZN(new_n25605_));
  INV_X1     g22507(.I(new_n25605_), .ZN(new_n25606_));
  NAND2_X1   g22508(.A1(new_n25606_), .A2(new_n12112_), .ZN(new_n25607_));
  NOR2_X1    g22509(.A1(new_n24795_), .A2(pi0680), .ZN(new_n25608_));
  OAI21_X1   g22510(.A1(new_n12226_), .A2(new_n12384_), .B(new_n5104_), .ZN(new_n25609_));
  AOI21_X1   g22511(.A1(new_n25607_), .A2(new_n25608_), .B(new_n25609_), .ZN(new_n25610_));
  OAI21_X1   g22512(.A1(new_n12220_), .A2(pi0642), .B(new_n25610_), .ZN(new_n25611_));
  AOI21_X1   g22513(.A1(new_n25611_), .A2(new_n25604_), .B(new_n12731_), .ZN(new_n25612_));
  NOR2_X1    g22514(.A1(new_n25421_), .A2(new_n25612_), .ZN(new_n25613_));
  MUX2_X1    g22515(.I0(new_n25613_), .I1(new_n25603_), .S(new_n6445_), .Z(new_n25614_));
  OAI21_X1   g22516(.A1(new_n25413_), .A2(new_n12731_), .B(new_n25513_), .ZN(new_n25615_));
  NAND2_X1   g22517(.A1(new_n25218_), .A2(new_n12187_), .ZN(new_n25616_));
  NAND3_X1   g22518(.A1(new_n25063_), .A2(new_n25215_), .A3(new_n25598_), .ZN(new_n25617_));
  NOR2_X1    g22519(.A1(pi0642), .A2(pi0680), .ZN(new_n25618_));
  NAND4_X1   g22520(.A1(new_n25616_), .A2(new_n25223_), .A3(new_n25617_), .A4(new_n25618_), .ZN(new_n25619_));
  NAND3_X1   g22521(.A1(new_n25415_), .A2(new_n25615_), .A3(new_n25619_), .ZN(new_n25620_));
  OAI21_X1   g22522(.A1(new_n24792_), .A2(new_n12111_), .B(new_n12384_), .ZN(new_n25621_));
  NAND2_X1   g22523(.A1(new_n25621_), .A2(new_n25606_), .ZN(new_n25622_));
  NOR2_X1    g22524(.A1(new_n5105_), .A2(pi0680), .ZN(new_n25623_));
  AOI22_X1   g22525(.A1(new_n25405_), .A2(new_n25513_), .B1(new_n25622_), .B2(new_n25623_), .ZN(new_n25624_));
  NAND2_X1   g22526(.A1(new_n25409_), .A2(new_n25624_), .ZN(new_n25625_));
  AOI21_X1   g22527(.A1(new_n25625_), .A2(new_n25620_), .B(pi0223), .ZN(new_n25626_));
  OAI22_X1   g22528(.A1(new_n25626_), .A2(new_n3284_), .B1(pi0223), .B2(new_n25614_), .ZN(new_n25627_));
  NAND2_X1   g22529(.A1(new_n13829_), .A2(new_n25521_), .ZN(new_n25628_));
  NAND3_X1   g22530(.A1(new_n25310_), .A2(pi0223), .A3(new_n25469_), .ZN(new_n25629_));
  NOR2_X1    g22531(.A1(new_n25471_), .A2(new_n25508_), .ZN(new_n25630_));
  NAND4_X1   g22532(.A1(new_n25628_), .A2(new_n13358_), .A3(new_n25629_), .A4(new_n25630_), .ZN(new_n25631_));
  NAND4_X1   g22533(.A1(new_n25475_), .A2(new_n13355_), .A3(new_n25315_), .A4(new_n25513_), .ZN(new_n25632_));
  NOR3_X1    g22534(.A1(new_n25474_), .A2(pi0223), .A3(new_n12731_), .ZN(new_n25633_));
  NAND3_X1   g22535(.A1(new_n25632_), .A2(new_n13844_), .A3(new_n25633_), .ZN(new_n25634_));
  NAND3_X1   g22536(.A1(new_n25631_), .A2(new_n25634_), .A3(new_n3154_), .ZN(new_n25635_));
  NAND2_X1   g22537(.A1(new_n25635_), .A2(new_n3172_), .ZN(new_n25636_));
  INV_X1     g22538(.I(new_n25451_), .ZN(new_n25637_));
  NAND3_X1   g22539(.A1(new_n25285_), .A2(pi0642), .A3(new_n5095_), .ZN(new_n25638_));
  AOI21_X1   g22540(.A1(new_n12465_), .A2(new_n25598_), .B(new_n25638_), .ZN(new_n25639_));
  INV_X1     g22541(.I(new_n12258_), .ZN(new_n25640_));
  OAI21_X1   g22542(.A1(new_n12467_), .A2(new_n25640_), .B(new_n12187_), .ZN(new_n25641_));
  NOR4_X1    g22543(.A1(new_n25288_), .A2(new_n12384_), .A3(pi0680), .A4(pi0681), .ZN(new_n25642_));
  NOR2_X1    g22544(.A1(new_n25642_), .A2(new_n5094_), .ZN(new_n25643_));
  OAI21_X1   g22545(.A1(new_n25639_), .A2(new_n25641_), .B(new_n25643_), .ZN(new_n25644_));
  INV_X1     g22546(.I(new_n25455_), .ZN(new_n25645_));
  NAND2_X1   g22547(.A1(new_n12468_), .A2(new_n25610_), .ZN(new_n25646_));
  NAND4_X1   g22548(.A1(new_n25645_), .A2(new_n25521_), .A3(new_n25604_), .A4(new_n25646_), .ZN(new_n25647_));
  AOI21_X1   g22549(.A1(new_n25644_), .A2(new_n25637_), .B(new_n25647_), .ZN(new_n25648_));
  INV_X1     g22550(.I(new_n25438_), .ZN(new_n25649_));
  NOR2_X1    g22551(.A1(new_n12355_), .A2(new_n5095_), .ZN(new_n25650_));
  INV_X1     g22552(.I(new_n25650_), .ZN(new_n25651_));
  NAND4_X1   g22553(.A1(new_n25288_), .A2(new_n5105_), .A3(new_n12302_), .A4(new_n12304_), .ZN(new_n25652_));
  NAND4_X1   g22554(.A1(new_n25651_), .A2(new_n12384_), .A3(new_n25267_), .A4(new_n25652_), .ZN(new_n25653_));
  NAND4_X1   g22555(.A1(new_n25653_), .A2(new_n5095_), .A3(new_n12731_), .A4(new_n25649_), .ZN(new_n25654_));
  NAND4_X1   g22556(.A1(new_n25649_), .A2(new_n12731_), .A3(new_n5099_), .A4(new_n25439_), .ZN(new_n25655_));
  NAND2_X1   g22557(.A1(new_n25654_), .A2(new_n25655_), .ZN(new_n25656_));
  NOR2_X1    g22558(.A1(new_n5098_), .A2(new_n12731_), .ZN(new_n25657_));
  NAND2_X1   g22559(.A1(new_n25445_), .A2(new_n5095_), .ZN(new_n25658_));
  INV_X1     g22560(.I(new_n12340_), .ZN(new_n25659_));
  NAND2_X1   g22561(.A1(new_n25659_), .A2(new_n25594_), .ZN(new_n25660_));
  AOI21_X1   g22562(.A1(new_n25660_), .A2(new_n5105_), .B(new_n5095_), .ZN(new_n25661_));
  INV_X1     g22563(.I(new_n12381_), .ZN(new_n25662_));
  NOR4_X1    g22564(.A1(new_n25662_), .A2(new_n12382_), .A3(pi0614), .A4(new_n12354_), .ZN(new_n25663_));
  OAI21_X1   g22565(.A1(new_n25663_), .A2(new_n25605_), .B(new_n12166_), .ZN(new_n25664_));
  AOI21_X1   g22566(.A1(new_n25664_), .A2(new_n25661_), .B(new_n12731_), .ZN(new_n25665_));
  AOI22_X1   g22567(.A1(new_n25658_), .A2(new_n25665_), .B1(new_n25445_), .B2(new_n25657_), .ZN(new_n25666_));
  MUX2_X1    g22568(.I0(new_n25666_), .I1(new_n25656_), .S(new_n6445_), .Z(new_n25667_));
  AOI21_X1   g22569(.A1(new_n25667_), .A2(pi0223), .B(new_n25648_), .ZN(new_n25668_));
  NOR2_X1    g22570(.A1(new_n25656_), .A2(new_n5141_), .ZN(new_n25669_));
  NOR2_X1    g22571(.A1(new_n25669_), .A2(pi0223), .ZN(new_n25670_));
  OAI21_X1   g22572(.A1(new_n6460_), .A2(new_n25666_), .B(new_n25670_), .ZN(new_n25671_));
  NOR2_X1    g22573(.A1(new_n25592_), .A2(new_n12133_), .ZN(new_n25672_));
  NOR3_X1    g22574(.A1(new_n25672_), .A2(new_n2614_), .A3(new_n3294_), .ZN(new_n25673_));
  OAI21_X1   g22575(.A1(new_n25613_), .A2(new_n6460_), .B(new_n25673_), .ZN(new_n25674_));
  AOI21_X1   g22576(.A1(new_n25603_), .A2(new_n5141_), .B(new_n25674_), .ZN(new_n25675_));
  AOI21_X1   g22577(.A1(new_n25671_), .A2(new_n25675_), .B(new_n3154_), .ZN(new_n25676_));
  NAND4_X1   g22578(.A1(new_n25672_), .A2(new_n2604_), .A3(new_n25517_), .A4(new_n25595_), .ZN(new_n25677_));
  NAND2_X1   g22579(.A1(new_n25677_), .A2(new_n4905_), .ZN(new_n25678_));
  NOR3_X1    g22580(.A1(new_n25676_), .A2(new_n25668_), .A3(new_n25678_), .ZN(new_n25679_));
  NAND3_X1   g22581(.A1(new_n25636_), .A2(new_n25627_), .A3(new_n25679_), .ZN(new_n25680_));
  AOI21_X1   g22582(.A1(new_n25680_), .A2(new_n25596_), .B(new_n3232_), .ZN(new_n25681_));
  XOR2_X1    g22583(.A1(new_n25681_), .A2(new_n25390_), .Z(new_n25682_));
  OAI21_X1   g22584(.A1(new_n25682_), .A2(pi0625), .B(new_n25587_), .ZN(new_n25683_));
  NAND3_X1   g22585(.A1(new_n25682_), .A2(new_n12970_), .A3(new_n25482_), .ZN(new_n25684_));
  NAND3_X1   g22586(.A1(new_n25683_), .A2(new_n25684_), .A3(new_n12977_), .ZN(new_n25685_));
  NOR4_X1    g22587(.A1(new_n25587_), .A2(new_n12970_), .A3(new_n25682_), .A4(pi1153), .ZN(new_n25686_));
  OAI21_X1   g22588(.A1(new_n25686_), .A2(new_n25555_), .B(new_n13657_), .ZN(new_n25687_));
  NAND2_X1   g22589(.A1(new_n25685_), .A2(new_n25687_), .ZN(new_n25688_));
  NOR2_X1    g22590(.A1(new_n25682_), .A2(pi0778), .ZN(new_n25689_));
  AOI21_X1   g22591(.A1(new_n25688_), .A2(pi0778), .B(new_n25689_), .ZN(new_n25690_));
  NOR2_X1    g22592(.A1(new_n25690_), .A2(pi0785), .ZN(new_n25691_));
  NOR3_X1    g22593(.A1(new_n25557_), .A2(new_n11903_), .A3(new_n11912_), .ZN(new_n25692_));
  OAI21_X1   g22594(.A1(new_n25486_), .A2(new_n11912_), .B(new_n11923_), .ZN(new_n25693_));
  INV_X1     g22595(.I(new_n25557_), .ZN(new_n25694_));
  NOR4_X1    g22596(.A1(new_n25690_), .A2(new_n11903_), .A3(pi1155), .A4(new_n25694_), .ZN(new_n25695_));
  NOR2_X1    g22597(.A1(new_n25695_), .A2(new_n25485_), .ZN(new_n25696_));
  OAI22_X1   g22598(.A1(new_n25696_), .A2(pi0660), .B1(new_n25692_), .B2(new_n25693_), .ZN(new_n25697_));
  AOI21_X1   g22599(.A1(new_n25697_), .A2(pi0785), .B(new_n25691_), .ZN(new_n25698_));
  NAND2_X1   g22600(.A1(new_n25698_), .A2(new_n11969_), .ZN(new_n25699_));
  NOR2_X1    g22601(.A1(new_n11934_), .A2(pi1154), .ZN(new_n25700_));
  NAND2_X1   g22602(.A1(new_n25698_), .A2(new_n25700_), .ZN(new_n25701_));
  AOI21_X1   g22603(.A1(pi0627), .A2(new_n25493_), .B(new_n25701_), .ZN(new_n25702_));
  NAND2_X1   g22604(.A1(new_n25558_), .A2(pi0618), .ZN(new_n25703_));
  NAND2_X1   g22605(.A1(new_n25703_), .A2(new_n11960_), .ZN(new_n25704_));
  AOI21_X1   g22606(.A1(new_n25698_), .A2(new_n11934_), .B(new_n25704_), .ZN(new_n25705_));
  OAI21_X1   g22607(.A1(new_n25702_), .A2(new_n25705_), .B(pi0781), .ZN(new_n25706_));
  XOR2_X1    g22608(.A1(new_n25706_), .A2(new_n25699_), .Z(new_n25707_));
  NAND2_X1   g22609(.A1(new_n25707_), .A2(pi0619), .ZN(new_n25708_));
  AND2_X2    g22610(.A1(new_n25559_), .A2(new_n14638_), .Z(new_n25709_));
  AOI21_X1   g22611(.A1(new_n25708_), .A2(new_n25709_), .B(new_n25499_), .ZN(new_n25710_));
  NOR3_X1    g22612(.A1(new_n25559_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n25711_));
  OAI21_X1   g22613(.A1(new_n25707_), .A2(pi0789), .B(new_n11998_), .ZN(new_n25712_));
  NAND4_X1   g22614(.A1(new_n25712_), .A2(new_n11966_), .A3(new_n11985_), .A4(new_n25711_), .ZN(new_n25713_));
  NOR2_X1    g22615(.A1(new_n25713_), .A2(new_n25710_), .ZN(new_n25714_));
  AOI21_X1   g22616(.A1(new_n25586_), .A2(pi0792), .B(new_n25714_), .ZN(new_n25715_));
  OAI21_X1   g22617(.A1(new_n25586_), .A2(new_n14732_), .B(new_n14726_), .ZN(new_n25716_));
  AOI21_X1   g22618(.A1(new_n25580_), .A2(new_n25715_), .B(new_n25716_), .ZN(new_n25717_));
  NOR2_X1    g22619(.A1(new_n25717_), .A2(new_n25572_), .ZN(new_n25718_));
  NAND2_X1   g22620(.A1(new_n25502_), .A2(new_n12092_), .ZN(new_n25719_));
  AOI21_X1   g22621(.A1(new_n25385_), .A2(new_n12091_), .B(new_n12082_), .ZN(new_n25720_));
  NAND2_X1   g22622(.A1(new_n25719_), .A2(new_n25720_), .ZN(new_n25721_));
  OAI21_X1   g22623(.A1(new_n12082_), .A2(new_n25384_), .B(new_n25721_), .ZN(new_n25722_));
  AOI21_X1   g22624(.A1(new_n25722_), .A2(pi0715), .B(pi1160), .ZN(new_n25723_));
  NOR4_X1    g22625(.A1(new_n25723_), .A2(pi0644), .A3(new_n12099_), .A4(new_n25718_), .ZN(new_n25726_));
  AOI21_X1   g22626(.A1(new_n25384_), .A2(new_n12082_), .B(pi0715), .ZN(new_n25727_));
  AOI21_X1   g22627(.A1(new_n25721_), .A2(new_n25727_), .B(new_n12081_), .ZN(new_n25728_));
  NAND2_X1   g22628(.A1(new_n12099_), .A2(pi0644), .ZN(new_n25729_));
  NOR3_X1    g22629(.A1(new_n25718_), .A2(new_n25728_), .A3(new_n25729_), .ZN(new_n25730_));
  NOR2_X1    g22630(.A1(new_n25726_), .A2(new_n25730_), .ZN(new_n25731_));
  MUX2_X1    g22631(.I0(new_n25731_), .I1(new_n25718_), .S(new_n11867_), .Z(new_n25732_));
  NAND2_X1   g22632(.A1(po1038), .A2(pi0223), .ZN(new_n25733_));
  OAI21_X1   g22633(.A1(new_n25732_), .A2(po1038), .B(new_n25733_), .ZN(po0380));
  NAND2_X1   g22634(.A1(new_n25018_), .A2(pi0224), .ZN(new_n25735_));
  INV_X1     g22635(.I(new_n25735_), .ZN(new_n25736_));
  NOR2_X1    g22636(.A1(new_n25736_), .A2(new_n12054_), .ZN(new_n25737_));
  NOR2_X1    g22637(.A1(new_n25735_), .A2(new_n14624_), .ZN(new_n25738_));
  NOR2_X1    g22638(.A1(new_n3231_), .A2(pi0224), .ZN(new_n25739_));
  NOR2_X1    g22639(.A1(new_n11875_), .A2(new_n12443_), .ZN(new_n25740_));
  INV_X1     g22640(.I(new_n25740_), .ZN(new_n25741_));
  AOI21_X1   g22641(.A1(new_n25741_), .A2(new_n12132_), .B(new_n5106_), .ZN(new_n25742_));
  AOI21_X1   g22642(.A1(new_n24957_), .A2(new_n12166_), .B(new_n25742_), .ZN(new_n25743_));
  NAND2_X1   g22643(.A1(new_n25743_), .A2(new_n12461_), .ZN(new_n25744_));
  INV_X1     g22644(.I(new_n25743_), .ZN(new_n25745_));
  NOR2_X1    g22645(.A1(new_n12231_), .A2(new_n25740_), .ZN(new_n25746_));
  INV_X1     g22646(.I(new_n25746_), .ZN(new_n25747_));
  MUX2_X1    g22647(.I0(new_n25747_), .I1(new_n25745_), .S(new_n5095_), .Z(new_n25748_));
  OAI21_X1   g22648(.A1(new_n25748_), .A2(new_n12461_), .B(new_n25744_), .ZN(new_n25749_));
  AOI21_X1   g22649(.A1(new_n12158_), .A2(pi0616), .B(pi0614), .ZN(new_n25750_));
  AOI21_X1   g22650(.A1(new_n12489_), .A2(pi0614), .B(new_n25750_), .ZN(new_n25751_));
  NAND3_X1   g22651(.A1(new_n12489_), .A2(new_n25750_), .A3(pi0614), .ZN(new_n25752_));
  AOI21_X1   g22652(.A1(new_n12156_), .A2(new_n5104_), .B(new_n5108_), .ZN(new_n25753_));
  NAND2_X1   g22653(.A1(new_n25752_), .A2(new_n25753_), .ZN(new_n25754_));
  NOR3_X1    g22654(.A1(new_n25754_), .A2(new_n12411_), .A3(new_n25751_), .ZN(new_n25755_));
  AOI21_X1   g22655(.A1(new_n12425_), .A2(pi0614), .B(new_n5095_), .ZN(new_n25756_));
  INV_X1     g22656(.I(new_n25756_), .ZN(new_n25757_));
  OAI22_X1   g22657(.A1(new_n25757_), .A2(new_n12156_), .B1(new_n5095_), .B2(new_n25741_), .ZN(new_n25758_));
  NAND2_X1   g22658(.A1(new_n25758_), .A2(new_n12461_), .ZN(new_n25759_));
  INV_X1     g22659(.I(new_n25759_), .ZN(new_n25760_));
  OAI21_X1   g22660(.A1(new_n25755_), .A2(pi0680), .B(new_n25760_), .ZN(new_n25761_));
  OAI21_X1   g22661(.A1(new_n12129_), .A2(new_n25755_), .B(new_n25761_), .ZN(new_n25762_));
  AOI21_X1   g22662(.A1(new_n25762_), .A2(new_n6445_), .B(pi0224), .ZN(new_n25763_));
  OAI21_X1   g22663(.A1(new_n25749_), .A2(new_n6445_), .B(new_n25763_), .ZN(new_n25764_));
  NAND2_X1   g22664(.A1(new_n12157_), .A2(new_n25740_), .ZN(new_n25765_));
  NAND2_X1   g22665(.A1(new_n25765_), .A2(new_n5095_), .ZN(new_n25766_));
  AOI21_X1   g22666(.A1(new_n25766_), .A2(new_n25757_), .B(new_n12461_), .ZN(new_n25767_));
  AOI21_X1   g22667(.A1(new_n12461_), .A2(new_n25765_), .B(new_n25767_), .ZN(new_n25768_));
  NAND2_X1   g22668(.A1(new_n25061_), .A2(pi0614), .ZN(new_n25769_));
  INV_X1     g22669(.I(new_n25769_), .ZN(new_n25770_));
  MUX2_X1    g22670(.I0(new_n25770_), .I1(new_n25768_), .S(new_n6445_), .Z(new_n25771_));
  AOI21_X1   g22671(.A1(new_n25771_), .A2(new_n2595_), .B(new_n3284_), .ZN(new_n25772_));
  AOI21_X1   g22672(.A1(new_n12133_), .A2(pi0224), .B(new_n3285_), .ZN(new_n25773_));
  NOR2_X1    g22673(.A1(new_n12209_), .A2(new_n12443_), .ZN(new_n25774_));
  INV_X1     g22674(.I(new_n25774_), .ZN(new_n25775_));
  NAND2_X1   g22675(.A1(new_n25775_), .A2(new_n25773_), .ZN(new_n25776_));
  NAND2_X1   g22676(.A1(new_n25776_), .A2(new_n2566_), .ZN(new_n25777_));
  AOI21_X1   g22677(.A1(new_n25764_), .A2(new_n25772_), .B(new_n25777_), .ZN(new_n25778_));
  OR2_X2     g22678(.A1(new_n25749_), .A2(new_n6460_), .Z(new_n25779_));
  AOI21_X1   g22679(.A1(new_n25762_), .A2(new_n6460_), .B(pi0224), .ZN(new_n25780_));
  NOR2_X1    g22680(.A1(new_n25025_), .A2(new_n25742_), .ZN(new_n25781_));
  INV_X1     g22681(.I(new_n25781_), .ZN(new_n25782_));
  NOR2_X1    g22682(.A1(new_n12725_), .A2(new_n25740_), .ZN(new_n25783_));
  MUX2_X1    g22683(.I0(new_n25783_), .I1(new_n25781_), .S(new_n5095_), .Z(new_n25784_));
  NAND2_X1   g22684(.A1(new_n25784_), .A2(new_n12129_), .ZN(new_n25785_));
  OAI21_X1   g22685(.A1(new_n12129_), .A2(new_n25782_), .B(new_n25785_), .ZN(new_n25786_));
  NOR2_X1    g22686(.A1(new_n25786_), .A2(new_n6460_), .ZN(new_n25787_));
  NAND2_X1   g22687(.A1(new_n12310_), .A2(pi0614), .ZN(new_n25788_));
  AND2_X2    g22688(.A1(new_n24857_), .A2(new_n25788_), .Z(new_n25789_));
  INV_X1     g22689(.I(new_n25789_), .ZN(new_n25790_));
  NOR2_X1    g22690(.A1(new_n25789_), .A2(pi0680), .ZN(new_n25791_));
  AOI21_X1   g22691(.A1(pi0614), .A2(new_n12308_), .B(new_n12262_), .ZN(new_n25792_));
  OAI21_X1   g22692(.A1(new_n25792_), .A2(new_n5095_), .B(new_n12461_), .ZN(new_n25793_));
  NOR2_X1    g22693(.A1(new_n25791_), .A2(new_n25793_), .ZN(new_n25794_));
  AOI21_X1   g22694(.A1(new_n12461_), .A2(new_n25790_), .B(new_n25794_), .ZN(new_n25795_));
  OAI21_X1   g22695(.A1(new_n25795_), .A2(new_n5141_), .B(new_n2595_), .ZN(new_n25796_));
  NOR2_X1    g22696(.A1(new_n25042_), .A2(new_n25775_), .ZN(new_n25797_));
  NAND2_X1   g22697(.A1(new_n25797_), .A2(new_n2595_), .ZN(new_n25798_));
  NOR3_X1    g22698(.A1(new_n25798_), .A2(pi0223), .A3(new_n12685_), .ZN(new_n25799_));
  OAI21_X1   g22699(.A1(new_n25796_), .A2(new_n25787_), .B(new_n25799_), .ZN(new_n25800_));
  AOI21_X1   g22700(.A1(new_n25769_), .A2(new_n25768_), .B(new_n6460_), .ZN(new_n25801_));
  NAND2_X1   g22701(.A1(new_n25801_), .A2(new_n4878_), .ZN(new_n25802_));
  NAND2_X1   g22702(.A1(new_n12506_), .A2(pi0614), .ZN(new_n25803_));
  NAND4_X1   g22703(.A1(new_n25800_), .A2(new_n2604_), .A3(new_n25802_), .A4(new_n25803_), .ZN(new_n25804_));
  AOI21_X1   g22704(.A1(new_n25779_), .A2(new_n25780_), .B(new_n25804_), .ZN(new_n25805_));
  NOR2_X1    g22705(.A1(new_n25786_), .A2(new_n6445_), .ZN(new_n25806_));
  OAI21_X1   g22706(.A1(new_n25795_), .A2(new_n5094_), .B(new_n2595_), .ZN(new_n25807_));
  NOR2_X1    g22707(.A1(new_n25807_), .A2(new_n25806_), .ZN(new_n25808_));
  AOI21_X1   g22708(.A1(new_n12676_), .A2(new_n25798_), .B(new_n25808_), .ZN(new_n25809_));
  NOR2_X1    g22709(.A1(new_n25809_), .A2(new_n24682_), .ZN(new_n25810_));
  OAI21_X1   g22710(.A1(new_n25805_), .A2(new_n6594_), .B(new_n25810_), .ZN(new_n25811_));
  NAND2_X1   g22711(.A1(new_n13831_), .A2(pi0614), .ZN(new_n25812_));
  INV_X1     g22712(.I(new_n25812_), .ZN(new_n25813_));
  NAND2_X1   g22713(.A1(new_n12627_), .A2(pi0224), .ZN(new_n25814_));
  OAI22_X1   g22714(.A1(new_n25813_), .A2(new_n25814_), .B1(new_n2595_), .B2(new_n12590_), .ZN(new_n25815_));
  OAI21_X1   g22715(.A1(new_n13858_), .A2(pi0614), .B(pi0224), .ZN(new_n25816_));
  NOR2_X1    g22716(.A1(new_n25816_), .A2(new_n13859_), .ZN(new_n25817_));
  NAND2_X1   g22717(.A1(new_n12610_), .A2(pi0614), .ZN(new_n25818_));
  OAI21_X1   g22718(.A1(new_n25818_), .A2(pi0224), .B(new_n2587_), .ZN(new_n25819_));
  NOR2_X1    g22719(.A1(pi0038), .A2(pi0039), .ZN(new_n25821_));
  OAI21_X1   g22720(.A1(new_n25817_), .A2(new_n25819_), .B(new_n25821_), .ZN(new_n25822_));
  AOI21_X1   g22721(.A1(pi0299), .A2(new_n25815_), .B(new_n25822_), .ZN(new_n25823_));
  OAI21_X1   g22722(.A1(new_n25811_), .A2(new_n25778_), .B(new_n25823_), .ZN(new_n25824_));
  NAND2_X1   g22723(.A1(new_n25824_), .A2(new_n3231_), .ZN(new_n25825_));
  XOR2_X1    g22724(.A1(new_n25825_), .A2(new_n25739_), .Z(new_n25826_));
  NAND2_X1   g22725(.A1(new_n25826_), .A2(new_n11924_), .ZN(new_n25827_));
  NAND2_X1   g22726(.A1(new_n25735_), .A2(new_n11914_), .ZN(new_n25828_));
  NAND2_X1   g22727(.A1(new_n25827_), .A2(new_n25828_), .ZN(new_n25829_));
  INV_X1     g22728(.I(new_n25829_), .ZN(new_n25830_));
  NAND3_X1   g22729(.A1(new_n25829_), .A2(new_n11903_), .A3(new_n25736_), .ZN(new_n25831_));
  OAI21_X1   g22730(.A1(new_n25829_), .A2(pi0609), .B(new_n25735_), .ZN(new_n25832_));
  NAND3_X1   g22731(.A1(new_n25832_), .A2(new_n25831_), .A3(new_n11912_), .ZN(new_n25833_));
  MUX2_X1    g22732(.I0(new_n25833_), .I1(new_n25830_), .S(new_n11870_), .Z(new_n25834_));
  NAND2_X1   g22733(.A1(new_n25834_), .A2(new_n11969_), .ZN(new_n25835_));
  NOR3_X1    g22734(.A1(new_n25834_), .A2(pi0618), .A3(new_n25735_), .ZN(new_n25836_));
  AOI21_X1   g22735(.A1(new_n25834_), .A2(new_n11934_), .B(new_n25736_), .ZN(new_n25837_));
  NOR3_X1    g22736(.A1(new_n25836_), .A2(new_n25837_), .A3(pi1154), .ZN(new_n25838_));
  NOR2_X1    g22737(.A1(new_n25838_), .A2(new_n11969_), .ZN(new_n25839_));
  XNOR2_X1   g22738(.A1(new_n25839_), .A2(new_n25835_), .ZN(new_n25840_));
  INV_X1     g22739(.I(new_n25840_), .ZN(new_n25841_));
  NAND3_X1   g22740(.A1(new_n25841_), .A2(new_n11967_), .A3(new_n25736_), .ZN(new_n25842_));
  OAI21_X1   g22741(.A1(new_n25841_), .A2(pi0619), .B(new_n25735_), .ZN(new_n25843_));
  NAND3_X1   g22742(.A1(new_n25843_), .A2(new_n25842_), .A3(new_n11869_), .ZN(new_n25844_));
  MUX2_X1    g22743(.I0(new_n25844_), .I1(new_n25840_), .S(new_n11985_), .Z(new_n25845_));
  AOI21_X1   g22744(.A1(new_n25845_), .A2(new_n14624_), .B(new_n25738_), .ZN(new_n25846_));
  AOI21_X1   g22745(.A1(new_n25846_), .A2(new_n12054_), .B(new_n25737_), .ZN(new_n25847_));
  NAND2_X1   g22746(.A1(new_n25847_), .A2(new_n15076_), .ZN(new_n25848_));
  NOR2_X1    g22747(.A1(new_n25736_), .A2(new_n12067_), .ZN(new_n25849_));
  AOI21_X1   g22748(.A1(new_n13368_), .A2(pi0224), .B(new_n3172_), .ZN(new_n25850_));
  NAND2_X1   g22749(.A1(new_n13402_), .A2(pi0662), .ZN(new_n25851_));
  NOR2_X1    g22750(.A1(new_n24848_), .A2(new_n5095_), .ZN(new_n25852_));
  INV_X1     g22751(.I(new_n25852_), .ZN(new_n25853_));
  OAI21_X1   g22752(.A1(new_n12160_), .A2(new_n25853_), .B(new_n25773_), .ZN(new_n25854_));
  NAND2_X1   g22753(.A1(new_n25118_), .A2(pi0662), .ZN(new_n25855_));
  OAI21_X1   g22754(.A1(new_n12879_), .A2(pi0662), .B(new_n25855_), .ZN(new_n25856_));
  NOR2_X1    g22755(.A1(new_n25856_), .A2(new_n6445_), .ZN(new_n25857_));
  AOI21_X1   g22756(.A1(new_n25128_), .A2(new_n5097_), .B(new_n12767_), .ZN(new_n25858_));
  OAI21_X1   g22757(.A1(new_n25858_), .A2(new_n5094_), .B(new_n2595_), .ZN(new_n25859_));
  NAND2_X1   g22758(.A1(new_n12944_), .A2(new_n25852_), .ZN(new_n25860_));
  NAND2_X1   g22759(.A1(new_n25860_), .A2(new_n5094_), .ZN(new_n25861_));
  NOR2_X1    g22760(.A1(new_n25143_), .A2(new_n24848_), .ZN(new_n25862_));
  NOR2_X1    g22761(.A1(new_n25862_), .A2(new_n5094_), .ZN(new_n25863_));
  NOR2_X1    g22762(.A1(new_n25863_), .A2(pi0224), .ZN(new_n25864_));
  AOI21_X1   g22763(.A1(new_n25864_), .A2(new_n25861_), .B(new_n3284_), .ZN(new_n25865_));
  OAI21_X1   g22764(.A1(new_n25857_), .A2(new_n25859_), .B(new_n25865_), .ZN(new_n25866_));
  AOI21_X1   g22765(.A1(new_n25866_), .A2(new_n25854_), .B(pi0215), .ZN(new_n25867_));
  NOR2_X1    g22766(.A1(new_n25856_), .A2(new_n6460_), .ZN(new_n25868_));
  OAI21_X1   g22767(.A1(new_n25858_), .A2(new_n5141_), .B(new_n2595_), .ZN(new_n25869_));
  NOR2_X1    g22768(.A1(new_n25868_), .A2(new_n25869_), .ZN(new_n25870_));
  NOR2_X1    g22769(.A1(new_n12913_), .A2(new_n24848_), .ZN(new_n25871_));
  AOI21_X1   g22770(.A1(new_n12886_), .A2(new_n24848_), .B(new_n25871_), .ZN(new_n25872_));
  NOR2_X1    g22771(.A1(new_n25135_), .A2(new_n24848_), .ZN(new_n25873_));
  AOI21_X1   g22772(.A1(new_n24990_), .A2(new_n24848_), .B(new_n25873_), .ZN(new_n25874_));
  AND3_X2    g22773(.A1(new_n25874_), .A2(new_n2595_), .A3(new_n5141_), .Z(new_n25875_));
  NOR2_X1    g22774(.A1(pi0223), .A2(pi0224), .ZN(new_n25876_));
  NAND3_X1   g22775(.A1(new_n12939_), .A2(pi0662), .A3(new_n25876_), .ZN(new_n25877_));
  AOI21_X1   g22776(.A1(new_n25875_), .A2(new_n25872_), .B(new_n25877_), .ZN(new_n25878_));
  NAND3_X1   g22777(.A1(new_n12504_), .A2(pi0662), .A3(new_n11884_), .ZN(new_n25879_));
  NAND2_X1   g22778(.A1(new_n4878_), .A2(new_n3154_), .ZN(new_n25880_));
  AOI21_X1   g22779(.A1(new_n25879_), .A2(new_n2604_), .B(new_n25880_), .ZN(new_n25881_));
  OAI21_X1   g22780(.A1(new_n25862_), .A2(new_n5141_), .B(new_n25881_), .ZN(new_n25882_));
  AOI21_X1   g22781(.A1(new_n5141_), .A2(new_n25860_), .B(new_n25882_), .ZN(new_n25883_));
  OAI21_X1   g22782(.A1(new_n25878_), .A2(pi0299), .B(new_n25883_), .ZN(new_n25884_));
  NAND3_X1   g22783(.A1(new_n12951_), .A2(new_n2595_), .A3(pi0662), .ZN(new_n25885_));
  NAND4_X1   g22784(.A1(new_n25872_), .A2(new_n25874_), .A3(new_n2595_), .A4(new_n5094_), .ZN(new_n25886_));
  AOI21_X1   g22785(.A1(new_n25886_), .A2(new_n25885_), .B(new_n24682_), .ZN(new_n25887_));
  OAI21_X1   g22786(.A1(new_n25884_), .A2(new_n25870_), .B(new_n25887_), .ZN(new_n25888_));
  MUX2_X1    g22787(.I0(new_n25853_), .I1(new_n2595_), .S(new_n12624_), .Z(new_n25889_));
  OAI21_X1   g22788(.A1(new_n12648_), .A2(new_n2595_), .B(new_n2587_), .ZN(new_n25890_));
  MUX2_X1    g22789(.I0(new_n12641_), .I1(new_n12655_), .S(pi0224), .Z(new_n25891_));
  NAND2_X1   g22790(.A1(new_n12641_), .A2(new_n25853_), .ZN(new_n25892_));
  AOI21_X1   g22791(.A1(new_n25891_), .A2(pi0299), .B(new_n25892_), .ZN(new_n25893_));
  OAI22_X1   g22792(.A1(new_n25893_), .A2(pi0039), .B1(new_n25889_), .B2(new_n25890_), .ZN(new_n25894_));
  OAI21_X1   g22793(.A1(new_n25888_), .A2(new_n25867_), .B(new_n25894_), .ZN(new_n25895_));
  AOI22_X1   g22794(.A1(new_n25895_), .A2(new_n3172_), .B1(new_n25850_), .B2(new_n25851_), .ZN(new_n25896_));
  NOR2_X1    g22795(.A1(new_n25896_), .A2(new_n3232_), .ZN(new_n25897_));
  XOR2_X1    g22796(.A1(new_n25897_), .A2(new_n25739_), .Z(new_n25898_));
  INV_X1     g22797(.I(new_n25898_), .ZN(new_n25899_));
  NOR2_X1    g22798(.A1(new_n25899_), .A2(pi0778), .ZN(new_n25900_));
  NAND3_X1   g22799(.A1(new_n25899_), .A2(new_n12970_), .A3(new_n25736_), .ZN(new_n25901_));
  OAI21_X1   g22800(.A1(new_n25899_), .A2(pi0625), .B(new_n25735_), .ZN(new_n25902_));
  NAND3_X1   g22801(.A1(new_n25902_), .A2(new_n25901_), .A3(new_n11893_), .ZN(new_n25903_));
  NAND2_X1   g22802(.A1(new_n25903_), .A2(pi0778), .ZN(new_n25904_));
  XNOR2_X1   g22803(.A1(new_n25904_), .A2(new_n25900_), .ZN(new_n25905_));
  INV_X1     g22804(.I(new_n25905_), .ZN(new_n25906_));
  NOR2_X1    g22805(.A1(new_n25736_), .A2(new_n11938_), .ZN(new_n25907_));
  AOI21_X1   g22806(.A1(new_n25906_), .A2(new_n11938_), .B(new_n25907_), .ZN(new_n25908_));
  INV_X1     g22807(.I(new_n25908_), .ZN(new_n25909_));
  NOR2_X1    g22808(.A1(new_n25736_), .A2(new_n11961_), .ZN(new_n25910_));
  AOI21_X1   g22809(.A1(new_n25909_), .A2(new_n11961_), .B(new_n25910_), .ZN(new_n25911_));
  INV_X1     g22810(.I(new_n25911_), .ZN(new_n25912_));
  NOR2_X1    g22811(.A1(new_n25912_), .A2(new_n13713_), .ZN(new_n25913_));
  NAND2_X1   g22812(.A1(new_n25736_), .A2(new_n13713_), .ZN(new_n25914_));
  XNOR2_X1   g22813(.A1(new_n25913_), .A2(new_n25914_), .ZN(new_n25915_));
  AOI21_X1   g22814(.A1(new_n25915_), .A2(new_n12067_), .B(new_n25849_), .ZN(new_n25916_));
  MUX2_X1    g22815(.I0(new_n25916_), .I1(new_n25736_), .S(pi0647), .Z(new_n25917_));
  NAND2_X1   g22816(.A1(new_n25917_), .A2(new_n12049_), .ZN(new_n25918_));
  NAND2_X1   g22817(.A1(new_n25918_), .A2(pi0630), .ZN(new_n25919_));
  MUX2_X1    g22818(.I0(new_n25916_), .I1(new_n25736_), .S(new_n12061_), .Z(new_n25920_));
  NAND2_X1   g22819(.A1(new_n25920_), .A2(pi1157), .ZN(new_n25921_));
  NAND2_X1   g22820(.A1(new_n25921_), .A2(new_n12060_), .ZN(new_n25922_));
  AOI21_X1   g22821(.A1(new_n25919_), .A2(new_n25922_), .B(pi0787), .ZN(new_n25923_));
  NAND2_X1   g22822(.A1(new_n25923_), .A2(new_n25848_), .ZN(new_n25924_));
  NAND2_X1   g22823(.A1(new_n25915_), .A2(new_n12031_), .ZN(new_n25925_));
  AOI21_X1   g22824(.A1(new_n25735_), .A2(pi0628), .B(new_n24207_), .ZN(new_n25926_));
  NAND2_X1   g22825(.A1(new_n25925_), .A2(new_n25926_), .ZN(new_n25927_));
  NOR2_X1    g22826(.A1(new_n12050_), .A2(new_n12031_), .ZN(new_n25928_));
  AOI21_X1   g22827(.A1(new_n25915_), .A2(new_n25928_), .B(new_n24358_), .ZN(new_n25929_));
  NAND2_X1   g22828(.A1(new_n25927_), .A2(new_n25929_), .ZN(new_n25930_));
  NOR2_X1    g22829(.A1(new_n25846_), .A2(new_n25930_), .ZN(new_n25931_));
  MUX2_X1    g22830(.I0(new_n25911_), .I1(new_n25736_), .S(new_n12013_), .Z(new_n25932_));
  INV_X1     g22831(.I(new_n25932_), .ZN(new_n25933_));
  NAND2_X1   g22832(.A1(new_n25845_), .A2(new_n11994_), .ZN(new_n25934_));
  AOI21_X1   g22833(.A1(new_n25736_), .A2(pi0626), .B(new_n17171_), .ZN(new_n25935_));
  AOI22_X1   g22834(.A1(new_n25934_), .A2(new_n25935_), .B1(new_n17173_), .B2(new_n25933_), .ZN(new_n25936_));
  NOR4_X1    g22835(.A1(new_n25845_), .A2(new_n11994_), .A3(new_n11988_), .A4(new_n25736_), .ZN(new_n25937_));
  NOR3_X1    g22836(.A1(new_n25937_), .A2(pi0788), .A3(new_n25936_), .ZN(new_n25938_));
  OAI21_X1   g22837(.A1(new_n12443_), .A2(new_n13367_), .B(new_n25850_), .ZN(new_n25939_));
  NOR3_X1    g22838(.A1(new_n13368_), .A2(new_n24848_), .A3(new_n12114_), .ZN(new_n25940_));
  NAND2_X1   g22839(.A1(new_n25268_), .A2(pi0614), .ZN(new_n25941_));
  AND2_X2    g22840(.A1(new_n12356_), .A2(new_n25941_), .Z(new_n25942_));
  OAI21_X1   g22841(.A1(new_n25942_), .A2(new_n5095_), .B(new_n24848_), .ZN(new_n25943_));
  NOR2_X1    g22842(.A1(new_n12127_), .A2(pi0662), .ZN(new_n25944_));
  AOI21_X1   g22843(.A1(new_n25790_), .A2(new_n25944_), .B(new_n25794_), .ZN(new_n25945_));
  OAI21_X1   g22844(.A1(new_n25791_), .A2(new_n25943_), .B(new_n25945_), .ZN(new_n25946_));
  NAND2_X1   g22845(.A1(new_n25797_), .A2(new_n12464_), .ZN(new_n25947_));
  INV_X1     g22846(.I(new_n12468_), .ZN(new_n25948_));
  OAI21_X1   g22847(.A1(new_n25948_), .A2(new_n12465_), .B(new_n5104_), .ZN(new_n25949_));
  NOR3_X1    g22848(.A1(new_n12250_), .A2(new_n12258_), .A3(new_n12443_), .ZN(new_n25950_));
  NOR4_X1    g22849(.A1(new_n25288_), .A2(new_n12443_), .A3(pi0662), .A4(pi0680), .ZN(new_n25951_));
  NAND3_X1   g22850(.A1(new_n12466_), .A2(pi0614), .A3(new_n5095_), .ZN(new_n25952_));
  NOR3_X1    g22851(.A1(new_n25952_), .A2(new_n25951_), .A3(new_n25950_), .ZN(new_n25953_));
  AOI22_X1   g22852(.A1(new_n25949_), .A2(new_n25953_), .B1(new_n24848_), .B2(new_n25947_), .ZN(new_n25954_));
  NAND2_X1   g22853(.A1(new_n5141_), .A2(pi0224), .ZN(new_n25955_));
  OAI21_X1   g22854(.A1(new_n25946_), .A2(new_n25955_), .B(pi0223), .ZN(new_n25956_));
  NOR2_X1    g22855(.A1(new_n25743_), .A2(pi0680), .ZN(new_n25957_));
  NAND2_X1   g22856(.A1(new_n17309_), .A2(new_n12443_), .ZN(new_n25958_));
  OAI21_X1   g22857(.A1(new_n12443_), .A2(new_n25588_), .B(new_n25958_), .ZN(new_n25959_));
  NAND2_X1   g22858(.A1(new_n25959_), .A2(new_n25659_), .ZN(new_n25960_));
  AOI22_X1   g22859(.A1(new_n25960_), .A2(pi0616), .B1(pi0614), .B2(new_n12331_), .ZN(new_n25961_));
  AOI21_X1   g22860(.A1(new_n25229_), .A2(new_n25961_), .B(new_n5095_), .ZN(new_n25962_));
  XNOR2_X1   g22861(.A1(new_n25962_), .A2(new_n25957_), .ZN(new_n25963_));
  NAND2_X1   g22862(.A1(new_n25963_), .A2(new_n24848_), .ZN(new_n25964_));
  AOI22_X1   g22863(.A1(new_n25748_), .A2(new_n12129_), .B1(new_n25745_), .B2(new_n25944_), .ZN(new_n25965_));
  NAND3_X1   g22864(.A1(new_n25964_), .A2(new_n5141_), .A3(new_n25965_), .ZN(new_n25966_));
  INV_X1     g22865(.I(new_n25755_), .ZN(new_n25967_));
  OAI21_X1   g22866(.A1(new_n25219_), .A2(new_n12166_), .B(new_n12443_), .ZN(new_n25968_));
  NAND2_X1   g22867(.A1(new_n25223_), .A2(pi0614), .ZN(new_n25969_));
  XNOR2_X1   g22868(.A1(new_n25968_), .A2(new_n25969_), .ZN(new_n25970_));
  NAND2_X1   g22869(.A1(new_n25222_), .A2(new_n25970_), .ZN(new_n25971_));
  MUX2_X1    g22870(.I0(new_n25971_), .I1(new_n25967_), .S(new_n5095_), .Z(new_n25972_));
  NOR2_X1    g22871(.A1(new_n25972_), .A2(pi0662), .ZN(new_n25973_));
  INV_X1     g22872(.I(new_n25944_), .ZN(new_n25974_));
  OAI21_X1   g22873(.A1(new_n25755_), .A2(new_n25974_), .B(new_n25761_), .ZN(new_n25975_));
  OR3_X2     g22874(.A1(new_n25973_), .A2(new_n5141_), .A3(new_n25975_), .Z(new_n25976_));
  NAND3_X1   g22875(.A1(new_n25976_), .A2(new_n2595_), .A3(new_n25966_), .ZN(new_n25977_));
  MUX2_X1    g22876(.I0(new_n12491_), .I1(new_n12164_), .S(new_n12443_), .Z(new_n25978_));
  OAI21_X1   g22877(.A1(new_n25978_), .A2(pi0680), .B(new_n25766_), .ZN(new_n25979_));
  AOI21_X1   g22878(.A1(new_n25765_), .A2(new_n25944_), .B(new_n25767_), .ZN(new_n25980_));
  NOR2_X1    g22879(.A1(new_n25980_), .A2(new_n24848_), .ZN(new_n25981_));
  NAND2_X1   g22880(.A1(new_n25979_), .A2(new_n25981_), .ZN(new_n25982_));
  NAND2_X1   g22881(.A1(new_n12478_), .A2(new_n12443_), .ZN(new_n25983_));
  NOR2_X1    g22882(.A1(new_n25239_), .A2(pi0616), .ZN(new_n25984_));
  AOI21_X1   g22883(.A1(new_n25983_), .A2(new_n25984_), .B(new_n5095_), .ZN(new_n25985_));
  AOI21_X1   g22884(.A1(new_n25240_), .A2(new_n25775_), .B(new_n25985_), .ZN(new_n25986_));
  MUX2_X1    g22885(.I0(new_n25986_), .I1(new_n25770_), .S(new_n24848_), .Z(new_n25987_));
  OAI21_X1   g22886(.A1(new_n25982_), .A2(new_n25987_), .B(new_n5141_), .ZN(new_n25988_));
  NOR2_X1    g22887(.A1(new_n25988_), .A2(new_n4879_), .ZN(new_n25989_));
  NOR2_X1    g22888(.A1(new_n12478_), .A2(new_n25853_), .ZN(new_n25990_));
  OAI21_X1   g22889(.A1(new_n25990_), .A2(new_n25774_), .B(new_n2595_), .ZN(new_n25991_));
  OAI21_X1   g22890(.A1(new_n25991_), .A2(pi0222), .B(new_n2604_), .ZN(new_n25992_));
  OAI21_X1   g22891(.A1(new_n25989_), .A2(new_n25992_), .B(new_n25977_), .ZN(new_n25993_));
  AOI21_X1   g22892(.A1(new_n25993_), .A2(new_n25956_), .B(pi0299), .ZN(new_n25994_));
  AOI21_X1   g22893(.A1(new_n25982_), .A2(new_n2595_), .B(new_n5094_), .ZN(new_n25995_));
  OAI21_X1   g22894(.A1(new_n25973_), .A2(new_n25975_), .B(pi0224), .ZN(new_n25996_));
  OAI21_X1   g22895(.A1(new_n25996_), .A2(new_n25995_), .B(new_n3285_), .ZN(new_n25997_));
  NOR2_X1    g22896(.A1(new_n25784_), .A2(new_n12461_), .ZN(new_n25998_));
  NOR2_X1    g22897(.A1(new_n12386_), .A2(pi0616), .ZN(new_n25999_));
  NAND2_X1   g22898(.A1(new_n25999_), .A2(new_n25961_), .ZN(new_n26000_));
  MUX2_X1    g22899(.I0(new_n26000_), .I1(new_n25782_), .S(new_n5095_), .Z(new_n26001_));
  OAI22_X1   g22900(.A1(new_n26001_), .A2(pi0662), .B1(new_n25781_), .B2(new_n25974_), .ZN(new_n26002_));
  NOR2_X1    g22901(.A1(new_n26002_), .A2(new_n25998_), .ZN(new_n26003_));
  MUX2_X1    g22902(.I0(new_n26003_), .I1(new_n25946_), .S(new_n6445_), .Z(new_n26004_));
  NAND2_X1   g22903(.A1(new_n25797_), .A2(new_n24848_), .ZN(new_n26005_));
  OAI21_X1   g22904(.A1(new_n12476_), .A2(new_n5095_), .B(new_n25775_), .ZN(new_n26006_));
  NOR2_X1    g22905(.A1(new_n25985_), .A2(new_n24848_), .ZN(new_n26007_));
  NAND2_X1   g22906(.A1(new_n26006_), .A2(new_n26007_), .ZN(new_n26008_));
  AOI22_X1   g22907(.A1(new_n6445_), .A2(new_n25954_), .B1(new_n26008_), .B2(new_n26005_), .ZN(new_n26009_));
  NAND2_X1   g22908(.A1(new_n26008_), .A2(new_n26005_), .ZN(new_n26010_));
  NOR3_X1    g22909(.A1(new_n26010_), .A2(new_n5094_), .A3(new_n25954_), .ZN(new_n26011_));
  NOR3_X1    g22910(.A1(new_n26011_), .A2(pi0224), .A3(new_n26009_), .ZN(new_n26012_));
  OAI21_X1   g22911(.A1(new_n26004_), .A2(new_n2595_), .B(new_n26012_), .ZN(new_n26013_));
  NOR3_X1    g22912(.A1(new_n24848_), .A2(new_n5095_), .A3(pi0224), .ZN(new_n26014_));
  NAND2_X1   g22913(.A1(new_n25959_), .A2(new_n26014_), .ZN(new_n26015_));
  AOI21_X1   g22914(.A1(new_n26015_), .A2(new_n25991_), .B(new_n25773_), .ZN(new_n26016_));
  OAI21_X1   g22915(.A1(new_n26016_), .A2(pi0215), .B(new_n3154_), .ZN(new_n26017_));
  AOI21_X1   g22916(.A1(new_n26013_), .A2(new_n4905_), .B(new_n26017_), .ZN(new_n26018_));
  NAND2_X1   g22917(.A1(new_n25997_), .A2(new_n26018_), .ZN(new_n26019_));
  OAI21_X1   g22918(.A1(new_n25994_), .A2(new_n26019_), .B(new_n3172_), .ZN(new_n26020_));
  INV_X1     g22919(.I(new_n25310_), .ZN(new_n26021_));
  OAI21_X1   g22920(.A1(new_n13830_), .A2(pi0614), .B(pi0224), .ZN(new_n26022_));
  NOR2_X1    g22921(.A1(new_n25813_), .A2(new_n13358_), .ZN(new_n26023_));
  OAI22_X1   g22922(.A1(new_n26023_), .A2(pi0224), .B1(new_n26021_), .B2(new_n26022_), .ZN(new_n26024_));
  MUX2_X1    g22923(.I0(new_n25815_), .I1(new_n26024_), .S(new_n25853_), .Z(new_n26025_));
  NAND2_X1   g22924(.A1(new_n13355_), .A2(new_n25852_), .ZN(new_n26026_));
  AOI21_X1   g22925(.A1(new_n26026_), .A2(new_n25818_), .B(pi0224), .ZN(new_n26027_));
  AND4_X2    g22926(.A1(new_n13355_), .A2(new_n25816_), .A3(new_n25315_), .A4(new_n25853_), .Z(new_n26028_));
  OAI21_X1   g22927(.A1(new_n26028_), .A2(new_n26027_), .B(new_n2587_), .ZN(new_n26029_));
  NAND2_X1   g22928(.A1(new_n26029_), .A2(new_n3154_), .ZN(new_n26030_));
  AOI21_X1   g22929(.A1(new_n26025_), .A2(new_n2587_), .B(new_n26030_), .ZN(new_n26031_));
  AOI22_X1   g22930(.A1(new_n26020_), .A2(new_n26031_), .B1(new_n25939_), .B2(new_n25940_), .ZN(new_n26032_));
  NOR2_X1    g22931(.A1(new_n26032_), .A2(new_n3232_), .ZN(new_n26033_));
  XOR2_X1    g22932(.A1(new_n26033_), .A2(new_n25739_), .Z(new_n26034_));
  NAND2_X1   g22933(.A1(new_n26034_), .A2(pi0625), .ZN(new_n26035_));
  AOI21_X1   g22934(.A1(new_n25826_), .A2(pi0625), .B(new_n12978_), .ZN(new_n26036_));
  NAND2_X1   g22935(.A1(new_n26035_), .A2(new_n26036_), .ZN(new_n26037_));
  OAI21_X1   g22936(.A1(new_n25826_), .A2(pi0625), .B(new_n11893_), .ZN(new_n26038_));
  AOI21_X1   g22937(.A1(new_n26034_), .A2(pi0625), .B(new_n26038_), .ZN(new_n26039_));
  OAI21_X1   g22938(.A1(new_n26039_), .A2(new_n25903_), .B(new_n13657_), .ZN(new_n26040_));
  AOI21_X1   g22939(.A1(new_n26040_), .A2(new_n26037_), .B(new_n11891_), .ZN(new_n26041_));
  AOI21_X1   g22940(.A1(new_n11891_), .A2(new_n26034_), .B(new_n26041_), .ZN(new_n26042_));
  NOR4_X1    g22941(.A1(new_n26042_), .A2(new_n11903_), .A3(pi1155), .A4(new_n25906_), .ZN(new_n26043_));
  NAND4_X1   g22942(.A1(new_n25832_), .A2(new_n25831_), .A3(pi0660), .A4(new_n11912_), .ZN(new_n26044_));
  NOR3_X1    g22943(.A1(new_n25905_), .A2(new_n11903_), .A3(new_n11912_), .ZN(new_n26045_));
  OAI22_X1   g22944(.A1(new_n26043_), .A2(new_n26044_), .B1(pi0660), .B2(new_n26045_), .ZN(new_n26046_));
  MUX2_X1    g22945(.I0(new_n26046_), .I1(new_n26042_), .S(new_n11870_), .Z(new_n26047_));
  NAND2_X1   g22946(.A1(new_n26047_), .A2(new_n11969_), .ZN(new_n26048_));
  NAND2_X1   g22947(.A1(new_n11950_), .A2(pi0618), .ZN(new_n26049_));
  AOI21_X1   g22948(.A1(new_n25838_), .A2(pi0627), .B(new_n26049_), .ZN(new_n26050_));
  NAND2_X1   g22949(.A1(new_n26047_), .A2(new_n11934_), .ZN(new_n26051_));
  AOI21_X1   g22950(.A1(new_n25909_), .A2(pi0618), .B(new_n14687_), .ZN(new_n26052_));
  AOI22_X1   g22951(.A1(new_n26051_), .A2(new_n26052_), .B1(new_n26047_), .B2(new_n26050_), .ZN(new_n26053_));
  OR3_X2     g22952(.A1(new_n26053_), .A2(new_n11969_), .A3(new_n26048_), .Z(new_n26054_));
  OAI21_X1   g22953(.A1(new_n26053_), .A2(new_n11969_), .B(new_n26048_), .ZN(new_n26055_));
  NAND2_X1   g22954(.A1(new_n26054_), .A2(new_n26055_), .ZN(new_n26056_));
  INV_X1     g22955(.I(new_n26056_), .ZN(new_n26057_));
  NOR3_X1    g22956(.A1(new_n25911_), .A2(new_n11967_), .A3(new_n11869_), .ZN(new_n26058_));
  NOR2_X1    g22957(.A1(new_n26058_), .A2(pi0648), .ZN(new_n26059_));
  NAND2_X1   g22958(.A1(new_n26057_), .A2(pi0619), .ZN(new_n26060_));
  NOR3_X1    g22959(.A1(new_n25912_), .A2(new_n11967_), .A3(pi1159), .ZN(new_n26061_));
  AOI21_X1   g22960(.A1(new_n26060_), .A2(new_n26061_), .B(new_n25844_), .ZN(new_n26062_));
  OAI21_X1   g22961(.A1(new_n26057_), .A2(pi0789), .B(new_n11998_), .ZN(new_n26063_));
  NAND2_X1   g22962(.A1(new_n26063_), .A2(new_n17372_), .ZN(new_n26064_));
  NOR4_X1    g22963(.A1(new_n26062_), .A2(new_n26064_), .A3(new_n25938_), .A4(new_n26059_), .ZN(new_n26065_));
  OAI21_X1   g22964(.A1(new_n26065_), .A2(new_n25931_), .B(new_n14726_), .ZN(new_n26066_));
  AND2_X2    g22965(.A1(new_n26066_), .A2(new_n25924_), .Z(new_n26067_));
  OAI21_X1   g22966(.A1(new_n25735_), .A2(new_n12092_), .B(pi0644), .ZN(new_n26068_));
  AOI21_X1   g22967(.A1(new_n25847_), .A2(new_n12092_), .B(new_n26068_), .ZN(new_n26069_));
  AOI21_X1   g22968(.A1(pi0644), .A2(new_n25736_), .B(new_n26069_), .ZN(new_n26070_));
  OAI21_X1   g22969(.A1(new_n26070_), .A2(new_n12099_), .B(new_n12081_), .ZN(new_n26071_));
  NAND2_X1   g22970(.A1(new_n12082_), .A2(pi0715), .ZN(new_n26075_));
  AOI21_X1   g22971(.A1(new_n26066_), .A2(new_n25924_), .B(new_n26075_), .ZN(new_n26076_));
  OAI21_X1   g22972(.A1(new_n25736_), .A2(pi0644), .B(new_n12099_), .ZN(new_n26077_));
  OAI21_X1   g22973(.A1(new_n26069_), .A2(new_n26077_), .B(pi1160), .ZN(new_n26078_));
  NAND2_X1   g22974(.A1(new_n12099_), .A2(pi0644), .ZN(new_n26079_));
  AOI21_X1   g22975(.A1(new_n26066_), .A2(new_n25924_), .B(new_n26079_), .ZN(new_n26080_));
  AOI22_X1   g22976(.A1(new_n26071_), .A2(new_n26076_), .B1(new_n26080_), .B2(new_n26078_), .ZN(new_n26081_));
  MUX2_X1    g22977(.I0(new_n26081_), .I1(new_n26067_), .S(new_n11867_), .Z(new_n26082_));
  NAND2_X1   g22978(.A1(po1038), .A2(pi0224), .ZN(new_n26083_));
  OAI21_X1   g22979(.A1(new_n26082_), .A2(po1038), .B(new_n26083_), .ZN(po0381));
  OAI21_X1   g22980(.A1(new_n2869_), .A2(new_n2871_), .B(pi0137), .ZN(new_n26085_));
  NAND2_X1   g22981(.A1(new_n26085_), .A2(new_n3033_), .ZN(new_n26086_));
  NOR2_X1    g22982(.A1(new_n2857_), .A2(new_n8646_), .ZN(new_n26087_));
  NOR3_X1    g22983(.A1(new_n26087_), .A2(new_n2863_), .A3(new_n3105_), .ZN(new_n26088_));
  NOR2_X1    g22984(.A1(new_n26088_), .A2(new_n3091_), .ZN(new_n26089_));
  NOR2_X1    g22985(.A1(new_n26089_), .A2(new_n2656_), .ZN(new_n26090_));
  AOI21_X1   g22986(.A1(new_n2483_), .A2(new_n8646_), .B(new_n2971_), .ZN(new_n26091_));
  NOR4_X1    g22987(.A1(new_n26091_), .A2(pi0095), .A3(pi0137), .A4(new_n2656_), .ZN(new_n26092_));
  OAI21_X1   g22988(.A1(new_n26090_), .A2(new_n3039_), .B(new_n26092_), .ZN(new_n26093_));
  MUX2_X1    g22989(.I0(new_n26093_), .I1(new_n26086_), .S(new_n2563_), .Z(new_n26094_));
  OAI21_X1   g22990(.A1(new_n2911_), .A2(new_n2871_), .B(pi0137), .ZN(new_n26095_));
  NOR2_X1    g22991(.A1(new_n2994_), .A2(new_n2957_), .ZN(new_n26096_));
  NOR2_X1    g22992(.A1(new_n5971_), .A2(new_n2633_), .ZN(new_n26097_));
  AOI21_X1   g22993(.A1(new_n2895_), .A2(new_n26097_), .B(pi0032), .ZN(new_n26098_));
  INV_X1     g22994(.I(new_n26098_), .ZN(new_n26099_));
  AOI21_X1   g22995(.A1(new_n26099_), .A2(new_n26096_), .B(pi1093), .ZN(new_n26100_));
  OAI21_X1   g22996(.A1(new_n2956_), .A2(new_n2997_), .B(new_n26100_), .ZN(new_n26101_));
  OAI21_X1   g22997(.A1(new_n2924_), .A2(new_n2996_), .B(new_n26101_), .ZN(new_n26102_));
  NAND2_X1   g22998(.A1(new_n26102_), .A2(new_n8734_), .ZN(new_n26103_));
  NOR4_X1    g22999(.A1(new_n2995_), .A2(pi1093), .A3(new_n2956_), .A4(new_n2994_), .ZN(new_n26105_));
  INV_X1     g23000(.I(new_n26105_), .ZN(new_n26106_));
  NAND2_X1   g23001(.A1(new_n26101_), .A2(new_n26106_), .ZN(new_n26107_));
  NOR2_X1    g23002(.A1(new_n2922_), .A2(pi0137), .ZN(new_n26108_));
  AND2_X2    g23003(.A1(new_n26107_), .A2(new_n26108_), .Z(new_n26109_));
  INV_X1     g23004(.I(new_n26109_), .ZN(new_n26110_));
  NAND4_X1   g23005(.A1(new_n26095_), .A2(new_n2563_), .A3(new_n26103_), .A4(new_n26110_), .ZN(new_n26111_));
  OAI21_X1   g23006(.A1(new_n26089_), .A2(new_n2909_), .B(new_n2437_), .ZN(new_n26112_));
  NAND3_X1   g23007(.A1(new_n26112_), .A2(pi0137), .A3(new_n2872_), .ZN(new_n26113_));
  INV_X1     g23008(.I(new_n26091_), .ZN(new_n26114_));
  NAND4_X1   g23009(.A1(new_n26097_), .A2(new_n2658_), .A3(new_n2671_), .A4(pi0070), .ZN(new_n26115_));
  MUX2_X1    g23010(.I0(new_n26114_), .I1(new_n26115_), .S(new_n2957_), .Z(new_n26116_));
  NOR2_X1    g23011(.A1(new_n26116_), .A2(new_n2993_), .ZN(new_n26117_));
  NAND2_X1   g23012(.A1(new_n26117_), .A2(new_n26100_), .ZN(new_n26118_));
  OAI21_X1   g23013(.A1(new_n26091_), .A2(new_n2994_), .B(pi1093), .ZN(new_n26119_));
  NAND3_X1   g23014(.A1(new_n26118_), .A2(new_n8734_), .A3(new_n26119_), .ZN(new_n26120_));
  NAND2_X1   g23015(.A1(new_n26109_), .A2(new_n26117_), .ZN(new_n26121_));
  NAND4_X1   g23016(.A1(new_n26113_), .A2(pi0332), .A3(new_n26120_), .A4(new_n26121_), .ZN(new_n26122_));
  XNOR2_X1   g23017(.A1(new_n26122_), .A2(new_n26111_), .ZN(new_n26123_));
  NAND2_X1   g23018(.A1(new_n26123_), .A2(new_n2577_), .ZN(new_n26124_));
  NAND4_X1   g23019(.A1(new_n26124_), .A2(new_n2631_), .A3(new_n2587_), .A4(new_n26094_), .ZN(new_n26125_));
  AND2_X2    g23020(.A1(new_n26123_), .A2(new_n5161_), .Z(new_n26126_));
  NOR4_X1    g23021(.A1(new_n26126_), .A2(pi0198), .A3(pi0299), .A4(new_n26094_), .ZN(new_n26127_));
  NAND2_X1   g23022(.A1(new_n3172_), .A2(new_n3154_), .ZN(new_n26128_));
  AOI21_X1   g23023(.A1(new_n26127_), .A2(new_n26125_), .B(new_n26128_), .ZN(new_n26129_));
  NOR2_X1    g23024(.A1(new_n2436_), .A2(pi0038), .ZN(new_n26130_));
  AOI21_X1   g23025(.A1(new_n5153_), .A2(new_n26130_), .B(pi0100), .ZN(new_n26131_));
  OAI21_X1   g23026(.A1(new_n5163_), .A2(new_n5081_), .B(new_n2436_), .ZN(new_n26132_));
  AOI21_X1   g23027(.A1(new_n5160_), .A2(new_n26132_), .B(pi0087), .ZN(new_n26133_));
  OAI21_X1   g23028(.A1(new_n26129_), .A2(new_n26131_), .B(new_n26133_), .ZN(new_n26134_));
  NOR3_X1    g23029(.A1(new_n2491_), .A2(new_n2436_), .A3(new_n3198_), .ZN(new_n26135_));
  NAND2_X1   g23030(.A1(new_n26135_), .A2(pi0087), .ZN(new_n26136_));
  AOI21_X1   g23031(.A1(new_n26134_), .A2(new_n2628_), .B(new_n26136_), .ZN(new_n26137_));
  NAND3_X1   g23032(.A1(new_n5875_), .A2(new_n2628_), .A3(new_n26132_), .ZN(new_n26138_));
  NAND2_X1   g23033(.A1(new_n26138_), .A2(new_n3203_), .ZN(new_n26139_));
  NAND3_X1   g23034(.A1(new_n26135_), .A2(pi0092), .A3(new_n2534_), .ZN(new_n26140_));
  NAND2_X1   g23035(.A1(new_n26135_), .A2(new_n5196_), .ZN(new_n26141_));
  NAND4_X1   g23036(.A1(new_n26139_), .A2(new_n2538_), .A3(new_n26140_), .A4(new_n26141_), .ZN(new_n26142_));
  NOR3_X1    g23037(.A1(new_n2537_), .A2(pi0054), .A3(new_n3202_), .ZN(new_n26143_));
  AOI21_X1   g23038(.A1(new_n26135_), .A2(new_n26143_), .B(pi0055), .ZN(new_n26144_));
  OAI21_X1   g23039(.A1(new_n26137_), .A2(new_n26142_), .B(new_n26144_), .ZN(new_n26145_));
  OAI21_X1   g23040(.A1(pi0056), .A2(new_n5889_), .B(new_n26145_), .ZN(new_n26146_));
  NOR2_X1    g23041(.A1(new_n2543_), .A2(new_n3335_), .ZN(new_n26147_));
  AOI21_X1   g23042(.A1(new_n26135_), .A2(new_n26147_), .B(pi0062), .ZN(new_n26148_));
  NAND2_X1   g23043(.A1(new_n26135_), .A2(new_n3341_), .ZN(new_n26149_));
  OAI21_X1   g23044(.A1(new_n26149_), .A2(new_n3240_), .B(new_n2571_), .ZN(new_n26151_));
  AOI21_X1   g23045(.A1(new_n26146_), .A2(new_n26148_), .B(new_n26151_), .ZN(po0382));
  NAND2_X1   g23046(.A1(pi0228), .A2(pi0231), .ZN(new_n26153_));
  INV_X1     g23047(.I(new_n26153_), .ZN(new_n26154_));
  NAND2_X1   g23048(.A1(new_n3405_), .A2(new_n26154_), .ZN(new_n26155_));
  NAND2_X1   g23049(.A1(new_n26153_), .A2(pi0092), .ZN(new_n26156_));
  OAI21_X1   g23050(.A1(new_n5907_), .A2(new_n26154_), .B(new_n3177_), .ZN(new_n26157_));
  AOI21_X1   g23051(.A1(pi0035), .A2(new_n2851_), .B(new_n3058_), .ZN(new_n26158_));
  NOR2_X1    g23052(.A1(new_n26158_), .A2(pi0070), .ZN(new_n26159_));
  NAND2_X1   g23053(.A1(new_n2658_), .A2(pi0096), .ZN(new_n26160_));
  OAI21_X1   g23054(.A1(new_n26159_), .A2(new_n26160_), .B(new_n3107_), .ZN(new_n26161_));
  AOI21_X1   g23055(.A1(new_n26161_), .A2(new_n5086_), .B(new_n3077_), .ZN(new_n26162_));
  OR3_X2     g23056(.A1(new_n26162_), .A2(new_n3154_), .A3(new_n2491_), .Z(new_n26163_));
  OAI21_X1   g23057(.A1(new_n3154_), .A2(new_n2490_), .B(new_n26162_), .ZN(new_n26164_));
  AOI21_X1   g23058(.A1(new_n26163_), .A2(new_n26164_), .B(pi0038), .ZN(new_n26165_));
  MUX2_X1    g23059(.I0(new_n26165_), .I1(pi0231), .S(pi0228), .Z(new_n26166_));
  NAND2_X1   g23060(.A1(new_n26166_), .A2(new_n3173_), .ZN(new_n26167_));
  NAND2_X1   g23061(.A1(new_n10248_), .A2(new_n26153_), .ZN(new_n26168_));
  AOI21_X1   g23062(.A1(new_n26168_), .A2(pi0100), .B(pi0087), .ZN(new_n26169_));
  AOI22_X1   g23063(.A1(new_n26167_), .A2(new_n26169_), .B1(new_n2628_), .B2(new_n26157_), .ZN(new_n26170_));
  OAI21_X1   g23064(.A1(new_n10222_), .A2(new_n26154_), .B(pi0075), .ZN(new_n26171_));
  NAND2_X1   g23065(.A1(new_n26171_), .A2(new_n3203_), .ZN(new_n26172_));
  OAI22_X1   g23066(.A1(new_n26170_), .A2(new_n26172_), .B1(new_n5910_), .B2(new_n26156_), .ZN(new_n26173_));
  MUX2_X1    g23067(.I0(new_n26173_), .I1(new_n26153_), .S(pi0054), .Z(new_n26174_));
  OAI21_X1   g23068(.A1(new_n3311_), .A2(new_n8423_), .B(new_n26153_), .ZN(new_n26175_));
  AOI21_X1   g23069(.A1(new_n26175_), .A2(pi0074), .B(pi0055), .ZN(new_n26176_));
  OAI21_X1   g23070(.A1(new_n26174_), .A2(pi0074), .B(new_n26176_), .ZN(new_n26177_));
  AOI21_X1   g23071(.A1(new_n26153_), .A2(pi0055), .B(pi0056), .ZN(new_n26178_));
  NAND3_X1   g23072(.A1(new_n5921_), .A2(new_n3335_), .A3(new_n26153_), .ZN(new_n26179_));
  NAND4_X1   g23073(.A1(new_n5925_), .A2(new_n3240_), .A3(new_n26153_), .A4(new_n26179_), .ZN(new_n26180_));
  AOI21_X1   g23074(.A1(new_n26177_), .A2(new_n26178_), .B(new_n26180_), .ZN(new_n26181_));
  OAI21_X1   g23075(.A1(new_n26181_), .A2(new_n3405_), .B(new_n26155_), .ZN(po0383));
  NAND2_X1   g23076(.A1(new_n2662_), .A2(pi0047), .ZN(new_n26183_));
  OAI21_X1   g23077(.A1(new_n2635_), .A2(new_n26183_), .B(new_n2660_), .ZN(new_n26184_));
  INV_X1     g23078(.I(new_n26184_), .ZN(new_n26185_));
  NOR2_X1    g23079(.A1(new_n5303_), .A2(new_n2652_), .ZN(new_n26186_));
  AOI21_X1   g23080(.A1(new_n26186_), .A2(new_n26185_), .B(pi0072), .ZN(new_n26187_));
  INV_X1     g23081(.I(new_n26187_), .ZN(new_n26188_));
  NAND3_X1   g23082(.A1(new_n8398_), .A2(new_n6005_), .A3(new_n26186_), .ZN(new_n26189_));
  AOI21_X1   g23083(.A1(new_n26189_), .A2(new_n6977_), .B(new_n26188_), .ZN(new_n26190_));
  NOR4_X1    g23084(.A1(new_n9692_), .A2(new_n2652_), .A3(new_n10561_), .A4(new_n6005_), .ZN(new_n26191_));
  NAND2_X1   g23085(.A1(new_n5365_), .A2(pi1093), .ZN(new_n26192_));
  OAI22_X1   g23086(.A1(new_n26191_), .A2(new_n26192_), .B1(new_n26190_), .B2(new_n10561_), .ZN(new_n26193_));
  NAND4_X1   g23087(.A1(new_n8407_), .A2(new_n5366_), .A3(new_n8437_), .A4(new_n8404_), .ZN(new_n26194_));
  NAND4_X1   g23088(.A1(new_n8398_), .A2(new_n2955_), .A3(new_n26185_), .A4(new_n26194_), .ZN(new_n26195_));
  AOI21_X1   g23089(.A1(new_n26195_), .A2(new_n26186_), .B(pi0072), .ZN(new_n26196_));
  NOR2_X1    g23090(.A1(new_n5113_), .A2(new_n2927_), .ZN(new_n26197_));
  OAI21_X1   g23091(.A1(new_n26196_), .A2(new_n10561_), .B(new_n26197_), .ZN(new_n26198_));
  NAND2_X1   g23092(.A1(new_n8398_), .A2(new_n26186_), .ZN(new_n26199_));
  NAND4_X1   g23093(.A1(new_n26199_), .A2(new_n10561_), .A3(new_n9859_), .A4(new_n26187_), .ZN(new_n26200_));
  NAND3_X1   g23094(.A1(new_n26193_), .A2(new_n26198_), .A3(new_n26200_), .ZN(new_n26201_));
  AOI21_X1   g23095(.A1(new_n26201_), .A2(new_n3154_), .B(new_n8676_), .ZN(po0384));
  NAND3_X1   g23096(.A1(new_n5362_), .A2(pi1091), .A3(new_n8655_), .ZN(new_n26203_));
  NOR2_X1    g23097(.A1(new_n5145_), .A2(new_n3296_), .ZN(new_n26204_));
  OAI21_X1   g23098(.A1(new_n8651_), .A2(new_n26204_), .B(pi0039), .ZN(new_n26205_));
  NOR2_X1    g23099(.A1(new_n26203_), .A2(new_n26205_), .ZN(new_n26206_));
  NOR2_X1    g23100(.A1(pi0039), .A2(pi0095), .ZN(new_n26207_));
  NAND2_X1   g23101(.A1(new_n8771_), .A2(new_n7756_), .ZN(new_n26208_));
  NAND4_X1   g23102(.A1(new_n2875_), .A2(new_n2632_), .A3(new_n26207_), .A4(new_n26208_), .ZN(new_n26209_));
  OAI21_X1   g23103(.A1(new_n26209_), .A2(new_n8697_), .B(new_n7855_), .ZN(new_n26210_));
  OAI22_X1   g23104(.A1(new_n26206_), .A2(new_n26210_), .B1(pi0039), .B2(new_n2523_), .ZN(po0385));
  NAND2_X1   g23105(.A1(new_n12593_), .A2(new_n2632_), .ZN(new_n26212_));
  NOR3_X1    g23106(.A1(new_n12534_), .A2(new_n2927_), .A3(new_n2918_), .ZN(new_n26213_));
  AOI21_X1   g23107(.A1(new_n26212_), .A2(new_n26213_), .B(pi0824), .ZN(new_n26214_));
  NOR3_X1    g23108(.A1(new_n26214_), .A2(new_n2927_), .A3(new_n2918_), .ZN(new_n26215_));
  INV_X1     g23109(.I(new_n12533_), .ZN(new_n26216_));
  NOR3_X1    g23110(.A1(new_n26216_), .A2(pi0824), .A3(new_n12534_), .ZN(new_n26217_));
  OR3_X2     g23111(.A1(new_n26217_), .A2(new_n2955_), .A3(new_n5081_), .Z(new_n26218_));
  OAI22_X1   g23112(.A1(new_n26218_), .A2(new_n26215_), .B1(new_n2918_), .B2(new_n2958_), .ZN(new_n26219_));
  NOR2_X1    g23113(.A1(new_n2958_), .A2(new_n2918_), .ZN(new_n26220_));
  NOR2_X1    g23114(.A1(new_n26217_), .A2(new_n26220_), .ZN(new_n26221_));
  AOI21_X1   g23115(.A1(new_n26221_), .A2(new_n26214_), .B(new_n12552_), .ZN(new_n26222_));
  INV_X1     g23116(.I(new_n12552_), .ZN(new_n26223_));
  OAI21_X1   g23117(.A1(new_n26223_), .A2(new_n6004_), .B(new_n12577_), .ZN(new_n26224_));
  NOR2_X1    g23118(.A1(new_n5081_), .A2(new_n26220_), .ZN(new_n26225_));
  AOI21_X1   g23119(.A1(new_n26224_), .A2(new_n26225_), .B(new_n2924_), .ZN(new_n26226_));
  NOR2_X1    g23120(.A1(new_n12524_), .A2(new_n5083_), .ZN(new_n26227_));
  OAI21_X1   g23121(.A1(pi0047), .A2(new_n12541_), .B(new_n26227_), .ZN(new_n26228_));
  AOI21_X1   g23122(.A1(new_n26228_), .A2(new_n12546_), .B(new_n3181_), .ZN(new_n26229_));
  OR2_X2     g23123(.A1(new_n26229_), .A2(new_n12549_), .Z(new_n26230_));
  NOR4_X1    g23124(.A1(new_n26230_), .A2(pi1093), .A3(new_n5181_), .A4(new_n26223_), .ZN(new_n26231_));
  NOR4_X1    g23125(.A1(new_n26222_), .A2(pi0039), .A3(new_n26226_), .A4(new_n26231_), .ZN(new_n26232_));
  NOR2_X1    g23126(.A1(new_n6037_), .A2(new_n5114_), .ZN(new_n26233_));
  NAND4_X1   g23127(.A1(new_n12149_), .A2(new_n2918_), .A3(new_n12173_), .A4(new_n26233_), .ZN(new_n26234_));
  INV_X1     g23128(.I(new_n26234_), .ZN(new_n26235_));
  NOR2_X1    g23129(.A1(new_n12339_), .A2(new_n5368_), .ZN(new_n26236_));
  NOR2_X1    g23130(.A1(pi0120), .A2(pi1091), .ZN(new_n26237_));
  NAND2_X1   g23131(.A1(new_n12138_), .A2(new_n5367_), .ZN(new_n26238_));
  NAND4_X1   g23132(.A1(new_n26238_), .A2(pi0120), .A3(new_n2490_), .A4(new_n26237_), .ZN(new_n26239_));
  NOR3_X1    g23133(.A1(new_n26235_), .A2(new_n26236_), .A3(new_n26239_), .ZN(new_n26240_));
  INV_X1     g23134(.I(new_n26240_), .ZN(new_n26241_));
  NOR2_X1    g23135(.A1(new_n12681_), .A2(new_n5143_), .ZN(new_n26242_));
  AOI21_X1   g23136(.A1(new_n26241_), .A2(new_n5143_), .B(new_n26242_), .ZN(new_n26243_));
  OR2_X2     g23137(.A1(new_n26243_), .A2(new_n6445_), .Z(new_n26244_));
  NOR2_X1    g23138(.A1(new_n6446_), .A2(new_n12681_), .ZN(new_n26245_));
  AOI21_X1   g23139(.A1(new_n26241_), .A2(new_n6446_), .B(new_n26245_), .ZN(new_n26246_));
  AOI21_X1   g23140(.A1(new_n26246_), .A2(new_n5094_), .B(new_n3284_), .ZN(new_n26247_));
  NAND4_X1   g23141(.A1(new_n6446_), .A2(pi0120), .A3(new_n5126_), .A4(new_n12680_), .ZN(new_n26248_));
  NOR4_X1    g23142(.A1(new_n6548_), .A2(new_n10267_), .A3(new_n2490_), .A4(new_n5129_), .ZN(new_n26249_));
  OAI21_X1   g23143(.A1(new_n26248_), .A2(new_n26249_), .B(new_n5094_), .ZN(new_n26250_));
  NAND2_X1   g23144(.A1(new_n12681_), .A2(new_n3284_), .ZN(new_n26251_));
  AOI21_X1   g23145(.A1(new_n26251_), .A2(new_n2566_), .B(pi0299), .ZN(new_n26252_));
  OAI21_X1   g23146(.A1(new_n26250_), .A2(new_n2566_), .B(new_n26252_), .ZN(new_n26253_));
  AOI21_X1   g23147(.A1(new_n26244_), .A2(new_n26247_), .B(new_n26253_), .ZN(new_n26254_));
  NOR2_X1    g23148(.A1(new_n26243_), .A2(new_n6460_), .ZN(new_n26255_));
  NAND2_X1   g23149(.A1(new_n26246_), .A2(new_n5141_), .ZN(new_n26256_));
  NOR3_X1    g23150(.A1(new_n2614_), .A2(pi0223), .A3(pi0299), .ZN(new_n26258_));
  NAND2_X1   g23151(.A1(new_n26256_), .A2(new_n26258_), .ZN(new_n26259_));
  OAI21_X1   g23152(.A1(new_n26259_), .A2(new_n26255_), .B(new_n3154_), .ZN(new_n26260_));
  NOR3_X1    g23153(.A1(new_n5154_), .A2(pi0038), .A3(new_n7832_), .ZN(new_n26261_));
  OAI21_X1   g23154(.A1(new_n26260_), .A2(new_n26254_), .B(new_n26261_), .ZN(new_n26262_));
  AOI21_X1   g23155(.A1(new_n26232_), .A2(new_n26219_), .B(new_n26262_), .ZN(po0387));
  INV_X1     g23156(.I(new_n11302_), .ZN(new_n26264_));
  INV_X1     g23157(.I(new_n5881_), .ZN(new_n26265_));
  NOR2_X1    g23158(.A1(new_n5146_), .A2(pi0299), .ZN(new_n26266_));
  AOI21_X1   g23159(.A1(new_n5866_), .A2(pi0299), .B(new_n26266_), .ZN(new_n26267_));
  NOR2_X1    g23160(.A1(new_n5117_), .A2(new_n2955_), .ZN(new_n26268_));
  NAND4_X1   g23161(.A1(new_n26267_), .A2(pi0835), .A3(new_n8648_), .A4(new_n26268_), .ZN(new_n26269_));
  NAND4_X1   g23162(.A1(new_n26269_), .A2(new_n8018_), .A3(new_n8648_), .A4(new_n8619_), .ZN(new_n26270_));
  NOR2_X1    g23163(.A1(new_n2669_), .A2(new_n2841_), .ZN(new_n26271_));
  INV_X1     g23164(.I(new_n2824_), .ZN(new_n26272_));
  MUX2_X1    g23165(.I0(new_n2805_), .I1(new_n2699_), .S(pi0081), .Z(new_n26273_));
  NOR2_X1    g23166(.A1(new_n26273_), .A2(pi0102), .ZN(new_n26274_));
  NAND3_X1   g23167(.A1(new_n2713_), .A2(new_n2709_), .A3(new_n2463_), .ZN(new_n26275_));
  NOR2_X1    g23168(.A1(new_n5279_), .A2(new_n2696_), .ZN(new_n26276_));
  OAI21_X1   g23169(.A1(new_n26274_), .A2(new_n26275_), .B(new_n26276_), .ZN(new_n26277_));
  NOR2_X1    g23170(.A1(new_n2694_), .A2(pi0086), .ZN(new_n26278_));
  AOI21_X1   g23171(.A1(new_n26277_), .A2(new_n26278_), .B(new_n26272_), .ZN(new_n26279_));
  OAI21_X1   g23172(.A1(new_n26279_), .A2(new_n2689_), .B(new_n2829_), .ZN(new_n26280_));
  AOI21_X1   g23173(.A1(new_n26280_), .A2(new_n2833_), .B(new_n2679_), .ZN(new_n26281_));
  OAI21_X1   g23174(.A1(new_n26281_), .A2(new_n2678_), .B(new_n3055_), .ZN(new_n26282_));
  NAND2_X1   g23175(.A1(new_n26282_), .A2(pi0093), .ZN(new_n26283_));
  XOR2_X1    g23176(.A1(new_n26283_), .A2(new_n2670_), .Z(new_n26284_));
  NAND2_X1   g23177(.A1(new_n26284_), .A2(new_n2876_), .ZN(new_n26285_));
  NAND2_X1   g23178(.A1(new_n26285_), .A2(new_n26271_), .ZN(new_n26286_));
  NOR2_X1    g23179(.A1(new_n26285_), .A2(new_n26271_), .ZN(new_n26287_));
  NOR2_X1    g23180(.A1(new_n26287_), .A2(new_n2849_), .ZN(new_n26288_));
  AOI21_X1   g23181(.A1(pi0070), .A2(new_n2671_), .B(new_n3105_), .ZN(new_n26289_));
  NAND4_X1   g23182(.A1(new_n2864_), .A2(new_n2658_), .A3(new_n2675_), .A4(new_n26289_), .ZN(new_n26290_));
  AOI21_X1   g23183(.A1(new_n26288_), .A2(new_n26286_), .B(new_n26290_), .ZN(new_n26291_));
  NOR2_X1    g23184(.A1(new_n2858_), .A2(pi1082), .ZN(new_n26292_));
  OAI21_X1   g23185(.A1(new_n26291_), .A2(new_n26292_), .B(new_n2632_), .ZN(new_n26293_));
  AOI21_X1   g23186(.A1(new_n2655_), .A2(pi0032), .B(pi0095), .ZN(new_n26294_));
  AOI21_X1   g23187(.A1(new_n26293_), .A2(new_n26294_), .B(new_n2871_), .ZN(new_n26295_));
  MUX2_X1    g23188(.I0(new_n26295_), .I1(new_n2490_), .S(pi0039), .Z(new_n26296_));
  NAND2_X1   g23189(.A1(new_n26296_), .A2(new_n26270_), .ZN(new_n26297_));
  MUX2_X1    g23190(.I0(new_n26297_), .I1(new_n5154_), .S(pi0038), .Z(new_n26298_));
  NOR2_X1    g23191(.A1(new_n26298_), .A2(pi0100), .ZN(new_n26299_));
  OAI21_X1   g23192(.A1(new_n26299_), .A2(new_n5160_), .B(new_n3177_), .ZN(new_n26300_));
  AOI21_X1   g23193(.A1(new_n5056_), .A2(pi0087), .B(new_n3228_), .ZN(new_n26301_));
  AOI21_X1   g23194(.A1(new_n26300_), .A2(new_n26301_), .B(new_n26265_), .ZN(new_n26302_));
  OAI21_X1   g23195(.A1(new_n26302_), .A2(pi0054), .B(new_n26264_), .ZN(new_n26303_));
  AOI21_X1   g23196(.A1(new_n26303_), .A2(new_n6962_), .B(new_n11295_), .ZN(new_n26304_));
  OAI21_X1   g23197(.A1(new_n26304_), .A2(pi0056), .B(new_n11294_), .ZN(new_n26305_));
  AOI21_X1   g23198(.A1(new_n26305_), .A2(new_n11308_), .B(new_n11309_), .ZN(po0389));
  INV_X1     g23199(.I(pi0230), .ZN(new_n26307_));
  NOR2_X1    g23200(.A1(pi0212), .A2(pi0214), .ZN(new_n26308_));
  NOR2_X1    g23201(.A1(new_n26308_), .A2(pi0211), .ZN(new_n26309_));
  NOR2_X1    g23202(.A1(new_n26309_), .A2(new_n8247_), .ZN(new_n26310_));
  NOR2_X1    g23203(.A1(new_n6845_), .A2(new_n26310_), .ZN(new_n26311_));
  NOR2_X1    g23204(.A1(pi0211), .A2(pi1144), .ZN(new_n26312_));
  AOI21_X1   g23205(.A1(pi0211), .A2(new_n3548_), .B(new_n26312_), .ZN(new_n26313_));
  NOR2_X1    g23206(.A1(new_n8248_), .A2(new_n26308_), .ZN(new_n26314_));
  NOR2_X1    g23207(.A1(new_n3548_), .A2(pi0211), .ZN(new_n26315_));
  AOI22_X1   g23208(.A1(new_n26314_), .A2(new_n26313_), .B1(new_n8248_), .B2(new_n26315_), .ZN(new_n26316_));
  OAI22_X1   g23209(.A1(new_n8082_), .A2(new_n3700_), .B1(new_n26316_), .B2(pi0219), .ZN(new_n26317_));
  AND2_X2    g23210(.A1(new_n26317_), .A2(new_n26311_), .Z(new_n26318_));
  INV_X1     g23211(.I(new_n26309_), .ZN(new_n26319_));
  NOR2_X1    g23212(.A1(new_n3548_), .A2(pi0199), .ZN(new_n26320_));
  INV_X1     g23213(.I(new_n26320_), .ZN(new_n26321_));
  NAND2_X1   g23214(.A1(new_n26321_), .A2(pi0200), .ZN(new_n26322_));
  AOI21_X1   g23215(.A1(pi0199), .A2(pi1142), .B(pi0200), .ZN(new_n26323_));
  NOR2_X1    g23216(.A1(new_n2552_), .A2(pi0199), .ZN(new_n26324_));
  INV_X1     g23217(.I(new_n26324_), .ZN(new_n26325_));
  OAI21_X1   g23218(.A1(new_n26323_), .A2(new_n26325_), .B(new_n26322_), .ZN(new_n26326_));
  AOI21_X1   g23219(.A1(new_n26326_), .A2(pi0207), .B(pi0208), .ZN(new_n26327_));
  NOR2_X1    g23220(.A1(new_n8087_), .A2(pi0299), .ZN(new_n26328_));
  NOR2_X1    g23221(.A1(new_n3700_), .A2(pi0199), .ZN(new_n26329_));
  INV_X1     g23222(.I(new_n26329_), .ZN(new_n26330_));
  NOR3_X1    g23223(.A1(new_n26330_), .A2(pi0200), .A3(new_n26328_), .ZN(new_n26331_));
  INV_X1     g23224(.I(new_n26323_), .ZN(new_n26332_));
  NAND2_X1   g23225(.A1(new_n26332_), .A2(new_n26320_), .ZN(new_n26333_));
  NOR2_X1    g23226(.A1(new_n26326_), .A2(pi0299), .ZN(new_n26334_));
  OAI22_X1   g23227(.A1(new_n26334_), .A2(pi0207), .B1(new_n26331_), .B2(new_n26333_), .ZN(new_n26335_));
  NAND2_X1   g23228(.A1(new_n26335_), .A2(pi0208), .ZN(new_n26336_));
  XNOR2_X1   g23229(.A1(new_n26336_), .A2(new_n26327_), .ZN(new_n26337_));
  MUX2_X1    g23230(.I0(new_n26337_), .I1(new_n3700_), .S(new_n2587_), .Z(new_n26338_));
  INV_X1     g23231(.I(new_n26337_), .ZN(new_n26339_));
  NOR2_X1    g23232(.A1(new_n26339_), .A2(pi0299), .ZN(new_n26340_));
  NAND4_X1   g23233(.A1(new_n26338_), .A2(new_n26340_), .A3(new_n8247_), .A4(new_n26319_), .ZN(new_n26341_));
  INV_X1     g23234(.I(new_n26308_), .ZN(new_n26342_));
  INV_X1     g23235(.I(new_n26340_), .ZN(new_n26343_));
  MUX2_X1    g23236(.I0(pi1143), .I1(pi1142), .S(pi0211), .Z(new_n26344_));
  NAND2_X1   g23237(.A1(new_n26344_), .A2(pi0299), .ZN(new_n26345_));
  AOI21_X1   g23238(.A1(new_n26343_), .A2(new_n26345_), .B(new_n26342_), .ZN(new_n26346_));
  INV_X1     g23239(.I(new_n26313_), .ZN(new_n26347_));
  NOR2_X1    g23240(.A1(new_n26347_), .A2(new_n2587_), .ZN(new_n26348_));
  NOR4_X1    g23241(.A1(new_n26346_), .A2(pi0214), .A3(new_n26340_), .A4(new_n26348_), .ZN(new_n26349_));
  AOI21_X1   g23242(.A1(pi0214), .A2(new_n26348_), .B(new_n26340_), .ZN(new_n26350_));
  NOR2_X1    g23243(.A1(po1038), .A2(pi0219), .ZN(new_n26351_));
  OAI21_X1   g23244(.A1(new_n26350_), .A2(pi0212), .B(new_n26351_), .ZN(new_n26352_));
  NOR2_X1    g23245(.A1(new_n26349_), .A2(new_n26352_), .ZN(new_n26353_));
  AOI21_X1   g23246(.A1(new_n26353_), .A2(new_n26341_), .B(new_n26318_), .ZN(new_n26354_));
  NOR2_X1    g23247(.A1(new_n8247_), .A2(pi0211), .ZN(new_n26355_));
  NOR2_X1    g23248(.A1(new_n2587_), .A2(new_n11950_), .ZN(new_n26356_));
  INV_X1     g23249(.I(new_n26356_), .ZN(new_n26357_));
  NOR2_X1    g23250(.A1(new_n2587_), .A2(new_n11893_), .ZN(new_n26358_));
  INV_X1     g23251(.I(new_n26358_), .ZN(new_n26359_));
  MUX2_X1    g23252(.I0(new_n26357_), .I1(new_n26359_), .S(pi0214), .Z(new_n26360_));
  NOR2_X1    g23253(.A1(new_n8078_), .A2(pi0212), .ZN(new_n26361_));
  INV_X1     g23254(.I(new_n26361_), .ZN(new_n26362_));
  NOR2_X1    g23255(.A1(new_n2587_), .A2(new_n11912_), .ZN(new_n26363_));
  INV_X1     g23256(.I(new_n26363_), .ZN(new_n26364_));
  OAI22_X1   g23257(.A1(new_n26360_), .A2(new_n8076_), .B1(new_n26362_), .B2(new_n26364_), .ZN(new_n26365_));
  NOR2_X1    g23258(.A1(new_n8077_), .A2(new_n12026_), .ZN(new_n26366_));
  NOR2_X1    g23259(.A1(new_n12049_), .A2(pi0211), .ZN(new_n26367_));
  NOR2_X1    g23260(.A1(new_n26366_), .A2(new_n26367_), .ZN(new_n26368_));
  OAI21_X1   g23261(.A1(new_n26368_), .A2(new_n8078_), .B(new_n8076_), .ZN(new_n26369_));
  NOR2_X1    g23262(.A1(new_n2587_), .A2(pi0219), .ZN(new_n26370_));
  AOI22_X1   g23263(.A1(new_n26365_), .A2(new_n26355_), .B1(new_n26369_), .B2(new_n26370_), .ZN(new_n26371_));
  AND2_X2    g23264(.A1(new_n26343_), .A2(new_n26371_), .Z(new_n26372_));
  NOR4_X1    g23265(.A1(new_n26372_), .A2(pi0209), .A3(new_n24753_), .A4(po1038), .ZN(new_n26373_));
  INV_X1     g23266(.I(pi0209), .ZN(new_n26374_));
  NOR2_X1    g23267(.A1(new_n26308_), .A2(pi0219), .ZN(new_n26375_));
  NOR2_X1    g23268(.A1(new_n26309_), .A2(new_n26375_), .ZN(new_n26376_));
  NOR2_X1    g23269(.A1(new_n8098_), .A2(pi1155), .ZN(new_n26377_));
  NOR3_X1    g23270(.A1(new_n8170_), .A2(new_n26377_), .A3(new_n12026_), .ZN(new_n26378_));
  NOR2_X1    g23271(.A1(new_n8098_), .A2(pi0299), .ZN(new_n26379_));
  INV_X1     g23272(.I(new_n26379_), .ZN(new_n26380_));
  NOR2_X1    g23273(.A1(new_n11912_), .A2(pi0199), .ZN(new_n26381_));
  INV_X1     g23274(.I(new_n26381_), .ZN(new_n26382_));
  NOR2_X1    g23275(.A1(new_n26380_), .A2(new_n26382_), .ZN(new_n26383_));
  NOR2_X1    g23276(.A1(new_n26383_), .A2(pi1154), .ZN(new_n26384_));
  NOR2_X1    g23277(.A1(new_n26381_), .A2(new_n8098_), .ZN(new_n26385_));
  OAI21_X1   g23278(.A1(new_n26384_), .A2(new_n26385_), .B(new_n8269_), .ZN(new_n26386_));
  INV_X1     g23279(.I(new_n26386_), .ZN(new_n26387_));
  NOR2_X1    g23280(.A1(new_n26387_), .A2(new_n26378_), .ZN(new_n26388_));
  NOR2_X1    g23281(.A1(pi0200), .A2(pi0299), .ZN(new_n26389_));
  INV_X1     g23282(.I(new_n26389_), .ZN(new_n26390_));
  NOR2_X1    g23283(.A1(new_n8094_), .A2(pi1153), .ZN(new_n26391_));
  NOR2_X1    g23284(.A1(pi0199), .A2(pi1155), .ZN(new_n26392_));
  NOR4_X1    g23285(.A1(new_n26390_), .A2(new_n26391_), .A3(pi1154), .A4(new_n26392_), .ZN(new_n26393_));
  NOR2_X1    g23286(.A1(new_n8098_), .A2(pi0199), .ZN(new_n26394_));
  NOR2_X1    g23287(.A1(new_n8094_), .A2(pi0200), .ZN(new_n26395_));
  NOR2_X1    g23288(.A1(new_n26394_), .A2(new_n26395_), .ZN(new_n26396_));
  NOR2_X1    g23289(.A1(new_n26396_), .A2(new_n11950_), .ZN(new_n26397_));
  INV_X1     g23290(.I(new_n26397_), .ZN(new_n26398_));
  NOR2_X1    g23291(.A1(new_n11912_), .A2(pi0200), .ZN(new_n26399_));
  NOR2_X1    g23292(.A1(new_n26397_), .A2(new_n26399_), .ZN(new_n26400_));
  OAI22_X1   g23293(.A1(new_n26400_), .A2(new_n8170_), .B1(new_n26398_), .B2(new_n11893_), .ZN(new_n26401_));
  NOR2_X1    g23294(.A1(new_n8094_), .A2(new_n8098_), .ZN(new_n26402_));
  NOR2_X1    g23295(.A1(new_n26402_), .A2(pi0299), .ZN(new_n26403_));
  NOR2_X1    g23296(.A1(new_n26403_), .A2(new_n11893_), .ZN(new_n26404_));
  OR2_X2     g23297(.A1(new_n26401_), .A2(new_n26404_), .Z(new_n26405_));
  AOI21_X1   g23298(.A1(new_n26405_), .A2(new_n11950_), .B(new_n26393_), .ZN(new_n26406_));
  MUX2_X1    g23299(.I0(new_n26406_), .I1(new_n26388_), .S(new_n8087_), .Z(new_n26407_));
  NOR2_X1    g23300(.A1(new_n26407_), .A2(new_n8088_), .ZN(new_n26408_));
  NOR3_X1    g23301(.A1(new_n8094_), .A2(new_n11912_), .A3(pi0200), .ZN(new_n26409_));
  AOI21_X1   g23302(.A1(new_n26409_), .A2(new_n2587_), .B(pi1156), .ZN(new_n26410_));
  NOR2_X1    g23303(.A1(new_n26396_), .A2(pi0299), .ZN(new_n26411_));
  INV_X1     g23304(.I(new_n26411_), .ZN(new_n26412_));
  NOR2_X1    g23305(.A1(pi0200), .A2(pi1155), .ZN(new_n26413_));
  NOR3_X1    g23306(.A1(new_n26412_), .A2(new_n26410_), .A3(new_n26413_), .ZN(new_n26414_));
  INV_X1     g23307(.I(new_n26414_), .ZN(new_n26415_));
  NOR2_X1    g23308(.A1(new_n26415_), .A2(new_n8087_), .ZN(new_n26416_));
  NOR2_X1    g23309(.A1(new_n26416_), .A2(pi0208), .ZN(new_n26417_));
  NOR2_X1    g23310(.A1(new_n8094_), .A2(pi1155), .ZN(new_n26418_));
  AOI21_X1   g23311(.A1(new_n26390_), .A2(new_n12026_), .B(new_n26418_), .ZN(new_n26419_));
  OAI21_X1   g23312(.A1(new_n12026_), .A2(new_n26403_), .B(new_n26419_), .ZN(new_n26420_));
  INV_X1     g23313(.I(new_n26420_), .ZN(new_n26421_));
  NOR2_X1    g23314(.A1(new_n26421_), .A2(new_n8087_), .ZN(new_n26422_));
  NOR2_X1    g23315(.A1(new_n12049_), .A2(pi0208), .ZN(new_n26423_));
  INV_X1     g23316(.I(new_n26423_), .ZN(new_n26424_));
  OAI22_X1   g23317(.A1(new_n26417_), .A2(new_n12049_), .B1(new_n26422_), .B2(new_n26424_), .ZN(new_n26425_));
  NOR2_X1    g23318(.A1(new_n26408_), .A2(new_n26425_), .ZN(new_n26426_));
  NOR2_X1    g23319(.A1(new_n8269_), .A2(pi1155), .ZN(new_n26427_));
  AOI21_X1   g23320(.A1(pi1155), .A2(new_n8626_), .B(new_n26427_), .ZN(new_n26428_));
  INV_X1     g23321(.I(new_n26428_), .ZN(new_n26429_));
  NOR2_X1    g23322(.A1(new_n26429_), .A2(new_n12026_), .ZN(new_n26430_));
  NOR2_X1    g23323(.A1(new_n26395_), .A2(pi0299), .ZN(new_n26431_));
  NOR2_X1    g23324(.A1(new_n26431_), .A2(pi1155), .ZN(new_n26432_));
  INV_X1     g23325(.I(new_n26396_), .ZN(new_n26433_));
  NOR2_X1    g23326(.A1(new_n26433_), .A2(pi0299), .ZN(new_n26434_));
  NOR2_X1    g23327(.A1(new_n26434_), .A2(new_n11912_), .ZN(new_n26435_));
  NOR2_X1    g23328(.A1(new_n26435_), .A2(new_n26432_), .ZN(new_n26436_));
  NOR2_X1    g23329(.A1(new_n26436_), .A2(new_n11950_), .ZN(new_n26437_));
  NOR2_X1    g23330(.A1(new_n26437_), .A2(new_n26430_), .ZN(new_n26438_));
  INV_X1     g23331(.I(new_n26438_), .ZN(new_n26439_));
  OAI21_X1   g23332(.A1(new_n2587_), .A2(pi1142), .B(new_n26439_), .ZN(new_n26440_));
  INV_X1     g23333(.I(new_n26383_), .ZN(new_n26441_));
  NAND2_X1   g23334(.A1(pi0299), .A2(pi1142), .ZN(new_n26442_));
  NAND2_X1   g23335(.A1(new_n26441_), .A2(new_n26442_), .ZN(new_n26443_));
  NOR2_X1    g23336(.A1(pi1154), .A2(pi1156), .ZN(new_n26444_));
  AOI21_X1   g23337(.A1(new_n26443_), .A2(new_n26444_), .B(pi0207), .ZN(new_n26445_));
  NAND3_X1   g23338(.A1(new_n3700_), .A2(pi0207), .A3(pi0299), .ZN(new_n26446_));
  NAND2_X1   g23339(.A1(new_n26446_), .A2(pi0208), .ZN(new_n26447_));
  AOI21_X1   g23340(.A1(new_n26440_), .A2(new_n26445_), .B(new_n26447_), .ZN(new_n26448_));
  NOR2_X1    g23341(.A1(new_n26394_), .A2(pi0299), .ZN(new_n26449_));
  INV_X1     g23342(.I(new_n26449_), .ZN(new_n26450_));
  AOI21_X1   g23343(.A1(new_n26450_), .A2(new_n26409_), .B(new_n26410_), .ZN(new_n26451_));
  NAND2_X1   g23344(.A1(new_n26451_), .A2(pi0207), .ZN(new_n26452_));
  AOI21_X1   g23345(.A1(new_n26452_), .A2(new_n2587_), .B(pi0208), .ZN(new_n26453_));
  NOR2_X1    g23346(.A1(new_n26453_), .A2(pi1157), .ZN(new_n26454_));
  NOR2_X1    g23347(.A1(pi0207), .A2(pi0299), .ZN(new_n26455_));
  NOR2_X1    g23348(.A1(new_n26455_), .A2(pi0208), .ZN(new_n26456_));
  INV_X1     g23349(.I(new_n26456_), .ZN(new_n26457_));
  AOI21_X1   g23350(.A1(pi1155), .A2(new_n26379_), .B(new_n26427_), .ZN(new_n26458_));
  INV_X1     g23351(.I(new_n26458_), .ZN(new_n26459_));
  INV_X1     g23352(.I(new_n8626_), .ZN(new_n26460_));
  NOR3_X1    g23353(.A1(new_n26460_), .A2(new_n12026_), .A3(new_n26399_), .ZN(new_n26461_));
  AOI21_X1   g23354(.A1(new_n26459_), .A2(new_n12026_), .B(new_n26461_), .ZN(new_n26462_));
  INV_X1     g23355(.I(new_n26462_), .ZN(new_n26463_));
  AOI21_X1   g23356(.A1(new_n26463_), .A2(pi0207), .B(new_n26457_), .ZN(new_n26464_));
  NOR2_X1    g23357(.A1(new_n26464_), .A2(new_n12049_), .ZN(new_n26465_));
  INV_X1     g23358(.I(new_n26465_), .ZN(new_n26466_));
  NOR2_X1    g23359(.A1(new_n2587_), .A2(pi1142), .ZN(new_n26467_));
  NOR4_X1    g23360(.A1(po1038), .A2(new_n8082_), .A3(new_n26376_), .A4(new_n26467_), .ZN(new_n26468_));
  NAND2_X1   g23361(.A1(new_n26466_), .A2(new_n26468_), .ZN(new_n26469_));
  NOR3_X1    g23362(.A1(new_n26448_), .A2(new_n26469_), .A3(new_n26454_), .ZN(new_n26470_));
  OAI21_X1   g23363(.A1(new_n26426_), .A2(new_n26376_), .B(new_n26470_), .ZN(new_n26471_));
  NOR2_X1    g23364(.A1(new_n8076_), .A2(pi0214), .ZN(new_n26472_));
  NOR2_X1    g23365(.A1(new_n26361_), .A2(new_n26472_), .ZN(new_n26473_));
  INV_X1     g23366(.I(new_n26406_), .ZN(new_n26474_));
  NAND2_X1   g23367(.A1(new_n26474_), .A2(pi0207), .ZN(new_n26475_));
  NOR2_X1    g23368(.A1(new_n2587_), .A2(new_n2552_), .ZN(new_n26476_));
  NOR2_X1    g23369(.A1(new_n26475_), .A2(new_n26476_), .ZN(new_n26477_));
  NOR2_X1    g23370(.A1(new_n2587_), .A2(pi1144), .ZN(new_n26478_));
  INV_X1     g23371(.I(new_n26478_), .ZN(new_n26479_));
  INV_X1     g23372(.I(new_n26476_), .ZN(new_n26480_));
  OAI21_X1   g23373(.A1(new_n26480_), .A2(pi1156), .B(new_n11950_), .ZN(new_n26482_));
  AOI21_X1   g23374(.A1(new_n26428_), .A2(new_n26479_), .B(new_n26482_), .ZN(new_n26483_));
  NOR3_X1    g23375(.A1(new_n8626_), .A2(pi1154), .A3(new_n26413_), .ZN(new_n26484_));
  INV_X1     g23376(.I(new_n26484_), .ZN(new_n26485_));
  NOR2_X1    g23377(.A1(pi1155), .A2(pi1156), .ZN(new_n26486_));
  NAND4_X1   g23378(.A1(new_n26384_), .A2(new_n26476_), .A3(new_n26485_), .A4(new_n26486_), .ZN(new_n26487_));
  AOI21_X1   g23379(.A1(new_n26435_), .A2(new_n26479_), .B(new_n26487_), .ZN(new_n26488_));
  NOR2_X1    g23380(.A1(pi0207), .A2(pi0208), .ZN(new_n26489_));
  OAI21_X1   g23381(.A1(new_n26488_), .A2(new_n26483_), .B(new_n26489_), .ZN(new_n26490_));
  NOR2_X1    g23382(.A1(new_n26478_), .A2(pi1157), .ZN(new_n26491_));
  INV_X1     g23383(.I(new_n26328_), .ZN(new_n26492_));
  INV_X1     g23384(.I(new_n26403_), .ZN(new_n26493_));
  NOR4_X1    g23385(.A1(new_n26459_), .A2(new_n12026_), .A3(new_n26493_), .A4(new_n26418_), .ZN(new_n26494_));
  NOR2_X1    g23386(.A1(new_n26494_), .A2(new_n26492_), .ZN(new_n26495_));
  NAND2_X1   g23387(.A1(new_n26495_), .A2(new_n26480_), .ZN(new_n26496_));
  NOR2_X1    g23388(.A1(new_n26495_), .A2(new_n26480_), .ZN(new_n26497_));
  NOR2_X1    g23389(.A1(new_n26497_), .A2(new_n26424_), .ZN(new_n26498_));
  AOI22_X1   g23390(.A1(new_n26498_), .A2(new_n26496_), .B1(new_n26453_), .B2(new_n26491_), .ZN(new_n26499_));
  OAI21_X1   g23391(.A1(new_n26477_), .A2(new_n26490_), .B(new_n26499_), .ZN(new_n26500_));
  AOI21_X1   g23392(.A1(new_n26500_), .A2(new_n8077_), .B(new_n26473_), .ZN(new_n26501_));
  NOR2_X1    g23393(.A1(new_n2587_), .A2(new_n3548_), .ZN(new_n26502_));
  NOR2_X1    g23394(.A1(new_n26475_), .A2(new_n26502_), .ZN(new_n26503_));
  INV_X1     g23395(.I(new_n26489_), .ZN(new_n26504_));
  NOR2_X1    g23396(.A1(new_n2587_), .A2(pi1143), .ZN(new_n26505_));
  OAI21_X1   g23397(.A1(new_n26429_), .A2(new_n26505_), .B(new_n11950_), .ZN(new_n26506_));
  NOR4_X1    g23398(.A1(new_n2587_), .A2(new_n3548_), .A3(pi1154), .A4(pi1156), .ZN(new_n26507_));
  NAND3_X1   g23399(.A1(new_n3548_), .A2(new_n11912_), .A3(pi0299), .ZN(new_n26508_));
  INV_X1     g23400(.I(new_n26502_), .ZN(new_n26509_));
  OAI21_X1   g23401(.A1(new_n26384_), .A2(new_n26509_), .B(new_n12026_), .ZN(new_n26510_));
  AOI22_X1   g23402(.A1(new_n26506_), .A2(new_n26507_), .B1(new_n26508_), .B2(new_n26510_), .ZN(new_n26511_));
  OR2_X2     g23403(.A1(new_n26511_), .A2(new_n26504_), .Z(new_n26512_));
  INV_X1     g23404(.I(new_n26505_), .ZN(new_n26513_));
  NOR3_X1    g23405(.A1(new_n26453_), .A2(pi1157), .A3(new_n26513_), .ZN(new_n26514_));
  XOR2_X1    g23406(.A1(new_n26495_), .A2(new_n26502_), .Z(new_n26515_));
  AOI21_X1   g23407(.A1(new_n26515_), .A2(new_n26424_), .B(new_n26514_), .ZN(new_n26516_));
  OAI21_X1   g23408(.A1(new_n26503_), .A2(new_n26512_), .B(new_n26516_), .ZN(new_n26517_));
  NAND3_X1   g23409(.A1(new_n26517_), .A2(new_n8077_), .A3(new_n8250_), .ZN(new_n26518_));
  OAI21_X1   g23410(.A1(new_n26518_), .A2(new_n26501_), .B(new_n8247_), .ZN(new_n26519_));
  AOI21_X1   g23411(.A1(new_n26519_), .A2(new_n26471_), .B(new_n26318_), .ZN(new_n26520_));
  OAI21_X1   g23412(.A1(new_n26520_), .A2(pi0213), .B(new_n26374_), .ZN(new_n26521_));
  NOR2_X1    g23413(.A1(new_n26449_), .A2(new_n11912_), .ZN(new_n26522_));
  NOR2_X1    g23414(.A1(new_n2587_), .A2(pi1155), .ZN(new_n26523_));
  NOR2_X1    g23415(.A1(new_n26522_), .A2(new_n26523_), .ZN(new_n26524_));
  INV_X1     g23416(.I(new_n26524_), .ZN(new_n26525_));
  NOR2_X1    g23417(.A1(new_n26439_), .A2(new_n26525_), .ZN(new_n26526_));
  INV_X1     g23418(.I(new_n26526_), .ZN(new_n26527_));
  NOR2_X1    g23419(.A1(new_n2587_), .A2(pi1153), .ZN(new_n26528_));
  INV_X1     g23420(.I(new_n26528_), .ZN(new_n26529_));
  AOI21_X1   g23421(.A1(new_n26527_), .A2(new_n26529_), .B(pi0207), .ZN(new_n26530_));
  OAI21_X1   g23422(.A1(new_n11893_), .A2(new_n26431_), .B(new_n26401_), .ZN(new_n26531_));
  NOR2_X1    g23423(.A1(new_n26531_), .A2(new_n8087_), .ZN(new_n26532_));
  NOR3_X1    g23424(.A1(new_n26530_), .A2(new_n8088_), .A3(new_n26532_), .ZN(new_n26533_));
  NOR2_X1    g23425(.A1(new_n8078_), .A2(pi0211), .ZN(new_n26534_));
  NAND2_X1   g23426(.A1(new_n26466_), .A2(new_n26529_), .ZN(new_n26535_));
  OAI21_X1   g23427(.A1(new_n26535_), .A2(new_n26454_), .B(new_n26534_), .ZN(new_n26536_));
  NOR2_X1    g23428(.A1(new_n26533_), .A2(new_n26536_), .ZN(new_n26537_));
  NOR2_X1    g23429(.A1(new_n26416_), .A2(new_n26356_), .ZN(new_n26538_));
  NOR2_X1    g23430(.A1(new_n26538_), .A2(pi0208), .ZN(new_n26539_));
  NAND2_X1   g23431(.A1(new_n26539_), .A2(new_n12049_), .ZN(new_n26540_));
  INV_X1     g23432(.I(new_n26393_), .ZN(new_n26541_));
  NOR2_X1    g23433(.A1(new_n26412_), .A2(new_n26391_), .ZN(new_n26542_));
  INV_X1     g23434(.I(new_n26542_), .ZN(new_n26543_));
  NOR2_X1    g23435(.A1(new_n8626_), .A2(new_n11912_), .ZN(new_n26544_));
  INV_X1     g23436(.I(new_n26544_), .ZN(new_n26545_));
  NAND4_X1   g23437(.A1(new_n26543_), .A2(new_n2587_), .A3(new_n11950_), .A4(new_n26545_), .ZN(new_n26546_));
  AOI21_X1   g23438(.A1(new_n26546_), .A2(new_n26541_), .B(new_n8087_), .ZN(new_n26547_));
  INV_X1     g23439(.I(new_n26547_), .ZN(new_n26548_));
  NOR2_X1    g23440(.A1(new_n8087_), .A2(pi0208), .ZN(new_n26549_));
  NOR2_X1    g23441(.A1(new_n26437_), .A2(new_n26388_), .ZN(new_n26550_));
  INV_X1     g23442(.I(new_n26550_), .ZN(new_n26551_));
  NAND3_X1   g23443(.A1(new_n26548_), .A2(new_n26551_), .A3(new_n26549_), .ZN(new_n26552_));
  NOR2_X1    g23444(.A1(new_n2587_), .A2(pi1154), .ZN(new_n26553_));
  INV_X1     g23445(.I(new_n26553_), .ZN(new_n26554_));
  NAND3_X1   g23446(.A1(new_n26464_), .A2(pi1157), .A3(new_n26554_), .ZN(new_n26555_));
  AND3_X2    g23447(.A1(new_n26552_), .A2(new_n26540_), .A3(new_n26555_), .Z(new_n26556_));
  NOR2_X1    g23448(.A1(pi0211), .A2(pi0214), .ZN(new_n26557_));
  INV_X1     g23449(.I(new_n26557_), .ZN(new_n26558_));
  NOR4_X1    g23450(.A1(new_n26537_), .A2(new_n26556_), .A3(pi0212), .A4(new_n26558_), .ZN(new_n26559_));
  NAND2_X1   g23451(.A1(new_n26426_), .A2(new_n8078_), .ZN(new_n26560_));
  NAND2_X1   g23452(.A1(new_n26560_), .A2(new_n8076_), .ZN(new_n26561_));
  AOI21_X1   g23453(.A1(new_n26364_), .A2(new_n8087_), .B(pi0208), .ZN(new_n26562_));
  INV_X1     g23454(.I(new_n26562_), .ZN(new_n26563_));
  NAND2_X1   g23455(.A1(new_n26380_), .A2(pi1155), .ZN(new_n26564_));
  NOR2_X1    g23456(.A1(new_n8169_), .A2(new_n12026_), .ZN(new_n26565_));
  OAI21_X1   g23457(.A1(new_n26431_), .A2(pi1155), .B(new_n26380_), .ZN(new_n26566_));
  AOI22_X1   g23458(.A1(new_n26566_), .A2(new_n12026_), .B1(new_n26564_), .B2(new_n26565_), .ZN(new_n26567_));
  NOR2_X1    g23459(.A1(new_n26563_), .A2(new_n12049_), .ZN(new_n26568_));
  OAI21_X1   g23460(.A1(new_n26567_), .A2(new_n8087_), .B(new_n26568_), .ZN(new_n26569_));
  NOR2_X1    g23461(.A1(new_n8169_), .A2(pi1155), .ZN(new_n26570_));
  INV_X1     g23462(.I(new_n26410_), .ZN(new_n26571_));
  NAND2_X1   g23463(.A1(new_n26571_), .A2(new_n26433_), .ZN(new_n26572_));
  AOI21_X1   g23464(.A1(new_n26572_), .A2(new_n2587_), .B(new_n26570_), .ZN(new_n26573_));
  INV_X1     g23465(.I(new_n26573_), .ZN(new_n26574_));
  OAI21_X1   g23466(.A1(new_n26563_), .A2(new_n26574_), .B(new_n26569_), .ZN(new_n26575_));
  AOI21_X1   g23467(.A1(new_n26534_), .A2(new_n26575_), .B(new_n26561_), .ZN(new_n26576_));
  AOI21_X1   g23468(.A1(new_n26426_), .A2(pi0211), .B(pi0219), .ZN(new_n26577_));
  OAI21_X1   g23469(.A1(new_n26576_), .A2(new_n26559_), .B(new_n26577_), .ZN(new_n26578_));
  OAI21_X1   g23470(.A1(new_n26408_), .A2(new_n26417_), .B(new_n12049_), .ZN(new_n26579_));
  NOR2_X1    g23471(.A1(new_n26527_), .A2(pi0207), .ZN(new_n26580_));
  NOR2_X1    g23472(.A1(new_n26531_), .A2(new_n26492_), .ZN(new_n26581_));
  NOR4_X1    g23473(.A1(new_n26580_), .A2(new_n8088_), .A3(new_n26465_), .A4(new_n26581_), .ZN(new_n26582_));
  NOR2_X1    g23474(.A1(new_n26430_), .A2(new_n26387_), .ZN(new_n26583_));
  NOR4_X1    g23475(.A1(new_n8087_), .A2(new_n2587_), .A3(new_n12026_), .A4(pi0208), .ZN(new_n26584_));
  NOR2_X1    g23476(.A1(new_n2587_), .A2(new_n12026_), .ZN(new_n26585_));
  OAI21_X1   g23477(.A1(new_n26422_), .A2(new_n26585_), .B(new_n26423_), .ZN(new_n26586_));
  NAND2_X1   g23478(.A1(new_n26453_), .A2(new_n26571_), .ZN(new_n26587_));
  NAND2_X1   g23479(.A1(new_n26587_), .A2(new_n26586_), .ZN(new_n26588_));
  AOI21_X1   g23480(.A1(new_n26406_), .A2(new_n26584_), .B(new_n26588_), .ZN(new_n26589_));
  NOR3_X1    g23481(.A1(new_n26582_), .A2(new_n26558_), .A3(new_n26589_), .ZN(new_n26590_));
  NAND3_X1   g23482(.A1(new_n26561_), .A2(new_n26579_), .A3(new_n26590_), .ZN(new_n26591_));
  NAND2_X1   g23483(.A1(new_n26589_), .A2(new_n8077_), .ZN(new_n26592_));
  XNOR2_X1   g23484(.A1(new_n26592_), .A2(new_n26575_), .ZN(new_n26593_));
  OAI22_X1   g23485(.A1(new_n26593_), .A2(pi0214), .B1(pi0211), .B2(new_n26575_), .ZN(new_n26594_));
  INV_X1     g23486(.I(new_n26556_), .ZN(new_n26595_));
  NOR4_X1    g23487(.A1(new_n26589_), .A2(pi0211), .A3(pi0214), .A4(new_n26575_), .ZN(new_n26596_));
  NAND2_X1   g23488(.A1(new_n8079_), .A2(new_n8076_), .ZN(new_n26597_));
  NOR3_X1    g23489(.A1(new_n26595_), .A2(new_n26596_), .A3(new_n26597_), .ZN(new_n26598_));
  NAND2_X1   g23490(.A1(new_n26594_), .A2(new_n26598_), .ZN(new_n26599_));
  NOR3_X1    g23491(.A1(po1038), .A2(new_n24753_), .A3(pi0219), .ZN(new_n26600_));
  NAND4_X1   g23492(.A1(new_n26578_), .A2(new_n26599_), .A3(new_n26591_), .A4(new_n26600_), .ZN(new_n26601_));
  AOI22_X1   g23493(.A1(new_n26601_), .A2(new_n26521_), .B1(new_n26354_), .B2(new_n26373_), .ZN(new_n26602_));
  MUX2_X1    g23494(.I0(new_n26602_), .I1(pi0233), .S(new_n26307_), .Z(po0390));
  INV_X1     g23495(.I(pi1152), .ZN(new_n26604_));
  NOR2_X1    g23496(.A1(new_n8161_), .A2(pi0299), .ZN(new_n26605_));
  INV_X1     g23497(.I(new_n26605_), .ZN(new_n26606_));
  OAI21_X1   g23498(.A1(new_n26606_), .A2(new_n26403_), .B(pi1153), .ZN(new_n26607_));
  NOR2_X1    g23499(.A1(new_n26607_), .A2(new_n11950_), .ZN(new_n26608_));
  NOR2_X1    g23500(.A1(pi0199), .A2(pi1153), .ZN(new_n26609_));
  NOR2_X1    g23501(.A1(new_n26412_), .A2(new_n26609_), .ZN(new_n26610_));
  NOR2_X1    g23502(.A1(new_n26608_), .A2(new_n26610_), .ZN(new_n26611_));
  NOR2_X1    g23503(.A1(new_n26611_), .A2(new_n8087_), .ZN(new_n26612_));
  NOR2_X1    g23504(.A1(new_n8161_), .A2(pi1153), .ZN(new_n26613_));
  NOR2_X1    g23505(.A1(new_n26493_), .A2(new_n26613_), .ZN(new_n26614_));
  NAND2_X1   g23506(.A1(new_n26614_), .A2(pi0207), .ZN(new_n26615_));
  XNOR2_X1   g23507(.A1(new_n26611_), .A2(new_n26615_), .ZN(new_n26616_));
  NAND2_X1   g23508(.A1(new_n26616_), .A2(new_n8088_), .ZN(new_n26617_));
  XOR2_X1    g23509(.A1(new_n26617_), .A2(new_n26612_), .Z(new_n26618_));
  AOI21_X1   g23510(.A1(new_n26618_), .A2(new_n26319_), .B(new_n8247_), .ZN(new_n26619_));
  INV_X1     g23511(.I(new_n26618_), .ZN(new_n26620_));
  NOR3_X1    g23512(.A1(new_n26620_), .A2(pi0212), .A3(pi0214), .ZN(new_n26621_));
  INV_X1     g23513(.I(new_n26585_), .ZN(new_n26622_));
  NAND2_X1   g23514(.A1(new_n26611_), .A2(new_n26622_), .ZN(new_n26623_));
  NOR2_X1    g23515(.A1(pi0200), .A2(pi1153), .ZN(new_n26624_));
  INV_X1     g23516(.I(new_n26624_), .ZN(new_n26625_));
  AOI21_X1   g23517(.A1(new_n26625_), .A2(new_n8094_), .B(pi0299), .ZN(new_n26626_));
  NOR2_X1    g23518(.A1(new_n26626_), .A2(new_n26395_), .ZN(new_n26627_));
  NOR4_X1    g23519(.A1(new_n26627_), .A2(pi0207), .A3(new_n2587_), .A4(pi1156), .ZN(new_n26628_));
  AOI21_X1   g23520(.A1(new_n26623_), .A2(new_n8087_), .B(new_n26628_), .ZN(new_n26629_));
  NOR3_X1    g23521(.A1(new_n26612_), .A2(pi0208), .A3(new_n26585_), .ZN(new_n26630_));
  OAI21_X1   g23522(.A1(new_n26630_), .A2(pi0211), .B(new_n8088_), .ZN(new_n26631_));
  NAND3_X1   g23523(.A1(new_n8160_), .A2(new_n26455_), .A3(new_n11950_), .ZN(new_n26632_));
  XOR2_X1    g23524(.A1(new_n26632_), .A2(new_n26523_), .Z(new_n26633_));
  INV_X1     g23525(.I(new_n26549_), .ZN(new_n26634_));
  INV_X1     g23526(.I(new_n26394_), .ZN(new_n26635_));
  NOR2_X1    g23527(.A1(new_n26635_), .A2(new_n11893_), .ZN(new_n26636_));
  INV_X1     g23528(.I(new_n26636_), .ZN(new_n26637_));
  NOR2_X1    g23529(.A1(new_n26637_), .A2(pi0299), .ZN(new_n26638_));
  NOR2_X1    g23530(.A1(new_n26638_), .A2(pi1154), .ZN(new_n26639_));
  INV_X1     g23531(.I(new_n26431_), .ZN(new_n26640_));
  INV_X1     g23532(.I(new_n26391_), .ZN(new_n26641_));
  NAND3_X1   g23533(.A1(new_n26641_), .A2(pi1154), .A3(new_n26379_), .ZN(new_n26642_));
  NAND2_X1   g23534(.A1(new_n26642_), .A2(new_n26640_), .ZN(new_n26643_));
  NOR2_X1    g23535(.A1(new_n26639_), .A2(new_n26643_), .ZN(new_n26644_));
  NOR3_X1    g23536(.A1(new_n26626_), .A2(new_n8087_), .A3(new_n26395_), .ZN(new_n26645_));
  NOR3_X1    g23537(.A1(new_n26644_), .A2(new_n26634_), .A3(new_n26645_), .ZN(new_n26646_));
  NOR2_X1    g23538(.A1(new_n26644_), .A2(new_n26563_), .ZN(new_n26647_));
  NOR2_X1    g23539(.A1(new_n26646_), .A2(new_n26647_), .ZN(new_n26648_));
  NOR2_X1    g23540(.A1(new_n26648_), .A2(new_n26633_), .ZN(new_n26649_));
  INV_X1     g23541(.I(new_n26314_), .ZN(new_n26650_));
  NOR2_X1    g23542(.A1(new_n26650_), .A2(pi0219), .ZN(new_n26651_));
  INV_X1     g23543(.I(new_n26651_), .ZN(new_n26652_));
  AOI21_X1   g23544(.A1(new_n26649_), .A2(pi0211), .B(new_n26652_), .ZN(new_n26653_));
  OAI21_X1   g23545(.A1(new_n26629_), .A2(new_n26631_), .B(new_n26653_), .ZN(new_n26654_));
  NOR3_X1    g23546(.A1(new_n26621_), .A2(new_n26619_), .A3(new_n26654_), .ZN(new_n26655_));
  AOI21_X1   g23547(.A1(new_n8160_), .A2(pi1153), .B(pi0299), .ZN(new_n26656_));
  NOR2_X1    g23548(.A1(new_n26656_), .A2(new_n26523_), .ZN(new_n26657_));
  INV_X1     g23549(.I(new_n26657_), .ZN(new_n26658_));
  AOI21_X1   g23550(.A1(new_n26658_), .A2(pi0207), .B(new_n8088_), .ZN(new_n26659_));
  INV_X1     g23551(.I(new_n26659_), .ZN(new_n26660_));
  MUX2_X1    g23552(.I0(new_n26637_), .I1(new_n11912_), .S(pi0299), .Z(new_n26661_));
  NOR4_X1    g23553(.A1(new_n8268_), .A2(new_n11893_), .A3(pi1154), .A4(new_n8626_), .ZN(new_n26662_));
  INV_X1     g23554(.I(new_n26662_), .ZN(new_n26663_));
  OAI22_X1   g23555(.A1(new_n26661_), .A2(pi1154), .B1(new_n26570_), .B2(new_n26663_), .ZN(new_n26664_));
  NOR2_X1    g23556(.A1(new_n26664_), .A2(pi0207), .ZN(new_n26665_));
  NOR3_X1    g23557(.A1(new_n26664_), .A2(new_n8087_), .A3(new_n26562_), .ZN(new_n26666_));
  AOI21_X1   g23558(.A1(new_n26660_), .A2(new_n26665_), .B(new_n26666_), .ZN(new_n26667_));
  INV_X1     g23559(.I(new_n26667_), .ZN(new_n26668_));
  NOR2_X1    g23560(.A1(new_n8268_), .A2(new_n11893_), .ZN(new_n26669_));
  NOR2_X1    g23561(.A1(new_n26492_), .A2(new_n8088_), .ZN(new_n26670_));
  AOI21_X1   g23562(.A1(pi0200), .A2(new_n11893_), .B(new_n8170_), .ZN(new_n26671_));
  INV_X1     g23563(.I(new_n26671_), .ZN(new_n26672_));
  NOR2_X1    g23564(.A1(new_n26672_), .A2(new_n11950_), .ZN(new_n26673_));
  AOI21_X1   g23565(.A1(new_n26638_), .A2(new_n11950_), .B(new_n26673_), .ZN(new_n26674_));
  INV_X1     g23566(.I(new_n26674_), .ZN(new_n26675_));
  NOR2_X1    g23567(.A1(new_n8088_), .A2(pi0207), .ZN(new_n26676_));
  NOR2_X1    g23568(.A1(new_n26549_), .A2(new_n26676_), .ZN(new_n26677_));
  INV_X1     g23569(.I(new_n26677_), .ZN(new_n26678_));
  AOI22_X1   g23570(.A1(new_n26675_), .A2(new_n26678_), .B1(new_n26669_), .B2(new_n26670_), .ZN(new_n26679_));
  OAI21_X1   g23571(.A1(pi0211), .A2(new_n26585_), .B(new_n26679_), .ZN(new_n26680_));
  NAND4_X1   g23572(.A1(new_n26668_), .A2(pi0211), .A3(new_n26314_), .A4(new_n26680_), .ZN(new_n26681_));
  NOR2_X1    g23573(.A1(new_n26667_), .A2(pi0211), .ZN(new_n26682_));
  NOR2_X1    g23574(.A1(new_n26638_), .A2(new_n26662_), .ZN(new_n26683_));
  MUX2_X1    g23575(.I0(new_n26683_), .I1(new_n26357_), .S(new_n8087_), .Z(new_n26684_));
  NAND2_X1   g23576(.A1(new_n26683_), .A2(new_n8087_), .ZN(new_n26685_));
  OAI21_X1   g23577(.A1(new_n26656_), .A2(new_n26553_), .B(pi0207), .ZN(new_n26686_));
  NAND2_X1   g23578(.A1(new_n26685_), .A2(new_n26686_), .ZN(new_n26687_));
  INV_X1     g23579(.I(new_n26687_), .ZN(new_n26688_));
  MUX2_X1    g23580(.I0(new_n26688_), .I1(new_n26684_), .S(new_n8088_), .Z(new_n26689_));
  OAI21_X1   g23581(.A1(new_n26689_), .A2(new_n8077_), .B(new_n8248_), .ZN(new_n26690_));
  NAND2_X1   g23582(.A1(new_n26690_), .A2(new_n26682_), .ZN(new_n26691_));
  NAND3_X1   g23583(.A1(new_n26691_), .A2(new_n8247_), .A3(new_n26681_), .ZN(new_n26692_));
  NOR2_X1    g23584(.A1(new_n26308_), .A2(new_n8247_), .ZN(new_n26693_));
  INV_X1     g23585(.I(new_n26693_), .ZN(new_n26694_));
  NAND4_X1   g23586(.A1(new_n26689_), .A2(pi0211), .A3(new_n26679_), .A4(new_n26694_), .ZN(new_n26695_));
  NAND2_X1   g23587(.A1(new_n26679_), .A2(new_n26308_), .ZN(new_n26696_));
  AND3_X2    g23588(.A1(new_n26692_), .A2(new_n26695_), .A3(new_n26696_), .Z(new_n26697_));
  INV_X1     g23589(.I(new_n26697_), .ZN(new_n26698_));
  AOI21_X1   g23590(.A1(new_n26698_), .A2(new_n26604_), .B(new_n26655_), .ZN(new_n26699_));
  NAND3_X1   g23591(.A1(new_n26697_), .A2(new_n26655_), .A3(new_n26604_), .ZN(new_n26700_));
  INV_X1     g23592(.I(new_n26700_), .ZN(new_n26701_));
  NOR3_X1    g23593(.A1(new_n26701_), .A2(new_n26699_), .A3(po1038), .ZN(new_n26702_));
  INV_X1     g23594(.I(new_n26702_), .ZN(new_n26703_));
  INV_X1     g23595(.I(new_n26473_), .ZN(new_n26704_));
  INV_X1     g23596(.I(new_n26689_), .ZN(new_n26705_));
  NOR2_X1    g23597(.A1(new_n26358_), .A2(pi0207), .ZN(new_n26706_));
  NOR2_X1    g23598(.A1(new_n26389_), .A2(pi1153), .ZN(new_n26707_));
  NAND2_X1   g23599(.A1(new_n26460_), .A2(pi1154), .ZN(new_n26708_));
  NOR2_X1    g23600(.A1(new_n26708_), .A2(new_n26707_), .ZN(new_n26709_));
  NOR2_X1    g23601(.A1(new_n11893_), .A2(pi1154), .ZN(new_n26710_));
  INV_X1     g23602(.I(new_n26710_), .ZN(new_n26711_));
  NOR2_X1    g23603(.A1(new_n26449_), .A2(new_n26711_), .ZN(new_n26712_));
  NOR3_X1    g23604(.A1(new_n26709_), .A2(new_n8087_), .A3(new_n26712_), .ZN(new_n26713_));
  NOR2_X1    g23605(.A1(new_n26713_), .A2(new_n26706_), .ZN(new_n26714_));
  NOR2_X1    g23606(.A1(new_n26714_), .A2(pi0208), .ZN(new_n26715_));
  MUX2_X1    g23607(.I0(new_n26715_), .I1(new_n26705_), .S(new_n8077_), .Z(new_n26716_));
  NAND2_X1   g23608(.A1(new_n26716_), .A2(new_n26704_), .ZN(new_n26717_));
  AOI21_X1   g23609(.A1(new_n26715_), .A2(new_n8251_), .B(pi0219), .ZN(new_n26718_));
  INV_X1     g23610(.I(new_n26375_), .ZN(new_n26719_));
  NOR2_X1    g23611(.A1(pi0211), .A2(pi1154), .ZN(new_n26720_));
  NOR2_X1    g23612(.A1(new_n8077_), .A2(pi1153), .ZN(new_n26721_));
  NOR2_X1    g23613(.A1(new_n26721_), .A2(new_n26720_), .ZN(new_n26722_));
  INV_X1     g23614(.I(new_n26722_), .ZN(new_n26723_));
  AOI21_X1   g23615(.A1(new_n26723_), .A2(new_n8250_), .B(new_n26719_), .ZN(new_n26724_));
  INV_X1     g23616(.I(new_n26724_), .ZN(new_n26725_));
  NOR2_X1    g23617(.A1(new_n11893_), .A2(pi0211), .ZN(new_n26726_));
  INV_X1     g23618(.I(new_n26726_), .ZN(new_n26727_));
  AOI21_X1   g23619(.A1(new_n8248_), .A2(new_n26727_), .B(new_n26725_), .ZN(new_n26728_));
  AOI21_X1   g23620(.A1(new_n26728_), .A2(po1038), .B(pi1152), .ZN(new_n26729_));
  INV_X1     g23621(.I(new_n26729_), .ZN(new_n26730_));
  NOR2_X1    g23622(.A1(new_n26704_), .A2(new_n26534_), .ZN(new_n26731_));
  INV_X1     g23623(.I(new_n26731_), .ZN(new_n26732_));
  AOI21_X1   g23624(.A1(new_n8247_), .A2(new_n26732_), .B(new_n26679_), .ZN(new_n26733_));
  OAI21_X1   g23625(.A1(new_n26733_), .A2(po1038), .B(new_n26730_), .ZN(new_n26734_));
  AOI21_X1   g23626(.A1(new_n26717_), .A2(new_n26718_), .B(new_n26734_), .ZN(new_n26735_));
  NOR2_X1    g23627(.A1(pi0211), .A2(pi1153), .ZN(new_n26736_));
  INV_X1     g23628(.I(new_n26736_), .ZN(new_n26737_));
  NOR2_X1    g23629(.A1(new_n26720_), .A2(pi1153), .ZN(new_n26738_));
  NOR3_X1    g23630(.A1(new_n11893_), .A2(pi0211), .A3(pi1154), .ZN(new_n26739_));
  OAI21_X1   g23631(.A1(new_n26738_), .A2(new_n26739_), .B(new_n8078_), .ZN(new_n26740_));
  OAI21_X1   g23632(.A1(new_n26740_), .A2(new_n26737_), .B(pi0212), .ZN(new_n26741_));
  AOI21_X1   g23633(.A1(new_n26740_), .A2(new_n26737_), .B(new_n26741_), .ZN(new_n26742_));
  INV_X1     g23634(.I(new_n26311_), .ZN(new_n26743_));
  NAND2_X1   g23635(.A1(new_n26722_), .A2(new_n26361_), .ZN(new_n26744_));
  NAND4_X1   g23636(.A1(new_n26743_), .A2(new_n8247_), .A3(new_n26604_), .A4(new_n26744_), .ZN(new_n26745_));
  NOR2_X1    g23637(.A1(new_n26745_), .A2(new_n26742_), .ZN(new_n26746_));
  NAND2_X1   g23638(.A1(new_n26620_), .A2(pi0211), .ZN(new_n26747_));
  INV_X1     g23639(.I(new_n26646_), .ZN(new_n26748_));
  OAI21_X1   g23640(.A1(new_n26457_), .A2(new_n26644_), .B(new_n26748_), .ZN(new_n26749_));
  NAND2_X1   g23641(.A1(new_n26749_), .A2(new_n8077_), .ZN(new_n26750_));
  NOR3_X1    g23642(.A1(new_n26620_), .A2(pi0219), .A3(new_n26342_), .ZN(new_n26751_));
  NAND3_X1   g23643(.A1(new_n26751_), .A2(new_n26747_), .A3(new_n26750_), .ZN(new_n26752_));
  AOI21_X1   g23644(.A1(new_n26434_), .A2(new_n26708_), .B(new_n26707_), .ZN(new_n26753_));
  NOR2_X1    g23645(.A1(new_n26753_), .A2(new_n8087_), .ZN(new_n26754_));
  OAI21_X1   g23646(.A1(new_n26754_), .A2(new_n26706_), .B(new_n8088_), .ZN(new_n26755_));
  NOR2_X1    g23647(.A1(new_n8268_), .A2(pi1153), .ZN(new_n26756_));
  NOR2_X1    g23648(.A1(new_n26380_), .A2(new_n8094_), .ZN(new_n26757_));
  NOR2_X1    g23649(.A1(new_n26757_), .A2(new_n26756_), .ZN(new_n26758_));
  MUX2_X1    g23650(.I0(new_n26758_), .I1(new_n26753_), .S(new_n8087_), .Z(new_n26759_));
  OAI21_X1   g23651(.A1(new_n8088_), .A2(new_n26759_), .B(new_n26755_), .ZN(new_n26760_));
  NAND4_X1   g23652(.A1(new_n26760_), .A2(pi0211), .A3(new_n8076_), .A4(new_n8078_), .ZN(new_n26762_));
  NOR2_X1    g23653(.A1(new_n8076_), .A2(new_n8078_), .ZN(new_n26763_));
  NAND3_X1   g23654(.A1(new_n26760_), .A2(pi0211), .A3(new_n26763_), .ZN(new_n26764_));
  NAND3_X1   g23655(.A1(new_n26762_), .A2(new_n26764_), .A3(new_n8247_), .ZN(new_n26765_));
  NAND3_X1   g23656(.A1(new_n26752_), .A2(new_n6845_), .A3(new_n26765_), .ZN(new_n26766_));
  AOI21_X1   g23657(.A1(new_n26766_), .A2(new_n26746_), .B(new_n26735_), .ZN(new_n26767_));
  NAND3_X1   g23658(.A1(new_n26703_), .A2(new_n24753_), .A3(new_n26767_), .ZN(new_n26768_));
  OAI21_X1   g23659(.A1(pi0213), .A2(new_n26767_), .B(new_n26702_), .ZN(new_n26769_));
  INV_X1     g23660(.I(new_n26746_), .ZN(new_n26770_));
  NOR2_X1    g23661(.A1(new_n8087_), .A2(new_n8088_), .ZN(new_n26771_));
  AOI21_X1   g23662(.A1(new_n26399_), .A2(new_n8169_), .B(pi1154), .ZN(new_n26772_));
  NOR2_X1    g23663(.A1(new_n8161_), .A2(pi1155), .ZN(new_n26773_));
  OR2_X2     g23664(.A1(new_n26773_), .A2(new_n26402_), .Z(new_n26774_));
  AOI21_X1   g23665(.A1(new_n26774_), .A2(new_n2587_), .B(new_n26772_), .ZN(new_n26775_));
  NAND3_X1   g23666(.A1(new_n26551_), .A2(new_n8087_), .A3(new_n26775_), .ZN(new_n26776_));
  OAI21_X1   g23667(.A1(pi0207), .A2(new_n26775_), .B(new_n26550_), .ZN(new_n26777_));
  NAND2_X1   g23668(.A1(new_n26776_), .A2(new_n26777_), .ZN(new_n26778_));
  AOI22_X1   g23669(.A1(new_n26778_), .A2(new_n8088_), .B1(new_n26550_), .B2(new_n26771_), .ZN(new_n26779_));
  NAND2_X1   g23670(.A1(new_n26779_), .A2(new_n8077_), .ZN(new_n26780_));
  NOR2_X1    g23671(.A1(new_n26527_), .A2(new_n8087_), .ZN(new_n26781_));
  INV_X1     g23672(.I(new_n26781_), .ZN(new_n26782_));
  OAI21_X1   g23673(.A1(new_n26775_), .A2(new_n26492_), .B(pi0208), .ZN(new_n26783_));
  AOI22_X1   g23674(.A1(new_n26782_), .A2(new_n26456_), .B1(new_n26580_), .B2(new_n26783_), .ZN(new_n26784_));
  AOI21_X1   g23675(.A1(new_n26784_), .A2(new_n26529_), .B(new_n8077_), .ZN(new_n26785_));
  INV_X1     g23676(.I(new_n26785_), .ZN(new_n26786_));
  NAND2_X1   g23677(.A1(new_n26786_), .A2(new_n26780_), .ZN(new_n26787_));
  NOR2_X1    g23678(.A1(new_n26529_), .A2(pi0211), .ZN(new_n26788_));
  NAND3_X1   g23679(.A1(new_n26784_), .A2(new_n8078_), .A3(new_n26788_), .ZN(new_n26789_));
  OAI21_X1   g23680(.A1(new_n26787_), .A2(pi0214), .B(new_n26789_), .ZN(new_n26790_));
  NAND2_X1   g23681(.A1(new_n26388_), .A2(pi0207), .ZN(new_n26791_));
  NOR2_X1    g23682(.A1(new_n26377_), .A2(pi0199), .ZN(new_n26792_));
  XOR2_X1    g23683(.A1(new_n26792_), .A2(pi0200), .Z(new_n26793_));
  NOR4_X1    g23684(.A1(new_n26793_), .A2(new_n8087_), .A3(pi0299), .A4(new_n26772_), .ZN(new_n26794_));
  XNOR2_X1   g23685(.A1(new_n26388_), .A2(new_n26794_), .ZN(new_n26795_));
  NAND2_X1   g23686(.A1(new_n26795_), .A2(new_n8088_), .ZN(new_n26796_));
  XNOR2_X1   g23687(.A1(new_n26796_), .A2(new_n26791_), .ZN(new_n26797_));
  NAND3_X1   g23688(.A1(new_n26787_), .A2(pi0212), .A3(pi0214), .ZN(new_n26798_));
  NAND2_X1   g23689(.A1(new_n26798_), .A2(new_n8247_), .ZN(new_n26799_));
  NAND3_X1   g23690(.A1(new_n26799_), .A2(pi0212), .A3(new_n26790_), .ZN(new_n26800_));
  INV_X1     g23691(.I(new_n26797_), .ZN(new_n26801_));
  AOI21_X1   g23692(.A1(new_n26801_), .A2(new_n26319_), .B(new_n8247_), .ZN(new_n26802_));
  NAND2_X1   g23693(.A1(new_n26784_), .A2(new_n26309_), .ZN(new_n26803_));
  AOI21_X1   g23694(.A1(new_n26802_), .A2(new_n26803_), .B(po1038), .ZN(new_n26804_));
  AOI21_X1   g23695(.A1(new_n26800_), .A2(new_n26804_), .B(new_n26770_), .ZN(new_n26805_));
  NOR2_X1    g23696(.A1(new_n26787_), .A2(pi0214), .ZN(new_n26806_));
  NAND2_X1   g23697(.A1(new_n26801_), .A2(pi0211), .ZN(new_n26807_));
  AOI21_X1   g23698(.A1(new_n26786_), .A2(new_n26807_), .B(new_n8078_), .ZN(new_n26808_));
  NOR2_X1    g23699(.A1(new_n26806_), .A2(new_n26808_), .ZN(new_n26809_));
  OAI21_X1   g23700(.A1(new_n26801_), .A2(new_n8247_), .B(new_n6845_), .ZN(new_n26810_));
  NAND4_X1   g23701(.A1(new_n26799_), .A2(pi0212), .A3(new_n26730_), .A4(new_n26810_), .ZN(new_n26811_));
  OAI21_X1   g23702(.A1(new_n26319_), .A2(new_n26779_), .B(new_n26802_), .ZN(new_n26812_));
  NOR3_X1    g23703(.A1(po1038), .A2(new_n24753_), .A3(new_n8247_), .ZN(new_n26813_));
  AOI21_X1   g23704(.A1(new_n26812_), .A2(new_n26813_), .B(pi0213), .ZN(new_n26814_));
  OAI21_X1   g23705(.A1(new_n26811_), .A2(new_n26809_), .B(new_n26814_), .ZN(new_n26815_));
  OAI21_X1   g23706(.A1(new_n26815_), .A2(new_n26805_), .B(new_n26374_), .ZN(new_n26816_));
  NOR2_X1    g23707(.A1(new_n8077_), .A2(new_n11912_), .ZN(new_n26817_));
  INV_X1     g23708(.I(new_n26817_), .ZN(new_n26818_));
  NOR2_X1    g23709(.A1(new_n12026_), .A2(pi0211), .ZN(new_n26819_));
  INV_X1     g23710(.I(new_n26819_), .ZN(new_n26820_));
  AOI21_X1   g23711(.A1(new_n26818_), .A2(new_n26820_), .B(new_n8078_), .ZN(new_n26821_));
  NOR2_X1    g23712(.A1(new_n11950_), .A2(pi0211), .ZN(new_n26822_));
  NOR4_X1    g23713(.A1(new_n26821_), .A2(pi0212), .A3(new_n24753_), .A4(pi0219), .ZN(new_n26823_));
  AOI21_X1   g23714(.A1(new_n26311_), .A2(new_n26823_), .B(pi0209), .ZN(new_n26824_));
  NAND4_X1   g23715(.A1(new_n26816_), .A2(new_n26768_), .A3(new_n26769_), .A4(new_n26824_), .ZN(new_n26825_));
  MUX2_X1    g23716(.I0(new_n26825_), .I1(pi0234), .S(new_n26307_), .Z(po0391));
  INV_X1     g23717(.I(new_n26451_), .ZN(new_n26827_));
  NOR2_X1    g23718(.A1(new_n26383_), .A2(pi1156), .ZN(new_n26828_));
  NAND4_X1   g23719(.A1(new_n26429_), .A2(pi0207), .A3(pi1156), .A4(new_n26828_), .ZN(new_n26829_));
  OAI21_X1   g23720(.A1(pi0207), .A2(new_n26827_), .B(new_n26829_), .ZN(new_n26830_));
  NAND2_X1   g23721(.A1(new_n26830_), .A2(pi0208), .ZN(new_n26831_));
  AOI21_X1   g23722(.A1(new_n26831_), .A2(new_n26587_), .B(pi1157), .ZN(new_n26832_));
  INV_X1     g23723(.I(new_n26832_), .ZN(new_n26833_));
  NOR2_X1    g23724(.A1(new_n8088_), .A2(new_n12049_), .ZN(new_n26834_));
  NOR3_X1    g23725(.A1(new_n26390_), .A2(new_n26418_), .A3(pi1156), .ZN(new_n26835_));
  NOR2_X1    g23726(.A1(new_n26460_), .A2(new_n26399_), .ZN(new_n26836_));
  NOR2_X1    g23727(.A1(new_n26836_), .A2(new_n12026_), .ZN(new_n26837_));
  OAI21_X1   g23728(.A1(new_n26837_), .A2(new_n26835_), .B(new_n8087_), .ZN(new_n26838_));
  NAND2_X1   g23729(.A1(new_n26829_), .A2(new_n26838_), .ZN(new_n26839_));
  NAND2_X1   g23730(.A1(new_n26839_), .A2(new_n26834_), .ZN(new_n26840_));
  NAND3_X1   g23731(.A1(new_n26833_), .A2(new_n26586_), .A3(new_n26840_), .ZN(new_n26841_));
  NOR2_X1    g23732(.A1(new_n26522_), .A2(new_n26378_), .ZN(new_n26842_));
  NOR2_X1    g23733(.A1(new_n26842_), .A2(new_n8087_), .ZN(new_n26843_));
  NAND2_X1   g23734(.A1(new_n26567_), .A2(new_n8087_), .ZN(new_n26844_));
  INV_X1     g23735(.I(new_n26844_), .ZN(new_n26845_));
  OAI21_X1   g23736(.A1(new_n26845_), .A2(new_n26843_), .B(new_n26834_), .ZN(new_n26846_));
  NOR2_X1    g23737(.A1(new_n26574_), .A2(pi0207), .ZN(new_n26847_));
  OAI21_X1   g23738(.A1(new_n26847_), .A2(new_n26843_), .B(pi0208), .ZN(new_n26848_));
  AOI21_X1   g23739(.A1(new_n26573_), .A2(new_n26562_), .B(pi1157), .ZN(new_n26849_));
  AOI22_X1   g23740(.A1(new_n26848_), .A2(new_n26849_), .B1(new_n26846_), .B2(new_n26569_), .ZN(new_n26850_));
  INV_X1     g23741(.I(new_n26850_), .ZN(new_n26851_));
  MUX2_X1    g23742(.I0(new_n26851_), .I1(new_n26841_), .S(new_n8077_), .Z(new_n26852_));
  OR2_X2     g23743(.A1(new_n26852_), .A2(new_n8250_), .Z(new_n26853_));
  NOR4_X1    g23744(.A1(new_n26383_), .A2(new_n12026_), .A3(new_n8089_), .A4(new_n26378_), .ZN(new_n26854_));
  INV_X1     g23745(.I(new_n26854_), .ZN(new_n26855_));
  NOR3_X1    g23746(.A1(new_n26415_), .A2(pi0207), .A3(new_n8088_), .ZN(new_n26856_));
  AOI21_X1   g23747(.A1(new_n26415_), .A2(new_n8088_), .B(new_n8087_), .ZN(new_n26857_));
  OAI21_X1   g23748(.A1(new_n26856_), .A2(new_n26857_), .B(new_n26855_), .ZN(new_n26858_));
  OAI21_X1   g23749(.A1(new_n8090_), .A2(new_n26421_), .B(new_n26855_), .ZN(new_n26859_));
  NAND3_X1   g23750(.A1(new_n26859_), .A2(pi1157), .A3(new_n26489_), .ZN(new_n26860_));
  OAI21_X1   g23751(.A1(new_n26858_), .A2(pi1157), .B(new_n26860_), .ZN(new_n26861_));
  NOR2_X1    g23752(.A1(new_n26861_), .A2(new_n26342_), .ZN(new_n26862_));
  AOI21_X1   g23753(.A1(new_n26858_), .A2(new_n12049_), .B(pi0211), .ZN(new_n26863_));
  AOI21_X1   g23754(.A1(new_n26463_), .A2(new_n8087_), .B(new_n8088_), .ZN(new_n26864_));
  NOR4_X1    g23755(.A1(new_n26864_), .A2(new_n8087_), .A3(new_n26430_), .A4(new_n26525_), .ZN(new_n26865_));
  NOR2_X1    g23756(.A1(new_n26865_), .A2(new_n26464_), .ZN(new_n26866_));
  INV_X1     g23757(.I(new_n26866_), .ZN(new_n26867_));
  OR3_X2     g23758(.A1(new_n26867_), .A2(new_n12049_), .A3(new_n26863_), .Z(new_n26868_));
  NOR3_X1    g23759(.A1(new_n26841_), .A2(pi0211), .A3(new_n26704_), .ZN(new_n26869_));
  AOI21_X1   g23760(.A1(new_n26868_), .A2(new_n26869_), .B(new_n26862_), .ZN(new_n26870_));
  AOI21_X1   g23761(.A1(new_n26853_), .A2(new_n26870_), .B(pi0219), .ZN(new_n26871_));
  NOR2_X1    g23762(.A1(new_n26861_), .A2(new_n8077_), .ZN(new_n26872_));
  NOR2_X1    g23763(.A1(new_n26872_), .A2(new_n26650_), .ZN(new_n26873_));
  AOI21_X1   g23764(.A1(new_n26861_), .A2(new_n26650_), .B(new_n8247_), .ZN(new_n26874_));
  NOR4_X1    g23765(.A1(new_n26873_), .A2(new_n26874_), .A3(pi0211), .A4(new_n26851_), .ZN(new_n26875_));
  OAI21_X1   g23766(.A1(new_n26871_), .A2(new_n26875_), .B(new_n26374_), .ZN(new_n26876_));
  NOR3_X1    g23767(.A1(new_n26531_), .A2(pi0207), .A3(pi0299), .ZN(new_n26877_));
  AOI21_X1   g23768(.A1(new_n26637_), .A2(new_n2587_), .B(pi1154), .ZN(new_n26878_));
  OAI21_X1   g23769(.A1(new_n26878_), .A2(new_n26662_), .B(new_n26549_), .ZN(new_n26879_));
  NOR2_X1    g23770(.A1(new_n26581_), .A2(new_n26457_), .ZN(new_n26880_));
  INV_X1     g23771(.I(new_n26880_), .ZN(new_n26881_));
  OAI21_X1   g23772(.A1(new_n26877_), .A2(new_n26879_), .B(new_n26881_), .ZN(new_n26882_));
  AOI21_X1   g23773(.A1(new_n26474_), .A2(new_n8090_), .B(new_n26489_), .ZN(new_n26883_));
  INV_X1     g23774(.I(new_n26883_), .ZN(new_n26884_));
  AOI21_X1   g23775(.A1(new_n8089_), .A2(new_n26674_), .B(new_n26884_), .ZN(new_n26885_));
  INV_X1     g23776(.I(new_n26885_), .ZN(new_n26886_));
  NOR3_X1    g23777(.A1(new_n26886_), .A2(pi1157), .A3(new_n26882_), .ZN(new_n26887_));
  OAI21_X1   g23778(.A1(new_n26885_), .A2(pi1157), .B(new_n26882_), .ZN(new_n26888_));
  NOR2_X1    g23779(.A1(new_n26885_), .A2(new_n26585_), .ZN(new_n26889_));
  NAND2_X1   g23780(.A1(new_n26888_), .A2(new_n8077_), .ZN(new_n26890_));
  OAI21_X1   g23781(.A1(new_n26890_), .A2(new_n26887_), .B(new_n26704_), .ZN(new_n26891_));
  OAI21_X1   g23782(.A1(new_n26886_), .A2(new_n26314_), .B(pi0219), .ZN(new_n26892_));
  AOI21_X1   g23783(.A1(new_n26886_), .A2(pi0211), .B(new_n26650_), .ZN(new_n26893_));
  OAI21_X1   g23784(.A1(new_n26664_), .A2(new_n8087_), .B(pi0208), .ZN(new_n26894_));
  INV_X1     g23785(.I(new_n26894_), .ZN(new_n26895_));
  NOR2_X1    g23786(.A1(new_n26894_), .A2(new_n8087_), .ZN(new_n26896_));
  NOR3_X1    g23787(.A1(new_n26896_), .A2(new_n26895_), .A3(new_n26562_), .ZN(new_n26897_));
  NOR3_X1    g23788(.A1(new_n26893_), .A2(pi0211), .A3(new_n26897_), .ZN(new_n26898_));
  AOI21_X1   g23789(.A1(new_n26898_), .A2(new_n26892_), .B(pi0209), .ZN(new_n26899_));
  AOI21_X1   g23790(.A1(new_n26885_), .A2(new_n26342_), .B(pi0219), .ZN(new_n26900_));
  INV_X1     g23791(.I(new_n26889_), .ZN(new_n26901_));
  INV_X1     g23792(.I(new_n26897_), .ZN(new_n26902_));
  OAI21_X1   g23793(.A1(new_n26901_), .A2(new_n26902_), .B(pi0211), .ZN(new_n26903_));
  OAI21_X1   g23794(.A1(new_n26903_), .A2(new_n8250_), .B(new_n26900_), .ZN(new_n26904_));
  NOR2_X1    g23795(.A1(new_n26899_), .A2(new_n26904_), .ZN(new_n26905_));
  AOI21_X1   g23796(.A1(new_n26905_), .A2(new_n26891_), .B(po1038), .ZN(new_n26906_));
  NOR2_X1    g23797(.A1(new_n26368_), .A2(pi0214), .ZN(new_n26907_));
  OAI21_X1   g23798(.A1(new_n26907_), .A2(new_n26821_), .B(pi0212), .ZN(new_n26908_));
  NAND2_X1   g23799(.A1(new_n26908_), .A2(new_n8247_), .ZN(new_n26909_));
  NOR2_X1    g23800(.A1(new_n11912_), .A2(pi0211), .ZN(new_n26910_));
  INV_X1     g23801(.I(new_n26910_), .ZN(new_n26911_));
  NOR4_X1    g23802(.A1(po1038), .A2(pi0219), .A3(new_n26473_), .A4(new_n26911_), .ZN(new_n26912_));
  OR3_X2     g23803(.A1(new_n26912_), .A2(new_n26362_), .A3(new_n26368_), .Z(new_n26913_));
  OAI21_X1   g23804(.A1(new_n26913_), .A2(new_n26909_), .B(pi0213), .ZN(new_n26914_));
  AOI21_X1   g23805(.A1(new_n26906_), .A2(new_n26876_), .B(new_n26914_), .ZN(new_n26915_));
  INV_X1     g23806(.I(new_n26874_), .ZN(new_n26916_));
  NAND3_X1   g23807(.A1(new_n26866_), .A2(pi0299), .A3(new_n12049_), .ZN(new_n26917_));
  OAI21_X1   g23808(.A1(pi0299), .A2(pi1157), .B(new_n26867_), .ZN(new_n26918_));
  NAND4_X1   g23809(.A1(new_n26918_), .A2(new_n26529_), .A3(new_n26833_), .A4(new_n26917_), .ZN(new_n26919_));
  NAND2_X1   g23810(.A1(new_n26919_), .A2(new_n8077_), .ZN(new_n26920_));
  NAND3_X1   g23811(.A1(new_n26920_), .A2(new_n26873_), .A3(new_n26916_), .ZN(new_n26921_));
  NOR2_X1    g23812(.A1(new_n26412_), .A2(new_n26413_), .ZN(new_n26922_));
  NOR2_X1    g23813(.A1(new_n26571_), .A2(pi0299), .ZN(new_n26923_));
  NOR4_X1    g23814(.A1(new_n26450_), .A2(pi1154), .A3(new_n12026_), .A4(new_n26409_), .ZN(new_n26924_));
  NOR4_X1    g23815(.A1(new_n26922_), .A2(pi0207), .A3(new_n26923_), .A4(new_n26924_), .ZN(new_n26925_));
  NOR2_X1    g23816(.A1(new_n26378_), .A2(pi0207), .ZN(new_n26926_));
  OAI21_X1   g23817(.A1(new_n26524_), .A2(new_n26384_), .B(new_n26926_), .ZN(new_n26927_));
  AOI21_X1   g23818(.A1(new_n26925_), .A2(new_n26927_), .B(new_n8088_), .ZN(new_n26928_));
  NOR2_X1    g23819(.A1(new_n26539_), .A2(new_n26928_), .ZN(new_n26929_));
  NOR2_X1    g23820(.A1(new_n26866_), .A2(new_n26553_), .ZN(new_n26930_));
  MUX2_X1    g23821(.I0(new_n26930_), .I1(new_n26929_), .S(new_n12049_), .Z(new_n26931_));
  OAI21_X1   g23822(.A1(new_n26850_), .A2(pi0211), .B(new_n26704_), .ZN(new_n26932_));
  AOI21_X1   g23823(.A1(new_n26931_), .A2(pi0211), .B(new_n26932_), .ZN(new_n26933_));
  OAI21_X1   g23824(.A1(new_n26933_), .A2(new_n26862_), .B(new_n8247_), .ZN(new_n26934_));
  AOI21_X1   g23825(.A1(new_n26921_), .A2(new_n26934_), .B(new_n26374_), .ZN(new_n26935_));
  NOR2_X1    g23826(.A1(new_n26706_), .A2(pi0208), .ZN(new_n26936_));
  INV_X1     g23827(.I(new_n26936_), .ZN(new_n26937_));
  NOR2_X1    g23828(.A1(new_n26713_), .A2(new_n26634_), .ZN(new_n26938_));
  AOI22_X1   g23829(.A1(new_n26532_), .A2(new_n26937_), .B1(new_n26531_), .B2(new_n26938_), .ZN(new_n26939_));
  NAND2_X1   g23830(.A1(new_n26939_), .A2(new_n8077_), .ZN(new_n26940_));
  AOI21_X1   g23831(.A1(new_n26893_), .A2(new_n26940_), .B(new_n26892_), .ZN(new_n26941_));
  INV_X1     g23832(.I(new_n26900_), .ZN(new_n26942_));
  AOI21_X1   g23833(.A1(new_n26357_), .A2(new_n8087_), .B(pi0208), .ZN(new_n26943_));
  NOR2_X1    g23834(.A1(new_n26548_), .A2(new_n26943_), .ZN(new_n26944_));
  NAND2_X1   g23835(.A1(new_n26546_), .A2(new_n26541_), .ZN(new_n26945_));
  NOR2_X1    g23836(.A1(new_n26945_), .A2(pi0207), .ZN(new_n26946_));
  NOR2_X1    g23837(.A1(new_n26683_), .A2(new_n8087_), .ZN(new_n26947_));
  NOR2_X1    g23838(.A1(new_n26946_), .A2(new_n26947_), .ZN(new_n26948_));
  NAND2_X1   g23839(.A1(new_n26946_), .A2(new_n26947_), .ZN(new_n26949_));
  NAND2_X1   g23840(.A1(new_n26949_), .A2(pi0208), .ZN(new_n26950_));
  NOR2_X1    g23841(.A1(new_n26950_), .A2(new_n26948_), .ZN(new_n26951_));
  OAI21_X1   g23842(.A1(new_n26951_), .A2(new_n26944_), .B(pi0211), .ZN(new_n26952_));
  NAND2_X1   g23843(.A1(new_n26939_), .A2(pi0211), .ZN(new_n26953_));
  AOI21_X1   g23844(.A1(new_n26952_), .A2(new_n26953_), .B(new_n8250_), .ZN(new_n26954_));
  NAND2_X1   g23845(.A1(new_n26952_), .A2(new_n26314_), .ZN(new_n26955_));
  AOI21_X1   g23846(.A1(new_n8077_), .A2(new_n26897_), .B(new_n26955_), .ZN(new_n26956_));
  NOR3_X1    g23847(.A1(new_n26956_), .A2(new_n26942_), .A3(new_n26954_), .ZN(new_n26957_));
  OAI21_X1   g23848(.A1(new_n26957_), .A2(new_n26941_), .B(new_n26374_), .ZN(new_n26958_));
  NAND2_X1   g23849(.A1(new_n26958_), .A2(new_n6845_), .ZN(new_n26959_));
  NAND2_X1   g23850(.A1(new_n26727_), .A2(pi0219), .ZN(new_n26960_));
  NAND2_X1   g23851(.A1(po1038), .A2(new_n26960_), .ZN(new_n26961_));
  INV_X1     g23852(.I(new_n26961_), .ZN(new_n26962_));
  NOR2_X1    g23853(.A1(new_n8077_), .A2(new_n11950_), .ZN(new_n26963_));
  NOR2_X1    g23854(.A1(new_n26963_), .A2(new_n26910_), .ZN(new_n26964_));
  NOR2_X1    g23855(.A1(new_n26473_), .A2(new_n26964_), .ZN(new_n26965_));
  NOR2_X1    g23856(.A1(new_n26723_), .A2(new_n8250_), .ZN(new_n26966_));
  NOR3_X1    g23857(.A1(new_n26966_), .A2(pi0219), .A3(new_n26965_), .ZN(new_n26967_));
  AOI21_X1   g23858(.A1(pi0219), .A2(new_n26473_), .B(new_n26967_), .ZN(new_n26968_));
  AOI21_X1   g23859(.A1(new_n26962_), .A2(new_n26968_), .B(pi0213), .ZN(new_n26969_));
  OAI21_X1   g23860(.A1(new_n26959_), .A2(new_n26935_), .B(new_n26969_), .ZN(new_n26970_));
  NOR2_X1    g23861(.A1(new_n26915_), .A2(new_n26970_), .ZN(new_n26971_));
  MUX2_X1    g23862(.I0(new_n26971_), .I1(pi0235), .S(new_n26307_), .Z(po0392));
  NAND2_X1   g23863(.A1(new_n26165_), .A2(new_n3173_), .ZN(new_n26973_));
  NOR3_X1    g23864(.A1(new_n5191_), .A2(pi0087), .A3(new_n5160_), .ZN(new_n26974_));
  AOI21_X1   g23865(.A1(new_n26973_), .A2(new_n26974_), .B(pi0075), .ZN(new_n26975_));
  NOR2_X1    g23866(.A1(new_n3214_), .A2(pi0092), .ZN(new_n26976_));
  OAI21_X1   g23867(.A1(new_n26975_), .A2(new_n5876_), .B(new_n26976_), .ZN(new_n26977_));
  AOI21_X1   g23868(.A1(new_n26977_), .A2(new_n5200_), .B(pi0056), .ZN(new_n26978_));
  OAI21_X1   g23869(.A1(new_n26978_), .A2(new_n5057_), .B(new_n5203_), .ZN(po0393));
  NOR2_X1    g23870(.A1(pi0211), .A2(pi1145), .ZN(new_n26980_));
  AOI21_X1   g23871(.A1(pi0211), .A2(new_n2552_), .B(new_n26980_), .ZN(new_n26981_));
  NOR3_X1    g23872(.A1(new_n26347_), .A2(new_n8076_), .A3(new_n8078_), .ZN(new_n26982_));
  AOI21_X1   g23873(.A1(new_n26704_), .A2(new_n26981_), .B(new_n26982_), .ZN(new_n26983_));
  OAI21_X1   g23874(.A1(new_n26983_), .A2(new_n26315_), .B(pi0219), .ZN(new_n26984_));
  NOR2_X1    g23875(.A1(new_n26984_), .A2(new_n26743_), .ZN(new_n26985_));
  INV_X1     g23876(.I(new_n26670_), .ZN(new_n26986_));
  OAI21_X1   g23877(.A1(pi0199), .A2(pi1144), .B(pi1143), .ZN(new_n26987_));
  INV_X1     g23878(.I(new_n26987_), .ZN(new_n26988_));
  NOR3_X1    g23879(.A1(new_n2552_), .A2(pi0199), .A3(pi1143), .ZN(new_n26989_));
  NAND2_X1   g23880(.A1(new_n26322_), .A2(new_n8098_), .ZN(new_n26990_));
  NOR4_X1    g23881(.A1(new_n26990_), .A2(new_n26986_), .A3(new_n26988_), .A4(new_n26989_), .ZN(new_n26991_));
  OAI21_X1   g23882(.A1(pi0199), .A2(pi1145), .B(pi1143), .ZN(new_n26992_));
  NAND3_X1   g23883(.A1(new_n8094_), .A2(new_n3548_), .A3(pi1145), .ZN(new_n26993_));
  NOR3_X1    g23884(.A1(new_n26678_), .A2(pi0200), .A3(new_n26325_), .ZN(new_n26994_));
  AND3_X2    g23885(.A1(new_n26994_), .A2(new_n26992_), .A3(new_n26993_), .Z(new_n26995_));
  OAI21_X1   g23886(.A1(new_n26995_), .A2(new_n26991_), .B(new_n2587_), .ZN(new_n26996_));
  NAND3_X1   g23887(.A1(new_n26693_), .A2(pi0299), .A3(new_n26315_), .ZN(new_n26997_));
  INV_X1     g23888(.I(new_n26370_), .ZN(new_n26998_));
  OR2_X2     g23889(.A1(new_n26983_), .A2(new_n26998_), .Z(new_n26999_));
  NAND3_X1   g23890(.A1(new_n26996_), .A2(new_n26999_), .A3(new_n26997_), .ZN(new_n27000_));
  AOI21_X1   g23891(.A1(new_n27000_), .A2(new_n6845_), .B(new_n26985_), .ZN(new_n27001_));
  NAND2_X1   g23892(.A1(new_n27001_), .A2(pi0213), .ZN(new_n27002_));
  MUX2_X1    g23893(.I0(pi1158), .I1(pi1157), .S(pi0211), .Z(new_n27003_));
  NAND2_X1   g23894(.A1(new_n27003_), .A2(new_n26361_), .ZN(new_n27004_));
  NAND2_X1   g23895(.A1(new_n26909_), .A2(new_n27004_), .ZN(new_n27005_));
  NAND4_X1   g23896(.A1(new_n6845_), .A2(new_n8247_), .A3(new_n26361_), .A4(new_n26819_), .ZN(new_n27006_));
  AOI21_X1   g23897(.A1(new_n11950_), .A2(pi0214), .B(pi0211), .ZN(new_n27007_));
  OAI21_X1   g23898(.A1(pi0214), .A2(pi1155), .B(new_n27007_), .ZN(new_n27008_));
  NAND4_X1   g23899(.A1(new_n27006_), .A2(pi0212), .A3(po1038), .A4(new_n27008_), .ZN(new_n27009_));
  AOI21_X1   g23900(.A1(new_n27009_), .A2(new_n27005_), .B(pi0213), .ZN(new_n27010_));
  NOR2_X1    g23901(.A1(new_n27005_), .A2(new_n26370_), .ZN(new_n27011_));
  OAI21_X1   g23902(.A1(new_n26364_), .A2(new_n26356_), .B(pi0214), .ZN(new_n27012_));
  OAI22_X1   g23903(.A1(new_n27012_), .A2(new_n8076_), .B1(new_n26362_), .B2(new_n26622_), .ZN(new_n27013_));
  AOI21_X1   g23904(.A1(new_n27013_), .A2(new_n26355_), .B(po1038), .ZN(new_n27014_));
  NAND2_X1   g23905(.A1(new_n26996_), .A2(new_n27014_), .ZN(new_n27015_));
  OAI21_X1   g23906(.A1(new_n27015_), .A2(new_n27011_), .B(new_n27010_), .ZN(new_n27016_));
  AOI21_X1   g23907(.A1(new_n27002_), .A2(pi0209), .B(new_n27016_), .ZN(new_n27017_));
  NAND2_X1   g23908(.A1(new_n26606_), .A2(new_n12026_), .ZN(new_n27018_));
  AOI22_X1   g23909(.A1(new_n27018_), .A2(pi1158), .B1(pi0199), .B2(pi1156), .ZN(new_n27019_));
  INV_X1     g23910(.I(new_n27019_), .ZN(new_n27020_));
  NOR2_X1    g23911(.A1(new_n8087_), .A2(pi0200), .ZN(new_n27021_));
  INV_X1     g23912(.I(new_n27021_), .ZN(new_n27022_));
  NOR2_X1    g23913(.A1(new_n27020_), .A2(new_n27022_), .ZN(new_n27023_));
  NOR3_X1    g23914(.A1(new_n27023_), .A2(pi0208), .A3(new_n26585_), .ZN(new_n27024_));
  NOR2_X1    g23915(.A1(new_n27024_), .A2(pi1157), .ZN(new_n27025_));
  NAND2_X1   g23916(.A1(new_n26583_), .A2(pi0207), .ZN(new_n27026_));
  INV_X1     g23917(.I(new_n27026_), .ZN(new_n27027_));
  NOR4_X1    g23918(.A1(new_n27025_), .A2(new_n27027_), .A3(new_n26451_), .A4(new_n26634_), .ZN(new_n27028_));
  INV_X1     g23919(.I(new_n26834_), .ZN(new_n27029_));
  AOI21_X1   g23920(.A1(new_n27026_), .A2(new_n26838_), .B(new_n27029_), .ZN(new_n27030_));
  NOR2_X1    g23921(.A1(new_n11987_), .A2(pi1156), .ZN(new_n27031_));
  INV_X1     g23922(.I(new_n27031_), .ZN(new_n27032_));
  AOI21_X1   g23923(.A1(new_n11987_), .A2(pi1156), .B(pi0200), .ZN(new_n27033_));
  AOI21_X1   g23924(.A1(new_n27032_), .A2(new_n27033_), .B(pi0199), .ZN(new_n27034_));
  OAI21_X1   g23925(.A1(new_n8098_), .A2(pi1156), .B(new_n27034_), .ZN(new_n27035_));
  NOR3_X1    g23926(.A1(new_n8094_), .A2(new_n8098_), .A3(pi1156), .ZN(new_n27036_));
  INV_X1     g23927(.I(new_n27036_), .ZN(new_n27037_));
  AND2_X2    g23928(.A1(new_n27035_), .A2(new_n27037_), .Z(new_n27038_));
  NAND2_X1   g23929(.A1(new_n27038_), .A2(new_n26328_), .ZN(new_n27039_));
  AOI21_X1   g23930(.A1(new_n27039_), .A2(new_n26622_), .B(new_n26424_), .ZN(new_n27040_));
  NOR3_X1    g23931(.A1(new_n27028_), .A2(new_n27030_), .A3(new_n27040_), .ZN(new_n27041_));
  NOR3_X1    g23932(.A1(new_n27020_), .A2(new_n26390_), .A3(new_n26634_), .ZN(new_n27042_));
  INV_X1     g23933(.I(new_n26388_), .ZN(new_n27043_));
  MUX2_X1    g23934(.I0(new_n26415_), .I1(new_n27043_), .S(pi0207), .Z(new_n27044_));
  NOR2_X1    g23935(.A1(new_n27044_), .A2(new_n8088_), .ZN(new_n27045_));
  OAI21_X1   g23936(.A1(new_n27045_), .A2(new_n27042_), .B(new_n12049_), .ZN(new_n27046_));
  INV_X1     g23937(.I(new_n27038_), .ZN(new_n27047_));
  AOI21_X1   g23938(.A1(new_n27047_), .A2(new_n2587_), .B(new_n26457_), .ZN(new_n27048_));
  INV_X1     g23939(.I(new_n26864_), .ZN(new_n27049_));
  NOR2_X1    g23940(.A1(new_n26781_), .A2(new_n27049_), .ZN(new_n27050_));
  OAI21_X1   g23941(.A1(new_n27050_), .A2(new_n27048_), .B(pi1157), .ZN(new_n27051_));
  NAND2_X1   g23942(.A1(new_n27051_), .A2(new_n27046_), .ZN(new_n27052_));
  NOR2_X1    g23943(.A1(new_n27052_), .A2(pi0211), .ZN(new_n27053_));
  XOR2_X1    g23944(.A1(new_n27053_), .A2(new_n27041_), .Z(new_n27054_));
  AOI22_X1   g23945(.A1(new_n27054_), .A2(new_n8078_), .B1(new_n8077_), .B2(new_n27041_), .ZN(new_n27055_));
  INV_X1     g23946(.I(new_n27041_), .ZN(new_n27056_));
  NOR4_X1    g23947(.A1(new_n27053_), .A2(pi0211), .A3(pi0214), .A4(new_n27056_), .ZN(new_n27057_));
  NOR2_X1    g23948(.A1(new_n26757_), .A2(new_n12026_), .ZN(new_n27058_));
  OAI21_X1   g23949(.A1(new_n26411_), .A2(pi1158), .B(new_n27058_), .ZN(new_n27059_));
  OAI21_X1   g23950(.A1(pi0200), .A2(pi1158), .B(new_n8094_), .ZN(new_n27060_));
  NAND3_X1   g23951(.A1(new_n27059_), .A2(new_n26328_), .A3(new_n27060_), .ZN(new_n27061_));
  NAND2_X1   g23952(.A1(new_n27061_), .A2(new_n26364_), .ZN(new_n27062_));
  NOR2_X1    g23953(.A1(new_n26388_), .A2(new_n26363_), .ZN(new_n27063_));
  OAI21_X1   g23954(.A1(new_n27063_), .A2(new_n8087_), .B(new_n26844_), .ZN(new_n27064_));
  AOI22_X1   g23955(.A1(new_n27064_), .A2(new_n26834_), .B1(new_n26423_), .B2(new_n27062_), .ZN(new_n27065_));
  NOR2_X1    g23956(.A1(new_n27063_), .A2(new_n8087_), .ZN(new_n27066_));
  NOR2_X1    g23957(.A1(new_n27066_), .A2(new_n26847_), .ZN(new_n27067_));
  NAND3_X1   g23958(.A1(new_n27067_), .A2(new_n8088_), .A3(new_n26363_), .ZN(new_n27068_));
  AOI21_X1   g23959(.A1(new_n8088_), .A2(new_n26364_), .B(new_n27067_), .ZN(new_n27069_));
  NOR3_X1    g23960(.A1(new_n27069_), .A2(pi1157), .A3(new_n27042_), .ZN(new_n27070_));
  AOI21_X1   g23961(.A1(new_n27070_), .A2(new_n27068_), .B(new_n27065_), .ZN(new_n27071_));
  OR3_X2     g23962(.A1(new_n27057_), .A2(new_n26597_), .A3(new_n27071_), .Z(new_n27072_));
  INV_X1     g23963(.I(new_n27046_), .ZN(new_n27073_));
  AOI21_X1   g23964(.A1(new_n26420_), .A2(new_n8087_), .B(pi0208), .ZN(new_n27074_));
  NAND2_X1   g23965(.A1(new_n26791_), .A2(new_n27074_), .ZN(new_n27075_));
  NOR3_X1    g23966(.A1(new_n27047_), .A2(pi0208), .A3(new_n26492_), .ZN(new_n27076_));
  INV_X1     g23967(.I(new_n27076_), .ZN(new_n27077_));
  AOI21_X1   g23968(.A1(new_n27077_), .A2(new_n27075_), .B(new_n12049_), .ZN(new_n27078_));
  NOR2_X1    g23969(.A1(new_n27073_), .A2(new_n27078_), .ZN(new_n27079_));
  OAI21_X1   g23970(.A1(new_n27079_), .A2(pi0214), .B(new_n8076_), .ZN(new_n27080_));
  INV_X1     g23971(.I(new_n27080_), .ZN(new_n27081_));
  NAND2_X1   g23972(.A1(new_n27052_), .A2(pi0211), .ZN(new_n27082_));
  MUX2_X1    g23973(.I0(new_n26827_), .I1(new_n11987_), .S(pi0299), .Z(new_n27083_));
  OAI21_X1   g23974(.A1(new_n27083_), .A2(pi0207), .B(pi0208), .ZN(new_n27084_));
  AOI21_X1   g23975(.A1(new_n26388_), .A2(new_n11987_), .B(pi0207), .ZN(new_n27085_));
  OAI21_X1   g23976(.A1(new_n26526_), .A2(new_n11987_), .B(new_n27085_), .ZN(new_n27086_));
  INV_X1     g23977(.I(new_n27086_), .ZN(new_n27087_));
  NAND2_X1   g23978(.A1(new_n27087_), .A2(new_n27084_), .ZN(new_n27088_));
  NAND2_X1   g23979(.A1(new_n11987_), .A2(pi0299), .ZN(new_n27089_));
  NAND4_X1   g23980(.A1(new_n27086_), .A2(new_n8087_), .A3(new_n26462_), .A4(new_n27089_), .ZN(new_n27090_));
  OAI21_X1   g23981(.A1(new_n8161_), .A2(new_n8087_), .B(new_n2587_), .ZN(new_n27091_));
  NAND2_X1   g23982(.A1(new_n27091_), .A2(pi1158), .ZN(new_n27092_));
  INV_X1     g23983(.I(new_n27092_), .ZN(new_n27093_));
  NOR2_X1    g23984(.A1(new_n26379_), .A2(pi1156), .ZN(new_n27094_));
  OAI22_X1   g23985(.A1(new_n26412_), .A2(new_n27094_), .B1(new_n11987_), .B2(new_n26606_), .ZN(new_n27095_));
  NOR2_X1    g23986(.A1(pi0207), .A2(pi1157), .ZN(new_n27096_));
  AOI21_X1   g23987(.A1(new_n27095_), .A2(new_n27096_), .B(new_n27093_), .ZN(new_n27097_));
  OAI21_X1   g23988(.A1(new_n27097_), .A2(new_n26424_), .B(new_n8077_), .ZN(new_n27098_));
  NAND3_X1   g23989(.A1(new_n26328_), .A2(new_n26395_), .A3(pi1156), .ZN(new_n27099_));
  NAND3_X1   g23990(.A1(new_n27092_), .A2(new_n8088_), .A3(new_n27099_), .ZN(new_n27100_));
  NOR4_X1    g23991(.A1(new_n27098_), .A2(pi1157), .A3(new_n27029_), .A4(new_n27100_), .ZN(new_n27101_));
  NAND3_X1   g23992(.A1(new_n27088_), .A2(new_n27090_), .A3(new_n27101_), .ZN(new_n27102_));
  NAND3_X1   g23993(.A1(new_n27082_), .A2(pi0214), .A3(new_n27102_), .ZN(new_n27103_));
  AOI21_X1   g23994(.A1(new_n27103_), .A2(new_n27081_), .B(pi0219), .ZN(new_n27104_));
  OAI21_X1   g23995(.A1(new_n27055_), .A2(new_n27072_), .B(new_n27104_), .ZN(new_n27105_));
  OAI21_X1   g23996(.A1(new_n27073_), .A2(new_n27078_), .B(new_n26319_), .ZN(new_n27106_));
  AOI21_X1   g23997(.A1(new_n8160_), .A2(pi1157), .B(pi0299), .ZN(new_n27107_));
  NAND2_X1   g23998(.A1(new_n26827_), .A2(new_n27107_), .ZN(new_n27108_));
  NAND3_X1   g23999(.A1(new_n27108_), .A2(new_n8087_), .A3(new_n26513_), .ZN(new_n27109_));
  NOR2_X1    g24000(.A1(new_n27023_), .A2(pi1157), .ZN(new_n27110_));
  NOR3_X1    g24001(.A1(new_n27110_), .A2(pi0208), .A3(new_n27061_), .ZN(new_n27111_));
  NOR2_X1    g24002(.A1(new_n27111_), .A2(pi0208), .ZN(new_n27112_));
  OAI22_X1   g24003(.A1(new_n27112_), .A2(new_n26509_), .B1(new_n26512_), .B2(new_n27109_), .ZN(new_n27113_));
  OAI21_X1   g24004(.A1(new_n26319_), .A2(new_n27113_), .B(new_n27106_), .ZN(new_n27114_));
  AOI21_X1   g24005(.A1(new_n27114_), .A2(pi0219), .B(po1038), .ZN(new_n27115_));
  NOR2_X1    g24006(.A1(new_n27080_), .A2(pi0214), .ZN(new_n27116_));
  NAND2_X1   g24007(.A1(new_n27113_), .A2(pi0211), .ZN(new_n27117_));
  NOR2_X1    g24008(.A1(new_n26478_), .A2(pi0207), .ZN(new_n27118_));
  AOI21_X1   g24009(.A1(new_n27108_), .A2(new_n27118_), .B(new_n26490_), .ZN(new_n27119_));
  NOR2_X1    g24010(.A1(new_n27112_), .A2(new_n26480_), .ZN(new_n27120_));
  NOR4_X1    g24011(.A1(new_n27120_), .A2(new_n8077_), .A3(pi0214), .A4(new_n27119_), .ZN(new_n27121_));
  AOI21_X1   g24012(.A1(new_n27121_), .A2(new_n27117_), .B(new_n8250_), .ZN(new_n27122_));
  NOR3_X1    g24013(.A1(new_n27116_), .A2(pi0219), .A3(new_n27122_), .ZN(new_n27123_));
  OAI22_X1   g24014(.A1(new_n27123_), .A2(new_n27115_), .B1(new_n26743_), .B2(new_n26984_), .ZN(new_n27124_));
  INV_X1     g24015(.I(new_n26925_), .ZN(new_n27125_));
  OAI21_X1   g24016(.A1(new_n27042_), .A2(new_n27125_), .B(new_n12049_), .ZN(new_n27126_));
  NAND4_X1   g24017(.A1(new_n26462_), .A2(new_n8087_), .A3(pi1157), .A4(new_n26554_), .ZN(new_n27127_));
  NAND4_X1   g24018(.A1(new_n27126_), .A2(new_n26550_), .A3(new_n26489_), .A4(new_n27127_), .ZN(new_n27128_));
  NOR2_X1    g24019(.A1(new_n27042_), .A2(pi1157), .ZN(new_n27129_));
  NOR2_X1    g24020(.A1(new_n27129_), .A2(new_n27061_), .ZN(new_n27130_));
  NOR4_X1    g24021(.A1(new_n27130_), .A2(pi0208), .A3(new_n8078_), .A4(new_n26356_), .ZN(new_n27131_));
  AOI21_X1   g24022(.A1(new_n27131_), .A2(new_n27128_), .B(new_n8076_), .ZN(new_n27132_));
  OAI21_X1   g24023(.A1(new_n27071_), .A2(pi0214), .B(new_n27132_), .ZN(new_n27133_));
  NAND2_X1   g24024(.A1(new_n27056_), .A2(new_n26361_), .ZN(new_n27134_));
  AOI21_X1   g24025(.A1(new_n27133_), .A2(new_n27134_), .B(pi0211), .ZN(new_n27135_));
  NAND2_X1   g24026(.A1(new_n27106_), .A2(new_n8247_), .ZN(new_n27136_));
  NOR3_X1    g24027(.A1(new_n27010_), .A2(pi0209), .A3(po1038), .ZN(new_n27137_));
  OAI21_X1   g24028(.A1(new_n27135_), .A2(new_n27136_), .B(new_n27137_), .ZN(new_n27138_));
  AOI21_X1   g24029(.A1(new_n27124_), .A2(new_n24753_), .B(new_n27138_), .ZN(new_n27139_));
  AOI21_X1   g24030(.A1(new_n27105_), .A2(new_n27139_), .B(new_n27017_), .ZN(new_n27140_));
  MUX2_X1    g24031(.I0(new_n27140_), .I1(pi0237), .S(new_n26307_), .Z(po0394));
  NAND2_X1   g24032(.A1(new_n26532_), .A2(new_n26937_), .ZN(new_n27142_));
  INV_X1     g24033(.I(new_n26608_), .ZN(new_n27143_));
  NOR2_X1    g24034(.A1(new_n26434_), .A2(new_n11893_), .ZN(new_n27144_));
  INV_X1     g24035(.I(new_n27144_), .ZN(new_n27145_));
  AOI21_X1   g24036(.A1(new_n27143_), .A2(new_n27145_), .B(new_n8087_), .ZN(new_n27146_));
  AOI21_X1   g24037(.A1(new_n8087_), .A2(new_n26531_), .B(new_n27146_), .ZN(new_n27147_));
  NAND3_X1   g24038(.A1(new_n27146_), .A2(new_n26531_), .A3(new_n8087_), .ZN(new_n27148_));
  NAND2_X1   g24039(.A1(new_n27148_), .A2(pi0208), .ZN(new_n27149_));
  OAI21_X1   g24040(.A1(new_n27147_), .A2(new_n27149_), .B(new_n27142_), .ZN(new_n27150_));
  NOR2_X1    g24041(.A1(new_n27150_), .A2(pi0211), .ZN(new_n27151_));
  NOR2_X1    g24042(.A1(new_n26412_), .A2(new_n26711_), .ZN(new_n27152_));
  INV_X1     g24043(.I(new_n27152_), .ZN(new_n27153_));
  AOI21_X1   g24044(.A1(new_n27143_), .A2(new_n27153_), .B(new_n8089_), .ZN(new_n27154_));
  NOR2_X1    g24045(.A1(new_n26884_), .A2(new_n27154_), .ZN(new_n27155_));
  INV_X1     g24046(.I(new_n27155_), .ZN(new_n27156_));
  NOR2_X1    g24047(.A1(new_n27156_), .A2(new_n8077_), .ZN(new_n27157_));
  NOR2_X1    g24048(.A1(new_n27157_), .A2(new_n27151_), .ZN(new_n27158_));
  INV_X1     g24049(.I(new_n27158_), .ZN(new_n27159_));
  NAND2_X1   g24050(.A1(new_n27159_), .A2(new_n26693_), .ZN(new_n27160_));
  NOR2_X1    g24051(.A1(new_n8268_), .A2(new_n11950_), .ZN(new_n27161_));
  NOR2_X1    g24052(.A1(new_n26608_), .A2(new_n27161_), .ZN(new_n27162_));
  NOR2_X1    g24053(.A1(new_n26396_), .A2(new_n11893_), .ZN(new_n27163_));
  OAI21_X1   g24054(.A1(new_n27163_), .A2(pi0299), .B(new_n11950_), .ZN(new_n27164_));
  NAND3_X1   g24055(.A1(new_n27162_), .A2(new_n26549_), .A3(new_n27164_), .ZN(new_n27165_));
  AOI21_X1   g24056(.A1(new_n26658_), .A2(new_n26493_), .B(pi0207), .ZN(new_n27166_));
  NAND2_X1   g24057(.A1(new_n27165_), .A2(new_n27166_), .ZN(new_n27167_));
  NAND3_X1   g24058(.A1(new_n27165_), .A2(pi0207), .A3(new_n27166_), .ZN(new_n27168_));
  NAND3_X1   g24059(.A1(new_n27168_), .A2(new_n27167_), .A3(new_n26563_), .ZN(new_n27169_));
  INV_X1     g24060(.I(new_n27169_), .ZN(new_n27170_));
  INV_X1     g24061(.I(new_n26945_), .ZN(new_n27171_));
  NAND2_X1   g24062(.A1(new_n27162_), .A2(new_n27153_), .ZN(new_n27172_));
  AOI21_X1   g24063(.A1(new_n27171_), .A2(new_n8087_), .B(new_n27172_), .ZN(new_n27173_));
  NAND3_X1   g24064(.A1(new_n26945_), .A2(new_n27172_), .A3(new_n8087_), .ZN(new_n27174_));
  NAND2_X1   g24065(.A1(new_n27174_), .A2(pi0208), .ZN(new_n27175_));
  OAI22_X1   g24066(.A1(new_n26548_), .A2(new_n26943_), .B1(new_n27173_), .B2(new_n27175_), .ZN(new_n27176_));
  MUX2_X1    g24067(.I0(new_n27176_), .I1(new_n27170_), .S(new_n8077_), .Z(new_n27177_));
  NOR2_X1    g24068(.A1(new_n27177_), .A2(new_n26362_), .ZN(new_n27178_));
  NOR2_X1    g24069(.A1(new_n8077_), .A2(pi0214), .ZN(new_n27179_));
  NOR2_X1    g24070(.A1(new_n26534_), .A2(new_n27179_), .ZN(new_n27180_));
  INV_X1     g24071(.I(new_n27180_), .ZN(new_n27181_));
  NAND2_X1   g24072(.A1(new_n27150_), .A2(new_n8079_), .ZN(new_n27182_));
  AOI21_X1   g24073(.A1(new_n27170_), .A2(new_n26557_), .B(new_n8076_), .ZN(new_n27183_));
  NAND2_X1   g24074(.A1(new_n27182_), .A2(new_n27183_), .ZN(new_n27184_));
  AOI21_X1   g24075(.A1(new_n27176_), .A2(new_n27181_), .B(new_n27184_), .ZN(new_n27185_));
  OAI21_X1   g24076(.A1(new_n27178_), .A2(new_n27185_), .B(new_n8247_), .ZN(new_n27186_));
  NOR2_X1    g24077(.A1(new_n27156_), .A2(new_n26342_), .ZN(new_n27187_));
  OAI21_X1   g24078(.A1(new_n27187_), .A2(po1038), .B(new_n26374_), .ZN(new_n27188_));
  AOI21_X1   g24079(.A1(new_n27160_), .A2(new_n27186_), .B(new_n27188_), .ZN(new_n27189_));
  NOR2_X1    g24080(.A1(new_n8161_), .A2(pi0207), .ZN(new_n27190_));
  NOR3_X1    g24081(.A1(new_n26493_), .A2(new_n8088_), .A3(new_n27190_), .ZN(new_n27191_));
  NOR2_X1    g24082(.A1(new_n26396_), .A2(new_n26492_), .ZN(new_n27192_));
  NOR2_X1    g24083(.A1(new_n27191_), .A2(new_n27192_), .ZN(new_n27193_));
  INV_X1     g24084(.I(new_n27193_), .ZN(new_n27194_));
  NOR2_X1    g24085(.A1(new_n27194_), .A2(pi0214), .ZN(new_n27195_));
  NOR2_X1    g24086(.A1(new_n26606_), .A2(new_n26677_), .ZN(new_n27196_));
  INV_X1     g24087(.I(new_n27196_), .ZN(new_n27197_));
  NOR2_X1    g24088(.A1(new_n27197_), .A2(new_n11893_), .ZN(new_n27198_));
  INV_X1     g24089(.I(new_n27198_), .ZN(new_n27199_));
  AOI21_X1   g24090(.A1(new_n27195_), .A2(new_n27199_), .B(pi0212), .ZN(new_n27200_));
  NAND2_X1   g24091(.A1(new_n27200_), .A2(new_n8078_), .ZN(new_n27201_));
  INV_X1     g24092(.I(new_n26626_), .ZN(new_n27202_));
  NAND2_X1   g24093(.A1(new_n27202_), .A2(new_n8087_), .ZN(new_n27203_));
  AOI21_X1   g24094(.A1(new_n8268_), .A2(pi0207), .B(new_n8088_), .ZN(new_n27204_));
  AOI22_X1   g24095(.A1(new_n27203_), .A2(new_n27204_), .B1(new_n26456_), .B2(new_n26626_), .ZN(new_n27205_));
  INV_X1     g24096(.I(new_n27205_), .ZN(new_n27206_));
  NOR3_X1    g24097(.A1(new_n27206_), .A2(pi0211), .A3(new_n26553_), .ZN(new_n27207_));
  NOR2_X1    g24098(.A1(new_n26677_), .A2(new_n8161_), .ZN(new_n27208_));
  NOR2_X1    g24099(.A1(new_n27208_), .A2(pi0299), .ZN(new_n27209_));
  NOR3_X1    g24100(.A1(new_n27209_), .A2(new_n8077_), .A3(new_n11893_), .ZN(new_n27210_));
  NOR2_X1    g24101(.A1(new_n27193_), .A2(new_n8248_), .ZN(new_n27211_));
  OAI21_X1   g24102(.A1(new_n27207_), .A2(new_n27210_), .B(new_n27211_), .ZN(new_n27212_));
  NAND3_X1   g24103(.A1(new_n27201_), .A2(new_n8247_), .A3(new_n27212_), .ZN(new_n27213_));
  INV_X1     g24104(.I(new_n27207_), .ZN(new_n27214_));
  OAI21_X1   g24105(.A1(new_n8161_), .A2(pi0207), .B(new_n2587_), .ZN(new_n27215_));
  NOR2_X1    g24106(.A1(new_n8098_), .A2(new_n8087_), .ZN(new_n27216_));
  NOR2_X1    g24107(.A1(new_n27216_), .A2(pi0199), .ZN(new_n27217_));
  INV_X1     g24108(.I(new_n27217_), .ZN(new_n27218_));
  AOI21_X1   g24109(.A1(new_n27218_), .A2(new_n2587_), .B(new_n8088_), .ZN(new_n27219_));
  INV_X1     g24110(.I(new_n27219_), .ZN(new_n27220_));
  AOI21_X1   g24111(.A1(new_n11893_), .A2(new_n27215_), .B(new_n27220_), .ZN(new_n27221_));
  NAND2_X1   g24112(.A1(new_n26460_), .A2(pi1153), .ZN(new_n27222_));
  NOR2_X1    g24113(.A1(new_n8662_), .A2(new_n8087_), .ZN(new_n27223_));
  AOI21_X1   g24114(.A1(new_n27223_), .A2(new_n27222_), .B(new_n26937_), .ZN(new_n27224_));
  OAI21_X1   g24115(.A1(new_n27221_), .A2(new_n27224_), .B(pi0211), .ZN(new_n27225_));
  AOI21_X1   g24116(.A1(new_n27214_), .A2(new_n27225_), .B(new_n8250_), .ZN(new_n27226_));
  NOR2_X1    g24117(.A1(new_n27206_), .A2(new_n26650_), .ZN(new_n27227_));
  NAND2_X1   g24118(.A1(new_n26964_), .A2(pi0299), .ZN(new_n27228_));
  OAI21_X1   g24119(.A1(new_n27227_), .A2(new_n27228_), .B(new_n8247_), .ZN(new_n27229_));
  NOR2_X1    g24120(.A1(po1038), .A2(pi1151), .ZN(new_n27230_));
  OAI21_X1   g24121(.A1(pi0200), .A2(pi0208), .B(pi0207), .ZN(new_n27231_));
  NOR2_X1    g24122(.A1(new_n8170_), .A2(new_n27231_), .ZN(new_n27232_));
  INV_X1     g24123(.I(new_n27232_), .ZN(new_n27233_));
  AOI21_X1   g24124(.A1(new_n8090_), .A2(new_n26624_), .B(new_n27233_), .ZN(new_n27234_));
  INV_X1     g24125(.I(new_n27234_), .ZN(new_n27235_));
  NOR2_X1    g24126(.A1(new_n26359_), .A2(pi0211), .ZN(new_n27236_));
  OAI21_X1   g24127(.A1(new_n26342_), .A2(new_n27236_), .B(new_n27235_), .ZN(new_n27237_));
  AOI21_X1   g24128(.A1(new_n27237_), .A2(new_n26719_), .B(new_n27230_), .ZN(new_n27238_));
  OAI21_X1   g24129(.A1(new_n27226_), .A2(new_n27229_), .B(new_n27238_), .ZN(new_n27239_));
  NOR3_X1    g24130(.A1(new_n26627_), .A2(new_n26634_), .A3(new_n26757_), .ZN(new_n27240_));
  AOI21_X1   g24131(.A1(new_n26645_), .A2(new_n26457_), .B(new_n27240_), .ZN(new_n27241_));
  OAI21_X1   g24132(.A1(pi0211), .A2(new_n26523_), .B(new_n26553_), .ZN(new_n27242_));
  NAND3_X1   g24133(.A1(new_n26554_), .A2(new_n8077_), .A3(new_n26523_), .ZN(new_n27243_));
  NAND4_X1   g24134(.A1(new_n27241_), .A2(new_n26314_), .A3(new_n27242_), .A4(new_n27243_), .ZN(new_n27244_));
  NOR2_X1    g24135(.A1(new_n27196_), .A2(pi0214), .ZN(new_n27245_));
  NOR2_X1    g24136(.A1(new_n8077_), .A2(new_n2587_), .ZN(new_n27246_));
  NOR2_X1    g24137(.A1(new_n27209_), .A2(new_n27246_), .ZN(new_n27247_));
  INV_X1     g24138(.I(new_n27247_), .ZN(new_n27248_));
  AOI21_X1   g24139(.A1(new_n8076_), .A2(new_n27245_), .B(new_n27248_), .ZN(new_n27249_));
  NOR2_X1    g24140(.A1(new_n27249_), .A2(new_n11893_), .ZN(new_n27250_));
  INV_X1     g24141(.I(pi1151), .ZN(new_n27251_));
  NOR2_X1    g24142(.A1(po1038), .A2(new_n27251_), .ZN(new_n27252_));
  NOR4_X1    g24143(.A1(new_n27250_), .A2(new_n8247_), .A3(new_n27194_), .A4(new_n27252_), .ZN(new_n27253_));
  NOR2_X1    g24144(.A1(new_n27253_), .A2(pi1152), .ZN(new_n27254_));
  NAND4_X1   g24145(.A1(new_n27254_), .A2(new_n27239_), .A3(new_n27213_), .A4(new_n27244_), .ZN(new_n27255_));
  AOI21_X1   g24146(.A1(new_n26396_), .A2(new_n26328_), .B(new_n8088_), .ZN(new_n27256_));
  NOR2_X1    g24147(.A1(new_n27256_), .A2(new_n26562_), .ZN(new_n27257_));
  NAND2_X1   g24148(.A1(new_n26379_), .A2(pi1153), .ZN(new_n27258_));
  OAI21_X1   g24149(.A1(new_n26640_), .A2(pi1153), .B(new_n27258_), .ZN(new_n27259_));
  OAI22_X1   g24150(.A1(new_n27259_), .A2(new_n11912_), .B1(new_n26390_), .B2(new_n26609_), .ZN(new_n27260_));
  OAI22_X1   g24151(.A1(new_n27260_), .A2(new_n27257_), .B1(new_n26396_), .B2(new_n26986_), .ZN(new_n27261_));
  OAI21_X1   g24152(.A1(new_n27261_), .A2(new_n2587_), .B(new_n27228_), .ZN(new_n27262_));
  NAND2_X1   g24153(.A1(new_n27262_), .A2(pi0214), .ZN(new_n27263_));
  INV_X1     g24154(.I(new_n26756_), .ZN(new_n27264_));
  NOR3_X1    g24155(.A1(new_n27256_), .A2(pi0200), .A3(new_n26455_), .ZN(new_n27265_));
  AOI21_X1   g24156(.A1(new_n27022_), .A2(new_n2587_), .B(pi0208), .ZN(new_n27266_));
  NOR2_X1    g24157(.A1(new_n27265_), .A2(new_n27266_), .ZN(new_n27267_));
  NOR2_X1    g24158(.A1(new_n26986_), .A2(new_n26396_), .ZN(new_n27268_));
  AOI21_X1   g24159(.A1(new_n26389_), .A2(new_n26678_), .B(new_n27268_), .ZN(new_n27269_));
  NOR2_X1    g24160(.A1(new_n27269_), .A2(new_n8077_), .ZN(new_n27270_));
  AOI21_X1   g24161(.A1(new_n8077_), .A2(new_n27267_), .B(new_n27270_), .ZN(new_n27271_));
  INV_X1     g24162(.I(new_n27269_), .ZN(new_n27272_));
  NOR2_X1    g24163(.A1(new_n27272_), .A2(new_n26613_), .ZN(new_n27273_));
  NAND2_X1   g24164(.A1(new_n27273_), .A2(new_n26342_), .ZN(new_n27274_));
  NAND3_X1   g24165(.A1(new_n27274_), .A2(new_n27271_), .A3(new_n27264_), .ZN(new_n27275_));
  OAI21_X1   g24166(.A1(new_n27275_), .A2(new_n8247_), .B(new_n27252_), .ZN(new_n27276_));
  NOR2_X1    g24167(.A1(new_n27267_), .A2(new_n26756_), .ZN(new_n27277_));
  INV_X1     g24168(.I(new_n27273_), .ZN(new_n27278_));
  NAND3_X1   g24169(.A1(new_n27261_), .A2(new_n8077_), .A3(new_n8078_), .ZN(new_n27281_));
  OAI21_X1   g24170(.A1(new_n27273_), .A2(pi0214), .B(new_n8076_), .ZN(new_n27282_));
  NOR2_X1    g24171(.A1(new_n27282_), .A2(pi0219), .ZN(new_n27283_));
  NAND4_X1   g24172(.A1(new_n27276_), .A2(new_n27263_), .A3(new_n27281_), .A4(new_n27283_), .ZN(new_n27284_));
  INV_X1     g24173(.I(new_n27210_), .ZN(new_n27285_));
  OAI21_X1   g24174(.A1(new_n27198_), .A2(new_n26356_), .B(new_n8077_), .ZN(new_n27286_));
  AOI21_X1   g24175(.A1(new_n27286_), .A2(new_n27285_), .B(new_n8248_), .ZN(new_n27287_));
  NOR3_X1    g24176(.A1(new_n26963_), .A2(new_n26910_), .A3(pi0299), .ZN(new_n27288_));
  NOR4_X1    g24177(.A1(new_n27287_), .A2(new_n26652_), .A3(new_n27198_), .A4(new_n27288_), .ZN(new_n27289_));
  OAI21_X1   g24178(.A1(new_n27250_), .A2(new_n26375_), .B(new_n27230_), .ZN(new_n27290_));
  OAI21_X1   g24179(.A1(new_n27290_), .A2(new_n27289_), .B(new_n26604_), .ZN(new_n27291_));
  NAND2_X1   g24180(.A1(new_n27284_), .A2(new_n27291_), .ZN(new_n27292_));
  AOI21_X1   g24181(.A1(new_n27292_), .A2(new_n27255_), .B(pi0209), .ZN(new_n27293_));
  NOR3_X1    g24182(.A1(new_n26311_), .A2(new_n8247_), .A3(new_n26737_), .ZN(new_n27294_));
  NOR2_X1    g24183(.A1(new_n27294_), .A2(pi0213), .ZN(new_n27295_));
  OAI21_X1   g24184(.A1(new_n27189_), .A2(new_n27293_), .B(new_n27295_), .ZN(new_n27296_));
  INV_X1     g24185(.I(new_n27157_), .ZN(new_n27297_));
  OAI21_X1   g24186(.A1(new_n26877_), .A2(new_n27165_), .B(new_n26881_), .ZN(new_n27298_));
  OAI21_X1   g24187(.A1(pi0211), .A2(new_n27298_), .B(new_n27297_), .ZN(new_n27299_));
  NAND2_X1   g24188(.A1(new_n27299_), .A2(new_n26342_), .ZN(new_n27300_));
  INV_X1     g24189(.I(new_n27300_), .ZN(new_n27301_));
  NOR2_X1    g24190(.A1(new_n27301_), .A2(new_n27187_), .ZN(new_n27302_));
  NAND2_X1   g24191(.A1(new_n27301_), .A2(new_n27187_), .ZN(new_n27303_));
  NAND2_X1   g24192(.A1(new_n27303_), .A2(pi0219), .ZN(new_n27304_));
  OAI21_X1   g24193(.A1(new_n27304_), .A2(new_n27302_), .B(new_n6845_), .ZN(new_n27305_));
  AOI21_X1   g24194(.A1(new_n27155_), .A2(new_n8078_), .B(pi0212), .ZN(new_n27306_));
  NOR2_X1    g24195(.A1(new_n27298_), .A2(new_n8077_), .ZN(new_n27307_));
  NOR2_X1    g24196(.A1(new_n27307_), .A2(new_n27151_), .ZN(new_n27308_));
  INV_X1     g24197(.I(new_n27308_), .ZN(new_n27309_));
  NAND2_X1   g24198(.A1(new_n27309_), .A2(pi0214), .ZN(new_n27310_));
  OAI21_X1   g24199(.A1(new_n27310_), .A2(new_n27306_), .B(new_n8247_), .ZN(new_n27311_));
  NOR2_X1    g24200(.A1(new_n8250_), .A2(new_n8077_), .ZN(new_n27312_));
  AOI21_X1   g24201(.A1(new_n8446_), .A2(new_n11893_), .B(new_n27312_), .ZN(new_n27313_));
  INV_X1     g24202(.I(new_n27313_), .ZN(new_n27314_));
  NOR2_X1    g24203(.A1(new_n8081_), .A2(new_n26719_), .ZN(new_n27315_));
  INV_X1     g24204(.I(new_n27315_), .ZN(new_n27316_));
  NOR2_X1    g24205(.A1(new_n27316_), .A2(new_n6845_), .ZN(new_n27317_));
  INV_X1     g24206(.I(new_n27317_), .ZN(new_n27318_));
  NOR2_X1    g24207(.A1(new_n27318_), .A2(new_n27314_), .ZN(new_n27319_));
  INV_X1     g24208(.I(new_n27319_), .ZN(new_n27320_));
  NOR2_X1    g24209(.A1(new_n26743_), .A2(new_n8082_), .ZN(new_n27321_));
  NOR2_X1    g24210(.A1(new_n27321_), .A2(pi1151), .ZN(new_n27322_));
  INV_X1     g24211(.I(new_n27322_), .ZN(new_n27323_));
  NOR2_X1    g24212(.A1(new_n27323_), .A2(new_n27320_), .ZN(new_n27324_));
  INV_X1     g24213(.I(new_n27324_), .ZN(new_n27325_));
  NAND4_X1   g24214(.A1(new_n27308_), .A2(new_n8076_), .A3(pi0214), .A4(new_n27298_), .ZN(new_n27326_));
  NAND2_X1   g24215(.A1(new_n27326_), .A2(new_n27325_), .ZN(new_n27327_));
  NOR2_X1    g24216(.A1(new_n27311_), .A2(new_n27327_), .ZN(new_n27328_));
  NOR2_X1    g24217(.A1(new_n27299_), .A2(new_n8078_), .ZN(new_n27329_));
  NOR2_X1    g24218(.A1(new_n27329_), .A2(pi0212), .ZN(new_n27330_));
  OAI21_X1   g24219(.A1(pi0214), .A2(new_n27309_), .B(new_n27330_), .ZN(new_n27331_));
  NOR2_X1    g24220(.A1(new_n27319_), .A2(pi1151), .ZN(new_n27332_));
  AOI21_X1   g24221(.A1(new_n27155_), .A2(pi0219), .B(po1038), .ZN(new_n27333_));
  NOR3_X1    g24222(.A1(new_n27311_), .A2(new_n27332_), .A3(new_n27333_), .ZN(new_n27334_));
  AOI22_X1   g24223(.A1(new_n27305_), .A2(new_n27328_), .B1(new_n27334_), .B2(new_n27331_), .ZN(new_n27335_));
  NAND2_X1   g24224(.A1(new_n26374_), .A2(new_n26604_), .ZN(new_n27336_));
  NAND3_X1   g24225(.A1(new_n27159_), .A2(new_n8078_), .A3(new_n27156_), .ZN(new_n27337_));
  OAI21_X1   g24226(.A1(pi0214), .A2(new_n27156_), .B(new_n27158_), .ZN(new_n27338_));
  NAND3_X1   g24227(.A1(new_n27337_), .A2(new_n27338_), .A3(new_n8076_), .ZN(new_n27342_));
  NOR2_X1    g24228(.A1(new_n6845_), .A2(pi0219), .ZN(new_n27343_));
  NOR2_X1    g24229(.A1(new_n26473_), .A2(pi0211), .ZN(new_n27344_));
  INV_X1     g24230(.I(new_n27344_), .ZN(new_n27345_));
  NOR2_X1    g24231(.A1(new_n27345_), .A2(new_n11893_), .ZN(new_n27346_));
  NOR2_X1    g24232(.A1(new_n6845_), .A2(pi0219), .ZN(new_n27347_));
  AOI21_X1   g24233(.A1(new_n27347_), .A2(new_n27346_), .B(pi1151), .ZN(new_n27348_));
  INV_X1     g24234(.I(new_n27348_), .ZN(new_n27349_));
  NOR2_X1    g24235(.A1(new_n26473_), .A2(pi0219), .ZN(new_n27350_));
  OAI21_X1   g24236(.A1(new_n27156_), .A2(new_n27350_), .B(new_n6845_), .ZN(new_n27351_));
  INV_X1     g24237(.I(new_n27350_), .ZN(new_n27352_));
  NOR2_X1    g24238(.A1(new_n27158_), .A2(new_n27352_), .ZN(new_n27353_));
  AOI21_X1   g24239(.A1(new_n27353_), .A2(new_n27351_), .B(new_n27349_), .ZN(new_n27354_));
  INV_X1     g24240(.I(new_n8082_), .ZN(new_n27355_));
  NOR4_X1    g24241(.A1(new_n26311_), .A2(new_n27346_), .A3(pi1151), .A4(new_n27355_), .ZN(new_n27356_));
  OAI21_X1   g24242(.A1(new_n27354_), .A2(pi1152), .B(new_n27356_), .ZN(new_n27357_));
  AOI21_X1   g24243(.A1(new_n27342_), .A2(new_n27343_), .B(new_n27357_), .ZN(new_n27358_));
  OAI21_X1   g24244(.A1(new_n27335_), .A2(new_n27336_), .B(new_n27358_), .ZN(new_n27359_));
  NOR2_X1    g24245(.A1(new_n27194_), .A2(new_n27198_), .ZN(new_n27360_));
  INV_X1     g24246(.I(new_n27360_), .ZN(new_n27361_));
  INV_X1     g24247(.I(new_n27241_), .ZN(new_n27362_));
  NOR2_X1    g24248(.A1(new_n27362_), .A2(pi0211), .ZN(new_n27363_));
  NOR2_X1    g24249(.A1(new_n27363_), .A2(new_n27361_), .ZN(new_n27364_));
  NOR2_X1    g24250(.A1(new_n27361_), .A2(pi0214), .ZN(new_n27365_));
  NOR3_X1    g24251(.A1(new_n27363_), .A2(new_n27361_), .A3(new_n8078_), .ZN(new_n27366_));
  NOR3_X1    g24252(.A1(new_n27366_), .A2(pi0212), .A3(new_n27365_), .ZN(new_n27367_));
  OR2_X2     g24253(.A1(new_n27367_), .A2(new_n27364_), .Z(new_n27368_));
  AOI21_X1   g24254(.A1(new_n27368_), .A2(pi0219), .B(po1038), .ZN(new_n27369_));
  OAI22_X1   g24255(.A1(new_n27362_), .A2(new_n8077_), .B1(new_n11893_), .B2(new_n27209_), .ZN(new_n27370_));
  NAND2_X1   g24256(.A1(new_n27370_), .A2(new_n27195_), .ZN(new_n27371_));
  NOR2_X1    g24257(.A1(new_n27241_), .A2(new_n8078_), .ZN(new_n27372_));
  NOR2_X1    g24258(.A1(new_n27372_), .A2(new_n8076_), .ZN(new_n27373_));
  INV_X1     g24259(.I(new_n27200_), .ZN(new_n27374_));
  NAND4_X1   g24260(.A1(new_n27374_), .A2(pi0214), .A3(new_n27370_), .A4(new_n27193_), .ZN(new_n27375_));
  NAND2_X1   g24261(.A1(new_n27375_), .A2(new_n8247_), .ZN(new_n27376_));
  AOI21_X1   g24262(.A1(new_n27371_), .A2(new_n27373_), .B(new_n27376_), .ZN(new_n27377_));
  AOI21_X1   g24263(.A1(new_n8251_), .A2(pi0299), .B(pi0219), .ZN(new_n27378_));
  NOR2_X1    g24264(.A1(new_n27235_), .A2(new_n26704_), .ZN(new_n27379_));
  NOR4_X1    g24265(.A1(new_n27227_), .A2(pi0211), .A3(new_n27221_), .A4(new_n27224_), .ZN(new_n27380_));
  OAI21_X1   g24266(.A1(new_n27378_), .A2(new_n27379_), .B(new_n27380_), .ZN(new_n27381_));
  NAND2_X1   g24267(.A1(new_n27234_), .A2(new_n8247_), .ZN(new_n27382_));
  NAND4_X1   g24268(.A1(new_n27381_), .A2(new_n6845_), .A3(new_n27332_), .A4(new_n27382_), .ZN(new_n27383_));
  AOI21_X1   g24269(.A1(new_n27383_), .A2(pi1152), .B(new_n27325_), .ZN(new_n27384_));
  OAI21_X1   g24270(.A1(new_n27369_), .A2(new_n27377_), .B(new_n27384_), .ZN(new_n27385_));
  AND3_X2    g24271(.A1(new_n27271_), .A2(new_n8078_), .A3(new_n27264_), .Z(new_n27386_));
  NOR2_X1    g24272(.A1(new_n27198_), .A2(new_n27246_), .ZN(new_n27387_));
  NAND3_X1   g24273(.A1(new_n27278_), .A2(new_n26308_), .A3(new_n27387_), .ZN(new_n27388_));
  OAI22_X1   g24274(.A1(new_n27386_), .A2(new_n27388_), .B1(new_n27275_), .B2(pi0212), .ZN(new_n27389_));
  NOR2_X1    g24275(.A1(new_n2587_), .A2(pi0211), .ZN(new_n27390_));
  NOR2_X1    g24276(.A1(new_n27198_), .A2(new_n27390_), .ZN(new_n27391_));
  OAI21_X1   g24277(.A1(new_n26308_), .A2(new_n27391_), .B(new_n27278_), .ZN(new_n27392_));
  INV_X1     g24278(.I(new_n27392_), .ZN(new_n27393_));
  MUX2_X1    g24279(.I0(new_n27393_), .I1(new_n27389_), .S(new_n8247_), .Z(new_n27394_));
  OR3_X2     g24280(.A1(new_n27394_), .A2(po1038), .A3(new_n27356_), .Z(new_n27395_));
  OAI21_X1   g24281(.A1(new_n27387_), .A2(new_n27245_), .B(new_n8076_), .ZN(new_n27396_));
  NAND2_X1   g24282(.A1(new_n27396_), .A2(new_n8247_), .ZN(new_n27397_));
  NAND2_X1   g24283(.A1(new_n27250_), .A2(new_n27245_), .ZN(new_n27398_));
  NAND2_X1   g24284(.A1(new_n27236_), .A2(new_n26361_), .ZN(new_n27399_));
  NAND4_X1   g24285(.A1(new_n27398_), .A2(new_n27197_), .A3(new_n27397_), .A4(new_n27399_), .ZN(new_n27400_));
  AOI21_X1   g24286(.A1(pi0219), .A2(new_n27197_), .B(po1038), .ZN(new_n27401_));
  NAND4_X1   g24287(.A1(new_n27400_), .A2(new_n27250_), .A3(new_n27349_), .A4(new_n27401_), .ZN(new_n27402_));
  NAND4_X1   g24288(.A1(new_n27395_), .A2(new_n26604_), .A3(new_n27385_), .A4(new_n27402_), .ZN(new_n27403_));
  NAND2_X1   g24289(.A1(new_n27403_), .A2(new_n26374_), .ZN(new_n27404_));
  NAND4_X1   g24290(.A1(new_n27359_), .A2(new_n24753_), .A3(new_n27296_), .A4(new_n27404_), .ZN(new_n27405_));
  MUX2_X1    g24291(.I0(new_n27405_), .I1(pi0238), .S(new_n26307_), .Z(po0395));
  NOR2_X1    g24292(.A1(new_n26585_), .A2(pi0211), .ZN(new_n27407_));
  OAI21_X1   g24293(.A1(new_n27027_), .A2(new_n26585_), .B(new_n8088_), .ZN(new_n27408_));
  NAND2_X1   g24294(.A1(new_n27408_), .A2(new_n27407_), .ZN(new_n27409_));
  NOR2_X1    g24295(.A1(new_n26363_), .A2(new_n8077_), .ZN(new_n27410_));
  OAI21_X1   g24296(.A1(new_n27063_), .A2(new_n26563_), .B(new_n27410_), .ZN(new_n27411_));
  NAND2_X1   g24297(.A1(new_n27409_), .A2(new_n27411_), .ZN(new_n27412_));
  NOR2_X1    g24298(.A1(pi0212), .A2(pi0219), .ZN(new_n27413_));
  NOR2_X1    g24299(.A1(new_n27043_), .A2(new_n26634_), .ZN(new_n27414_));
  INV_X1     g24300(.I(new_n27414_), .ZN(new_n27415_));
  OAI21_X1   g24301(.A1(new_n27415_), .A2(pi0214), .B(new_n27413_), .ZN(new_n27416_));
  NOR2_X1    g24302(.A1(new_n27416_), .A2(pi0214), .ZN(new_n27417_));
  AOI21_X1   g24303(.A1(new_n27415_), .A2(pi0212), .B(po1038), .ZN(new_n27418_));
  INV_X1     g24304(.I(new_n27418_), .ZN(new_n27419_));
  NAND3_X1   g24305(.A1(new_n27414_), .A2(new_n8078_), .A3(new_n27413_), .ZN(new_n27420_));
  AOI21_X1   g24306(.A1(new_n27415_), .A2(pi0211), .B(new_n8078_), .ZN(new_n27421_));
  NAND2_X1   g24307(.A1(new_n26550_), .A2(new_n26771_), .ZN(new_n27422_));
  NAND2_X1   g24308(.A1(new_n27422_), .A2(new_n26357_), .ZN(new_n27423_));
  NAND4_X1   g24309(.A1(new_n27419_), .A2(new_n27420_), .A3(new_n27421_), .A4(new_n27423_), .ZN(new_n27424_));
  AOI21_X1   g24310(.A1(new_n27412_), .A2(new_n27417_), .B(new_n27424_), .ZN(new_n27425_));
  INV_X1     g24311(.I(new_n27410_), .ZN(new_n27426_));
  NOR2_X1    g24312(.A1(new_n27077_), .A2(new_n27129_), .ZN(new_n27427_));
  INV_X1     g24313(.I(new_n27427_), .ZN(new_n27428_));
  AOI21_X1   g24314(.A1(new_n27428_), .A2(new_n27407_), .B(new_n8078_), .ZN(new_n27429_));
  OAI21_X1   g24315(.A1(new_n27428_), .A2(pi0214), .B(new_n27413_), .ZN(new_n27430_));
  NOR4_X1    g24316(.A1(new_n27429_), .A2(new_n27430_), .A3(new_n27111_), .A4(new_n27426_), .ZN(new_n27431_));
  NAND3_X1   g24317(.A1(new_n27427_), .A2(new_n8078_), .A3(new_n27413_), .ZN(new_n27432_));
  AOI21_X1   g24318(.A1(new_n27428_), .A2(pi0212), .B(po1038), .ZN(new_n27433_));
  INV_X1     g24319(.I(new_n27433_), .ZN(new_n27434_));
  OR3_X2     g24320(.A1(new_n27111_), .A2(pi0211), .A3(new_n26356_), .Z(new_n27435_));
  NOR4_X1    g24321(.A1(new_n27428_), .A2(new_n26374_), .A3(pi0211), .A4(pi0214), .ZN(new_n27436_));
  NAND4_X1   g24322(.A1(new_n27434_), .A2(new_n27432_), .A3(new_n27435_), .A4(new_n27436_), .ZN(new_n27437_));
  NOR2_X1    g24323(.A1(new_n26822_), .A2(new_n8247_), .ZN(new_n27438_));
  NOR2_X1    g24324(.A1(new_n6845_), .A2(new_n27438_), .ZN(new_n27439_));
  OR2_X2     g24325(.A1(new_n26821_), .A2(pi0219), .Z(new_n27440_));
  NAND3_X1   g24326(.A1(new_n27439_), .A2(new_n27440_), .A3(new_n26361_), .ZN(new_n27441_));
  AOI21_X1   g24327(.A1(new_n27441_), .A2(new_n24753_), .B(new_n26374_), .ZN(new_n27442_));
  OAI21_X1   g24328(.A1(new_n27437_), .A2(new_n27431_), .B(new_n27442_), .ZN(new_n27443_));
  NOR2_X1    g24329(.A1(new_n27443_), .A2(new_n27425_), .ZN(new_n27444_));
  NAND2_X1   g24330(.A1(new_n27086_), .A2(pi0208), .ZN(new_n27445_));
  NAND2_X1   g24331(.A1(pi0299), .A2(pi1158), .ZN(new_n27446_));
  AOI21_X1   g24332(.A1(new_n26676_), .A2(new_n27446_), .B(pi0211), .ZN(new_n27447_));
  NOR3_X1    g24333(.A1(new_n8088_), .A2(new_n2587_), .A3(pi1157), .ZN(new_n27448_));
  OAI21_X1   g24334(.A1(new_n27414_), .A2(pi1157), .B(pi0211), .ZN(new_n27449_));
  OAI21_X1   g24335(.A1(new_n27449_), .A2(new_n27448_), .B(new_n8078_), .ZN(new_n27450_));
  AOI21_X1   g24336(.A1(new_n27445_), .A2(new_n27447_), .B(new_n27450_), .ZN(new_n27451_));
  NAND2_X1   g24337(.A1(new_n27428_), .A2(pi0211), .ZN(new_n27452_));
  NAND3_X1   g24338(.A1(new_n27429_), .A2(new_n27452_), .A3(new_n27432_), .ZN(new_n27453_));
  NOR2_X1    g24339(.A1(new_n27434_), .A2(new_n26374_), .ZN(new_n27454_));
  NOR3_X1    g24340(.A1(new_n8088_), .A2(new_n2587_), .A3(pi1157), .ZN(new_n27455_));
  OAI21_X1   g24341(.A1(new_n27129_), .A2(new_n27455_), .B(pi0211), .ZN(new_n27456_));
  MUX2_X1    g24342(.I0(pi1157), .I1(new_n27446_), .S(pi0208), .Z(new_n27457_));
  NOR3_X1    g24343(.A1(new_n27100_), .A2(pi0214), .A3(new_n27457_), .ZN(new_n27458_));
  NAND3_X1   g24344(.A1(new_n27456_), .A2(new_n27098_), .A3(new_n27458_), .ZN(new_n27459_));
  NAND2_X1   g24345(.A1(new_n27004_), .A2(new_n8247_), .ZN(new_n27460_));
  NAND3_X1   g24346(.A1(new_n27006_), .A2(new_n24753_), .A3(new_n27460_), .ZN(new_n27461_));
  NAND3_X1   g24347(.A1(new_n27430_), .A2(new_n27459_), .A3(new_n27461_), .ZN(new_n27462_));
  AOI21_X1   g24348(.A1(new_n27454_), .A2(new_n27453_), .B(new_n27462_), .ZN(new_n27463_));
  AOI21_X1   g24349(.A1(new_n27409_), .A2(new_n27421_), .B(new_n27420_), .ZN(new_n27464_));
  NAND2_X1   g24350(.A1(new_n27418_), .A2(new_n26374_), .ZN(new_n27465_));
  OAI21_X1   g24351(.A1(new_n27464_), .A2(new_n27465_), .B(new_n27416_), .ZN(new_n27466_));
  NOR3_X1    g24352(.A1(new_n27463_), .A2(new_n27451_), .A3(new_n27466_), .ZN(new_n27467_));
  NOR2_X1    g24353(.A1(new_n27444_), .A2(new_n27467_), .ZN(new_n27468_));
  MUX2_X1    g24354(.I0(new_n27468_), .I1(pi0239), .S(new_n26307_), .Z(po0396));
  INV_X1     g24355(.I(pi1149), .ZN(new_n27470_));
  NOR4_X1    g24356(.A1(po1038), .A2(pi0211), .A3(pi0219), .A4(new_n3414_), .ZN(new_n27471_));
  NOR2_X1    g24357(.A1(new_n8077_), .A2(new_n3258_), .ZN(new_n27472_));
  INV_X1     g24358(.I(new_n27472_), .ZN(new_n27473_));
  NOR2_X1    g24359(.A1(new_n27473_), .A2(new_n8076_), .ZN(new_n27474_));
  NOR2_X1    g24360(.A1(new_n8077_), .A2(pi1145), .ZN(new_n27475_));
  AOI21_X1   g24361(.A1(new_n8077_), .A2(new_n3258_), .B(new_n27475_), .ZN(new_n27476_));
  NAND2_X1   g24362(.A1(new_n27476_), .A2(pi0212), .ZN(new_n27477_));
  XOR2_X1    g24363(.A1(new_n27477_), .A2(new_n27473_), .Z(new_n27478_));
  NAND2_X1   g24364(.A1(new_n27478_), .A2(pi0214), .ZN(new_n27479_));
  XOR2_X1    g24365(.A1(new_n27479_), .A2(new_n27474_), .Z(new_n27480_));
  INV_X1     g24366(.I(new_n27480_), .ZN(new_n27481_));
  AOI21_X1   g24367(.A1(new_n27481_), .A2(new_n26694_), .B(new_n27471_), .ZN(new_n27482_));
  NOR2_X1    g24368(.A1(new_n27482_), .A2(pi1147), .ZN(new_n27483_));
  INV_X1     g24369(.I(new_n27483_), .ZN(new_n27484_));
  NOR3_X1    g24370(.A1(new_n27481_), .A2(po1038), .A3(new_n26998_), .ZN(new_n27485_));
  INV_X1     g24371(.I(new_n27485_), .ZN(new_n27486_));
  NOR2_X1    g24372(.A1(po1038), .A2(new_n26310_), .ZN(new_n27487_));
  NOR2_X1    g24373(.A1(new_n2587_), .A2(new_n3414_), .ZN(new_n27488_));
  INV_X1     g24374(.I(new_n27488_), .ZN(new_n27489_));
  NOR4_X1    g24375(.A1(new_n27487_), .A2(pi0211), .A3(pi0219), .A4(new_n27489_), .ZN(new_n27490_));
  INV_X1     g24376(.I(new_n27490_), .ZN(new_n27491_));
  OAI21_X1   g24377(.A1(new_n8247_), .A2(new_n27491_), .B(new_n27486_), .ZN(new_n27492_));
  NOR2_X1    g24378(.A1(new_n27492_), .A2(new_n27484_), .ZN(new_n27493_));
  INV_X1     g24379(.I(pi1147), .ZN(new_n27494_));
  NOR2_X1    g24380(.A1(new_n8447_), .A2(new_n26719_), .ZN(new_n27495_));
  INV_X1     g24381(.I(new_n27495_), .ZN(new_n27496_));
  NOR2_X1    g24382(.A1(new_n27496_), .A2(new_n6845_), .ZN(new_n27497_));
  NOR3_X1    g24383(.A1(new_n27482_), .A2(new_n27494_), .A3(new_n27497_), .ZN(new_n27498_));
  INV_X1     g24384(.I(new_n27498_), .ZN(new_n27499_));
  AOI21_X1   g24385(.A1(new_n27194_), .A2(new_n26308_), .B(pi0219), .ZN(new_n27500_));
  INV_X1     g24386(.I(new_n27500_), .ZN(new_n27501_));
  INV_X1     g24387(.I(new_n27476_), .ZN(new_n27502_));
  NOR2_X1    g24388(.A1(new_n27502_), .A2(new_n2587_), .ZN(new_n27503_));
  INV_X1     g24389(.I(new_n27503_), .ZN(new_n27504_));
  AOI21_X1   g24390(.A1(new_n27193_), .A2(new_n27504_), .B(new_n8250_), .ZN(new_n27505_));
  NOR2_X1    g24391(.A1(new_n2587_), .A2(new_n3258_), .ZN(new_n27506_));
  INV_X1     g24392(.I(new_n27506_), .ZN(new_n27507_));
  NOR2_X1    g24393(.A1(new_n27507_), .A2(new_n8077_), .ZN(new_n27508_));
  NOR2_X1    g24394(.A1(new_n27508_), .A2(new_n27390_), .ZN(new_n27509_));
  INV_X1     g24395(.I(new_n27509_), .ZN(new_n27510_));
  NOR4_X1    g24396(.A1(new_n27505_), .A2(new_n26704_), .A3(new_n27194_), .A4(new_n27510_), .ZN(new_n27511_));
  NOR2_X1    g24397(.A1(new_n27193_), .A2(po1038), .ZN(new_n27512_));
  INV_X1     g24398(.I(new_n27512_), .ZN(new_n27513_));
  AOI22_X1   g24399(.A1(new_n27491_), .A2(new_n27513_), .B1(new_n27501_), .B2(new_n27511_), .ZN(new_n27514_));
  INV_X1     g24400(.I(pi1148), .ZN(new_n27515_));
  NOR3_X1    g24401(.A1(new_n8268_), .A2(new_n8087_), .A3(new_n8088_), .ZN(new_n27516_));
  AOI21_X1   g24402(.A1(new_n26678_), .A2(new_n26450_), .B(new_n27516_), .ZN(new_n27517_));
  NAND3_X1   g24403(.A1(new_n27517_), .A2(new_n2587_), .A3(new_n27190_), .ZN(new_n27518_));
  NOR2_X1    g24404(.A1(new_n27518_), .A2(po1038), .ZN(new_n27519_));
  INV_X1     g24405(.I(new_n27519_), .ZN(new_n27520_));
  NAND2_X1   g24406(.A1(new_n27520_), .A2(new_n27515_), .ZN(new_n27521_));
  AOI21_X1   g24407(.A1(new_n27499_), .A2(new_n27514_), .B(new_n27521_), .ZN(new_n27522_));
  OAI21_X1   g24408(.A1(new_n8098_), .A2(new_n8087_), .B(new_n26431_), .ZN(new_n27523_));
  AOI21_X1   g24409(.A1(new_n27523_), .A2(pi0208), .B(pi0199), .ZN(new_n27524_));
  NOR2_X1    g24410(.A1(new_n27193_), .A2(new_n27524_), .ZN(new_n27525_));
  NOR2_X1    g24411(.A1(new_n27525_), .A2(pi0299), .ZN(new_n27526_));
  NOR2_X1    g24412(.A1(new_n27526_), .A2(pi0219), .ZN(new_n27527_));
  INV_X1     g24413(.I(new_n27246_), .ZN(new_n27528_));
  NOR2_X1    g24414(.A1(new_n27528_), .A2(pi1146), .ZN(new_n27529_));
  NOR2_X1    g24415(.A1(new_n27529_), .A2(new_n26473_), .ZN(new_n27530_));
  NOR3_X1    g24416(.A1(new_n27527_), .A2(new_n27505_), .A3(new_n27530_), .ZN(new_n27531_));
  INV_X1     g24417(.I(new_n27525_), .ZN(new_n27532_));
  NAND4_X1   g24418(.A1(new_n26693_), .A2(new_n8077_), .A3(pi0299), .A4(pi1145), .ZN(new_n27533_));
  OAI21_X1   g24419(.A1(new_n27532_), .A2(new_n26375_), .B(new_n27533_), .ZN(new_n27534_));
  OAI21_X1   g24420(.A1(new_n27531_), .A2(new_n27534_), .B(new_n6845_), .ZN(new_n27535_));
  NAND2_X1   g24421(.A1(new_n27498_), .A2(new_n27535_), .ZN(new_n27536_));
  NOR2_X1    g24422(.A1(new_n27493_), .A2(pi1148), .ZN(new_n27537_));
  AOI22_X1   g24423(.A1(new_n27537_), .A2(new_n27536_), .B1(new_n27493_), .B2(new_n27522_), .ZN(new_n27538_));
  NAND2_X1   g24424(.A1(new_n26549_), .A2(new_n8169_), .ZN(new_n27539_));
  NAND3_X1   g24425(.A1(new_n27220_), .A2(new_n2587_), .A3(new_n27539_), .ZN(new_n27540_));
  INV_X1     g24426(.I(new_n27540_), .ZN(new_n27541_));
  AOI21_X1   g24427(.A1(new_n27232_), .A2(new_n26319_), .B(new_n8247_), .ZN(new_n27542_));
  OAI21_X1   g24428(.A1(new_n27541_), .A2(new_n26319_), .B(new_n27542_), .ZN(new_n27543_));
  INV_X1     g24429(.I(new_n27543_), .ZN(new_n27544_));
  NOR2_X1    g24430(.A1(new_n27544_), .A2(po1038), .ZN(new_n27545_));
  INV_X1     g24431(.I(new_n27545_), .ZN(new_n27546_));
  NOR2_X1    g24432(.A1(new_n27546_), .A2(new_n8170_), .ZN(new_n27547_));
  NOR2_X1    g24433(.A1(new_n27547_), .A2(new_n27490_), .ZN(new_n27548_));
  NOR2_X1    g24434(.A1(new_n27232_), .A2(pi0214), .ZN(new_n27549_));
  NOR2_X1    g24435(.A1(new_n27549_), .A2(pi0212), .ZN(new_n27550_));
  INV_X1     g24436(.I(new_n27550_), .ZN(new_n27551_));
  NOR2_X1    g24437(.A1(new_n27541_), .A2(new_n8076_), .ZN(new_n27552_));
  NOR2_X1    g24438(.A1(new_n27472_), .A2(pi0214), .ZN(new_n27553_));
  AOI21_X1   g24439(.A1(new_n27502_), .A2(pi0214), .B(new_n27553_), .ZN(new_n27554_));
  NOR3_X1    g24440(.A1(new_n27552_), .A2(new_n27232_), .A3(new_n27554_), .ZN(new_n27555_));
  NOR2_X1    g24441(.A1(new_n27508_), .A2(new_n27232_), .ZN(new_n27556_));
  NOR4_X1    g24442(.A1(new_n27555_), .A2(pi0219), .A3(new_n27551_), .A4(new_n27556_), .ZN(new_n27557_));
  NOR2_X1    g24443(.A1(new_n26493_), .A2(new_n26489_), .ZN(new_n27558_));
  INV_X1     g24444(.I(new_n27558_), .ZN(new_n27559_));
  AOI21_X1   g24445(.A1(pi0219), .A2(new_n27559_), .B(po1038), .ZN(new_n27560_));
  NOR3_X1    g24446(.A1(new_n26557_), .A2(new_n8076_), .A3(new_n2587_), .ZN(new_n27561_));
  OAI21_X1   g24447(.A1(new_n27558_), .A2(pi0299), .B(pi0212), .ZN(new_n27562_));
  NOR2_X1    g24448(.A1(new_n8078_), .A2(new_n2587_), .ZN(new_n27563_));
  INV_X1     g24449(.I(new_n27563_), .ZN(new_n27564_));
  AOI21_X1   g24450(.A1(new_n27559_), .A2(new_n27564_), .B(pi0212), .ZN(new_n27565_));
  NOR2_X1    g24451(.A1(new_n27558_), .A2(new_n8077_), .ZN(new_n27566_));
  INV_X1     g24452(.I(new_n27566_), .ZN(new_n27567_));
  AOI21_X1   g24453(.A1(new_n27565_), .A2(new_n27567_), .B(pi0219), .ZN(new_n27568_));
  OAI21_X1   g24454(.A1(new_n27561_), .A2(new_n27562_), .B(new_n27568_), .ZN(new_n27569_));
  NAND2_X1   g24455(.A1(new_n27569_), .A2(new_n27560_), .ZN(new_n27570_));
  INV_X1     g24456(.I(new_n27570_), .ZN(new_n27571_));
  NOR2_X1    g24457(.A1(new_n27482_), .A2(pi1147), .ZN(new_n27573_));
  OAI21_X1   g24458(.A1(new_n27548_), .A2(new_n27557_), .B(new_n27573_), .ZN(new_n27574_));
  INV_X1     g24459(.I(new_n27267_), .ZN(new_n27575_));
  NOR2_X1    g24460(.A1(new_n26634_), .A2(pi0200), .ZN(new_n27576_));
  OAI21_X1   g24461(.A1(new_n27265_), .A2(new_n27576_), .B(new_n2587_), .ZN(new_n27577_));
  INV_X1     g24462(.I(new_n27577_), .ZN(new_n27578_));
  AOI21_X1   g24463(.A1(new_n27578_), .A2(new_n27507_), .B(new_n8077_), .ZN(new_n27579_));
  AOI21_X1   g24464(.A1(new_n8077_), .A2(new_n27575_), .B(new_n27579_), .ZN(new_n27580_));
  INV_X1     g24465(.I(new_n27580_), .ZN(new_n27581_));
  NAND2_X1   g24466(.A1(new_n8076_), .A2(new_n8078_), .ZN(new_n27582_));
  NOR2_X1    g24467(.A1(new_n27581_), .A2(new_n27582_), .ZN(new_n27583_));
  NOR2_X1    g24468(.A1(new_n27269_), .A2(pi0214), .ZN(new_n27584_));
  NOR2_X1    g24469(.A1(new_n27584_), .A2(pi0212), .ZN(new_n27585_));
  INV_X1     g24470(.I(new_n27585_), .ZN(new_n27586_));
  NOR2_X1    g24471(.A1(new_n27581_), .A2(new_n8078_), .ZN(new_n27587_));
  OAI22_X1   g24472(.A1(pi0219), .A2(new_n27583_), .B1(new_n27587_), .B2(new_n27586_), .ZN(new_n27588_));
  AOI21_X1   g24473(.A1(new_n27272_), .A2(pi0219), .B(po1038), .ZN(new_n27589_));
  INV_X1     g24474(.I(new_n27589_), .ZN(new_n27590_));
  NAND2_X1   g24475(.A1(new_n27590_), .A2(new_n27491_), .ZN(new_n27591_));
  NAND3_X1   g24476(.A1(new_n27499_), .A2(new_n27588_), .A3(new_n27591_), .ZN(new_n27592_));
  NAND2_X1   g24477(.A1(new_n11749_), .A2(new_n27208_), .ZN(new_n27593_));
  AOI21_X1   g24478(.A1(new_n27493_), .A2(new_n27593_), .B(pi1148), .ZN(new_n27594_));
  AND3_X2    g24479(.A1(new_n27594_), .A2(new_n27574_), .A3(new_n27592_), .Z(new_n27595_));
  MUX2_X1    g24480(.I0(new_n27595_), .I1(new_n27538_), .S(new_n27470_), .Z(new_n27596_));
  NOR2_X1    g24481(.A1(new_n27355_), .A2(new_n27344_), .ZN(new_n27597_));
  NOR2_X1    g24482(.A1(new_n26743_), .A2(new_n27597_), .ZN(new_n27598_));
  OAI21_X1   g24483(.A1(new_n27269_), .A2(new_n27267_), .B(pi0211), .ZN(new_n27599_));
  NOR2_X1    g24484(.A1(new_n27599_), .A2(new_n8078_), .ZN(new_n27600_));
  INV_X1     g24485(.I(new_n27600_), .ZN(new_n27601_));
  NOR2_X1    g24486(.A1(new_n27271_), .A2(new_n8078_), .ZN(new_n27602_));
  NOR2_X1    g24487(.A1(new_n27602_), .A2(new_n27586_), .ZN(new_n27603_));
  AOI21_X1   g24488(.A1(new_n27601_), .A2(new_n27271_), .B(pi0212), .ZN(new_n27604_));
  OAI21_X1   g24489(.A1(new_n27603_), .A2(pi0219), .B(new_n27604_), .ZN(new_n27605_));
  AOI21_X1   g24490(.A1(new_n8248_), .A2(new_n27601_), .B(new_n27605_), .ZN(new_n27606_));
  INV_X1     g24491(.I(new_n27413_), .ZN(new_n27607_));
  NOR3_X1    g24492(.A1(new_n27603_), .A2(new_n27271_), .A3(new_n27607_), .ZN(new_n27608_));
  NOR2_X1    g24493(.A1(new_n27608_), .A2(po1038), .ZN(new_n27609_));
  INV_X1     g24494(.I(new_n27609_), .ZN(new_n27610_));
  NOR2_X1    g24495(.A1(new_n27610_), .A2(new_n27606_), .ZN(new_n27611_));
  NOR2_X1    g24496(.A1(new_n27611_), .A2(new_n27598_), .ZN(new_n27612_));
  INV_X1     g24497(.I(new_n27593_), .ZN(new_n27613_));
  NOR2_X1    g24498(.A1(new_n11749_), .A2(pi0219), .ZN(new_n27614_));
  INV_X1     g24499(.I(new_n27614_), .ZN(new_n27615_));
  NOR2_X1    g24500(.A1(new_n27615_), .A2(new_n27345_), .ZN(new_n27616_));
  NOR2_X1    g24501(.A1(new_n27616_), .A2(new_n27613_), .ZN(new_n27617_));
  INV_X1     g24502(.I(new_n27617_), .ZN(new_n27618_));
  AOI21_X1   g24503(.A1(new_n27618_), .A2(new_n27494_), .B(pi1149), .ZN(new_n27619_));
  OAI21_X1   g24504(.A1(new_n27612_), .A2(new_n27494_), .B(new_n27619_), .ZN(new_n27620_));
  INV_X1     g24505(.I(new_n27321_), .ZN(new_n27621_));
  INV_X1     g24506(.I(new_n27390_), .ZN(new_n27622_));
  NOR3_X1    g24507(.A1(new_n27194_), .A2(new_n8078_), .A3(new_n27246_), .ZN(new_n27624_));
  AOI21_X1   g24508(.A1(pi0214), .A2(new_n27390_), .B(new_n27194_), .ZN(new_n27625_));
  INV_X1     g24509(.I(new_n27625_), .ZN(new_n27626_));
  AOI21_X1   g24510(.A1(new_n27626_), .A2(new_n8076_), .B(pi0219), .ZN(new_n27627_));
  INV_X1     g24511(.I(new_n27627_), .ZN(new_n27628_));
  NOR2_X1    g24512(.A1(new_n27628_), .A2(new_n27624_), .ZN(new_n27629_));
  INV_X1     g24513(.I(new_n27487_), .ZN(new_n27630_));
  AOI21_X1   g24514(.A1(pi0219), .A2(new_n27622_), .B(new_n27630_), .ZN(new_n27631_));
  INV_X1     g24515(.I(new_n27631_), .ZN(new_n27632_));
  AOI21_X1   g24516(.A1(new_n27513_), .A2(new_n27632_), .B(new_n27629_), .ZN(new_n27633_));
  INV_X1     g24517(.I(new_n27633_), .ZN(new_n27634_));
  NOR2_X1    g24518(.A1(new_n27634_), .A2(new_n27526_), .ZN(new_n27635_));
  NOR2_X1    g24519(.A1(new_n8080_), .A2(new_n2587_), .ZN(new_n27636_));
  NOR3_X1    g24520(.A1(new_n27194_), .A2(pi0212), .A3(new_n27636_), .ZN(new_n27637_));
  AOI21_X1   g24521(.A1(new_n27246_), .A2(new_n8078_), .B(new_n8076_), .ZN(new_n27638_));
  AOI21_X1   g24522(.A1(new_n27625_), .A2(new_n27638_), .B(new_n27637_), .ZN(new_n27639_));
  NOR2_X1    g24523(.A1(new_n27639_), .A2(new_n27526_), .ZN(new_n27640_));
  NOR2_X1    g24524(.A1(new_n27640_), .A2(pi0219), .ZN(new_n27641_));
  NAND2_X1   g24525(.A1(new_n27641_), .A2(new_n8077_), .ZN(new_n27642_));
  NAND2_X1   g24526(.A1(new_n27635_), .A2(new_n27642_), .ZN(new_n27643_));
  NAND2_X1   g24527(.A1(new_n27643_), .A2(new_n27621_), .ZN(new_n27644_));
  NAND2_X1   g24528(.A1(new_n27644_), .A2(new_n27470_), .ZN(new_n27645_));
  NAND2_X1   g24529(.A1(new_n27645_), .A2(new_n27494_), .ZN(new_n27646_));
  NAND3_X1   g24530(.A1(new_n27646_), .A2(new_n27515_), .A3(new_n27620_), .ZN(new_n27647_));
  NOR2_X1    g24531(.A1(po1038), .A2(new_n27233_), .ZN(new_n27648_));
  MUX2_X1    g24532(.I0(new_n27540_), .I1(new_n27232_), .S(pi0211), .Z(new_n27649_));
  NOR2_X1    g24533(.A1(new_n27649_), .A2(new_n8078_), .ZN(new_n27650_));
  NOR2_X1    g24534(.A1(new_n27650_), .A2(new_n8076_), .ZN(new_n27651_));
  NOR2_X1    g24535(.A1(new_n27540_), .A2(new_n8078_), .ZN(new_n27652_));
  AOI21_X1   g24536(.A1(new_n27652_), .A2(new_n27551_), .B(pi0219), .ZN(new_n27653_));
  NAND3_X1   g24537(.A1(new_n27651_), .A2(new_n27540_), .A3(new_n27653_), .ZN(new_n27654_));
  OAI21_X1   g24538(.A1(new_n27401_), .A2(new_n27648_), .B(new_n27654_), .ZN(new_n27655_));
  OR2_X2     g24539(.A1(new_n27655_), .A2(new_n27317_), .Z(new_n27656_));
  NOR2_X1    g24540(.A1(new_n26308_), .A2(new_n2587_), .ZN(new_n27657_));
  INV_X1     g24541(.I(new_n27657_), .ZN(new_n27658_));
  NOR2_X1    g24542(.A1(new_n27630_), .A2(new_n27658_), .ZN(new_n27659_));
  NOR2_X1    g24543(.A1(new_n8077_), .A2(new_n8247_), .ZN(new_n27660_));
  INV_X1     g24544(.I(new_n27660_), .ZN(new_n27661_));
  NOR3_X1    g24545(.A1(po1038), .A2(new_n26308_), .A3(new_n27661_), .ZN(new_n27662_));
  NOR2_X1    g24546(.A1(new_n6845_), .A2(new_n27558_), .ZN(new_n27663_));
  NOR3_X1    g24547(.A1(new_n27659_), .A2(new_n27662_), .A3(new_n27663_), .ZN(new_n27664_));
  NAND4_X1   g24548(.A1(new_n27656_), .A2(pi1147), .A3(new_n27470_), .A4(new_n27664_), .ZN(new_n27665_));
  XOR2_X1    g24549(.A1(pi0211), .A2(pi0212), .Z(new_n27666_));
  XOR2_X1    g24550(.A1(new_n27666_), .A2(new_n8078_), .Z(new_n27667_));
  AOI21_X1   g24551(.A1(new_n27347_), .A2(new_n26558_), .B(new_n27667_), .ZN(new_n27668_));
  INV_X1     g24552(.I(new_n27518_), .ZN(new_n27669_));
  NOR2_X1    g24553(.A1(new_n27669_), .A2(new_n27636_), .ZN(new_n27670_));
  INV_X1     g24554(.I(new_n27670_), .ZN(new_n27671_));
  AOI21_X1   g24555(.A1(new_n27671_), .A2(new_n8076_), .B(pi0219), .ZN(new_n27672_));
  INV_X1     g24556(.I(new_n27672_), .ZN(new_n27673_));
  NAND2_X1   g24557(.A1(new_n27517_), .A2(new_n2587_), .ZN(new_n27674_));
  INV_X1     g24558(.I(new_n27674_), .ZN(new_n27675_));
  NOR2_X1    g24559(.A1(new_n27675_), .A2(new_n8078_), .ZN(new_n27676_));
  AOI21_X1   g24560(.A1(new_n27518_), .A2(new_n27528_), .B(pi0212), .ZN(new_n27677_));
  NAND2_X1   g24561(.A1(new_n27676_), .A2(new_n27677_), .ZN(new_n27678_));
  INV_X1     g24562(.I(new_n27678_), .ZN(new_n27679_));
  INV_X1     g24563(.I(new_n27676_), .ZN(new_n27680_));
  AOI21_X1   g24564(.A1(new_n27669_), .A2(new_n8078_), .B(pi0212), .ZN(new_n27681_));
  NOR2_X1    g24565(.A1(new_n27675_), .A2(pi0211), .ZN(new_n27682_));
  NOR2_X1    g24566(.A1(new_n27682_), .A2(new_n27669_), .ZN(new_n27683_));
  NOR2_X1    g24567(.A1(new_n27683_), .A2(new_n26362_), .ZN(new_n27684_));
  INV_X1     g24568(.I(new_n27684_), .ZN(new_n27685_));
  NOR2_X1    g24569(.A1(new_n27675_), .A2(pi0214), .ZN(new_n27686_));
  OAI22_X1   g24570(.A1(new_n27685_), .A2(new_n27686_), .B1(new_n27680_), .B2(new_n27681_), .ZN(new_n27687_));
  AOI21_X1   g24571(.A1(new_n27687_), .A2(new_n27679_), .B(new_n27673_), .ZN(new_n27688_));
  AOI21_X1   g24572(.A1(new_n27518_), .A2(pi0219), .B(po1038), .ZN(new_n27689_));
  INV_X1     g24573(.I(new_n27689_), .ZN(new_n27690_));
  NOR2_X1    g24574(.A1(new_n27688_), .A2(new_n27690_), .ZN(new_n27691_));
  NOR2_X1    g24575(.A1(new_n27691_), .A2(new_n27668_), .ZN(new_n27692_));
  INV_X1     g24576(.I(new_n27692_), .ZN(new_n27693_));
  NAND2_X1   g24577(.A1(new_n27693_), .A2(pi1147), .ZN(new_n27694_));
  INV_X1     g24578(.I(new_n27659_), .ZN(new_n27695_));
  NAND2_X1   g24579(.A1(new_n26342_), .A2(pi0211), .ZN(new_n27696_));
  NAND3_X1   g24580(.A1(new_n27696_), .A2(new_n8250_), .A3(new_n8247_), .ZN(new_n27697_));
  AOI21_X1   g24581(.A1(new_n27695_), .A2(new_n26743_), .B(new_n27697_), .ZN(new_n27698_));
  NOR2_X1    g24582(.A1(new_n27698_), .A2(new_n27512_), .ZN(new_n27699_));
  INV_X1     g24583(.I(new_n27699_), .ZN(new_n27700_));
  NAND2_X1   g24584(.A1(new_n27700_), .A2(pi1147), .ZN(new_n27701_));
  NAND4_X1   g24585(.A1(new_n27694_), .A2(new_n27470_), .A3(new_n27665_), .A4(new_n27701_), .ZN(new_n27702_));
  NAND2_X1   g24586(.A1(new_n27702_), .A2(pi1148), .ZN(new_n27703_));
  XNOR2_X1   g24587(.A1(new_n27647_), .A2(new_n27703_), .ZN(new_n27704_));
  MUX2_X1    g24588(.I0(new_n27704_), .I1(new_n27596_), .S(new_n24753_), .Z(new_n27705_));
  NOR2_X1    g24589(.A1(new_n3258_), .A2(pi0199), .ZN(new_n27706_));
  INV_X1     g24590(.I(new_n27706_), .ZN(new_n27707_));
  AOI21_X1   g24591(.A1(new_n27707_), .A2(pi0200), .B(pi0299), .ZN(new_n27708_));
  INV_X1     g24592(.I(new_n27708_), .ZN(new_n27709_));
  AOI21_X1   g24593(.A1(new_n8098_), .A2(new_n3414_), .B(pi0199), .ZN(new_n27710_));
  NAND2_X1   g24594(.A1(new_n27709_), .A2(new_n27710_), .ZN(new_n27711_));
  AOI21_X1   g24595(.A1(pi0199), .A2(pi1145), .B(pi0200), .ZN(new_n27712_));
  NOR2_X1    g24596(.A1(new_n3414_), .A2(pi0199), .ZN(new_n27713_));
  NOR2_X1    g24597(.A1(new_n27713_), .A2(new_n8098_), .ZN(new_n27714_));
  NOR4_X1    g24598(.A1(new_n27714_), .A2(new_n27707_), .A3(new_n26328_), .A4(new_n27712_), .ZN(new_n27715_));
  NOR2_X1    g24599(.A1(new_n27711_), .A2(new_n26504_), .ZN(new_n27716_));
  OAI21_X1   g24600(.A1(new_n27506_), .A2(new_n27715_), .B(new_n27716_), .ZN(new_n27717_));
  OAI21_X1   g24601(.A1(new_n26634_), .A2(new_n27711_), .B(new_n27717_), .ZN(new_n27718_));
  NOR2_X1    g24602(.A1(new_n27718_), .A2(pi0299), .ZN(new_n27719_));
  INV_X1     g24603(.I(new_n27719_), .ZN(new_n27720_));
  NOR2_X1    g24604(.A1(new_n27715_), .A2(new_n26678_), .ZN(new_n27721_));
  AOI21_X1   g24605(.A1(new_n27711_), .A2(new_n8090_), .B(new_n27721_), .ZN(new_n27722_));
  NAND4_X1   g24606(.A1(new_n27720_), .A2(new_n8077_), .A3(new_n8247_), .A4(new_n26342_), .ZN(new_n27723_));
  NAND2_X1   g24607(.A1(new_n27723_), .A2(new_n6845_), .ZN(new_n27724_));
  NAND2_X1   g24608(.A1(new_n27720_), .A2(pi0211), .ZN(new_n27725_));
  INV_X1     g24609(.I(new_n27711_), .ZN(new_n27726_));
  NAND4_X1   g24610(.A1(new_n27717_), .A2(new_n8087_), .A3(new_n27712_), .A4(new_n27726_), .ZN(new_n27727_));
  INV_X1     g24611(.I(new_n27712_), .ZN(new_n27728_));
  NAND3_X1   g24612(.A1(new_n27708_), .A2(new_n26549_), .A3(new_n27728_), .ZN(new_n27729_));
  NAND2_X1   g24613(.A1(new_n27727_), .A2(new_n27729_), .ZN(new_n27730_));
  INV_X1     g24614(.I(new_n27730_), .ZN(new_n27731_));
  NOR2_X1    g24615(.A1(new_n27731_), .A2(pi0299), .ZN(new_n27732_));
  INV_X1     g24616(.I(new_n27732_), .ZN(new_n27733_));
  NAND2_X1   g24617(.A1(new_n27733_), .A2(pi0214), .ZN(new_n27734_));
  AOI21_X1   g24618(.A1(new_n27734_), .A2(new_n27725_), .B(new_n8076_), .ZN(new_n27735_));
  NOR2_X1    g24619(.A1(new_n27719_), .A2(new_n8080_), .ZN(new_n27736_));
  NOR4_X1    g24620(.A1(new_n27735_), .A2(pi0219), .A3(new_n27722_), .A4(new_n27736_), .ZN(new_n27737_));
  NAND2_X1   g24621(.A1(new_n27737_), .A2(new_n27724_), .ZN(new_n27738_));
  INV_X1     g24622(.I(new_n27738_), .ZN(new_n27739_));
  NOR2_X1    g24623(.A1(new_n26743_), .A2(new_n27697_), .ZN(new_n27740_));
  OAI21_X1   g24624(.A1(new_n27739_), .A2(new_n27740_), .B(new_n27494_), .ZN(new_n27741_));
  AOI21_X1   g24625(.A1(new_n27708_), .A2(new_n27728_), .B(new_n8089_), .ZN(new_n27742_));
  NOR2_X1    g24626(.A1(new_n27721_), .A2(new_n27742_), .ZN(new_n27743_));
  NAND3_X1   g24627(.A1(new_n27732_), .A2(new_n8078_), .A3(new_n27743_), .ZN(new_n27744_));
  OAI21_X1   g24628(.A1(pi0214), .A2(new_n27743_), .B(new_n27733_), .ZN(new_n27745_));
  INV_X1     g24629(.I(new_n27722_), .ZN(new_n27746_));
  OAI21_X1   g24630(.A1(new_n27719_), .A2(pi0211), .B(new_n27746_), .ZN(new_n27747_));
  NAND2_X1   g24631(.A1(new_n27747_), .A2(new_n8078_), .ZN(new_n27748_));
  NAND3_X1   g24632(.A1(new_n27733_), .A2(new_n27748_), .A3(pi0212), .ZN(new_n27749_));
  NAND4_X1   g24633(.A1(new_n27745_), .A2(new_n8076_), .A3(new_n27749_), .A4(new_n27744_), .ZN(new_n27750_));
  AND3_X2    g24634(.A1(new_n27750_), .A2(pi0219), .A3(new_n27743_), .Z(new_n27751_));
  INV_X1     g24635(.I(new_n27743_), .ZN(new_n27752_));
  AOI21_X1   g24636(.A1(pi0219), .A2(new_n27752_), .B(new_n27750_), .ZN(new_n27753_));
  OAI21_X1   g24637(.A1(new_n27751_), .A2(new_n27753_), .B(new_n6845_), .ZN(new_n27754_));
  NAND4_X1   g24638(.A1(new_n27754_), .A2(new_n26308_), .A3(new_n27737_), .A4(new_n27743_), .ZN(new_n27755_));
  NOR2_X1    g24639(.A1(new_n27668_), .A2(pi1147), .ZN(new_n27756_));
  AOI22_X1   g24640(.A1(new_n27755_), .A2(new_n27756_), .B1(new_n27470_), .B2(new_n27741_), .ZN(new_n27757_));
  NOR2_X1    g24641(.A1(new_n27317_), .A2(pi1147), .ZN(new_n27758_));
  INV_X1     g24642(.I(new_n27724_), .ZN(new_n27759_));
  NOR3_X1    g24643(.A1(new_n27722_), .A2(pi0219), .A3(new_n27657_), .ZN(new_n27760_));
  NOR2_X1    g24644(.A1(new_n27759_), .A2(new_n27760_), .ZN(new_n27761_));
  NOR2_X1    g24645(.A1(pi1147), .A2(pi1149), .ZN(new_n27762_));
  OAI21_X1   g24646(.A1(new_n27761_), .A2(new_n27662_), .B(new_n27762_), .ZN(new_n27763_));
  AOI21_X1   g24647(.A1(new_n27754_), .A2(new_n27758_), .B(new_n27763_), .ZN(new_n27764_));
  NOR2_X1    g24648(.A1(new_n27757_), .A2(new_n27764_), .ZN(new_n27765_));
  NAND2_X1   g24649(.A1(new_n27743_), .A2(new_n6845_), .ZN(new_n27766_));
  OAI21_X1   g24650(.A1(new_n27747_), .A2(pi0214), .B(pi0212), .ZN(new_n27767_));
  NAND2_X1   g24651(.A1(new_n27725_), .A2(new_n27746_), .ZN(new_n27768_));
  NAND3_X1   g24652(.A1(new_n27768_), .A2(new_n8078_), .A3(new_n27767_), .ZN(new_n27769_));
  NOR2_X1    g24653(.A1(new_n27719_), .A2(pi0211), .ZN(new_n27770_));
  NAND2_X1   g24654(.A1(new_n27770_), .A2(pi0214), .ZN(new_n27771_));
  AOI21_X1   g24655(.A1(new_n27771_), .A2(new_n27746_), .B(pi0212), .ZN(new_n27772_));
  NOR2_X1    g24656(.A1(new_n27772_), .A2(pi0219), .ZN(new_n27773_));
  NAND2_X1   g24657(.A1(new_n27773_), .A2(new_n27769_), .ZN(new_n27774_));
  AOI21_X1   g24658(.A1(new_n27739_), .A2(new_n27774_), .B(new_n27321_), .ZN(new_n27775_));
  NOR2_X1    g24659(.A1(new_n27766_), .A2(pi1147), .ZN(new_n27776_));
  NOR2_X1    g24660(.A1(new_n27766_), .A2(pi1147), .ZN(new_n27777_));
  NOR3_X1    g24661(.A1(new_n27775_), .A2(new_n27494_), .A3(new_n27777_), .ZN(new_n27778_));
  NOR3_X1    g24662(.A1(new_n27778_), .A2(pi1149), .A3(new_n27776_), .ZN(new_n27779_));
  AOI21_X1   g24663(.A1(new_n27773_), .A2(new_n27769_), .B(new_n27759_), .ZN(new_n27780_));
  OAI21_X1   g24664(.A1(new_n27780_), .A2(new_n27598_), .B(pi1147), .ZN(new_n27781_));
  NAND2_X1   g24665(.A1(new_n27766_), .A2(new_n27496_), .ZN(new_n27782_));
  INV_X1     g24666(.I(new_n11749_), .ZN(new_n27783_));
  NOR2_X1    g24667(.A1(new_n27783_), .A2(new_n27496_), .ZN(new_n27784_));
  AOI22_X1   g24668(.A1(new_n27730_), .A2(new_n27784_), .B1(new_n27494_), .B2(new_n27782_), .ZN(new_n27785_));
  AOI21_X1   g24669(.A1(new_n27781_), .A2(new_n27785_), .B(new_n27470_), .ZN(new_n27786_));
  OAI21_X1   g24670(.A1(new_n27786_), .A2(pi1148), .B(new_n24753_), .ZN(new_n27787_));
  OAI21_X1   g24671(.A1(new_n27779_), .A2(new_n27787_), .B(new_n27515_), .ZN(new_n27788_));
  AOI21_X1   g24672(.A1(new_n27752_), .A2(new_n8078_), .B(pi0212), .ZN(new_n27789_));
  INV_X1     g24673(.I(new_n27508_), .ZN(new_n27790_));
  NAND2_X1   g24674(.A1(new_n27752_), .A2(new_n27790_), .ZN(new_n27791_));
  AOI21_X1   g24675(.A1(new_n27789_), .A2(new_n27791_), .B(pi0219), .ZN(new_n27792_));
  NOR2_X1    g24676(.A1(new_n27730_), .A2(pi0299), .ZN(new_n27793_));
  INV_X1     g24677(.I(new_n27793_), .ZN(new_n27794_));
  NOR3_X1    g24678(.A1(new_n27503_), .A2(pi0212), .A3(new_n8078_), .ZN(new_n27795_));
  NAND3_X1   g24679(.A1(new_n27794_), .A2(new_n27792_), .A3(new_n27795_), .ZN(new_n27796_));
  NAND3_X1   g24680(.A1(new_n27794_), .A2(new_n8077_), .A3(new_n27489_), .ZN(new_n27797_));
  OAI21_X1   g24681(.A1(new_n27752_), .A2(new_n26342_), .B(pi0219), .ZN(new_n27798_));
  AOI21_X1   g24682(.A1(new_n27752_), .A2(pi0211), .B(new_n26308_), .ZN(new_n27799_));
  NAND3_X1   g24683(.A1(new_n27797_), .A2(new_n27798_), .A3(new_n27799_), .ZN(new_n27800_));
  NAND4_X1   g24684(.A1(new_n27800_), .A2(new_n6845_), .A3(new_n27483_), .A4(new_n27796_), .ZN(new_n27801_));
  NAND2_X1   g24685(.A1(new_n27509_), .A2(new_n26308_), .ZN(new_n27802_));
  OAI21_X1   g24686(.A1(new_n27718_), .A2(new_n27802_), .B(new_n27792_), .ZN(new_n27803_));
  NOR3_X1    g24687(.A1(new_n27718_), .A2(new_n8078_), .A3(new_n27503_), .ZN(new_n27804_));
  NOR2_X1    g24688(.A1(new_n2587_), .A2(pi1145), .ZN(new_n27805_));
  OAI22_X1   g24689(.A1(new_n27725_), .A2(new_n27805_), .B1(new_n27736_), .B2(new_n27804_), .ZN(new_n27806_));
  NOR3_X1    g24690(.A1(new_n27806_), .A2(new_n27772_), .A3(new_n27803_), .ZN(new_n27807_));
  AOI21_X1   g24691(.A1(new_n27722_), .A2(new_n26319_), .B(new_n8247_), .ZN(new_n27808_));
  NOR3_X1    g24692(.A1(new_n27808_), .A2(new_n26308_), .A3(new_n27805_), .ZN(new_n27809_));
  AOI21_X1   g24693(.A1(new_n27770_), .A2(new_n27809_), .B(po1038), .ZN(new_n27810_));
  NAND2_X1   g24694(.A1(new_n27498_), .A2(new_n27810_), .ZN(new_n27811_));
  OAI21_X1   g24695(.A1(new_n27807_), .A2(new_n27811_), .B(new_n27801_), .ZN(new_n27812_));
  AOI21_X1   g24696(.A1(new_n27812_), .A2(new_n24753_), .B(pi0209), .ZN(new_n27813_));
  OAI21_X1   g24697(.A1(new_n27788_), .A2(new_n27765_), .B(new_n27813_), .ZN(new_n27814_));
  AOI21_X1   g24698(.A1(new_n27705_), .A2(pi0209), .B(new_n27814_), .ZN(new_n27815_));
  MUX2_X1    g24699(.I0(new_n27815_), .I1(pi0240), .S(new_n26307_), .Z(po0397));
  INV_X1     g24700(.I(pi1150), .ZN(new_n27817_));
  INV_X1     g24701(.I(new_n27230_), .ZN(new_n27818_));
  NOR2_X1    g24702(.A1(new_n27818_), .A2(new_n26604_), .ZN(new_n27819_));
  AOI21_X1   g24703(.A1(po1038), .A2(new_n27496_), .B(new_n27251_), .ZN(new_n27820_));
  NAND4_X1   g24704(.A1(new_n27361_), .A2(new_n26604_), .A3(new_n27241_), .A4(new_n27495_), .ZN(new_n27821_));
  NAND2_X1   g24705(.A1(new_n27821_), .A2(new_n6845_), .ZN(new_n27822_));
  AOI22_X1   g24706(.A1(new_n27822_), .A2(new_n27820_), .B1(new_n27234_), .B2(new_n27819_), .ZN(new_n27823_));
  INV_X1     g24707(.I(new_n27820_), .ZN(new_n27824_));
  NOR2_X1    g24708(.A1(new_n27345_), .A2(new_n26998_), .ZN(new_n27825_));
  INV_X1     g24709(.I(new_n27825_), .ZN(new_n27826_));
  AOI21_X1   g24710(.A1(new_n27278_), .A2(new_n27826_), .B(new_n27824_), .ZN(new_n27827_));
  NOR2_X1    g24711(.A1(new_n27818_), .A2(new_n27199_), .ZN(new_n27828_));
  OAI21_X1   g24712(.A1(new_n27827_), .A2(new_n27828_), .B(new_n26604_), .ZN(new_n27829_));
  NOR2_X1    g24713(.A1(new_n27823_), .A2(new_n27829_), .ZN(new_n27830_));
  NOR2_X1    g24714(.A1(new_n27277_), .A2(pi0299), .ZN(new_n27831_));
  AOI21_X1   g24715(.A1(new_n27267_), .A2(new_n8078_), .B(new_n8076_), .ZN(new_n27832_));
  OAI21_X1   g24716(.A1(new_n27271_), .A2(new_n8078_), .B(new_n27832_), .ZN(new_n27833_));
  NAND3_X1   g24717(.A1(new_n27272_), .A2(pi0219), .A3(pi1152), .ZN(new_n27835_));
  AOI21_X1   g24718(.A1(new_n27241_), .A2(new_n8078_), .B(pi0212), .ZN(new_n27836_));
  OAI21_X1   g24719(.A1(new_n27364_), .A2(new_n8078_), .B(new_n27836_), .ZN(new_n27837_));
  AOI21_X1   g24720(.A1(new_n27374_), .A2(new_n27372_), .B(pi0219), .ZN(new_n27838_));
  NOR2_X1    g24721(.A1(new_n27838_), .A2(pi1152), .ZN(new_n27839_));
  NAND2_X1   g24722(.A1(new_n27839_), .A2(new_n27837_), .ZN(new_n27840_));
  NOR2_X1    g24723(.A1(new_n27317_), .A2(new_n27251_), .ZN(new_n27841_));
  INV_X1     g24724(.I(new_n27841_), .ZN(new_n27842_));
  AOI21_X1   g24725(.A1(new_n27199_), .A2(pi0219), .B(po1038), .ZN(new_n27843_));
  INV_X1     g24726(.I(new_n27843_), .ZN(new_n27844_));
  NAND2_X1   g24727(.A1(new_n27844_), .A2(new_n27513_), .ZN(new_n27845_));
  NAND4_X1   g24728(.A1(new_n27840_), .A2(new_n27835_), .A3(new_n27842_), .A4(new_n27845_), .ZN(new_n27846_));
  NOR2_X1    g24729(.A1(new_n27209_), .A2(pi0212), .ZN(new_n27847_));
  INV_X1     g24730(.I(new_n27847_), .ZN(new_n27848_));
  NOR2_X1    g24731(.A1(new_n27848_), .A2(new_n27245_), .ZN(new_n27849_));
  AOI21_X1   g24732(.A1(new_n27849_), .A2(new_n27622_), .B(pi0219), .ZN(new_n27850_));
  INV_X1     g24733(.I(new_n27850_), .ZN(new_n27851_));
  INV_X1     g24734(.I(new_n27245_), .ZN(new_n27852_));
  NOR4_X1    g24735(.A1(new_n27852_), .A2(new_n27209_), .A3(pi0211), .A4(pi0212), .ZN(new_n27853_));
  NOR3_X1    g24736(.A1(new_n27853_), .A2(new_n8078_), .A3(new_n27247_), .ZN(new_n27854_));
  NOR2_X1    g24737(.A1(new_n27851_), .A2(new_n27854_), .ZN(new_n27855_));
  AOI21_X1   g24738(.A1(new_n2587_), .A2(new_n27199_), .B(new_n27397_), .ZN(new_n27856_));
  NOR2_X1    g24739(.A1(new_n27856_), .A2(new_n27855_), .ZN(new_n27857_));
  OAI21_X1   g24740(.A1(new_n27857_), .A2(new_n27844_), .B(new_n26604_), .ZN(new_n27858_));
  INV_X1     g24741(.I(new_n27858_), .ZN(new_n27859_));
  OAI21_X1   g24742(.A1(new_n27857_), .A2(pi0219), .B(new_n27235_), .ZN(new_n27860_));
  AOI21_X1   g24743(.A1(new_n27860_), .A2(new_n6845_), .B(new_n26604_), .ZN(new_n27861_));
  NOR2_X1    g24744(.A1(new_n27668_), .A2(pi1151), .ZN(new_n27862_));
  OAI21_X1   g24745(.A1(new_n27861_), .A2(new_n27859_), .B(new_n27862_), .ZN(new_n27863_));
  NAND2_X1   g24746(.A1(new_n27863_), .A2(new_n27846_), .ZN(new_n27864_));
  OAI21_X1   g24747(.A1(new_n27864_), .A2(new_n27817_), .B(new_n27830_), .ZN(new_n27865_));
  INV_X1     g24748(.I(new_n27830_), .ZN(new_n27866_));
  NAND3_X1   g24749(.A1(new_n27864_), .A2(pi1150), .A3(new_n27866_), .ZN(new_n27867_));
  NAND3_X1   g24750(.A1(new_n27865_), .A2(new_n27867_), .A3(new_n27470_), .ZN(new_n27868_));
  NOR2_X1    g24751(.A1(new_n27631_), .A2(new_n27843_), .ZN(new_n27869_));
  INV_X1     g24752(.I(new_n27869_), .ZN(new_n27870_));
  AOI21_X1   g24753(.A1(new_n27235_), .A2(pi0219), .B(po1038), .ZN(new_n27871_));
  NOR2_X1    g24754(.A1(new_n27870_), .A2(new_n27871_), .ZN(new_n27872_));
  NOR3_X1    g24755(.A1(new_n27872_), .A2(new_n8247_), .A3(pi1152), .ZN(new_n27873_));
  AOI21_X1   g24756(.A1(new_n27199_), .A2(new_n27397_), .B(new_n27869_), .ZN(new_n27874_));
  NOR2_X1    g24757(.A1(new_n27858_), .A2(new_n27874_), .ZN(new_n27875_));
  NOR2_X1    g24758(.A1(new_n27740_), .A2(pi1151), .ZN(new_n27876_));
  OAI21_X1   g24759(.A1(new_n27875_), .A2(new_n27873_), .B(new_n27876_), .ZN(new_n27877_));
  INV_X1     g24760(.I(new_n27369_), .ZN(new_n27878_));
  NOR2_X1    g24761(.A1(new_n27662_), .A2(new_n27251_), .ZN(new_n27879_));
  AOI21_X1   g24762(.A1(new_n27278_), .A2(new_n26308_), .B(new_n27831_), .ZN(new_n27880_));
  NOR2_X1    g24763(.A1(po1038), .A2(pi1152), .ZN(new_n27881_));
  OAI21_X1   g24764(.A1(new_n27393_), .A2(pi0219), .B(new_n27881_), .ZN(new_n27882_));
  OAI21_X1   g24765(.A1(new_n27880_), .A2(pi0219), .B(new_n27882_), .ZN(new_n27883_));
  NAND4_X1   g24766(.A1(new_n27838_), .A2(pi0212), .A3(new_n26604_), .A4(new_n27241_), .ZN(new_n27884_));
  AOI21_X1   g24767(.A1(new_n27883_), .A2(new_n27879_), .B(new_n27884_), .ZN(new_n27885_));
  NAND2_X1   g24768(.A1(new_n27885_), .A2(new_n27878_), .ZN(new_n27886_));
  AOI21_X1   g24769(.A1(pi1150), .A2(new_n27877_), .B(new_n27886_), .ZN(new_n27887_));
  NAND2_X1   g24770(.A1(new_n27241_), .A2(new_n27180_), .ZN(new_n27888_));
  NAND4_X1   g24771(.A1(new_n27367_), .A2(pi0212), .A3(new_n27360_), .A4(new_n27888_), .ZN(new_n27889_));
  NAND2_X1   g24772(.A1(new_n27889_), .A2(new_n8247_), .ZN(new_n27890_));
  AOI21_X1   g24773(.A1(new_n27278_), .A2(new_n27391_), .B(pi0214), .ZN(new_n27891_));
  NOR4_X1    g24774(.A1(new_n27392_), .A2(new_n27891_), .A3(new_n27388_), .A4(pi0212), .ZN(new_n27892_));
  OR2_X2     g24775(.A1(new_n27892_), .A2(pi0219), .Z(new_n27893_));
  NOR2_X1    g24776(.A1(new_n27598_), .A2(new_n27251_), .ZN(new_n27894_));
  INV_X1     g24777(.I(new_n27894_), .ZN(new_n27895_));
  NAND3_X1   g24778(.A1(new_n27893_), .A2(new_n27882_), .A3(new_n27895_), .ZN(new_n27896_));
  NAND4_X1   g24779(.A1(new_n27896_), .A2(pi1152), .A3(new_n27878_), .A4(new_n27890_), .ZN(new_n27897_));
  INV_X1     g24780(.I(new_n27872_), .ZN(new_n27898_));
  NAND4_X1   g24781(.A1(new_n27898_), .A2(new_n26604_), .A3(new_n27235_), .A4(new_n27397_), .ZN(new_n27899_));
  AND3_X2    g24782(.A1(new_n27874_), .A2(new_n26604_), .A3(new_n27323_), .Z(new_n27900_));
  AOI21_X1   g24783(.A1(new_n27899_), .A2(new_n27900_), .B(pi1150), .ZN(new_n27901_));
  NAND2_X1   g24784(.A1(new_n27897_), .A2(new_n27901_), .ZN(new_n27902_));
  OAI21_X1   g24785(.A1(new_n27887_), .A2(new_n27902_), .B(pi1149), .ZN(new_n27903_));
  AND2_X2    g24786(.A1(new_n27868_), .A2(new_n27903_), .Z(new_n27904_));
  OAI21_X1   g24787(.A1(new_n27868_), .A2(new_n27903_), .B(pi0213), .ZN(new_n27905_));
  NAND2_X1   g24788(.A1(new_n27403_), .A2(pi0213), .ZN(new_n27906_));
  OAI21_X1   g24789(.A1(new_n27904_), .A2(new_n27905_), .B(new_n27906_), .ZN(new_n27907_));
  AOI21_X1   g24790(.A1(new_n27575_), .A2(new_n26529_), .B(pi0211), .ZN(new_n27908_));
  OAI22_X1   g24791(.A1(new_n27600_), .A2(new_n8250_), .B1(new_n27270_), .B2(new_n27908_), .ZN(new_n27909_));
  AOI21_X1   g24792(.A1(new_n27601_), .A2(pi0212), .B(new_n27585_), .ZN(new_n27910_));
  INV_X1     g24793(.I(new_n27910_), .ZN(new_n27911_));
  AOI21_X1   g24794(.A1(new_n27911_), .A2(new_n27909_), .B(pi0219), .ZN(new_n27912_));
  NOR3_X1    g24795(.A1(new_n27610_), .A2(new_n27356_), .A3(new_n27912_), .ZN(new_n27913_));
  INV_X1     g24796(.I(new_n27913_), .ZN(new_n27914_));
  NOR2_X1    g24797(.A1(new_n27600_), .A2(new_n27584_), .ZN(new_n27915_));
  OAI22_X1   g24798(.A1(new_n27525_), .A2(new_n27657_), .B1(new_n26411_), .B2(new_n27313_), .ZN(new_n27916_));
  NAND2_X1   g24799(.A1(new_n27916_), .A2(new_n8247_), .ZN(new_n27917_));
  NOR2_X1    g24800(.A1(new_n27332_), .A2(pi1152), .ZN(new_n27918_));
  AOI21_X1   g24801(.A1(new_n27532_), .A2(pi0219), .B(po1038), .ZN(new_n27919_));
  NAND3_X1   g24802(.A1(new_n27918_), .A2(new_n27917_), .A3(new_n27919_), .ZN(new_n27920_));
  INV_X1     g24803(.I(new_n27920_), .ZN(new_n27921_));
  INV_X1     g24804(.I(new_n27561_), .ZN(new_n27922_));
  NAND3_X1   g24805(.A1(new_n27325_), .A2(new_n8247_), .A3(new_n27922_), .ZN(new_n27923_));
  NOR4_X1    g24806(.A1(new_n27923_), .A2(new_n27921_), .A3(new_n27275_), .A4(new_n27915_), .ZN(new_n27924_));
  NAND2_X1   g24807(.A1(new_n27924_), .A2(new_n27609_), .ZN(new_n27925_));
  AOI21_X1   g24808(.A1(new_n27532_), .A2(new_n27826_), .B(po1038), .ZN(new_n27926_));
  NOR2_X1    g24809(.A1(new_n26737_), .A2(new_n2587_), .ZN(new_n27927_));
  NOR2_X1    g24810(.A1(new_n27348_), .A2(new_n27927_), .ZN(new_n27928_));
  NOR2_X1    g24811(.A1(pi1150), .A2(pi1152), .ZN(new_n27929_));
  INV_X1     g24812(.I(new_n27929_), .ZN(new_n27930_));
  AOI21_X1   g24813(.A1(new_n27926_), .A2(new_n27928_), .B(new_n27930_), .ZN(new_n27931_));
  AND3_X2    g24814(.A1(new_n27914_), .A2(new_n27925_), .A3(new_n27931_), .Z(new_n27932_));
  INV_X1     g24815(.I(new_n27932_), .ZN(new_n27933_));
  NOR2_X1    g24816(.A1(new_n27558_), .A2(pi0219), .ZN(new_n27934_));
  NAND3_X1   g24817(.A1(new_n27934_), .A2(new_n8077_), .A3(new_n27922_), .ZN(new_n27935_));
  NOR2_X1    g24818(.A1(po1038), .A2(new_n27559_), .ZN(new_n27936_));
  OAI21_X1   g24819(.A1(new_n27659_), .A2(new_n27936_), .B(new_n27935_), .ZN(new_n27937_));
  INV_X1     g24820(.I(new_n8081_), .ZN(new_n27938_));
  NOR2_X1    g24821(.A1(new_n27938_), .A2(new_n2587_), .ZN(new_n27939_));
  NOR2_X1    g24822(.A1(new_n27939_), .A2(pi0219), .ZN(new_n27940_));
  INV_X1     g24823(.I(new_n27940_), .ZN(new_n27941_));
  NOR2_X1    g24824(.A1(new_n27632_), .A2(new_n27941_), .ZN(new_n27942_));
  NOR2_X1    g24825(.A1(new_n27571_), .A2(new_n27942_), .ZN(new_n27943_));
  AOI21_X1   g24826(.A1(new_n11893_), .A2(new_n27922_), .B(new_n27934_), .ZN(new_n27944_));
  NOR2_X1    g24827(.A1(new_n27943_), .A2(new_n27944_), .ZN(new_n27945_));
  AOI21_X1   g24828(.A1(new_n27193_), .A2(new_n27622_), .B(new_n8250_), .ZN(new_n27946_));
  NOR2_X1    g24829(.A1(new_n26650_), .A2(new_n27927_), .ZN(new_n27947_));
  OAI21_X1   g24830(.A1(new_n27193_), .A2(new_n2587_), .B(new_n27947_), .ZN(new_n27948_));
  NOR3_X1    g24831(.A1(new_n27501_), .A2(new_n27948_), .A3(new_n27946_), .ZN(new_n27949_));
  AOI21_X1   g24832(.A1(new_n27193_), .A2(pi0219), .B(po1038), .ZN(new_n27950_));
  NAND2_X1   g24833(.A1(new_n27918_), .A2(new_n27950_), .ZN(new_n27951_));
  OAI21_X1   g24834(.A1(new_n27951_), .A2(new_n27949_), .B(new_n27325_), .ZN(new_n27952_));
  AOI21_X1   g24835(.A1(new_n27945_), .A2(new_n27937_), .B(new_n27952_), .ZN(new_n27953_));
  INV_X1     g24836(.I(new_n27953_), .ZN(new_n27954_));
  NAND2_X1   g24837(.A1(new_n27825_), .A2(pi1153), .ZN(new_n27955_));
  OAI21_X1   g24838(.A1(new_n27348_), .A2(new_n27955_), .B(new_n26604_), .ZN(new_n27956_));
  INV_X1     g24839(.I(new_n27956_), .ZN(new_n27957_));
  NOR2_X1    g24840(.A1(new_n27512_), .A2(pi1151), .ZN(new_n27958_));
  NOR2_X1    g24841(.A1(new_n27958_), .A2(pi1152), .ZN(new_n27959_));
  INV_X1     g24842(.I(new_n27959_), .ZN(new_n27960_));
  NAND4_X1   g24843(.A1(new_n27945_), .A2(new_n27356_), .A3(new_n27957_), .A4(new_n27960_), .ZN(new_n27961_));
  NOR2_X1    g24844(.A1(pi1149), .A2(pi1150), .ZN(new_n27962_));
  INV_X1     g24845(.I(new_n27962_), .ZN(new_n27963_));
  AOI21_X1   g24846(.A1(new_n27954_), .A2(new_n27961_), .B(new_n27963_), .ZN(new_n27964_));
  AOI21_X1   g24847(.A1(new_n27249_), .A2(pi0219), .B(po1038), .ZN(new_n27965_));
  NAND2_X1   g24848(.A1(new_n27400_), .A2(new_n27965_), .ZN(new_n27966_));
  INV_X1     g24849(.I(new_n27356_), .ZN(new_n27967_));
  NOR2_X1    g24850(.A1(new_n27956_), .A2(new_n27967_), .ZN(new_n27968_));
  AOI21_X1   g24851(.A1(new_n27966_), .A2(new_n27968_), .B(pi1150), .ZN(new_n27969_));
  INV_X1     g24852(.I(new_n27853_), .ZN(new_n27970_));
  INV_X1     g24853(.I(new_n27965_), .ZN(new_n27971_));
  AOI21_X1   g24854(.A1(new_n27850_), .A2(new_n27970_), .B(new_n27971_), .ZN(new_n27972_));
  INV_X1     g24855(.I(new_n27972_), .ZN(new_n27973_));
  INV_X1     g24856(.I(new_n27332_), .ZN(new_n27974_));
  NOR4_X1    g24857(.A1(new_n27314_), .A2(new_n2587_), .A3(pi1152), .A4(new_n27316_), .ZN(new_n27975_));
  AOI21_X1   g24858(.A1(new_n27974_), .A2(new_n27975_), .B(new_n27324_), .ZN(new_n27976_));
  INV_X1     g24859(.I(new_n27976_), .ZN(new_n27977_));
  AOI21_X1   g24860(.A1(new_n27966_), .A2(new_n27973_), .B(new_n27977_), .ZN(new_n27978_));
  OAI21_X1   g24861(.A1(new_n27978_), .A2(new_n27969_), .B(new_n27470_), .ZN(new_n27979_));
  NOR2_X1    g24862(.A1(new_n27675_), .A2(new_n27927_), .ZN(new_n27980_));
  INV_X1     g24863(.I(new_n27980_), .ZN(new_n27981_));
  NOR3_X1    g24864(.A1(new_n27981_), .A2(new_n8078_), .A3(new_n27681_), .ZN(new_n27982_));
  NAND3_X1   g24865(.A1(new_n27685_), .A2(new_n8078_), .A3(new_n27980_), .ZN(new_n27983_));
  NAND2_X1   g24866(.A1(new_n27983_), .A2(new_n8247_), .ZN(new_n27984_));
  NOR2_X1    g24867(.A1(new_n27332_), .A2(new_n27690_), .ZN(new_n27985_));
  OAI21_X1   g24868(.A1(new_n27984_), .A2(new_n27982_), .B(new_n27985_), .ZN(new_n27986_));
  OAI21_X1   g24869(.A1(new_n8626_), .A2(new_n26457_), .B(new_n27220_), .ZN(new_n27987_));
  NAND3_X1   g24870(.A1(new_n27987_), .A2(new_n8077_), .A3(new_n26529_), .ZN(new_n27988_));
  INV_X1     g24871(.I(new_n27988_), .ZN(new_n27989_));
  NOR2_X1    g24872(.A1(new_n27541_), .A2(new_n8077_), .ZN(new_n27990_));
  NOR2_X1    g24873(.A1(new_n27989_), .A2(new_n27990_), .ZN(new_n27991_));
  INV_X1     g24874(.I(new_n27991_), .ZN(new_n27992_));
  NOR2_X1    g24875(.A1(new_n27992_), .A2(new_n8078_), .ZN(new_n27993_));
  INV_X1     g24876(.I(new_n27993_), .ZN(new_n27994_));
  OR3_X2     g24877(.A1(new_n27992_), .A2(pi0214), .A3(new_n27552_), .Z(new_n27995_));
  NOR2_X1    g24878(.A1(new_n27551_), .A2(pi0219), .ZN(new_n27996_));
  NAND4_X1   g24879(.A1(new_n27995_), .A2(new_n27994_), .A3(new_n27546_), .A4(new_n27996_), .ZN(new_n27997_));
  AND4_X2    g24880(.A1(new_n26604_), .A2(new_n27997_), .A3(new_n27324_), .A4(new_n27986_), .Z(new_n27998_));
  NOR2_X1    g24881(.A1(new_n27518_), .A2(new_n27350_), .ZN(new_n27999_));
  INV_X1     g24882(.I(new_n27999_), .ZN(new_n28000_));
  AOI21_X1   g24883(.A1(new_n27674_), .A2(new_n26529_), .B(pi0211), .ZN(new_n28001_));
  INV_X1     g24884(.I(new_n28001_), .ZN(new_n28002_));
  NOR2_X1    g24885(.A1(new_n27683_), .A2(new_n27352_), .ZN(new_n28003_));
  NAND2_X1   g24886(.A1(new_n28003_), .A2(new_n28002_), .ZN(new_n28004_));
  AOI21_X1   g24887(.A1(new_n28004_), .A2(new_n28000_), .B(po1038), .ZN(new_n28005_));
  NOR4_X1    g24888(.A1(new_n27990_), .A2(pi0212), .A3(new_n8078_), .A4(new_n27232_), .ZN(new_n28007_));
  NOR2_X1    g24889(.A1(new_n27992_), .A2(new_n28007_), .ZN(new_n28008_));
  NOR2_X1    g24890(.A1(new_n27233_), .A2(new_n8077_), .ZN(new_n28009_));
  OAI21_X1   g24891(.A1(new_n27989_), .A2(new_n28009_), .B(new_n27550_), .ZN(new_n28010_));
  NAND4_X1   g24892(.A1(new_n27545_), .A2(new_n8247_), .A3(new_n28010_), .A4(new_n27967_), .ZN(new_n28011_));
  NOR2_X1    g24893(.A1(new_n27349_), .A2(new_n27930_), .ZN(new_n28012_));
  OAI21_X1   g24894(.A1(new_n28011_), .A2(new_n28008_), .B(new_n28012_), .ZN(new_n28013_));
  NOR3_X1    g24895(.A1(new_n27998_), .A2(new_n28005_), .A3(new_n28013_), .ZN(new_n28014_));
  AOI22_X1   g24896(.A1(new_n27933_), .A2(new_n27964_), .B1(new_n27979_), .B2(new_n28014_), .ZN(new_n28015_));
  NOR2_X1    g24897(.A1(new_n27693_), .A2(pi1151), .ZN(new_n28016_));
  NOR2_X1    g24898(.A1(new_n27655_), .A2(new_n27842_), .ZN(new_n28017_));
  NOR2_X1    g24899(.A1(new_n28016_), .A2(new_n28017_), .ZN(new_n28018_));
  OAI21_X1   g24900(.A1(new_n27617_), .A2(pi1150), .B(new_n27251_), .ZN(new_n28019_));
  NAND2_X1   g24901(.A1(new_n28019_), .A2(new_n27962_), .ZN(new_n28020_));
  NOR2_X1    g24902(.A1(new_n27611_), .A2(new_n27895_), .ZN(new_n28021_));
  NAND2_X1   g24903(.A1(new_n27643_), .A2(new_n27322_), .ZN(new_n28022_));
  NAND2_X1   g24904(.A1(new_n28022_), .A2(new_n27817_), .ZN(new_n28023_));
  INV_X1     g24905(.I(new_n27879_), .ZN(new_n28024_));
  NAND3_X1   g24906(.A1(new_n27695_), .A2(new_n27663_), .A3(new_n28024_), .ZN(new_n28025_));
  NAND3_X1   g24907(.A1(new_n28025_), .A2(new_n27817_), .A3(new_n27251_), .ZN(new_n28026_));
  OAI22_X1   g24908(.A1(new_n28023_), .A2(new_n28021_), .B1(new_n27699_), .B2(new_n28026_), .ZN(new_n28027_));
  INV_X1     g24909(.I(new_n28027_), .ZN(new_n28028_));
  OAI22_X1   g24910(.A1(new_n28028_), .A2(pi1149), .B1(new_n28018_), .B2(new_n28020_), .ZN(new_n28029_));
  INV_X1     g24911(.I(new_n28029_), .ZN(new_n28030_));
  OR3_X2     g24912(.A1(new_n28030_), .A2(pi0213), .A3(new_n28015_), .Z(new_n28031_));
  OAI21_X1   g24913(.A1(new_n28029_), .A2(pi0213), .B(new_n28015_), .ZN(new_n28032_));
  NAND3_X1   g24914(.A1(new_n28031_), .A2(new_n26374_), .A3(new_n28032_), .ZN(new_n28033_));
  AOI21_X1   g24915(.A1(pi0209), .A2(new_n27907_), .B(new_n28033_), .ZN(new_n28034_));
  MUX2_X1    g24916(.I0(new_n28034_), .I1(pi0241), .S(new_n26307_), .Z(po0398));
  NAND3_X1   g24917(.A1(new_n26345_), .A2(pi0212), .A3(pi0214), .ZN(new_n28036_));
  AOI21_X1   g24918(.A1(pi0199), .A2(pi1144), .B(pi0200), .ZN(new_n28037_));
  NOR2_X1    g24919(.A1(new_n27707_), .A2(new_n28037_), .ZN(new_n28038_));
  NOR3_X1    g24920(.A1(new_n28038_), .A2(pi0299), .A3(new_n27714_), .ZN(new_n28039_));
  NOR2_X1    g24921(.A1(new_n28039_), .A2(new_n26634_), .ZN(new_n28040_));
  INV_X1     g24922(.I(new_n28040_), .ZN(new_n28041_));
  OAI21_X1   g24923(.A1(new_n2587_), .A2(new_n26347_), .B(new_n26704_), .ZN(new_n28042_));
  NAND4_X1   g24924(.A1(new_n28041_), .A2(new_n8247_), .A3(new_n28042_), .A4(new_n28036_), .ZN(new_n28043_));
  NOR2_X1    g24925(.A1(new_n28039_), .A2(new_n26677_), .ZN(new_n28044_));
  OAI21_X1   g24926(.A1(new_n26342_), .A2(new_n28044_), .B(new_n28043_), .ZN(new_n28045_));
  NAND3_X1   g24927(.A1(new_n28041_), .A2(new_n26309_), .A3(new_n26442_), .ZN(new_n28046_));
  OAI21_X1   g24928(.A1(new_n28039_), .A2(new_n26677_), .B(pi0211), .ZN(new_n28047_));
  NAND4_X1   g24929(.A1(new_n28045_), .A2(pi0219), .A3(new_n28046_), .A4(new_n28047_), .ZN(new_n28048_));
  OR2_X2     g24930(.A1(new_n26318_), .A2(pi0213), .Z(new_n28049_));
  NAND2_X1   g24931(.A1(new_n28039_), .A2(pi0207), .ZN(new_n28050_));
  INV_X1     g24932(.I(new_n28037_), .ZN(new_n28051_));
  AOI21_X1   g24933(.A1(new_n26324_), .A2(new_n8098_), .B(pi0299), .ZN(new_n28052_));
  NAND4_X1   g24934(.A1(new_n28052_), .A2(pi0207), .A3(new_n27713_), .A4(new_n28051_), .ZN(new_n28053_));
  AOI21_X1   g24935(.A1(new_n28050_), .A2(new_n28053_), .B(new_n8088_), .ZN(new_n28054_));
  INV_X1     g24936(.I(new_n28054_), .ZN(new_n28055_));
  NAND4_X1   g24937(.A1(new_n28048_), .A2(new_n6845_), .A3(new_n28049_), .A4(new_n28055_), .ZN(new_n28056_));
  NOR2_X1    g24938(.A1(new_n26981_), .A2(new_n8078_), .ZN(new_n28057_));
  AOI21_X1   g24939(.A1(new_n27502_), .A2(new_n8078_), .B(new_n28057_), .ZN(new_n28058_));
  NAND2_X1   g24940(.A1(new_n27476_), .A2(pi0214), .ZN(new_n28059_));
  NOR3_X1    g24941(.A1(new_n28058_), .A2(pi0212), .A3(new_n28059_), .ZN(new_n28060_));
  INV_X1     g24942(.I(new_n28058_), .ZN(new_n28061_));
  AOI21_X1   g24943(.A1(new_n8076_), .A2(new_n28059_), .B(new_n28061_), .ZN(new_n28062_));
  NOR3_X1    g24944(.A1(new_n28062_), .A2(pi0219), .A3(new_n28060_), .ZN(new_n28063_));
  OAI21_X1   g24945(.A1(new_n2552_), .A2(pi0211), .B(pi0219), .ZN(new_n28064_));
  NAND3_X1   g24946(.A1(new_n28063_), .A2(new_n26311_), .A3(new_n28064_), .ZN(new_n28065_));
  NOR2_X1    g24947(.A1(new_n28054_), .A2(new_n28040_), .ZN(new_n28066_));
  INV_X1     g24948(.I(new_n28066_), .ZN(new_n28067_));
  NOR2_X1    g24949(.A1(new_n28067_), .A2(new_n27506_), .ZN(new_n28068_));
  NOR2_X1    g24950(.A1(new_n28067_), .A2(new_n27488_), .ZN(new_n28069_));
  INV_X1     g24951(.I(new_n28069_), .ZN(new_n28070_));
  NOR2_X1    g24952(.A1(new_n28070_), .A2(new_n8077_), .ZN(new_n28071_));
  AOI21_X1   g24953(.A1(new_n8077_), .A2(new_n28068_), .B(new_n28071_), .ZN(new_n28072_));
  NOR2_X1    g24954(.A1(new_n28054_), .A2(new_n28044_), .ZN(new_n28073_));
  INV_X1     g24955(.I(new_n28073_), .ZN(new_n28074_));
  NOR2_X1    g24956(.A1(new_n28074_), .A2(pi0214), .ZN(new_n28075_));
  NOR2_X1    g24957(.A1(new_n28075_), .A2(pi0212), .ZN(new_n28076_));
  NOR3_X1    g24958(.A1(new_n28072_), .A2(new_n8078_), .A3(new_n28076_), .ZN(new_n28077_));
  NOR2_X1    g24959(.A1(new_n28077_), .A2(pi0219), .ZN(new_n28078_));
  NAND3_X1   g24960(.A1(new_n28055_), .A2(new_n26480_), .A3(new_n28041_), .ZN(new_n28079_));
  NOR3_X1    g24961(.A1(new_n28072_), .A2(pi0212), .A3(pi0214), .ZN(new_n28081_));
  AOI21_X1   g24962(.A1(new_n28074_), .A2(new_n26319_), .B(new_n8247_), .ZN(new_n28082_));
  NOR3_X1    g24963(.A1(new_n28082_), .A2(new_n26319_), .A3(new_n28079_), .ZN(new_n28083_));
  OR3_X2     g24964(.A1(new_n28081_), .A2(po1038), .A3(new_n28083_), .Z(new_n28084_));
  OAI21_X1   g24965(.A1(new_n28084_), .A2(new_n28078_), .B(new_n28065_), .ZN(new_n28085_));
  NAND2_X1   g24966(.A1(new_n28085_), .A2(pi0213), .ZN(new_n28086_));
  AOI21_X1   g24967(.A1(new_n28086_), .A2(new_n28056_), .B(new_n26374_), .ZN(new_n28087_));
  NAND2_X1   g24968(.A1(new_n26308_), .A2(pi0219), .ZN(new_n28088_));
  AND4_X2    g24969(.A1(new_n2587_), .A2(new_n28063_), .A3(new_n28064_), .A4(new_n28088_), .Z(new_n28089_));
  NAND2_X1   g24970(.A1(new_n26339_), .A2(new_n11749_), .ZN(new_n28090_));
  OAI21_X1   g24971(.A1(new_n28090_), .A2(new_n28089_), .B(new_n28065_), .ZN(new_n28091_));
  MUX2_X1    g24972(.I0(new_n28091_), .I1(new_n26354_), .S(new_n24753_), .Z(new_n28092_));
  AOI21_X1   g24973(.A1(new_n28092_), .A2(new_n26374_), .B(new_n28087_), .ZN(new_n28093_));
  MUX2_X1    g24974(.I0(new_n28093_), .I1(pi0242), .S(new_n26307_), .Z(po0399));
  INV_X1     g24975(.I(pi0273), .ZN(new_n28095_));
  INV_X1     g24976(.I(pi0271), .ZN(new_n28096_));
  INV_X1     g24977(.I(pi0802), .ZN(new_n28097_));
  NOR2_X1    g24978(.A1(new_n3272_), .A2(new_n28097_), .ZN(new_n28098_));
  INV_X1     g24979(.I(new_n28098_), .ZN(new_n28099_));
  NOR2_X1    g24980(.A1(pi0083), .A2(pi0085), .ZN(new_n28100_));
  NOR2_X1    g24981(.A1(new_n28100_), .A2(new_n5276_), .ZN(new_n28101_));
  INV_X1     g24982(.I(new_n28101_), .ZN(new_n28102_));
  NOR2_X1    g24983(.A1(new_n28102_), .A2(new_n28099_), .ZN(new_n28103_));
  INV_X1     g24984(.I(new_n28103_), .ZN(new_n28104_));
  NOR2_X1    g24985(.A1(new_n28104_), .A2(new_n28096_), .ZN(new_n28105_));
  INV_X1     g24986(.I(new_n28105_), .ZN(new_n28106_));
  AOI21_X1   g24987(.A1(new_n28106_), .A2(new_n2918_), .B(new_n28095_), .ZN(new_n28107_));
  NOR2_X1    g24988(.A1(new_n28107_), .A2(pi1091), .ZN(new_n28108_));
  NOR2_X1    g24989(.A1(new_n28108_), .A2(new_n8094_), .ZN(new_n28109_));
  NAND2_X1   g24990(.A1(new_n28100_), .A2(new_n2441_), .ZN(new_n28110_));
  NAND2_X1   g24991(.A1(new_n28110_), .A2(pi0314), .ZN(new_n28111_));
  NOR2_X1    g24992(.A1(new_n28111_), .A2(new_n28099_), .ZN(new_n28112_));
  NAND2_X1   g24993(.A1(new_n28112_), .A2(new_n2918_), .ZN(new_n28113_));
  INV_X1     g24994(.I(new_n28113_), .ZN(new_n28114_));
  NOR2_X1    g24995(.A1(new_n28113_), .A2(new_n28096_), .ZN(new_n28115_));
  NAND2_X1   g24996(.A1(new_n28115_), .A2(pi0273), .ZN(new_n28116_));
  INV_X1     g24997(.I(new_n28116_), .ZN(new_n28117_));
  NOR2_X1    g24998(.A1(new_n28117_), .A2(new_n28107_), .ZN(new_n28118_));
  NAND2_X1   g24999(.A1(new_n28118_), .A2(new_n2918_), .ZN(new_n28119_));
  INV_X1     g25000(.I(new_n28119_), .ZN(new_n28120_));
  NOR2_X1    g25001(.A1(new_n28120_), .A2(pi0199), .ZN(new_n28121_));
  NOR2_X1    g25002(.A1(new_n28121_), .A2(new_n28109_), .ZN(new_n28122_));
  INV_X1     g25003(.I(new_n28122_), .ZN(new_n28123_));
  AOI21_X1   g25004(.A1(new_n28123_), .A2(new_n28114_), .B(pi0299), .ZN(new_n28124_));
  INV_X1     g25005(.I(new_n28124_), .ZN(new_n28125_));
  NOR2_X1    g25006(.A1(new_n28125_), .A2(new_n28109_), .ZN(new_n28126_));
  INV_X1     g25007(.I(new_n28126_), .ZN(new_n28127_));
  NOR2_X1    g25008(.A1(new_n28108_), .A2(pi0200), .ZN(new_n28128_));
  NOR2_X1    g25009(.A1(new_n28127_), .A2(new_n28128_), .ZN(new_n28129_));
  INV_X1     g25010(.I(new_n28129_), .ZN(new_n28130_));
  NOR2_X1    g25011(.A1(new_n28114_), .A2(pi0200), .ZN(new_n28131_));
  INV_X1     g25012(.I(new_n28131_), .ZN(new_n28132_));
  AOI21_X1   g25013(.A1(new_n28123_), .A2(new_n28132_), .B(pi0299), .ZN(new_n28133_));
  INV_X1     g25014(.I(new_n28133_), .ZN(new_n28134_));
  NOR2_X1    g25015(.A1(new_n28117_), .A2(new_n2587_), .ZN(new_n28135_));
  NOR2_X1    g25016(.A1(new_n28134_), .A2(new_n28135_), .ZN(new_n28136_));
  INV_X1     g25017(.I(new_n28136_), .ZN(new_n28137_));
  NOR2_X1    g25018(.A1(new_n28137_), .A2(pi0243), .ZN(new_n28138_));
  NOR2_X1    g25019(.A1(new_n28125_), .A2(new_n28128_), .ZN(new_n28139_));
  INV_X1     g25020(.I(new_n28108_), .ZN(new_n28140_));
  NOR2_X1    g25021(.A1(new_n28140_), .A2(new_n2587_), .ZN(new_n28141_));
  NOR2_X1    g25022(.A1(new_n28139_), .A2(new_n28141_), .ZN(new_n28142_));
  NOR2_X1    g25023(.A1(new_n28133_), .A2(new_n28109_), .ZN(new_n28143_));
  NOR2_X1    g25024(.A1(new_n28104_), .A2(pi1091), .ZN(new_n28144_));
  INV_X1     g25025(.I(new_n28144_), .ZN(new_n28145_));
  NOR3_X1    g25026(.A1(new_n28145_), .A2(new_n28096_), .A3(new_n28095_), .ZN(new_n28146_));
  NOR2_X1    g25027(.A1(new_n28146_), .A2(new_n2587_), .ZN(new_n28147_));
  INV_X1     g25028(.I(new_n28139_), .ZN(new_n28148_));
  NOR2_X1    g25029(.A1(new_n28148_), .A2(new_n28121_), .ZN(new_n28149_));
  NOR2_X1    g25030(.A1(new_n28149_), .A2(new_n28147_), .ZN(new_n28150_));
  INV_X1     g25031(.I(new_n28150_), .ZN(new_n28151_));
  NOR2_X1    g25032(.A1(new_n28151_), .A2(new_n28143_), .ZN(new_n28152_));
  NOR2_X1    g25033(.A1(pi0243), .A2(pi1155), .ZN(new_n28153_));
  OAI21_X1   g25034(.A1(new_n28152_), .A2(new_n28142_), .B(new_n28153_), .ZN(new_n28154_));
  INV_X1     g25035(.I(new_n28135_), .ZN(new_n28155_));
  NOR2_X1    g25036(.A1(new_n28155_), .A2(new_n28140_), .ZN(new_n28156_));
  NOR2_X1    g25037(.A1(new_n28149_), .A2(new_n28156_), .ZN(new_n28157_));
  INV_X1     g25038(.I(new_n28157_), .ZN(new_n28158_));
  NOR2_X1    g25039(.A1(new_n28158_), .A2(new_n11912_), .ZN(new_n28159_));
  INV_X1     g25040(.I(new_n28159_), .ZN(new_n28160_));
  AOI22_X1   g25041(.A1(new_n28154_), .A2(new_n28160_), .B1(new_n28130_), .B2(new_n28138_), .ZN(new_n28161_));
  NOR2_X1    g25042(.A1(new_n28161_), .A2(new_n11912_), .ZN(new_n28162_));
  INV_X1     g25043(.I(pi0243), .ZN(new_n28163_));
  NOR2_X1    g25044(.A1(new_n28163_), .A2(pi1091), .ZN(new_n28164_));
  INV_X1     g25045(.I(new_n28164_), .ZN(new_n28165_));
  NOR2_X1    g25046(.A1(new_n28129_), .A2(new_n28135_), .ZN(new_n28166_));
  INV_X1     g25047(.I(new_n28166_), .ZN(new_n28167_));
  AOI21_X1   g25048(.A1(new_n28167_), .A2(new_n28165_), .B(pi1156), .ZN(new_n28168_));
  NAND2_X1   g25049(.A1(new_n28162_), .A2(new_n28168_), .ZN(new_n28169_));
  NAND2_X1   g25050(.A1(new_n28148_), .A2(new_n28155_), .ZN(new_n28170_));
  NOR3_X1    g25051(.A1(new_n28170_), .A2(new_n28126_), .A3(new_n28163_), .ZN(new_n28171_));
  NOR2_X1    g25052(.A1(new_n28133_), .A2(new_n28121_), .ZN(new_n28172_));
  NOR2_X1    g25053(.A1(new_n28172_), .A2(new_n28141_), .ZN(new_n28173_));
  INV_X1     g25054(.I(new_n28173_), .ZN(new_n28174_));
  NOR2_X1    g25055(.A1(new_n28124_), .A2(new_n28135_), .ZN(new_n28175_));
  NOR2_X1    g25056(.A1(new_n28175_), .A2(pi0243), .ZN(new_n28176_));
  AOI21_X1   g25057(.A1(new_n28174_), .A2(new_n28176_), .B(pi1155), .ZN(new_n28177_));
  NOR2_X1    g25058(.A1(new_n28171_), .A2(new_n28177_), .ZN(new_n28178_));
  NOR2_X1    g25059(.A1(new_n28134_), .A2(new_n28156_), .ZN(new_n28179_));
  INV_X1     g25060(.I(new_n28179_), .ZN(new_n28180_));
  NOR2_X1    g25061(.A1(new_n28163_), .A2(new_n11912_), .ZN(new_n28181_));
  NAND3_X1   g25062(.A1(new_n28180_), .A2(new_n28163_), .A3(new_n28181_), .ZN(new_n28182_));
  NOR2_X1    g25063(.A1(new_n28182_), .A2(new_n28170_), .ZN(new_n28183_));
  NOR4_X1    g25064(.A1(new_n28178_), .A2(pi1156), .A3(pi1157), .A4(new_n28183_), .ZN(new_n28184_));
  NOR4_X1    g25065(.A1(new_n28108_), .A2(new_n8094_), .A3(new_n11912_), .A4(new_n28164_), .ZN(new_n28185_));
  NOR2_X1    g25066(.A1(new_n28124_), .A2(new_n28147_), .ZN(new_n28186_));
  INV_X1     g25067(.I(new_n28186_), .ZN(new_n28187_));
  NAND3_X1   g25068(.A1(new_n28187_), .A2(new_n28163_), .A3(new_n2918_), .ZN(new_n28188_));
  INV_X1     g25069(.I(new_n28175_), .ZN(new_n28189_));
  OAI21_X1   g25070(.A1(new_n28189_), .A2(new_n28163_), .B(new_n26486_), .ZN(new_n28190_));
  AOI21_X1   g25071(.A1(new_n28175_), .A2(new_n28188_), .B(new_n28190_), .ZN(new_n28191_));
  OAI21_X1   g25072(.A1(new_n28183_), .A2(new_n28185_), .B(new_n28191_), .ZN(new_n28192_));
  NOR2_X1    g25073(.A1(new_n28125_), .A2(new_n28121_), .ZN(new_n28193_));
  NOR2_X1    g25074(.A1(new_n28193_), .A2(new_n28156_), .ZN(new_n28194_));
  NOR2_X1    g25075(.A1(new_n28126_), .A2(new_n28135_), .ZN(new_n28195_));
  NOR2_X1    g25076(.A1(new_n28195_), .A2(pi0243), .ZN(new_n28196_));
  AOI21_X1   g25077(.A1(pi0243), .A2(new_n28194_), .B(new_n28196_), .ZN(new_n28197_));
  NOR3_X1    g25078(.A1(new_n28170_), .A2(pi1155), .A3(new_n28114_), .ZN(new_n28198_));
  OR3_X2     g25079(.A1(new_n28197_), .A2(new_n12026_), .A3(new_n28198_), .Z(new_n28199_));
  NAND4_X1   g25080(.A1(new_n28199_), .A2(pi0211), .A3(new_n12049_), .A4(new_n28192_), .ZN(new_n28200_));
  AOI21_X1   g25081(.A1(new_n28169_), .A2(new_n28184_), .B(new_n28200_), .ZN(new_n28201_));
  NOR2_X1    g25082(.A1(new_n28139_), .A2(new_n28156_), .ZN(new_n28202_));
  AOI21_X1   g25083(.A1(new_n11912_), .A2(new_n28137_), .B(new_n28202_), .ZN(new_n28203_));
  NAND2_X1   g25084(.A1(new_n28199_), .A2(new_n28203_), .ZN(new_n28204_));
  NOR2_X1    g25085(.A1(new_n28136_), .A2(pi0243), .ZN(new_n28205_));
  AOI21_X1   g25086(.A1(pi0243), .A2(new_n28202_), .B(new_n28205_), .ZN(new_n28206_));
  NOR4_X1    g25087(.A1(new_n28197_), .A2(new_n28206_), .A3(new_n28191_), .A4(pi1155), .ZN(new_n28207_));
  NOR2_X1    g25088(.A1(new_n28207_), .A2(pi1157), .ZN(new_n28208_));
  AOI21_X1   g25089(.A1(new_n28204_), .A2(new_n28208_), .B(pi0211), .ZN(new_n28209_));
  OR3_X2     g25090(.A1(new_n28162_), .A2(new_n12026_), .A3(pi1157), .Z(new_n28210_));
  OAI21_X1   g25091(.A1(new_n28210_), .A2(new_n28209_), .B(new_n8247_), .ZN(new_n28211_));
  NOR2_X1    g25092(.A1(new_n28211_), .A2(new_n28201_), .ZN(new_n28212_));
  NAND2_X1   g25093(.A1(pi0211), .A2(pi1157), .ZN(new_n28213_));
  NOR2_X1    g25094(.A1(new_n28173_), .A2(pi0243), .ZN(new_n28214_));
  NOR2_X1    g25095(.A1(new_n28139_), .A2(new_n28147_), .ZN(new_n28215_));
  INV_X1     g25096(.I(new_n28215_), .ZN(new_n28216_));
  NOR4_X1    g25097(.A1(new_n28216_), .A2(new_n28179_), .A3(new_n28163_), .A4(pi1155), .ZN(new_n28217_));
  NOR2_X1    g25098(.A1(new_n28216_), .A2(new_n28126_), .ZN(new_n28218_));
  INV_X1     g25099(.I(new_n28218_), .ZN(new_n28219_));
  NOR2_X1    g25100(.A1(new_n28219_), .A2(new_n28163_), .ZN(new_n28220_));
  OAI21_X1   g25101(.A1(new_n28214_), .A2(new_n28217_), .B(new_n28220_), .ZN(new_n28221_));
  AOI21_X1   g25102(.A1(new_n28221_), .A2(new_n12026_), .B(new_n28213_), .ZN(new_n28222_));
  NAND2_X1   g25103(.A1(new_n28152_), .A2(pi0243), .ZN(new_n28223_));
  NOR2_X1    g25104(.A1(new_n28129_), .A2(new_n28141_), .ZN(new_n28224_));
  OAI21_X1   g25105(.A1(pi0243), .A2(new_n28224_), .B(new_n28223_), .ZN(new_n28225_));
  OAI22_X1   g25106(.A1(new_n28151_), .A2(new_n28182_), .B1(pi1155), .B2(new_n28214_), .ZN(new_n28226_));
  OAI21_X1   g25107(.A1(new_n28225_), .A2(new_n28226_), .B(pi1156), .ZN(new_n28227_));
  NOR2_X1    g25108(.A1(new_n28186_), .A2(new_n28164_), .ZN(new_n28228_));
  XOR2_X1    g25109(.A1(new_n28228_), .A2(new_n28163_), .Z(new_n28229_));
  NAND2_X1   g25110(.A1(new_n28229_), .A2(new_n11912_), .ZN(new_n28230_));
  NOR2_X1    g25111(.A1(new_n28143_), .A2(new_n28141_), .ZN(new_n28231_));
  INV_X1     g25112(.I(new_n28231_), .ZN(new_n28232_));
  NAND2_X1   g25113(.A1(new_n28232_), .A2(new_n28163_), .ZN(new_n28233_));
  NOR2_X1    g25114(.A1(new_n28193_), .A2(new_n28163_), .ZN(new_n28234_));
  AOI21_X1   g25115(.A1(new_n28215_), .A2(new_n28234_), .B(new_n11912_), .ZN(new_n28235_));
  AOI21_X1   g25116(.A1(new_n28235_), .A2(new_n28233_), .B(pi1156), .ZN(new_n28236_));
  AOI21_X1   g25117(.A1(new_n28230_), .A2(new_n28236_), .B(pi1157), .ZN(new_n28237_));
  NOR2_X1    g25118(.A1(new_n28126_), .A2(new_n28141_), .ZN(new_n28238_));
  OAI21_X1   g25119(.A1(new_n28198_), .A2(new_n28238_), .B(new_n28163_), .ZN(new_n28239_));
  NOR2_X1    g25120(.A1(new_n28193_), .A2(new_n28147_), .ZN(new_n28240_));
  INV_X1     g25121(.I(new_n28240_), .ZN(new_n28241_));
  NOR2_X1    g25122(.A1(new_n28133_), .A2(pi1155), .ZN(new_n28242_));
  OAI21_X1   g25123(.A1(new_n28241_), .A2(new_n28242_), .B(pi0243), .ZN(new_n28243_));
  NAND3_X1   g25124(.A1(new_n28239_), .A2(pi1156), .A3(new_n28243_), .ZN(new_n28244_));
  OAI22_X1   g25125(.A1(new_n28227_), .A2(new_n28222_), .B1(new_n28237_), .B2(new_n28244_), .ZN(new_n28245_));
  NOR2_X1    g25126(.A1(new_n28172_), .A2(new_n28147_), .ZN(new_n28246_));
  INV_X1     g25127(.I(new_n28246_), .ZN(new_n28247_));
  MUX2_X1    g25128(.I0(new_n28247_), .I1(new_n28127_), .S(pi0243), .Z(new_n28248_));
  INV_X1     g25129(.I(new_n28142_), .ZN(new_n28249_));
  NOR2_X1    g25130(.A1(new_n28134_), .A2(new_n28147_), .ZN(new_n28250_));
  INV_X1     g25131(.I(new_n28250_), .ZN(new_n28251_));
  NOR3_X1    g25132(.A1(new_n28251_), .A2(pi0243), .A3(new_n11912_), .ZN(new_n28252_));
  NOR4_X1    g25133(.A1(new_n28252_), .A2(new_n28249_), .A3(pi0243), .A4(pi1156), .ZN(new_n28253_));
  OAI21_X1   g25134(.A1(new_n28248_), .A2(pi1155), .B(new_n28253_), .ZN(new_n28254_));
  OAI22_X1   g25135(.A1(new_n28166_), .A2(new_n28164_), .B1(pi0243), .B2(new_n28173_), .ZN(new_n28255_));
  OAI21_X1   g25136(.A1(new_n28225_), .A2(new_n28255_), .B(new_n11912_), .ZN(new_n28256_));
  NAND4_X1   g25137(.A1(new_n28154_), .A2(new_n28163_), .A3(new_n28224_), .A4(new_n28250_), .ZN(new_n28257_));
  NOR2_X1    g25138(.A1(new_n26367_), .A2(pi1156), .ZN(new_n28258_));
  NAND4_X1   g25139(.A1(new_n28256_), .A2(new_n28254_), .A3(new_n28257_), .A4(new_n28258_), .ZN(new_n28259_));
  INV_X1     g25140(.I(pi0267), .ZN(new_n28260_));
  INV_X1     g25141(.I(pi0253), .ZN(new_n28261_));
  INV_X1     g25142(.I(pi0254), .ZN(new_n28262_));
  NOR2_X1    g25143(.A1(new_n28261_), .A2(new_n28262_), .ZN(new_n28263_));
  INV_X1     g25144(.I(new_n28263_), .ZN(new_n28264_));
  NOR2_X1    g25145(.A1(new_n28264_), .A2(new_n28260_), .ZN(new_n28265_));
  INV_X1     g25146(.I(new_n28265_), .ZN(new_n28266_));
  NOR2_X1    g25147(.A1(new_n28266_), .A2(pi0263), .ZN(new_n28267_));
  INV_X1     g25148(.I(new_n28267_), .ZN(new_n28268_));
  NOR2_X1    g25149(.A1(new_n26366_), .A2(new_n26910_), .ZN(new_n28269_));
  AOI21_X1   g25150(.A1(new_n28269_), .A2(pi1091), .B(pi0219), .ZN(new_n28270_));
  OAI21_X1   g25151(.A1(new_n28116_), .A2(pi0243), .B(new_n28270_), .ZN(new_n28271_));
  NAND2_X1   g25152(.A1(new_n28118_), .A2(new_n28164_), .ZN(new_n28272_));
  NAND2_X1   g25153(.A1(new_n28140_), .A2(pi0243), .ZN(new_n28273_));
  NAND2_X1   g25154(.A1(new_n28165_), .A2(new_n26367_), .ZN(new_n28274_));
  OAI21_X1   g25155(.A1(new_n28144_), .A2(new_n28274_), .B(pi0219), .ZN(new_n28275_));
  AOI21_X1   g25156(.A1(new_n28146_), .A2(pi0243), .B(new_n28275_), .ZN(new_n28276_));
  AOI22_X1   g25157(.A1(new_n28273_), .A2(new_n28276_), .B1(new_n28271_), .B2(new_n28272_), .ZN(new_n28277_));
  MUX2_X1    g25158(.I0(new_n28277_), .I1(new_n28164_), .S(new_n28268_), .Z(new_n28278_));
  NAND2_X1   g25159(.A1(new_n28267_), .A2(new_n6845_), .ZN(new_n28279_));
  INV_X1     g25160(.I(pi0268), .ZN(new_n28280_));
  INV_X1     g25161(.I(pi0272), .ZN(new_n28281_));
  INV_X1     g25162(.I(pi0275), .ZN(new_n28282_));
  INV_X1     g25163(.I(pi0283), .ZN(new_n28283_));
  NOR3_X1    g25164(.A1(new_n28281_), .A2(new_n28282_), .A3(new_n28283_), .ZN(new_n28284_));
  INV_X1     g25165(.I(new_n28284_), .ZN(new_n28285_));
  NOR2_X1    g25166(.A1(new_n28285_), .A2(new_n28280_), .ZN(new_n28286_));
  INV_X1     g25167(.I(new_n28286_), .ZN(new_n28287_));
  NAND4_X1   g25168(.A1(new_n28279_), .A2(new_n28268_), .A3(new_n8247_), .A4(new_n28287_), .ZN(new_n28288_));
  AOI21_X1   g25169(.A1(new_n28278_), .A2(po1038), .B(new_n28288_), .ZN(new_n28289_));
  NAND3_X1   g25170(.A1(new_n28245_), .A2(new_n28259_), .A3(new_n28289_), .ZN(new_n28290_));
  NOR2_X1    g25171(.A1(new_n6845_), .A2(new_n28165_), .ZN(new_n28291_));
  NAND2_X1   g25172(.A1(new_n28287_), .A2(new_n26307_), .ZN(new_n28292_));
  NOR3_X1    g25173(.A1(new_n28291_), .A2(new_n28292_), .A3(po1038), .ZN(new_n28293_));
  OAI21_X1   g25174(.A1(new_n28212_), .A2(new_n28290_), .B(new_n28293_), .ZN(po0400));
  NAND3_X1   g25175(.A1(new_n27510_), .A2(new_n8250_), .A3(new_n27503_), .ZN(new_n28295_));
  OAI21_X1   g25176(.A1(new_n27503_), .A2(new_n8248_), .B(new_n27509_), .ZN(new_n28296_));
  AOI21_X1   g25177(.A1(new_n28295_), .A2(new_n28296_), .B(new_n26375_), .ZN(new_n28297_));
  NOR4_X1    g25178(.A1(new_n27483_), .A2(new_n2587_), .A3(new_n27481_), .A4(new_n28297_), .ZN(new_n28298_));
  NAND2_X1   g25179(.A1(new_n26996_), .A2(new_n27533_), .ZN(new_n28299_));
  NOR2_X1    g25180(.A1(new_n28298_), .A2(new_n28299_), .ZN(new_n28300_));
  NOR2_X1    g25181(.A1(new_n27484_), .A2(new_n27485_), .ZN(new_n28301_));
  OAI22_X1   g25182(.A1(new_n28300_), .A2(po1038), .B1(new_n28301_), .B2(new_n27498_), .ZN(new_n28302_));
  OAI21_X1   g25183(.A1(new_n27001_), .A2(pi0213), .B(new_n26374_), .ZN(new_n28303_));
  AOI21_X1   g25184(.A1(new_n28302_), .A2(pi0213), .B(new_n28303_), .ZN(new_n28304_));
  NOR2_X1    g25185(.A1(new_n26315_), .A2(new_n8247_), .ZN(new_n28305_));
  AOI21_X1   g25186(.A1(new_n28305_), .A2(pi0299), .B(new_n27494_), .ZN(new_n28306_));
  INV_X1     g25187(.I(new_n27805_), .ZN(new_n28307_));
  MUX2_X1    g25188(.I0(new_n28307_), .I1(new_n26479_), .S(pi0211), .Z(new_n28308_));
  NAND2_X1   g25189(.A1(new_n27720_), .A2(new_n28308_), .ZN(new_n28309_));
  INV_X1     g25190(.I(new_n28309_), .ZN(new_n28310_));
  NAND2_X1   g25191(.A1(pi0212), .A2(pi0214), .ZN(new_n28311_));
  OAI21_X1   g25192(.A1(new_n28310_), .A2(new_n28311_), .B(new_n8247_), .ZN(new_n28312_));
  OAI21_X1   g25193(.A1(new_n27564_), .A2(new_n26313_), .B(pi0212), .ZN(new_n28313_));
  AOI21_X1   g25194(.A1(new_n28309_), .A2(new_n8078_), .B(new_n28313_), .ZN(new_n28314_));
  NAND3_X1   g25195(.A1(new_n28312_), .A2(new_n27720_), .A3(new_n28314_), .ZN(new_n28315_));
  AOI21_X1   g25196(.A1(new_n27724_), .A2(new_n28306_), .B(new_n28315_), .ZN(new_n28316_));
  AND2_X2    g25197(.A1(new_n28314_), .A2(new_n27733_), .Z(new_n28317_));
  NOR3_X1    g25198(.A1(new_n8077_), .A2(new_n2587_), .A3(new_n3548_), .ZN(new_n28318_));
  NAND2_X1   g25199(.A1(pi0212), .A2(pi0214), .ZN(new_n28319_));
  AOI21_X1   g25200(.A1(new_n28310_), .A2(new_n27733_), .B(new_n28319_), .ZN(new_n28320_));
  NOR2_X1    g25201(.A1(po1038), .A2(pi1147), .ZN(new_n28321_));
  INV_X1     g25202(.I(new_n28321_), .ZN(new_n28322_));
  NAND4_X1   g25203(.A1(new_n27799_), .A2(new_n27798_), .A3(new_n8247_), .A4(new_n28322_), .ZN(new_n28323_));
  NOR4_X1    g25204(.A1(new_n28317_), .A2(new_n28318_), .A3(new_n28320_), .A4(new_n28323_), .ZN(new_n28324_));
  NOR4_X1    g25205(.A1(new_n28316_), .A2(pi0213), .A3(new_n28324_), .A4(new_n26985_), .ZN(new_n28325_));
  OAI21_X1   g25206(.A1(new_n27812_), .A2(new_n24753_), .B(new_n28325_), .ZN(new_n28326_));
  AOI21_X1   g25207(.A1(new_n28326_), .A2(pi0209), .B(new_n28304_), .ZN(new_n28327_));
  MUX2_X1    g25208(.I0(new_n28327_), .I1(pi0244), .S(new_n26307_), .Z(po0401));
  NAND2_X1   g25209(.A1(new_n28072_), .A2(new_n2587_), .ZN(new_n28329_));
  NOR2_X1    g25210(.A1(new_n27508_), .A2(new_n8078_), .ZN(new_n28330_));
  NAND3_X1   g25211(.A1(new_n28329_), .A2(new_n8076_), .A3(new_n28330_), .ZN(new_n28331_));
  OAI21_X1   g25212(.A1(new_n28073_), .A2(pi0212), .B(new_n8247_), .ZN(new_n28332_));
  NAND3_X1   g25213(.A1(new_n28331_), .A2(new_n28075_), .A3(new_n28332_), .ZN(new_n28333_));
  NOR2_X1    g25214(.A1(new_n27621_), .A2(new_n3258_), .ZN(new_n28334_));
  NOR2_X1    g25215(.A1(new_n28334_), .A2(pi1147), .ZN(new_n28335_));
  INV_X1     g25216(.I(new_n28335_), .ZN(new_n28336_));
  INV_X1     g25217(.I(new_n28068_), .ZN(new_n28337_));
  NAND2_X1   g25218(.A1(new_n28337_), .A2(new_n26309_), .ZN(new_n28338_));
  AOI21_X1   g25219(.A1(new_n28338_), .A2(new_n28082_), .B(po1038), .ZN(new_n28339_));
  AND3_X2    g25220(.A1(new_n28333_), .A2(new_n28336_), .A3(new_n28339_), .Z(new_n28340_));
  INV_X1     g25221(.I(new_n27740_), .ZN(new_n28341_));
  NAND2_X1   g25222(.A1(new_n28334_), .A2(new_n27758_), .ZN(new_n28342_));
  INV_X1     g25223(.I(new_n28342_), .ZN(new_n28343_));
  AOI21_X1   g25224(.A1(pi1147), .A2(new_n28341_), .B(new_n28343_), .ZN(new_n28344_));
  NOR2_X1    g25225(.A1(new_n28070_), .A2(pi0299), .ZN(new_n28345_));
  INV_X1     g25226(.I(new_n28345_), .ZN(new_n28346_));
  NOR2_X1    g25227(.A1(new_n28346_), .A2(pi0211), .ZN(new_n28347_));
  NOR2_X1    g25228(.A1(new_n28337_), .A2(new_n8077_), .ZN(new_n28348_));
  NOR3_X1    g25229(.A1(new_n28074_), .A2(pi0214), .A3(new_n27246_), .ZN(new_n28349_));
  OAI21_X1   g25230(.A1(new_n28347_), .A2(new_n28348_), .B(pi0214), .ZN(new_n28350_));
  NOR2_X1    g25231(.A1(new_n28074_), .A2(new_n27246_), .ZN(new_n28351_));
  AOI21_X1   g25232(.A1(new_n8078_), .A2(new_n28351_), .B(new_n28350_), .ZN(new_n28352_));
  OAI21_X1   g25233(.A1(pi0212), .A2(new_n28075_), .B(new_n28351_), .ZN(new_n28353_));
  NAND3_X1   g25234(.A1(new_n28353_), .A2(pi0212), .A3(new_n8247_), .ZN(new_n28354_));
  NOR4_X1    g25235(.A1(new_n28352_), .A2(new_n28339_), .A3(new_n28349_), .A4(new_n28354_), .ZN(new_n28355_));
  OAI22_X1   g25236(.A1(new_n28340_), .A2(pi1148), .B1(new_n28344_), .B2(new_n28355_), .ZN(new_n28356_));
  AOI21_X1   g25237(.A1(new_n28346_), .A2(new_n8077_), .B(new_n28074_), .ZN(new_n28357_));
  NAND4_X1   g25238(.A1(new_n28329_), .A2(new_n8076_), .A3(pi0214), .A4(new_n27790_), .ZN(new_n28358_));
  INV_X1     g25239(.I(new_n28357_), .ZN(new_n28359_));
  NAND2_X1   g25240(.A1(new_n28359_), .A2(new_n28076_), .ZN(new_n28360_));
  NAND3_X1   g25241(.A1(new_n28336_), .A2(new_n27318_), .A3(new_n27597_), .ZN(new_n28361_));
  INV_X1     g25242(.I(new_n28361_), .ZN(new_n28362_));
  NOR3_X1    g25243(.A1(new_n28362_), .A2(pi0219), .A3(new_n28339_), .ZN(new_n28363_));
  NAND3_X1   g25244(.A1(new_n28358_), .A2(new_n28360_), .A3(new_n28363_), .ZN(new_n28364_));
  INV_X1     g25245(.I(new_n28350_), .ZN(new_n28365_));
  AOI21_X1   g25246(.A1(new_n28346_), .A2(new_n28076_), .B(pi0219), .ZN(new_n28366_));
  NAND2_X1   g25247(.A1(new_n28345_), .A2(new_n8078_), .ZN(new_n28367_));
  NAND4_X1   g25248(.A1(new_n28367_), .A2(pi0212), .A3(new_n27515_), .A4(new_n28342_), .ZN(new_n28368_));
  NOR4_X1    g25249(.A1(new_n28365_), .A2(new_n28366_), .A3(new_n28368_), .A4(new_n28339_), .ZN(new_n28369_));
  AOI21_X1   g25250(.A1(new_n28369_), .A2(new_n28364_), .B(new_n24753_), .ZN(new_n28370_));
  OAI21_X1   g25251(.A1(new_n28085_), .A2(pi0213), .B(new_n26374_), .ZN(new_n28371_));
  AOI21_X1   g25252(.A1(new_n28356_), .A2(new_n28370_), .B(new_n28371_), .ZN(new_n28372_));
  INV_X1     g25253(.I(new_n28344_), .ZN(new_n28373_));
  NOR3_X1    g25254(.A1(new_n8094_), .A2(pi0200), .A3(pi1146), .ZN(new_n28374_));
  NOR2_X1    g25255(.A1(new_n27709_), .A2(new_n28374_), .ZN(new_n28375_));
  INV_X1     g25256(.I(new_n28375_), .ZN(new_n28376_));
  NOR3_X1    g25257(.A1(new_n8094_), .A2(new_n3258_), .A3(pi0200), .ZN(new_n28377_));
  NOR2_X1    g25258(.A1(new_n8098_), .A2(pi0199), .ZN(new_n28378_));
  OAI21_X1   g25259(.A1(new_n28377_), .A2(new_n28378_), .B(new_n2587_), .ZN(new_n28379_));
  INV_X1     g25260(.I(new_n28379_), .ZN(new_n28380_));
  NOR3_X1    g25261(.A1(new_n28376_), .A2(new_n8087_), .A3(new_n8088_), .ZN(new_n28381_));
  NOR2_X1    g25262(.A1(new_n28376_), .A2(new_n8087_), .ZN(new_n28382_));
  NAND2_X1   g25263(.A1(new_n28382_), .A2(pi0208), .ZN(new_n28383_));
  INV_X1     g25264(.I(new_n28383_), .ZN(new_n28384_));
  NOR3_X1    g25265(.A1(new_n28384_), .A2(new_n26677_), .A3(new_n28379_), .ZN(new_n28385_));
  NOR2_X1    g25266(.A1(new_n28385_), .A2(new_n28381_), .ZN(new_n28386_));
  NOR2_X1    g25267(.A1(new_n28386_), .A2(pi0214), .ZN(new_n28387_));
  NOR2_X1    g25268(.A1(new_n28387_), .A2(pi0212), .ZN(new_n28388_));
  INV_X1     g25269(.I(new_n28388_), .ZN(new_n28389_));
  AOI21_X1   g25270(.A1(new_n28386_), .A2(new_n27528_), .B(new_n8078_), .ZN(new_n28390_));
  NOR4_X1    g25271(.A1(new_n28376_), .A2(new_n8087_), .A3(pi0208), .A4(new_n27507_), .ZN(new_n28391_));
  AOI21_X1   g25272(.A1(new_n28380_), .A2(pi0207), .B(new_n27506_), .ZN(new_n28392_));
  NOR3_X1    g25273(.A1(new_n28391_), .A2(pi0208), .A3(new_n28392_), .ZN(new_n28393_));
  INV_X1     g25274(.I(new_n28393_), .ZN(new_n28394_));
  NOR2_X1    g25275(.A1(new_n28394_), .A2(pi0299), .ZN(new_n28395_));
  NOR2_X1    g25276(.A1(new_n28395_), .A2(new_n8078_), .ZN(new_n28396_));
  NOR2_X1    g25277(.A1(new_n26493_), .A2(new_n28374_), .ZN(new_n28397_));
  NAND2_X1   g25278(.A1(new_n28397_), .A2(new_n26678_), .ZN(new_n28398_));
  XNOR2_X1   g25279(.A1(new_n28383_), .A2(new_n28398_), .ZN(new_n28399_));
  INV_X1     g25280(.I(new_n28399_), .ZN(new_n28400_));
  NOR2_X1    g25281(.A1(new_n28376_), .A2(new_n8088_), .ZN(new_n28401_));
  NAND2_X1   g25282(.A1(new_n28397_), .A2(new_n26549_), .ZN(new_n28402_));
  XOR2_X1    g25283(.A1(new_n28401_), .A2(new_n28402_), .Z(new_n28403_));
  AOI21_X1   g25284(.A1(new_n2587_), .A2(new_n28391_), .B(new_n28403_), .ZN(new_n28404_));
  INV_X1     g25285(.I(new_n28404_), .ZN(new_n28405_));
  NOR2_X1    g25286(.A1(new_n28405_), .A2(pi0299), .ZN(new_n28406_));
  INV_X1     g25287(.I(new_n28406_), .ZN(new_n28407_));
  AOI21_X1   g25288(.A1(new_n28407_), .A2(new_n8077_), .B(new_n28400_), .ZN(new_n28408_));
  INV_X1     g25289(.I(new_n28408_), .ZN(new_n28409_));
  AOI21_X1   g25290(.A1(new_n28409_), .A2(new_n28396_), .B(new_n8076_), .ZN(new_n28410_));
  INV_X1     g25291(.I(new_n28386_), .ZN(new_n28411_));
  OAI21_X1   g25292(.A1(new_n28411_), .A2(new_n27246_), .B(new_n8078_), .ZN(new_n28412_));
  AOI22_X1   g25293(.A1(new_n28410_), .A2(new_n28412_), .B1(new_n28389_), .B2(new_n28390_), .ZN(new_n28413_));
  OAI21_X1   g25294(.A1(new_n27181_), .A2(pi1146), .B(new_n27561_), .ZN(new_n28414_));
  AND3_X2    g25295(.A1(new_n28413_), .A2(new_n8247_), .A3(new_n28414_), .Z(new_n28415_));
  NOR2_X1    g25296(.A1(new_n28411_), .A2(new_n26719_), .ZN(new_n28416_));
  NAND2_X1   g25297(.A1(new_n28386_), .A2(pi0211), .ZN(new_n28417_));
  NAND3_X1   g25298(.A1(new_n28417_), .A2(new_n26342_), .A3(new_n28394_), .ZN(new_n28418_));
  AOI21_X1   g25299(.A1(new_n28418_), .A2(new_n28416_), .B(po1038), .ZN(new_n28419_));
  OAI21_X1   g25300(.A1(new_n28415_), .A2(new_n28419_), .B(new_n28373_), .ZN(new_n28420_));
  NOR2_X1    g25301(.A1(new_n26412_), .A2(new_n3258_), .ZN(new_n28421_));
  AOI22_X1   g25302(.A1(new_n28421_), .A2(pi0207), .B1(pi1146), .B2(new_n26640_), .ZN(new_n28422_));
  OR3_X2     g25303(.A1(new_n28422_), .A2(pi0208), .A3(new_n27507_), .Z(new_n28423_));
  NOR3_X1    g25304(.A1(new_n8089_), .A2(new_n28374_), .A3(new_n26390_), .ZN(new_n28424_));
  OAI21_X1   g25305(.A1(new_n28401_), .A2(pi0207), .B(new_n28424_), .ZN(new_n28425_));
  OAI21_X1   g25306(.A1(pi0208), .A2(new_n27506_), .B(new_n28422_), .ZN(new_n28426_));
  NAND3_X1   g25307(.A1(new_n28423_), .A2(new_n28425_), .A3(new_n28426_), .ZN(new_n28427_));
  MUX2_X1    g25308(.I0(new_n28427_), .I1(new_n27938_), .S(new_n2587_), .Z(new_n28428_));
  NAND2_X1   g25309(.A1(new_n28428_), .A2(new_n28422_), .ZN(new_n28429_));
  XOR2_X1    g25310(.A1(new_n26389_), .A2(pi0208), .Z(new_n28430_));
  NAND2_X1   g25311(.A1(new_n28430_), .A2(pi0207), .ZN(new_n28431_));
  NAND2_X1   g25312(.A1(new_n26389_), .A2(pi0208), .ZN(new_n28432_));
  XOR2_X1    g25313(.A1(new_n28431_), .A2(new_n28432_), .Z(new_n28433_));
  NAND2_X1   g25314(.A1(new_n28433_), .A2(new_n28421_), .ZN(new_n28434_));
  NOR2_X1    g25315(.A1(new_n28421_), .A2(pi0299), .ZN(new_n28437_));
  NOR2_X1    g25316(.A1(new_n28427_), .A2(new_n28437_), .ZN(new_n28438_));
  NOR2_X1    g25317(.A1(new_n6845_), .A2(pi0219), .ZN(new_n28441_));
  NAND2_X1   g25318(.A1(new_n28429_), .A2(new_n28441_), .ZN(new_n28442_));
  AOI21_X1   g25319(.A1(new_n28442_), .A2(new_n28335_), .B(pi1148), .ZN(new_n28443_));
  NAND2_X1   g25320(.A1(new_n28420_), .A2(new_n28443_), .ZN(new_n28444_));
  NOR2_X1    g25321(.A1(new_n28427_), .A2(pi0299), .ZN(new_n28445_));
  INV_X1     g25322(.I(new_n28445_), .ZN(new_n28446_));
  NOR2_X1    g25323(.A1(new_n28438_), .A2(pi0299), .ZN(new_n28447_));
  NOR3_X1    g25324(.A1(new_n28446_), .A2(new_n8077_), .A3(new_n28434_), .ZN(new_n28448_));
  INV_X1     g25325(.I(new_n28448_), .ZN(new_n28449_));
  NAND2_X1   g25326(.A1(new_n28449_), .A2(new_n8076_), .ZN(new_n28450_));
  NOR2_X1    g25327(.A1(new_n28445_), .A2(pi0214), .ZN(new_n28451_));
  AOI21_X1   g25328(.A1(new_n28450_), .A2(new_n28451_), .B(pi0219), .ZN(new_n28452_));
  OAI21_X1   g25329(.A1(new_n28449_), .A2(pi0214), .B(pi0212), .ZN(new_n28453_));
  NAND3_X1   g25330(.A1(new_n28453_), .A2(new_n28330_), .A3(new_n28446_), .ZN(new_n28454_));
  AOI21_X1   g25331(.A1(new_n28445_), .A2(new_n26319_), .B(new_n8247_), .ZN(new_n28455_));
  INV_X1     g25332(.I(new_n28427_), .ZN(new_n28456_));
  NAND2_X1   g25333(.A1(new_n28456_), .A2(new_n26309_), .ZN(new_n28457_));
  AOI21_X1   g25334(.A1(new_n28455_), .A2(new_n28457_), .B(po1038), .ZN(new_n28458_));
  OAI21_X1   g25335(.A1(new_n28454_), .A2(new_n28452_), .B(new_n28458_), .ZN(new_n28459_));
  NOR2_X1    g25336(.A1(new_n28400_), .A2(pi0214), .ZN(new_n28460_));
  INV_X1     g25337(.I(new_n28460_), .ZN(new_n28461_));
  NAND2_X1   g25338(.A1(new_n28461_), .A2(new_n8076_), .ZN(new_n28462_));
  NOR2_X1    g25339(.A1(new_n28462_), .A2(new_n28406_), .ZN(new_n28463_));
  NOR4_X1    g25340(.A1(new_n28405_), .A2(new_n2587_), .A3(pi1146), .A4(new_n26597_), .ZN(new_n28464_));
  NOR2_X1    g25341(.A1(new_n28405_), .A2(new_n27506_), .ZN(new_n28465_));
  NAND2_X1   g25342(.A1(new_n26309_), .A2(new_n8247_), .ZN(new_n28466_));
  NOR2_X1    g25343(.A1(new_n28343_), .A2(po1038), .ZN(new_n28467_));
  OAI21_X1   g25344(.A1(new_n28465_), .A2(new_n28466_), .B(new_n28467_), .ZN(new_n28468_));
  NOR4_X1    g25345(.A1(new_n28463_), .A2(pi0219), .A3(new_n28464_), .A4(new_n28468_), .ZN(new_n28469_));
  AOI21_X1   g25346(.A1(new_n28459_), .A2(new_n28362_), .B(new_n28469_), .ZN(new_n28470_));
  OAI21_X1   g25347(.A1(pi1148), .A2(new_n28470_), .B(new_n28444_), .ZN(new_n28471_));
  NOR2_X1    g25348(.A1(new_n28447_), .A2(new_n8078_), .ZN(new_n28472_));
  NAND2_X1   g25349(.A1(new_n28446_), .A2(new_n27504_), .ZN(new_n28473_));
  NOR2_X1    g25350(.A1(new_n28434_), .A2(pi0214), .ZN(new_n28474_));
  AOI21_X1   g25351(.A1(new_n28472_), .A2(new_n28473_), .B(new_n28474_), .ZN(new_n28475_));
  OAI21_X1   g25352(.A1(new_n28434_), .A2(new_n26342_), .B(pi0219), .ZN(new_n28476_));
  INV_X1     g25353(.I(new_n28447_), .ZN(new_n28477_));
  NAND2_X1   g25354(.A1(new_n28477_), .A2(new_n26479_), .ZN(new_n28478_));
  NOR2_X1    g25355(.A1(new_n26342_), .A2(pi0211), .ZN(new_n28479_));
  AOI21_X1   g25356(.A1(new_n28478_), .A2(new_n28479_), .B(new_n28476_), .ZN(new_n28480_));
  NOR2_X1    g25357(.A1(new_n28061_), .A2(new_n2587_), .ZN(new_n28481_));
  NOR2_X1    g25358(.A1(new_n28445_), .A2(new_n28481_), .ZN(new_n28482_));
  NAND3_X1   g25359(.A1(new_n28322_), .A2(new_n8076_), .A3(new_n8247_), .ZN(new_n28483_));
  OR3_X2     g25360(.A1(new_n28480_), .A2(new_n28475_), .A3(new_n28483_), .Z(new_n28484_));
  NOR2_X1    g25361(.A1(po1038), .A2(new_n27494_), .ZN(new_n28485_));
  NOR2_X1    g25362(.A1(new_n28405_), .A2(new_n26476_), .ZN(new_n28486_));
  NOR2_X1    g25363(.A1(new_n28486_), .A2(new_n28395_), .ZN(new_n28487_));
  NOR2_X1    g25364(.A1(new_n28487_), .A2(pi0211), .ZN(new_n28488_));
  NAND3_X1   g25365(.A1(new_n28416_), .A2(new_n26342_), .A3(new_n28417_), .ZN(new_n28489_));
  OAI21_X1   g25366(.A1(new_n28488_), .A2(new_n28489_), .B(new_n28485_), .ZN(new_n28490_));
  NOR2_X1    g25367(.A1(new_n28405_), .A2(new_n27503_), .ZN(new_n28491_));
  INV_X1     g25368(.I(new_n28491_), .ZN(new_n28492_));
  AOI21_X1   g25369(.A1(new_n28492_), .A2(new_n28396_), .B(new_n28387_), .ZN(new_n28493_));
  OAI21_X1   g25370(.A1(new_n28405_), .A2(new_n28481_), .B(pi0212), .ZN(new_n28494_));
  AOI21_X1   g25371(.A1(new_n28494_), .A2(new_n28395_), .B(pi0219), .ZN(new_n28495_));
  OAI21_X1   g25372(.A1(new_n28493_), .A2(pi0212), .B(new_n28495_), .ZN(new_n28496_));
  NAND2_X1   g25373(.A1(new_n28490_), .A2(new_n28496_), .ZN(new_n28497_));
  NAND3_X1   g25374(.A1(new_n28497_), .A2(new_n27515_), .A3(new_n28065_), .ZN(new_n28498_));
  NAND2_X1   g25375(.A1(new_n27503_), .A2(pi0214), .ZN(new_n28499_));
  AOI21_X1   g25376(.A1(new_n28446_), .A2(new_n28499_), .B(pi0212), .ZN(new_n28500_));
  OAI21_X1   g25377(.A1(new_n28482_), .A2(new_n8076_), .B(new_n8247_), .ZN(new_n28501_));
  NOR2_X1    g25378(.A1(new_n28501_), .A2(new_n28500_), .ZN(new_n28502_));
  INV_X1     g25379(.I(new_n28455_), .ZN(new_n28503_));
  NOR2_X1    g25380(.A1(new_n28456_), .A2(pi0299), .ZN(new_n28504_));
  NOR2_X1    g25381(.A1(new_n28504_), .A2(new_n26319_), .ZN(new_n28505_));
  NAND4_X1   g25382(.A1(new_n28503_), .A2(new_n28505_), .A3(new_n26479_), .A4(new_n28322_), .ZN(new_n28506_));
  NAND3_X1   g25383(.A1(new_n28462_), .A2(pi0214), .A3(new_n28491_), .ZN(new_n28507_));
  NAND3_X1   g25384(.A1(new_n28507_), .A2(new_n8247_), .A3(new_n28494_), .ZN(new_n28508_));
  AOI21_X1   g25385(.A1(new_n28400_), .A2(new_n26319_), .B(new_n8247_), .ZN(new_n28509_));
  NOR4_X1    g25386(.A1(new_n28486_), .A2(new_n28509_), .A3(new_n26319_), .A4(new_n28485_), .ZN(new_n28510_));
  NAND2_X1   g25387(.A1(new_n28065_), .A2(pi1148), .ZN(new_n28511_));
  AOI21_X1   g25388(.A1(new_n28508_), .A2(new_n28510_), .B(new_n28511_), .ZN(new_n28512_));
  OAI21_X1   g25389(.A1(new_n28502_), .A2(new_n28506_), .B(new_n28512_), .ZN(new_n28513_));
  NAND3_X1   g25390(.A1(new_n28513_), .A2(new_n26374_), .A3(new_n24753_), .ZN(new_n28514_));
  AOI21_X1   g25391(.A1(new_n28484_), .A2(new_n28498_), .B(new_n28514_), .ZN(new_n28515_));
  AOI21_X1   g25392(.A1(new_n28471_), .A2(new_n28515_), .B(new_n28372_), .ZN(new_n28516_));
  MUX2_X1    g25393(.I0(new_n28516_), .I1(pi0245), .S(new_n26307_), .Z(po0402));
  NOR2_X1    g25394(.A1(new_n27272_), .A2(pi0212), .ZN(new_n28518_));
  OAI21_X1   g25395(.A1(new_n27849_), .A2(pi0219), .B(new_n28518_), .ZN(new_n28519_));
  INV_X1     g25396(.I(new_n28519_), .ZN(new_n28520_));
  OAI21_X1   g25397(.A1(new_n27581_), .A2(new_n8078_), .B(new_n27832_), .ZN(new_n28521_));
  AOI21_X1   g25398(.A1(pi0219), .A2(new_n27507_), .B(new_n27630_), .ZN(new_n28522_));
  OAI21_X1   g25399(.A1(new_n27589_), .A2(new_n28522_), .B(new_n28342_), .ZN(new_n28523_));
  AOI21_X1   g25400(.A1(new_n28521_), .A2(new_n28520_), .B(new_n28523_), .ZN(new_n28524_));
  NOR2_X1    g25401(.A1(new_n28522_), .A2(new_n27589_), .ZN(new_n28525_));
  INV_X1     g25402(.I(new_n28525_), .ZN(new_n28526_));
  NOR3_X1    g25403(.A1(new_n27271_), .A2(pi0212), .A3(pi0214), .ZN(new_n28528_));
  NOR4_X1    g25404(.A1(new_n27603_), .A2(pi0219), .A3(new_n28526_), .A4(new_n28528_), .ZN(new_n28529_));
  NOR4_X1    g25405(.A1(new_n28524_), .A2(pi1150), .A3(new_n28361_), .A4(new_n28529_), .ZN(new_n28530_));
  INV_X1     g25406(.I(new_n28522_), .ZN(new_n28531_));
  NOR2_X1    g25407(.A1(new_n27526_), .A2(new_n27529_), .ZN(new_n28532_));
  OAI22_X1   g25408(.A1(new_n28532_), .A2(new_n26314_), .B1(new_n27525_), .B2(new_n27657_), .ZN(new_n28533_));
  INV_X1     g25409(.I(new_n27524_), .ZN(new_n28534_));
  NAND2_X1   g25410(.A1(new_n27512_), .A2(new_n28534_), .ZN(new_n28535_));
  AOI22_X1   g25411(.A1(new_n28533_), .A2(new_n8247_), .B1(new_n28531_), .B2(new_n28535_), .ZN(new_n28536_));
  AOI21_X1   g25412(.A1(new_n8247_), .A2(new_n27526_), .B(new_n27629_), .ZN(new_n28537_));
  AOI21_X1   g25413(.A1(new_n28361_), .A2(new_n28342_), .B(pi1150), .ZN(new_n28538_));
  OAI21_X1   g25414(.A1(new_n28361_), .A2(new_n28537_), .B(new_n28538_), .ZN(new_n28539_));
  OAI21_X1   g25415(.A1(new_n28539_), .A2(new_n28536_), .B(pi1148), .ZN(new_n28540_));
  NOR4_X1    g25416(.A1(new_n28531_), .A2(pi0219), .A3(new_n27473_), .A4(new_n27939_), .ZN(new_n28541_));
  OAI22_X1   g25417(.A1(new_n28344_), .A2(new_n28522_), .B1(new_n28336_), .B2(new_n28541_), .ZN(new_n28542_));
  NAND2_X1   g25418(.A1(new_n27613_), .A2(pi1150), .ZN(new_n28543_));
  OAI21_X1   g25419(.A1(new_n27528_), .A2(new_n26362_), .B(new_n8247_), .ZN(new_n28544_));
  AND2_X2    g25420(.A1(new_n28414_), .A2(new_n28544_), .Z(new_n28545_));
  NOR3_X1    g25421(.A1(new_n28545_), .A2(new_n27817_), .A3(new_n27197_), .ZN(new_n28546_));
  AOI22_X1   g25422(.A1(new_n28542_), .A2(new_n28543_), .B1(new_n28373_), .B2(new_n28546_), .ZN(new_n28547_));
  OAI22_X1   g25423(.A1(new_n28540_), .A2(new_n28530_), .B1(pi1148), .B2(new_n28547_), .ZN(new_n28548_));
  NAND2_X1   g25424(.A1(new_n8088_), .A2(pi0299), .ZN(new_n28549_));
  NAND3_X1   g25425(.A1(new_n27507_), .A2(new_n27539_), .A3(new_n28549_), .ZN(new_n28550_));
  INV_X1     g25426(.I(new_n27651_), .ZN(new_n28551_));
  NOR3_X1    g25427(.A1(new_n27990_), .A2(pi0214), .A3(new_n27232_), .ZN(new_n28552_));
  AOI21_X1   g25428(.A1(new_n28551_), .A2(new_n28552_), .B(pi0219), .ZN(new_n28553_));
  NOR2_X1    g25429(.A1(new_n27990_), .A2(new_n27232_), .ZN(new_n28554_));
  NOR2_X1    g25430(.A1(new_n28554_), .A2(new_n27549_), .ZN(new_n28555_));
  AOI21_X1   g25431(.A1(new_n8076_), .A2(new_n28555_), .B(new_n28553_), .ZN(new_n28556_));
  OAI22_X1   g25432(.A1(new_n28553_), .A2(new_n28555_), .B1(new_n27547_), .B2(new_n28522_), .ZN(new_n28557_));
  AOI21_X1   g25433(.A1(new_n28550_), .A2(new_n28556_), .B(new_n28557_), .ZN(new_n28558_));
  AOI21_X1   g25434(.A1(new_n28558_), .A2(new_n28373_), .B(new_n27817_), .ZN(new_n28559_));
  OAI21_X1   g25435(.A1(po1038), .A2(new_n27233_), .B(new_n28558_), .ZN(new_n28560_));
  NOR2_X1    g25436(.A1(new_n28007_), .A2(pi0219), .ZN(new_n28561_));
  OAI21_X1   g25437(.A1(new_n27551_), .A2(new_n27650_), .B(new_n28561_), .ZN(new_n28562_));
  INV_X1     g25438(.I(new_n28562_), .ZN(new_n28563_));
  NAND4_X1   g25439(.A1(new_n28560_), .A2(new_n27545_), .A3(new_n28336_), .A4(new_n28563_), .ZN(new_n28564_));
  AOI21_X1   g25440(.A1(new_n27487_), .A2(new_n27674_), .B(new_n27689_), .ZN(new_n28565_));
  NOR2_X1    g25441(.A1(new_n27669_), .A2(pi1146), .ZN(new_n28566_));
  NOR2_X1    g25442(.A1(new_n28566_), .A2(pi0219), .ZN(new_n28567_));
  AOI21_X1   g25443(.A1(new_n27472_), .A2(new_n27563_), .B(new_n27669_), .ZN(new_n28568_));
  OR4_X2     g25444(.A1(new_n27688_), .A2(new_n28565_), .A3(new_n28567_), .A4(new_n28568_), .Z(new_n28569_));
  NAND2_X1   g25445(.A1(new_n27671_), .A2(new_n27848_), .ZN(new_n28570_));
  AOI21_X1   g25446(.A1(new_n28570_), .A2(new_n8247_), .B(new_n28565_), .ZN(new_n28571_));
  OR3_X2     g25447(.A1(new_n28571_), .A2(new_n28335_), .A3(new_n28566_), .Z(new_n28572_));
  AOI21_X1   g25448(.A1(new_n28572_), .A2(new_n27817_), .B(new_n28344_), .ZN(new_n28573_));
  OAI21_X1   g25449(.A1(new_n27194_), .A2(new_n27390_), .B(new_n27624_), .ZN(new_n28575_));
  INV_X1     g25450(.I(new_n27560_), .ZN(new_n28583_));
  AOI21_X1   g25451(.A1(pi0214), .A2(new_n27566_), .B(new_n27562_), .ZN(new_n28584_));
  NOR4_X1    g25452(.A1(new_n28583_), .A2(pi0219), .A3(new_n27565_), .A4(new_n28584_), .ZN(new_n28585_));
  AOI21_X1   g25453(.A1(new_n28569_), .A2(new_n28573_), .B(pi1148), .ZN(new_n28589_));
  OAI21_X1   g25454(.A1(new_n28564_), .A2(new_n28559_), .B(new_n28589_), .ZN(new_n28590_));
  MUX2_X1    g25455(.I0(new_n28590_), .I1(new_n28548_), .S(new_n27470_), .Z(new_n28591_));
  NAND4_X1   g25456(.A1(new_n27693_), .A2(new_n27470_), .A3(pi1150), .A4(new_n27656_), .ZN(new_n28592_));
  NAND2_X1   g25457(.A1(new_n27618_), .A2(new_n27470_), .ZN(new_n28593_));
  AOI21_X1   g25458(.A1(new_n28593_), .A2(new_n27817_), .B(pi1148), .ZN(new_n28594_));
  NAND2_X1   g25459(.A1(new_n28592_), .A2(new_n28594_), .ZN(new_n28595_));
  INV_X1     g25460(.I(new_n27612_), .ZN(new_n28596_));
  AOI21_X1   g25461(.A1(new_n27644_), .A2(new_n27817_), .B(new_n28596_), .ZN(new_n28597_));
  NOR3_X1    g25462(.A1(new_n27644_), .A2(new_n27612_), .A3(pi1150), .ZN(new_n28598_));
  NOR2_X1    g25463(.A1(new_n27700_), .A2(pi1150), .ZN(new_n28599_));
  NOR4_X1    g25464(.A1(new_n27659_), .A2(new_n27817_), .A3(new_n27662_), .A4(new_n27663_), .ZN(new_n28600_));
  OAI21_X1   g25465(.A1(new_n28599_), .A2(new_n28600_), .B(new_n27470_), .ZN(new_n28601_));
  NOR3_X1    g25466(.A1(new_n28597_), .A2(new_n28598_), .A3(new_n28601_), .ZN(new_n28602_));
  NOR2_X1    g25467(.A1(new_n28602_), .A2(new_n27515_), .ZN(new_n28603_));
  XOR2_X1    g25468(.A1(new_n28603_), .A2(new_n28595_), .Z(new_n28604_));
  MUX2_X1    g25469(.I0(new_n28604_), .I1(new_n28591_), .S(new_n24753_), .Z(new_n28605_));
  NOR3_X1    g25470(.A1(new_n28471_), .A2(new_n26374_), .A3(pi0213), .ZN(new_n28677_));
  AOI21_X1   g25471(.A1(new_n28605_), .A2(pi0209), .B(new_n28677_), .ZN(new_n28678_));
  MUX2_X1    g25472(.I0(new_n28678_), .I1(pi0246), .S(new_n26307_), .Z(po0403));
  INV_X1     g25473(.I(new_n27950_), .ZN(new_n28680_));
  AOI21_X1   g25474(.A1(new_n27627_), .A2(new_n28575_), .B(new_n28680_), .ZN(new_n28681_));
  AOI21_X1   g25475(.A1(new_n27639_), .A2(new_n8247_), .B(new_n28680_), .ZN(new_n28682_));
  NOR2_X1    g25476(.A1(new_n28681_), .A2(new_n28682_), .ZN(new_n28683_));
  NAND2_X1   g25477(.A1(new_n28683_), .A2(new_n27841_), .ZN(new_n28684_));
  INV_X1     g25478(.I(new_n28682_), .ZN(new_n28685_));
  AOI21_X1   g25479(.A1(new_n28685_), .A2(new_n27862_), .B(new_n27494_), .ZN(new_n28686_));
  AOI21_X1   g25480(.A1(new_n28684_), .A2(new_n28686_), .B(new_n27817_), .ZN(new_n28687_));
  AOI21_X1   g25481(.A1(new_n27687_), .A2(new_n27689_), .B(new_n27842_), .ZN(new_n28688_));
  NOR4_X1    g25482(.A1(new_n28016_), .A2(pi1147), .A3(new_n28687_), .A4(new_n28688_), .ZN(new_n28689_));
  NAND2_X1   g25483(.A1(new_n27520_), .A2(new_n27251_), .ZN(new_n28690_));
  NAND2_X1   g25484(.A1(new_n28690_), .A2(new_n27494_), .ZN(new_n28691_));
  INV_X1     g25485(.I(new_n27497_), .ZN(new_n28692_));
  NOR2_X1    g25486(.A1(new_n28003_), .A2(new_n27999_), .ZN(new_n28693_));
  OAI21_X1   g25487(.A1(new_n28693_), .A2(po1038), .B(new_n28692_), .ZN(new_n28694_));
  INV_X1     g25488(.I(new_n28694_), .ZN(new_n28695_));
  NOR2_X1    g25489(.A1(new_n28695_), .A2(new_n28691_), .ZN(new_n28696_));
  NOR3_X1    g25490(.A1(new_n28681_), .A2(new_n27251_), .A3(new_n27497_), .ZN(new_n28697_));
  NOR3_X1    g25491(.A1(new_n28697_), .A2(new_n27494_), .A3(new_n27958_), .ZN(new_n28698_));
  NAND2_X1   g25492(.A1(new_n27817_), .A2(pi1149), .ZN(new_n28699_));
  OR3_X2     g25493(.A1(new_n28698_), .A2(new_n28696_), .A3(new_n28699_), .Z(new_n28700_));
  NOR2_X1    g25494(.A1(new_n28553_), .A2(new_n28555_), .ZN(new_n28701_));
  NOR2_X1    g25495(.A1(new_n28701_), .A2(new_n27546_), .ZN(new_n28702_));
  NOR2_X1    g25496(.A1(new_n28702_), .A2(new_n27740_), .ZN(new_n28703_));
  NAND2_X1   g25497(.A1(new_n28703_), .A2(new_n27251_), .ZN(new_n28704_));
  NOR4_X1    g25498(.A1(new_n27545_), .A2(new_n27653_), .A3(new_n27552_), .A4(new_n27879_), .ZN(new_n28705_));
  NOR2_X1    g25499(.A1(new_n28705_), .A2(pi1147), .ZN(new_n28706_));
  NAND2_X1   g25500(.A1(new_n27937_), .A2(new_n28341_), .ZN(new_n28707_));
  INV_X1     g25501(.I(new_n28707_), .ZN(new_n28708_));
  NAND4_X1   g25502(.A1(new_n28708_), .A2(new_n27494_), .A3(new_n27251_), .A4(new_n28025_), .ZN(new_n28709_));
  NAND2_X1   g25503(.A1(new_n28709_), .A2(pi1150), .ZN(new_n28710_));
  AOI21_X1   g25504(.A1(new_n28704_), .A2(new_n28706_), .B(new_n28710_), .ZN(new_n28711_));
  NOR3_X1    g25505(.A1(new_n28701_), .A2(new_n27546_), .A3(new_n28562_), .ZN(new_n28712_));
  NOR2_X1    g25506(.A1(new_n28712_), .A2(new_n27323_), .ZN(new_n28713_));
  INV_X1     g25507(.I(new_n27598_), .ZN(new_n28714_));
  OAI21_X1   g25508(.A1(new_n28562_), .A2(new_n27546_), .B(new_n28714_), .ZN(new_n28715_));
  NOR2_X1    g25509(.A1(new_n27942_), .A2(new_n27323_), .ZN(new_n28716_));
  INV_X1     g25510(.I(new_n27943_), .ZN(new_n28717_));
  NOR2_X1    g25511(.A1(new_n28717_), .A2(new_n27895_), .ZN(new_n28718_));
  NOR2_X1    g25512(.A1(pi1147), .A2(pi1150), .ZN(new_n28719_));
  OAI21_X1   g25513(.A1(new_n28715_), .A2(new_n27251_), .B(new_n28719_), .ZN(new_n28720_));
  NOR2_X1    g25514(.A1(new_n28713_), .A2(new_n28720_), .ZN(new_n28721_));
  NOR2_X1    g25515(.A1(new_n28711_), .A2(new_n28721_), .ZN(new_n28722_));
  OAI22_X1   g25516(.A1(new_n28689_), .A2(new_n28700_), .B1(new_n27470_), .B2(new_n28722_), .ZN(new_n28723_));
  NAND4_X1   g25517(.A1(new_n27610_), .A2(pi0212), .A3(new_n27575_), .A4(new_n28519_), .ZN(new_n28724_));
  NAND2_X1   g25518(.A1(new_n28724_), .A2(new_n27879_), .ZN(new_n28725_));
  NAND2_X1   g25519(.A1(new_n27970_), .A2(new_n8247_), .ZN(new_n28726_));
  OAI21_X1   g25520(.A1(new_n27915_), .A2(new_n28726_), .B(new_n27609_), .ZN(new_n28727_));
  AND2_X2    g25521(.A1(new_n28727_), .A2(new_n28341_), .Z(new_n28728_));
  NAND2_X1   g25522(.A1(new_n28728_), .A2(new_n27251_), .ZN(new_n28729_));
  NAND3_X1   g25523(.A1(new_n28729_), .A2(pi1147), .A3(new_n28725_), .ZN(new_n28730_));
  NOR2_X1    g25524(.A1(new_n27972_), .A2(new_n27740_), .ZN(new_n28731_));
  NAND2_X1   g25525(.A1(new_n28731_), .A2(new_n27251_), .ZN(new_n28732_));
  INV_X1     g25526(.I(new_n27401_), .ZN(new_n28733_));
  NOR4_X1    g25527(.A1(new_n27972_), .A2(new_n27249_), .A3(new_n28733_), .A4(new_n27879_), .ZN(new_n28734_));
  NOR2_X1    g25528(.A1(new_n28734_), .A2(pi1147), .ZN(new_n28735_));
  NAND2_X1   g25529(.A1(new_n28735_), .A2(new_n28732_), .ZN(new_n28736_));
  AOI21_X1   g25530(.A1(new_n28730_), .A2(new_n28736_), .B(pi1150), .ZN(new_n28737_));
  INV_X1     g25531(.I(new_n28021_), .ZN(new_n28738_));
  OAI21_X1   g25532(.A1(new_n28727_), .A2(new_n27606_), .B(new_n27322_), .ZN(new_n28739_));
  NAND3_X1   g25533(.A1(new_n28738_), .A2(pi1147), .A3(new_n28739_), .ZN(new_n28740_));
  NOR2_X1    g25534(.A1(new_n27926_), .A2(new_n27497_), .ZN(new_n28741_));
  INV_X1     g25535(.I(new_n28741_), .ZN(new_n28742_));
  INV_X1     g25536(.I(new_n27616_), .ZN(new_n28743_));
  NAND2_X1   g25537(.A1(new_n27494_), .A2(pi1151), .ZN(new_n28744_));
  OAI21_X1   g25538(.A1(new_n28743_), .A2(new_n28744_), .B(new_n27817_), .ZN(new_n28745_));
  NAND2_X1   g25539(.A1(new_n28535_), .A2(new_n27251_), .ZN(new_n28746_));
  NAND4_X1   g25540(.A1(new_n28745_), .A2(pi1147), .A3(new_n28742_), .A4(new_n28746_), .ZN(new_n28747_));
  INV_X1     g25541(.I(new_n27668_), .ZN(new_n28748_));
  INV_X1     g25542(.I(new_n27919_), .ZN(new_n28749_));
  OAI21_X1   g25543(.A1(new_n27641_), .A2(new_n28749_), .B(new_n28748_), .ZN(new_n28750_));
  NOR4_X1    g25544(.A1(new_n27919_), .A2(new_n27526_), .A3(new_n26650_), .A4(new_n27625_), .ZN(new_n28751_));
  NOR2_X1    g25545(.A1(new_n28751_), .A2(new_n27842_), .ZN(new_n28752_));
  NOR4_X1    g25546(.A1(new_n28750_), .A2(pi1147), .A3(pi1151), .A4(new_n28752_), .ZN(new_n28753_));
  AOI21_X1   g25547(.A1(new_n27614_), .A2(new_n26558_), .B(new_n27667_), .ZN(new_n28754_));
  NOR2_X1    g25548(.A1(new_n28754_), .A2(pi1151), .ZN(new_n28755_));
  NOR2_X1    g25549(.A1(new_n28755_), .A2(pi1147), .ZN(new_n28756_));
  OAI21_X1   g25550(.A1(new_n11749_), .A2(new_n27316_), .B(pi1151), .ZN(new_n28757_));
  NAND3_X1   g25551(.A1(new_n28756_), .A2(new_n27817_), .A3(new_n28757_), .ZN(new_n28758_));
  OAI21_X1   g25552(.A1(new_n28753_), .A2(new_n28758_), .B(new_n28747_), .ZN(new_n28759_));
  AOI21_X1   g25553(.A1(new_n27197_), .A2(new_n27941_), .B(new_n27971_), .ZN(new_n28760_));
  NOR3_X1    g25554(.A1(new_n27249_), .A2(new_n28733_), .A3(new_n8248_), .ZN(new_n28761_));
  NOR2_X1    g25555(.A1(new_n28760_), .A2(new_n28761_), .ZN(new_n28762_));
  NAND2_X1   g25556(.A1(new_n27494_), .A2(new_n27817_), .ZN(new_n28763_));
  NOR2_X1    g25557(.A1(new_n28760_), .A2(new_n27323_), .ZN(new_n28764_));
  NOR4_X1    g25558(.A1(new_n28764_), .A2(pi1148), .A3(new_n27470_), .A4(new_n28763_), .ZN(new_n28765_));
  OAI21_X1   g25559(.A1(new_n27895_), .A2(new_n28762_), .B(new_n28765_), .ZN(new_n28766_));
  AOI21_X1   g25560(.A1(new_n27470_), .A2(new_n28759_), .B(new_n28766_), .ZN(new_n28767_));
  NAND2_X1   g25561(.A1(new_n28740_), .A2(new_n28767_), .ZN(new_n28768_));
  OAI21_X1   g25562(.A1(new_n28737_), .A2(new_n28768_), .B(pi0213), .ZN(new_n28769_));
  AOI21_X1   g25563(.A1(new_n28723_), .A2(pi1148), .B(new_n28769_), .ZN(new_n28770_));
  OAI21_X1   g25564(.A1(new_n27704_), .A2(pi0213), .B(new_n26374_), .ZN(new_n28771_));
  NOR2_X1    g25565(.A1(new_n28771_), .A2(new_n28770_), .ZN(new_n28772_));
  NAND2_X1   g25566(.A1(new_n28703_), .A2(pi1151), .ZN(new_n28773_));
  AOI21_X1   g25567(.A1(new_n27672_), .A2(new_n27678_), .B(new_n28565_), .ZN(new_n28774_));
  NOR2_X1    g25568(.A1(new_n28774_), .A2(new_n27740_), .ZN(new_n28775_));
  NAND4_X1   g25569(.A1(new_n28773_), .A2(new_n27494_), .A3(new_n27251_), .A4(new_n28775_), .ZN(new_n28776_));
  NOR2_X1    g25570(.A1(new_n28016_), .A2(pi1147), .ZN(new_n28777_));
  NOR2_X1    g25571(.A1(new_n27401_), .A2(new_n27648_), .ZN(new_n28778_));
  NOR2_X1    g25572(.A1(new_n27668_), .A2(new_n27251_), .ZN(new_n28779_));
  OAI21_X1   g25573(.A1(new_n28556_), .A2(new_n28778_), .B(new_n28779_), .ZN(new_n28780_));
  NAND2_X1   g25574(.A1(new_n28777_), .A2(new_n28780_), .ZN(new_n28781_));
  NOR2_X1    g25575(.A1(new_n27317_), .A2(pi1151), .ZN(new_n28782_));
  INV_X1     g25576(.I(new_n28025_), .ZN(new_n28783_));
  NOR2_X1    g25577(.A1(new_n27662_), .A2(pi1151), .ZN(new_n28784_));
  INV_X1     g25578(.I(new_n28784_), .ZN(new_n28785_));
  NOR4_X1    g25579(.A1(new_n28783_), .A2(new_n27512_), .A3(new_n27659_), .A4(new_n28785_), .ZN(new_n28786_));
  NOR2_X1    g25580(.A1(new_n28585_), .A2(new_n27842_), .ZN(new_n28787_));
  INV_X1     g25581(.I(new_n28787_), .ZN(new_n28788_));
  NAND4_X1   g25582(.A1(new_n28786_), .A2(new_n28788_), .A3(new_n27817_), .A4(new_n27762_), .ZN(new_n28789_));
  AOI21_X1   g25583(.A1(new_n28683_), .A2(new_n28782_), .B(new_n28789_), .ZN(new_n28790_));
  NAND3_X1   g25584(.A1(new_n28781_), .A2(new_n28776_), .A3(new_n28790_), .ZN(new_n28791_));
  NAND3_X1   g25585(.A1(new_n28520_), .A2(new_n27590_), .A3(new_n27833_), .ZN(new_n28792_));
  NAND2_X1   g25586(.A1(new_n28792_), .A2(new_n27318_), .ZN(new_n28793_));
  NAND2_X1   g25587(.A1(new_n28793_), .A2(pi1151), .ZN(new_n28794_));
  NOR3_X1    g25588(.A1(new_n27635_), .A2(new_n28751_), .A3(new_n28785_), .ZN(new_n28795_));
  NOR3_X1    g25589(.A1(new_n28751_), .A2(pi1151), .A3(new_n27317_), .ZN(new_n28796_));
  INV_X1     g25590(.I(new_n28796_), .ZN(new_n28797_));
  AND3_X2    g25591(.A1(new_n28795_), .A2(new_n27762_), .A3(new_n28797_), .Z(new_n28798_));
  NAND4_X1   g25592(.A1(new_n28798_), .A2(pi1147), .A3(new_n28725_), .A4(new_n28794_), .ZN(new_n28799_));
  OAI21_X1   g25593(.A1(new_n27698_), .A2(pi1151), .B(new_n27494_), .ZN(new_n28800_));
  INV_X1     g25594(.I(new_n28779_), .ZN(new_n28801_));
  NOR2_X1    g25595(.A1(new_n27855_), .A2(new_n28733_), .ZN(new_n28802_));
  NOR4_X1    g25596(.A1(new_n28802_), .A2(pi1149), .A3(new_n28756_), .A4(new_n28801_), .ZN(new_n28803_));
  AOI21_X1   g25597(.A1(new_n28803_), .A2(new_n28800_), .B(pi1150), .ZN(new_n28804_));
  AOI21_X1   g25598(.A1(new_n28799_), .A2(new_n28804_), .B(new_n27515_), .ZN(new_n28805_));
  NAND2_X1   g25599(.A1(new_n28805_), .A2(new_n28791_), .ZN(new_n28806_));
  NOR2_X1    g25600(.A1(new_n27598_), .A2(pi1151), .ZN(new_n28807_));
  INV_X1     g25601(.I(new_n28807_), .ZN(new_n28808_));
  NOR2_X1    g25602(.A1(new_n27635_), .A2(new_n28808_), .ZN(new_n28809_));
  OR3_X2     g25603(.A1(new_n28021_), .A2(new_n28809_), .A3(new_n27494_), .Z(new_n28810_));
  AOI21_X1   g25604(.A1(new_n27605_), .A2(new_n27589_), .B(new_n27497_), .ZN(new_n28811_));
  INV_X1     g25605(.I(new_n28811_), .ZN(new_n28812_));
  NOR2_X1    g25606(.A1(new_n28812_), .A2(new_n27251_), .ZN(new_n28813_));
  OR3_X2     g25607(.A1(new_n28681_), .A2(pi1151), .A3(new_n27497_), .Z(new_n28814_));
  NOR2_X1    g25608(.A1(new_n27497_), .A2(new_n27251_), .ZN(new_n28815_));
  AOI21_X1   g25609(.A1(new_n27570_), .A2(new_n28815_), .B(pi1147), .ZN(new_n28816_));
  AOI21_X1   g25610(.A1(new_n28814_), .A2(new_n28816_), .B(new_n27817_), .ZN(new_n28817_));
  NAND4_X1   g25611(.A1(new_n27634_), .A2(new_n27494_), .A3(new_n27251_), .A4(new_n28714_), .ZN(new_n28818_));
  NOR2_X1    g25612(.A1(new_n28818_), .A2(new_n28817_), .ZN(new_n28819_));
  NOR2_X1    g25613(.A1(new_n28742_), .A2(pi1151), .ZN(new_n28820_));
  NOR4_X1    g25614(.A1(new_n28819_), .A2(new_n28763_), .A3(new_n28813_), .A4(new_n28820_), .ZN(new_n28821_));
  AOI21_X1   g25615(.A1(new_n28810_), .A2(new_n28821_), .B(new_n27470_), .ZN(new_n28822_));
  NAND2_X1   g25616(.A1(new_n27621_), .A2(pi1151), .ZN(new_n28823_));
  NOR2_X1    g25617(.A1(new_n28760_), .A2(new_n28823_), .ZN(new_n28824_));
  NAND3_X1   g25618(.A1(new_n27613_), .A2(new_n27494_), .A3(pi1151), .ZN(new_n28825_));
  AOI21_X1   g25619(.A1(new_n28825_), .A2(new_n27817_), .B(pi1147), .ZN(new_n28826_));
  OAI21_X1   g25620(.A1(new_n28824_), .A2(new_n28716_), .B(new_n28826_), .ZN(new_n28827_));
  NAND4_X1   g25621(.A1(new_n28571_), .A2(new_n27494_), .A3(new_n27251_), .A4(new_n27621_), .ZN(new_n28828_));
  NOR2_X1    g25622(.A1(new_n27648_), .A2(new_n27251_), .ZN(new_n28829_));
  NAND4_X1   g25623(.A1(new_n28828_), .A2(new_n27817_), .A3(new_n28691_), .A4(new_n28829_), .ZN(new_n28830_));
  AOI21_X1   g25624(.A1(new_n28827_), .A2(new_n28830_), .B(pi1149), .ZN(new_n28831_));
  OAI21_X1   g25625(.A1(new_n28822_), .A2(new_n28831_), .B(new_n27515_), .ZN(new_n28832_));
  NAND2_X1   g25626(.A1(new_n28806_), .A2(new_n28832_), .ZN(new_n28833_));
  MUX2_X1    g25627(.I0(new_n28833_), .I1(new_n28030_), .S(pi0213), .Z(new_n28834_));
  AOI21_X1   g25628(.A1(pi0209), .A2(new_n28834_), .B(new_n28772_), .ZN(new_n28835_));
  MUX2_X1    g25629(.I0(new_n28835_), .I1(pi0247), .S(new_n26307_), .Z(po0404));
  NAND2_X1   g25630(.A1(new_n27251_), .A2(new_n26604_), .ZN(new_n28837_));
  NOR3_X1    g25631(.A1(new_n28715_), .A2(new_n28705_), .A3(new_n28837_), .ZN(new_n28838_));
  NOR2_X1    g25632(.A1(new_n28713_), .A2(pi1152), .ZN(new_n28839_));
  AOI21_X1   g25633(.A1(new_n28839_), .A2(new_n28773_), .B(new_n28838_), .ZN(new_n28840_));
  NOR2_X1    g25634(.A1(new_n27691_), .A2(new_n28801_), .ZN(new_n28841_));
  NOR2_X1    g25635(.A1(new_n28841_), .A2(pi1152), .ZN(new_n28842_));
  NOR2_X1    g25636(.A1(new_n28694_), .A2(pi1151), .ZN(new_n28843_));
  OR2_X2     g25637(.A1(new_n28688_), .A2(new_n26604_), .Z(new_n28844_));
  OAI21_X1   g25638(.A1(new_n28844_), .A2(new_n28843_), .B(new_n27817_), .ZN(new_n28845_));
  AOI21_X1   g25639(.A1(new_n28842_), .A2(new_n28690_), .B(new_n28845_), .ZN(new_n28846_));
  OAI21_X1   g25640(.A1(new_n28840_), .A2(new_n27963_), .B(new_n28846_), .ZN(new_n28847_));
  NOR2_X1    g25641(.A1(new_n27611_), .A2(new_n28808_), .ZN(new_n28848_));
  NOR2_X1    g25642(.A1(new_n28848_), .A2(new_n26604_), .ZN(new_n28849_));
  NAND2_X1   g25643(.A1(new_n28728_), .A2(pi1151), .ZN(new_n28850_));
  AOI21_X1   g25644(.A1(new_n28724_), .A2(new_n27879_), .B(new_n27930_), .ZN(new_n28851_));
  NAND4_X1   g25645(.A1(new_n28850_), .A2(new_n28739_), .A3(new_n28849_), .A4(new_n28851_), .ZN(new_n28852_));
  OAI21_X1   g25646(.A1(new_n28820_), .A2(new_n28752_), .B(new_n26604_), .ZN(new_n28853_));
  NAND3_X1   g25647(.A1(new_n27817_), .A2(pi1151), .A3(pi1152), .ZN(new_n28854_));
  NOR2_X1    g25648(.A1(new_n28750_), .A2(new_n28854_), .ZN(new_n28855_));
  AOI21_X1   g25649(.A1(new_n28855_), .A2(new_n28853_), .B(pi1149), .ZN(new_n28856_));
  NAND2_X1   g25650(.A1(new_n27960_), .A2(new_n28779_), .ZN(new_n28857_));
  OAI21_X1   g25651(.A1(new_n28857_), .A2(new_n28682_), .B(new_n27929_), .ZN(new_n28858_));
  AOI21_X1   g25652(.A1(new_n28684_), .A2(new_n28814_), .B(new_n28858_), .ZN(new_n28859_));
  NAND2_X1   g25653(.A1(new_n28708_), .A2(pi1151), .ZN(new_n28860_));
  INV_X1     g25654(.I(new_n27936_), .ZN(new_n28861_));
  AOI21_X1   g25655(.A1(new_n28716_), .A2(new_n28861_), .B(pi1152), .ZN(new_n28862_));
  AOI21_X1   g25656(.A1(new_n28862_), .A2(new_n28860_), .B(new_n27817_), .ZN(new_n28863_));
  NOR2_X1    g25657(.A1(new_n28783_), .A2(new_n26604_), .ZN(new_n28864_));
  NOR4_X1    g25658(.A1(new_n28863_), .A2(new_n28717_), .A3(new_n28808_), .A4(new_n28864_), .ZN(new_n28865_));
  NOR2_X1    g25659(.A1(pi1148), .A2(pi1149), .ZN(new_n28866_));
  OAI21_X1   g25660(.A1(new_n28865_), .A2(new_n28859_), .B(new_n28866_), .ZN(new_n28867_));
  INV_X1     g25661(.I(new_n28764_), .ZN(new_n28868_));
  NAND2_X1   g25662(.A1(new_n28868_), .A2(new_n26604_), .ZN(new_n28869_));
  AOI21_X1   g25663(.A1(pi1151), .A2(new_n28731_), .B(new_n28869_), .ZN(new_n28870_));
  NOR4_X1    g25664(.A1(new_n28734_), .A2(pi1152), .A3(new_n28762_), .A4(new_n28808_), .ZN(new_n28871_));
  OAI21_X1   g25665(.A1(new_n28870_), .A2(new_n27817_), .B(new_n28871_), .ZN(new_n28872_));
  NAND2_X1   g25666(.A1(new_n28743_), .A2(new_n27251_), .ZN(new_n28873_));
  NAND2_X1   g25667(.A1(new_n28873_), .A2(new_n28757_), .ZN(new_n28874_));
  NOR2_X1    g25668(.A1(new_n27251_), .A2(pi1152), .ZN(new_n28875_));
  AOI21_X1   g25669(.A1(new_n28754_), .A2(new_n28875_), .B(new_n27930_), .ZN(new_n28876_));
  NAND2_X1   g25670(.A1(new_n28874_), .A2(new_n28876_), .ZN(new_n28877_));
  NOR3_X1    g25671(.A1(pi0213), .A2(pi1148), .A3(pi1149), .ZN(new_n28878_));
  NAND4_X1   g25672(.A1(new_n28872_), .A2(new_n28867_), .A3(new_n28877_), .A4(new_n28878_), .ZN(new_n28879_));
  AOI21_X1   g25673(.A1(new_n28852_), .A2(new_n28856_), .B(new_n28879_), .ZN(new_n28880_));
  AOI21_X1   g25674(.A1(new_n28880_), .A2(new_n28847_), .B(pi0209), .ZN(new_n28881_));
  NOR3_X1    g25675(.A1(new_n28604_), .A2(pi0213), .A3(new_n28881_), .ZN(new_n28882_));
  INV_X1     g25676(.I(new_n28848_), .ZN(new_n28883_));
  INV_X1     g25677(.I(new_n28864_), .ZN(new_n28884_));
  NAND2_X1   g25678(.A1(new_n27700_), .A2(pi1151), .ZN(new_n28885_));
  NAND4_X1   g25679(.A1(new_n28022_), .A2(new_n27929_), .A3(new_n28884_), .A4(new_n28885_), .ZN(new_n28886_));
  NOR4_X1    g25680(.A1(new_n28017_), .A2(pi1152), .A3(new_n27613_), .A4(new_n28873_), .ZN(new_n28887_));
  NAND2_X1   g25681(.A1(new_n27693_), .A2(new_n28875_), .ZN(new_n28888_));
  NAND2_X1   g25682(.A1(new_n28888_), .A2(new_n27817_), .ZN(new_n28889_));
  OAI22_X1   g25683(.A1(new_n28886_), .A2(new_n28883_), .B1(new_n28887_), .B2(new_n28889_), .ZN(new_n28890_));
  AOI21_X1   g25684(.A1(pi1152), .A2(new_n28732_), .B(new_n28773_), .ZN(new_n28891_));
  NAND2_X1   g25685(.A1(new_n28724_), .A2(new_n28784_), .ZN(new_n28892_));
  NOR2_X1    g25686(.A1(new_n28024_), .A2(new_n27512_), .ZN(new_n28893_));
  AOI21_X1   g25687(.A1(new_n28893_), .A2(new_n27695_), .B(pi1152), .ZN(new_n28894_));
  NAND2_X1   g25688(.A1(new_n28795_), .A2(new_n28894_), .ZN(new_n28895_));
  NAND2_X1   g25689(.A1(new_n28895_), .A2(pi1150), .ZN(new_n28896_));
  NAND2_X1   g25690(.A1(new_n28775_), .A2(pi1151), .ZN(new_n28897_));
  NAND3_X1   g25691(.A1(new_n27515_), .A2(new_n27817_), .A3(new_n26604_), .ZN(new_n28898_));
  NOR4_X1    g25692(.A1(new_n28884_), .A2(pi1151), .A3(new_n27698_), .A4(new_n28898_), .ZN(new_n28899_));
  NAND4_X1   g25693(.A1(new_n28896_), .A2(new_n28892_), .A3(new_n28897_), .A4(new_n28899_), .ZN(new_n28900_));
  NOR2_X1    g25694(.A1(new_n28900_), .A2(new_n28891_), .ZN(new_n28901_));
  INV_X1     g25695(.I(new_n28802_), .ZN(new_n28902_));
  AOI21_X1   g25696(.A1(new_n28902_), .A2(new_n27862_), .B(new_n26604_), .ZN(new_n28903_));
  AOI21_X1   g25697(.A1(new_n28780_), .A2(new_n28903_), .B(pi1150), .ZN(new_n28904_));
  OAI21_X1   g25698(.A1(pi1151), .A2(new_n28754_), .B(new_n28842_), .ZN(new_n28905_));
  NAND3_X1   g25699(.A1(new_n28684_), .A2(new_n26604_), .A3(new_n28797_), .ZN(new_n28906_));
  NOR2_X1    g25700(.A1(pi1151), .A2(pi1152), .ZN(new_n28907_));
  AOI21_X1   g25701(.A1(new_n28793_), .A2(new_n28907_), .B(new_n27817_), .ZN(new_n28908_));
  AOI21_X1   g25702(.A1(new_n28906_), .A2(new_n28908_), .B(pi1148), .ZN(new_n28909_));
  OAI21_X1   g25703(.A1(new_n28905_), .A2(new_n28904_), .B(new_n28909_), .ZN(new_n28910_));
  OAI21_X1   g25704(.A1(new_n28901_), .A2(new_n28910_), .B(pi1149), .ZN(new_n28911_));
  OR2_X2     g25705(.A1(new_n28712_), .A2(new_n28823_), .Z(new_n28912_));
  AOI21_X1   g25706(.A1(new_n28912_), .A2(new_n28868_), .B(new_n26604_), .ZN(new_n28913_));
  AND3_X2    g25707(.A1(new_n28571_), .A2(pi1151), .A3(new_n27621_), .Z(new_n28914_));
  OAI21_X1   g25708(.A1(new_n28914_), .A2(new_n28716_), .B(new_n26604_), .ZN(new_n28915_));
  NAND2_X1   g25709(.A1(new_n28915_), .A2(new_n27817_), .ZN(new_n28916_));
  OAI21_X1   g25710(.A1(new_n28913_), .A2(new_n28916_), .B(pi1148), .ZN(new_n28917_));
  NAND2_X1   g25711(.A1(new_n28883_), .A2(pi1152), .ZN(new_n28918_));
  NOR3_X1    g25712(.A1(new_n27633_), .A2(new_n27251_), .A3(new_n27598_), .ZN(new_n28919_));
  NOR3_X1    g25713(.A1(new_n28809_), .A2(new_n28919_), .A3(pi1152), .ZN(new_n28920_));
  OAI21_X1   g25714(.A1(new_n28918_), .A2(new_n28718_), .B(new_n28920_), .ZN(new_n28921_));
  NAND3_X1   g25715(.A1(new_n28921_), .A2(new_n28917_), .A3(pi1150), .ZN(new_n28922_));
  NOR2_X1    g25716(.A1(new_n28829_), .A2(new_n26604_), .ZN(new_n28923_));
  OAI21_X1   g25717(.A1(pi1151), .A2(new_n27613_), .B(new_n28923_), .ZN(new_n28924_));
  NAND4_X1   g25718(.A1(new_n28924_), .A2(new_n27817_), .A3(new_n27519_), .A4(new_n28875_), .ZN(new_n28925_));
  NAND2_X1   g25719(.A1(new_n27251_), .A2(new_n26604_), .ZN(new_n28926_));
  NOR2_X1    g25720(.A1(new_n28812_), .A2(new_n28926_), .ZN(new_n28927_));
  OAI21_X1   g25721(.A1(new_n28742_), .A2(pi1151), .B(new_n26604_), .ZN(new_n28928_));
  OAI21_X1   g25722(.A1(new_n28697_), .A2(new_n28928_), .B(pi1150), .ZN(new_n28929_));
  OAI21_X1   g25723(.A1(new_n28927_), .A2(new_n28929_), .B(new_n28925_), .ZN(new_n28930_));
  NAND2_X1   g25724(.A1(new_n28930_), .A2(new_n27515_), .ZN(new_n28931_));
  NAND4_X1   g25725(.A1(new_n28911_), .A2(new_n27470_), .A3(new_n28922_), .A4(new_n28931_), .ZN(new_n28932_));
  MUX2_X1    g25726(.I0(new_n28932_), .I1(new_n28890_), .S(pi0213), .Z(new_n28933_));
  AOI21_X1   g25727(.A1(new_n28933_), .A2(pi0209), .B(new_n28882_), .ZN(new_n28934_));
  MUX2_X1    g25728(.I0(new_n28934_), .I1(pi0248), .S(new_n26307_), .Z(po0405));
  NAND3_X1   g25729(.A1(new_n27195_), .A2(pi0299), .A3(new_n26723_), .ZN(new_n28936_));
  NOR2_X1    g25730(.A1(new_n26722_), .A2(new_n2587_), .ZN(new_n28937_));
  OAI21_X1   g25731(.A1(new_n27525_), .A2(pi0299), .B(new_n8078_), .ZN(new_n28938_));
  NOR2_X1    g25732(.A1(new_n27525_), .A2(new_n27390_), .ZN(new_n28939_));
  NOR3_X1    g25733(.A1(new_n28939_), .A2(new_n8078_), .A3(new_n27927_), .ZN(new_n28940_));
  AOI21_X1   g25734(.A1(new_n28937_), .A2(new_n28938_), .B(new_n28940_), .ZN(new_n28941_));
  AOI21_X1   g25735(.A1(new_n28941_), .A2(pi0212), .B(new_n28936_), .ZN(new_n28942_));
  INV_X1     g25736(.I(new_n28936_), .ZN(new_n28943_));
  NOR3_X1    g25737(.A1(new_n28941_), .A2(new_n28943_), .A3(new_n8076_), .ZN(new_n28944_));
  NOR3_X1    g25738(.A1(new_n28944_), .A2(new_n28942_), .A3(new_n8247_), .ZN(new_n28945_));
  AOI21_X1   g25739(.A1(pi0219), .A2(new_n27525_), .B(new_n28945_), .ZN(new_n28946_));
  NOR2_X1    g25740(.A1(new_n28946_), .A2(new_n5223_), .ZN(new_n28947_));
  NOR2_X1    g25741(.A1(new_n26723_), .A2(new_n2587_), .ZN(new_n28948_));
  AOI21_X1   g25742(.A1(new_n27194_), .A2(new_n2587_), .B(new_n28948_), .ZN(new_n28949_));
  NOR3_X1    g25743(.A1(new_n28949_), .A2(pi0214), .A3(new_n27194_), .ZN(new_n28950_));
  INV_X1     g25744(.I(new_n28949_), .ZN(new_n28951_));
  AOI21_X1   g25745(.A1(new_n8078_), .A2(new_n27194_), .B(new_n28951_), .ZN(new_n28952_));
  OAI21_X1   g25746(.A1(new_n26359_), .A2(pi0211), .B(new_n26361_), .ZN(new_n28953_));
  OAI21_X1   g25747(.A1(new_n27194_), .A2(new_n28953_), .B(new_n8078_), .ZN(new_n28954_));
  NOR4_X1    g25748(.A1(new_n27194_), .A2(new_n8247_), .A3(new_n5224_), .A4(new_n27607_), .ZN(new_n28955_));
  OAI21_X1   g25749(.A1(new_n28951_), .A2(new_n28954_), .B(new_n28955_), .ZN(new_n28956_));
  NOR3_X1    g25750(.A1(new_n28952_), .A2(new_n28950_), .A3(new_n28956_), .ZN(new_n28957_));
  NAND2_X1   g25751(.A1(new_n26728_), .A2(new_n5223_), .ZN(new_n28958_));
  NAND3_X1   g25752(.A1(new_n28958_), .A2(new_n5055_), .A3(pi1151), .ZN(new_n28959_));
  NOR3_X1    g25753(.A1(pi0057), .A2(pi1151), .A3(pi1152), .ZN(new_n28960_));
  NAND2_X1   g25754(.A1(new_n28958_), .A2(new_n28960_), .ZN(new_n28961_));
  AOI21_X1   g25755(.A1(new_n5055_), .A2(new_n26728_), .B(new_n28961_), .ZN(new_n28962_));
  OAI21_X1   g25756(.A1(new_n28957_), .A2(new_n28959_), .B(new_n28962_), .ZN(new_n28963_));
  NOR3_X1    g25757(.A1(new_n26723_), .A2(new_n2587_), .A3(new_n8248_), .ZN(new_n28964_));
  NOR2_X1    g25758(.A1(new_n27934_), .A2(new_n27658_), .ZN(new_n28965_));
  OAI21_X1   g25759(.A1(new_n26742_), .A2(new_n28964_), .B(new_n28965_), .ZN(new_n28966_));
  AOI21_X1   g25760(.A1(new_n27632_), .A2(new_n28583_), .B(new_n27251_), .ZN(new_n28967_));
  OAI21_X1   g25761(.A1(pi0211), .A2(new_n26529_), .B(new_n27575_), .ZN(new_n28968_));
  INV_X1     g25762(.I(new_n28937_), .ZN(new_n28969_));
  AOI21_X1   g25763(.A1(new_n27575_), .A2(new_n28969_), .B(pi0214), .ZN(new_n28970_));
  AOI21_X1   g25764(.A1(pi0214), .A2(new_n28968_), .B(new_n28970_), .ZN(new_n28971_));
  INV_X1     g25765(.I(new_n28971_), .ZN(new_n28972_));
  NAND2_X1   g25766(.A1(new_n27849_), .A2(new_n28969_), .ZN(new_n28973_));
  NAND2_X1   g25767(.A1(new_n28973_), .A2(new_n8247_), .ZN(new_n28974_));
  AOI21_X1   g25768(.A1(new_n28974_), .A2(new_n27269_), .B(pi0212), .ZN(new_n28975_));
  AOI21_X1   g25769(.A1(new_n28975_), .A2(new_n28972_), .B(pi1151), .ZN(new_n28976_));
  AOI22_X1   g25770(.A1(new_n27609_), .A2(new_n28976_), .B1(new_n28966_), .B2(new_n28967_), .ZN(new_n28977_));
  NOR3_X1    g25771(.A1(new_n28977_), .A2(pi1150), .A3(new_n26746_), .ZN(new_n28978_));
  OAI21_X1   g25772(.A1(new_n28947_), .A2(new_n28963_), .B(new_n28978_), .ZN(new_n28979_));
  NOR2_X1    g25773(.A1(new_n28002_), .A2(new_n26704_), .ZN(new_n28980_));
  NOR2_X1    g25774(.A1(new_n28002_), .A2(new_n8250_), .ZN(new_n28981_));
  NOR2_X1    g25775(.A1(new_n27669_), .A2(new_n26732_), .ZN(new_n28982_));
  NAND2_X1   g25776(.A1(new_n27682_), .A2(new_n26554_), .ZN(new_n28983_));
  NOR4_X1    g25777(.A1(new_n28980_), .A2(new_n28981_), .A3(new_n28983_), .A4(new_n28982_), .ZN(new_n28984_));
  NOR2_X1    g25778(.A1(new_n27690_), .A2(new_n27251_), .ZN(new_n28985_));
  OAI21_X1   g25779(.A1(new_n28984_), .A2(pi0219), .B(new_n28985_), .ZN(new_n28986_));
  OAI21_X1   g25780(.A1(new_n27236_), .A2(new_n28964_), .B(new_n26724_), .ZN(new_n28987_));
  NOR2_X1    g25781(.A1(new_n27818_), .A2(new_n28987_), .ZN(new_n28988_));
  NOR2_X1    g25782(.A1(new_n26730_), .A2(new_n28988_), .ZN(new_n28989_));
  AOI21_X1   g25783(.A1(new_n27232_), .A2(new_n8076_), .B(pi0219), .ZN(new_n28990_));
  NOR4_X1    g25784(.A1(new_n27549_), .A2(pi0212), .A3(new_n2587_), .A4(new_n26723_), .ZN(new_n28991_));
  AOI22_X1   g25785(.A1(new_n27994_), .A2(new_n28991_), .B1(new_n28973_), .B2(new_n28990_), .ZN(new_n28992_));
  INV_X1     g25786(.I(new_n28992_), .ZN(new_n28993_));
  NOR3_X1    g25787(.A1(new_n26746_), .A2(pi1151), .A3(new_n28988_), .ZN(new_n28994_));
  NAND2_X1   g25788(.A1(new_n27543_), .A2(new_n27252_), .ZN(new_n28995_));
  AOI21_X1   g25789(.A1(new_n28760_), .A2(new_n28994_), .B(new_n28995_), .ZN(new_n28996_));
  AOI21_X1   g25790(.A1(new_n28993_), .A2(new_n28996_), .B(pi1150), .ZN(new_n28997_));
  INV_X1     g25791(.I(new_n28997_), .ZN(new_n28998_));
  AOI21_X1   g25792(.A1(new_n28986_), .A2(new_n28989_), .B(new_n28998_), .ZN(new_n28999_));
  AND2_X2    g25793(.A1(new_n28999_), .A2(new_n28979_), .Z(new_n29000_));
  NOR3_X1    g25794(.A1(new_n29000_), .A2(new_n28890_), .A3(pi0213), .ZN(new_n29001_));
  INV_X1     g25795(.I(new_n29000_), .ZN(new_n29002_));
  AOI21_X1   g25796(.A1(new_n28890_), .A2(new_n24753_), .B(new_n29002_), .ZN(new_n29003_));
  NOR3_X1    g25797(.A1(new_n29003_), .A2(pi0209), .A3(new_n29001_), .ZN(new_n29004_));
  MUX2_X1    g25798(.I0(new_n29004_), .I1(pi0249), .S(new_n26307_), .Z(po0406));
  NOR3_X1    g25799(.A1(new_n6967_), .A2(pi0087), .A3(pi0250), .ZN(po0407));
  NAND3_X1   g25800(.A1(pi0199), .A2(pi0200), .A3(pi0476), .ZN(new_n29007_));
  INV_X1     g25801(.I(new_n29007_), .ZN(new_n29008_));
  NAND2_X1   g25802(.A1(new_n29008_), .A2(pi0251), .ZN(new_n29009_));
  OAI21_X1   g25803(.A1(pi0200), .A2(pi1053), .B(pi1039), .ZN(new_n29010_));
  INV_X1     g25804(.I(pi1039), .ZN(new_n29011_));
  NAND3_X1   g25805(.A1(new_n8098_), .A2(new_n29011_), .A3(pi1053), .ZN(new_n29012_));
  NAND4_X1   g25806(.A1(new_n29012_), .A2(new_n8094_), .A3(new_n29007_), .A4(new_n29010_), .ZN(new_n29013_));
  NAND2_X1   g25807(.A1(new_n29013_), .A2(new_n29009_), .ZN(po0408));
  NOR2_X1    g25808(.A1(pi0979), .A2(pi0984), .ZN(new_n29015_));
  NAND4_X1   g25809(.A1(new_n29015_), .A2(pi0835), .A3(pi0950), .A4(pi1001), .ZN(new_n29016_));
  NOR4_X1    g25810(.A1(new_n15500_), .A2(new_n5117_), .A3(new_n8533_), .A4(new_n29016_), .ZN(new_n29017_));
  NAND3_X1   g25811(.A1(new_n26267_), .A2(new_n5358_), .A3(new_n29017_), .ZN(new_n29018_));
  NOR2_X1    g25812(.A1(pi0057), .A2(pi0252), .ZN(new_n29019_));
  NAND3_X1   g25813(.A1(pi0057), .A2(pi0252), .A3(pi1092), .ZN(new_n29020_));
  OAI21_X1   g25814(.A1(new_n6953_), .A2(new_n29020_), .B(new_n2923_), .ZN(new_n29021_));
  AOI21_X1   g25815(.A1(new_n29018_), .A2(new_n29019_), .B(new_n29021_), .ZN(new_n29022_));
  NOR2_X1    g25816(.A1(new_n6446_), .A2(new_n8736_), .ZN(new_n29023_));
  NOR2_X1    g25817(.A1(new_n29016_), .A2(new_n5114_), .ZN(new_n29024_));
  AOI21_X1   g25818(.A1(new_n5358_), .A2(new_n29024_), .B(pi0252), .ZN(new_n29025_));
  NOR4_X1    g25819(.A1(new_n26203_), .A2(new_n2923_), .A3(pi1093), .A4(new_n29025_), .ZN(new_n29026_));
  AOI21_X1   g25820(.A1(new_n29026_), .A2(new_n6446_), .B(new_n29023_), .ZN(new_n29027_));
  NOR2_X1    g25821(.A1(new_n5143_), .A2(new_n8736_), .ZN(new_n29028_));
  AOI21_X1   g25822(.A1(new_n29026_), .A2(new_n5143_), .B(new_n29028_), .ZN(new_n29029_));
  MUX2_X1    g25823(.I0(new_n29029_), .I1(new_n29027_), .S(new_n6445_), .Z(new_n29030_));
  NAND2_X1   g25824(.A1(new_n29027_), .A2(new_n6460_), .ZN(new_n29031_));
  AOI21_X1   g25825(.A1(new_n29029_), .A2(new_n5141_), .B(pi0299), .ZN(new_n29032_));
  AOI21_X1   g25826(.A1(new_n29032_), .A2(new_n29031_), .B(new_n8371_), .ZN(new_n29033_));
  OAI21_X1   g25827(.A1(new_n2587_), .A2(new_n29030_), .B(new_n29033_), .ZN(new_n29034_));
  AOI21_X1   g25828(.A1(new_n8371_), .A2(new_n8736_), .B(new_n6953_), .ZN(new_n29035_));
  AOI21_X1   g25829(.A1(new_n29034_), .A2(new_n29035_), .B(new_n29022_), .ZN(po0409));
  OAI21_X1   g25830(.A1(new_n8269_), .A2(pi1153), .B(new_n27258_), .ZN(new_n29037_));
  NAND2_X1   g25831(.A1(new_n29037_), .A2(new_n9658_), .ZN(new_n29038_));
  AOI21_X1   g25832(.A1(new_n26641_), .A2(new_n26389_), .B(new_n8077_), .ZN(new_n29039_));
  XOR2_X1    g25833(.A1(new_n29038_), .A2(new_n29039_), .Z(new_n29040_));
  NOR2_X1    g25834(.A1(new_n8169_), .A2(pi1153), .ZN(new_n29041_));
  NOR4_X1    g25835(.A1(po1038), .A2(new_n26379_), .A3(new_n26355_), .A4(new_n29041_), .ZN(new_n29042_));
  NAND2_X1   g25836(.A1(new_n29040_), .A2(new_n29042_), .ZN(new_n29043_));
  NOR3_X1    g25837(.A1(new_n26961_), .A2(pi1151), .A3(new_n8663_), .ZN(new_n29044_));
  NOR3_X1    g25838(.A1(new_n26431_), .A2(new_n26370_), .A3(new_n27246_), .ZN(new_n29045_));
  INV_X1     g25839(.I(new_n29045_), .ZN(new_n29046_));
  NOR3_X1    g25840(.A1(po1038), .A2(new_n29046_), .A3(new_n26355_), .ZN(new_n29047_));
  INV_X1     g25841(.I(new_n26355_), .ZN(new_n29048_));
  AOI21_X1   g25842(.A1(new_n6845_), .A2(new_n29046_), .B(new_n29048_), .ZN(new_n29049_));
  NOR2_X1    g25843(.A1(new_n29047_), .A2(new_n29049_), .ZN(new_n29050_));
  NAND2_X1   g25844(.A1(new_n29050_), .A2(pi1153), .ZN(new_n29051_));
  AOI22_X1   g25845(.A1(new_n29051_), .A2(new_n27251_), .B1(new_n29043_), .B2(new_n29044_), .ZN(new_n29052_));
  INV_X1     g25846(.I(new_n8665_), .ZN(new_n29053_));
  NAND4_X1   g25847(.A1(new_n6845_), .A2(new_n27251_), .A3(new_n29053_), .A4(new_n26355_), .ZN(new_n29054_));
  NOR3_X1    g25848(.A1(new_n26370_), .A2(new_n27251_), .A3(new_n8169_), .ZN(new_n29055_));
  NOR2_X1    g25849(.A1(new_n27390_), .A2(new_n26389_), .ZN(new_n29056_));
  INV_X1     g25850(.I(new_n29056_), .ZN(new_n29057_));
  NAND2_X1   g25851(.A1(new_n29057_), .A2(pi1153), .ZN(new_n29058_));
  NOR2_X1    g25852(.A1(new_n27145_), .A2(new_n26542_), .ZN(new_n29059_));
  OAI21_X1   g25853(.A1(new_n29055_), .A2(new_n29058_), .B(new_n29059_), .ZN(new_n29060_));
  NAND2_X1   g25854(.A1(new_n27251_), .A2(pi1153), .ZN(new_n29061_));
  AOI21_X1   g25855(.A1(new_n11893_), .A2(pi1151), .B(pi0211), .ZN(new_n29062_));
  AOI21_X1   g25856(.A1(new_n29062_), .A2(new_n29061_), .B(pi0219), .ZN(new_n29063_));
  XNOR2_X1   g25857(.A1(new_n29063_), .A2(new_n26721_), .ZN(new_n29064_));
  OAI22_X1   g25858(.A1(new_n29060_), .A2(new_n29054_), .B1(new_n6845_), .B2(new_n29064_), .ZN(new_n29065_));
  MUX2_X1    g25859(.I0(new_n29065_), .I1(new_n29052_), .S(new_n26604_), .Z(new_n29066_));
  NAND2_X1   g25860(.A1(new_n29066_), .A2(pi0230), .ZN(new_n29067_));
  NOR2_X1    g25861(.A1(new_n2918_), .A2(pi0299), .ZN(new_n29068_));
  INV_X1     g25862(.I(new_n29068_), .ZN(new_n29069_));
  NOR4_X1    g25863(.A1(new_n26542_), .A2(pi0253), .A3(new_n8664_), .A4(new_n29069_), .ZN(new_n29070_));
  NOR2_X1    g25864(.A1(new_n26433_), .A2(new_n29069_), .ZN(new_n29071_));
  INV_X1     g25865(.I(new_n29071_), .ZN(new_n29072_));
  NOR3_X1    g25866(.A1(new_n29072_), .A2(pi1153), .A3(new_n26355_), .ZN(new_n29073_));
  NOR2_X1    g25867(.A1(new_n8662_), .A2(new_n2918_), .ZN(new_n29074_));
  OAI21_X1   g25868(.A1(pi1153), .A2(new_n29074_), .B(new_n29073_), .ZN(new_n29075_));
  NOR2_X1    g25869(.A1(new_n2918_), .A2(pi0211), .ZN(new_n29076_));
  INV_X1     g25870(.I(new_n29076_), .ZN(new_n29077_));
  AOI21_X1   g25871(.A1(new_n26543_), .A2(new_n2587_), .B(new_n29077_), .ZN(new_n29078_));
  NOR2_X1    g25872(.A1(new_n27145_), .A2(new_n2918_), .ZN(new_n29079_));
  NOR2_X1    g25873(.A1(new_n26380_), .A2(new_n2918_), .ZN(new_n29080_));
  NAND2_X1   g25874(.A1(new_n29080_), .A2(new_n26609_), .ZN(new_n29081_));
  NAND2_X1   g25875(.A1(new_n29081_), .A2(new_n26355_), .ZN(new_n29082_));
  OAI21_X1   g25876(.A1(new_n29079_), .A2(new_n29082_), .B(new_n28261_), .ZN(new_n29083_));
  OAI22_X1   g25877(.A1(new_n29083_), .A2(new_n29078_), .B1(new_n29070_), .B2(new_n29075_), .ZN(new_n29084_));
  NOR2_X1    g25878(.A1(pi0253), .A2(pi1091), .ZN(new_n29085_));
  NOR2_X1    g25879(.A1(new_n27660_), .A2(new_n9658_), .ZN(new_n29086_));
  INV_X1     g25880(.I(new_n29086_), .ZN(new_n29087_));
  NOR2_X1    g25881(.A1(new_n29087_), .A2(new_n29085_), .ZN(new_n29088_));
  OAI21_X1   g25882(.A1(new_n26542_), .A2(new_n2918_), .B(new_n29088_), .ZN(new_n29089_));
  NAND2_X1   g25883(.A1(new_n29084_), .A2(new_n29089_), .ZN(new_n29090_));
  NOR2_X1    g25884(.A1(new_n26960_), .A2(new_n2918_), .ZN(new_n29091_));
  NOR3_X1    g25885(.A1(new_n6845_), .A2(new_n29085_), .A3(new_n29091_), .ZN(new_n29092_));
  INV_X1     g25886(.I(new_n29085_), .ZN(new_n29093_));
  NOR2_X1    g25887(.A1(new_n29057_), .A2(pi1153), .ZN(new_n29094_));
  AOI21_X1   g25888(.A1(new_n29056_), .A2(new_n28261_), .B(pi1091), .ZN(new_n29095_));
  NOR2_X1    g25889(.A1(new_n26370_), .A2(new_n8169_), .ZN(new_n29096_));
  OAI21_X1   g25890(.A1(new_n29094_), .A2(new_n29095_), .B(new_n29096_), .ZN(new_n29097_));
  AOI21_X1   g25891(.A1(new_n29097_), .A2(new_n6845_), .B(new_n29093_), .ZN(new_n29098_));
  NOR4_X1    g25892(.A1(new_n29092_), .A2(pi0219), .A3(pi1152), .A4(new_n29077_), .ZN(new_n29099_));
  NOR2_X1    g25893(.A1(new_n29099_), .A2(new_n27251_), .ZN(new_n29100_));
  OAI21_X1   g25894(.A1(new_n29092_), .A2(new_n29098_), .B(new_n29100_), .ZN(new_n29101_));
  NAND3_X1   g25895(.A1(new_n29090_), .A2(new_n27818_), .A3(new_n29101_), .ZN(new_n29102_));
  AOI21_X1   g25896(.A1(new_n26606_), .A2(pi1091), .B(pi1153), .ZN(new_n29103_));
  NOR2_X1    g25897(.A1(new_n29080_), .A2(new_n11893_), .ZN(new_n29104_));
  NOR3_X1    g25898(.A1(new_n29103_), .A2(new_n29048_), .A3(new_n29104_), .ZN(new_n29105_));
  AOI21_X1   g25899(.A1(new_n29040_), .A2(pi1091), .B(new_n29105_), .ZN(new_n29106_));
  NAND2_X1   g25900(.A1(new_n29058_), .A2(new_n9660_), .ZN(new_n29107_));
  AOI21_X1   g25901(.A1(new_n29107_), .A2(pi1091), .B(pi0253), .ZN(new_n29108_));
  AOI21_X1   g25902(.A1(new_n11893_), .A2(pi0219), .B(pi0211), .ZN(new_n29109_));
  NOR4_X1    g25903(.A1(new_n6845_), .A2(new_n2918_), .A3(new_n29085_), .A4(new_n29109_), .ZN(new_n29110_));
  NOR3_X1    g25904(.A1(new_n29110_), .A2(new_n28261_), .A3(pi1151), .ZN(new_n29111_));
  OAI21_X1   g25905(.A1(new_n29108_), .A2(po1038), .B(new_n29111_), .ZN(new_n29112_));
  NOR2_X1    g25906(.A1(new_n2918_), .A2(new_n11893_), .ZN(new_n29113_));
  INV_X1     g25907(.I(new_n29113_), .ZN(new_n29114_));
  NOR3_X1    g25908(.A1(po1038), .A2(new_n29046_), .A3(new_n29114_), .ZN(new_n29115_));
  NOR2_X1    g25909(.A1(new_n28261_), .A2(pi1091), .ZN(new_n29116_));
  NOR4_X1    g25910(.A1(new_n29115_), .A2(new_n8247_), .A3(pi1151), .A4(new_n29116_), .ZN(new_n29117_));
  AOI21_X1   g25911(.A1(new_n29117_), .A2(new_n29092_), .B(pi1152), .ZN(new_n29118_));
  OAI21_X1   g25912(.A1(new_n29112_), .A2(new_n29106_), .B(new_n29118_), .ZN(new_n29119_));
  AOI21_X1   g25913(.A1(new_n29102_), .A2(new_n28287_), .B(new_n29119_), .ZN(new_n29120_));
  NOR2_X1    g25914(.A1(new_n28172_), .A2(new_n28156_), .ZN(new_n29121_));
  NOR2_X1    g25915(.A1(new_n29121_), .A2(pi1153), .ZN(new_n29122_));
  NOR2_X1    g25916(.A1(new_n28143_), .A2(new_n28156_), .ZN(new_n29123_));
  INV_X1     g25917(.I(new_n29123_), .ZN(new_n29124_));
  AOI21_X1   g25918(.A1(new_n8077_), .A2(new_n28135_), .B(new_n29124_), .ZN(new_n29125_));
  INV_X1     g25919(.I(new_n29125_), .ZN(new_n29126_));
  NOR3_X1    g25920(.A1(new_n29126_), .A2(new_n28149_), .A3(new_n29122_), .ZN(new_n29127_));
  INV_X1     g25921(.I(new_n28238_), .ZN(new_n29128_));
  NOR2_X1    g25922(.A1(new_n29128_), .A2(new_n28139_), .ZN(new_n29129_));
  INV_X1     g25923(.I(new_n29129_), .ZN(new_n29130_));
  NOR2_X1    g25924(.A1(new_n29130_), .A2(pi0211), .ZN(new_n29131_));
  NOR2_X1    g25925(.A1(new_n29131_), .A2(new_n28150_), .ZN(new_n29132_));
  INV_X1     g25926(.I(new_n29132_), .ZN(new_n29133_));
  AOI21_X1   g25927(.A1(new_n29133_), .A2(pi1153), .B(new_n28240_), .ZN(new_n29134_));
  NOR2_X1    g25928(.A1(new_n29134_), .A2(new_n28143_), .ZN(new_n29135_));
  MUX2_X1    g25929(.I0(new_n29135_), .I1(new_n29127_), .S(new_n8247_), .Z(new_n29136_));
  NOR3_X1    g25930(.A1(new_n29126_), .A2(new_n28129_), .A3(new_n28174_), .ZN(new_n29137_));
  NOR2_X1    g25931(.A1(new_n29137_), .A2(new_n28246_), .ZN(new_n29138_));
  NAND2_X1   g25932(.A1(new_n28224_), .A2(pi0219), .ZN(new_n29139_));
  NAND2_X1   g25933(.A1(new_n29139_), .A2(new_n11893_), .ZN(new_n29140_));
  INV_X1     g25934(.I(new_n29131_), .ZN(new_n29141_));
  NOR2_X1    g25935(.A1(new_n28120_), .A2(pi0219), .ZN(new_n29142_));
  INV_X1     g25936(.I(new_n29142_), .ZN(new_n29143_));
  AOI21_X1   g25937(.A1(new_n29141_), .A2(new_n28167_), .B(new_n29143_), .ZN(new_n29144_));
  INV_X1     g25938(.I(new_n29144_), .ZN(new_n29145_));
  NOR2_X1    g25939(.A1(new_n28129_), .A2(new_n28172_), .ZN(new_n29146_));
  NOR2_X1    g25940(.A1(new_n29146_), .A2(new_n29122_), .ZN(new_n29147_));
  OAI22_X1   g25941(.A1(new_n29145_), .A2(new_n29147_), .B1(new_n29138_), .B2(new_n29140_), .ZN(new_n29148_));
  MUX2_X1    g25942(.I0(new_n29148_), .I1(new_n29136_), .S(new_n28261_), .Z(new_n29149_));
  MUX2_X1    g25943(.I0(new_n29137_), .I1(new_n28238_), .S(new_n11893_), .Z(new_n29150_));
  INV_X1     g25944(.I(new_n28195_), .ZN(new_n29151_));
  NAND2_X1   g25945(.A1(new_n29151_), .A2(new_n11893_), .ZN(new_n29152_));
  OAI21_X1   g25946(.A1(new_n28167_), .A2(new_n28180_), .B(pi1153), .ZN(new_n29153_));
  AND2_X2    g25947(.A1(new_n29153_), .A2(new_n8247_), .Z(new_n29154_));
  OAI21_X1   g25948(.A1(new_n29154_), .A2(new_n29152_), .B(pi0253), .ZN(new_n29155_));
  AOI21_X1   g25949(.A1(new_n29150_), .A2(pi0219), .B(new_n29155_), .ZN(new_n29156_));
  INV_X1     g25950(.I(new_n28194_), .ZN(new_n29157_));
  AOI21_X1   g25951(.A1(new_n11893_), .A2(new_n29157_), .B(new_n28158_), .ZN(new_n29158_));
  NOR3_X1    g25952(.A1(new_n28157_), .A2(pi1153), .A3(new_n29157_), .ZN(new_n29159_));
  NOR3_X1    g25953(.A1(new_n29158_), .A2(pi0219), .A3(new_n29159_), .ZN(new_n29160_));
  NAND2_X1   g25954(.A1(new_n29134_), .A2(pi0219), .ZN(new_n29161_));
  NAND3_X1   g25955(.A1(new_n29161_), .A2(new_n29160_), .A3(new_n28261_), .ZN(new_n29162_));
  OAI21_X1   g25956(.A1(new_n29162_), .A2(new_n29156_), .B(new_n6845_), .ZN(new_n29163_));
  INV_X1     g25957(.I(new_n29091_), .ZN(new_n29164_));
  MUX2_X1    g25958(.I0(new_n28146_), .I1(new_n28140_), .S(new_n8077_), .Z(new_n29165_));
  NOR2_X1    g25959(.A1(new_n29165_), .A2(new_n8247_), .ZN(new_n29166_));
  NOR2_X1    g25960(.A1(new_n28117_), .A2(pi0219), .ZN(new_n29167_));
  NOR2_X1    g25961(.A1(new_n29166_), .A2(new_n29167_), .ZN(new_n29168_));
  NAND2_X1   g25962(.A1(new_n29168_), .A2(new_n29164_), .ZN(new_n29169_));
  INV_X1     g25963(.I(new_n28146_), .ZN(new_n29170_));
  NAND3_X1   g25964(.A1(new_n29143_), .A2(new_n29170_), .A3(new_n29164_), .ZN(new_n29171_));
  MUX2_X1    g25965(.I0(new_n29171_), .I1(new_n29169_), .S(new_n28261_), .Z(new_n29172_));
  NOR2_X1    g25966(.A1(new_n29172_), .A2(new_n6845_), .ZN(new_n29173_));
  AOI21_X1   g25967(.A1(new_n8077_), .A2(new_n28116_), .B(new_n29143_), .ZN(new_n29174_));
  NOR4_X1    g25968(.A1(new_n29174_), .A2(pi0219), .A3(new_n6845_), .A4(new_n28108_), .ZN(new_n29175_));
  NOR3_X1    g25969(.A1(new_n29173_), .A2(new_n27251_), .A3(new_n29175_), .ZN(new_n29176_));
  NAND3_X1   g25970(.A1(new_n29163_), .A2(new_n27251_), .A3(new_n29176_), .ZN(new_n29177_));
  AOI21_X1   g25971(.A1(new_n29149_), .A2(new_n6845_), .B(new_n29177_), .ZN(new_n29178_));
  OAI21_X1   g25972(.A1(pi0211), .A2(new_n28108_), .B(new_n29167_), .ZN(new_n29179_));
  INV_X1     g25973(.I(new_n29179_), .ZN(new_n29180_));
  NOR2_X1    g25974(.A1(new_n29143_), .A2(new_n29180_), .ZN(new_n29181_));
  NAND2_X1   g25975(.A1(new_n28108_), .A2(new_n26351_), .ZN(new_n29182_));
  NOR2_X1    g25976(.A1(new_n29181_), .A2(new_n29182_), .ZN(new_n29183_));
  AOI21_X1   g25977(.A1(new_n29183_), .A2(new_n28140_), .B(new_n26604_), .ZN(new_n29184_));
  OAI21_X1   g25978(.A1(new_n29172_), .A2(new_n6845_), .B(new_n29184_), .ZN(new_n29185_));
  NAND2_X1   g25979(.A1(new_n29144_), .A2(new_n29160_), .ZN(new_n29186_));
  OR2_X2     g25980(.A1(new_n29134_), .A2(new_n8247_), .Z(new_n29187_));
  AOI21_X1   g25981(.A1(new_n29187_), .A2(new_n29186_), .B(new_n28139_), .ZN(new_n29188_));
  NOR2_X1    g25982(.A1(new_n29137_), .A2(new_n28250_), .ZN(new_n29189_));
  NOR2_X1    g25983(.A1(new_n28231_), .A2(pi1153), .ZN(new_n29190_));
  NAND4_X1   g25984(.A1(new_n29189_), .A2(pi0219), .A3(pi1153), .A4(new_n29190_), .ZN(new_n29191_));
  NOR2_X1    g25985(.A1(new_n29126_), .A2(new_n29143_), .ZN(new_n29192_));
  INV_X1     g25986(.I(new_n29192_), .ZN(new_n29193_));
  NOR2_X1    g25987(.A1(new_n28179_), .A2(new_n11893_), .ZN(new_n29194_));
  NAND2_X1   g25988(.A1(new_n29193_), .A2(new_n29194_), .ZN(new_n29195_));
  NAND2_X1   g25989(.A1(new_n29191_), .A2(new_n29195_), .ZN(new_n29196_));
  MUX2_X1    g25990(.I0(new_n29196_), .I1(new_n29188_), .S(new_n28261_), .Z(new_n29197_));
  NOR2_X1    g25991(.A1(new_n29174_), .A2(pi0219), .ZN(new_n29198_));
  NOR2_X1    g25992(.A1(po1038), .A2(pi1151), .ZN(new_n29199_));
  NOR2_X1    g25993(.A1(new_n29134_), .A2(new_n28126_), .ZN(new_n29200_));
  INV_X1     g25994(.I(new_n29138_), .ZN(new_n29201_));
  NOR2_X1    g25995(.A1(new_n28240_), .A2(pi1091), .ZN(new_n29202_));
  NOR2_X1    g25996(.A1(new_n29202_), .A2(pi1153), .ZN(new_n29203_));
  INV_X1     g25997(.I(new_n29121_), .ZN(new_n29204_));
  NOR2_X1    g25998(.A1(new_n29204_), .A2(pi0219), .ZN(new_n29205_));
  OR3_X2     g25999(.A1(new_n29203_), .A2(pi0253), .A3(new_n29205_), .Z(new_n29206_));
  NOR2_X1    g26000(.A1(new_n28175_), .A2(pi1153), .ZN(new_n29207_));
  NOR2_X1    g26001(.A1(new_n29207_), .A2(new_n28139_), .ZN(new_n29208_));
  INV_X1     g26002(.I(new_n29208_), .ZN(new_n29209_));
  NOR2_X1    g26003(.A1(new_n29151_), .A2(pi0219), .ZN(new_n29210_));
  INV_X1     g26004(.I(new_n29210_), .ZN(new_n29211_));
  NOR2_X1    g26005(.A1(new_n29211_), .A2(new_n29209_), .ZN(new_n29212_));
  NOR4_X1    g26006(.A1(new_n29212_), .A2(pi0219), .A3(pi0253), .A4(po1038), .ZN(new_n29213_));
  OAI21_X1   g26007(.A1(new_n29201_), .A2(new_n29206_), .B(new_n29213_), .ZN(new_n29214_));
  NOR2_X1    g26008(.A1(new_n29173_), .A2(new_n28837_), .ZN(new_n29215_));
  OAI21_X1   g26009(.A1(new_n29200_), .A2(new_n29214_), .B(new_n29215_), .ZN(new_n29216_));
  AOI21_X1   g26010(.A1(new_n29197_), .A2(new_n29199_), .B(new_n29216_), .ZN(new_n29217_));
  OAI21_X1   g26011(.A1(new_n29178_), .A2(new_n29185_), .B(new_n29217_), .ZN(new_n29218_));
  AOI21_X1   g26012(.A1(new_n29218_), .A2(new_n28286_), .B(new_n29120_), .ZN(new_n29219_));
  OAI21_X1   g26013(.A1(new_n29219_), .A2(pi0230), .B(new_n29067_), .ZN(po0410));
  NOR3_X1    g26014(.A1(new_n26434_), .A2(new_n11950_), .A3(new_n26707_), .ZN(new_n29221_));
  OAI21_X1   g26015(.A1(new_n29221_), .A2(new_n26712_), .B(new_n8663_), .ZN(new_n29222_));
  NAND3_X1   g26016(.A1(new_n8077_), .A2(new_n2587_), .A3(pi0219), .ZN(new_n29223_));
  OAI22_X1   g26017(.A1(new_n26610_), .A2(new_n29223_), .B1(pi1154), .B2(new_n26638_), .ZN(new_n29224_));
  NAND3_X1   g26018(.A1(new_n29224_), .A2(new_n29222_), .A3(new_n6845_), .ZN(new_n29225_));
  AOI21_X1   g26019(.A1(new_n8664_), .A2(new_n29048_), .B(new_n26723_), .ZN(new_n29226_));
  NAND2_X1   g26020(.A1(po1038), .A2(new_n29226_), .ZN(new_n29227_));
  AOI21_X1   g26021(.A1(new_n29225_), .A2(new_n26604_), .B(new_n29227_), .ZN(new_n29228_));
  OAI21_X1   g26022(.A1(new_n26404_), .A2(new_n26707_), .B(new_n26963_), .ZN(new_n29229_));
  NAND2_X1   g26023(.A1(new_n26672_), .A2(new_n11950_), .ZN(new_n29230_));
  AOI21_X1   g26024(.A1(new_n26642_), .A2(new_n29229_), .B(new_n29230_), .ZN(new_n29231_));
  NAND2_X1   g26025(.A1(new_n29231_), .A2(new_n8247_), .ZN(new_n29232_));
  OAI21_X1   g26026(.A1(pi0219), .A2(pi1153), .B(new_n8077_), .ZN(new_n29233_));
  NOR2_X1    g26027(.A1(new_n27439_), .A2(new_n29233_), .ZN(new_n29234_));
  NAND2_X1   g26028(.A1(new_n8098_), .A2(pi1154), .ZN(new_n29235_));
  AOI22_X1   g26029(.A1(new_n27622_), .A2(new_n26707_), .B1(new_n8626_), .B2(new_n29235_), .ZN(new_n29236_));
  NOR2_X1    g26030(.A1(new_n29236_), .A2(pi0219), .ZN(new_n29237_));
  NOR3_X1    g26031(.A1(new_n29234_), .A2(po1038), .A3(new_n29237_), .ZN(new_n29238_));
  AOI21_X1   g26032(.A1(new_n29238_), .A2(new_n29232_), .B(pi1152), .ZN(new_n29239_));
  OAI21_X1   g26033(.A1(new_n29228_), .A2(new_n29239_), .B(pi0230), .ZN(new_n29240_));
  AOI21_X1   g26034(.A1(new_n26610_), .A2(pi1091), .B(new_n11950_), .ZN(new_n29241_));
  NOR2_X1    g26035(.A1(new_n26822_), .A2(pi1091), .ZN(new_n29242_));
  OAI21_X1   g26036(.A1(pi1153), .A2(new_n26431_), .B(new_n29242_), .ZN(new_n29243_));
  AOI21_X1   g26037(.A1(new_n8662_), .A2(new_n29113_), .B(pi1154), .ZN(new_n29244_));
  NAND4_X1   g26038(.A1(new_n29079_), .A2(new_n8247_), .A3(new_n29243_), .A4(new_n29244_), .ZN(new_n29245_));
  AOI21_X1   g26039(.A1(pi0211), .A2(new_n29241_), .B(new_n29245_), .ZN(new_n29246_));
  NOR2_X1    g26040(.A1(new_n26460_), .A2(new_n2918_), .ZN(new_n29247_));
  NOR2_X1    g26041(.A1(new_n29247_), .A2(new_n11893_), .ZN(new_n29248_));
  NOR2_X1    g26042(.A1(new_n29248_), .A2(pi1154), .ZN(new_n29249_));
  NOR2_X1    g26043(.A1(new_n29249_), .A2(new_n8077_), .ZN(new_n29250_));
  INV_X1     g26044(.I(new_n29250_), .ZN(new_n29251_));
  INV_X1     g26045(.I(new_n29241_), .ZN(new_n29252_));
  NAND3_X1   g26046(.A1(new_n29252_), .A2(new_n8077_), .A3(new_n29244_), .ZN(new_n29253_));
  AOI21_X1   g26047(.A1(new_n29253_), .A2(new_n29251_), .B(pi0219), .ZN(new_n29254_));
  NOR2_X1    g26048(.A1(new_n29246_), .A2(new_n29254_), .ZN(new_n29255_));
  INV_X1     g26049(.I(new_n29255_), .ZN(new_n29256_));
  NOR2_X1    g26050(.A1(new_n26411_), .A2(new_n2918_), .ZN(new_n29257_));
  NOR3_X1    g26051(.A1(new_n8094_), .A2(pi0200), .A3(pi0299), .ZN(new_n29258_));
  NOR2_X1    g26052(.A1(new_n29258_), .A2(new_n2918_), .ZN(new_n29259_));
  INV_X1     g26053(.I(new_n29259_), .ZN(new_n29260_));
  MUX2_X1    g26054(.I0(new_n29260_), .I1(new_n29072_), .S(pi1153), .Z(new_n29261_));
  INV_X1     g26055(.I(new_n29261_), .ZN(new_n29262_));
  NAND3_X1   g26056(.A1(new_n29073_), .A2(pi1091), .A3(new_n26431_), .ZN(new_n29263_));
  AOI21_X1   g26057(.A1(new_n29263_), .A2(pi1154), .B(new_n29086_), .ZN(new_n29264_));
  OAI21_X1   g26058(.A1(new_n29257_), .A2(new_n29262_), .B(new_n29264_), .ZN(new_n29265_));
  NOR2_X1    g26059(.A1(new_n8663_), .A2(new_n2918_), .ZN(new_n29266_));
  INV_X1     g26060(.I(new_n29266_), .ZN(new_n29267_));
  OAI21_X1   g26061(.A1(new_n26638_), .A2(new_n29267_), .B(new_n11950_), .ZN(new_n29268_));
  NOR2_X1    g26062(.A1(new_n2918_), .A2(pi1154), .ZN(new_n29269_));
  INV_X1     g26063(.I(new_n29269_), .ZN(new_n29270_));
  OAI21_X1   g26064(.A1(new_n26450_), .A2(new_n29270_), .B(new_n29261_), .ZN(new_n29271_));
  AOI22_X1   g26065(.A1(new_n29265_), .A2(new_n29268_), .B1(new_n8663_), .B2(new_n29271_), .ZN(new_n29272_));
  MUX2_X1    g26066(.I0(new_n29272_), .I1(new_n29256_), .S(new_n28262_), .Z(new_n29273_));
  MUX2_X1    g26067(.I0(new_n29226_), .I1(pi0254), .S(new_n2918_), .Z(new_n29274_));
  NAND2_X1   g26068(.A1(new_n29274_), .A2(po1038), .ZN(new_n29275_));
  AOI21_X1   g26069(.A1(new_n29275_), .A2(new_n26604_), .B(po1038), .ZN(new_n29276_));
  NAND2_X1   g26070(.A1(new_n29057_), .A2(pi1154), .ZN(new_n29277_));
  NAND2_X1   g26071(.A1(new_n29277_), .A2(new_n26672_), .ZN(new_n29278_));
  AOI21_X1   g26072(.A1(new_n29278_), .A2(new_n8247_), .B(new_n29237_), .ZN(new_n29279_));
  NOR3_X1    g26073(.A1(new_n29279_), .A2(pi0254), .A3(new_n2918_), .ZN(new_n29280_));
  NOR2_X1    g26074(.A1(new_n29077_), .A2(new_n11950_), .ZN(new_n29281_));
  AOI21_X1   g26075(.A1(pi0219), .A2(pi1091), .B(new_n29281_), .ZN(new_n29282_));
  INV_X1     g26076(.I(new_n26963_), .ZN(new_n29283_));
  NOR3_X1    g26077(.A1(new_n29283_), .A2(new_n2918_), .A3(new_n26389_), .ZN(new_n29284_));
  NOR4_X1    g26078(.A1(new_n29249_), .A2(new_n27264_), .A3(pi0211), .A4(new_n29103_), .ZN(new_n29285_));
  AOI21_X1   g26079(.A1(new_n27222_), .A2(new_n29284_), .B(new_n29285_), .ZN(new_n29286_));
  OAI22_X1   g26080(.A1(new_n29286_), .A2(pi0219), .B1(new_n29231_), .B2(new_n29282_), .ZN(new_n29287_));
  NAND2_X1   g26081(.A1(new_n29287_), .A2(pi0254), .ZN(new_n29288_));
  XOR2_X1    g26082(.A1(new_n29288_), .A2(new_n29280_), .Z(new_n29289_));
  NOR2_X1    g26083(.A1(new_n29289_), .A2(po1038), .ZN(new_n29290_));
  NAND3_X1   g26084(.A1(po1038), .A2(new_n8247_), .A3(new_n29076_), .ZN(new_n29291_));
  NAND2_X1   g26085(.A1(new_n29275_), .A2(new_n29291_), .ZN(new_n29292_));
  NAND2_X1   g26086(.A1(new_n29292_), .A2(pi1152), .ZN(new_n29293_));
  OAI21_X1   g26087(.A1(new_n29290_), .A2(new_n29293_), .B(new_n28287_), .ZN(new_n29294_));
  AOI21_X1   g26088(.A1(new_n29273_), .A2(new_n29276_), .B(new_n29294_), .ZN(new_n29295_));
  NOR2_X1    g26089(.A1(new_n28149_), .A2(new_n28232_), .ZN(new_n29296_));
  INV_X1     g26090(.I(new_n29296_), .ZN(new_n29297_));
  NOR2_X1    g26091(.A1(new_n28151_), .A2(new_n11893_), .ZN(new_n29308_));
  NOR2_X1    g26092(.A1(new_n28186_), .A2(pi1153), .ZN(new_n29310_));
  NOR2_X1    g26093(.A1(new_n29310_), .A2(new_n28134_), .ZN(new_n29311_));
  NOR2_X1    g26094(.A1(new_n28238_), .A2(pi1153), .ZN(new_n29314_));
  NAND3_X1   g26095(.A1(new_n29289_), .A2(new_n28261_), .A3(po1038), .ZN(new_n29322_));
  OAI21_X1   g26096(.A1(new_n28261_), .A2(new_n6845_), .B(new_n29292_), .ZN(new_n29323_));
  INV_X1     g26097(.I(new_n29166_), .ZN(new_n29324_));
  NOR3_X1    g26098(.A1(new_n26822_), .A2(new_n8247_), .A3(new_n2918_), .ZN(new_n29325_));
  NOR3_X1    g26099(.A1(new_n29325_), .A2(new_n29114_), .A3(pi0254), .ZN(new_n29326_));
  NAND3_X1   g26100(.A1(new_n29324_), .A2(new_n29179_), .A3(new_n29326_), .ZN(new_n29327_));
  NOR2_X1    g26101(.A1(new_n28108_), .A2(new_n8247_), .ZN(new_n29328_));
  OAI21_X1   g26102(.A1(pi0211), .A2(new_n28144_), .B(new_n29328_), .ZN(new_n29329_));
  INV_X1     g26103(.I(new_n29329_), .ZN(new_n29330_));
  NOR2_X1    g26104(.A1(new_n28116_), .A2(pi0219), .ZN(new_n29331_));
  NAND4_X1   g26105(.A1(new_n8663_), .A2(new_n28262_), .A3(pi1091), .A4(new_n11893_), .ZN(new_n29332_));
  NOR4_X1    g26106(.A1(new_n29330_), .A2(new_n29325_), .A3(new_n29331_), .A4(new_n29332_), .ZN(new_n29333_));
  INV_X1     g26107(.I(new_n29333_), .ZN(new_n29334_));
  NAND2_X1   g26108(.A1(new_n29327_), .A2(new_n29334_), .ZN(new_n29335_));
  NAND2_X1   g26109(.A1(new_n29335_), .A2(new_n28261_), .ZN(new_n29336_));
  NAND3_X1   g26110(.A1(new_n29336_), .A2(new_n29322_), .A3(new_n29323_), .ZN(new_n29337_));
  AOI21_X1   g26111(.A1(new_n28129_), .A2(pi1153), .B(new_n28174_), .ZN(new_n29338_));
  NOR2_X1    g26112(.A1(new_n28219_), .A2(pi1154), .ZN(new_n29339_));
  AOI21_X1   g26113(.A1(new_n28247_), .A2(new_n26822_), .B(new_n8247_), .ZN(new_n29340_));
  OAI21_X1   g26114(.A1(new_n29339_), .A2(new_n29338_), .B(new_n29340_), .ZN(new_n29341_));
  NOR2_X1    g26115(.A1(new_n28174_), .A2(pi1153), .ZN(new_n29342_));
  NAND2_X1   g26116(.A1(new_n28172_), .A2(pi1154), .ZN(new_n29343_));
  NAND3_X1   g26117(.A1(new_n29343_), .A2(new_n8247_), .A3(pi0254), .ZN(new_n29344_));
  NOR4_X1    g26118(.A1(new_n29131_), .A2(new_n28166_), .A3(new_n29342_), .A4(new_n29344_), .ZN(new_n29345_));
  NOR2_X1    g26119(.A1(new_n29314_), .A2(new_n26963_), .ZN(new_n29346_));
  AOI21_X1   g26120(.A1(new_n28152_), .A2(new_n29346_), .B(new_n8247_), .ZN(new_n29347_));
  OAI21_X1   g26121(.A1(new_n29311_), .A2(new_n28240_), .B(new_n11950_), .ZN(new_n29348_));
  NOR2_X1    g26122(.A1(new_n29314_), .A2(new_n26822_), .ZN(new_n29349_));
  AOI21_X1   g26123(.A1(new_n29296_), .A2(new_n29349_), .B(new_n29348_), .ZN(new_n29350_));
  INV_X1     g26124(.I(new_n29207_), .ZN(new_n29351_));
  NOR2_X1    g26125(.A1(new_n29157_), .A2(new_n28134_), .ZN(new_n29352_));
  NOR2_X1    g26126(.A1(new_n29151_), .A2(new_n28139_), .ZN(new_n29353_));
  AOI22_X1   g26127(.A1(pi1154), .A2(new_n29353_), .B1(new_n29352_), .B2(new_n29351_), .ZN(new_n29354_));
  AOI21_X1   g26128(.A1(new_n28143_), .A2(pi1154), .B(new_n28135_), .ZN(new_n29355_));
  OAI21_X1   g26129(.A1(new_n29355_), .A2(pi0211), .B(new_n8247_), .ZN(new_n29356_));
  NOR2_X1    g26130(.A1(new_n29354_), .A2(new_n29356_), .ZN(new_n29357_));
  AOI21_X1   g26131(.A1(new_n29347_), .A2(new_n29350_), .B(new_n29357_), .ZN(new_n29358_));
  INV_X1     g26132(.I(new_n29358_), .ZN(new_n29359_));
  AOI22_X1   g26133(.A1(new_n29359_), .A2(new_n28262_), .B1(new_n29341_), .B2(new_n29345_), .ZN(new_n29360_));
  OR3_X2     g26134(.A1(new_n29360_), .A2(pi0253), .A3(new_n29273_), .Z(new_n29361_));
  INV_X1     g26135(.I(new_n29273_), .ZN(new_n29362_));
  OAI21_X1   g26136(.A1(pi0253), .A2(new_n29362_), .B(new_n29360_), .ZN(new_n29363_));
  OAI21_X1   g26137(.A1(new_n29198_), .A2(new_n29327_), .B(pi0253), .ZN(new_n29364_));
  NOR2_X1    g26138(.A1(new_n29334_), .A2(new_n29181_), .ZN(new_n29365_));
  OAI21_X1   g26139(.A1(new_n28261_), .A2(new_n6845_), .B(new_n29275_), .ZN(new_n29366_));
  NAND2_X1   g26140(.A1(new_n29366_), .A2(new_n27881_), .ZN(new_n29367_));
  AOI21_X1   g26141(.A1(new_n29364_), .A2(new_n29365_), .B(new_n29367_), .ZN(new_n29368_));
  NAND3_X1   g26142(.A1(new_n29361_), .A2(new_n29363_), .A3(new_n29368_), .ZN(new_n29369_));
  AOI21_X1   g26143(.A1(new_n29369_), .A2(new_n28286_), .B(pi1152), .ZN(new_n29370_));
  AOI21_X1   g26144(.A1(new_n29370_), .A2(new_n29337_), .B(new_n29295_), .ZN(new_n29371_));
  OAI21_X1   g26145(.A1(new_n29371_), .A2(pi0230), .B(new_n29240_), .ZN(po0411));
  NAND2_X1   g26146(.A1(new_n29008_), .A2(pi0255), .ZN(new_n29373_));
  INV_X1     g26147(.I(pi1036), .ZN(new_n29374_));
  NAND2_X1   g26148(.A1(new_n29374_), .A2(pi0200), .ZN(new_n29375_));
  OAI21_X1   g26149(.A1(pi0200), .A2(pi1049), .B(new_n29375_), .ZN(new_n29376_));
  OAI21_X1   g26150(.A1(new_n29008_), .A2(new_n29376_), .B(new_n29373_), .ZN(po0412));
  NAND2_X1   g26151(.A1(new_n29008_), .A2(pi0256), .ZN(new_n29378_));
  INV_X1     g26152(.I(pi1070), .ZN(new_n29379_));
  NOR2_X1    g26153(.A1(pi0200), .A2(pi1048), .ZN(new_n29380_));
  AOI21_X1   g26154(.A1(pi0200), .A2(new_n29379_), .B(new_n29380_), .ZN(new_n29381_));
  NAND2_X1   g26155(.A1(new_n29381_), .A2(new_n29007_), .ZN(new_n29382_));
  NAND2_X1   g26156(.A1(new_n29382_), .A2(new_n29378_), .ZN(po0413));
  NAND2_X1   g26157(.A1(new_n29008_), .A2(pi0257), .ZN(new_n29384_));
  INV_X1     g26158(.I(pi1065), .ZN(new_n29385_));
  NOR2_X1    g26159(.A1(pi0200), .A2(pi1084), .ZN(new_n29386_));
  AOI21_X1   g26160(.A1(pi0200), .A2(new_n29385_), .B(new_n29386_), .ZN(new_n29387_));
  NAND2_X1   g26161(.A1(new_n29387_), .A2(new_n29007_), .ZN(new_n29388_));
  NAND2_X1   g26162(.A1(new_n29388_), .A2(new_n29384_), .ZN(po0414));
  NAND2_X1   g26163(.A1(new_n29008_), .A2(pi0258), .ZN(new_n29390_));
  INV_X1     g26164(.I(pi1062), .ZN(new_n29391_));
  NOR2_X1    g26165(.A1(pi0200), .A2(pi1072), .ZN(new_n29392_));
  AOI21_X1   g26166(.A1(pi0200), .A2(new_n29391_), .B(new_n29392_), .ZN(new_n29393_));
  NAND2_X1   g26167(.A1(new_n29393_), .A2(new_n29007_), .ZN(new_n29394_));
  NAND2_X1   g26168(.A1(new_n29394_), .A2(new_n29390_), .ZN(po0415));
  NAND2_X1   g26169(.A1(new_n29008_), .A2(pi0259), .ZN(new_n29396_));
  INV_X1     g26170(.I(pi1069), .ZN(new_n29397_));
  NOR2_X1    g26171(.A1(pi0200), .A2(pi1059), .ZN(new_n29398_));
  AOI21_X1   g26172(.A1(pi0200), .A2(new_n29397_), .B(new_n29398_), .ZN(new_n29399_));
  NAND2_X1   g26173(.A1(new_n29399_), .A2(new_n29007_), .ZN(new_n29400_));
  NAND2_X1   g26174(.A1(new_n29400_), .A2(new_n29396_), .ZN(po0416));
  NAND2_X1   g26175(.A1(new_n29008_), .A2(pi0260), .ZN(new_n29402_));
  OAI21_X1   g26176(.A1(pi0200), .A2(pi1044), .B(pi1067), .ZN(new_n29403_));
  INV_X1     g26177(.I(pi1067), .ZN(new_n29404_));
  NAND3_X1   g26178(.A1(new_n8098_), .A2(new_n29404_), .A3(pi1044), .ZN(new_n29405_));
  NAND4_X1   g26179(.A1(new_n29405_), .A2(new_n8094_), .A3(new_n29007_), .A4(new_n29403_), .ZN(new_n29406_));
  NAND2_X1   g26180(.A1(new_n29406_), .A2(new_n29402_), .ZN(po0417));
  NAND2_X1   g26181(.A1(new_n29008_), .A2(pi0261), .ZN(new_n29408_));
  OAI21_X1   g26182(.A1(pi0200), .A2(pi1037), .B(pi1040), .ZN(new_n29409_));
  INV_X1     g26183(.I(pi1040), .ZN(new_n29410_));
  NAND3_X1   g26184(.A1(new_n8098_), .A2(new_n29410_), .A3(pi1037), .ZN(new_n29411_));
  NAND4_X1   g26185(.A1(new_n29411_), .A2(new_n8094_), .A3(new_n29007_), .A4(new_n29409_), .ZN(new_n29412_));
  NAND2_X1   g26186(.A1(new_n29412_), .A2(new_n29408_), .ZN(po0418));
  NOR3_X1    g26187(.A1(new_n3712_), .A2(new_n3700_), .A3(pi1093), .ZN(new_n29414_));
  AOI21_X1   g26188(.A1(new_n3712_), .A2(new_n2924_), .B(pi1142), .ZN(new_n29415_));
  NOR3_X1    g26189(.A1(new_n29415_), .A2(new_n29414_), .A3(pi0228), .ZN(new_n29416_));
  NOR2_X1    g26190(.A1(new_n2924_), .A2(pi0228), .ZN(new_n29417_));
  NOR2_X1    g26191(.A1(new_n2523_), .A2(pi0123), .ZN(new_n29418_));
  NOR2_X1    g26192(.A1(new_n29417_), .A2(new_n29418_), .ZN(new_n29419_));
  INV_X1     g26193(.I(new_n29419_), .ZN(new_n29420_));
  NOR4_X1    g26194(.A1(po1038), .A2(new_n27316_), .A3(new_n29416_), .A4(new_n29420_), .ZN(new_n29421_));
  NOR2_X1    g26195(.A1(new_n27316_), .A2(new_n2587_), .ZN(new_n29422_));
  AOI21_X1   g26196(.A1(new_n3712_), .A2(new_n29419_), .B(new_n29422_), .ZN(new_n29423_));
  NOR4_X1    g26197(.A1(new_n29423_), .A2(new_n8094_), .A3(new_n26328_), .A4(new_n29419_), .ZN(new_n29424_));
  NOR2_X1    g26198(.A1(pi0207), .A2(pi0262), .ZN(new_n29425_));
  AOI21_X1   g26199(.A1(new_n29419_), .A2(new_n29425_), .B(pi0208), .ZN(new_n29426_));
  OAI22_X1   g26200(.A1(new_n29424_), .A2(new_n29416_), .B1(new_n29422_), .B2(new_n29426_), .ZN(new_n29427_));
  INV_X1     g26201(.I(new_n29416_), .ZN(new_n29428_));
  INV_X1     g26202(.I(new_n29423_), .ZN(new_n29429_));
  NOR2_X1    g26203(.A1(new_n29420_), .A2(new_n27218_), .ZN(new_n29430_));
  NOR4_X1    g26204(.A1(new_n29429_), .A2(pi0208), .A3(pi0299), .A4(new_n29430_), .ZN(new_n29431_));
  AOI21_X1   g26205(.A1(new_n29431_), .A2(new_n29428_), .B(po1038), .ZN(new_n29432_));
  AOI21_X1   g26206(.A1(new_n29432_), .A2(new_n29427_), .B(new_n29421_), .ZN(po0419));
  INV_X1     g26207(.I(pi0263), .ZN(new_n29434_));
  NOR2_X1    g26208(.A1(new_n28137_), .A2(new_n28193_), .ZN(new_n29435_));
  INV_X1     g26209(.I(new_n29435_), .ZN(new_n29436_));
  AOI21_X1   g26210(.A1(new_n11912_), .A2(new_n28189_), .B(new_n29436_), .ZN(new_n29437_));
  NOR3_X1    g26211(.A1(new_n29435_), .A2(pi1155), .A3(new_n28189_), .ZN(new_n29438_));
  NOR3_X1    g26212(.A1(new_n29437_), .A2(new_n29438_), .A3(pi1154), .ZN(new_n29439_));
  NOR2_X1    g26213(.A1(new_n28157_), .A2(new_n11912_), .ZN(new_n29440_));
  INV_X1     g26214(.I(new_n29440_), .ZN(new_n29441_));
  INV_X1     g26215(.I(new_n28202_), .ZN(new_n29442_));
  AOI21_X1   g26216(.A1(new_n29442_), .A2(new_n11912_), .B(pi1154), .ZN(new_n29443_));
  AOI21_X1   g26217(.A1(new_n29441_), .A2(new_n29443_), .B(new_n12026_), .ZN(new_n29444_));
  OAI21_X1   g26218(.A1(new_n29353_), .A2(new_n29439_), .B(new_n29444_), .ZN(new_n29445_));
  NAND2_X1   g26219(.A1(new_n29441_), .A2(new_n29443_), .ZN(new_n29446_));
  NAND3_X1   g26220(.A1(new_n29446_), .A2(new_n12026_), .A3(new_n29343_), .ZN(new_n29447_));
  NAND2_X1   g26221(.A1(new_n29447_), .A2(new_n29439_), .ZN(new_n29448_));
  AOI21_X1   g26222(.A1(new_n8077_), .A2(new_n29445_), .B(new_n29448_), .ZN(new_n29449_));
  OR3_X2     g26223(.A1(new_n29352_), .A2(pi1155), .A3(new_n28189_), .Z(new_n29450_));
  NAND2_X1   g26224(.A1(new_n29450_), .A2(new_n11950_), .ZN(new_n29451_));
  OAI21_X1   g26225(.A1(pi1155), .A2(new_n28175_), .B(new_n29352_), .ZN(new_n29452_));
  OAI21_X1   g26226(.A1(new_n29447_), .A2(pi1156), .B(new_n29452_), .ZN(new_n29453_));
  AOI21_X1   g26227(.A1(new_n28170_), .A2(new_n11912_), .B(pi1154), .ZN(new_n29454_));
  AOI22_X1   g26228(.A1(new_n29441_), .A2(new_n29454_), .B1(pi1156), .B2(new_n29353_), .ZN(new_n29455_));
  OAI21_X1   g26229(.A1(new_n29453_), .A2(new_n29451_), .B(new_n29455_), .ZN(new_n29456_));
  NAND2_X1   g26230(.A1(new_n29456_), .A2(new_n8663_), .ZN(new_n29457_));
  INV_X1     g26231(.I(new_n26366_), .ZN(new_n29458_));
  AOI21_X1   g26232(.A1(pi1155), .A2(new_n28240_), .B(new_n28142_), .ZN(new_n29459_));
  NAND3_X1   g26233(.A1(new_n28151_), .A2(pi1154), .A3(new_n28143_), .ZN(new_n29460_));
  INV_X1     g26234(.I(new_n28143_), .ZN(new_n29461_));
  OAI21_X1   g26235(.A1(pi1154), .A2(new_n29461_), .B(new_n28150_), .ZN(new_n29462_));
  AOI21_X1   g26236(.A1(new_n29460_), .A2(new_n29462_), .B(new_n29459_), .ZN(new_n29463_));
  OAI21_X1   g26237(.A1(new_n29463_), .A2(new_n29458_), .B(pi0219), .ZN(new_n29464_));
  INV_X1     g26238(.I(new_n28193_), .ZN(new_n29465_));
  NAND2_X1   g26239(.A1(new_n29463_), .A2(new_n29465_), .ZN(new_n29466_));
  NAND2_X1   g26240(.A1(new_n29466_), .A2(new_n12026_), .ZN(new_n29467_));
  MUX2_X1    g26241(.I0(new_n29296_), .I1(new_n29129_), .S(new_n11912_), .Z(new_n29468_));
  NOR2_X1    g26242(.A1(new_n26819_), .A2(pi1154), .ZN(new_n29469_));
  NAND4_X1   g26243(.A1(new_n29467_), .A2(new_n29464_), .A3(new_n29468_), .A4(new_n29469_), .ZN(new_n29470_));
  OAI21_X1   g26244(.A1(new_n29457_), .A2(new_n29449_), .B(new_n29470_), .ZN(new_n29471_));
  NOR2_X1    g26245(.A1(new_n28232_), .A2(new_n11950_), .ZN(new_n29472_));
  OAI21_X1   g26246(.A1(new_n28130_), .A2(new_n11912_), .B(new_n29472_), .ZN(new_n29473_));
  INV_X1     g26247(.I(new_n28224_), .ZN(new_n29474_));
  INV_X1     g26248(.I(new_n29202_), .ZN(new_n29475_));
  NOR3_X1    g26249(.A1(new_n29474_), .A2(pi1155), .A3(new_n29475_), .ZN(new_n29476_));
  AOI21_X1   g26250(.A1(new_n11912_), .A2(new_n29475_), .B(new_n28224_), .ZN(new_n29477_));
  NOR3_X1    g26251(.A1(new_n29476_), .A2(pi1154), .A3(new_n29477_), .ZN(new_n29478_));
  AOI21_X1   g26252(.A1(new_n29478_), .A2(new_n29473_), .B(pi1156), .ZN(new_n29479_));
  NOR2_X1    g26253(.A1(pi1154), .A2(pi1155), .ZN(new_n29480_));
  NAND3_X1   g26254(.A1(new_n28224_), .A2(new_n28174_), .A3(new_n29480_), .ZN(new_n29481_));
  OAI21_X1   g26255(.A1(new_n28134_), .A2(new_n29473_), .B(new_n29481_), .ZN(new_n29482_));
  NAND2_X1   g26256(.A1(new_n29482_), .A2(new_n26366_), .ZN(new_n29483_));
  OAI21_X1   g26257(.A1(new_n28241_), .A2(pi1154), .B(new_n28251_), .ZN(new_n29484_));
  AOI21_X1   g26258(.A1(new_n28129_), .A2(pi1155), .B(new_n26820_), .ZN(new_n29485_));
  AOI21_X1   g26259(.A1(new_n29485_), .A2(new_n29484_), .B(new_n8247_), .ZN(new_n29486_));
  NAND2_X1   g26260(.A1(new_n29483_), .A2(new_n29486_), .ZN(new_n29487_));
  NOR2_X1    g26261(.A1(new_n29487_), .A2(new_n29479_), .ZN(new_n29488_));
  AOI21_X1   g26262(.A1(new_n29151_), .A2(pi1155), .B(new_n11950_), .ZN(new_n29489_));
  INV_X1     g26263(.I(new_n29489_), .ZN(new_n29490_));
  NOR3_X1    g26264(.A1(new_n29490_), .A2(new_n28135_), .A3(new_n28143_), .ZN(new_n29491_));
  NOR4_X1    g26265(.A1(new_n29491_), .A2(new_n29476_), .A3(pi1154), .A4(new_n29477_), .ZN(new_n29492_));
  NAND2_X1   g26266(.A1(new_n29491_), .A2(new_n28132_), .ZN(new_n29493_));
  NAND2_X1   g26267(.A1(new_n29146_), .A2(new_n28155_), .ZN(new_n29494_));
  AOI21_X1   g26268(.A1(new_n28173_), .A2(new_n11912_), .B(pi1154), .ZN(new_n29495_));
  AOI21_X1   g26269(.A1(new_n29494_), .A2(new_n29495_), .B(new_n12026_), .ZN(new_n29496_));
  INV_X1     g26270(.I(new_n29496_), .ZN(new_n29497_));
  AOI21_X1   g26271(.A1(new_n29493_), .A2(new_n29481_), .B(new_n29497_), .ZN(new_n29498_));
  NAND2_X1   g26272(.A1(new_n28166_), .A2(new_n11912_), .ZN(new_n29499_));
  NAND3_X1   g26273(.A1(new_n29202_), .A2(new_n29157_), .A3(new_n11912_), .ZN(new_n29500_));
  NAND3_X1   g26274(.A1(new_n29499_), .A2(new_n26444_), .A3(new_n29500_), .ZN(new_n29501_));
  OAI21_X1   g26275(.A1(new_n29498_), .A2(pi0211), .B(new_n29501_), .ZN(new_n29502_));
  OAI21_X1   g26276(.A1(new_n28180_), .A2(new_n29490_), .B(new_n29496_), .ZN(new_n29503_));
  AND4_X2    g26277(.A1(new_n8077_), .A2(new_n29501_), .A3(new_n29123_), .A4(new_n29489_), .Z(new_n29504_));
  NAND2_X1   g26278(.A1(new_n8247_), .A2(new_n29434_), .ZN(new_n29505_));
  AOI21_X1   g26279(.A1(new_n29504_), .A2(new_n29503_), .B(new_n29505_), .ZN(new_n29506_));
  OAI21_X1   g26280(.A1(new_n29502_), .A2(new_n29492_), .B(new_n29506_), .ZN(new_n29507_));
  OAI21_X1   g26281(.A1(new_n29507_), .A2(new_n29488_), .B(new_n28265_), .ZN(new_n29508_));
  NAND3_X1   g26282(.A1(new_n29471_), .A2(new_n29434_), .A3(new_n29508_), .ZN(new_n29509_));
  INV_X1     g26283(.I(new_n27161_), .ZN(new_n29510_));
  NAND2_X1   g26284(.A1(new_n26441_), .A2(new_n29510_), .ZN(new_n29511_));
  NOR2_X1    g26285(.A1(new_n29511_), .A2(new_n29077_), .ZN(new_n29512_));
  OAI21_X1   g26286(.A1(new_n26606_), .A2(new_n11950_), .B(pi1091), .ZN(new_n29513_));
  NOR2_X1    g26287(.A1(new_n29513_), .A2(new_n26522_), .ZN(new_n29514_));
  NAND2_X1   g26288(.A1(new_n29514_), .A2(pi0211), .ZN(new_n29515_));
  OAI21_X1   g26289(.A1(new_n29515_), .A2(new_n29512_), .B(new_n12026_), .ZN(new_n29516_));
  AOI21_X1   g26290(.A1(new_n29512_), .A2(new_n29515_), .B(new_n29516_), .ZN(new_n29517_));
  NOR2_X1    g26291(.A1(pi0199), .A2(pi1154), .ZN(new_n29518_));
  NOR2_X1    g26292(.A1(new_n8077_), .A2(new_n2918_), .ZN(new_n29519_));
  NOR4_X1    g26293(.A1(new_n26522_), .A2(new_n26390_), .A3(new_n29518_), .A4(new_n29519_), .ZN(new_n29520_));
  NOR2_X1    g26294(.A1(new_n26757_), .A2(new_n11912_), .ZN(new_n29521_));
  INV_X1     g26295(.I(new_n29521_), .ZN(new_n29522_));
  AOI22_X1   g26296(.A1(new_n29522_), .A2(new_n29080_), .B1(new_n11950_), .B2(new_n29257_), .ZN(new_n29523_));
  AOI21_X1   g26297(.A1(new_n29523_), .A2(new_n8077_), .B(new_n29520_), .ZN(new_n29524_));
  OAI21_X1   g26298(.A1(new_n29524_), .A2(new_n12026_), .B(new_n8247_), .ZN(new_n29525_));
  NAND4_X1   g26299(.A1(new_n29523_), .A2(pi0299), .A3(pi1091), .A4(new_n29458_), .ZN(new_n29526_));
  OAI21_X1   g26300(.A1(new_n26435_), .A2(new_n26432_), .B(new_n11950_), .ZN(new_n29527_));
  INV_X1     g26301(.I(new_n29513_), .ZN(new_n29528_));
  NAND3_X1   g26302(.A1(new_n29528_), .A2(new_n8247_), .A3(new_n26828_), .ZN(new_n29529_));
  NOR3_X1    g26303(.A1(new_n26382_), .A2(pi1154), .A3(new_n26379_), .ZN(new_n29530_));
  NOR3_X1    g26304(.A1(new_n29530_), .A2(new_n2918_), .A3(new_n26820_), .ZN(new_n29531_));
  NAND4_X1   g26305(.A1(new_n29526_), .A2(new_n29527_), .A3(new_n29529_), .A4(new_n29531_), .ZN(new_n29532_));
  OAI21_X1   g26306(.A1(new_n29517_), .A2(new_n29525_), .B(new_n29532_), .ZN(new_n29533_));
  NAND3_X1   g26307(.A1(new_n29527_), .A2(new_n11912_), .A3(new_n8269_), .ZN(new_n29534_));
  NAND4_X1   g26308(.A1(new_n29534_), .A2(new_n26390_), .A3(new_n26444_), .A4(new_n26545_), .ZN(new_n29535_));
  NAND4_X1   g26309(.A1(new_n29535_), .A2(new_n8077_), .A3(new_n12026_), .A4(new_n29514_), .ZN(new_n29536_));
  NAND2_X1   g26310(.A1(new_n12026_), .A2(pi1154), .ZN(new_n29537_));
  OAI21_X1   g26311(.A1(new_n26385_), .A2(new_n29537_), .B(new_n2587_), .ZN(new_n29538_));
  NAND2_X1   g26312(.A1(new_n8268_), .A2(new_n11950_), .ZN(new_n29539_));
  OAI21_X1   g26313(.A1(new_n29539_), .A2(new_n26385_), .B(new_n27622_), .ZN(new_n29540_));
  OAI21_X1   g26314(.A1(new_n29540_), .A2(new_n29538_), .B(pi1156), .ZN(new_n29541_));
  AOI21_X1   g26315(.A1(new_n29511_), .A2(new_n29538_), .B(new_n8247_), .ZN(new_n29542_));
  NAND2_X1   g26316(.A1(pi0263), .A2(pi1091), .ZN(new_n29543_));
  AOI21_X1   g26317(.A1(new_n29542_), .A2(new_n29541_), .B(new_n29543_), .ZN(new_n29544_));
  NOR2_X1    g26318(.A1(new_n26412_), .A2(new_n27094_), .ZN(new_n29545_));
  NOR3_X1    g26319(.A1(new_n29545_), .A2(new_n8098_), .A3(pi1155), .ZN(new_n29546_));
  NAND2_X1   g26320(.A1(new_n29510_), .A2(new_n8077_), .ZN(new_n29547_));
  OAI21_X1   g26321(.A1(new_n29546_), .A2(new_n29547_), .B(new_n8247_), .ZN(new_n29548_));
  NOR2_X1    g26322(.A1(new_n29548_), .A2(new_n29544_), .ZN(new_n29549_));
  AOI22_X1   g26323(.A1(new_n29533_), .A2(new_n29434_), .B1(new_n29536_), .B2(new_n29549_), .ZN(new_n29550_));
  NAND2_X1   g26324(.A1(new_n29550_), .A2(new_n28266_), .ZN(new_n29551_));
  AOI21_X1   g26325(.A1(new_n29509_), .A2(new_n6845_), .B(new_n29551_), .ZN(new_n29552_));
  OAI22_X1   g26326(.A1(new_n28140_), .A2(new_n8077_), .B1(new_n26817_), .B2(new_n29281_), .ZN(new_n29553_));
  NAND4_X1   g26327(.A1(new_n29324_), .A2(new_n29434_), .A3(new_n29167_), .A4(new_n29553_), .ZN(new_n29554_));
  NAND2_X1   g26328(.A1(new_n29329_), .A2(new_n29434_), .ZN(new_n29555_));
  NAND3_X1   g26329(.A1(new_n28108_), .A2(pi0211), .A3(pi1155), .ZN(new_n29556_));
  NAND3_X1   g26330(.A1(new_n29555_), .A2(new_n29167_), .A3(new_n29556_), .ZN(new_n29557_));
  NAND3_X1   g26331(.A1(new_n26820_), .A2(pi0219), .A3(pi1091), .ZN(new_n29558_));
  NAND2_X1   g26332(.A1(new_n28265_), .A2(new_n29558_), .ZN(new_n29559_));
  AOI21_X1   g26333(.A1(new_n29554_), .A2(new_n29557_), .B(new_n29559_), .ZN(new_n29560_));
  NOR2_X1    g26334(.A1(new_n26820_), .A2(new_n8247_), .ZN(new_n29561_));
  OAI21_X1   g26335(.A1(pi0211), .A2(new_n11950_), .B(new_n26818_), .ZN(new_n29562_));
  AOI21_X1   g26336(.A1(new_n29562_), .A2(new_n8247_), .B(new_n29561_), .ZN(new_n29563_));
  NOR2_X1    g26337(.A1(new_n29563_), .A2(new_n2918_), .ZN(new_n29564_));
  AOI21_X1   g26338(.A1(new_n29434_), .A2(new_n2918_), .B(new_n29564_), .ZN(new_n29565_));
  INV_X1     g26339(.I(new_n29565_), .ZN(new_n29566_));
  NAND3_X1   g26340(.A1(new_n29566_), .A2(new_n6845_), .A3(new_n28266_), .ZN(new_n29567_));
  OAI21_X1   g26341(.A1(new_n29560_), .A2(new_n29567_), .B(new_n28286_), .ZN(new_n29568_));
  NOR3_X1    g26342(.A1(new_n29550_), .A2(po1038), .A3(new_n29565_), .ZN(new_n29569_));
  AOI21_X1   g26343(.A1(new_n29550_), .A2(new_n6845_), .B(new_n29566_), .ZN(new_n29570_));
  NOR3_X1    g26344(.A1(new_n29569_), .A2(new_n29570_), .A3(new_n28292_), .ZN(new_n29571_));
  OAI21_X1   g26345(.A1(new_n29552_), .A2(new_n29568_), .B(new_n29571_), .ZN(po0420));
  OAI21_X1   g26346(.A1(pi0211), .A2(pi1141), .B(pi1142), .ZN(new_n29573_));
  INV_X1     g26347(.I(new_n29573_), .ZN(new_n29574_));
  NOR3_X1    g26348(.A1(new_n3831_), .A2(pi0211), .A3(pi1142), .ZN(new_n29575_));
  NOR4_X1    g26349(.A1(new_n28305_), .A2(pi0219), .A3(new_n29574_), .A4(new_n29575_), .ZN(new_n29576_));
  OAI21_X1   g26350(.A1(pi0199), .A2(pi1141), .B(pi1143), .ZN(new_n29577_));
  NAND3_X1   g26351(.A1(new_n8094_), .A2(new_n3548_), .A3(pi1141), .ZN(new_n29578_));
  NAND4_X1   g26352(.A1(new_n26330_), .A2(new_n8098_), .A3(new_n29577_), .A4(new_n29578_), .ZN(new_n29579_));
  MUX2_X1    g26353(.I0(new_n29576_), .I1(new_n29579_), .S(new_n11749_), .Z(new_n29580_));
  NAND2_X1   g26354(.A1(new_n29580_), .A2(pi0230), .ZN(new_n29581_));
  NAND3_X1   g26355(.A1(new_n28111_), .A2(pi0264), .A3(pi0796), .ZN(new_n29582_));
  INV_X1     g26356(.I(pi0796), .ZN(new_n29583_));
  INV_X1     g26357(.I(new_n28111_), .ZN(new_n29584_));
  OAI21_X1   g26358(.A1(new_n29584_), .A2(pi0264), .B(new_n29583_), .ZN(new_n29585_));
  NAND3_X1   g26359(.A1(new_n29585_), .A2(new_n2918_), .A3(new_n29582_), .ZN(new_n29586_));
  AOI21_X1   g26360(.A1(pi1091), .A2(pi1141), .B(new_n29586_), .ZN(new_n29587_));
  AOI21_X1   g26361(.A1(pi1091), .A2(pi1142), .B(new_n29586_), .ZN(new_n29588_));
  XNOR2_X1   g26362(.A1(new_n29587_), .A2(new_n29588_), .ZN(new_n29589_));
  NOR2_X1    g26363(.A1(new_n29589_), .A2(new_n8077_), .ZN(new_n29590_));
  XNOR2_X1   g26364(.A1(new_n29590_), .A2(new_n29587_), .ZN(new_n29591_));
  OAI21_X1   g26365(.A1(new_n29591_), .A2(pi0219), .B(new_n27783_), .ZN(new_n29592_));
  INV_X1     g26366(.I(pi0264), .ZN(new_n29593_));
  NOR3_X1    g26367(.A1(new_n28101_), .A2(new_n29593_), .A3(new_n29583_), .ZN(new_n29594_));
  AOI21_X1   g26368(.A1(new_n28102_), .A2(new_n29593_), .B(pi0796), .ZN(new_n29595_));
  AOI21_X1   g26369(.A1(pi0219), .A2(new_n29077_), .B(new_n28305_), .ZN(new_n29596_));
  NOR4_X1    g26370(.A1(new_n29596_), .A2(new_n29595_), .A3(pi1091), .A4(new_n29594_), .ZN(new_n29597_));
  MUX2_X1    g26371(.I0(new_n29588_), .I1(new_n29587_), .S(new_n8098_), .Z(new_n29598_));
  NAND2_X1   g26372(.A1(new_n29598_), .A2(new_n8094_), .ZN(new_n29599_));
  NOR3_X1    g26373(.A1(new_n29595_), .A2(pi1091), .A3(new_n29594_), .ZN(new_n29600_));
  NOR2_X1    g26374(.A1(new_n2918_), .A2(pi0200), .ZN(new_n29601_));
  INV_X1     g26375(.I(new_n29601_), .ZN(new_n29602_));
  NOR2_X1    g26376(.A1(new_n26321_), .A2(new_n29602_), .ZN(new_n29603_));
  NOR3_X1    g26377(.A1(new_n11749_), .A2(new_n29600_), .A3(new_n29603_), .ZN(new_n29604_));
  AOI22_X1   g26378(.A1(new_n29592_), .A2(new_n29597_), .B1(new_n29599_), .B2(new_n29604_), .ZN(new_n29605_));
  OAI21_X1   g26379(.A1(new_n29605_), .A2(pi0230), .B(new_n29581_), .ZN(po0421));
  INV_X1     g26380(.I(pi0265), .ZN(new_n29607_));
  INV_X1     g26381(.I(pi0819), .ZN(new_n29608_));
  NOR3_X1    g26382(.A1(new_n29584_), .A2(new_n29607_), .A3(new_n29608_), .ZN(new_n29609_));
  AOI21_X1   g26383(.A1(new_n28111_), .A2(new_n29607_), .B(pi0819), .ZN(new_n29610_));
  NOR3_X1    g26384(.A1(new_n29609_), .A2(pi1091), .A3(new_n29610_), .ZN(new_n29611_));
  OAI21_X1   g26385(.A1(new_n2918_), .A2(new_n3700_), .B(new_n29611_), .ZN(new_n29612_));
  NAND2_X1   g26386(.A1(pi1091), .A2(pi1143), .ZN(new_n29613_));
  NAND2_X1   g26387(.A1(new_n29611_), .A2(new_n29613_), .ZN(new_n29614_));
  MUX2_X1    g26388(.I0(new_n29614_), .I1(new_n29612_), .S(new_n8077_), .Z(new_n29615_));
  NOR2_X1    g26389(.A1(new_n29615_), .A2(pi0219), .ZN(new_n29616_));
  NOR3_X1    g26390(.A1(new_n28101_), .A2(new_n29607_), .A3(new_n29608_), .ZN(new_n29617_));
  AOI21_X1   g26391(.A1(new_n28102_), .A2(new_n29607_), .B(pi0819), .ZN(new_n29618_));
  NOR3_X1    g26392(.A1(new_n29618_), .A2(pi1091), .A3(new_n29617_), .ZN(new_n29619_));
  OAI21_X1   g26393(.A1(new_n8247_), .A2(new_n29076_), .B(new_n28064_), .ZN(new_n29620_));
  AOI21_X1   g26394(.A1(new_n29619_), .A2(new_n29620_), .B(new_n11749_), .ZN(new_n29621_));
  MUX2_X1    g26395(.I0(new_n29614_), .I1(new_n29612_), .S(new_n8098_), .Z(new_n29622_));
  NOR2_X1    g26396(.A1(new_n26325_), .A2(new_n29602_), .ZN(new_n29623_));
  AOI21_X1   g26397(.A1(new_n29619_), .A2(new_n29623_), .B(new_n27783_), .ZN(new_n29624_));
  OAI21_X1   g26398(.A1(new_n29622_), .A2(pi0199), .B(new_n29624_), .ZN(new_n29625_));
  OAI21_X1   g26399(.A1(new_n29616_), .A2(new_n29621_), .B(new_n29625_), .ZN(new_n29626_));
  OAI21_X1   g26400(.A1(pi0211), .A2(pi1142), .B(pi1143), .ZN(new_n29627_));
  NAND3_X1   g26401(.A1(new_n8077_), .A2(new_n3548_), .A3(pi1142), .ZN(new_n29628_));
  NAND4_X1   g26402(.A1(new_n29628_), .A2(new_n28064_), .A3(new_n8247_), .A4(new_n29627_), .ZN(new_n29629_));
  NAND2_X1   g26403(.A1(new_n27783_), .A2(new_n29629_), .ZN(new_n29630_));
  AOI22_X1   g26404(.A1(pi0200), .A2(new_n26321_), .B1(new_n26330_), .B2(new_n28037_), .ZN(new_n29631_));
  OAI21_X1   g26405(.A1(new_n27783_), .A2(new_n29631_), .B(new_n29630_), .ZN(new_n29632_));
  MUX2_X1    g26406(.I0(new_n29632_), .I1(new_n29626_), .S(new_n26307_), .Z(po0422));
  INV_X1     g26407(.I(pi1134), .ZN(new_n29634_));
  NOR2_X1    g26408(.A1(new_n29584_), .A2(pi0266), .ZN(new_n29635_));
  NOR2_X1    g26409(.A1(new_n28111_), .A2(pi0948), .ZN(new_n29636_));
  NOR3_X1    g26410(.A1(new_n29635_), .A2(pi1091), .A3(new_n29636_), .ZN(new_n29637_));
  INV_X1     g26411(.I(new_n29637_), .ZN(new_n29638_));
  OAI21_X1   g26412(.A1(new_n28102_), .A2(pi0948), .B(new_n2918_), .ZN(new_n29639_));
  AOI21_X1   g26413(.A1(new_n4559_), .A2(new_n28102_), .B(new_n29639_), .ZN(new_n29640_));
  NAND2_X1   g26414(.A1(pi1091), .A2(pi1135), .ZN(new_n29641_));
  NAND4_X1   g26415(.A1(new_n29638_), .A2(new_n8160_), .A3(new_n29640_), .A4(new_n29641_), .ZN(new_n29642_));
  INV_X1     g26416(.I(new_n29642_), .ZN(new_n29643_));
  INV_X1     g26417(.I(new_n29640_), .ZN(new_n29644_));
  OAI21_X1   g26418(.A1(new_n2918_), .A2(new_n4543_), .B(new_n29644_), .ZN(new_n29645_));
  MUX2_X1    g26419(.I0(new_n29645_), .I1(new_n29637_), .S(new_n8094_), .Z(new_n29646_));
  AOI21_X1   g26420(.A1(new_n29646_), .A2(new_n8098_), .B(new_n29643_), .ZN(new_n29647_));
  NOR2_X1    g26421(.A1(new_n29637_), .A2(pi0219), .ZN(new_n29648_));
  INV_X1     g26422(.I(new_n29648_), .ZN(new_n29649_));
  NAND3_X1   g26423(.A1(new_n29076_), .A2(new_n8247_), .A3(pi1136), .ZN(new_n29650_));
  AOI21_X1   g26424(.A1(new_n29644_), .A2(new_n29650_), .B(new_n11749_), .ZN(new_n29651_));
  NOR4_X1    g26425(.A1(new_n29651_), .A2(new_n8077_), .A3(new_n2918_), .A4(new_n4696_), .ZN(new_n29652_));
  AOI21_X1   g26426(.A1(new_n29652_), .A2(new_n29649_), .B(pi0230), .ZN(new_n29653_));
  OAI21_X1   g26427(.A1(new_n29647_), .A2(new_n27783_), .B(new_n29653_), .ZN(new_n29654_));
  AOI21_X1   g26428(.A1(new_n8094_), .A2(pi1091), .B(new_n29646_), .ZN(new_n29655_));
  OAI21_X1   g26429(.A1(new_n29655_), .A2(pi0200), .B(new_n29642_), .ZN(new_n29656_));
  INV_X1     g26430(.I(new_n29651_), .ZN(new_n29657_));
  NOR4_X1    g26431(.A1(new_n29648_), .A2(new_n8077_), .A3(pi1091), .A4(pi1135), .ZN(new_n29658_));
  NOR2_X1    g26432(.A1(new_n8077_), .A2(pi1136), .ZN(new_n29659_));
  AOI21_X1   g26433(.A1(new_n4696_), .A2(pi0211), .B(pi0219), .ZN(new_n29660_));
  OAI21_X1   g26434(.A1(new_n29659_), .A2(new_n29660_), .B(new_n27783_), .ZN(new_n29661_));
  NOR2_X1    g26435(.A1(new_n8094_), .A2(pi1136), .ZN(new_n29662_));
  OAI22_X1   g26436(.A1(new_n29662_), .A2(pi0200), .B1(new_n8094_), .B2(pi1135), .ZN(new_n29663_));
  NAND2_X1   g26437(.A1(new_n11749_), .A2(new_n29663_), .ZN(new_n29664_));
  AOI21_X1   g26438(.A1(new_n29661_), .A2(new_n29664_), .B(pi0230), .ZN(new_n29665_));
  OAI21_X1   g26439(.A1(new_n29657_), .A2(new_n29658_), .B(new_n29665_), .ZN(new_n29666_));
  AOI21_X1   g26440(.A1(new_n29656_), .A2(new_n11749_), .B(new_n29666_), .ZN(new_n29667_));
  MUX2_X1    g26441(.I0(new_n29667_), .I1(new_n29654_), .S(new_n29634_), .Z(po0423));
  AOI21_X1   g26442(.A1(new_n29157_), .A2(pi1153), .B(pi1155), .ZN(new_n29669_));
  OAI21_X1   g26443(.A1(pi1153), .A2(new_n29435_), .B(new_n29669_), .ZN(new_n29670_));
  NOR2_X1    g26444(.A1(new_n28249_), .A2(new_n11893_), .ZN(new_n29671_));
  OAI21_X1   g26445(.A1(new_n29353_), .A2(new_n29671_), .B(pi1155), .ZN(new_n29672_));
  NAND2_X1   g26446(.A1(new_n29435_), .A2(pi1155), .ZN(new_n29673_));
  NAND4_X1   g26447(.A1(new_n29670_), .A2(pi1154), .A3(new_n29672_), .A4(new_n29673_), .ZN(new_n29674_));
  NOR2_X1    g26448(.A1(new_n29157_), .A2(pi1153), .ZN(new_n29675_));
  NAND3_X1   g26449(.A1(new_n29675_), .A2(new_n11912_), .A3(new_n29209_), .ZN(new_n29676_));
  AND2_X2    g26450(.A1(new_n29672_), .A2(new_n11950_), .Z(new_n29677_));
  AOI21_X1   g26451(.A1(new_n29677_), .A2(new_n29676_), .B(pi0211), .ZN(new_n29678_));
  AOI21_X1   g26452(.A1(new_n29678_), .A2(new_n29674_), .B(pi0267), .ZN(new_n29679_));
  AOI21_X1   g26453(.A1(new_n29152_), .A2(new_n29480_), .B(new_n28170_), .ZN(new_n29680_));
  INV_X1     g26454(.I(new_n29675_), .ZN(new_n29681_));
  AOI21_X1   g26455(.A1(new_n29124_), .A2(new_n29681_), .B(new_n29474_), .ZN(new_n29682_));
  NOR3_X1    g26456(.A1(new_n28166_), .A2(new_n29296_), .A3(pi1155), .ZN(new_n29683_));
  NAND2_X1   g26457(.A1(new_n29682_), .A2(new_n29683_), .ZN(new_n29684_));
  AOI21_X1   g26458(.A1(new_n29684_), .A2(pi1154), .B(new_n29680_), .ZN(new_n29685_));
  NOR3_X1    g26459(.A1(new_n28241_), .A2(new_n28139_), .A3(new_n29310_), .ZN(new_n29686_));
  NOR3_X1    g26460(.A1(new_n29686_), .A2(new_n29352_), .A3(pi1155), .ZN(new_n29687_));
  NOR4_X1    g26461(.A1(new_n29679_), .A2(new_n8077_), .A3(new_n29685_), .A4(new_n29687_), .ZN(new_n29688_));
  OAI21_X1   g26462(.A1(pi1153), .A2(new_n29442_), .B(new_n29151_), .ZN(new_n29689_));
  NAND2_X1   g26463(.A1(new_n29689_), .A2(new_n11912_), .ZN(new_n29690_));
  NOR2_X1    g26464(.A1(new_n29194_), .A2(new_n11912_), .ZN(new_n29691_));
  NOR4_X1    g26465(.A1(new_n28129_), .A2(pi1154), .A3(new_n28135_), .A4(new_n28172_), .ZN(new_n29692_));
  AOI21_X1   g26466(.A1(new_n29692_), .A2(new_n29691_), .B(new_n28166_), .ZN(new_n29693_));
  NAND2_X1   g26467(.A1(new_n29681_), .A2(new_n11950_), .ZN(new_n29694_));
  NOR2_X1    g26468(.A1(new_n28143_), .A2(new_n28135_), .ZN(new_n29695_));
  OAI21_X1   g26469(.A1(new_n29694_), .A2(new_n29695_), .B(new_n11912_), .ZN(new_n29696_));
  NAND2_X1   g26470(.A1(new_n29696_), .A2(new_n28180_), .ZN(new_n29697_));
  AOI22_X1   g26471(.A1(new_n29697_), .A2(new_n29694_), .B1(new_n29690_), .B2(new_n29693_), .ZN(new_n29698_));
  NOR2_X1    g26472(.A1(new_n29689_), .A2(new_n11950_), .ZN(new_n29699_));
  OAI21_X1   g26473(.A1(new_n28174_), .A2(pi1153), .B(new_n28137_), .ZN(new_n29700_));
  AOI21_X1   g26474(.A1(new_n28129_), .A2(pi1154), .B(new_n11912_), .ZN(new_n29701_));
  NAND2_X1   g26475(.A1(new_n8077_), .A2(new_n28260_), .ZN(new_n29702_));
  AOI21_X1   g26476(.A1(new_n29701_), .A2(new_n29700_), .B(new_n29702_), .ZN(new_n29703_));
  OAI21_X1   g26477(.A1(new_n29696_), .A2(new_n29699_), .B(new_n29703_), .ZN(new_n29704_));
  NOR2_X1    g26478(.A1(new_n29698_), .A2(new_n29704_), .ZN(new_n29705_));
  OAI21_X1   g26479(.A1(new_n29688_), .A2(new_n29705_), .B(new_n8247_), .ZN(new_n29706_));
  OAI21_X1   g26480(.A1(pi1154), .A2(new_n28241_), .B(new_n28129_), .ZN(new_n29707_));
  OAI21_X1   g26481(.A1(new_n29194_), .A2(new_n11912_), .B(new_n28260_), .ZN(new_n29708_));
  AOI21_X1   g26482(.A1(new_n29201_), .A2(new_n29707_), .B(new_n29708_), .ZN(new_n29709_));
  NAND2_X1   g26483(.A1(new_n28232_), .A2(new_n11950_), .ZN(new_n29710_));
  OAI21_X1   g26484(.A1(new_n29203_), .A2(new_n29710_), .B(new_n11912_), .ZN(new_n29711_));
  NOR2_X1    g26485(.A1(new_n29682_), .A2(new_n11950_), .ZN(new_n29712_));
  NAND2_X1   g26486(.A1(new_n29712_), .A2(new_n29711_), .ZN(new_n29713_));
  INV_X1     g26487(.I(new_n29686_), .ZN(new_n29714_));
  NOR2_X1    g26488(.A1(new_n28241_), .A2(new_n28134_), .ZN(new_n29715_));
  AOI21_X1   g26489(.A1(new_n29715_), .A2(pi1154), .B(pi1155), .ZN(new_n29716_));
  AOI21_X1   g26490(.A1(new_n29716_), .A2(new_n29714_), .B(pi0267), .ZN(new_n29717_));
  NOR4_X1    g26491(.A1(new_n29129_), .A2(new_n11893_), .A3(new_n26910_), .A4(new_n28249_), .ZN(new_n29718_));
  NOR4_X1    g26492(.A1(new_n29717_), .A2(new_n11950_), .A3(new_n29297_), .A4(new_n29718_), .ZN(new_n29719_));
  NOR4_X1    g26493(.A1(new_n28152_), .A2(new_n29308_), .A3(new_n11950_), .A4(new_n11912_), .ZN(new_n29720_));
  NOR3_X1    g26494(.A1(new_n29686_), .A2(new_n28218_), .A3(pi1154), .ZN(new_n29721_));
  OAI21_X1   g26495(.A1(new_n29720_), .A2(new_n29721_), .B(pi0211), .ZN(new_n29722_));
  OAI22_X1   g26496(.A1(new_n29709_), .A2(new_n29713_), .B1(new_n29722_), .B2(new_n29719_), .ZN(new_n29723_));
  AOI21_X1   g26497(.A1(new_n29723_), .A2(pi0219), .B(new_n28264_), .ZN(new_n29724_));
  AOI22_X1   g26498(.A1(new_n27202_), .A2(new_n11912_), .B1(pi0219), .B2(pi0299), .ZN(new_n29725_));
  INV_X1     g26499(.I(new_n29725_), .ZN(new_n29726_));
  AOI21_X1   g26500(.A1(pi1155), .A2(new_n26434_), .B(new_n29726_), .ZN(new_n29727_));
  NOR2_X1    g26501(.A1(new_n26432_), .A2(new_n29259_), .ZN(new_n29728_));
  AOI21_X1   g26502(.A1(new_n26605_), .A2(pi1153), .B(new_n29270_), .ZN(new_n29729_));
  NAND2_X1   g26503(.A1(new_n29729_), .A2(new_n8077_), .ZN(new_n29730_));
  NOR2_X1    g26504(.A1(new_n29728_), .A2(new_n29730_), .ZN(new_n29731_));
  AOI21_X1   g26505(.A1(new_n26614_), .A2(pi1155), .B(new_n11950_), .ZN(new_n29732_));
  INV_X1     g26506(.I(new_n29732_), .ZN(new_n29733_));
  NOR4_X1    g26507(.A1(new_n29727_), .A2(new_n2918_), .A3(new_n29731_), .A4(new_n29733_), .ZN(new_n29734_));
  NOR4_X1    g26508(.A1(new_n27259_), .A2(new_n29729_), .A3(pi0219), .A4(new_n11912_), .ZN(new_n29735_));
  NOR3_X1    g26509(.A1(new_n29522_), .A2(new_n29103_), .A3(new_n29270_), .ZN(new_n29736_));
  NOR2_X1    g26510(.A1(new_n26625_), .A2(new_n8169_), .ZN(new_n29737_));
  INV_X1     g26511(.I(new_n29737_), .ZN(new_n29738_));
  NAND3_X1   g26512(.A1(new_n29736_), .A2(pi1091), .A3(new_n29738_), .ZN(new_n29739_));
  OAI21_X1   g26513(.A1(new_n29260_), .A2(new_n29080_), .B(pi1153), .ZN(new_n29740_));
  NOR2_X1    g26514(.A1(new_n26669_), .A2(pi1155), .ZN(new_n29741_));
  INV_X1     g26515(.I(new_n29741_), .ZN(new_n29742_));
  OAI22_X1   g26516(.A1(new_n2918_), .A2(new_n29742_), .B1(new_n29740_), .B2(new_n11912_), .ZN(new_n29743_));
  MUX2_X1    g26517(.I0(new_n29247_), .I1(new_n29074_), .S(new_n11893_), .Z(new_n29744_));
  NOR2_X1    g26518(.A1(new_n29104_), .A2(new_n11912_), .ZN(new_n29745_));
  AOI22_X1   g26519(.A1(new_n29744_), .A2(new_n11912_), .B1(new_n29257_), .B2(new_n29745_), .ZN(new_n29746_));
  MUX2_X1    g26520(.I0(new_n29746_), .I1(new_n29743_), .S(new_n11950_), .Z(new_n29747_));
  OAI22_X1   g26521(.A1(new_n29747_), .A2(pi0219), .B1(new_n29735_), .B2(new_n29739_), .ZN(new_n29748_));
  AOI21_X1   g26522(.A1(new_n29748_), .A2(new_n8077_), .B(new_n29734_), .ZN(new_n29749_));
  NOR2_X1    g26523(.A1(new_n29749_), .A2(new_n28260_), .ZN(new_n29750_));
  NOR4_X1    g26524(.A1(new_n29736_), .A2(new_n2918_), .A3(pi1155), .A4(new_n29738_), .ZN(new_n29751_));
  NOR2_X1    g26525(.A1(new_n29733_), .A2(new_n29522_), .ZN(new_n29752_));
  OAI21_X1   g26526(.A1(new_n29751_), .A2(new_n29752_), .B(pi0211), .ZN(new_n29753_));
  OAI21_X1   g26527(.A1(new_n27259_), .A2(new_n26432_), .B(new_n29270_), .ZN(new_n29754_));
  NOR3_X1    g26528(.A1(new_n29751_), .A2(new_n11950_), .A3(new_n9659_), .ZN(new_n29755_));
  NAND3_X1   g26529(.A1(new_n29755_), .A2(new_n29753_), .A3(new_n29754_), .ZN(new_n29756_));
  NOR2_X1    g26530(.A1(new_n26380_), .A2(pi1154), .ZN(new_n29757_));
  NOR3_X1    g26531(.A1(new_n26836_), .A2(new_n29757_), .A3(new_n26756_), .ZN(new_n29758_));
  OAI21_X1   g26532(.A1(new_n29758_), .A2(new_n2918_), .B(new_n8077_), .ZN(new_n29759_));
  NOR2_X1    g26533(.A1(new_n26963_), .A2(pi1091), .ZN(new_n29760_));
  OAI21_X1   g26534(.A1(new_n27202_), .A2(pi1155), .B(new_n29760_), .ZN(new_n29761_));
  NOR3_X1    g26535(.A1(new_n29522_), .A2(new_n2918_), .A3(new_n29103_), .ZN(new_n29762_));
  AOI21_X1   g26536(.A1(new_n29762_), .A2(new_n29761_), .B(pi0219), .ZN(new_n29763_));
  AOI21_X1   g26537(.A1(new_n29258_), .A2(new_n26390_), .B(new_n11893_), .ZN(new_n29764_));
  AOI21_X1   g26538(.A1(new_n29764_), .A2(pi1091), .B(new_n29741_), .ZN(new_n29765_));
  NOR3_X1    g26539(.A1(new_n29765_), .A2(new_n8077_), .A3(pi1154), .ZN(new_n29766_));
  AOI21_X1   g26540(.A1(new_n29763_), .A2(new_n29759_), .B(new_n29766_), .ZN(new_n29767_));
  AOI21_X1   g26541(.A1(new_n29756_), .A2(new_n29767_), .B(pi0267), .ZN(new_n29768_));
  NOR2_X1    g26542(.A1(new_n29750_), .A2(new_n29768_), .ZN(new_n29769_));
  NAND2_X1   g26543(.A1(new_n29769_), .A2(new_n28264_), .ZN(new_n29770_));
  NAND2_X1   g26544(.A1(new_n29770_), .A2(new_n6845_), .ZN(new_n29771_));
  AOI21_X1   g26545(.A1(new_n29706_), .A2(new_n29724_), .B(new_n29771_), .ZN(new_n29772_));
  NOR2_X1    g26546(.A1(new_n29330_), .A2(new_n29331_), .ZN(new_n29773_));
  NAND2_X1   g26547(.A1(new_n28119_), .A2(new_n28260_), .ZN(new_n29774_));
  OAI21_X1   g26548(.A1(new_n29166_), .A2(new_n29774_), .B(new_n28263_), .ZN(new_n29775_));
  NOR2_X1    g26549(.A1(new_n26911_), .A2(new_n8247_), .ZN(new_n29776_));
  AOI21_X1   g26550(.A1(new_n29283_), .A2(new_n26727_), .B(pi0219), .ZN(new_n29777_));
  OAI21_X1   g26551(.A1(new_n29777_), .A2(new_n29776_), .B(pi1091), .ZN(new_n29778_));
  AOI21_X1   g26552(.A1(new_n28264_), .A2(new_n28260_), .B(pi1091), .ZN(new_n29779_));
  NOR4_X1    g26553(.A1(po1038), .A2(new_n28260_), .A3(new_n28286_), .A4(new_n29779_), .ZN(new_n29780_));
  NAND4_X1   g26554(.A1(new_n29775_), .A2(new_n29773_), .A3(new_n29778_), .A4(new_n29780_), .ZN(new_n29781_));
  OAI21_X1   g26555(.A1(new_n28260_), .A2(pi1091), .B(new_n29778_), .ZN(new_n29782_));
  INV_X1     g26556(.I(new_n29782_), .ZN(new_n29783_));
  NOR3_X1    g26557(.A1(new_n29769_), .A2(po1038), .A3(new_n29783_), .ZN(new_n29784_));
  AOI21_X1   g26558(.A1(new_n29769_), .A2(new_n6845_), .B(new_n29782_), .ZN(new_n29785_));
  NOR3_X1    g26559(.A1(new_n29784_), .A2(new_n29785_), .A3(new_n28292_), .ZN(new_n29786_));
  OAI21_X1   g26560(.A1(new_n29772_), .A2(new_n29781_), .B(new_n29786_), .ZN(po0424));
  INV_X1     g26561(.I(new_n29050_), .ZN(new_n29788_));
  MUX2_X1    g26562(.I0(new_n29087_), .I1(new_n26396_), .S(new_n11749_), .Z(new_n29789_));
  NAND3_X1   g26563(.A1(new_n29789_), .A2(pi1151), .A3(pi1152), .ZN(new_n29790_));
  NOR2_X1    g26564(.A1(new_n6845_), .A2(new_n8663_), .ZN(new_n29791_));
  AOI21_X1   g26565(.A1(new_n6845_), .A2(new_n8666_), .B(new_n29791_), .ZN(new_n29792_));
  INV_X1     g26566(.I(new_n29792_), .ZN(new_n29793_));
  OAI21_X1   g26567(.A1(new_n29793_), .A2(new_n27251_), .B(new_n26604_), .ZN(new_n29794_));
  NAND2_X1   g26568(.A1(new_n29794_), .A2(new_n27817_), .ZN(new_n29795_));
  NAND4_X1   g26569(.A1(new_n29795_), .A2(new_n29790_), .A3(new_n27251_), .A4(new_n29788_), .ZN(new_n29796_));
  NAND2_X1   g26570(.A1(new_n27783_), .A2(new_n8077_), .ZN(new_n29797_));
  OAI21_X1   g26571(.A1(po1038), .A2(new_n26390_), .B(new_n29797_), .ZN(new_n29798_));
  NOR2_X1    g26572(.A1(new_n29798_), .A2(pi1151), .ZN(new_n29799_));
  INV_X1     g26573(.I(new_n29799_), .ZN(new_n29800_));
  NOR2_X1    g26574(.A1(new_n27783_), .A2(pi0199), .ZN(new_n29801_));
  NOR2_X1    g26575(.A1(new_n29801_), .A2(new_n27614_), .ZN(new_n29802_));
  INV_X1     g26576(.I(new_n29802_), .ZN(new_n29803_));
  NAND3_X1   g26577(.A1(new_n29803_), .A2(pi1152), .A3(new_n29798_), .ZN(new_n29804_));
  AOI21_X1   g26578(.A1(new_n29800_), .A2(pi1150), .B(new_n29804_), .ZN(new_n29805_));
  NOR2_X1    g26579(.A1(new_n29805_), .A2(new_n26307_), .ZN(new_n29806_));
  INV_X1     g26580(.I(new_n29168_), .ZN(new_n29807_));
  AOI21_X1   g26581(.A1(new_n28158_), .A2(new_n8247_), .B(po1038), .ZN(new_n29808_));
  NOR3_X1    g26582(.A1(new_n29133_), .A2(new_n29808_), .A3(new_n8247_), .ZN(new_n29809_));
  AOI21_X1   g26583(.A1(new_n28170_), .A2(new_n8247_), .B(new_n28126_), .ZN(new_n29810_));
  AOI22_X1   g26584(.A1(new_n29809_), .A2(new_n29810_), .B1(new_n6845_), .B2(new_n29807_), .ZN(new_n29811_));
  INV_X1     g26585(.I(new_n29811_), .ZN(new_n29812_));
  NOR3_X1    g26586(.A1(new_n29132_), .A2(new_n8247_), .A3(new_n28143_), .ZN(new_n29813_));
  NOR2_X1    g26587(.A1(new_n29193_), .A2(new_n28149_), .ZN(new_n29814_));
  NOR2_X1    g26588(.A1(new_n29813_), .A2(new_n29814_), .ZN(new_n29815_));
  INV_X1     g26589(.I(new_n29815_), .ZN(new_n29816_));
  NOR2_X1    g26590(.A1(new_n29198_), .A2(new_n29166_), .ZN(new_n29817_));
  MUX2_X1    g26591(.I0(new_n29817_), .I1(new_n29816_), .S(new_n6845_), .Z(new_n29818_));
  AOI21_X1   g26592(.A1(new_n29818_), .A2(new_n29812_), .B(new_n27251_), .ZN(new_n29819_));
  NOR2_X1    g26593(.A1(new_n29205_), .A2(new_n28250_), .ZN(new_n29820_));
  OAI21_X1   g26594(.A1(new_n29815_), .A2(new_n29820_), .B(new_n6845_), .ZN(new_n29821_));
  INV_X1     g26595(.I(new_n29821_), .ZN(new_n29822_));
  NOR2_X1    g26596(.A1(new_n6845_), .A2(new_n8247_), .ZN(new_n29823_));
  AOI22_X1   g26597(.A1(new_n29198_), .A2(po1038), .B1(new_n29170_), .B2(new_n29823_), .ZN(new_n29824_));
  NAND2_X1   g26598(.A1(new_n29822_), .A2(new_n29824_), .ZN(new_n29825_));
  AOI21_X1   g26599(.A1(new_n28116_), .A2(new_n8247_), .B(po1038), .ZN(new_n29826_));
  NAND3_X1   g26600(.A1(new_n29211_), .A2(new_n28187_), .A3(new_n29826_), .ZN(new_n29827_));
  INV_X1     g26601(.I(new_n29827_), .ZN(new_n29828_));
  OAI21_X1   g26602(.A1(pi1151), .A2(new_n29828_), .B(new_n29825_), .ZN(new_n29829_));
  INV_X1     g26603(.I(new_n29825_), .ZN(new_n29830_));
  NAND3_X1   g26604(.A1(new_n29830_), .A2(new_n27251_), .A3(new_n29828_), .ZN(new_n29831_));
  NAND3_X1   g26605(.A1(new_n29831_), .A2(new_n26604_), .A3(new_n29829_), .ZN(new_n29832_));
  AOI21_X1   g26606(.A1(pi1152), .A2(new_n29819_), .B(new_n29832_), .ZN(new_n29833_));
  OAI21_X1   g26607(.A1(new_n28195_), .A2(new_n8247_), .B(new_n6845_), .ZN(new_n29834_));
  AOI21_X1   g26608(.A1(pi0219), .A2(new_n28238_), .B(new_n29834_), .ZN(new_n29835_));
  NAND4_X1   g26609(.A1(new_n28108_), .A2(new_n28116_), .A3(pi0219), .A4(new_n6845_), .ZN(new_n29836_));
  NAND2_X1   g26610(.A1(new_n29835_), .A2(new_n29836_), .ZN(new_n29837_));
  INV_X1     g26611(.I(new_n29837_), .ZN(new_n29838_));
  NOR2_X1    g26612(.A1(new_n29838_), .A2(new_n28140_), .ZN(new_n29839_));
  OAI21_X1   g26613(.A1(new_n29839_), .A2(pi1151), .B(new_n26604_), .ZN(new_n29840_));
  NAND2_X1   g26614(.A1(new_n29139_), .A2(new_n6845_), .ZN(new_n29841_));
  OAI22_X1   g26615(.A1(new_n29144_), .A2(new_n29841_), .B1(new_n29181_), .B2(new_n29182_), .ZN(new_n29842_));
  INV_X1     g26616(.I(new_n29842_), .ZN(new_n29843_));
  NAND3_X1   g26617(.A1(new_n29843_), .A2(pi1151), .A3(new_n29840_), .ZN(new_n29844_));
  NOR2_X1    g26618(.A1(new_n29138_), .A2(new_n8247_), .ZN(new_n29845_));
  OAI21_X1   g26619(.A1(new_n29144_), .A2(new_n29845_), .B(new_n29146_), .ZN(new_n29846_));
  NOR2_X1    g26620(.A1(new_n29181_), .A2(new_n29330_), .ZN(new_n29847_));
  MUX2_X1    g26621(.I0(new_n29847_), .I1(new_n29846_), .S(new_n6845_), .Z(new_n29848_));
  INV_X1     g26622(.I(new_n29848_), .ZN(new_n29849_));
  AOI21_X1   g26623(.A1(new_n29121_), .A2(new_n8247_), .B(po1038), .ZN(new_n29850_));
  OAI21_X1   g26624(.A1(new_n29201_), .A2(pi0219), .B(new_n29850_), .ZN(new_n29851_));
  AOI21_X1   g26625(.A1(new_n29851_), .A2(new_n27251_), .B(pi1152), .ZN(new_n29852_));
  OAI21_X1   g26626(.A1(new_n29849_), .A2(new_n27251_), .B(new_n29852_), .ZN(new_n29853_));
  NAND4_X1   g26627(.A1(new_n29853_), .A2(new_n28280_), .A3(new_n27817_), .A4(new_n29844_), .ZN(new_n29854_));
  NOR2_X1    g26628(.A1(new_n29833_), .A2(new_n29854_), .ZN(new_n29855_));
  NOR2_X1    g26629(.A1(new_n29330_), .A2(new_n6845_), .ZN(new_n29856_));
  NOR3_X1    g26630(.A1(new_n29166_), .A2(new_n6845_), .A3(new_n29180_), .ZN(new_n29857_));
  INV_X1     g26631(.I(new_n29857_), .ZN(new_n29858_));
  AOI21_X1   g26632(.A1(new_n29143_), .A2(new_n29856_), .B(new_n29858_), .ZN(new_n29859_));
  OAI21_X1   g26633(.A1(new_n28146_), .A2(new_n2587_), .B(pi0219), .ZN(new_n29860_));
  AOI21_X1   g26634(.A1(new_n29145_), .A2(new_n29860_), .B(new_n28139_), .ZN(new_n29861_));
  AOI21_X1   g26635(.A1(new_n6845_), .A2(new_n29465_), .B(new_n29861_), .ZN(new_n29862_));
  NOR2_X1    g26636(.A1(new_n29862_), .A2(new_n29859_), .ZN(new_n29863_));
  INV_X1     g26637(.I(new_n29863_), .ZN(new_n29864_));
  NOR2_X1    g26638(.A1(new_n29864_), .A2(new_n27251_), .ZN(new_n29865_));
  NOR2_X1    g26639(.A1(new_n29137_), .A2(po1038), .ZN(new_n29866_));
  OAI22_X1   g26640(.A1(new_n29815_), .A2(new_n29866_), .B1(new_n29174_), .B2(new_n29182_), .ZN(new_n29867_));
  NOR4_X1    g26641(.A1(new_n29867_), .A2(pi0268), .A3(new_n27251_), .A4(new_n29838_), .ZN(new_n29868_));
  AOI21_X1   g26642(.A1(new_n29837_), .A2(new_n28140_), .B(new_n29828_), .ZN(new_n29869_));
  AOI21_X1   g26643(.A1(new_n29869_), .A2(pi1151), .B(pi0268), .ZN(new_n29870_));
  INV_X1     g26644(.I(new_n29870_), .ZN(new_n29871_));
  NOR3_X1    g26645(.A1(new_n29865_), .A2(new_n29868_), .A3(new_n29871_), .ZN(new_n29872_));
  INV_X1     g26646(.I(new_n29872_), .ZN(new_n29873_));
  INV_X1     g26647(.I(new_n29856_), .ZN(new_n29874_));
  NOR2_X1    g26648(.A1(new_n29189_), .A2(new_n28146_), .ZN(new_n29875_));
  OAI22_X1   g26649(.A1(new_n29822_), .A2(new_n29875_), .B1(new_n29174_), .B2(new_n29874_), .ZN(new_n29876_));
  NAND2_X1   g26650(.A1(new_n29876_), .A2(pi1151), .ZN(new_n29877_));
  NAND2_X1   g26651(.A1(new_n29874_), .A2(new_n29331_), .ZN(new_n29878_));
  NAND2_X1   g26652(.A1(new_n29835_), .A2(new_n29878_), .ZN(new_n29879_));
  OAI21_X1   g26653(.A1(pi1091), .A2(new_n28103_), .B(new_n29866_), .ZN(new_n29880_));
  NAND2_X1   g26654(.A1(new_n29880_), .A2(new_n29879_), .ZN(new_n29881_));
  INV_X1     g26655(.I(new_n29881_), .ZN(new_n29882_));
  NAND2_X1   g26656(.A1(new_n29882_), .A2(pi1151), .ZN(new_n29883_));
  AOI21_X1   g26657(.A1(new_n29877_), .A2(new_n29883_), .B(new_n28280_), .ZN(new_n29884_));
  OAI21_X1   g26658(.A1(new_n29861_), .A2(new_n29131_), .B(new_n6845_), .ZN(new_n29885_));
  NAND2_X1   g26659(.A1(new_n29885_), .A2(new_n29858_), .ZN(new_n29886_));
  NOR2_X1    g26660(.A1(new_n29817_), .A2(po1038), .ZN(new_n29887_));
  NOR2_X1    g26661(.A1(new_n29887_), .A2(new_n29859_), .ZN(new_n29888_));
  NOR2_X1    g26662(.A1(new_n29809_), .A2(new_n29888_), .ZN(new_n29889_));
  MUX2_X1    g26663(.I0(new_n29889_), .I1(new_n29886_), .S(new_n27251_), .Z(new_n29890_));
  AOI21_X1   g26664(.A1(new_n28280_), .A2(new_n29890_), .B(new_n29884_), .ZN(new_n29891_));
  AOI21_X1   g26665(.A1(new_n29891_), .A2(pi1152), .B(new_n29873_), .ZN(new_n29892_));
  NOR3_X1    g26666(.A1(new_n29891_), .A2(new_n26604_), .A3(new_n29872_), .ZN(new_n29893_));
  NOR3_X1    g26667(.A1(new_n29892_), .A2(new_n29893_), .A3(new_n27817_), .ZN(new_n29894_));
  OAI21_X1   g26668(.A1(new_n29894_), .A2(new_n29855_), .B(new_n28284_), .ZN(new_n29895_));
  NAND4_X1   g26669(.A1(new_n29805_), .A2(new_n28280_), .A3(new_n2918_), .A4(pi1152), .ZN(new_n29896_));
  NOR3_X1    g26670(.A1(new_n29805_), .A2(new_n28280_), .A3(new_n26604_), .ZN(new_n29897_));
  NAND2_X1   g26671(.A1(new_n29796_), .A2(pi1091), .ZN(new_n29898_));
  OAI21_X1   g26672(.A1(new_n29897_), .A2(new_n29898_), .B(new_n29896_), .ZN(new_n29899_));
  AOI21_X1   g26673(.A1(new_n29899_), .A2(new_n28285_), .B(pi0230), .ZN(new_n29900_));
  AOI22_X1   g26674(.A1(new_n29895_), .A2(new_n29900_), .B1(new_n29796_), .B2(new_n29806_), .ZN(po0425));
  NOR2_X1    g26675(.A1(new_n11749_), .A2(new_n8247_), .ZN(new_n29902_));
  NOR3_X1    g26676(.A1(new_n29902_), .A2(new_n4261_), .A3(new_n29077_), .ZN(new_n29903_));
  NAND2_X1   g26677(.A1(new_n11749_), .A2(pi0199), .ZN(new_n29904_));
  AOI21_X1   g26678(.A1(pi1138), .A2(new_n29601_), .B(new_n29904_), .ZN(new_n29905_));
  AND3_X2    g26679(.A1(new_n28102_), .A2(pi0269), .A3(pi0817), .Z(new_n29906_));
  INV_X1     g26680(.I(pi0817), .ZN(new_n29907_));
  OAI21_X1   g26681(.A1(new_n28101_), .A2(pi0269), .B(new_n29907_), .ZN(new_n29908_));
  NAND2_X1   g26682(.A1(new_n29908_), .A2(new_n2918_), .ZN(new_n29909_));
  NOR4_X1    g26683(.A1(new_n29905_), .A2(new_n29903_), .A3(new_n29906_), .A4(new_n29909_), .ZN(new_n29910_));
  NOR2_X1    g26684(.A1(new_n8077_), .A2(pi1137), .ZN(new_n29911_));
  NOR2_X1    g26685(.A1(pi0211), .A2(pi1136), .ZN(new_n29912_));
  NOR3_X1    g26686(.A1(new_n29911_), .A2(new_n2918_), .A3(new_n29912_), .ZN(new_n29913_));
  NOR2_X1    g26687(.A1(new_n27615_), .A2(new_n29913_), .ZN(new_n29914_));
  NAND3_X1   g26688(.A1(new_n4543_), .A2(pi0200), .A3(pi1137), .ZN(new_n29915_));
  OAI21_X1   g26689(.A1(new_n8098_), .A2(pi1137), .B(pi1136), .ZN(new_n29916_));
  AOI21_X1   g26690(.A1(new_n29916_), .A2(new_n29915_), .B(new_n2918_), .ZN(new_n29917_));
  NAND2_X1   g26691(.A1(new_n29801_), .A2(new_n29917_), .ZN(new_n29918_));
  NAND3_X1   g26692(.A1(new_n28111_), .A2(pi0269), .A3(pi0817), .ZN(new_n29919_));
  OAI21_X1   g26693(.A1(new_n29584_), .A2(pi0269), .B(new_n29907_), .ZN(new_n29920_));
  NAND4_X1   g26694(.A1(new_n29918_), .A2(new_n2918_), .A3(new_n29919_), .A4(new_n29920_), .ZN(new_n29921_));
  OAI21_X1   g26695(.A1(new_n29921_), .A2(new_n29914_), .B(new_n26307_), .ZN(new_n29922_));
  OAI21_X1   g26696(.A1(pi0199), .A2(pi1136), .B(pi1138), .ZN(new_n29923_));
  NAND3_X1   g26697(.A1(new_n8094_), .A2(new_n4261_), .A3(pi1136), .ZN(new_n29924_));
  NAND2_X1   g26698(.A1(new_n8160_), .A2(pi1137), .ZN(new_n29925_));
  NAND4_X1   g26699(.A1(new_n29925_), .A2(new_n29924_), .A3(new_n8098_), .A4(new_n29923_), .ZN(new_n29926_));
  NOR2_X1    g26700(.A1(new_n27783_), .A2(new_n29926_), .ZN(new_n29927_));
  OAI22_X1   g26701(.A1(new_n29922_), .A2(new_n29910_), .B1(new_n26307_), .B2(new_n29927_), .ZN(po0426));
  OAI21_X1   g26702(.A1(pi0199), .A2(pi1139), .B(pi1141), .ZN(new_n29929_));
  NOR3_X1    g26703(.A1(new_n4115_), .A2(pi0199), .A3(pi1141), .ZN(new_n29930_));
  NOR2_X1    g26704(.A1(new_n3973_), .A2(pi0199), .ZN(new_n29931_));
  NOR3_X1    g26705(.A1(new_n29930_), .A2(new_n29931_), .A3(pi0200), .ZN(new_n29932_));
  AOI21_X1   g26706(.A1(new_n29929_), .A2(new_n29932_), .B(new_n27783_), .ZN(new_n29933_));
  NOR3_X1    g26707(.A1(new_n29902_), .A2(new_n3831_), .A3(new_n29077_), .ZN(new_n29934_));
  NOR4_X1    g26708(.A1(new_n27783_), .A2(pi0199), .A3(new_n3831_), .A4(new_n29602_), .ZN(new_n29935_));
  INV_X1     g26709(.I(pi0270), .ZN(new_n29936_));
  INV_X1     g26710(.I(pi0805), .ZN(new_n29937_));
  NOR3_X1    g26711(.A1(new_n28101_), .A2(new_n29936_), .A3(new_n29937_), .ZN(new_n29938_));
  AOI21_X1   g26712(.A1(new_n28102_), .A2(new_n29936_), .B(pi0805), .ZN(new_n29939_));
  NOR3_X1    g26713(.A1(new_n29939_), .A2(pi1091), .A3(new_n29938_), .ZN(new_n29940_));
  OAI21_X1   g26714(.A1(new_n29934_), .A2(new_n29935_), .B(new_n29940_), .ZN(new_n29941_));
  INV_X1     g26715(.I(new_n29801_), .ZN(new_n29942_));
  NOR2_X1    g26716(.A1(new_n8077_), .A2(pi1140), .ZN(new_n29943_));
  NOR2_X1    g26717(.A1(pi0211), .A2(pi1139), .ZN(new_n29944_));
  NOR3_X1    g26718(.A1(new_n29943_), .A2(new_n2918_), .A3(new_n29944_), .ZN(new_n29945_));
  MUX2_X1    g26719(.I0(pi1139), .I1(pi1140), .S(pi0200), .Z(new_n29946_));
  NAND2_X1   g26720(.A1(new_n29946_), .A2(pi1091), .ZN(new_n29947_));
  OAI22_X1   g26721(.A1(new_n29942_), .A2(new_n29947_), .B1(new_n27615_), .B2(new_n29945_), .ZN(new_n29948_));
  NOR3_X1    g26722(.A1(new_n29584_), .A2(new_n29936_), .A3(new_n29937_), .ZN(new_n29949_));
  AOI21_X1   g26723(.A1(new_n28111_), .A2(new_n29936_), .B(pi0805), .ZN(new_n29950_));
  NOR3_X1    g26724(.A1(new_n29949_), .A2(pi1091), .A3(new_n29950_), .ZN(new_n29951_));
  AOI21_X1   g26725(.A1(new_n29948_), .A2(new_n29951_), .B(pi0230), .ZN(new_n29952_));
  AOI22_X1   g26726(.A1(new_n29952_), .A2(new_n29941_), .B1(pi0230), .B2(new_n29933_), .ZN(po0427));
  NOR2_X1    g26727(.A1(new_n28104_), .A2(pi0271), .ZN(new_n29954_));
  NOR2_X1    g26728(.A1(new_n28103_), .A2(new_n28096_), .ZN(new_n29955_));
  OAI21_X1   g26729(.A1(new_n29954_), .A2(new_n29955_), .B(new_n2918_), .ZN(new_n29956_));
  INV_X1     g26730(.I(new_n29956_), .ZN(new_n29957_));
  XOR2_X1    g26731(.A1(new_n28112_), .A2(pi0271), .Z(new_n29958_));
  NAND2_X1   g26732(.A1(new_n29958_), .A2(new_n2918_), .ZN(new_n29959_));
  OAI21_X1   g26733(.A1(new_n2918_), .A2(new_n3258_), .B(new_n29959_), .ZN(new_n29960_));
  MUX2_X1    g26734(.I0(new_n29960_), .I1(new_n29957_), .S(pi0199), .Z(new_n29961_));
  NOR2_X1    g26735(.A1(new_n29961_), .A2(new_n8098_), .ZN(new_n29962_));
  NAND3_X1   g26736(.A1(pi0199), .A2(pi1091), .A3(pi1147), .ZN(new_n29963_));
  NAND2_X1   g26737(.A1(new_n29956_), .A2(pi0199), .ZN(new_n29964_));
  NAND2_X1   g26738(.A1(pi1091), .A2(pi1145), .ZN(new_n29965_));
  AND3_X2    g26739(.A1(new_n29959_), .A2(new_n8094_), .A3(new_n29965_), .Z(new_n29966_));
  AOI22_X1   g26740(.A1(new_n29966_), .A2(new_n29964_), .B1(new_n8098_), .B2(new_n29963_), .ZN(new_n29967_));
  OAI21_X1   g26741(.A1(new_n29962_), .A2(new_n29967_), .B(new_n11749_), .ZN(new_n29968_));
  NOR2_X1    g26742(.A1(new_n29077_), .A2(new_n3258_), .ZN(new_n29969_));
  INV_X1     g26743(.I(new_n29969_), .ZN(new_n29970_));
  AOI22_X1   g26744(.A1(new_n29960_), .A2(new_n29970_), .B1(pi1145), .B2(new_n29076_), .ZN(new_n29971_));
  NOR4_X1    g26745(.A1(new_n8247_), .A2(new_n2918_), .A3(new_n27494_), .A4(pi0211), .ZN(new_n29972_));
  AOI21_X1   g26746(.A1(new_n29957_), .A2(pi0219), .B(new_n29972_), .ZN(new_n29973_));
  OAI21_X1   g26747(.A1(new_n29971_), .A2(pi0219), .B(new_n29973_), .ZN(new_n29974_));
  AOI21_X1   g26748(.A1(new_n29974_), .A2(new_n27783_), .B(pi0230), .ZN(new_n29975_));
  NAND2_X1   g26749(.A1(new_n29968_), .A2(new_n29975_), .ZN(po0428));
  OAI21_X1   g26750(.A1(new_n29788_), .A2(new_n27817_), .B(new_n27470_), .ZN(new_n29977_));
  NAND2_X1   g26751(.A1(new_n29977_), .A2(new_n27515_), .ZN(new_n29978_));
  AND2_X2    g26752(.A1(new_n6845_), .A2(new_n9660_), .Z(new_n29979_));
  NOR2_X1    g26753(.A1(new_n6845_), .A2(new_n9658_), .ZN(new_n29980_));
  XOR2_X1    g26754(.A1(new_n29979_), .A2(new_n29980_), .Z(new_n29981_));
  INV_X1     g26755(.I(new_n29981_), .ZN(new_n29982_));
  NAND2_X1   g26756(.A1(new_n29982_), .A2(new_n27817_), .ZN(new_n29983_));
  AOI21_X1   g26757(.A1(new_n29983_), .A2(new_n29798_), .B(pi1149), .ZN(new_n29984_));
  NAND2_X1   g26758(.A1(po1038), .A2(new_n26493_), .ZN(new_n29985_));
  NAND4_X1   g26759(.A1(new_n27615_), .A2(new_n29797_), .A3(pi1150), .A4(new_n29985_), .ZN(new_n29986_));
  NAND4_X1   g26760(.A1(new_n29986_), .A2(new_n27515_), .A3(pi1149), .A4(new_n29802_), .ZN(new_n29987_));
  NOR2_X1    g26761(.A1(new_n29984_), .A2(new_n29987_), .ZN(new_n29988_));
  OAI21_X1   g26762(.A1(new_n29986_), .A2(new_n29789_), .B(pi1149), .ZN(new_n29989_));
  NOR2_X1    g26763(.A1(new_n29793_), .A2(pi1150), .ZN(new_n29990_));
  NOR4_X1    g26764(.A1(new_n29988_), .A2(pi0230), .A3(new_n29989_), .A4(new_n29990_), .ZN(new_n29991_));
  NAND2_X1   g26765(.A1(new_n29991_), .A2(new_n29978_), .ZN(new_n29992_));
  INV_X1     g26766(.I(new_n29818_), .ZN(new_n29993_));
  MUX2_X1    g26767(.I0(new_n29830_), .I1(new_n29993_), .S(pi1150), .Z(new_n29994_));
  NAND2_X1   g26768(.A1(pi1149), .A2(pi1150), .ZN(new_n29995_));
  OAI22_X1   g26769(.A1(new_n29994_), .A2(new_n27470_), .B1(new_n29811_), .B2(new_n29995_), .ZN(new_n29996_));
  NAND3_X1   g26770(.A1(new_n29863_), .A2(pi1150), .A3(new_n29886_), .ZN(new_n29997_));
  OAI21_X1   g26771(.A1(new_n27817_), .A2(new_n29886_), .B(new_n29864_), .ZN(new_n29998_));
  AOI21_X1   g26772(.A1(new_n29998_), .A2(new_n29997_), .B(pi1149), .ZN(new_n29999_));
  INV_X1     g26773(.I(new_n29869_), .ZN(new_n30000_));
  INV_X1     g26774(.I(new_n29889_), .ZN(new_n30001_));
  MUX2_X1    g26775(.I0(new_n30001_), .I1(new_n30000_), .S(new_n27817_), .Z(new_n30002_));
  OAI21_X1   g26776(.A1(new_n30002_), .A2(new_n27470_), .B(pi1148), .ZN(new_n30003_));
  INV_X1     g26777(.I(new_n29789_), .ZN(new_n30004_));
  NOR2_X1    g26778(.A1(new_n28283_), .A2(pi0272), .ZN(new_n30008_));
  OAI21_X1   g26779(.A1(new_n29999_), .A2(new_n30003_), .B(new_n30008_), .ZN(new_n30009_));
  AOI21_X1   g26780(.A1(new_n29996_), .A2(new_n27515_), .B(new_n30009_), .ZN(new_n30010_));
  INV_X1     g26781(.I(new_n29867_), .ZN(new_n30011_));
  AOI21_X1   g26782(.A1(new_n27817_), .A2(new_n30011_), .B(new_n29876_), .ZN(new_n30012_));
  AND3_X2    g26783(.A1(new_n29876_), .A2(new_n27817_), .A3(new_n29867_), .Z(new_n30013_));
  NOR2_X1    g26784(.A1(new_n29882_), .A2(new_n27817_), .ZN(new_n30014_));
  NOR2_X1    g26785(.A1(new_n29838_), .A2(pi1150), .ZN(new_n30015_));
  OAI21_X1   g26786(.A1(new_n30014_), .A2(new_n30015_), .B(new_n27470_), .ZN(new_n30016_));
  NOR3_X1    g26787(.A1(new_n30013_), .A2(new_n30012_), .A3(new_n30016_), .ZN(new_n30017_));
  NAND2_X1   g26788(.A1(new_n29848_), .A2(pi1150), .ZN(new_n30018_));
  AOI21_X1   g26789(.A1(new_n29842_), .A2(new_n27817_), .B(pi1149), .ZN(new_n30019_));
  OAI21_X1   g26790(.A1(new_n29839_), .A2(pi1150), .B(new_n27470_), .ZN(new_n30020_));
  NOR2_X1    g26791(.A1(new_n29851_), .A2(new_n27817_), .ZN(new_n30021_));
  AOI22_X1   g26792(.A1(new_n30018_), .A2(new_n30019_), .B1(new_n30020_), .B2(new_n30021_), .ZN(new_n30022_));
  NAND2_X1   g26793(.A1(new_n28283_), .A2(new_n27515_), .ZN(new_n30023_));
  OAI21_X1   g26794(.A1(new_n30022_), .A2(new_n30023_), .B(pi1148), .ZN(new_n30024_));
  AOI21_X1   g26795(.A1(new_n28699_), .A2(new_n29798_), .B(new_n29803_), .ZN(new_n30025_));
  NOR2_X1    g26796(.A1(new_n2918_), .A2(pi1148), .ZN(new_n30026_));
  OAI21_X1   g26797(.A1(new_n29984_), .A2(new_n30025_), .B(new_n30026_), .ZN(new_n30027_));
  NOR2_X1    g26798(.A1(new_n30004_), .A2(new_n2918_), .ZN(new_n30028_));
  NAND2_X1   g26799(.A1(new_n26635_), .A2(new_n29068_), .ZN(new_n30029_));
  OAI22_X1   g26800(.A1(new_n11749_), .A2(new_n29267_), .B1(po1038), .B2(new_n30029_), .ZN(new_n30030_));
  INV_X1     g26801(.I(new_n30030_), .ZN(new_n30031_));
  NAND4_X1   g26802(.A1(new_n30028_), .A2(new_n27470_), .A3(pi1150), .A4(new_n30031_), .ZN(new_n30032_));
  NOR4_X1    g26803(.A1(new_n29050_), .A2(pi1091), .A3(pi1149), .A4(pi1150), .ZN(new_n30033_));
  NOR2_X1    g26804(.A1(new_n30033_), .A2(pi1148), .ZN(new_n30034_));
  AOI21_X1   g26805(.A1(new_n30032_), .A2(new_n30034_), .B(pi0283), .ZN(new_n30035_));
  NAND2_X1   g26806(.A1(new_n26307_), .A2(pi0272), .ZN(new_n30036_));
  AOI21_X1   g26807(.A1(new_n30035_), .A2(new_n30027_), .B(new_n30036_), .ZN(new_n30037_));
  OAI21_X1   g26808(.A1(new_n30017_), .A2(new_n30024_), .B(new_n30037_), .ZN(new_n30038_));
  OAI21_X1   g26809(.A1(new_n30010_), .A2(new_n30038_), .B(new_n29992_), .ZN(po0429));
  OAI21_X1   g26810(.A1(pi1146), .A2(new_n8161_), .B(new_n29801_), .ZN(new_n30040_));
  OAI21_X1   g26811(.A1(pi0211), .A2(new_n27506_), .B(new_n27614_), .ZN(new_n30041_));
  AOI21_X1   g26812(.A1(new_n30040_), .A2(new_n30041_), .B(pi1147), .ZN(new_n30042_));
  NOR3_X1    g26813(.A1(new_n29982_), .A2(new_n3258_), .A3(new_n28485_), .ZN(new_n30043_));
  NAND2_X1   g26814(.A1(new_n9658_), .A2(new_n3258_), .ZN(new_n30044_));
  NAND3_X1   g26815(.A1(new_n30044_), .A2(new_n26307_), .A3(new_n27515_), .ZN(new_n30045_));
  NAND2_X1   g26816(.A1(new_n27494_), .A2(pi0199), .ZN(new_n30046_));
  NAND2_X1   g26817(.A1(new_n3258_), .A2(pi1147), .ZN(new_n30047_));
  AOI21_X1   g26818(.A1(new_n27494_), .A2(pi1146), .B(pi0199), .ZN(new_n30048_));
  AOI21_X1   g26819(.A1(new_n30048_), .A2(new_n30047_), .B(pi0200), .ZN(new_n30049_));
  XOR2_X1    g26820(.A1(new_n30049_), .A2(new_n30046_), .Z(new_n30050_));
  OAI21_X1   g26821(.A1(new_n27783_), .A2(new_n30050_), .B(pi1148), .ZN(new_n30051_));
  OAI21_X1   g26822(.A1(new_n27494_), .A2(new_n27615_), .B(new_n29797_), .ZN(new_n30052_));
  NAND2_X1   g26823(.A1(new_n30052_), .A2(new_n30051_), .ZN(new_n30053_));
  NOR4_X1    g26824(.A1(new_n30042_), .A2(new_n30043_), .A3(new_n30053_), .A4(new_n30045_), .ZN(new_n30054_));
  INV_X1     g26825(.I(new_n28107_), .ZN(new_n30055_));
  XOR2_X1    g26826(.A1(new_n28115_), .A2(pi0273), .Z(new_n30056_));
  NAND2_X1   g26827(.A1(new_n30056_), .A2(new_n30055_), .ZN(new_n30057_));
  OAI21_X1   g26828(.A1(new_n29602_), .A2(new_n3258_), .B(new_n8094_), .ZN(new_n30058_));
  NAND2_X1   g26829(.A1(new_n28105_), .A2(new_n28095_), .ZN(new_n30059_));
  NAND2_X1   g26830(.A1(new_n28106_), .A2(pi0273), .ZN(new_n30060_));
  AOI21_X1   g26831(.A1(new_n30060_), .A2(new_n30059_), .B(pi1091), .ZN(new_n30061_));
  OAI21_X1   g26832(.A1(new_n30061_), .A2(new_n8094_), .B(new_n2587_), .ZN(new_n30062_));
  AOI21_X1   g26833(.A1(new_n30057_), .A2(new_n30058_), .B(new_n30062_), .ZN(new_n30063_));
  NAND2_X1   g26834(.A1(new_n30061_), .A2(pi0219), .ZN(new_n30064_));
  AOI21_X1   g26835(.A1(new_n30056_), .A2(new_n30055_), .B(new_n29969_), .ZN(new_n30065_));
  OAI21_X1   g26836(.A1(new_n30065_), .A2(pi0219), .B(new_n30064_), .ZN(new_n30066_));
  AOI21_X1   g26837(.A1(new_n30066_), .A2(pi0299), .B(new_n30063_), .ZN(new_n30067_));
  OR3_X2     g26838(.A1(new_n30067_), .A2(new_n2918_), .A3(new_n8665_), .Z(new_n30068_));
  AOI21_X1   g26839(.A1(new_n29183_), .A2(pi1091), .B(po1038), .ZN(new_n30069_));
  OAI21_X1   g26840(.A1(new_n29715_), .A2(new_n30068_), .B(new_n30069_), .ZN(new_n30070_));
  NAND2_X1   g26841(.A1(new_n30070_), .A2(pi1147), .ZN(new_n30071_));
  NOR3_X1    g26842(.A1(new_n29961_), .A2(new_n8098_), .A3(new_n29247_), .ZN(new_n30072_));
  AOI21_X1   g26843(.A1(pi1091), .A2(new_n26355_), .B(new_n30066_), .ZN(new_n30073_));
  NOR2_X1    g26844(.A1(new_n30063_), .A2(po1038), .ZN(new_n30074_));
  OAI21_X1   g26845(.A1(new_n30073_), .A2(new_n2587_), .B(new_n30074_), .ZN(new_n30075_));
  NOR2_X1    g26846(.A1(new_n29077_), .A2(new_n8247_), .ZN(new_n30076_));
  AOI21_X1   g26847(.A1(po1038), .A2(new_n30076_), .B(new_n27515_), .ZN(new_n30077_));
  OAI21_X1   g26848(.A1(new_n30075_), .A2(new_n30072_), .B(new_n30077_), .ZN(new_n30078_));
  OAI21_X1   g26849(.A1(new_n30067_), .A2(new_n28322_), .B(new_n27515_), .ZN(new_n30079_));
  AOI22_X1   g26850(.A1(new_n30078_), .A2(new_n30079_), .B1(po1038), .B2(new_n30066_), .ZN(new_n30080_));
  NAND2_X1   g26851(.A1(new_n30071_), .A2(new_n30080_), .ZN(new_n30081_));
  AOI21_X1   g26852(.A1(new_n30081_), .A2(new_n26307_), .B(new_n30054_), .ZN(po0430));
  NOR2_X1    g26853(.A1(new_n26321_), .A2(new_n27712_), .ZN(new_n30083_));
  OAI21_X1   g26854(.A1(new_n27489_), .A2(pi0211), .B(new_n26998_), .ZN(new_n30084_));
  OAI21_X1   g26855(.A1(pi0211), .A2(pi1143), .B(pi1144), .ZN(new_n30085_));
  INV_X1     g26856(.I(new_n30085_), .ZN(new_n30086_));
  NOR3_X1    g26857(.A1(new_n3548_), .A2(pi0211), .A3(pi1144), .ZN(new_n30087_));
  NOR3_X1    g26858(.A1(new_n30086_), .A2(new_n30087_), .A3(pi0219), .ZN(new_n30088_));
  AOI22_X1   g26859(.A1(new_n30084_), .A2(new_n30088_), .B1(new_n28052_), .B2(new_n30083_), .ZN(new_n30089_));
  INV_X1     g26860(.I(new_n30088_), .ZN(new_n30090_));
  NOR2_X1    g26861(.A1(new_n27471_), .A2(new_n30090_), .ZN(new_n30091_));
  NOR4_X1    g26862(.A1(new_n30091_), .A2(new_n26307_), .A3(po1038), .A4(new_n30089_), .ZN(new_n30092_));
  INV_X1     g26863(.I(pi0659), .ZN(new_n30093_));
  NOR3_X1    g26864(.A1(new_n29584_), .A2(new_n3434_), .A3(new_n30093_), .ZN(new_n30094_));
  AOI21_X1   g26865(.A1(new_n28111_), .A2(new_n3434_), .B(pi0659), .ZN(new_n30095_));
  NOR3_X1    g26866(.A1(new_n30094_), .A2(pi1091), .A3(new_n30095_), .ZN(new_n30096_));
  AOI21_X1   g26867(.A1(new_n30096_), .A2(new_n29613_), .B(pi0200), .ZN(new_n30097_));
  OAI21_X1   g26868(.A1(new_n2918_), .A2(new_n2552_), .B(new_n30096_), .ZN(new_n30098_));
  NAND2_X1   g26869(.A1(new_n30098_), .A2(pi0200), .ZN(new_n30099_));
  NAND2_X1   g26870(.A1(new_n30099_), .A2(new_n8094_), .ZN(new_n30100_));
  NOR3_X1    g26871(.A1(new_n28101_), .A2(new_n3434_), .A3(new_n30093_), .ZN(new_n30101_));
  AOI21_X1   g26872(.A1(new_n28102_), .A2(new_n3434_), .B(pi0659), .ZN(new_n30102_));
  NOR3_X1    g26873(.A1(new_n30102_), .A2(pi1091), .A3(new_n30101_), .ZN(new_n30103_));
  NOR3_X1    g26874(.A1(new_n29602_), .A2(pi0199), .A3(new_n3414_), .ZN(new_n30104_));
  NOR3_X1    g26875(.A1(new_n11749_), .A2(new_n30103_), .A3(new_n30104_), .ZN(new_n30105_));
  OAI21_X1   g26876(.A1(new_n30100_), .A2(new_n30097_), .B(new_n30105_), .ZN(new_n30106_));
  NAND2_X1   g26877(.A1(new_n30096_), .A2(new_n29613_), .ZN(new_n30107_));
  NAND2_X1   g26878(.A1(new_n30107_), .A2(new_n8077_), .ZN(new_n30108_));
  AOI21_X1   g26879(.A1(new_n30098_), .A2(pi0211), .B(pi0219), .ZN(new_n30109_));
  AOI21_X1   g26880(.A1(new_n29076_), .A2(pi1145), .B(new_n8247_), .ZN(new_n30110_));
  NOR2_X1    g26881(.A1(new_n11749_), .A2(pi0230), .ZN(new_n30111_));
  OAI21_X1   g26882(.A1(new_n30103_), .A2(new_n30110_), .B(new_n30111_), .ZN(new_n30112_));
  AOI21_X1   g26883(.A1(new_n30109_), .A2(new_n30108_), .B(new_n30112_), .ZN(new_n30113_));
  AOI21_X1   g26884(.A1(new_n30106_), .A2(new_n30113_), .B(new_n30092_), .ZN(po0431));
  NAND3_X1   g26885(.A1(new_n29800_), .A2(pi1149), .A3(new_n29802_), .ZN(new_n30115_));
  OAI21_X1   g26886(.A1(new_n28699_), .A2(new_n29798_), .B(new_n30115_), .ZN(new_n30116_));
  NAND2_X1   g26887(.A1(new_n29050_), .A2(new_n27817_), .ZN(new_n30117_));
  AOI21_X1   g26888(.A1(new_n30117_), .A2(new_n27251_), .B(pi1149), .ZN(new_n30118_));
  NOR4_X1    g26889(.A1(new_n29789_), .A2(new_n29793_), .A3(pi1150), .A4(new_n27251_), .ZN(new_n30119_));
  OAI21_X1   g26890(.A1(new_n30118_), .A2(new_n30119_), .B(new_n30116_), .ZN(new_n30120_));
  OR2_X2     g26891(.A1(new_n30120_), .A2(new_n26307_), .Z(new_n30121_));
  INV_X1     g26892(.I(new_n29851_), .ZN(new_n30122_));
  MUX2_X1    g26893(.I0(new_n30122_), .I1(new_n29849_), .S(pi1150), .Z(new_n30123_));
  NAND3_X1   g26894(.A1(new_n29843_), .A2(new_n27817_), .A3(new_n29839_), .ZN(new_n30124_));
  OAI21_X1   g26895(.A1(new_n29839_), .A2(pi1150), .B(new_n29842_), .ZN(new_n30125_));
  NAND3_X1   g26896(.A1(new_n30124_), .A2(new_n27251_), .A3(new_n30125_), .ZN(new_n30126_));
  AOI21_X1   g26897(.A1(new_n30123_), .A2(pi1151), .B(new_n30126_), .ZN(new_n30127_));
  NAND4_X1   g26898(.A1(new_n29818_), .A2(pi1150), .A3(new_n27251_), .A4(new_n29811_), .ZN(new_n30128_));
  AOI21_X1   g26899(.A1(new_n29827_), .A2(new_n27817_), .B(pi1151), .ZN(new_n30129_));
  OAI21_X1   g26900(.A1(new_n29825_), .A2(new_n27817_), .B(new_n30129_), .ZN(new_n30130_));
  NAND2_X1   g26901(.A1(new_n30130_), .A2(new_n30128_), .ZN(new_n30131_));
  NAND4_X1   g26902(.A1(new_n30127_), .A2(new_n28282_), .A3(new_n27470_), .A4(new_n30131_), .ZN(new_n30132_));
  NAND2_X1   g26903(.A1(pi0272), .A2(pi0283), .ZN(new_n30133_));
  NAND3_X1   g26904(.A1(new_n29863_), .A2(pi1150), .A3(new_n29869_), .ZN(new_n30134_));
  OAI21_X1   g26905(.A1(new_n27817_), .A2(new_n29869_), .B(new_n29864_), .ZN(new_n30135_));
  AOI21_X1   g26906(.A1(new_n30135_), .A2(new_n30134_), .B(pi1151), .ZN(new_n30136_));
  INV_X1     g26907(.I(new_n29886_), .ZN(new_n30137_));
  OAI21_X1   g26908(.A1(new_n30137_), .A2(new_n29889_), .B(pi1150), .ZN(new_n30138_));
  OAI21_X1   g26909(.A1(new_n30138_), .A2(new_n27251_), .B(new_n28282_), .ZN(new_n30139_));
  OAI21_X1   g26910(.A1(new_n30136_), .A2(new_n30139_), .B(pi1149), .ZN(new_n30140_));
  AOI21_X1   g26911(.A1(new_n30011_), .A2(new_n27251_), .B(pi1150), .ZN(new_n30141_));
  MUX2_X1    g26912(.I0(new_n29882_), .I1(new_n29838_), .S(new_n27251_), .Z(new_n30142_));
  AOI22_X1   g26913(.A1(new_n29877_), .A2(new_n30141_), .B1(pi1150), .B2(new_n30142_), .ZN(new_n30143_));
  NOR2_X1    g26914(.A1(new_n30143_), .A2(pi0275), .ZN(new_n30144_));
  AOI21_X1   g26915(.A1(new_n30140_), .A2(new_n30144_), .B(new_n30133_), .ZN(new_n30145_));
  OAI21_X1   g26916(.A1(new_n30120_), .A2(new_n2918_), .B(new_n28282_), .ZN(new_n30146_));
  NOR4_X1    g26917(.A1(new_n30030_), .A2(pi1149), .A3(new_n27817_), .A4(pi1151), .ZN(new_n30147_));
  OAI21_X1   g26918(.A1(new_n30004_), .A2(pi1149), .B(new_n27251_), .ZN(new_n30148_));
  AOI21_X1   g26919(.A1(new_n30115_), .A2(new_n30148_), .B(new_n27817_), .ZN(new_n30149_));
  NAND4_X1   g26920(.A1(new_n29982_), .A2(new_n29798_), .A3(new_n27470_), .A4(new_n27251_), .ZN(new_n30150_));
  NAND3_X1   g26921(.A1(new_n29050_), .A2(new_n27470_), .A3(pi1151), .ZN(new_n30151_));
  AOI21_X1   g26922(.A1(new_n30150_), .A2(new_n30151_), .B(pi1150), .ZN(new_n30152_));
  NOR3_X1    g26923(.A1(new_n30149_), .A2(new_n2918_), .A3(new_n30152_), .ZN(new_n30153_));
  OAI21_X1   g26924(.A1(new_n30153_), .A2(new_n30147_), .B(pi0275), .ZN(new_n30154_));
  NAND3_X1   g26925(.A1(new_n30146_), .A2(new_n30133_), .A3(new_n30154_), .ZN(new_n30155_));
  AOI21_X1   g26926(.A1(new_n30145_), .A2(new_n30132_), .B(new_n30155_), .ZN(new_n30156_));
  OAI21_X1   g26927(.A1(new_n30156_), .A2(pi0230), .B(new_n30121_), .ZN(po0432));
  INV_X1     g26928(.I(new_n27714_), .ZN(new_n30158_));
  OAI21_X1   g26929(.A1(pi0199), .A2(pi1144), .B(pi1146), .ZN(new_n30159_));
  NAND3_X1   g26930(.A1(new_n8094_), .A2(new_n3258_), .A3(pi1144), .ZN(new_n30160_));
  NAND4_X1   g26931(.A1(new_n30158_), .A2(new_n8098_), .A3(new_n30159_), .A4(new_n30160_), .ZN(new_n30161_));
  NOR3_X1    g26932(.A1(new_n27783_), .A2(pi0230), .A3(new_n30161_), .ZN(new_n30162_));
  NOR2_X1    g26933(.A1(new_n28111_), .A2(new_n28097_), .ZN(new_n30163_));
  XOR2_X1    g26934(.A1(new_n30163_), .A2(new_n3272_), .Z(new_n30164_));
  NOR3_X1    g26935(.A1(new_n27475_), .A2(new_n2918_), .A3(new_n26312_), .ZN(new_n30165_));
  MUX2_X1    g26936(.I0(pi1144), .I1(pi1145), .S(pi0200), .Z(new_n30166_));
  NAND2_X1   g26937(.A1(new_n30166_), .A2(pi1091), .ZN(new_n30167_));
  OAI22_X1   g26938(.A1(new_n29942_), .A2(new_n30167_), .B1(new_n27615_), .B2(new_n30165_), .ZN(new_n30168_));
  OAI21_X1   g26939(.A1(pi1091), .A2(new_n30164_), .B(new_n30168_), .ZN(new_n30169_));
  NOR3_X1    g26940(.A1(new_n28102_), .A2(pi0276), .A3(new_n28097_), .ZN(new_n30170_));
  AOI21_X1   g26941(.A1(new_n28101_), .A2(pi0802), .B(new_n3272_), .ZN(new_n30171_));
  OAI21_X1   g26942(.A1(new_n30170_), .A2(new_n30171_), .B(new_n2918_), .ZN(new_n30172_));
  NAND4_X1   g26943(.A1(new_n11749_), .A2(new_n8094_), .A3(pi1146), .A4(new_n29601_), .ZN(new_n30173_));
  NAND2_X1   g26944(.A1(new_n29902_), .A2(new_n29970_), .ZN(new_n30174_));
  NAND2_X1   g26945(.A1(new_n30174_), .A2(new_n30173_), .ZN(new_n30175_));
  AOI21_X1   g26946(.A1(new_n30175_), .A2(new_n30172_), .B(pi0230), .ZN(new_n30176_));
  AOI21_X1   g26947(.A1(new_n30169_), .A2(new_n30176_), .B(new_n30162_), .ZN(po0433));
  OAI21_X1   g26948(.A1(pi0211), .A2(pi1140), .B(pi1141), .ZN(new_n30178_));
  NAND3_X1   g26949(.A1(new_n8077_), .A2(new_n3831_), .A3(pi1140), .ZN(new_n30179_));
  NAND2_X1   g26950(.A1(new_n9658_), .A2(pi1142), .ZN(new_n30180_));
  NAND4_X1   g26951(.A1(new_n30180_), .A2(new_n30179_), .A3(new_n8247_), .A4(new_n30178_), .ZN(new_n30181_));
  INV_X1     g26952(.I(new_n29931_), .ZN(new_n30182_));
  NOR2_X1    g26953(.A1(new_n3831_), .A2(pi0199), .ZN(new_n30183_));
  OAI22_X1   g26954(.A1(new_n30182_), .A2(new_n26323_), .B1(new_n8098_), .B2(new_n30183_), .ZN(new_n30184_));
  MUX2_X1    g26955(.I0(new_n30181_), .I1(new_n30184_), .S(new_n11749_), .Z(new_n30185_));
  NAND2_X1   g26956(.A1(new_n30185_), .A2(pi0230), .ZN(new_n30186_));
  NAND3_X1   g26957(.A1(new_n28111_), .A2(pi0277), .A3(pi0820), .ZN(new_n30187_));
  INV_X1     g26958(.I(pi0820), .ZN(new_n30188_));
  OAI21_X1   g26959(.A1(new_n29584_), .A2(pi0277), .B(new_n30188_), .ZN(new_n30189_));
  NAND3_X1   g26960(.A1(new_n30189_), .A2(new_n2918_), .A3(new_n30187_), .ZN(new_n30190_));
  AOI21_X1   g26961(.A1(pi1091), .A2(pi1140), .B(new_n30190_), .ZN(new_n30191_));
  AOI21_X1   g26962(.A1(pi1091), .A2(pi1141), .B(new_n30190_), .ZN(new_n30192_));
  XNOR2_X1   g26963(.A1(new_n30191_), .A2(new_n30192_), .ZN(new_n30193_));
  NOR2_X1    g26964(.A1(new_n30193_), .A2(new_n8077_), .ZN(new_n30194_));
  XNOR2_X1   g26965(.A1(new_n30194_), .A2(new_n30191_), .ZN(new_n30195_));
  OAI21_X1   g26966(.A1(new_n30195_), .A2(pi0219), .B(new_n27783_), .ZN(new_n30196_));
  NOR3_X1    g26967(.A1(new_n29077_), .A2(pi0219), .A3(new_n3700_), .ZN(new_n30197_));
  INV_X1     g26968(.I(pi0277), .ZN(new_n30198_));
  NOR3_X1    g26969(.A1(new_n28101_), .A2(new_n30198_), .A3(new_n30188_), .ZN(new_n30199_));
  AOI21_X1   g26970(.A1(new_n28102_), .A2(new_n30198_), .B(pi0820), .ZN(new_n30200_));
  NOR4_X1    g26971(.A1(new_n30200_), .A2(pi1091), .A3(new_n30197_), .A4(new_n30199_), .ZN(new_n30201_));
  MUX2_X1    g26972(.I0(new_n30192_), .I1(new_n30191_), .S(new_n8098_), .Z(new_n30202_));
  NAND2_X1   g26973(.A1(new_n30202_), .A2(new_n8094_), .ZN(new_n30203_));
  NOR3_X1    g26974(.A1(new_n30200_), .A2(pi1091), .A3(new_n30199_), .ZN(new_n30204_));
  NOR2_X1    g26975(.A1(new_n26330_), .A2(new_n29602_), .ZN(new_n30205_));
  NOR3_X1    g26976(.A1(new_n11749_), .A2(new_n30204_), .A3(new_n30205_), .ZN(new_n30206_));
  AOI22_X1   g26977(.A1(new_n30196_), .A2(new_n30201_), .B1(new_n30203_), .B2(new_n30206_), .ZN(new_n30207_));
  OAI21_X1   g26978(.A1(new_n30207_), .A2(pi0230), .B(new_n30186_), .ZN(po0434));
  INV_X1     g26979(.I(pi1132), .ZN(new_n30209_));
  INV_X1     g26980(.I(pi0278), .ZN(po1130));
  INV_X1     g26981(.I(pi0976), .ZN(new_n30211_));
  AOI21_X1   g26982(.A1(new_n28111_), .A2(po1130), .B(new_n30211_), .ZN(new_n30212_));
  NOR3_X1    g26983(.A1(new_n29584_), .A2(po1130), .A3(pi0976), .ZN(new_n30213_));
  NOR3_X1    g26984(.A1(new_n30213_), .A2(pi1091), .A3(new_n30212_), .ZN(new_n30214_));
  INV_X1     g26985(.I(new_n30214_), .ZN(new_n30215_));
  AOI21_X1   g26986(.A1(pi1091), .A2(new_n30209_), .B(new_n30215_), .ZN(new_n30216_));
  NOR2_X1    g26987(.A1(new_n28101_), .A2(pi0278), .ZN(new_n30217_));
  OAI21_X1   g26988(.A1(new_n28102_), .A2(pi0976), .B(new_n2918_), .ZN(new_n30218_));
  NOR3_X1    g26989(.A1(new_n30218_), .A2(new_n8094_), .A3(new_n30217_), .ZN(new_n30219_));
  NOR2_X1    g26990(.A1(new_n30219_), .A2(pi0200), .ZN(new_n30220_));
  OAI21_X1   g26991(.A1(new_n30216_), .A2(new_n8094_), .B(new_n30220_), .ZN(new_n30221_));
  INV_X1     g26992(.I(new_n30219_), .ZN(new_n30222_));
  NOR2_X1    g26993(.A1(new_n2918_), .A2(pi1133), .ZN(new_n30223_));
  NOR4_X1    g26994(.A1(new_n30215_), .A2(pi0199), .A3(new_n30222_), .A4(new_n30223_), .ZN(new_n30224_));
  OAI21_X1   g26995(.A1(new_n30224_), .A2(new_n8098_), .B(new_n2587_), .ZN(new_n30225_));
  OAI21_X1   g26996(.A1(new_n30221_), .A2(new_n30225_), .B(new_n6845_), .ZN(new_n30226_));
  NOR2_X1    g26997(.A1(new_n30209_), .A2(pi0211), .ZN(new_n30227_));
  AOI21_X1   g26998(.A1(pi0211), .A2(pi1133), .B(new_n30227_), .ZN(new_n30228_));
  NOR3_X1    g26999(.A1(new_n6845_), .A2(pi0219), .A3(new_n30228_), .ZN(new_n30229_));
  AOI21_X1   g27000(.A1(new_n8160_), .A2(pi1133), .B(pi0299), .ZN(new_n30230_));
  AOI21_X1   g27001(.A1(new_n8094_), .A2(pi1132), .B(pi0200), .ZN(new_n30231_));
  OAI22_X1   g27002(.A1(new_n30228_), .A2(new_n26998_), .B1(new_n30230_), .B2(new_n30231_), .ZN(new_n30232_));
  NAND3_X1   g27003(.A1(new_n6845_), .A2(new_n30232_), .A3(new_n26307_), .ZN(new_n30233_));
  OAI21_X1   g27004(.A1(new_n30229_), .A2(new_n30233_), .B(new_n29634_), .ZN(new_n30234_));
  AOI21_X1   g27005(.A1(new_n30226_), .A2(new_n26307_), .B(new_n30234_), .ZN(new_n30235_));
  INV_X1     g27006(.I(new_n30225_), .ZN(new_n30236_));
  NAND4_X1   g27007(.A1(new_n30216_), .A2(pi0199), .A3(pi1091), .A4(new_n30220_), .ZN(new_n30237_));
  AOI21_X1   g27008(.A1(pi0299), .A2(new_n30076_), .B(po1038), .ZN(new_n30238_));
  OAI21_X1   g27009(.A1(new_n30236_), .A2(new_n30237_), .B(new_n30238_), .ZN(new_n30239_));
  AOI21_X1   g27010(.A1(po1038), .A2(new_n30076_), .B(pi0230), .ZN(new_n30240_));
  OAI21_X1   g27011(.A1(pi0219), .A2(pi1132), .B(new_n8077_), .ZN(new_n30241_));
  OR3_X2     g27012(.A1(new_n30228_), .A2(new_n8077_), .A3(pi0219), .Z(new_n30242_));
  AOI21_X1   g27013(.A1(new_n30242_), .A2(new_n30241_), .B(new_n6845_), .ZN(new_n30243_));
  AOI21_X1   g27014(.A1(new_n30209_), .A2(new_n8160_), .B(new_n30230_), .ZN(new_n30244_));
  OAI22_X1   g27015(.A1(new_n30228_), .A2(new_n26998_), .B1(new_n2587_), .B2(new_n29048_), .ZN(new_n30245_));
  NOR3_X1    g27016(.A1(po1038), .A2(new_n30244_), .A3(new_n30245_), .ZN(new_n30246_));
  NOR3_X1    g27017(.A1(new_n30246_), .A2(new_n26307_), .A3(new_n30243_), .ZN(new_n30247_));
  AOI21_X1   g27018(.A1(new_n30239_), .A2(new_n30240_), .B(new_n30247_), .ZN(new_n30248_));
  NOR2_X1    g27019(.A1(new_n30248_), .A2(new_n29634_), .ZN(new_n30249_));
  XNOR2_X1   g27020(.A1(new_n30249_), .A2(new_n30235_), .ZN(po0435));
  OAI21_X1   g27021(.A1(pi0199), .A2(pi1135), .B(pi1137), .ZN(new_n30252_));
  NAND3_X1   g27022(.A1(new_n8094_), .A2(new_n4402_), .A3(pi1135), .ZN(new_n30253_));
  AOI21_X1   g27023(.A1(new_n8094_), .A2(pi1136), .B(pi0200), .ZN(new_n30254_));
  NAND3_X1   g27024(.A1(new_n30253_), .A2(new_n30254_), .A3(new_n30252_), .ZN(new_n30255_));
  AND3_X2    g27025(.A1(new_n11749_), .A2(new_n26307_), .A3(new_n30255_), .Z(new_n30256_));
  INV_X1     g27026(.I(pi0914), .ZN(new_n30257_));
  INV_X1     g27027(.I(pi0280), .ZN(new_n30258_));
  AOI21_X1   g27028(.A1(new_n28111_), .A2(new_n30258_), .B(pi1091), .ZN(new_n30259_));
  NOR3_X1    g27029(.A1(new_n30259_), .A2(new_n30257_), .A3(new_n28111_), .ZN(new_n30260_));
  INV_X1     g27030(.I(new_n30260_), .ZN(new_n30261_));
  NOR2_X1    g27031(.A1(pi0211), .A2(pi1135), .ZN(new_n30262_));
  OAI21_X1   g27032(.A1(new_n29659_), .A2(new_n30262_), .B(pi1091), .ZN(new_n30263_));
  NAND2_X1   g27033(.A1(new_n30261_), .A2(new_n30263_), .ZN(new_n30264_));
  NAND3_X1   g27034(.A1(new_n29076_), .A2(new_n8247_), .A3(pi1137), .ZN(new_n30265_));
  NOR3_X1    g27035(.A1(new_n28101_), .A2(new_n30258_), .A3(new_n30257_), .ZN(new_n30266_));
  AOI21_X1   g27036(.A1(new_n28102_), .A2(new_n30258_), .B(pi0914), .ZN(new_n30267_));
  NOR3_X1    g27037(.A1(new_n30267_), .A2(pi1091), .A3(new_n30266_), .ZN(new_n30268_));
  AOI22_X1   g27038(.A1(new_n30264_), .A2(new_n8247_), .B1(new_n30265_), .B2(new_n30268_), .ZN(new_n30269_));
  OAI21_X1   g27039(.A1(new_n4402_), .A2(new_n29602_), .B(new_n30268_), .ZN(new_n30270_));
  NOR2_X1    g27040(.A1(pi0200), .A2(pi1135), .ZN(new_n30271_));
  INV_X1     g27041(.I(new_n30271_), .ZN(new_n30272_));
  AOI21_X1   g27042(.A1(new_n4543_), .A2(pi0200), .B(pi1091), .ZN(new_n30273_));
  AOI21_X1   g27043(.A1(new_n30273_), .A2(new_n30272_), .B(pi0199), .ZN(new_n30274_));
  AOI22_X1   g27044(.A1(new_n30270_), .A2(pi0199), .B1(new_n30261_), .B2(new_n30274_), .ZN(new_n30275_));
  INV_X1     g27045(.I(new_n30275_), .ZN(new_n30276_));
  OAI21_X1   g27046(.A1(new_n30276_), .A2(new_n27783_), .B(new_n30269_), .ZN(new_n30277_));
  NOR3_X1    g27047(.A1(new_n30269_), .A2(new_n27783_), .A3(new_n30275_), .ZN(new_n30278_));
  NOR2_X1    g27048(.A1(new_n30278_), .A2(pi0230), .ZN(new_n30279_));
  AOI21_X1   g27049(.A1(new_n30279_), .A2(new_n30277_), .B(new_n30256_), .ZN(po0437));
  NOR3_X1    g27050(.A1(new_n29902_), .A2(new_n4115_), .A3(new_n29077_), .ZN(new_n30281_));
  AOI21_X1   g27051(.A1(pi1139), .A2(new_n29601_), .B(new_n29904_), .ZN(new_n30282_));
  INV_X1     g27052(.I(pi0830), .ZN(new_n30283_));
  NOR3_X1    g27053(.A1(new_n28101_), .A2(new_n4119_), .A3(new_n30283_), .ZN(new_n30284_));
  OAI21_X1   g27054(.A1(new_n28101_), .A2(pi0281), .B(new_n30283_), .ZN(new_n30285_));
  NAND2_X1   g27055(.A1(new_n30285_), .A2(new_n2918_), .ZN(new_n30286_));
  NOR4_X1    g27056(.A1(new_n30282_), .A2(new_n30281_), .A3(new_n30284_), .A4(new_n30286_), .ZN(new_n30287_));
  NOR2_X1    g27057(.A1(new_n8077_), .A2(pi1138), .ZN(new_n30288_));
  NOR2_X1    g27058(.A1(pi0211), .A2(pi1137), .ZN(new_n30289_));
  NOR3_X1    g27059(.A1(new_n30288_), .A2(new_n2918_), .A3(new_n30289_), .ZN(new_n30290_));
  NOR2_X1    g27060(.A1(new_n27615_), .A2(new_n30290_), .ZN(new_n30291_));
  NAND3_X1   g27061(.A1(new_n4402_), .A2(pi0200), .A3(pi1138), .ZN(new_n30292_));
  OAI21_X1   g27062(.A1(new_n8098_), .A2(pi1138), .B(pi1137), .ZN(new_n30293_));
  AOI21_X1   g27063(.A1(new_n30293_), .A2(new_n30292_), .B(new_n2918_), .ZN(new_n30294_));
  NAND2_X1   g27064(.A1(new_n29801_), .A2(new_n30294_), .ZN(new_n30295_));
  NAND3_X1   g27065(.A1(new_n28111_), .A2(pi0281), .A3(pi0830), .ZN(new_n30296_));
  OAI21_X1   g27066(.A1(new_n29584_), .A2(pi0281), .B(new_n30283_), .ZN(new_n30297_));
  NAND4_X1   g27067(.A1(new_n30295_), .A2(new_n2918_), .A3(new_n30296_), .A4(new_n30297_), .ZN(new_n30298_));
  OAI21_X1   g27068(.A1(new_n30298_), .A2(new_n30291_), .B(new_n26307_), .ZN(new_n30299_));
  OAI21_X1   g27069(.A1(pi0199), .A2(pi1137), .B(pi1139), .ZN(new_n30300_));
  NAND3_X1   g27070(.A1(new_n8094_), .A2(new_n4115_), .A3(pi1137), .ZN(new_n30301_));
  NAND2_X1   g27071(.A1(new_n8160_), .A2(pi1138), .ZN(new_n30302_));
  NAND4_X1   g27072(.A1(new_n30302_), .A2(new_n30301_), .A3(new_n8098_), .A4(new_n30300_), .ZN(new_n30303_));
  NOR2_X1    g27073(.A1(new_n27783_), .A2(new_n30303_), .ZN(new_n30304_));
  OAI22_X1   g27074(.A1(new_n30299_), .A2(new_n30287_), .B1(new_n26307_), .B2(new_n30304_), .ZN(po0438));
  NOR2_X1    g27075(.A1(new_n29982_), .A2(new_n27494_), .ZN(new_n30307_));
  NOR3_X1    g27076(.A1(new_n30307_), .A2(new_n27470_), .A3(new_n30004_), .ZN(new_n30308_));
  NOR4_X1    g27077(.A1(new_n29803_), .A2(pi1147), .A3(pi1149), .A4(new_n29793_), .ZN(new_n30309_));
  NOR2_X1    g27078(.A1(new_n30308_), .A2(new_n30309_), .ZN(new_n30310_));
  NAND2_X1   g27079(.A1(new_n29050_), .A2(pi1149), .ZN(new_n30311_));
  NOR2_X1    g27080(.A1(new_n30307_), .A2(pi1148), .ZN(new_n30312_));
  AOI21_X1   g27081(.A1(new_n30312_), .A2(new_n30311_), .B(new_n26307_), .ZN(new_n30313_));
  NOR3_X1    g27082(.A1(new_n30310_), .A2(new_n30313_), .A3(pi1148), .ZN(new_n30314_));
  AOI21_X1   g27083(.A1(new_n27494_), .A2(new_n29851_), .B(new_n29876_), .ZN(new_n30315_));
  NAND3_X1   g27084(.A1(new_n29876_), .A2(new_n27494_), .A3(new_n30122_), .ZN(new_n30316_));
  NAND4_X1   g27085(.A1(new_n29848_), .A2(pi1147), .A3(new_n27515_), .A4(new_n29881_), .ZN(new_n30317_));
  NAND3_X1   g27086(.A1(new_n30316_), .A2(new_n27515_), .A3(new_n30317_), .ZN(new_n30318_));
  NOR2_X1    g27087(.A1(new_n29839_), .A2(pi1147), .ZN(new_n30319_));
  NOR2_X1    g27088(.A1(new_n30319_), .A2(pi1148), .ZN(new_n30320_));
  NAND2_X1   g27089(.A1(new_n29867_), .A2(pi1147), .ZN(new_n30321_));
  NOR3_X1    g27090(.A1(new_n29838_), .A2(new_n27494_), .A3(pi1148), .ZN(new_n30322_));
  AOI21_X1   g27091(.A1(new_n29842_), .A2(new_n30322_), .B(pi1149), .ZN(new_n30323_));
  OAI21_X1   g27092(.A1(new_n30321_), .A2(new_n30320_), .B(new_n30323_), .ZN(new_n30324_));
  AOI21_X1   g27093(.A1(new_n30324_), .A2(pi0283), .B(pi1149), .ZN(new_n30325_));
  OAI21_X1   g27094(.A1(new_n30318_), .A2(new_n30315_), .B(new_n30325_), .ZN(new_n30326_));
  NOR4_X1    g27095(.A1(new_n29993_), .A2(new_n27494_), .A3(pi1149), .A4(new_n29889_), .ZN(new_n30327_));
  AOI21_X1   g27096(.A1(new_n29830_), .A2(new_n27494_), .B(pi1149), .ZN(new_n30328_));
  NOR3_X1    g27097(.A1(new_n30328_), .A2(new_n27494_), .A3(new_n30000_), .ZN(new_n30329_));
  OAI21_X1   g27098(.A1(new_n30329_), .A2(new_n30327_), .B(new_n27515_), .ZN(new_n30330_));
  NAND4_X1   g27099(.A1(new_n30137_), .A2(pi1147), .A3(new_n27470_), .A4(new_n29811_), .ZN(new_n30331_));
  NOR2_X1    g27100(.A1(new_n27494_), .A2(new_n27470_), .ZN(new_n30332_));
  AOI21_X1   g27101(.A1(new_n29864_), .A2(new_n30332_), .B(pi1148), .ZN(new_n30333_));
  AOI22_X1   g27102(.A1(new_n30330_), .A2(new_n28283_), .B1(new_n30331_), .B2(new_n30333_), .ZN(new_n30334_));
  NOR2_X1    g27103(.A1(new_n30334_), .A2(pi0230), .ZN(new_n30335_));
  AOI21_X1   g27104(.A1(new_n30335_), .A2(new_n30326_), .B(new_n30314_), .ZN(po0440));
  INV_X1     g27105(.I(pi0285), .ZN(new_n30338_));
  INV_X1     g27106(.I(pi0289), .ZN(new_n30339_));
  INV_X1     g27107(.I(pi0286), .ZN(new_n30340_));
  NAND2_X1   g27108(.A1(new_n8005_), .A2(new_n3233_), .ZN(new_n30341_));
  NOR2_X1    g27109(.A1(new_n30341_), .A2(new_n6428_), .ZN(new_n30342_));
  INV_X1     g27110(.I(new_n30342_), .ZN(new_n30343_));
  NOR2_X1    g27111(.A1(new_n30343_), .A2(new_n30340_), .ZN(new_n30344_));
  INV_X1     g27112(.I(new_n30344_), .ZN(new_n30345_));
  NOR3_X1    g27113(.A1(new_n30345_), .A2(new_n6536_), .A3(new_n30339_), .ZN(new_n30346_));
  NOR3_X1    g27114(.A1(new_n6429_), .A2(pi0286), .A3(pi0288), .ZN(new_n30347_));
  NAND2_X1   g27115(.A1(new_n30347_), .A2(new_n30339_), .ZN(new_n30348_));
  NAND4_X1   g27116(.A1(new_n30346_), .A2(new_n30338_), .A3(new_n6845_), .A4(new_n30348_), .ZN(new_n30349_));
  INV_X1     g27117(.I(new_n30341_), .ZN(new_n30350_));
  OAI21_X1   g27118(.A1(new_n30346_), .A2(new_n30350_), .B(pi0285), .ZN(new_n30351_));
  XNOR2_X1   g27119(.A1(new_n30351_), .A2(new_n30346_), .ZN(new_n30352_));
  NAND2_X1   g27120(.A1(new_n30352_), .A2(new_n6845_), .ZN(new_n30353_));
  AOI21_X1   g27121(.A1(new_n30353_), .A2(new_n30349_), .B(pi0793), .ZN(po0442));
  NOR2_X1    g27122(.A1(new_n30343_), .A2(pi0286), .ZN(new_n30355_));
  NOR2_X1    g27123(.A1(new_n30342_), .A2(new_n30340_), .ZN(new_n30356_));
  OAI21_X1   g27124(.A1(new_n30355_), .A2(new_n30356_), .B(pi0288), .ZN(new_n30357_));
  NOR2_X1    g27125(.A1(new_n6537_), .A2(pi0288), .ZN(new_n30358_));
  NAND2_X1   g27126(.A1(new_n30341_), .A2(new_n6428_), .ZN(new_n30359_));
  XOR2_X1    g27127(.A1(new_n30359_), .A2(new_n30340_), .Z(new_n30360_));
  AOI21_X1   g27128(.A1(new_n30360_), .A2(new_n30358_), .B(po1038), .ZN(new_n30361_));
  INV_X1     g27129(.I(pi0793), .ZN(new_n30362_));
  NAND2_X1   g27130(.A1(new_n6428_), .A2(new_n30358_), .ZN(new_n30363_));
  XOR2_X1    g27131(.A1(new_n30363_), .A2(pi0286), .Z(new_n30364_));
  OAI21_X1   g27132(.A1(new_n30364_), .A2(po1038), .B(new_n30362_), .ZN(new_n30365_));
  AOI21_X1   g27133(.A1(new_n30361_), .A2(new_n30357_), .B(new_n30365_), .ZN(po0443));
  AOI21_X1   g27134(.A1(new_n8018_), .A2(pi0457), .B(pi0332), .ZN(po0444));
  NAND2_X1   g27135(.A1(new_n6429_), .A2(new_n6536_), .ZN(new_n30368_));
  OAI21_X1   g27136(.A1(new_n6429_), .A2(new_n30358_), .B(new_n30368_), .ZN(new_n30369_));
  NOR2_X1    g27137(.A1(new_n30341_), .A2(po1038), .ZN(po0637));
  XOR2_X1    g27138(.A1(po0637), .A2(new_n30369_), .Z(new_n30371_));
  NOR2_X1    g27139(.A1(new_n30371_), .A2(pi0793), .ZN(po0445));
  NAND2_X1   g27140(.A1(new_n30345_), .A2(pi0289), .ZN(new_n30373_));
  NAND2_X1   g27141(.A1(new_n30344_), .A2(new_n30339_), .ZN(new_n30374_));
  AOI21_X1   g27142(.A1(new_n30373_), .A2(new_n30374_), .B(pi0288), .ZN(new_n30375_));
  NOR3_X1    g27143(.A1(new_n30350_), .A2(pi0286), .A3(new_n6429_), .ZN(new_n30376_));
  AOI21_X1   g27144(.A1(new_n30376_), .A2(new_n30338_), .B(pi0289), .ZN(new_n30377_));
  AND2_X2    g27145(.A1(new_n30377_), .A2(new_n30376_), .Z(new_n30378_));
  NOR2_X1    g27146(.A1(new_n30377_), .A2(new_n30376_), .ZN(new_n30379_));
  INV_X1     g27147(.I(new_n30347_), .ZN(new_n30380_));
  NAND2_X1   g27148(.A1(new_n30380_), .A2(pi0289), .ZN(new_n30381_));
  OAI21_X1   g27149(.A1(new_n30380_), .A2(pi0285), .B(new_n6845_), .ZN(new_n30382_));
  AOI21_X1   g27150(.A1(new_n30348_), .A2(new_n30381_), .B(new_n30382_), .ZN(new_n30383_));
  NOR2_X1    g27151(.A1(po1038), .A2(pi0288), .ZN(new_n30384_));
  OAI21_X1   g27152(.A1(new_n30383_), .A2(pi0793), .B(new_n30384_), .ZN(new_n30385_));
  NOR4_X1    g27153(.A1(new_n30375_), .A2(new_n30378_), .A3(new_n30379_), .A4(new_n30385_), .ZN(po0446));
  INV_X1     g27154(.I(pi1048), .ZN(new_n30387_));
  NAND2_X1   g27155(.A1(pi0290), .A2(pi0476), .ZN(new_n30388_));
  OAI21_X1   g27156(.A1(pi0476), .A2(new_n30387_), .B(new_n30388_), .ZN(po0447));
  INV_X1     g27157(.I(pi1049), .ZN(new_n30390_));
  NAND2_X1   g27158(.A1(pi0291), .A2(pi0476), .ZN(new_n30391_));
  OAI21_X1   g27159(.A1(pi0476), .A2(new_n30390_), .B(new_n30391_), .ZN(po0448));
  INV_X1     g27160(.I(pi1084), .ZN(new_n30393_));
  NAND2_X1   g27161(.A1(pi0292), .A2(pi0476), .ZN(new_n30394_));
  OAI21_X1   g27162(.A1(pi0476), .A2(new_n30393_), .B(new_n30394_), .ZN(po0449));
  INV_X1     g27163(.I(pi1059), .ZN(new_n30396_));
  NAND2_X1   g27164(.A1(pi0293), .A2(pi0476), .ZN(new_n30397_));
  OAI21_X1   g27165(.A1(pi0476), .A2(new_n30396_), .B(new_n30397_), .ZN(po0450));
  INV_X1     g27166(.I(pi1072), .ZN(new_n30399_));
  NAND2_X1   g27167(.A1(pi0294), .A2(pi0476), .ZN(new_n30400_));
  OAI21_X1   g27168(.A1(pi0476), .A2(new_n30399_), .B(new_n30400_), .ZN(po0451));
  INV_X1     g27169(.I(pi1053), .ZN(new_n30402_));
  NAND2_X1   g27170(.A1(pi0295), .A2(pi0476), .ZN(new_n30403_));
  OAI21_X1   g27171(.A1(pi0476), .A2(new_n30402_), .B(new_n30403_), .ZN(po0452));
  INV_X1     g27172(.I(pi1037), .ZN(new_n30405_));
  NAND2_X1   g27173(.A1(pi0296), .A2(pi0476), .ZN(new_n30406_));
  OAI21_X1   g27174(.A1(pi0476), .A2(new_n30405_), .B(new_n30406_), .ZN(po0453));
  INV_X1     g27175(.I(pi1044), .ZN(new_n30408_));
  NAND2_X1   g27176(.A1(pi0297), .A2(pi0476), .ZN(new_n30409_));
  OAI21_X1   g27177(.A1(pi0476), .A2(new_n30408_), .B(new_n30409_), .ZN(po0454));
  NAND2_X1   g27178(.A1(pi0298), .A2(pi0478), .ZN(new_n30411_));
  OAI21_X1   g27179(.A1(pi0478), .A2(new_n30408_), .B(new_n30411_), .ZN(po0455));
  NAND4_X1   g27180(.A1(new_n9873_), .A2(new_n3214_), .A3(new_n2889_), .A4(new_n8548_), .ZN(new_n30413_));
  NOR2_X1    g27181(.A1(new_n2491_), .A2(new_n3214_), .ZN(new_n30414_));
  NOR2_X1    g27182(.A1(new_n2491_), .A2(new_n3214_), .ZN(new_n30415_));
  NOR4_X1    g27183(.A1(new_n30415_), .A2(new_n3208_), .A3(new_n3228_), .A4(new_n6965_), .ZN(new_n30416_));
  OAI21_X1   g27184(.A1(new_n30413_), .A2(new_n30414_), .B(new_n30416_), .ZN(new_n30417_));
  AOI21_X1   g27185(.A1(new_n30417_), .A2(new_n3154_), .B(new_n8553_), .ZN(po0456));
  INV_X1     g27186(.I(pi0300), .ZN(new_n30419_));
  NOR4_X1    g27187(.A1(new_n7807_), .A2(new_n5055_), .A3(pi0059), .A4(pi0312), .ZN(new_n30420_));
  XOR2_X1    g27188(.A1(new_n30420_), .A2(new_n30419_), .Z(new_n30421_));
  NAND2_X1   g27189(.A1(new_n30421_), .A2(new_n3227_), .ZN(po0457));
  INV_X1     g27190(.I(pi0301), .ZN(new_n30423_));
  NAND2_X1   g27191(.A1(new_n30420_), .A2(new_n30419_), .ZN(new_n30424_));
  NAND2_X1   g27192(.A1(new_n30424_), .A2(new_n30423_), .ZN(new_n30425_));
  NOR2_X1    g27193(.A1(new_n30424_), .A2(new_n30423_), .ZN(new_n30426_));
  INV_X1     g27194(.I(new_n30426_), .ZN(new_n30427_));
  AOI21_X1   g27195(.A1(new_n30427_), .A2(new_n30425_), .B(pi0055), .ZN(po0458));
  NOR2_X1    g27196(.A1(new_n11749_), .A2(new_n3287_), .ZN(new_n30429_));
  INV_X1     g27197(.I(new_n30429_), .ZN(new_n30430_));
  INV_X1     g27198(.I(new_n4989_), .ZN(new_n30431_));
  NOR2_X1    g27199(.A1(po1038), .A2(new_n30431_), .ZN(new_n30432_));
  INV_X1     g27200(.I(new_n30432_), .ZN(new_n30433_));
  NAND2_X1   g27201(.A1(new_n2598_), .A2(pi0937), .ZN(new_n30434_));
  NAND4_X1   g27202(.A1(new_n30433_), .A2(pi0273), .A3(new_n3299_), .A4(new_n30434_), .ZN(new_n30435_));
  AOI21_X1   g27203(.A1(new_n30435_), .A2(new_n30430_), .B(new_n24070_), .ZN(new_n30436_));
  NOR2_X1    g27204(.A1(new_n11749_), .A2(new_n4981_), .ZN(new_n30437_));
  NOR2_X1    g27205(.A1(new_n30437_), .A2(new_n30432_), .ZN(new_n30438_));
  INV_X1     g27206(.I(new_n30438_), .ZN(new_n30439_));
  INV_X1     g27207(.I(pi0937), .ZN(new_n30440_));
  NAND3_X1   g27208(.A1(new_n6452_), .A2(pi0833), .A3(new_n30440_), .ZN(new_n30441_));
  NOR2_X1    g27209(.A1(new_n2531_), .A2(new_n2562_), .ZN(new_n30442_));
  NAND2_X1   g27210(.A1(new_n30442_), .A2(new_n28095_), .ZN(new_n30443_));
  NAND4_X1   g27211(.A1(new_n27783_), .A2(new_n3155_), .A3(new_n30441_), .A4(new_n30443_), .ZN(new_n30444_));
  NOR2_X1    g27212(.A1(new_n30435_), .A2(new_n30444_), .ZN(new_n30445_));
  NOR4_X1    g27213(.A1(new_n30436_), .A2(new_n30445_), .A3(pi1148), .A4(new_n30439_), .ZN(po0459));
  NAND2_X1   g27214(.A1(pi0303), .A2(pi0478), .ZN(new_n30447_));
  OAI21_X1   g27215(.A1(pi0478), .A2(new_n30390_), .B(new_n30447_), .ZN(po0460));
  NAND2_X1   g27216(.A1(pi0304), .A2(pi0478), .ZN(new_n30449_));
  OAI21_X1   g27217(.A1(pi0478), .A2(new_n30387_), .B(new_n30449_), .ZN(po0461));
  NAND2_X1   g27218(.A1(pi0305), .A2(pi0478), .ZN(new_n30451_));
  OAI21_X1   g27219(.A1(pi0478), .A2(new_n30393_), .B(new_n30451_), .ZN(po0462));
  NAND2_X1   g27220(.A1(pi0306), .A2(pi0478), .ZN(new_n30453_));
  OAI21_X1   g27221(.A1(pi0478), .A2(new_n30396_), .B(new_n30453_), .ZN(po0463));
  NAND2_X1   g27222(.A1(pi0307), .A2(pi0478), .ZN(new_n30455_));
  OAI21_X1   g27223(.A1(pi0478), .A2(new_n30402_), .B(new_n30455_), .ZN(po0464));
  NAND2_X1   g27224(.A1(pi0308), .A2(pi0478), .ZN(new_n30457_));
  OAI21_X1   g27225(.A1(pi0478), .A2(new_n30405_), .B(new_n30457_), .ZN(po0465));
  NAND2_X1   g27226(.A1(pi0309), .A2(pi0478), .ZN(new_n30459_));
  OAI21_X1   g27227(.A1(pi0478), .A2(new_n30399_), .B(new_n30459_), .ZN(po0466));
  AOI22_X1   g27228(.A1(new_n2531_), .A2(pi0934), .B1(new_n3278_), .B2(pi0271), .ZN(new_n30461_));
  NOR3_X1    g27229(.A1(new_n11749_), .A2(new_n4981_), .A3(new_n30461_), .ZN(new_n30462_));
  NOR2_X1    g27230(.A1(new_n27783_), .A2(new_n3590_), .ZN(new_n30463_));
  NAND2_X1   g27231(.A1(new_n3299_), .A2(new_n28096_), .ZN(new_n30464_));
  NOR2_X1    g27232(.A1(new_n2588_), .A2(pi0934), .ZN(new_n30465_));
  XOR2_X1    g27233(.A1(new_n30464_), .A2(new_n30465_), .Z(new_n30466_));
  AND2_X2    g27234(.A1(new_n30432_), .A2(new_n30466_), .Z(new_n30467_));
  NOR4_X1    g27235(.A1(new_n30463_), .A2(new_n30467_), .A3(new_n27494_), .A4(new_n30462_), .ZN(new_n30468_));
  AOI22_X1   g27236(.A1(new_n30437_), .A2(new_n3285_), .B1(new_n3155_), .B2(new_n30432_), .ZN(new_n30469_));
  AND3_X2    g27237(.A1(new_n30437_), .A2(new_n3285_), .A3(new_n30461_), .Z(new_n30470_));
  NOR2_X1    g27238(.A1(new_n30433_), .A2(new_n30466_), .ZN(new_n30471_));
  NOR4_X1    g27239(.A1(new_n30470_), .A2(pi1147), .A3(new_n30429_), .A4(new_n30471_), .ZN(new_n30472_));
  AOI21_X1   g27240(.A1(new_n30472_), .A2(new_n30469_), .B(new_n30468_), .ZN(new_n30473_));
  NOR3_X1    g27241(.A1(new_n30470_), .A2(new_n30429_), .A3(new_n30471_), .ZN(new_n30474_));
  NOR2_X1    g27242(.A1(new_n30439_), .A2(new_n27494_), .ZN(new_n30475_));
  OAI21_X1   g27243(.A1(new_n30474_), .A2(new_n30475_), .B(new_n24069_), .ZN(new_n30476_));
  OAI21_X1   g27244(.A1(new_n30473_), .A2(new_n24069_), .B(new_n30476_), .ZN(po0467));
  INV_X1     g27245(.I(pi0311), .ZN(new_n30478_));
  AOI21_X1   g27246(.A1(new_n30426_), .A2(new_n30478_), .B(pi0055), .ZN(new_n30479_));
  OAI21_X1   g27247(.A1(new_n30478_), .A2(new_n30426_), .B(new_n30479_), .ZN(po0468));
  NAND3_X1   g27248(.A1(new_n7806_), .A2(pi0057), .A3(new_n5205_), .ZN(new_n30481_));
  OAI21_X1   g27249(.A1(new_n30481_), .A2(pi0312), .B(new_n3227_), .ZN(new_n30482_));
  AOI21_X1   g27250(.A1(pi0312), .A2(new_n30481_), .B(new_n30482_), .ZN(po0469));
  INV_X1     g27251(.I(pi0313), .ZN(new_n30484_));
  NAND2_X1   g27252(.A1(new_n30484_), .A2(pi0954), .ZN(new_n30485_));
  NAND2_X1   g27253(.A1(new_n9902_), .A2(new_n7990_), .ZN(new_n30486_));
  NAND2_X1   g27254(.A1(new_n9905_), .A2(po0740), .ZN(new_n30487_));
  NAND3_X1   g27255(.A1(new_n30487_), .A2(new_n30486_), .A3(new_n7828_), .ZN(po0634));
  OAI21_X1   g27256(.A1(po0634), .A2(pi0954), .B(new_n30485_), .ZN(po0470));
  NAND2_X1   g27257(.A1(new_n10504_), .A2(new_n2622_), .ZN(new_n30490_));
  OAI21_X1   g27258(.A1(new_n11245_), .A2(new_n10978_), .B(pi0039), .ZN(new_n30491_));
  OAI21_X1   g27259(.A1(new_n30491_), .A2(new_n2622_), .B(new_n30490_), .ZN(new_n30492_));
  NOR2_X1    g27260(.A1(new_n7823_), .A2(new_n2537_), .ZN(new_n30493_));
  OAI21_X1   g27261(.A1(new_n5582_), .A2(new_n6965_), .B(new_n10506_), .ZN(new_n30494_));
  NAND3_X1   g27262(.A1(new_n30494_), .A2(new_n10499_), .A3(new_n10501_), .ZN(new_n30495_));
  AOI21_X1   g27263(.A1(new_n30492_), .A2(new_n30493_), .B(new_n30495_), .ZN(po0471));
  INV_X1     g27264(.I(pi1080), .ZN(new_n30497_));
  INV_X1     g27265(.I(pi0340), .ZN(new_n30498_));
  NAND3_X1   g27266(.A1(new_n30350_), .A2(new_n30498_), .A3(new_n6845_), .ZN(new_n30499_));
  NAND2_X1   g27267(.A1(new_n30499_), .A2(pi0315), .ZN(new_n30500_));
  OAI21_X1   g27268(.A1(new_n30497_), .A2(new_n30499_), .B(new_n30500_), .ZN(po0472));
  INV_X1     g27269(.I(pi1047), .ZN(new_n30502_));
  NAND2_X1   g27270(.A1(new_n30499_), .A2(pi0316), .ZN(new_n30503_));
  OAI21_X1   g27271(.A1(new_n30502_), .A2(new_n30499_), .B(new_n30503_), .ZN(po0473));
  INV_X1     g27272(.I(po0637), .ZN(new_n30505_));
  NOR2_X1    g27273(.A1(new_n30505_), .A2(pi0330), .ZN(new_n30506_));
  NAND2_X1   g27274(.A1(new_n30506_), .A2(pi1078), .ZN(new_n30507_));
  OAI21_X1   g27275(.A1(new_n6356_), .A2(new_n30506_), .B(new_n30507_), .ZN(po0474));
  INV_X1     g27276(.I(pi1074), .ZN(new_n30509_));
  INV_X1     g27277(.I(pi0341), .ZN(new_n30510_));
  NAND3_X1   g27278(.A1(new_n30350_), .A2(new_n30510_), .A3(new_n6845_), .ZN(new_n30511_));
  NAND2_X1   g27279(.A1(new_n30511_), .A2(pi0318), .ZN(new_n30512_));
  OAI21_X1   g27280(.A1(new_n30509_), .A2(new_n30511_), .B(new_n30512_), .ZN(po0475));
  NAND2_X1   g27281(.A1(new_n30511_), .A2(pi0319), .ZN(new_n30514_));
  OAI21_X1   g27282(.A1(new_n30399_), .A2(new_n30511_), .B(new_n30514_), .ZN(po0476));
  NAND2_X1   g27283(.A1(new_n30499_), .A2(pi0320), .ZN(new_n30516_));
  OAI21_X1   g27284(.A1(new_n30387_), .A2(new_n30499_), .B(new_n30516_), .ZN(po0477));
  INV_X1     g27285(.I(pi1058), .ZN(new_n30518_));
  NAND2_X1   g27286(.A1(new_n30499_), .A2(pi0321), .ZN(new_n30519_));
  OAI21_X1   g27287(.A1(new_n30518_), .A2(new_n30499_), .B(new_n30519_), .ZN(po0478));
  INV_X1     g27288(.I(pi1051), .ZN(new_n30521_));
  NAND2_X1   g27289(.A1(new_n30499_), .A2(pi0322), .ZN(new_n30522_));
  OAI21_X1   g27290(.A1(new_n30521_), .A2(new_n30499_), .B(new_n30522_), .ZN(po0479));
  NAND2_X1   g27291(.A1(new_n30499_), .A2(pi0323), .ZN(new_n30524_));
  OAI21_X1   g27292(.A1(new_n29385_), .A2(new_n30499_), .B(new_n30524_), .ZN(po0480));
  INV_X1     g27293(.I(pi1086), .ZN(new_n30526_));
  NAND2_X1   g27294(.A1(new_n30511_), .A2(pi0324), .ZN(new_n30527_));
  OAI21_X1   g27295(.A1(new_n30526_), .A2(new_n30511_), .B(new_n30527_), .ZN(po0481));
  INV_X1     g27296(.I(pi1063), .ZN(new_n30529_));
  NAND2_X1   g27297(.A1(new_n30511_), .A2(pi0325), .ZN(new_n30530_));
  OAI21_X1   g27298(.A1(new_n30529_), .A2(new_n30511_), .B(new_n30530_), .ZN(po0482));
  INV_X1     g27299(.I(pi1057), .ZN(new_n30532_));
  NAND2_X1   g27300(.A1(new_n30511_), .A2(pi0326), .ZN(new_n30533_));
  OAI21_X1   g27301(.A1(new_n30532_), .A2(new_n30511_), .B(new_n30533_), .ZN(po0483));
  NAND2_X1   g27302(.A1(new_n30499_), .A2(pi0327), .ZN(new_n30535_));
  OAI21_X1   g27303(.A1(new_n29410_), .A2(new_n30499_), .B(new_n30535_), .ZN(po0484));
  NAND2_X1   g27304(.A1(new_n30511_), .A2(pi0328), .ZN(new_n30537_));
  OAI21_X1   g27305(.A1(new_n30518_), .A2(new_n30511_), .B(new_n30537_), .ZN(po0485));
  INV_X1     g27306(.I(pi1043), .ZN(new_n30539_));
  NAND2_X1   g27307(.A1(new_n30511_), .A2(pi0329), .ZN(new_n30540_));
  OAI21_X1   g27308(.A1(new_n30539_), .A2(new_n30511_), .B(new_n30540_), .ZN(po0486));
  NAND2_X1   g27309(.A1(new_n30341_), .A2(pi0330), .ZN(new_n30542_));
  NOR2_X1    g27310(.A1(new_n2959_), .A2(new_n2923_), .ZN(new_n30543_));
  NOR3_X1    g27311(.A1(new_n6845_), .A2(pi0330), .A3(new_n30543_), .ZN(new_n30544_));
  NAND2_X1   g27312(.A1(new_n30542_), .A2(new_n30544_), .ZN(new_n30545_));
  AOI21_X1   g27313(.A1(pi0340), .A2(new_n30350_), .B(new_n30545_), .ZN(po0487));
  NOR2_X1    g27314(.A1(new_n30341_), .A2(new_n30510_), .ZN(new_n30547_));
  INV_X1     g27315(.I(pi0331), .ZN(new_n30548_));
  NOR2_X1    g27316(.A1(new_n30350_), .A2(new_n30548_), .ZN(new_n30549_));
  INV_X1     g27317(.I(new_n30543_), .ZN(new_n30550_));
  NAND3_X1   g27318(.A1(po1038), .A2(new_n30548_), .A3(new_n30550_), .ZN(new_n30551_));
  NOR3_X1    g27319(.A1(new_n30549_), .A2(new_n30547_), .A3(new_n30551_), .ZN(po0488));
  NOR3_X1    g27320(.A1(new_n8164_), .A2(new_n3172_), .A3(new_n3154_), .ZN(new_n30557_));
  NOR4_X1    g27321(.A1(new_n5154_), .A2(pi0038), .A3(new_n30557_), .A4(new_n7832_), .ZN(po0489));
  NAND2_X1   g27322(.A1(new_n30511_), .A2(pi0333), .ZN(new_n30559_));
  OAI21_X1   g27323(.A1(new_n29410_), .A2(new_n30511_), .B(new_n30559_), .ZN(po0490));
  NAND2_X1   g27324(.A1(new_n30511_), .A2(pi0334), .ZN(new_n30561_));
  OAI21_X1   g27325(.A1(new_n29385_), .A2(new_n30511_), .B(new_n30561_), .ZN(po0491));
  NAND2_X1   g27326(.A1(new_n30511_), .A2(pi0335), .ZN(new_n30563_));
  OAI21_X1   g27327(.A1(new_n29397_), .A2(new_n30511_), .B(new_n30563_), .ZN(po0492));
  INV_X1     g27328(.I(pi0336), .ZN(new_n30565_));
  NAND2_X1   g27329(.A1(new_n30506_), .A2(pi1070), .ZN(new_n30566_));
  OAI21_X1   g27330(.A1(new_n30565_), .A2(new_n30506_), .B(new_n30566_), .ZN(po0493));
  INV_X1     g27331(.I(new_n30506_), .ZN(new_n30568_));
  NAND2_X1   g27332(.A1(new_n30568_), .A2(pi0337), .ZN(new_n30569_));
  OAI21_X1   g27333(.A1(new_n30408_), .A2(new_n30568_), .B(new_n30569_), .ZN(po0494));
  INV_X1     g27334(.I(pi0338), .ZN(new_n30571_));
  NAND2_X1   g27335(.A1(new_n30506_), .A2(pi1072), .ZN(new_n30572_));
  OAI21_X1   g27336(.A1(new_n30571_), .A2(new_n30506_), .B(new_n30572_), .ZN(po0495));
  NAND2_X1   g27337(.A1(new_n30568_), .A2(pi0339), .ZN(new_n30574_));
  OAI21_X1   g27338(.A1(new_n30526_), .A2(new_n30568_), .B(new_n30574_), .ZN(po0496));
  MUX2_X1    g27339(.I0(new_n30548_), .I1(new_n30498_), .S(new_n30341_), .Z(new_n30576_));
  NAND2_X1   g27340(.A1(new_n6845_), .A2(new_n30543_), .ZN(new_n30577_));
  NAND2_X1   g27341(.A1(new_n30543_), .A2(pi0340), .ZN(new_n30578_));
  OAI22_X1   g27342(.A1(new_n30576_), .A2(new_n30577_), .B1(new_n6845_), .B2(new_n30578_), .ZN(po0497));
  NOR2_X1    g27343(.A1(po0637), .A2(pi0341), .ZN(new_n30580_));
  NOR3_X1    g27344(.A1(new_n30506_), .A2(new_n30543_), .A3(new_n30580_), .ZN(po0498));
  NAND2_X1   g27345(.A1(new_n30499_), .A2(pi0342), .ZN(new_n30582_));
  OAI21_X1   g27346(.A1(new_n30390_), .A2(new_n30499_), .B(new_n30582_), .ZN(po0499));
  NAND2_X1   g27347(.A1(new_n30499_), .A2(pi0343), .ZN(new_n30584_));
  OAI21_X1   g27348(.A1(new_n29391_), .A2(new_n30499_), .B(new_n30584_), .ZN(po0500));
  NAND2_X1   g27349(.A1(new_n30499_), .A2(pi0344), .ZN(new_n30586_));
  OAI21_X1   g27350(.A1(new_n29397_), .A2(new_n30499_), .B(new_n30586_), .ZN(po0501));
  NAND2_X1   g27351(.A1(new_n30499_), .A2(pi0345), .ZN(new_n30588_));
  OAI21_X1   g27352(.A1(new_n29011_), .A2(new_n30499_), .B(new_n30588_), .ZN(po0502));
  NAND2_X1   g27353(.A1(new_n30499_), .A2(pi0346), .ZN(new_n30590_));
  OAI21_X1   g27354(.A1(new_n29404_), .A2(new_n30499_), .B(new_n30590_), .ZN(po0503));
  INV_X1     g27355(.I(pi1055), .ZN(new_n30592_));
  NAND2_X1   g27356(.A1(new_n30499_), .A2(pi0347), .ZN(new_n30593_));
  OAI21_X1   g27357(.A1(new_n30592_), .A2(new_n30499_), .B(new_n30593_), .ZN(po0504));
  INV_X1     g27358(.I(pi1087), .ZN(new_n30595_));
  NAND2_X1   g27359(.A1(new_n30499_), .A2(pi0348), .ZN(new_n30596_));
  OAI21_X1   g27360(.A1(new_n30595_), .A2(new_n30499_), .B(new_n30596_), .ZN(po0505));
  NAND2_X1   g27361(.A1(new_n30499_), .A2(pi0349), .ZN(new_n30598_));
  OAI21_X1   g27362(.A1(new_n30539_), .A2(new_n30499_), .B(new_n30598_), .ZN(po0506));
  INV_X1     g27363(.I(pi1035), .ZN(new_n30600_));
  NAND2_X1   g27364(.A1(new_n30499_), .A2(pi0350), .ZN(new_n30601_));
  OAI21_X1   g27365(.A1(new_n30600_), .A2(new_n30499_), .B(new_n30601_), .ZN(po0507));
  INV_X1     g27366(.I(pi1079), .ZN(new_n30603_));
  NAND2_X1   g27367(.A1(new_n30499_), .A2(pi0351), .ZN(new_n30604_));
  OAI21_X1   g27368(.A1(new_n30603_), .A2(new_n30499_), .B(new_n30604_), .ZN(po0508));
  INV_X1     g27369(.I(pi1078), .ZN(new_n30606_));
  NAND2_X1   g27370(.A1(new_n30499_), .A2(pi0352), .ZN(new_n30607_));
  OAI21_X1   g27371(.A1(new_n30606_), .A2(new_n30499_), .B(new_n30607_), .ZN(po0509));
  NAND2_X1   g27372(.A1(new_n30499_), .A2(pi0353), .ZN(new_n30609_));
  OAI21_X1   g27373(.A1(new_n30529_), .A2(new_n30499_), .B(new_n30609_), .ZN(po0510));
  INV_X1     g27374(.I(pi1045), .ZN(new_n30611_));
  NAND2_X1   g27375(.A1(new_n30499_), .A2(pi0354), .ZN(new_n30612_));
  OAI21_X1   g27376(.A1(new_n30611_), .A2(new_n30499_), .B(new_n30612_), .ZN(po0511));
  NAND2_X1   g27377(.A1(new_n30499_), .A2(pi0355), .ZN(new_n30614_));
  OAI21_X1   g27378(.A1(new_n30393_), .A2(new_n30499_), .B(new_n30614_), .ZN(po0512));
  INV_X1     g27379(.I(pi1081), .ZN(new_n30616_));
  NAND2_X1   g27380(.A1(new_n30499_), .A2(pi0356), .ZN(new_n30617_));
  OAI21_X1   g27381(.A1(new_n30616_), .A2(new_n30499_), .B(new_n30617_), .ZN(po0513));
  INV_X1     g27382(.I(pi1076), .ZN(new_n30619_));
  NAND2_X1   g27383(.A1(new_n30499_), .A2(pi0357), .ZN(new_n30620_));
  OAI21_X1   g27384(.A1(new_n30619_), .A2(new_n30499_), .B(new_n30620_), .ZN(po0514));
  INV_X1     g27385(.I(pi1071), .ZN(new_n30622_));
  NAND2_X1   g27386(.A1(new_n30499_), .A2(pi0358), .ZN(new_n30623_));
  OAI21_X1   g27387(.A1(new_n30622_), .A2(new_n30499_), .B(new_n30623_), .ZN(po0515));
  INV_X1     g27388(.I(pi1068), .ZN(new_n30625_));
  NAND2_X1   g27389(.A1(new_n30499_), .A2(pi0359), .ZN(new_n30626_));
  OAI21_X1   g27390(.A1(new_n30625_), .A2(new_n30499_), .B(new_n30626_), .ZN(po0516));
  INV_X1     g27391(.I(pi1042), .ZN(new_n30628_));
  NAND2_X1   g27392(.A1(new_n30499_), .A2(pi0360), .ZN(new_n30629_));
  OAI21_X1   g27393(.A1(new_n30628_), .A2(new_n30499_), .B(new_n30629_), .ZN(po0517));
  NAND2_X1   g27394(.A1(new_n30499_), .A2(pi0361), .ZN(new_n30631_));
  OAI21_X1   g27395(.A1(new_n30396_), .A2(new_n30499_), .B(new_n30631_), .ZN(po0518));
  NAND2_X1   g27396(.A1(new_n30499_), .A2(pi0362), .ZN(new_n30633_));
  OAI21_X1   g27397(.A1(new_n29379_), .A2(new_n30499_), .B(new_n30633_), .ZN(po0519));
  NAND2_X1   g27398(.A1(new_n30568_), .A2(pi0363), .ZN(new_n30635_));
  OAI21_X1   g27399(.A1(new_n30390_), .A2(new_n30568_), .B(new_n30635_), .ZN(po0520));
  INV_X1     g27400(.I(pi0364), .ZN(new_n30637_));
  NAND2_X1   g27401(.A1(new_n30506_), .A2(pi1062), .ZN(new_n30638_));
  OAI21_X1   g27402(.A1(new_n30637_), .A2(new_n30506_), .B(new_n30638_), .ZN(po0521));
  NAND2_X1   g27403(.A1(new_n30568_), .A2(pi0365), .ZN(new_n30640_));
  OAI21_X1   g27404(.A1(new_n29385_), .A2(new_n30568_), .B(new_n30640_), .ZN(po0522));
  NAND2_X1   g27405(.A1(new_n30568_), .A2(pi0366), .ZN(new_n30642_));
  OAI21_X1   g27406(.A1(new_n29397_), .A2(new_n30568_), .B(new_n30642_), .ZN(po0523));
  INV_X1     g27407(.I(pi0367), .ZN(new_n30644_));
  NAND2_X1   g27408(.A1(new_n30506_), .A2(pi1039), .ZN(new_n30645_));
  OAI21_X1   g27409(.A1(new_n30644_), .A2(new_n30506_), .B(new_n30645_), .ZN(po0524));
  NAND2_X1   g27410(.A1(new_n30506_), .A2(pi1067), .ZN(new_n30647_));
  OAI21_X1   g27411(.A1(new_n6321_), .A2(new_n30506_), .B(new_n30647_), .ZN(po0525));
  NAND2_X1   g27412(.A1(new_n30506_), .A2(pi1080), .ZN(new_n30649_));
  OAI21_X1   g27413(.A1(new_n9228_), .A2(new_n30506_), .B(new_n30649_), .ZN(po0526));
  NAND2_X1   g27414(.A1(new_n30568_), .A2(pi0370), .ZN(new_n30651_));
  OAI21_X1   g27415(.A1(new_n30592_), .A2(new_n30568_), .B(new_n30651_), .ZN(po0527));
  NAND2_X1   g27416(.A1(new_n30506_), .A2(pi1051), .ZN(new_n30653_));
  OAI21_X1   g27417(.A1(new_n6672_), .A2(new_n30506_), .B(new_n30653_), .ZN(po0528));
  NAND2_X1   g27418(.A1(new_n30506_), .A2(pi1048), .ZN(new_n30655_));
  OAI21_X1   g27419(.A1(new_n6331_), .A2(new_n30506_), .B(new_n30655_), .ZN(po0529));
  NAND2_X1   g27420(.A1(new_n30506_), .A2(pi1087), .ZN(new_n30657_));
  OAI21_X1   g27421(.A1(new_n6396_), .A2(new_n30506_), .B(new_n30657_), .ZN(po0530));
  NAND2_X1   g27422(.A1(new_n30506_), .A2(pi1035), .ZN(new_n30659_));
  OAI21_X1   g27423(.A1(new_n6689_), .A2(new_n30506_), .B(new_n30659_), .ZN(po0531));
  NAND2_X1   g27424(.A1(new_n30568_), .A2(pi0375), .ZN(new_n30661_));
  OAI21_X1   g27425(.A1(new_n30502_), .A2(new_n30568_), .B(new_n30661_), .ZN(po0532));
  NAND2_X1   g27426(.A1(new_n30506_), .A2(pi1079), .ZN(new_n30663_));
  OAI21_X1   g27427(.A1(new_n6355_), .A2(new_n30506_), .B(new_n30663_), .ZN(po0533));
  NAND2_X1   g27428(.A1(new_n30506_), .A2(pi1074), .ZN(new_n30665_));
  OAI21_X1   g27429(.A1(new_n6354_), .A2(new_n30506_), .B(new_n30665_), .ZN(po0534));
  NAND2_X1   g27430(.A1(new_n30506_), .A2(pi1063), .ZN(new_n30667_));
  OAI21_X1   g27431(.A1(new_n6358_), .A2(new_n30506_), .B(new_n30667_), .ZN(po0535));
  INV_X1     g27432(.I(pi0379), .ZN(new_n30669_));
  NAND2_X1   g27433(.A1(new_n30506_), .A2(pi1045), .ZN(new_n30670_));
  OAI21_X1   g27434(.A1(new_n30669_), .A2(new_n30506_), .B(new_n30670_), .ZN(po0536));
  INV_X1     g27435(.I(pi0380), .ZN(new_n30672_));
  NAND2_X1   g27436(.A1(new_n30506_), .A2(pi1084), .ZN(new_n30673_));
  OAI21_X1   g27437(.A1(new_n30672_), .A2(new_n30506_), .B(new_n30673_), .ZN(po0537));
  NAND2_X1   g27438(.A1(new_n30568_), .A2(pi0381), .ZN(new_n30675_));
  OAI21_X1   g27439(.A1(new_n30616_), .A2(new_n30568_), .B(new_n30675_), .ZN(po0538));
  NAND2_X1   g27440(.A1(new_n30568_), .A2(pi0382), .ZN(new_n30677_));
  OAI21_X1   g27441(.A1(new_n30619_), .A2(new_n30568_), .B(new_n30677_), .ZN(po0539));
  NAND2_X1   g27442(.A1(new_n30506_), .A2(pi1071), .ZN(new_n30679_));
  OAI21_X1   g27443(.A1(new_n6314_), .A2(new_n30506_), .B(new_n30679_), .ZN(po0540));
  NAND2_X1   g27444(.A1(new_n30506_), .A2(pi1068), .ZN(new_n30681_));
  OAI21_X1   g27445(.A1(new_n6409_), .A2(new_n30506_), .B(new_n30681_), .ZN(po0541));
  NAND2_X1   g27446(.A1(new_n30506_), .A2(pi1042), .ZN(new_n30683_));
  OAI21_X1   g27447(.A1(new_n6359_), .A2(new_n30506_), .B(new_n30683_), .ZN(po0542));
  NAND2_X1   g27448(.A1(new_n30506_), .A2(pi1059), .ZN(new_n30685_));
  OAI21_X1   g27449(.A1(new_n6333_), .A2(new_n30506_), .B(new_n30685_), .ZN(po0543));
  NAND2_X1   g27450(.A1(new_n30506_), .A2(pi1053), .ZN(new_n30687_));
  OAI21_X1   g27451(.A1(new_n6337_), .A2(new_n30506_), .B(new_n30687_), .ZN(po0544));
  INV_X1     g27452(.I(pi0388), .ZN(new_n30689_));
  NAND2_X1   g27453(.A1(new_n30506_), .A2(pi1037), .ZN(new_n30690_));
  OAI21_X1   g27454(.A1(new_n30689_), .A2(new_n30506_), .B(new_n30690_), .ZN(po0545));
  NAND2_X1   g27455(.A1(new_n30506_), .A2(pi1036), .ZN(new_n30692_));
  OAI21_X1   g27456(.A1(new_n6319_), .A2(new_n30506_), .B(new_n30692_), .ZN(po0546));
  NAND2_X1   g27457(.A1(new_n30511_), .A2(pi0390), .ZN(new_n30694_));
  OAI21_X1   g27458(.A1(new_n30390_), .A2(new_n30511_), .B(new_n30694_), .ZN(po0547));
  NAND2_X1   g27459(.A1(new_n30511_), .A2(pi0391), .ZN(new_n30696_));
  OAI21_X1   g27460(.A1(new_n29391_), .A2(new_n30511_), .B(new_n30696_), .ZN(po0548));
  NAND2_X1   g27461(.A1(new_n30511_), .A2(pi0392), .ZN(new_n30698_));
  OAI21_X1   g27462(.A1(new_n29011_), .A2(new_n30511_), .B(new_n30698_), .ZN(po0549));
  NAND2_X1   g27463(.A1(new_n30511_), .A2(pi0393), .ZN(new_n30700_));
  OAI21_X1   g27464(.A1(new_n29404_), .A2(new_n30511_), .B(new_n30700_), .ZN(po0550));
  NAND2_X1   g27465(.A1(new_n30511_), .A2(pi0394), .ZN(new_n30702_));
  OAI21_X1   g27466(.A1(new_n30497_), .A2(new_n30511_), .B(new_n30702_), .ZN(po0551));
  NAND2_X1   g27467(.A1(new_n30511_), .A2(pi0395), .ZN(new_n30704_));
  OAI21_X1   g27468(.A1(new_n30592_), .A2(new_n30511_), .B(new_n30704_), .ZN(po0552));
  NAND2_X1   g27469(.A1(new_n30511_), .A2(pi0396), .ZN(new_n30706_));
  OAI21_X1   g27470(.A1(new_n30521_), .A2(new_n30511_), .B(new_n30706_), .ZN(po0553));
  NAND2_X1   g27471(.A1(new_n30511_), .A2(pi0397), .ZN(new_n30708_));
  OAI21_X1   g27472(.A1(new_n30387_), .A2(new_n30511_), .B(new_n30708_), .ZN(po0554));
  NAND2_X1   g27473(.A1(new_n30511_), .A2(pi0398), .ZN(new_n30710_));
  OAI21_X1   g27474(.A1(new_n30595_), .A2(new_n30511_), .B(new_n30710_), .ZN(po0555));
  NAND2_X1   g27475(.A1(new_n30511_), .A2(pi0399), .ZN(new_n30712_));
  OAI21_X1   g27476(.A1(new_n30502_), .A2(new_n30511_), .B(new_n30712_), .ZN(po0556));
  NAND2_X1   g27477(.A1(new_n30511_), .A2(pi0400), .ZN(new_n30714_));
  OAI21_X1   g27478(.A1(new_n30600_), .A2(new_n30511_), .B(new_n30714_), .ZN(po0557));
  NAND2_X1   g27479(.A1(new_n30511_), .A2(pi0401), .ZN(new_n30716_));
  OAI21_X1   g27480(.A1(new_n30603_), .A2(new_n30511_), .B(new_n30716_), .ZN(po0558));
  NAND2_X1   g27481(.A1(new_n30511_), .A2(pi0402), .ZN(new_n30718_));
  OAI21_X1   g27482(.A1(new_n30606_), .A2(new_n30511_), .B(new_n30718_), .ZN(po0559));
  NAND2_X1   g27483(.A1(new_n30511_), .A2(pi0403), .ZN(new_n30720_));
  OAI21_X1   g27484(.A1(new_n30611_), .A2(new_n30511_), .B(new_n30720_), .ZN(po0560));
  NAND2_X1   g27485(.A1(new_n30511_), .A2(pi0404), .ZN(new_n30722_));
  OAI21_X1   g27486(.A1(new_n30393_), .A2(new_n30511_), .B(new_n30722_), .ZN(po0561));
  NAND2_X1   g27487(.A1(new_n30511_), .A2(pi0405), .ZN(new_n30724_));
  OAI21_X1   g27488(.A1(new_n30616_), .A2(new_n30511_), .B(new_n30724_), .ZN(po0562));
  NAND2_X1   g27489(.A1(new_n30511_), .A2(pi0406), .ZN(new_n30726_));
  OAI21_X1   g27490(.A1(new_n30619_), .A2(new_n30511_), .B(new_n30726_), .ZN(po0563));
  NAND2_X1   g27491(.A1(new_n30511_), .A2(pi0407), .ZN(new_n30728_));
  OAI21_X1   g27492(.A1(new_n30622_), .A2(new_n30511_), .B(new_n30728_), .ZN(po0564));
  NAND2_X1   g27493(.A1(new_n30511_), .A2(pi0408), .ZN(new_n30730_));
  OAI21_X1   g27494(.A1(new_n30625_), .A2(new_n30511_), .B(new_n30730_), .ZN(po0565));
  NAND2_X1   g27495(.A1(new_n30511_), .A2(pi0409), .ZN(new_n30732_));
  OAI21_X1   g27496(.A1(new_n30628_), .A2(new_n30511_), .B(new_n30732_), .ZN(po0566));
  NAND2_X1   g27497(.A1(new_n30511_), .A2(pi0410), .ZN(new_n30734_));
  OAI21_X1   g27498(.A1(new_n30396_), .A2(new_n30511_), .B(new_n30734_), .ZN(po0567));
  NAND2_X1   g27499(.A1(new_n30511_), .A2(pi0411), .ZN(new_n30736_));
  OAI21_X1   g27500(.A1(new_n30402_), .A2(new_n30511_), .B(new_n30736_), .ZN(po0568));
  NAND2_X1   g27501(.A1(new_n30511_), .A2(pi0412), .ZN(new_n30738_));
  OAI21_X1   g27502(.A1(new_n30405_), .A2(new_n30511_), .B(new_n30738_), .ZN(po0569));
  NAND2_X1   g27503(.A1(new_n30511_), .A2(pi0413), .ZN(new_n30740_));
  OAI21_X1   g27504(.A1(new_n29374_), .A2(new_n30511_), .B(new_n30740_), .ZN(po0570));
  NAND3_X1   g27505(.A1(new_n30350_), .A2(new_n30548_), .A3(new_n6845_), .ZN(new_n30742_));
  NAND2_X1   g27506(.A1(new_n30742_), .A2(pi0414), .ZN(new_n30743_));
  OAI21_X1   g27507(.A1(new_n30390_), .A2(new_n30742_), .B(new_n30743_), .ZN(po0571));
  NAND2_X1   g27508(.A1(new_n30742_), .A2(pi0415), .ZN(new_n30745_));
  OAI21_X1   g27509(.A1(new_n29391_), .A2(new_n30742_), .B(new_n30745_), .ZN(po0572));
  NAND2_X1   g27510(.A1(new_n30742_), .A2(pi0416), .ZN(new_n30747_));
  OAI21_X1   g27511(.A1(new_n29397_), .A2(new_n30742_), .B(new_n30747_), .ZN(po0573));
  NAND2_X1   g27512(.A1(new_n30742_), .A2(pi0417), .ZN(new_n30749_));
  OAI21_X1   g27513(.A1(new_n29011_), .A2(new_n30742_), .B(new_n30749_), .ZN(po0574));
  NAND2_X1   g27514(.A1(new_n30742_), .A2(pi0418), .ZN(new_n30751_));
  OAI21_X1   g27515(.A1(new_n29404_), .A2(new_n30742_), .B(new_n30751_), .ZN(po0575));
  NAND2_X1   g27516(.A1(new_n30742_), .A2(pi0419), .ZN(new_n30753_));
  OAI21_X1   g27517(.A1(new_n30497_), .A2(new_n30742_), .B(new_n30753_), .ZN(po0576));
  NAND2_X1   g27518(.A1(new_n30742_), .A2(pi0420), .ZN(new_n30755_));
  OAI21_X1   g27519(.A1(new_n30592_), .A2(new_n30742_), .B(new_n30755_), .ZN(po0577));
  NAND2_X1   g27520(.A1(new_n30742_), .A2(pi0421), .ZN(new_n30757_));
  OAI21_X1   g27521(.A1(new_n30521_), .A2(new_n30742_), .B(new_n30757_), .ZN(po0578));
  NAND2_X1   g27522(.A1(new_n30742_), .A2(pi0422), .ZN(new_n30759_));
  OAI21_X1   g27523(.A1(new_n30387_), .A2(new_n30742_), .B(new_n30759_), .ZN(po0579));
  NAND2_X1   g27524(.A1(new_n30742_), .A2(pi0423), .ZN(new_n30761_));
  OAI21_X1   g27525(.A1(new_n30595_), .A2(new_n30742_), .B(new_n30761_), .ZN(po0580));
  NAND2_X1   g27526(.A1(new_n30742_), .A2(pi0424), .ZN(new_n30763_));
  OAI21_X1   g27527(.A1(new_n30502_), .A2(new_n30742_), .B(new_n30763_), .ZN(po0581));
  NAND2_X1   g27528(.A1(new_n30742_), .A2(pi0425), .ZN(new_n30765_));
  OAI21_X1   g27529(.A1(new_n30600_), .A2(new_n30742_), .B(new_n30765_), .ZN(po0582));
  NAND2_X1   g27530(.A1(new_n30742_), .A2(pi0426), .ZN(new_n30767_));
  OAI21_X1   g27531(.A1(new_n30603_), .A2(new_n30742_), .B(new_n30767_), .ZN(po0583));
  NAND2_X1   g27532(.A1(new_n30742_), .A2(pi0427), .ZN(new_n30769_));
  OAI21_X1   g27533(.A1(new_n30606_), .A2(new_n30742_), .B(new_n30769_), .ZN(po0584));
  NAND2_X1   g27534(.A1(new_n30742_), .A2(pi0428), .ZN(new_n30771_));
  OAI21_X1   g27535(.A1(new_n30611_), .A2(new_n30742_), .B(new_n30771_), .ZN(po0585));
  NAND2_X1   g27536(.A1(new_n30742_), .A2(pi0429), .ZN(new_n30773_));
  OAI21_X1   g27537(.A1(new_n30393_), .A2(new_n30742_), .B(new_n30773_), .ZN(po0586));
  NAND2_X1   g27538(.A1(new_n30742_), .A2(pi0430), .ZN(new_n30775_));
  OAI21_X1   g27539(.A1(new_n30619_), .A2(new_n30742_), .B(new_n30775_), .ZN(po0587));
  NAND2_X1   g27540(.A1(new_n30742_), .A2(pi0431), .ZN(new_n30777_));
  OAI21_X1   g27541(.A1(new_n30622_), .A2(new_n30742_), .B(new_n30777_), .ZN(po0588));
  NAND2_X1   g27542(.A1(new_n30742_), .A2(pi0432), .ZN(new_n30779_));
  OAI21_X1   g27543(.A1(new_n30625_), .A2(new_n30742_), .B(new_n30779_), .ZN(po0589));
  NAND2_X1   g27544(.A1(new_n30742_), .A2(pi0433), .ZN(new_n30781_));
  OAI21_X1   g27545(.A1(new_n30628_), .A2(new_n30742_), .B(new_n30781_), .ZN(po0590));
  NAND2_X1   g27546(.A1(new_n30742_), .A2(pi0434), .ZN(new_n30783_));
  OAI21_X1   g27547(.A1(new_n30396_), .A2(new_n30742_), .B(new_n30783_), .ZN(po0591));
  NAND2_X1   g27548(.A1(new_n30742_), .A2(pi0435), .ZN(new_n30785_));
  OAI21_X1   g27549(.A1(new_n30402_), .A2(new_n30742_), .B(new_n30785_), .ZN(po0592));
  NAND2_X1   g27550(.A1(new_n30742_), .A2(pi0436), .ZN(new_n30787_));
  OAI21_X1   g27551(.A1(new_n30405_), .A2(new_n30742_), .B(new_n30787_), .ZN(po0593));
  NAND2_X1   g27552(.A1(new_n30742_), .A2(pi0437), .ZN(new_n30789_));
  OAI21_X1   g27553(.A1(new_n29379_), .A2(new_n30742_), .B(new_n30789_), .ZN(po0594));
  NAND2_X1   g27554(.A1(new_n30742_), .A2(pi0438), .ZN(new_n30791_));
  OAI21_X1   g27555(.A1(new_n29374_), .A2(new_n30742_), .B(new_n30791_), .ZN(po0595));
  NAND2_X1   g27556(.A1(new_n30568_), .A2(pi0439), .ZN(new_n30793_));
  OAI21_X1   g27557(.A1(new_n30532_), .A2(new_n30568_), .B(new_n30793_), .ZN(po0596));
  NAND2_X1   g27558(.A1(new_n30506_), .A2(pi1043), .ZN(new_n30795_));
  OAI21_X1   g27559(.A1(new_n6410_), .A2(new_n30506_), .B(new_n30795_), .ZN(po0597));
  NAND2_X1   g27560(.A1(new_n30499_), .A2(pi0441), .ZN(new_n30797_));
  OAI21_X1   g27561(.A1(new_n30408_), .A2(new_n30499_), .B(new_n30797_), .ZN(po0598));
  NAND2_X1   g27562(.A1(new_n30506_), .A2(pi1058), .ZN(new_n30799_));
  OAI21_X1   g27563(.A1(new_n6412_), .A2(new_n30506_), .B(new_n30799_), .ZN(po0599));
  NAND2_X1   g27564(.A1(new_n30742_), .A2(pi0443), .ZN(new_n30801_));
  OAI21_X1   g27565(.A1(new_n30408_), .A2(new_n30742_), .B(new_n30801_), .ZN(po0600));
  NAND2_X1   g27566(.A1(new_n30742_), .A2(pi0444), .ZN(new_n30803_));
  OAI21_X1   g27567(.A1(new_n30399_), .A2(new_n30742_), .B(new_n30803_), .ZN(po0601));
  NAND2_X1   g27568(.A1(new_n30742_), .A2(pi0445), .ZN(new_n30805_));
  OAI21_X1   g27569(.A1(new_n30616_), .A2(new_n30742_), .B(new_n30805_), .ZN(po0602));
  NAND2_X1   g27570(.A1(new_n30742_), .A2(pi0446), .ZN(new_n30807_));
  OAI21_X1   g27571(.A1(new_n30526_), .A2(new_n30742_), .B(new_n30807_), .ZN(po0603));
  NAND2_X1   g27572(.A1(new_n30568_), .A2(pi0447), .ZN(new_n30809_));
  OAI21_X1   g27573(.A1(new_n29410_), .A2(new_n30568_), .B(new_n30809_), .ZN(po0604));
  NAND2_X1   g27574(.A1(new_n30742_), .A2(pi0448), .ZN(new_n30811_));
  OAI21_X1   g27575(.A1(new_n30509_), .A2(new_n30742_), .B(new_n30811_), .ZN(po0605));
  NAND2_X1   g27576(.A1(new_n30742_), .A2(pi0449), .ZN(new_n30813_));
  OAI21_X1   g27577(.A1(new_n30532_), .A2(new_n30742_), .B(new_n30813_), .ZN(po0606));
  NAND2_X1   g27578(.A1(new_n30499_), .A2(pi0450), .ZN(new_n30815_));
  OAI21_X1   g27579(.A1(new_n29374_), .A2(new_n30499_), .B(new_n30815_), .ZN(po0607));
  NAND2_X1   g27580(.A1(new_n30742_), .A2(pi0451), .ZN(new_n30817_));
  OAI21_X1   g27581(.A1(new_n30529_), .A2(new_n30742_), .B(new_n30817_), .ZN(po0608));
  NAND2_X1   g27582(.A1(new_n30499_), .A2(pi0452), .ZN(new_n30819_));
  OAI21_X1   g27583(.A1(new_n30402_), .A2(new_n30499_), .B(new_n30819_), .ZN(po0609));
  NAND2_X1   g27584(.A1(new_n30742_), .A2(pi0453), .ZN(new_n30821_));
  OAI21_X1   g27585(.A1(new_n29410_), .A2(new_n30742_), .B(new_n30821_), .ZN(po0610));
  NAND2_X1   g27586(.A1(new_n30742_), .A2(pi0454), .ZN(new_n30823_));
  OAI21_X1   g27587(.A1(new_n30539_), .A2(new_n30742_), .B(new_n30823_), .ZN(po0611));
  NAND2_X1   g27588(.A1(new_n30499_), .A2(pi0455), .ZN(new_n30825_));
  OAI21_X1   g27589(.A1(new_n30405_), .A2(new_n30499_), .B(new_n30825_), .ZN(po0612));
  NAND2_X1   g27590(.A1(new_n30511_), .A2(pi0456), .ZN(new_n30827_));
  OAI21_X1   g27591(.A1(new_n30408_), .A2(new_n30511_), .B(new_n30827_), .ZN(po0613));
  INV_X1     g27592(.I(pi0821), .ZN(new_n30829_));
  INV_X1     g27593(.I(pi0815), .ZN(new_n30830_));
  AND2_X2    g27594(.A1(pi0594), .A2(pi0600), .Z(new_n30831_));
  INV_X1     g27595(.I(pi0804), .ZN(new_n30832_));
  INV_X1     g27596(.I(pi0810), .ZN(new_n30833_));
  AOI21_X1   g27597(.A1(pi0600), .A2(new_n30833_), .B(new_n30832_), .ZN(new_n30834_));
  NAND4_X1   g27598(.A1(new_n30834_), .A2(new_n30830_), .A3(new_n30831_), .A4(pi0990), .ZN(new_n30835_));
  INV_X1     g27599(.I(pi0595), .ZN(new_n30836_));
  NOR2_X1    g27600(.A1(pi0596), .A2(pi0599), .ZN(new_n30837_));
  NAND3_X1   g27601(.A1(new_n30837_), .A2(new_n30832_), .A3(pi0810), .ZN(new_n30838_));
  NAND2_X1   g27602(.A1(new_n30838_), .A2(pi0815), .ZN(new_n30839_));
  NAND2_X1   g27603(.A1(new_n30832_), .A2(new_n30833_), .ZN(new_n30840_));
  AOI21_X1   g27604(.A1(new_n30836_), .A2(new_n30840_), .B(new_n30839_), .ZN(new_n30841_));
  NAND4_X1   g27605(.A1(new_n30836_), .A2(new_n30832_), .A3(new_n30833_), .A4(new_n30830_), .ZN(new_n30842_));
  NAND4_X1   g27606(.A1(new_n30842_), .A2(pi0597), .A3(pi0601), .A4(new_n30831_), .ZN(new_n30843_));
  INV_X1     g27607(.I(pi0605), .ZN(new_n30844_));
  INV_X1     g27608(.I(pi0601), .ZN(new_n30845_));
  NAND2_X1   g27609(.A1(new_n30840_), .A2(new_n30845_), .ZN(new_n30846_));
  NOR2_X1    g27610(.A1(new_n30834_), .A2(pi0815), .ZN(new_n30847_));
  AOI21_X1   g27611(.A1(new_n30847_), .A2(new_n30846_), .B(new_n30844_), .ZN(new_n30848_));
  OAI21_X1   g27612(.A1(new_n30841_), .A2(new_n30843_), .B(new_n30848_), .ZN(new_n30849_));
  AOI21_X1   g27613(.A1(new_n30849_), .A2(new_n30835_), .B(new_n30829_), .ZN(po0614));
  NAND2_X1   g27614(.A1(new_n30499_), .A2(pi0458), .ZN(new_n30851_));
  OAI21_X1   g27615(.A1(new_n30399_), .A2(new_n30499_), .B(new_n30851_), .ZN(po0615));
  NAND2_X1   g27616(.A1(new_n30742_), .A2(pi0459), .ZN(new_n30853_));
  OAI21_X1   g27617(.A1(new_n30518_), .A2(new_n30742_), .B(new_n30853_), .ZN(po0616));
  NAND2_X1   g27618(.A1(new_n30499_), .A2(pi0460), .ZN(new_n30855_));
  OAI21_X1   g27619(.A1(new_n30526_), .A2(new_n30499_), .B(new_n30855_), .ZN(po0617));
  NAND2_X1   g27620(.A1(new_n30499_), .A2(pi0461), .ZN(new_n30857_));
  OAI21_X1   g27621(.A1(new_n30532_), .A2(new_n30499_), .B(new_n30857_), .ZN(po0618));
  NAND2_X1   g27622(.A1(new_n30499_), .A2(pi0462), .ZN(new_n30859_));
  OAI21_X1   g27623(.A1(new_n30509_), .A2(new_n30499_), .B(new_n30859_), .ZN(po0619));
  NAND2_X1   g27624(.A1(new_n30511_), .A2(pi0463), .ZN(new_n30861_));
  OAI21_X1   g27625(.A1(new_n29379_), .A2(new_n30511_), .B(new_n30861_), .ZN(po0620));
  NAND2_X1   g27626(.A1(new_n30742_), .A2(pi0464), .ZN(new_n30863_));
  OAI21_X1   g27627(.A1(new_n29385_), .A2(new_n30742_), .B(new_n30863_), .ZN(po0621));
  NOR2_X1    g27628(.A1(new_n8636_), .A2(new_n8634_), .ZN(new_n30866_));
  NOR2_X1    g27629(.A1(po1038), .A2(new_n30866_), .ZN(new_n30867_));
  AOI21_X1   g27630(.A1(po1038), .A2(new_n30442_), .B(new_n30867_), .ZN(new_n30868_));
  NOR3_X1    g27631(.A1(new_n30469_), .A2(pi0943), .A3(new_n30868_), .ZN(new_n30869_));
  INV_X1     g27632(.I(pi0943), .ZN(new_n30870_));
  INV_X1     g27633(.I(new_n30469_), .ZN(new_n30871_));
  AOI21_X1   g27634(.A1(new_n30870_), .A2(new_n30868_), .B(new_n30871_), .ZN(new_n30872_));
  INV_X1     g27635(.I(new_n30868_), .ZN(new_n30873_));
  NOR2_X1    g27636(.A1(new_n30873_), .A2(new_n30438_), .ZN(new_n30874_));
  NOR2_X1    g27637(.A1(new_n11749_), .A2(new_n3286_), .ZN(new_n30875_));
  AOI21_X1   g27638(.A1(new_n3590_), .A2(new_n11749_), .B(new_n30875_), .ZN(new_n30876_));
  NOR2_X1    g27639(.A1(new_n30870_), .A2(new_n27251_), .ZN(new_n30877_));
  AOI22_X1   g27640(.A1(new_n30874_), .A2(new_n30870_), .B1(new_n30876_), .B2(new_n30877_), .ZN(new_n30878_));
  MUX2_X1    g27641(.I0(new_n2598_), .I1(new_n2531_), .S(pi0299), .Z(new_n30879_));
  MUX2_X1    g27642(.I0(new_n2530_), .I1(new_n30879_), .S(new_n6845_), .Z(new_n30880_));
  NAND3_X1   g27643(.A1(new_n30880_), .A2(new_n28282_), .A3(new_n27251_), .ZN(new_n30881_));
  NOR4_X1    g27644(.A1(new_n30872_), .A2(new_n30878_), .A3(new_n30869_), .A4(new_n30881_), .ZN(po0623));
  NAND2_X1   g27645(.A1(new_n29015_), .A2(pi1001), .ZN(new_n30883_));
  NOR3_X1    g27646(.A1(new_n30883_), .A2(new_n3364_), .A3(pi0287), .ZN(new_n30884_));
  INV_X1     g27647(.I(new_n30884_), .ZN(new_n30885_));
  NOR2_X1    g27648(.A1(new_n26268_), .A2(new_n30885_), .ZN(new_n30886_));
  NAND2_X1   g27649(.A1(new_n9852_), .A2(new_n2462_), .ZN(new_n30887_));
  NAND4_X1   g27650(.A1(new_n30887_), .A2(new_n6988_), .A3(new_n8548_), .A4(new_n12539_), .ZN(new_n30888_));
  NOR2_X1    g27651(.A1(new_n30888_), .A2(new_n12538_), .ZN(new_n30889_));
  AOI21_X1   g27652(.A1(new_n5182_), .A2(new_n30884_), .B(new_n30889_), .ZN(new_n30890_));
  NOR4_X1    g27653(.A1(new_n30888_), .A2(new_n5181_), .A3(new_n12538_), .A4(new_n30885_), .ZN(new_n30891_));
  NOR2_X1    g27654(.A1(new_n30890_), .A2(new_n30891_), .ZN(new_n30892_));
  NOR4_X1    g27655(.A1(new_n30885_), .A2(pi0824), .A3(new_n2927_), .A4(new_n2955_), .ZN(new_n30893_));
  NAND2_X1   g27656(.A1(new_n30893_), .A2(pi1093), .ZN(new_n30894_));
  XOR2_X1    g27657(.A1(new_n30892_), .A2(new_n30894_), .Z(new_n30895_));
  NOR3_X1    g27658(.A1(new_n30885_), .A2(new_n5182_), .A3(new_n6000_), .ZN(new_n30896_));
  XOR2_X1    g27659(.A1(new_n30892_), .A2(new_n30896_), .Z(new_n30897_));
  NOR2_X1    g27660(.A1(new_n30897_), .A2(new_n2918_), .ZN(new_n30898_));
  AOI21_X1   g27661(.A1(new_n2918_), .A2(new_n30895_), .B(new_n30898_), .ZN(new_n30899_));
  NAND3_X1   g27662(.A1(new_n6964_), .A2(new_n2625_), .A3(new_n5226_), .ZN(new_n30900_));
  OAI22_X1   g27663(.A1(new_n30899_), .A2(new_n30900_), .B1(new_n7824_), .B2(new_n30886_), .ZN(po0624));
  INV_X1     g27664(.I(new_n8597_), .ZN(new_n30902_));
  NOR4_X1    g27665(.A1(new_n7793_), .A2(new_n3172_), .A3(pi0039), .A4(new_n7833_), .ZN(new_n30903_));
  OAI22_X1   g27666(.A1(new_n30903_), .A2(new_n9909_), .B1(new_n7856_), .B2(new_n30902_), .ZN(po0625));
  NOR3_X1    g27667(.A1(new_n30469_), .A2(pi0922), .A3(new_n30868_), .ZN(new_n30909_));
  INV_X1     g27668(.I(pi0922), .ZN(new_n30910_));
  AOI21_X1   g27669(.A1(new_n30910_), .A2(new_n30868_), .B(new_n30871_), .ZN(new_n30911_));
  NOR2_X1    g27670(.A1(new_n30910_), .A2(new_n26604_), .ZN(new_n30912_));
  AOI22_X1   g27671(.A1(new_n30874_), .A2(new_n30910_), .B1(new_n30876_), .B2(new_n30912_), .ZN(new_n30913_));
  NAND3_X1   g27672(.A1(new_n30880_), .A2(new_n28280_), .A3(new_n26604_), .ZN(new_n30914_));
  NOR4_X1    g27673(.A1(new_n30911_), .A2(new_n30913_), .A3(new_n30909_), .A4(new_n30914_), .ZN(po0630));
  NOR3_X1    g27674(.A1(new_n30469_), .A2(pi0931), .A3(new_n30868_), .ZN(new_n30916_));
  INV_X1     g27675(.I(pi0931), .ZN(new_n30917_));
  AOI21_X1   g27676(.A1(new_n30917_), .A2(new_n30868_), .B(new_n30871_), .ZN(new_n30918_));
  NOR2_X1    g27677(.A1(new_n30917_), .A2(new_n27817_), .ZN(new_n30919_));
  AOI22_X1   g27678(.A1(new_n30874_), .A2(new_n30917_), .B1(new_n30876_), .B2(new_n30919_), .ZN(new_n30920_));
  NAND3_X1   g27679(.A1(new_n30880_), .A2(new_n28281_), .A3(new_n27817_), .ZN(new_n30921_));
  NOR4_X1    g27680(.A1(new_n30918_), .A2(new_n30920_), .A3(new_n30916_), .A4(new_n30921_), .ZN(po0631));
  NOR3_X1    g27681(.A1(new_n30469_), .A2(pi0936), .A3(new_n30868_), .ZN(new_n30923_));
  INV_X1     g27682(.I(pi0936), .ZN(new_n30924_));
  AOI21_X1   g27683(.A1(new_n30924_), .A2(new_n30868_), .B(new_n30871_), .ZN(new_n30925_));
  NOR2_X1    g27684(.A1(new_n30924_), .A2(new_n27470_), .ZN(new_n30926_));
  AOI22_X1   g27685(.A1(new_n30874_), .A2(new_n30924_), .B1(new_n30876_), .B2(new_n30926_), .ZN(new_n30927_));
  NAND3_X1   g27686(.A1(new_n30880_), .A2(new_n28283_), .A3(new_n27470_), .ZN(new_n30928_));
  NOR4_X1    g27687(.A1(new_n30925_), .A2(new_n30927_), .A3(new_n30923_), .A4(new_n30928_), .ZN(po0632));
  NOR3_X1    g27688(.A1(new_n7819_), .A2(new_n10509_), .A3(new_n8666_), .ZN(new_n30930_));
  NOR3_X1    g27689(.A1(new_n7819_), .A2(new_n10509_), .A3(new_n8666_), .ZN(new_n30931_));
  NOR4_X1    g27690(.A1(new_n30931_), .A2(new_n6999_), .A3(new_n8439_), .A4(new_n8667_), .ZN(new_n30932_));
  NAND4_X1   g27691(.A1(new_n9652_), .A2(new_n2449_), .A3(new_n3233_), .A4(new_n8548_), .ZN(new_n30933_));
  NOR3_X1    g27692(.A1(new_n30932_), .A2(new_n30933_), .A3(new_n30930_), .ZN(new_n30934_));
  NAND3_X1   g27693(.A1(new_n6845_), .A2(pi0071), .A3(new_n8663_), .ZN(new_n30935_));
  NOR2_X1    g27694(.A1(new_n8666_), .A2(new_n5250_), .ZN(new_n30936_));
  OAI21_X1   g27695(.A1(new_n30934_), .A2(new_n30936_), .B(po1038), .ZN(new_n30938_));
  NAND2_X1   g27696(.A1(new_n30938_), .A2(new_n30935_), .ZN(po0633));
  NOR2_X1    g27697(.A1(new_n29982_), .A2(new_n5250_), .ZN(po0635));
  INV_X1     g27698(.I(pi0481), .ZN(new_n30941_));
  NAND2_X1   g27699(.A1(new_n24077_), .A2(pi0248), .ZN(new_n30942_));
  OAI21_X1   g27700(.A1(new_n30941_), .A2(new_n24077_), .B(new_n30942_), .ZN(po0638));
  INV_X1     g27701(.I(pi0482), .ZN(new_n30944_));
  NAND2_X1   g27702(.A1(new_n24089_), .A2(pi0249), .ZN(new_n30945_));
  OAI21_X1   g27703(.A1(new_n30944_), .A2(new_n24089_), .B(new_n30945_), .ZN(po0639));
  INV_X1     g27704(.I(pi0483), .ZN(new_n30947_));
  NAND2_X1   g27705(.A1(new_n24125_), .A2(pi0242), .ZN(new_n30948_));
  OAI21_X1   g27706(.A1(new_n30947_), .A2(new_n24125_), .B(new_n30948_), .ZN(po0640));
  INV_X1     g27707(.I(pi0484), .ZN(new_n30950_));
  NAND2_X1   g27708(.A1(new_n24125_), .A2(pi0249), .ZN(new_n30951_));
  OAI21_X1   g27709(.A1(new_n30950_), .A2(new_n24125_), .B(new_n30951_), .ZN(po0641));
  INV_X1     g27710(.I(pi0485), .ZN(new_n30953_));
  NAND2_X1   g27711(.A1(new_n24931_), .A2(pi0234), .ZN(new_n30954_));
  OAI21_X1   g27712(.A1(new_n30953_), .A2(new_n24931_), .B(new_n30954_), .ZN(po0642));
  INV_X1     g27713(.I(pi0486), .ZN(new_n30956_));
  NAND2_X1   g27714(.A1(new_n24931_), .A2(pi0244), .ZN(new_n30957_));
  OAI21_X1   g27715(.A1(new_n30956_), .A2(new_n24931_), .B(new_n30957_), .ZN(po0643));
  INV_X1     g27716(.I(pi0487), .ZN(new_n30959_));
  NAND2_X1   g27717(.A1(new_n24077_), .A2(pi0246), .ZN(new_n30960_));
  OAI21_X1   g27718(.A1(new_n30959_), .A2(new_n24077_), .B(new_n30960_), .ZN(po0644));
  NAND2_X1   g27719(.A1(new_n24077_), .A2(pi0239), .ZN(new_n30962_));
  OAI21_X1   g27720(.A1(pi0488), .A2(new_n24077_), .B(new_n30962_), .ZN(po0645));
  INV_X1     g27721(.I(pi0489), .ZN(new_n30964_));
  NAND2_X1   g27722(.A1(new_n24931_), .A2(pi0242), .ZN(new_n30965_));
  OAI21_X1   g27723(.A1(new_n30964_), .A2(new_n24931_), .B(new_n30965_), .ZN(po0646));
  INV_X1     g27724(.I(pi0490), .ZN(new_n30967_));
  NAND2_X1   g27725(.A1(new_n24125_), .A2(pi0241), .ZN(new_n30968_));
  OAI21_X1   g27726(.A1(new_n30967_), .A2(new_n24125_), .B(new_n30968_), .ZN(po0647));
  INV_X1     g27727(.I(pi0491), .ZN(new_n30970_));
  NAND2_X1   g27728(.A1(new_n24125_), .A2(pi0238), .ZN(new_n30971_));
  OAI21_X1   g27729(.A1(new_n30970_), .A2(new_n24125_), .B(new_n30971_), .ZN(po0648));
  INV_X1     g27730(.I(pi0492), .ZN(new_n30973_));
  NAND2_X1   g27731(.A1(new_n24125_), .A2(pi0240), .ZN(new_n30974_));
  OAI21_X1   g27732(.A1(new_n30973_), .A2(new_n24125_), .B(new_n30974_), .ZN(po0649));
  INV_X1     g27733(.I(pi0493), .ZN(new_n30976_));
  NAND2_X1   g27734(.A1(new_n24125_), .A2(pi0244), .ZN(new_n30977_));
  OAI21_X1   g27735(.A1(new_n30976_), .A2(new_n24125_), .B(new_n30977_), .ZN(po0650));
  NAND2_X1   g27736(.A1(new_n24125_), .A2(pi0239), .ZN(new_n30979_));
  OAI21_X1   g27737(.A1(pi0494), .A2(new_n24125_), .B(new_n30979_), .ZN(po0651));
  INV_X1     g27738(.I(pi0495), .ZN(new_n30981_));
  NAND2_X1   g27739(.A1(new_n24125_), .A2(pi0235), .ZN(new_n30982_));
  OAI21_X1   g27740(.A1(new_n30981_), .A2(new_n24125_), .B(new_n30982_), .ZN(po0652));
  INV_X1     g27741(.I(pi0496), .ZN(new_n30984_));
  NAND2_X1   g27742(.A1(new_n24119_), .A2(pi0249), .ZN(new_n30985_));
  OAI21_X1   g27743(.A1(new_n30984_), .A2(new_n24119_), .B(new_n30985_), .ZN(po0653));
  NAND2_X1   g27744(.A1(new_n24119_), .A2(pi0239), .ZN(new_n30987_));
  OAI21_X1   g27745(.A1(pi0497), .A2(new_n24119_), .B(new_n30987_), .ZN(po0654));
  INV_X1     g27746(.I(pi0498), .ZN(new_n30989_));
  NAND2_X1   g27747(.A1(new_n24089_), .A2(pi0238), .ZN(new_n30990_));
  OAI21_X1   g27748(.A1(new_n30989_), .A2(new_n24089_), .B(new_n30990_), .ZN(po0655));
  INV_X1     g27749(.I(pi0499), .ZN(new_n30992_));
  NAND2_X1   g27750(.A1(new_n24119_), .A2(pi0246), .ZN(new_n30993_));
  OAI21_X1   g27751(.A1(new_n30992_), .A2(new_n24119_), .B(new_n30993_), .ZN(po0656));
  INV_X1     g27752(.I(pi0500), .ZN(new_n30995_));
  NAND2_X1   g27753(.A1(new_n24119_), .A2(pi0241), .ZN(new_n30996_));
  OAI21_X1   g27754(.A1(new_n30995_), .A2(new_n24119_), .B(new_n30996_), .ZN(po0657));
  INV_X1     g27755(.I(pi0501), .ZN(new_n30998_));
  NAND2_X1   g27756(.A1(new_n24119_), .A2(pi0248), .ZN(new_n30999_));
  OAI21_X1   g27757(.A1(new_n30998_), .A2(new_n24119_), .B(new_n30999_), .ZN(po0658));
  INV_X1     g27758(.I(pi0502), .ZN(new_n31001_));
  NAND2_X1   g27759(.A1(new_n24119_), .A2(pi0247), .ZN(new_n31002_));
  OAI21_X1   g27760(.A1(new_n31001_), .A2(new_n24119_), .B(new_n31002_), .ZN(po0659));
  INV_X1     g27761(.I(pi0503), .ZN(new_n31004_));
  NAND2_X1   g27762(.A1(new_n24119_), .A2(pi0245), .ZN(new_n31005_));
  OAI21_X1   g27763(.A1(new_n31004_), .A2(new_n24119_), .B(new_n31005_), .ZN(po0660));
  INV_X1     g27764(.I(pi0504), .ZN(new_n31007_));
  NAND2_X1   g27765(.A1(new_n24115_), .A2(pi0242), .ZN(new_n31008_));
  OAI21_X1   g27766(.A1(new_n31007_), .A2(new_n24115_), .B(new_n31008_), .ZN(po0661));
  INV_X1     g27767(.I(pi0505), .ZN(new_n31010_));
  NOR2_X1    g27768(.A1(new_n24114_), .A2(new_n2440_), .ZN(new_n31011_));
  NAND3_X1   g27769(.A1(new_n31011_), .A2(new_n31010_), .A3(new_n24080_), .ZN(new_n31012_));
  NOR3_X1    g27770(.A1(new_n5238_), .A2(new_n5220_), .A3(new_n11749_), .ZN(new_n31013_));
  AOI21_X1   g27771(.A1(new_n5238_), .A2(new_n27783_), .B(new_n5219_), .ZN(new_n31014_));
  NOR2_X1    g27772(.A1(new_n31013_), .A2(new_n31014_), .ZN(new_n31015_));
  INV_X1     g27773(.I(new_n31015_), .ZN(new_n31016_));
  NAND2_X1   g27774(.A1(new_n31016_), .A2(new_n2440_), .ZN(new_n31017_));
  NAND2_X1   g27775(.A1(new_n24119_), .A2(new_n31010_), .ZN(new_n31018_));
  OAI21_X1   g27776(.A1(new_n31017_), .A2(new_n31018_), .B(new_n31012_), .ZN(po0662));
  INV_X1     g27777(.I(pi0506), .ZN(new_n31020_));
  NAND2_X1   g27778(.A1(new_n24115_), .A2(pi0241), .ZN(new_n31021_));
  OAI21_X1   g27779(.A1(new_n31020_), .A2(new_n24115_), .B(new_n31021_), .ZN(po0663));
  INV_X1     g27780(.I(pi0507), .ZN(new_n31023_));
  NAND2_X1   g27781(.A1(new_n24115_), .A2(pi0238), .ZN(new_n31024_));
  OAI21_X1   g27782(.A1(new_n31023_), .A2(new_n24115_), .B(new_n31024_), .ZN(po0664));
  INV_X1     g27783(.I(pi0508), .ZN(new_n31026_));
  NAND2_X1   g27784(.A1(new_n24115_), .A2(pi0247), .ZN(new_n31027_));
  OAI21_X1   g27785(.A1(new_n31026_), .A2(new_n24115_), .B(new_n31027_), .ZN(po0665));
  INV_X1     g27786(.I(pi0509), .ZN(new_n31029_));
  NAND2_X1   g27787(.A1(new_n24115_), .A2(pi0245), .ZN(new_n31030_));
  OAI21_X1   g27788(.A1(new_n31029_), .A2(new_n24115_), .B(new_n31030_), .ZN(po0666));
  INV_X1     g27789(.I(pi0510), .ZN(new_n31032_));
  NAND2_X1   g27790(.A1(new_n24077_), .A2(pi0242), .ZN(new_n31033_));
  OAI21_X1   g27791(.A1(new_n31032_), .A2(new_n24077_), .B(new_n31033_), .ZN(po0667));
  NOR3_X1    g27792(.A1(new_n5430_), .A2(new_n5446_), .A3(new_n11749_), .ZN(new_n31035_));
  AOI21_X1   g27793(.A1(new_n5446_), .A2(new_n27783_), .B(new_n5429_), .ZN(new_n31036_));
  NOR2_X1    g27794(.A1(new_n31035_), .A2(new_n31036_), .ZN(new_n31037_));
  INV_X1     g27795(.I(new_n31037_), .ZN(new_n31038_));
  NAND2_X1   g27796(.A1(new_n31038_), .A2(new_n2440_), .ZN(new_n31039_));
  MUX2_X1    g27797(.I0(pi0511), .I1(new_n31039_), .S(new_n24077_), .Z(po0668));
  INV_X1     g27798(.I(pi0512), .ZN(new_n31041_));
  NAND2_X1   g27799(.A1(new_n24077_), .A2(pi0235), .ZN(new_n31042_));
  OAI21_X1   g27800(.A1(new_n31041_), .A2(new_n24077_), .B(new_n31042_), .ZN(po0669));
  INV_X1     g27801(.I(pi0513), .ZN(new_n31044_));
  NAND2_X1   g27802(.A1(new_n24077_), .A2(pi0244), .ZN(new_n31045_));
  OAI21_X1   g27803(.A1(new_n31044_), .A2(new_n24077_), .B(new_n31045_), .ZN(po0670));
  INV_X1     g27804(.I(pi0514), .ZN(new_n31047_));
  NAND2_X1   g27805(.A1(new_n24077_), .A2(pi0245), .ZN(new_n31048_));
  OAI21_X1   g27806(.A1(new_n31047_), .A2(new_n24077_), .B(new_n31048_), .ZN(po0671));
  INV_X1     g27807(.I(pi0515), .ZN(new_n31050_));
  NAND2_X1   g27808(.A1(new_n24077_), .A2(pi0240), .ZN(new_n31051_));
  OAI21_X1   g27809(.A1(new_n31050_), .A2(new_n24077_), .B(new_n31051_), .ZN(po0672));
  INV_X1     g27810(.I(pi0516), .ZN(new_n31053_));
  NAND2_X1   g27811(.A1(new_n24077_), .A2(pi0247), .ZN(new_n31054_));
  OAI21_X1   g27812(.A1(new_n31053_), .A2(new_n24077_), .B(new_n31054_), .ZN(po0673));
  INV_X1     g27813(.I(pi0517), .ZN(new_n31056_));
  NAND2_X1   g27814(.A1(new_n24077_), .A2(pi0238), .ZN(new_n31057_));
  OAI21_X1   g27815(.A1(new_n31056_), .A2(new_n24077_), .B(new_n31057_), .ZN(po0674));
  INV_X1     g27816(.I(pi0518), .ZN(new_n31059_));
  NOR2_X1    g27817(.A1(new_n24076_), .A2(new_n2440_), .ZN(new_n31060_));
  NAND3_X1   g27818(.A1(new_n31060_), .A2(new_n31059_), .A3(new_n24080_), .ZN(new_n31061_));
  NAND2_X1   g27819(.A1(new_n24083_), .A2(new_n31059_), .ZN(new_n31062_));
  OAI21_X1   g27820(.A1(new_n31039_), .A2(new_n31062_), .B(new_n31061_), .ZN(po0675));
  NAND2_X1   g27821(.A1(new_n24083_), .A2(pi0239), .ZN(new_n31064_));
  OAI21_X1   g27822(.A1(pi0519), .A2(new_n24083_), .B(new_n31064_), .ZN(po0676));
  INV_X1     g27823(.I(pi0520), .ZN(new_n31066_));
  NAND2_X1   g27824(.A1(new_n24083_), .A2(pi0246), .ZN(new_n31067_));
  OAI21_X1   g27825(.A1(new_n31066_), .A2(new_n24083_), .B(new_n31067_), .ZN(po0677));
  INV_X1     g27826(.I(pi0521), .ZN(new_n31069_));
  NAND2_X1   g27827(.A1(new_n24083_), .A2(pi0248), .ZN(new_n31070_));
  OAI21_X1   g27828(.A1(new_n31069_), .A2(new_n24083_), .B(new_n31070_), .ZN(po0678));
  INV_X1     g27829(.I(pi0522), .ZN(new_n31072_));
  NAND2_X1   g27830(.A1(new_n24083_), .A2(pi0238), .ZN(new_n31073_));
  OAI21_X1   g27831(.A1(new_n31072_), .A2(new_n24083_), .B(new_n31073_), .ZN(po0679));
  INV_X1     g27832(.I(pi0523), .ZN(new_n31075_));
  NAND3_X1   g27833(.A1(new_n31060_), .A2(new_n31075_), .A3(new_n24122_), .ZN(new_n31076_));
  NAND2_X1   g27834(.A1(new_n24947_), .A2(new_n31075_), .ZN(new_n31077_));
  OAI21_X1   g27835(.A1(new_n31039_), .A2(new_n31077_), .B(new_n31076_), .ZN(po0680));
  NAND2_X1   g27836(.A1(new_n24947_), .A2(pi0239), .ZN(new_n31079_));
  OAI21_X1   g27837(.A1(pi0524), .A2(new_n24947_), .B(new_n31079_), .ZN(po0681));
  INV_X1     g27838(.I(pi0525), .ZN(new_n31081_));
  NAND2_X1   g27839(.A1(new_n24947_), .A2(pi0245), .ZN(new_n31082_));
  OAI21_X1   g27840(.A1(new_n31081_), .A2(new_n24947_), .B(new_n31082_), .ZN(po0682));
  INV_X1     g27841(.I(pi0526), .ZN(new_n31084_));
  NAND2_X1   g27842(.A1(new_n24947_), .A2(pi0246), .ZN(new_n31085_));
  OAI21_X1   g27843(.A1(new_n31084_), .A2(new_n24947_), .B(new_n31085_), .ZN(po0683));
  INV_X1     g27844(.I(pi0527), .ZN(new_n31087_));
  NAND2_X1   g27845(.A1(new_n24947_), .A2(pi0247), .ZN(new_n31088_));
  OAI21_X1   g27846(.A1(new_n31087_), .A2(new_n24947_), .B(new_n31088_), .ZN(po0684));
  INV_X1     g27847(.I(pi0528), .ZN(new_n31090_));
  NAND2_X1   g27848(.A1(new_n24947_), .A2(pi0249), .ZN(new_n31091_));
  OAI21_X1   g27849(.A1(new_n31090_), .A2(new_n24947_), .B(new_n31091_), .ZN(po0685));
  INV_X1     g27850(.I(pi0529), .ZN(new_n31093_));
  NAND2_X1   g27851(.A1(new_n24947_), .A2(pi0238), .ZN(new_n31094_));
  OAI21_X1   g27852(.A1(new_n31093_), .A2(new_n24947_), .B(new_n31094_), .ZN(po0686));
  INV_X1     g27853(.I(pi0530), .ZN(new_n31096_));
  NAND2_X1   g27854(.A1(new_n24947_), .A2(pi0240), .ZN(new_n31097_));
  OAI21_X1   g27855(.A1(new_n31096_), .A2(new_n24947_), .B(new_n31097_), .ZN(po0687));
  INV_X1     g27856(.I(pi0531), .ZN(new_n31099_));
  NAND2_X1   g27857(.A1(new_n24089_), .A2(pi0235), .ZN(new_n31100_));
  OAI21_X1   g27858(.A1(new_n31099_), .A2(new_n24089_), .B(new_n31100_), .ZN(po0688));
  INV_X1     g27859(.I(pi0532), .ZN(new_n31102_));
  NAND2_X1   g27860(.A1(new_n24089_), .A2(pi0247), .ZN(new_n31103_));
  OAI21_X1   g27861(.A1(new_n31102_), .A2(new_n24089_), .B(new_n31103_), .ZN(po0689));
  INV_X1     g27862(.I(pi0533), .ZN(new_n31105_));
  NAND2_X1   g27863(.A1(new_n24115_), .A2(pi0235), .ZN(new_n31106_));
  OAI21_X1   g27864(.A1(new_n31105_), .A2(new_n24115_), .B(new_n31106_), .ZN(po0690));
  NAND2_X1   g27865(.A1(new_n24115_), .A2(pi0239), .ZN(new_n31108_));
  OAI21_X1   g27866(.A1(pi0534), .A2(new_n24115_), .B(new_n31108_), .ZN(po0691));
  INV_X1     g27867(.I(pi0535), .ZN(new_n31110_));
  NAND2_X1   g27868(.A1(new_n24115_), .A2(pi0240), .ZN(new_n31111_));
  OAI21_X1   g27869(.A1(new_n31110_), .A2(new_n24115_), .B(new_n31111_), .ZN(po0692));
  INV_X1     g27870(.I(pi0536), .ZN(new_n31113_));
  NAND2_X1   g27871(.A1(new_n24115_), .A2(pi0246), .ZN(new_n31114_));
  OAI21_X1   g27872(.A1(new_n31113_), .A2(new_n24115_), .B(new_n31114_), .ZN(po0693));
  INV_X1     g27873(.I(pi0537), .ZN(new_n31116_));
  NAND2_X1   g27874(.A1(new_n24115_), .A2(pi0248), .ZN(new_n31117_));
  OAI21_X1   g27875(.A1(new_n31116_), .A2(new_n24115_), .B(new_n31117_), .ZN(po0694));
  INV_X1     g27876(.I(pi0538), .ZN(new_n31119_));
  NAND2_X1   g27877(.A1(new_n24115_), .A2(pi0249), .ZN(new_n31120_));
  OAI21_X1   g27878(.A1(new_n31119_), .A2(new_n24115_), .B(new_n31120_), .ZN(po0695));
  INV_X1     g27879(.I(pi0539), .ZN(new_n31122_));
  NAND2_X1   g27880(.A1(new_n24119_), .A2(pi0242), .ZN(new_n31123_));
  OAI21_X1   g27881(.A1(new_n31122_), .A2(new_n24119_), .B(new_n31123_), .ZN(po0696));
  INV_X1     g27882(.I(pi0540), .ZN(new_n31125_));
  NAND2_X1   g27883(.A1(new_n24119_), .A2(pi0235), .ZN(new_n31126_));
  OAI21_X1   g27884(.A1(new_n31125_), .A2(new_n24119_), .B(new_n31126_), .ZN(po0697));
  INV_X1     g27885(.I(pi0541), .ZN(new_n31128_));
  NAND2_X1   g27886(.A1(new_n24119_), .A2(pi0244), .ZN(new_n31129_));
  OAI21_X1   g27887(.A1(new_n31128_), .A2(new_n24119_), .B(new_n31129_), .ZN(po0698));
  INV_X1     g27888(.I(pi0542), .ZN(new_n31131_));
  NAND2_X1   g27889(.A1(new_n24119_), .A2(pi0240), .ZN(new_n31132_));
  OAI21_X1   g27890(.A1(new_n31131_), .A2(new_n24119_), .B(new_n31132_), .ZN(po0699));
  INV_X1     g27891(.I(pi0543), .ZN(new_n31134_));
  NAND2_X1   g27892(.A1(new_n24119_), .A2(pi0238), .ZN(new_n31135_));
  OAI21_X1   g27893(.A1(new_n31134_), .A2(new_n24119_), .B(new_n31135_), .ZN(po0700));
  INV_X1     g27894(.I(pi0544), .ZN(new_n31137_));
  NAND3_X1   g27895(.A1(new_n31011_), .A2(new_n31137_), .A3(new_n24122_), .ZN(new_n31138_));
  NAND2_X1   g27896(.A1(new_n24125_), .A2(new_n31137_), .ZN(new_n31139_));
  OAI21_X1   g27897(.A1(new_n31017_), .A2(new_n31139_), .B(new_n31138_), .ZN(po0701));
  INV_X1     g27898(.I(pi0545), .ZN(new_n31141_));
  NAND2_X1   g27899(.A1(new_n24125_), .A2(pi0245), .ZN(new_n31142_));
  OAI21_X1   g27900(.A1(new_n31141_), .A2(new_n24125_), .B(new_n31142_), .ZN(po0702));
  INV_X1     g27901(.I(pi0546), .ZN(new_n31144_));
  NAND2_X1   g27902(.A1(new_n24125_), .A2(pi0246), .ZN(new_n31145_));
  OAI21_X1   g27903(.A1(new_n31144_), .A2(new_n24125_), .B(new_n31145_), .ZN(po0703));
  INV_X1     g27904(.I(pi0547), .ZN(new_n31147_));
  NAND2_X1   g27905(.A1(new_n24125_), .A2(pi0247), .ZN(new_n31148_));
  OAI21_X1   g27906(.A1(new_n31147_), .A2(new_n24125_), .B(new_n31148_), .ZN(po0704));
  INV_X1     g27907(.I(pi0548), .ZN(new_n31150_));
  NAND2_X1   g27908(.A1(new_n24125_), .A2(pi0248), .ZN(new_n31151_));
  OAI21_X1   g27909(.A1(new_n31150_), .A2(new_n24125_), .B(new_n31151_), .ZN(po0705));
  INV_X1     g27910(.I(pi0549), .ZN(new_n31153_));
  NAND2_X1   g27911(.A1(new_n24931_), .A2(pi0235), .ZN(new_n31154_));
  OAI21_X1   g27912(.A1(new_n31153_), .A2(new_n24931_), .B(new_n31154_), .ZN(po0706));
  NAND2_X1   g27913(.A1(new_n24931_), .A2(pi0239), .ZN(new_n31156_));
  OAI21_X1   g27914(.A1(pi0550), .A2(new_n24931_), .B(new_n31156_), .ZN(po0707));
  INV_X1     g27915(.I(pi0551), .ZN(new_n31158_));
  NAND2_X1   g27916(.A1(new_n24931_), .A2(pi0240), .ZN(new_n31159_));
  OAI21_X1   g27917(.A1(new_n31158_), .A2(new_n24931_), .B(new_n31159_), .ZN(po0708));
  INV_X1     g27918(.I(pi0552), .ZN(new_n31161_));
  NAND2_X1   g27919(.A1(new_n24931_), .A2(pi0247), .ZN(new_n31162_));
  OAI21_X1   g27920(.A1(new_n31161_), .A2(new_n24931_), .B(new_n31162_), .ZN(po0709));
  INV_X1     g27921(.I(pi0553), .ZN(new_n31164_));
  NAND2_X1   g27922(.A1(new_n24931_), .A2(pi0241), .ZN(new_n31165_));
  OAI21_X1   g27923(.A1(new_n31164_), .A2(new_n24931_), .B(new_n31165_), .ZN(po0710));
  INV_X1     g27924(.I(pi0554), .ZN(new_n31167_));
  NAND2_X1   g27925(.A1(new_n24931_), .A2(pi0248), .ZN(new_n31168_));
  OAI21_X1   g27926(.A1(new_n31167_), .A2(new_n24931_), .B(new_n31168_), .ZN(po0711));
  INV_X1     g27927(.I(pi0555), .ZN(new_n31170_));
  NAND2_X1   g27928(.A1(new_n24931_), .A2(pi0249), .ZN(new_n31171_));
  OAI21_X1   g27929(.A1(new_n31170_), .A2(new_n24931_), .B(new_n31171_), .ZN(po0712));
  INV_X1     g27930(.I(pi0556), .ZN(new_n31173_));
  NAND2_X1   g27931(.A1(new_n24089_), .A2(pi0242), .ZN(new_n31174_));
  OAI21_X1   g27932(.A1(new_n31173_), .A2(new_n24089_), .B(new_n31174_), .ZN(po0713));
  INV_X1     g27933(.I(pi0557), .ZN(new_n31176_));
  NAND3_X1   g27934(.A1(new_n31011_), .A2(new_n31176_), .A3(new_n24071_), .ZN(new_n31177_));
  NAND2_X1   g27935(.A1(new_n24115_), .A2(new_n31176_), .ZN(new_n31178_));
  OAI21_X1   g27936(.A1(new_n31017_), .A2(new_n31178_), .B(new_n31177_), .ZN(po0714));
  INV_X1     g27937(.I(pi0558), .ZN(new_n31180_));
  NAND2_X1   g27938(.A1(new_n24115_), .A2(pi0244), .ZN(new_n31181_));
  OAI21_X1   g27939(.A1(new_n31180_), .A2(new_n24115_), .B(new_n31181_), .ZN(po0715));
  INV_X1     g27940(.I(pi0559), .ZN(new_n31183_));
  NAND2_X1   g27941(.A1(new_n24077_), .A2(pi0241), .ZN(new_n31184_));
  OAI21_X1   g27942(.A1(new_n31183_), .A2(new_n24077_), .B(new_n31184_), .ZN(po0716));
  INV_X1     g27943(.I(pi0560), .ZN(new_n31186_));
  NAND2_X1   g27944(.A1(new_n24089_), .A2(pi0240), .ZN(new_n31187_));
  OAI21_X1   g27945(.A1(new_n31186_), .A2(new_n24089_), .B(new_n31187_), .ZN(po0717));
  INV_X1     g27946(.I(pi0561), .ZN(new_n31189_));
  NAND2_X1   g27947(.A1(new_n24083_), .A2(pi0247), .ZN(new_n31190_));
  OAI21_X1   g27948(.A1(new_n31189_), .A2(new_n24083_), .B(new_n31190_), .ZN(po0718));
  INV_X1     g27949(.I(pi0562), .ZN(new_n31192_));
  NAND2_X1   g27950(.A1(new_n24089_), .A2(pi0241), .ZN(new_n31193_));
  OAI21_X1   g27951(.A1(new_n31192_), .A2(new_n24089_), .B(new_n31193_), .ZN(po0719));
  INV_X1     g27952(.I(pi0563), .ZN(new_n31195_));
  NAND2_X1   g27953(.A1(new_n24931_), .A2(pi0246), .ZN(new_n31196_));
  OAI21_X1   g27954(.A1(new_n31195_), .A2(new_n24931_), .B(new_n31196_), .ZN(po0720));
  INV_X1     g27955(.I(pi0564), .ZN(new_n31198_));
  NAND2_X1   g27956(.A1(new_n24089_), .A2(pi0246), .ZN(new_n31199_));
  OAI21_X1   g27957(.A1(new_n31198_), .A2(new_n24089_), .B(new_n31199_), .ZN(po0721));
  INV_X1     g27958(.I(pi0565), .ZN(new_n31201_));
  NAND2_X1   g27959(.A1(new_n24089_), .A2(pi0248), .ZN(new_n31202_));
  OAI21_X1   g27960(.A1(new_n31201_), .A2(new_n24089_), .B(new_n31202_), .ZN(po0722));
  INV_X1     g27961(.I(pi0566), .ZN(new_n31204_));
  NAND2_X1   g27962(.A1(new_n24089_), .A2(pi0244), .ZN(new_n31205_));
  OAI21_X1   g27963(.A1(new_n31204_), .A2(new_n24089_), .B(new_n31205_), .ZN(po0723));
  NAND3_X1   g27964(.A1(new_n26307_), .A2(new_n6267_), .A3(pi1092), .ZN(new_n31207_));
  NOR3_X1    g27965(.A1(new_n2923_), .A2(pi0567), .A3(pi1093), .ZN(new_n31208_));
  NAND4_X1   g27966(.A1(new_n14637_), .A2(pi0603), .A3(new_n12307_), .A4(new_n14626_), .ZN(new_n31209_));
  NOR2_X1    g27967(.A1(new_n31209_), .A2(pi0619), .ZN(new_n31210_));
  OAI21_X1   g27968(.A1(new_n31210_), .A2(new_n31208_), .B(pi1159), .ZN(new_n31211_));
  NOR2_X1    g27969(.A1(new_n31208_), .A2(new_n11869_), .ZN(new_n31212_));
  OAI21_X1   g27970(.A1(new_n31209_), .A2(new_n11967_), .B(new_n31212_), .ZN(new_n31213_));
  AOI21_X1   g27971(.A1(new_n31211_), .A2(new_n31213_), .B(new_n11985_), .ZN(new_n31214_));
  INV_X1     g27972(.I(new_n31214_), .ZN(new_n31215_));
  INV_X1     g27973(.I(new_n31208_), .ZN(new_n31216_));
  NAND3_X1   g27974(.A1(new_n31209_), .A2(new_n11985_), .A3(new_n31216_), .ZN(new_n31217_));
  NAND2_X1   g27975(.A1(new_n31215_), .A2(new_n31217_), .ZN(new_n31218_));
  NOR3_X1    g27976(.A1(new_n2926_), .A2(new_n12223_), .A3(new_n5095_), .ZN(new_n31219_));
  AOI21_X1   g27977(.A1(new_n13637_), .A2(new_n31219_), .B(new_n31208_), .ZN(new_n31220_));
  INV_X1     g27978(.I(new_n31220_), .ZN(new_n31221_));
  NOR2_X1    g27979(.A1(new_n31221_), .A2(new_n13716_), .ZN(new_n31222_));
  OAI21_X1   g27980(.A1(new_n31215_), .A2(new_n12012_), .B(new_n31222_), .ZN(new_n31223_));
  AOI21_X1   g27981(.A1(new_n31223_), .A2(new_n31218_), .B(new_n11999_), .ZN(new_n31224_));
  NAND3_X1   g27982(.A1(new_n31215_), .A2(new_n24404_), .A3(new_n31217_), .ZN(new_n31225_));
  NOR3_X1    g27983(.A1(new_n31221_), .A2(new_n12013_), .A3(new_n13716_), .ZN(new_n31226_));
  NAND2_X1   g27984(.A1(new_n31226_), .A2(pi0641), .ZN(new_n31227_));
  NAND2_X1   g27985(.A1(new_n31227_), .A2(new_n31216_), .ZN(new_n31228_));
  NAND2_X1   g27986(.A1(new_n31226_), .A2(new_n11989_), .ZN(new_n31229_));
  NAND2_X1   g27987(.A1(new_n31229_), .A2(new_n31216_), .ZN(new_n31230_));
  AOI22_X1   g27988(.A1(new_n11993_), .A2(new_n31228_), .B1(new_n31230_), .B2(new_n11995_), .ZN(new_n31231_));
  AOI21_X1   g27989(.A1(new_n31225_), .A2(new_n31231_), .B(new_n11986_), .ZN(new_n31232_));
  OAI21_X1   g27990(.A1(new_n31232_), .A2(new_n31224_), .B(new_n14732_), .ZN(new_n31233_));
  NAND2_X1   g27991(.A1(new_n31218_), .A2(new_n14624_), .ZN(new_n31234_));
  OAI21_X1   g27992(.A1(new_n14624_), .A2(new_n31208_), .B(new_n31234_), .ZN(new_n31235_));
  NOR2_X1    g27993(.A1(new_n13717_), .A2(new_n31221_), .ZN(new_n31236_));
  INV_X1     g27994(.I(new_n31236_), .ZN(new_n31237_));
  OAI21_X1   g27995(.A1(new_n31237_), .A2(pi0628), .B(new_n31216_), .ZN(new_n31238_));
  NAND2_X1   g27996(.A1(new_n31238_), .A2(new_n12026_), .ZN(new_n31239_));
  NAND4_X1   g27997(.A1(new_n31235_), .A2(new_n12030_), .A3(new_n17150_), .A4(new_n31239_), .ZN(new_n31240_));
  NAND2_X1   g27998(.A1(new_n31235_), .A2(new_n16559_), .ZN(new_n31241_));
  OAI21_X1   g27999(.A1(new_n31237_), .A2(new_n12031_), .B(new_n31216_), .ZN(new_n31242_));
  NAND2_X1   g28000(.A1(new_n31242_), .A2(pi1156), .ZN(new_n31243_));
  NAND4_X1   g28001(.A1(new_n31240_), .A2(new_n12030_), .A3(new_n31241_), .A4(new_n31243_), .ZN(new_n31244_));
  NAND2_X1   g28002(.A1(new_n31244_), .A2(new_n11868_), .ZN(new_n31245_));
  NAND2_X1   g28003(.A1(new_n31245_), .A2(new_n31233_), .ZN(new_n31246_));
  NAND2_X1   g28004(.A1(new_n31246_), .A2(new_n12048_), .ZN(new_n31247_));
  INV_X1     g28005(.I(new_n31247_), .ZN(new_n31248_));
  INV_X1     g28006(.I(new_n31235_), .ZN(new_n31249_));
  NAND2_X1   g28007(.A1(new_n12053_), .A2(new_n31216_), .ZN(new_n31250_));
  OAI21_X1   g28008(.A1(new_n31249_), .A2(new_n12053_), .B(new_n31250_), .ZN(new_n31251_));
  XOR2_X1    g28009(.A1(new_n31246_), .A2(new_n31251_), .Z(new_n31252_));
  NAND2_X1   g28010(.A1(new_n31252_), .A2(pi0647), .ZN(new_n31253_));
  XNOR2_X1   g28011(.A1(new_n31253_), .A2(new_n31246_), .ZN(new_n31254_));
  NOR2_X1    g28012(.A1(new_n31237_), .A2(new_n12066_), .ZN(new_n31255_));
  NAND3_X1   g28013(.A1(new_n31255_), .A2(new_n13736_), .A3(new_n31216_), .ZN(new_n31256_));
  NAND2_X1   g28014(.A1(new_n31256_), .A2(new_n12060_), .ZN(new_n31257_));
  AOI21_X1   g28015(.A1(new_n31254_), .A2(new_n12049_), .B(new_n31257_), .ZN(new_n31258_));
  XOR2_X1    g28016(.A1(new_n31253_), .A2(new_n31251_), .Z(new_n31259_));
  NAND2_X1   g28017(.A1(new_n31216_), .A2(new_n12089_), .ZN(new_n31260_));
  AOI21_X1   g28018(.A1(new_n31255_), .A2(new_n12061_), .B(new_n31260_), .ZN(new_n31261_));
  OAI21_X1   g28019(.A1(new_n31259_), .A2(new_n12049_), .B(new_n31261_), .ZN(new_n31262_));
  NAND2_X1   g28020(.A1(new_n31262_), .A2(pi0787), .ZN(new_n31263_));
  NOR2_X1    g28021(.A1(new_n31258_), .A2(new_n31263_), .ZN(new_n31264_));
  NOR2_X1    g28022(.A1(new_n31264_), .A2(new_n31248_), .ZN(new_n31265_));
  INV_X1     g28023(.I(new_n31265_), .ZN(new_n31266_));
  NOR2_X1    g28024(.A1(new_n31266_), .A2(new_n12082_), .ZN(new_n31267_));
  AOI21_X1   g28025(.A1(new_n31255_), .A2(new_n13748_), .B(new_n31208_), .ZN(new_n31268_));
  OAI21_X1   g28026(.A1(new_n31268_), .A2(pi0644), .B(new_n12099_), .ZN(new_n31269_));
  NAND2_X1   g28027(.A1(new_n31249_), .A2(new_n16840_), .ZN(new_n31270_));
  OAI21_X1   g28028(.A1(new_n31270_), .A2(new_n12082_), .B(new_n31216_), .ZN(new_n31271_));
  AOI21_X1   g28029(.A1(new_n31271_), .A2(new_n12099_), .B(new_n12081_), .ZN(new_n31272_));
  OAI21_X1   g28030(.A1(new_n31267_), .A2(new_n31269_), .B(new_n31272_), .ZN(new_n31273_));
  NAND2_X1   g28031(.A1(new_n31216_), .A2(new_n14739_), .ZN(new_n31274_));
  INV_X1     g28032(.I(new_n31268_), .ZN(new_n31275_));
  MUX2_X1    g28033(.I0(new_n31275_), .I1(new_n31265_), .S(new_n12082_), .Z(new_n31276_));
  OAI22_X1   g28034(.A1(new_n31276_), .A2(pi0715), .B1(new_n31270_), .B2(new_n31274_), .ZN(new_n31277_));
  NAND2_X1   g28035(.A1(new_n31277_), .A2(new_n12081_), .ZN(new_n31278_));
  NAND2_X1   g28036(.A1(new_n31278_), .A2(new_n31273_), .ZN(new_n31279_));
  OAI21_X1   g28037(.A1(new_n31279_), .A2(new_n11867_), .B(new_n31266_), .ZN(new_n31280_));
  NAND3_X1   g28038(.A1(new_n31279_), .A2(pi0790), .A3(new_n31265_), .ZN(new_n31281_));
  NAND3_X1   g28039(.A1(new_n31280_), .A2(new_n31281_), .A3(pi0230), .ZN(new_n31282_));
  XOR2_X1    g28040(.A1(new_n31282_), .A2(new_n31207_), .Z(po0724));
  INV_X1     g28041(.I(pi0568), .ZN(new_n31284_));
  NAND2_X1   g28042(.A1(new_n24089_), .A2(pi0245), .ZN(new_n31285_));
  OAI21_X1   g28043(.A1(new_n31284_), .A2(new_n24089_), .B(new_n31285_), .ZN(po0725));
  NAND2_X1   g28044(.A1(new_n24089_), .A2(pi0239), .ZN(new_n31287_));
  OAI21_X1   g28045(.A1(pi0569), .A2(new_n24089_), .B(new_n31287_), .ZN(po0726));
  INV_X1     g28046(.I(pi0570), .ZN(new_n31289_));
  NAND3_X1   g28047(.A1(new_n31060_), .A2(new_n31289_), .A3(new_n24086_), .ZN(new_n31290_));
  NAND2_X1   g28048(.A1(new_n24089_), .A2(new_n31289_), .ZN(new_n31291_));
  OAI21_X1   g28049(.A1(new_n31039_), .A2(new_n31291_), .B(new_n31290_), .ZN(po0727));
  INV_X1     g28050(.I(pi0571), .ZN(new_n31293_));
  NAND2_X1   g28051(.A1(new_n24947_), .A2(pi0241), .ZN(new_n31294_));
  OAI21_X1   g28052(.A1(new_n31293_), .A2(new_n24947_), .B(new_n31294_), .ZN(po0728));
  INV_X1     g28053(.I(pi0572), .ZN(new_n31296_));
  NAND2_X1   g28054(.A1(new_n24947_), .A2(pi0244), .ZN(new_n31297_));
  OAI21_X1   g28055(.A1(new_n31296_), .A2(new_n24947_), .B(new_n31297_), .ZN(po0729));
  INV_X1     g28056(.I(pi0573), .ZN(new_n31299_));
  NAND2_X1   g28057(.A1(new_n24947_), .A2(pi0242), .ZN(new_n31300_));
  OAI21_X1   g28058(.A1(new_n31299_), .A2(new_n24947_), .B(new_n31300_), .ZN(po0730));
  INV_X1     g28059(.I(pi0574), .ZN(new_n31302_));
  NAND2_X1   g28060(.A1(new_n24083_), .A2(pi0241), .ZN(new_n31303_));
  OAI21_X1   g28061(.A1(new_n31302_), .A2(new_n24083_), .B(new_n31303_), .ZN(po0731));
  INV_X1     g28062(.I(pi0575), .ZN(new_n31305_));
  NAND2_X1   g28063(.A1(new_n24947_), .A2(pi0235), .ZN(new_n31306_));
  OAI21_X1   g28064(.A1(new_n31305_), .A2(new_n24947_), .B(new_n31306_), .ZN(po0732));
  INV_X1     g28065(.I(pi0576), .ZN(new_n31308_));
  NAND2_X1   g28066(.A1(new_n24947_), .A2(pi0248), .ZN(new_n31309_));
  OAI21_X1   g28067(.A1(new_n31308_), .A2(new_n24947_), .B(new_n31309_), .ZN(po0733));
  INV_X1     g28068(.I(pi0577), .ZN(new_n31311_));
  NAND2_X1   g28069(.A1(new_n24931_), .A2(pi0238), .ZN(new_n31312_));
  OAI21_X1   g28070(.A1(new_n31311_), .A2(new_n24931_), .B(new_n31312_), .ZN(po0734));
  INV_X1     g28071(.I(pi0578), .ZN(new_n31314_));
  NAND2_X1   g28072(.A1(new_n24083_), .A2(pi0249), .ZN(new_n31315_));
  OAI21_X1   g28073(.A1(new_n31314_), .A2(new_n24083_), .B(new_n31315_), .ZN(po0735));
  INV_X1     g28074(.I(pi0579), .ZN(new_n31317_));
  NAND2_X1   g28075(.A1(new_n24077_), .A2(pi0249), .ZN(new_n31318_));
  OAI21_X1   g28076(.A1(new_n31317_), .A2(new_n24077_), .B(new_n31318_), .ZN(po0736));
  INV_X1     g28077(.I(pi0580), .ZN(new_n31320_));
  NAND2_X1   g28078(.A1(new_n24931_), .A2(pi0245), .ZN(new_n31321_));
  OAI21_X1   g28079(.A1(new_n31320_), .A2(new_n24931_), .B(new_n31321_), .ZN(po0737));
  INV_X1     g28080(.I(pi0581), .ZN(new_n31323_));
  NAND2_X1   g28081(.A1(new_n24083_), .A2(pi0235), .ZN(new_n31324_));
  OAI21_X1   g28082(.A1(new_n31323_), .A2(new_n24083_), .B(new_n31324_), .ZN(po0738));
  INV_X1     g28083(.I(pi0582), .ZN(new_n31326_));
  NAND2_X1   g28084(.A1(new_n24083_), .A2(pi0240), .ZN(new_n31327_));
  OAI21_X1   g28085(.A1(new_n31326_), .A2(new_n24083_), .B(new_n31327_), .ZN(po0739));
  INV_X1     g28086(.I(pi0584), .ZN(new_n31329_));
  NAND2_X1   g28087(.A1(new_n24083_), .A2(pi0245), .ZN(new_n31330_));
  OAI21_X1   g28088(.A1(new_n31329_), .A2(new_n24083_), .B(new_n31330_), .ZN(po0741));
  INV_X1     g28089(.I(pi0585), .ZN(new_n31332_));
  NAND2_X1   g28090(.A1(new_n24083_), .A2(pi0244), .ZN(new_n31333_));
  OAI21_X1   g28091(.A1(new_n31332_), .A2(new_n24083_), .B(new_n31333_), .ZN(po0742));
  INV_X1     g28092(.I(pi0586), .ZN(new_n31335_));
  NAND2_X1   g28093(.A1(new_n24083_), .A2(pi0242), .ZN(new_n31336_));
  OAI21_X1   g28094(.A1(new_n31335_), .A2(new_n24083_), .B(new_n31336_), .ZN(po0743));
  NOR3_X1    g28095(.A1(new_n11997_), .A2(new_n11875_), .A3(new_n26307_), .ZN(new_n31338_));
  NAND4_X1   g28096(.A1(new_n31338_), .A2(new_n16840_), .A3(new_n14626_), .A4(new_n24570_), .ZN(new_n31339_));
  OAI22_X1   g28097(.A1(new_n14644_), .A2(new_n31339_), .B1(pi0230), .B2(new_n5468_), .ZN(po0744));
  NOR3_X1    g28098(.A1(new_n5366_), .A2(new_n2928_), .A3(pi0123), .ZN(new_n31341_));
  NAND3_X1   g28099(.A1(new_n31341_), .A2(new_n6711_), .A3(pi0591), .ZN(new_n31342_));
  INV_X1     g28100(.I(new_n31341_), .ZN(new_n31343_));
  OAI21_X1   g28101(.A1(new_n31343_), .A2(pi0591), .B(pi0588), .ZN(new_n31344_));
  AOI21_X1   g28102(.A1(new_n31344_), .A2(new_n31342_), .B(new_n30550_), .ZN(po0745));
  NOR2_X1    g28103(.A1(new_n31015_), .A2(pi0218), .ZN(new_n31346_));
  OAI21_X1   g28104(.A1(new_n31037_), .A2(pi0203), .B(new_n24069_), .ZN(new_n31347_));
  NOR2_X1    g28105(.A1(new_n31346_), .A2(new_n31347_), .ZN(new_n31348_));
  AOI21_X1   g28106(.A1(new_n31038_), .A2(new_n24945_), .B(new_n24069_), .ZN(new_n31349_));
  NOR3_X1    g28107(.A1(new_n31349_), .A2(new_n31015_), .A3(pi0206), .ZN(new_n31350_));
  OAI21_X1   g28108(.A1(new_n31348_), .A2(new_n31350_), .B(new_n24070_), .ZN(new_n31351_));
  NOR2_X1    g28109(.A1(new_n31015_), .A2(pi0205), .ZN(new_n31352_));
  OAI21_X1   g28110(.A1(new_n31037_), .A2(pi0202), .B(new_n24069_), .ZN(new_n31353_));
  NOR2_X1    g28111(.A1(new_n31352_), .A2(new_n31353_), .ZN(new_n31354_));
  AOI21_X1   g28112(.A1(new_n31038_), .A2(new_n24048_), .B(new_n24069_), .ZN(new_n31355_));
  NOR3_X1    g28113(.A1(new_n31355_), .A2(new_n31015_), .A3(pi0204), .ZN(new_n31356_));
  OAI21_X1   g28114(.A1(new_n31354_), .A2(new_n31356_), .B(pi0237), .ZN(new_n31357_));
  NAND2_X1   g28115(.A1(new_n31351_), .A2(new_n31357_), .ZN(po0746));
  OAI21_X1   g28116(.A1(pi0588), .A2(new_n31343_), .B(new_n30550_), .ZN(new_n31359_));
  AOI21_X1   g28117(.A1(new_n6203_), .A2(new_n31343_), .B(new_n31359_), .ZN(po0747));
  NAND3_X1   g28118(.A1(new_n31341_), .A2(new_n5940_), .A3(pi0592), .ZN(new_n31361_));
  OAI21_X1   g28119(.A1(new_n31343_), .A2(pi0592), .B(pi0591), .ZN(new_n31362_));
  AOI21_X1   g28120(.A1(new_n31362_), .A2(new_n31361_), .B(new_n30550_), .ZN(po0748));
  NAND3_X1   g28121(.A1(new_n31341_), .A2(pi0590), .A3(new_n6084_), .ZN(new_n31364_));
  OAI21_X1   g28122(.A1(new_n31343_), .A2(pi0590), .B(pi0592), .ZN(new_n31365_));
  AOI21_X1   g28123(.A1(new_n31365_), .A2(new_n31364_), .B(new_n30550_), .ZN(po0749));
  INV_X1     g28124(.I(pi0497), .ZN(new_n31367_));
  INV_X1     g28125(.I(pi0240), .ZN(new_n31368_));
  NOR2_X1    g28126(.A1(new_n31302_), .A2(pi0241), .ZN(new_n31369_));
  INV_X1     g28127(.I(pi0241), .ZN(new_n31370_));
  NOR2_X1    g28128(.A1(new_n31370_), .A2(pi0574), .ZN(new_n31371_));
  NOR2_X1    g28129(.A1(new_n31314_), .A2(pi0249), .ZN(new_n31372_));
  NOR2_X1    g28130(.A1(new_n3828_), .A2(pi0578), .ZN(new_n31373_));
  NOR4_X1    g28131(.A1(new_n31369_), .A2(new_n31371_), .A3(new_n31372_), .A4(new_n31373_), .ZN(new_n31374_));
  NOR2_X1    g28132(.A1(new_n31066_), .A2(pi0246), .ZN(new_n31375_));
  INV_X1     g28133(.I(pi0246), .ZN(new_n31376_));
  NOR2_X1    g28134(.A1(new_n31376_), .A2(pi0520), .ZN(new_n31377_));
  NOR2_X1    g28135(.A1(new_n31069_), .A2(pi0248), .ZN(new_n31378_));
  INV_X1     g28136(.I(pi0248), .ZN(new_n31379_));
  NOR2_X1    g28137(.A1(new_n31379_), .A2(pi0521), .ZN(new_n31380_));
  NOR4_X1    g28138(.A1(new_n31375_), .A2(new_n31377_), .A3(new_n31378_), .A4(new_n31380_), .ZN(new_n31381_));
  NOR2_X1    g28139(.A1(new_n31059_), .A2(pi0234), .ZN(new_n31382_));
  NOR2_X1    g28140(.A1(new_n2440_), .A2(pi0518), .ZN(new_n31383_));
  NOR4_X1    g28141(.A1(new_n31374_), .A2(new_n31381_), .A3(new_n31382_), .A4(new_n31383_), .ZN(new_n31384_));
  NAND2_X1   g28142(.A1(new_n31038_), .A2(new_n31384_), .ZN(new_n31385_));
  NOR2_X1    g28143(.A1(new_n30992_), .A2(pi0246), .ZN(new_n31386_));
  NOR2_X1    g28144(.A1(new_n31376_), .A2(pi0499), .ZN(new_n31387_));
  NOR2_X1    g28145(.A1(new_n3828_), .A2(pi0496), .ZN(new_n31388_));
  NOR2_X1    g28146(.A1(new_n30984_), .A2(pi0249), .ZN(new_n31389_));
  NOR4_X1    g28147(.A1(new_n31386_), .A2(new_n31387_), .A3(new_n31388_), .A4(new_n31389_), .ZN(new_n31390_));
  XOR2_X1    g28148(.A1(pi0248), .A2(pi0501), .Z(new_n31391_));
  NOR2_X1    g28149(.A1(new_n31010_), .A2(pi0234), .ZN(new_n31392_));
  NOR2_X1    g28150(.A1(new_n2440_), .A2(pi0505), .ZN(new_n31393_));
  NOR4_X1    g28151(.A1(new_n31390_), .A2(new_n31391_), .A3(new_n31392_), .A4(new_n31393_), .ZN(new_n31394_));
  NAND2_X1   g28152(.A1(new_n31016_), .A2(new_n31394_), .ZN(new_n31395_));
  INV_X1     g28153(.I(new_n31395_), .ZN(new_n31396_));
  XNOR2_X1   g28154(.A1(pi0241), .A2(pi0500), .ZN(new_n31397_));
  OAI21_X1   g28155(.A1(new_n31396_), .A2(new_n31397_), .B(new_n31385_), .ZN(new_n31398_));
  OAI21_X1   g28156(.A1(new_n31398_), .A2(pi0582), .B(new_n31368_), .ZN(new_n31399_));
  XOR2_X1    g28157(.A1(pi0241), .A2(pi0500), .Z(new_n31400_));
  NOR2_X1    g28158(.A1(new_n31395_), .A2(new_n31400_), .ZN(new_n31401_));
  NAND3_X1   g28159(.A1(new_n31399_), .A2(pi0582), .A3(new_n31401_), .ZN(new_n31402_));
  NAND4_X1   g28160(.A1(new_n31038_), .A2(new_n31368_), .A3(pi0582), .A4(new_n31384_), .ZN(new_n31403_));
  AOI21_X1   g28161(.A1(new_n31402_), .A2(new_n31403_), .B(pi0542), .ZN(new_n31404_));
  MUX2_X1    g28162(.I0(new_n31401_), .I1(new_n31398_), .S(new_n31326_), .Z(new_n31405_));
  OAI21_X1   g28163(.A1(new_n31385_), .A2(pi0582), .B(new_n31368_), .ZN(new_n31406_));
  NAND2_X1   g28164(.A1(new_n31406_), .A2(pi0542), .ZN(new_n31407_));
  AOI21_X1   g28165(.A1(new_n31405_), .A2(new_n31368_), .B(new_n31407_), .ZN(new_n31408_));
  NOR2_X1    g28166(.A1(new_n31404_), .A2(new_n31408_), .ZN(new_n31409_));
  XOR2_X1    g28167(.A1(pi0240), .A2(pi0582), .Z(new_n31410_));
  NOR2_X1    g28168(.A1(new_n31385_), .A2(new_n31410_), .ZN(new_n31411_));
  INV_X1     g28169(.I(new_n31411_), .ZN(new_n31412_));
  AOI21_X1   g28170(.A1(new_n31367_), .A2(new_n31412_), .B(new_n31409_), .ZN(new_n31413_));
  NAND3_X1   g28171(.A1(new_n31409_), .A2(new_n31367_), .A3(new_n31411_), .ZN(new_n31414_));
  XOR2_X1    g28172(.A1(pi0240), .A2(pi0542), .Z(new_n31415_));
  NOR3_X1    g28173(.A1(new_n31395_), .A2(new_n31400_), .A3(new_n31415_), .ZN(new_n31416_));
  AOI21_X1   g28174(.A1(new_n31416_), .A2(new_n31367_), .B(pi0239), .ZN(new_n31417_));
  NAND2_X1   g28175(.A1(new_n31414_), .A2(new_n31417_), .ZN(new_n31418_));
  OAI21_X1   g28176(.A1(new_n31418_), .A2(new_n31413_), .B(pi0519), .ZN(new_n31419_));
  NAND4_X1   g28177(.A1(new_n31409_), .A2(new_n3409_), .A3(pi0497), .A4(new_n31412_), .ZN(new_n31420_));
  NAND2_X1   g28178(.A1(new_n31416_), .A2(pi0497), .ZN(new_n31421_));
  AOI21_X1   g28179(.A1(new_n31421_), .A2(new_n3409_), .B(pi0519), .ZN(new_n31422_));
  AOI21_X1   g28180(.A1(new_n31420_), .A2(new_n31422_), .B(new_n31122_), .ZN(new_n31423_));
  NAND2_X1   g28181(.A1(new_n31419_), .A2(new_n31423_), .ZN(new_n31424_));
  XNOR2_X1   g28182(.A1(pi0239), .A2(pi0519), .ZN(new_n31425_));
  NOR2_X1    g28183(.A1(new_n31412_), .A2(new_n31425_), .ZN(new_n31426_));
  INV_X1     g28184(.I(new_n31426_), .ZN(new_n31427_));
  AOI21_X1   g28185(.A1(new_n31427_), .A2(new_n31122_), .B(pi0242), .ZN(new_n31428_));
  XNOR2_X1   g28186(.A1(pi0239), .A2(pi0497), .ZN(new_n31429_));
  NOR4_X1    g28187(.A1(new_n31395_), .A2(new_n31400_), .A3(new_n31415_), .A4(new_n31429_), .ZN(new_n31430_));
  INV_X1     g28188(.I(new_n31430_), .ZN(new_n31431_));
  OAI21_X1   g28189(.A1(new_n31431_), .A2(pi0539), .B(new_n4929_), .ZN(new_n31432_));
  NAND2_X1   g28190(.A1(new_n31432_), .A2(pi0586), .ZN(new_n31433_));
  AOI21_X1   g28191(.A1(new_n31424_), .A2(new_n31428_), .B(new_n31433_), .ZN(new_n31434_));
  INV_X1     g28192(.I(new_n31424_), .ZN(new_n31435_));
  NAND3_X1   g28193(.A1(new_n31430_), .A2(new_n4929_), .A3(pi0539), .ZN(new_n31436_));
  AOI21_X1   g28194(.A1(new_n31426_), .A2(pi0539), .B(pi0242), .ZN(new_n31437_));
  NAND2_X1   g28195(.A1(new_n31436_), .A2(new_n31437_), .ZN(new_n31438_));
  OAI21_X1   g28196(.A1(new_n31435_), .A2(new_n31438_), .B(new_n31335_), .ZN(new_n31439_));
  NAND2_X1   g28197(.A1(new_n31439_), .A2(pi0540), .ZN(new_n31440_));
  NOR2_X1    g28198(.A1(new_n31440_), .A2(new_n31434_), .ZN(new_n31441_));
  XOR2_X1    g28199(.A1(pi0242), .A2(pi0586), .Z(new_n31442_));
  NOR2_X1    g28200(.A1(new_n31427_), .A2(new_n31442_), .ZN(new_n31443_));
  OAI21_X1   g28201(.A1(new_n31443_), .A2(pi0540), .B(new_n3511_), .ZN(new_n31444_));
  XOR2_X1    g28202(.A1(pi0242), .A2(pi0539), .Z(new_n31445_));
  NOR2_X1    g28203(.A1(new_n31431_), .A2(new_n31445_), .ZN(new_n31446_));
  NAND2_X1   g28204(.A1(new_n31446_), .A2(new_n31125_), .ZN(new_n31447_));
  AOI21_X1   g28205(.A1(new_n31447_), .A2(new_n3511_), .B(new_n31323_), .ZN(new_n31448_));
  OAI21_X1   g28206(.A1(new_n31441_), .A2(new_n31444_), .B(new_n31448_), .ZN(new_n31449_));
  NAND3_X1   g28207(.A1(new_n31446_), .A2(new_n3511_), .A3(pi0540), .ZN(new_n31450_));
  NAND2_X1   g28208(.A1(new_n31443_), .A2(pi0540), .ZN(new_n31451_));
  NAND3_X1   g28209(.A1(new_n31450_), .A2(new_n3511_), .A3(new_n31451_), .ZN(new_n31452_));
  OAI21_X1   g28210(.A1(new_n31441_), .A2(new_n31452_), .B(new_n31323_), .ZN(new_n31453_));
  NAND3_X1   g28211(.A1(new_n31449_), .A2(new_n31453_), .A3(pi0585), .ZN(new_n31454_));
  XOR2_X1    g28212(.A1(pi0235), .A2(pi0540), .Z(new_n31455_));
  NOR3_X1    g28213(.A1(new_n31431_), .A2(new_n31445_), .A3(new_n31455_), .ZN(new_n31456_));
  INV_X1     g28214(.I(new_n31456_), .ZN(new_n31457_));
  AOI21_X1   g28215(.A1(new_n31457_), .A2(new_n31332_), .B(pi0244), .ZN(new_n31458_));
  INV_X1     g28216(.I(new_n31443_), .ZN(new_n31459_));
  XOR2_X1    g28217(.A1(pi0235), .A2(pi0581), .Z(new_n31460_));
  NOR3_X1    g28218(.A1(new_n31459_), .A2(pi0585), .A3(new_n31460_), .ZN(new_n31461_));
  OAI21_X1   g28219(.A1(new_n31461_), .A2(pi0244), .B(pi0541), .ZN(new_n31462_));
  AOI21_X1   g28220(.A1(new_n31454_), .A2(new_n31458_), .B(new_n31462_), .ZN(new_n31463_));
  NAND2_X1   g28221(.A1(new_n31456_), .A2(pi0585), .ZN(new_n31464_));
  NOR2_X1    g28222(.A1(new_n31459_), .A2(new_n31460_), .ZN(new_n31465_));
  AOI21_X1   g28223(.A1(new_n31465_), .A2(pi0585), .B(pi0244), .ZN(new_n31466_));
  AND3_X2    g28224(.A1(new_n31454_), .A2(new_n31464_), .A3(new_n31466_), .Z(new_n31467_));
  NOR2_X1    g28225(.A1(new_n31467_), .A2(pi0541), .ZN(new_n31468_));
  OR3_X2     g28226(.A1(new_n31468_), .A2(new_n31329_), .A3(new_n31463_), .Z(new_n31469_));
  XOR2_X1    g28227(.A1(pi0244), .A2(pi0541), .Z(new_n31470_));
  NOR2_X1    g28228(.A1(new_n31457_), .A2(new_n31470_), .ZN(new_n31471_));
  XNOR2_X1   g28229(.A1(pi0244), .A2(pi0585), .ZN(new_n31472_));
  NAND2_X1   g28230(.A1(new_n31465_), .A2(new_n31472_), .ZN(new_n31473_));
  OAI21_X1   g28231(.A1(new_n31473_), .A2(new_n31329_), .B(new_n4693_), .ZN(new_n31474_));
  AOI21_X1   g28232(.A1(new_n31471_), .A2(pi0584), .B(new_n31474_), .ZN(new_n31475_));
  NAND2_X1   g28233(.A1(new_n31469_), .A2(new_n31475_), .ZN(new_n31476_));
  INV_X1     g28234(.I(new_n31471_), .ZN(new_n31477_));
  AOI21_X1   g28235(.A1(new_n31477_), .A2(new_n31329_), .B(pi0245), .ZN(new_n31478_));
  NAND2_X1   g28236(.A1(new_n31469_), .A2(new_n31478_), .ZN(new_n31479_));
  NAND3_X1   g28237(.A1(new_n31465_), .A2(new_n31329_), .A3(new_n31472_), .ZN(new_n31480_));
  AOI21_X1   g28238(.A1(new_n31480_), .A2(new_n4693_), .B(new_n31004_), .ZN(new_n31481_));
  AOI22_X1   g28239(.A1(new_n31004_), .A2(new_n31476_), .B1(new_n31479_), .B2(new_n31481_), .ZN(new_n31482_));
  XOR2_X1    g28240(.A1(pi0245), .A2(pi0584), .Z(new_n31483_));
  NOR2_X1    g28241(.A1(new_n31473_), .A2(new_n31483_), .ZN(new_n31484_));
  INV_X1     g28242(.I(new_n31484_), .ZN(new_n31485_));
  XOR2_X1    g28243(.A1(new_n31482_), .A2(new_n31485_), .Z(new_n31486_));
  NAND2_X1   g28244(.A1(new_n31486_), .A2(pi0502), .ZN(new_n31487_));
  XNOR2_X1   g28245(.A1(new_n31487_), .A2(new_n31482_), .ZN(new_n31488_));
  XOR2_X1    g28246(.A1(pi0245), .A2(pi0503), .Z(new_n31489_));
  NOR2_X1    g28247(.A1(new_n31477_), .A2(new_n31489_), .ZN(new_n31490_));
  NOR2_X1    g28248(.A1(new_n31189_), .A2(pi0502), .ZN(new_n31491_));
  AOI21_X1   g28249(.A1(new_n31490_), .A2(new_n31491_), .B(pi0247), .ZN(new_n31492_));
  OAI21_X1   g28250(.A1(new_n31488_), .A2(pi0561), .B(new_n31492_), .ZN(new_n31493_));
  XOR2_X1    g28251(.A1(new_n31487_), .A2(new_n31484_), .Z(new_n31494_));
  NAND4_X1   g28252(.A1(new_n31490_), .A2(new_n4258_), .A3(pi0502), .A4(new_n31189_), .ZN(new_n31495_));
  OAI21_X1   g28253(.A1(new_n31494_), .A2(new_n31189_), .B(new_n31495_), .ZN(new_n31496_));
  AND2_X2    g28254(.A1(new_n31493_), .A2(new_n31496_), .Z(new_n31497_));
  NAND2_X1   g28255(.A1(new_n31497_), .A2(pi0238), .ZN(new_n31498_));
  XOR2_X1    g28256(.A1(pi0247), .A2(pi0502), .Z(new_n31499_));
  NOR3_X1    g28257(.A1(new_n31477_), .A2(new_n31489_), .A3(new_n31499_), .ZN(new_n31500_));
  XOR2_X1    g28258(.A1(pi0247), .A2(pi0561), .Z(new_n31501_));
  NOR2_X1    g28259(.A1(new_n31485_), .A2(new_n31501_), .ZN(new_n31502_));
  OAI21_X1   g28260(.A1(new_n31502_), .A2(pi0238), .B(new_n31500_), .ZN(new_n31503_));
  INV_X1     g28261(.I(new_n31502_), .ZN(new_n31504_));
  OR3_X2     g28262(.A1(new_n31504_), .A2(pi0238), .A3(new_n31500_), .Z(new_n31505_));
  NAND4_X1   g28263(.A1(new_n31505_), .A2(new_n31072_), .A3(pi0543), .A4(new_n31503_), .ZN(new_n31506_));
  AOI21_X1   g28264(.A1(new_n31498_), .A2(pi0522), .B(new_n31506_), .ZN(new_n31507_));
  NAND2_X1   g28265(.A1(new_n31497_), .A2(new_n3647_), .ZN(new_n31508_));
  NAND3_X1   g28266(.A1(new_n31504_), .A2(pi0238), .A3(new_n31072_), .ZN(new_n31509_));
  OAI21_X1   g28267(.A1(new_n31509_), .A2(new_n31500_), .B(new_n31134_), .ZN(new_n31510_));
  AOI21_X1   g28268(.A1(new_n31508_), .A2(new_n31072_), .B(new_n31510_), .ZN(new_n31511_));
  NOR2_X1    g28269(.A1(new_n31507_), .A2(new_n31511_), .ZN(new_n31512_));
  XNOR2_X1   g28270(.A1(pi0246), .A2(pi0487), .ZN(new_n31513_));
  XNOR2_X1   g28271(.A1(pi0234), .A2(pi0511), .ZN(new_n31514_));
  AOI21_X1   g28272(.A1(new_n31038_), .A2(new_n31513_), .B(new_n31514_), .ZN(new_n31515_));
  INV_X1     g28273(.I(new_n31515_), .ZN(new_n31516_));
  XOR2_X1    g28274(.A1(pi0249), .A2(pi0579), .Z(new_n31517_));
  NOR2_X1    g28275(.A1(new_n31516_), .A2(new_n31517_), .ZN(new_n31518_));
  XNOR2_X1   g28276(.A1(pi0246), .A2(pi0536), .ZN(new_n31519_));
  XNOR2_X1   g28277(.A1(pi0234), .A2(pi0557), .ZN(new_n31520_));
  AOI21_X1   g28278(.A1(new_n31016_), .A2(new_n31519_), .B(new_n31520_), .ZN(new_n31521_));
  AOI21_X1   g28279(.A1(new_n31521_), .A2(new_n31119_), .B(pi0249), .ZN(new_n31522_));
  NOR3_X1    g28280(.A1(new_n31522_), .A2(new_n31317_), .A3(new_n31516_), .ZN(new_n31523_));
  XOR2_X1    g28281(.A1(pi0249), .A2(pi0538), .Z(new_n31524_));
  INV_X1     g28282(.I(new_n31524_), .ZN(new_n31525_));
  AND2_X2    g28283(.A1(new_n31521_), .A2(new_n31525_), .Z(new_n31526_));
  NOR2_X1    g28284(.A1(new_n31518_), .A2(new_n31317_), .ZN(new_n31527_));
  NOR3_X1    g28285(.A1(new_n31523_), .A2(new_n31526_), .A3(new_n31527_), .ZN(new_n31528_));
  NAND3_X1   g28286(.A1(new_n31518_), .A2(pi0248), .A3(pi0537), .ZN(new_n31529_));
  NAND3_X1   g28287(.A1(new_n31526_), .A2(new_n31379_), .A3(pi0537), .ZN(new_n31530_));
  AOI21_X1   g28288(.A1(new_n31530_), .A2(new_n31529_), .B(pi0481), .ZN(new_n31531_));
  NOR4_X1    g28289(.A1(new_n31528_), .A2(pi0248), .A3(new_n31116_), .A4(new_n31518_), .ZN(new_n31532_));
  AOI21_X1   g28290(.A1(new_n31526_), .A2(new_n31116_), .B(pi0248), .ZN(new_n31533_));
  NOR3_X1    g28291(.A1(new_n31532_), .A2(new_n30941_), .A3(new_n31533_), .ZN(new_n31534_));
  OR3_X2     g28292(.A1(new_n31534_), .A2(new_n31183_), .A3(new_n31531_), .Z(new_n31535_));
  INV_X1     g28293(.I(new_n31526_), .ZN(new_n31536_));
  XOR2_X1    g28294(.A1(pi0248), .A2(pi0537), .Z(new_n31537_));
  NOR2_X1    g28295(.A1(new_n31536_), .A2(new_n31537_), .ZN(new_n31538_));
  INV_X1     g28296(.I(new_n31538_), .ZN(new_n31539_));
  AOI21_X1   g28297(.A1(new_n31539_), .A2(new_n31183_), .B(pi0241), .ZN(new_n31540_));
  XOR2_X1    g28298(.A1(pi0248), .A2(pi0481), .Z(new_n31541_));
  NOR3_X1    g28299(.A1(new_n31516_), .A2(new_n31517_), .A3(new_n31541_), .ZN(new_n31542_));
  INV_X1     g28300(.I(new_n31542_), .ZN(new_n31543_));
  OAI21_X1   g28301(.A1(new_n31543_), .A2(pi0559), .B(new_n31370_), .ZN(new_n31544_));
  NAND2_X1   g28302(.A1(new_n31544_), .A2(pi0506), .ZN(new_n31545_));
  AOI21_X1   g28303(.A1(new_n31535_), .A2(new_n31540_), .B(new_n31545_), .ZN(new_n31546_));
  OAI21_X1   g28304(.A1(new_n31543_), .A2(new_n31183_), .B(new_n31370_), .ZN(new_n31547_));
  AOI21_X1   g28305(.A1(new_n31538_), .A2(pi0559), .B(new_n31547_), .ZN(new_n31548_));
  AOI21_X1   g28306(.A1(new_n31535_), .A2(new_n31548_), .B(pi0506), .ZN(new_n31549_));
  OR3_X2     g28307(.A1(new_n31546_), .A2(new_n31549_), .A3(new_n31050_), .Z(new_n31550_));
  XOR2_X1    g28308(.A1(pi0241), .A2(pi0506), .Z(new_n31551_));
  NOR2_X1    g28309(.A1(new_n31539_), .A2(new_n31551_), .ZN(new_n31552_));
  XOR2_X1    g28310(.A1(pi0241), .A2(pi0559), .Z(new_n31553_));
  NOR2_X1    g28311(.A1(new_n31543_), .A2(new_n31553_), .ZN(new_n31554_));
  INV_X1     g28312(.I(new_n31554_), .ZN(new_n31555_));
  OAI21_X1   g28313(.A1(new_n31555_), .A2(new_n31050_), .B(new_n31368_), .ZN(new_n31556_));
  AOI21_X1   g28314(.A1(new_n31552_), .A2(pi0515), .B(new_n31556_), .ZN(new_n31557_));
  AOI21_X1   g28315(.A1(new_n31550_), .A2(new_n31557_), .B(pi0535), .ZN(new_n31558_));
  INV_X1     g28316(.I(new_n31552_), .ZN(new_n31559_));
  AOI21_X1   g28317(.A1(new_n31559_), .A2(new_n31050_), .B(pi0240), .ZN(new_n31560_));
  OAI21_X1   g28318(.A1(new_n31555_), .A2(pi0515), .B(new_n31368_), .ZN(new_n31561_));
  NAND2_X1   g28319(.A1(new_n31561_), .A2(pi0535), .ZN(new_n31562_));
  AOI21_X1   g28320(.A1(new_n31550_), .A2(new_n31560_), .B(new_n31562_), .ZN(new_n31563_));
  NOR2_X1    g28321(.A1(new_n31558_), .A2(new_n31563_), .ZN(new_n31564_));
  INV_X1     g28322(.I(new_n31564_), .ZN(new_n31565_));
  XOR2_X1    g28323(.A1(pi0240), .A2(pi0515), .Z(new_n31566_));
  NOR2_X1    g28324(.A1(new_n31555_), .A2(new_n31566_), .ZN(new_n31567_));
  OAI21_X1   g28325(.A1(pi0534), .A2(new_n31567_), .B(new_n31565_), .ZN(new_n31568_));
  INV_X1     g28326(.I(pi0534), .ZN(new_n31569_));
  NAND3_X1   g28327(.A1(new_n31564_), .A2(new_n31569_), .A3(new_n31567_), .ZN(new_n31570_));
  XOR2_X1    g28328(.A1(pi0240), .A2(pi0535), .Z(new_n31571_));
  NOR2_X1    g28329(.A1(new_n31559_), .A2(new_n31571_), .ZN(new_n31572_));
  AOI21_X1   g28330(.A1(new_n31572_), .A2(new_n31569_), .B(pi0239), .ZN(new_n31573_));
  NAND3_X1   g28331(.A1(new_n31568_), .A2(new_n31570_), .A3(new_n31573_), .ZN(new_n31574_));
  NOR4_X1    g28332(.A1(new_n31565_), .A2(pi0239), .A3(new_n31569_), .A4(new_n31567_), .ZN(new_n31575_));
  AOI21_X1   g28333(.A1(new_n31572_), .A2(pi0534), .B(pi0239), .ZN(new_n31576_));
  OR2_X2     g28334(.A1(new_n31576_), .A2(pi0488), .Z(new_n31577_));
  OAI21_X1   g28335(.A1(new_n31575_), .A2(new_n31577_), .B(pi0504), .ZN(new_n31578_));
  AOI21_X1   g28336(.A1(pi0488), .A2(new_n31574_), .B(new_n31578_), .ZN(new_n31579_));
  XNOR2_X1   g28337(.A1(pi0239), .A2(pi0488), .ZN(new_n31580_));
  NOR3_X1    g28338(.A1(new_n31555_), .A2(new_n31566_), .A3(new_n31580_), .ZN(new_n31581_));
  OAI21_X1   g28339(.A1(new_n31581_), .A2(pi0504), .B(new_n4929_), .ZN(new_n31582_));
  XNOR2_X1   g28340(.A1(pi0239), .A2(pi0534), .ZN(new_n31583_));
  NOR3_X1    g28341(.A1(new_n31559_), .A2(new_n31571_), .A3(new_n31583_), .ZN(new_n31584_));
  NAND2_X1   g28342(.A1(new_n31584_), .A2(new_n31007_), .ZN(new_n31585_));
  AOI21_X1   g28343(.A1(new_n31585_), .A2(new_n4929_), .B(new_n31032_), .ZN(new_n31586_));
  OAI21_X1   g28344(.A1(new_n31579_), .A2(new_n31582_), .B(new_n31586_), .ZN(new_n31587_));
  NAND3_X1   g28345(.A1(new_n31584_), .A2(new_n4929_), .A3(pi0504), .ZN(new_n31588_));
  AOI21_X1   g28346(.A1(new_n31581_), .A2(pi0504), .B(pi0242), .ZN(new_n31589_));
  NAND2_X1   g28347(.A1(new_n31588_), .A2(new_n31589_), .ZN(new_n31590_));
  OAI21_X1   g28348(.A1(new_n31579_), .A2(new_n31590_), .B(new_n31032_), .ZN(new_n31591_));
  NAND3_X1   g28349(.A1(new_n31587_), .A2(new_n31591_), .A3(pi0533), .ZN(new_n31592_));
  XNOR2_X1   g28350(.A1(pi0242), .A2(pi0510), .ZN(new_n31593_));
  NAND2_X1   g28351(.A1(new_n31581_), .A2(new_n31593_), .ZN(new_n31594_));
  AOI21_X1   g28352(.A1(new_n31594_), .A2(new_n31105_), .B(pi0235), .ZN(new_n31595_));
  XNOR2_X1   g28353(.A1(pi0242), .A2(pi0504), .ZN(new_n31596_));
  NAND2_X1   g28354(.A1(new_n31584_), .A2(new_n31596_), .ZN(new_n31597_));
  OAI21_X1   g28355(.A1(new_n31597_), .A2(pi0533), .B(new_n3511_), .ZN(new_n31598_));
  NAND2_X1   g28356(.A1(new_n31598_), .A2(pi0512), .ZN(new_n31599_));
  AOI21_X1   g28357(.A1(new_n31592_), .A2(new_n31595_), .B(new_n31599_), .ZN(new_n31600_));
  NOR3_X1    g28358(.A1(new_n31597_), .A2(pi0235), .A3(new_n31105_), .ZN(new_n31601_));
  OAI21_X1   g28359(.A1(new_n31594_), .A2(new_n31105_), .B(new_n3511_), .ZN(new_n31602_));
  NOR2_X1    g28360(.A1(new_n31601_), .A2(new_n31602_), .ZN(new_n31603_));
  AOI21_X1   g28361(.A1(new_n31592_), .A2(new_n31603_), .B(pi0512), .ZN(new_n31604_));
  NOR3_X1    g28362(.A1(new_n31600_), .A2(new_n31604_), .A3(new_n31180_), .ZN(new_n31605_));
  XOR2_X1    g28363(.A1(pi0235), .A2(pi0512), .Z(new_n31606_));
  NOR2_X1    g28364(.A1(new_n31594_), .A2(new_n31606_), .ZN(new_n31607_));
  OAI21_X1   g28365(.A1(new_n31607_), .A2(pi0558), .B(new_n4842_), .ZN(new_n31608_));
  XOR2_X1    g28366(.A1(pi0235), .A2(pi0533), .Z(new_n31609_));
  NOR2_X1    g28367(.A1(new_n31597_), .A2(new_n31609_), .ZN(new_n31610_));
  NAND2_X1   g28368(.A1(new_n31610_), .A2(new_n31180_), .ZN(new_n31611_));
  AOI21_X1   g28369(.A1(new_n31611_), .A2(new_n4842_), .B(new_n31044_), .ZN(new_n31612_));
  OAI21_X1   g28370(.A1(new_n31605_), .A2(new_n31608_), .B(new_n31612_), .ZN(new_n31613_));
  NAND3_X1   g28371(.A1(new_n31610_), .A2(new_n4842_), .A3(pi0558), .ZN(new_n31614_));
  AOI21_X1   g28372(.A1(new_n31607_), .A2(pi0558), .B(pi0244), .ZN(new_n31615_));
  NAND2_X1   g28373(.A1(new_n31614_), .A2(new_n31615_), .ZN(new_n31616_));
  OAI21_X1   g28374(.A1(new_n31605_), .A2(new_n31616_), .B(new_n31044_), .ZN(new_n31617_));
  NAND3_X1   g28375(.A1(new_n31613_), .A2(new_n31617_), .A3(pi0509), .ZN(new_n31618_));
  XNOR2_X1   g28376(.A1(pi0244), .A2(pi0513), .ZN(new_n31619_));
  NAND2_X1   g28377(.A1(new_n31607_), .A2(new_n31619_), .ZN(new_n31620_));
  AOI21_X1   g28378(.A1(new_n31620_), .A2(new_n31029_), .B(pi0245), .ZN(new_n31621_));
  XNOR2_X1   g28379(.A1(pi0244), .A2(pi0558), .ZN(new_n31622_));
  NAND2_X1   g28380(.A1(new_n31610_), .A2(new_n31622_), .ZN(new_n31623_));
  OAI21_X1   g28381(.A1(new_n31623_), .A2(pi0509), .B(new_n4693_), .ZN(new_n31624_));
  NAND2_X1   g28382(.A1(new_n31624_), .A2(pi0514), .ZN(new_n31625_));
  AOI21_X1   g28383(.A1(new_n31618_), .A2(new_n31621_), .B(new_n31625_), .ZN(new_n31626_));
  NAND4_X1   g28384(.A1(new_n31610_), .A2(new_n4693_), .A3(pi0509), .A4(new_n31622_), .ZN(new_n31627_));
  INV_X1     g28385(.I(new_n31620_), .ZN(new_n31628_));
  AOI21_X1   g28386(.A1(new_n31628_), .A2(pi0509), .B(pi0245), .ZN(new_n31629_));
  AND3_X2    g28387(.A1(new_n31618_), .A2(new_n31627_), .A3(new_n31629_), .Z(new_n31630_));
  OAI21_X1   g28388(.A1(new_n31630_), .A2(pi0514), .B(pi0508), .ZN(new_n31631_));
  NOR2_X1    g28389(.A1(new_n31631_), .A2(new_n31626_), .ZN(new_n31632_));
  INV_X1     g28390(.I(new_n31632_), .ZN(new_n31633_));
  XOR2_X1    g28391(.A1(pi0245), .A2(pi0509), .Z(new_n31634_));
  NOR2_X1    g28392(.A1(new_n31623_), .A2(new_n31634_), .ZN(new_n31635_));
  NAND3_X1   g28393(.A1(new_n31635_), .A2(new_n4258_), .A3(pi0508), .ZN(new_n31636_));
  XOR2_X1    g28394(.A1(pi0245), .A2(pi0514), .Z(new_n31637_));
  NOR2_X1    g28395(.A1(new_n31620_), .A2(new_n31637_), .ZN(new_n31638_));
  NAND2_X1   g28396(.A1(new_n31638_), .A2(pi0508), .ZN(new_n31639_));
  NAND4_X1   g28397(.A1(new_n31633_), .A2(new_n4258_), .A3(new_n31636_), .A4(new_n31639_), .ZN(new_n31640_));
  NOR2_X1    g28398(.A1(new_n31638_), .A2(pi0508), .ZN(new_n31641_));
  OR3_X2     g28399(.A1(new_n31632_), .A2(pi0247), .A3(new_n31641_), .Z(new_n31642_));
  NAND2_X1   g28400(.A1(new_n31635_), .A2(new_n31026_), .ZN(new_n31643_));
  AOI21_X1   g28401(.A1(new_n31643_), .A2(new_n4258_), .B(new_n31053_), .ZN(new_n31644_));
  AOI22_X1   g28402(.A1(new_n31640_), .A2(new_n31053_), .B1(new_n31642_), .B2(new_n31644_), .ZN(new_n31645_));
  OAI21_X1   g28403(.A1(new_n31645_), .A2(new_n3647_), .B(pi0517), .ZN(new_n31646_));
  XNOR2_X1   g28404(.A1(pi0247), .A2(pi0508), .ZN(new_n31647_));
  NAND2_X1   g28405(.A1(new_n31635_), .A2(new_n31647_), .ZN(new_n31648_));
  XNOR2_X1   g28406(.A1(pi0247), .A2(pi0516), .ZN(new_n31649_));
  NAND2_X1   g28407(.A1(new_n31638_), .A2(new_n31649_), .ZN(new_n31650_));
  AOI21_X1   g28408(.A1(new_n3647_), .A2(new_n31650_), .B(new_n31648_), .ZN(new_n31651_));
  INV_X1     g28409(.I(new_n31648_), .ZN(new_n31652_));
  NOR3_X1    g28410(.A1(new_n31652_), .A2(pi0238), .A3(new_n31650_), .ZN(new_n31653_));
  NOR4_X1    g28411(.A1(new_n31653_), .A2(new_n31023_), .A3(pi0517), .A4(new_n31651_), .ZN(new_n31654_));
  OAI21_X1   g28412(.A1(new_n31645_), .A2(pi0238), .B(new_n31056_), .ZN(new_n31655_));
  NAND3_X1   g28413(.A1(new_n31638_), .A2(pi0238), .A3(new_n31649_), .ZN(new_n31656_));
  NOR3_X1    g28414(.A1(new_n31652_), .A2(new_n3647_), .A3(pi0517), .ZN(new_n31657_));
  AOI21_X1   g28415(.A1(new_n31657_), .A2(new_n31656_), .B(pi0507), .ZN(new_n31658_));
  AOI22_X1   g28416(.A1(new_n31646_), .A2(new_n31654_), .B1(new_n31655_), .B2(new_n31658_), .ZN(new_n31659_));
  MUX2_X1    g28417(.I0(new_n31659_), .I1(new_n31512_), .S(new_n24069_), .Z(new_n31660_));
  INV_X1     g28418(.I(pi0524), .ZN(new_n31661_));
  INV_X1     g28419(.I(pi0494), .ZN(new_n31662_));
  NOR2_X1    g28420(.A1(new_n31084_), .A2(pi0246), .ZN(new_n31663_));
  NOR2_X1    g28421(.A1(new_n31376_), .A2(pi0526), .ZN(new_n31664_));
  NOR2_X1    g28422(.A1(new_n31308_), .A2(pi0248), .ZN(new_n31665_));
  NOR2_X1    g28423(.A1(new_n31379_), .A2(pi0576), .ZN(new_n31666_));
  NOR4_X1    g28424(.A1(new_n31663_), .A2(new_n31664_), .A3(new_n31665_), .A4(new_n31666_), .ZN(new_n31667_));
  XOR2_X1    g28425(.A1(pi0249), .A2(pi0528), .Z(new_n31668_));
  NOR2_X1    g28426(.A1(new_n31075_), .A2(pi0234), .ZN(new_n31669_));
  NOR2_X1    g28427(.A1(new_n2440_), .A2(pi0523), .ZN(new_n31670_));
  NOR4_X1    g28428(.A1(new_n31667_), .A2(new_n31668_), .A3(new_n31669_), .A4(new_n31670_), .ZN(new_n31671_));
  NAND2_X1   g28429(.A1(new_n31038_), .A2(new_n31671_), .ZN(new_n31672_));
  INV_X1     g28430(.I(new_n31672_), .ZN(new_n31673_));
  XNOR2_X1   g28431(.A1(pi0241), .A2(pi0571), .ZN(new_n31674_));
  NOR2_X1    g28432(.A1(new_n31673_), .A2(new_n31674_), .ZN(new_n31675_));
  NOR2_X1    g28433(.A1(new_n31144_), .A2(pi0246), .ZN(new_n31676_));
  NOR2_X1    g28434(.A1(new_n31376_), .A2(pi0546), .ZN(new_n31677_));
  NOR2_X1    g28435(.A1(new_n31150_), .A2(pi0248), .ZN(new_n31678_));
  NOR2_X1    g28436(.A1(new_n31379_), .A2(pi0548), .ZN(new_n31679_));
  NOR4_X1    g28437(.A1(new_n31676_), .A2(new_n31677_), .A3(new_n31678_), .A4(new_n31679_), .ZN(new_n31680_));
  XOR2_X1    g28438(.A1(pi0249), .A2(pi0484), .Z(new_n31681_));
  NOR2_X1    g28439(.A1(new_n31137_), .A2(pi0234), .ZN(new_n31682_));
  NOR2_X1    g28440(.A1(new_n2440_), .A2(pi0544), .ZN(new_n31683_));
  NOR4_X1    g28441(.A1(new_n31680_), .A2(new_n31681_), .A3(new_n31682_), .A4(new_n31683_), .ZN(new_n31684_));
  NAND2_X1   g28442(.A1(new_n31016_), .A2(new_n31684_), .ZN(new_n31685_));
  AOI21_X1   g28443(.A1(pi0241), .A2(new_n31685_), .B(new_n31675_), .ZN(new_n31686_));
  OAI22_X1   g28444(.A1(new_n31685_), .A2(new_n31370_), .B1(new_n31673_), .B2(new_n31674_), .ZN(new_n31687_));
  NAND2_X1   g28445(.A1(new_n31687_), .A2(pi0490), .ZN(new_n31688_));
  OAI21_X1   g28446(.A1(new_n31686_), .A2(pi0490), .B(new_n31688_), .ZN(new_n31689_));
  XOR2_X1    g28447(.A1(pi0241), .A2(pi0490), .Z(new_n31690_));
  NOR2_X1    g28448(.A1(new_n31685_), .A2(new_n31690_), .ZN(new_n31691_));
  XOR2_X1    g28449(.A1(new_n31689_), .A2(new_n31691_), .Z(new_n31692_));
  NAND2_X1   g28450(.A1(new_n31692_), .A2(pi0530), .ZN(new_n31693_));
  XNOR2_X1   g28451(.A1(new_n31693_), .A2(new_n31689_), .ZN(new_n31694_));
  XOR2_X1    g28452(.A1(pi0241), .A2(pi0571), .Z(new_n31695_));
  NOR2_X1    g28453(.A1(new_n31672_), .A2(new_n31695_), .ZN(new_n31696_));
  INV_X1     g28454(.I(new_n31696_), .ZN(new_n31697_));
  NAND2_X1   g28455(.A1(new_n31096_), .A2(pi0492), .ZN(new_n31698_));
  OAI21_X1   g28456(.A1(new_n31697_), .A2(new_n31698_), .B(new_n31368_), .ZN(new_n31699_));
  AOI21_X1   g28457(.A1(new_n31694_), .A2(new_n30973_), .B(new_n31699_), .ZN(new_n31700_));
  INV_X1     g28458(.I(new_n31691_), .ZN(new_n31701_));
  XOR2_X1    g28459(.A1(new_n31693_), .A2(new_n31701_), .Z(new_n31702_));
  NOR4_X1    g28460(.A1(new_n31697_), .A2(pi0240), .A3(pi0492), .A4(new_n31096_), .ZN(new_n31703_));
  AOI21_X1   g28461(.A1(new_n31702_), .A2(pi0492), .B(new_n31703_), .ZN(new_n31704_));
  NOR2_X1    g28462(.A1(new_n31700_), .A2(new_n31704_), .ZN(new_n31705_));
  INV_X1     g28463(.I(new_n31705_), .ZN(new_n31706_));
  XNOR2_X1   g28464(.A1(pi0240), .A2(pi0530), .ZN(new_n31707_));
  NAND2_X1   g28465(.A1(new_n31696_), .A2(new_n31707_), .ZN(new_n31708_));
  AOI21_X1   g28466(.A1(new_n31662_), .A2(new_n31708_), .B(new_n31706_), .ZN(new_n31709_));
  NOR3_X1    g28467(.A1(new_n31705_), .A2(pi0494), .A3(new_n31708_), .ZN(new_n31710_));
  XOR2_X1    g28468(.A1(pi0240), .A2(pi0492), .Z(new_n31711_));
  NOR2_X1    g28469(.A1(new_n31701_), .A2(new_n31711_), .ZN(new_n31712_));
  INV_X1     g28470(.I(new_n31712_), .ZN(new_n31713_));
  OAI21_X1   g28471(.A1(new_n31713_), .A2(pi0494), .B(new_n3409_), .ZN(new_n31714_));
  NOR3_X1    g28472(.A1(new_n31709_), .A2(new_n31710_), .A3(new_n31714_), .ZN(new_n31715_));
  NAND4_X1   g28473(.A1(new_n31706_), .A2(new_n3409_), .A3(pi0494), .A4(new_n31708_), .ZN(new_n31716_));
  NAND2_X1   g28474(.A1(new_n31712_), .A2(pi0494), .ZN(new_n31717_));
  AOI21_X1   g28475(.A1(new_n31717_), .A2(new_n3409_), .B(pi0524), .ZN(new_n31718_));
  AOI21_X1   g28476(.A1(new_n31716_), .A2(new_n31718_), .B(new_n30947_), .ZN(new_n31719_));
  OAI21_X1   g28477(.A1(new_n31715_), .A2(new_n31661_), .B(new_n31719_), .ZN(new_n31720_));
  XOR2_X1    g28478(.A1(pi0239), .A2(pi0524), .Z(new_n31721_));
  NAND3_X1   g28479(.A1(new_n31696_), .A2(new_n31707_), .A3(new_n31721_), .ZN(new_n31722_));
  AOI21_X1   g28480(.A1(new_n31722_), .A2(new_n30947_), .B(pi0242), .ZN(new_n31723_));
  XNOR2_X1   g28481(.A1(pi0239), .A2(pi0494), .ZN(new_n31724_));
  NOR2_X1    g28482(.A1(new_n31713_), .A2(new_n31724_), .ZN(new_n31725_));
  INV_X1     g28483(.I(new_n31725_), .ZN(new_n31726_));
  OAI21_X1   g28484(.A1(new_n31726_), .A2(pi0483), .B(new_n4929_), .ZN(new_n31727_));
  NAND2_X1   g28485(.A1(new_n31727_), .A2(pi0573), .ZN(new_n31728_));
  AOI21_X1   g28486(.A1(new_n31720_), .A2(new_n31723_), .B(new_n31728_), .ZN(new_n31729_));
  NOR2_X1    g28487(.A1(new_n30947_), .A2(pi0242), .ZN(new_n31730_));
  OAI21_X1   g28488(.A1(new_n31722_), .A2(new_n30947_), .B(new_n4929_), .ZN(new_n31731_));
  AOI21_X1   g28489(.A1(new_n31725_), .A2(new_n31730_), .B(new_n31731_), .ZN(new_n31732_));
  AOI21_X1   g28490(.A1(new_n31720_), .A2(new_n31732_), .B(pi0573), .ZN(new_n31733_));
  NOR3_X1    g28491(.A1(new_n31729_), .A2(new_n31733_), .A3(new_n30981_), .ZN(new_n31734_));
  XOR2_X1    g28492(.A1(pi0242), .A2(pi0573), .Z(new_n31735_));
  NOR2_X1    g28493(.A1(new_n31722_), .A2(new_n31735_), .ZN(new_n31736_));
  OAI21_X1   g28494(.A1(new_n31736_), .A2(pi0495), .B(new_n3511_), .ZN(new_n31737_));
  XOR2_X1    g28495(.A1(pi0242), .A2(pi0483), .Z(new_n31738_));
  NOR2_X1    g28496(.A1(new_n31726_), .A2(new_n31738_), .ZN(new_n31739_));
  NAND2_X1   g28497(.A1(new_n31739_), .A2(new_n30981_), .ZN(new_n31740_));
  AOI21_X1   g28498(.A1(new_n31740_), .A2(new_n3511_), .B(new_n31305_), .ZN(new_n31741_));
  OAI21_X1   g28499(.A1(new_n31734_), .A2(new_n31737_), .B(new_n31741_), .ZN(new_n31742_));
  INV_X1     g28500(.I(new_n31739_), .ZN(new_n31743_));
  NAND2_X1   g28501(.A1(new_n3511_), .A2(pi0495), .ZN(new_n31744_));
  AOI21_X1   g28502(.A1(new_n31736_), .A2(pi0495), .B(pi0235), .ZN(new_n31745_));
  OAI21_X1   g28503(.A1(new_n31743_), .A2(new_n31744_), .B(new_n31745_), .ZN(new_n31746_));
  OAI21_X1   g28504(.A1(new_n31734_), .A2(new_n31746_), .B(new_n31305_), .ZN(new_n31747_));
  NAND3_X1   g28505(.A1(new_n31742_), .A2(new_n31747_), .A3(pi0572), .ZN(new_n31748_));
  XOR2_X1    g28506(.A1(pi0235), .A2(pi0495), .Z(new_n31749_));
  NOR2_X1    g28507(.A1(new_n31743_), .A2(new_n31749_), .ZN(new_n31750_));
  INV_X1     g28508(.I(new_n31750_), .ZN(new_n31751_));
  AOI21_X1   g28509(.A1(new_n31751_), .A2(new_n31296_), .B(pi0244), .ZN(new_n31752_));
  XNOR2_X1   g28510(.A1(pi0235), .A2(pi0575), .ZN(new_n31753_));
  NAND2_X1   g28511(.A1(new_n31736_), .A2(new_n31753_), .ZN(new_n31754_));
  OAI21_X1   g28512(.A1(new_n31754_), .A2(pi0572), .B(new_n4842_), .ZN(new_n31755_));
  NAND2_X1   g28513(.A1(new_n31755_), .A2(pi0493), .ZN(new_n31756_));
  AOI21_X1   g28514(.A1(new_n31748_), .A2(new_n31752_), .B(new_n31756_), .ZN(new_n31757_));
  OAI21_X1   g28515(.A1(new_n31754_), .A2(new_n31296_), .B(new_n4842_), .ZN(new_n31758_));
  AOI21_X1   g28516(.A1(new_n31750_), .A2(pi0572), .B(new_n31758_), .ZN(new_n31759_));
  AOI21_X1   g28517(.A1(new_n31748_), .A2(new_n31759_), .B(pi0493), .ZN(new_n31760_));
  NOR3_X1    g28518(.A1(new_n31757_), .A2(new_n31760_), .A3(new_n31141_), .ZN(new_n31761_));
  XOR2_X1    g28519(.A1(pi0244), .A2(pi0572), .Z(new_n31762_));
  NOR2_X1    g28520(.A1(new_n31754_), .A2(new_n31762_), .ZN(new_n31763_));
  OAI21_X1   g28521(.A1(new_n31763_), .A2(pi0545), .B(new_n4693_), .ZN(new_n31764_));
  XOR2_X1    g28522(.A1(pi0244), .A2(pi0493), .Z(new_n31765_));
  NOR2_X1    g28523(.A1(new_n31751_), .A2(new_n31765_), .ZN(new_n31766_));
  NAND2_X1   g28524(.A1(new_n31766_), .A2(new_n31141_), .ZN(new_n31767_));
  AOI21_X1   g28525(.A1(new_n31767_), .A2(new_n4693_), .B(new_n31081_), .ZN(new_n31768_));
  OAI21_X1   g28526(.A1(new_n31761_), .A2(new_n31764_), .B(new_n31768_), .ZN(new_n31769_));
  INV_X1     g28527(.I(new_n31766_), .ZN(new_n31770_));
  NOR3_X1    g28528(.A1(new_n31770_), .A2(pi0245), .A3(new_n31141_), .ZN(new_n31771_));
  INV_X1     g28529(.I(new_n31763_), .ZN(new_n31772_));
  OAI21_X1   g28530(.A1(new_n31772_), .A2(new_n31141_), .B(new_n4693_), .ZN(new_n31773_));
  OR3_X2     g28531(.A1(new_n31761_), .A2(new_n31771_), .A3(new_n31773_), .Z(new_n31774_));
  NAND2_X1   g28532(.A1(new_n31774_), .A2(new_n31081_), .ZN(new_n31775_));
  NAND3_X1   g28533(.A1(new_n31775_), .A2(pi0547), .A3(new_n31769_), .ZN(new_n31776_));
  INV_X1     g28534(.I(new_n31776_), .ZN(new_n31777_));
  XOR2_X1    g28535(.A1(pi0245), .A2(pi0545), .Z(new_n31778_));
  NOR2_X1    g28536(.A1(new_n31770_), .A2(new_n31778_), .ZN(new_n31779_));
  INV_X1     g28537(.I(new_n31779_), .ZN(new_n31780_));
  NOR3_X1    g28538(.A1(new_n31780_), .A2(pi0247), .A3(new_n31147_), .ZN(new_n31781_));
  XOR2_X1    g28539(.A1(pi0245), .A2(pi0525), .Z(new_n31782_));
  NOR2_X1    g28540(.A1(new_n31772_), .A2(new_n31782_), .ZN(new_n31783_));
  INV_X1     g28541(.I(new_n31783_), .ZN(new_n31784_));
  NOR2_X1    g28542(.A1(new_n31784_), .A2(new_n31147_), .ZN(new_n31785_));
  NOR4_X1    g28543(.A1(new_n31777_), .A2(pi0247), .A3(new_n31781_), .A4(new_n31785_), .ZN(new_n31786_));
  OAI21_X1   g28544(.A1(new_n31783_), .A2(pi0547), .B(new_n4258_), .ZN(new_n31787_));
  NOR2_X1    g28545(.A1(new_n31777_), .A2(new_n31787_), .ZN(new_n31788_));
  OAI21_X1   g28546(.A1(new_n31780_), .A2(pi0547), .B(new_n4258_), .ZN(new_n31789_));
  NAND2_X1   g28547(.A1(new_n31789_), .A2(pi0527), .ZN(new_n31790_));
  OAI22_X1   g28548(.A1(new_n31786_), .A2(pi0527), .B1(new_n31788_), .B2(new_n31790_), .ZN(new_n31791_));
  AOI21_X1   g28549(.A1(new_n31791_), .A2(pi0238), .B(new_n31093_), .ZN(new_n31792_));
  XOR2_X1    g28550(.A1(pi0247), .A2(pi0547), .Z(new_n31793_));
  NOR2_X1    g28551(.A1(new_n31780_), .A2(new_n31793_), .ZN(new_n31794_));
  XOR2_X1    g28552(.A1(pi0247), .A2(pi0527), .Z(new_n31795_));
  NOR2_X1    g28553(.A1(new_n31784_), .A2(new_n31795_), .ZN(new_n31796_));
  OAI21_X1   g28554(.A1(pi0238), .A2(new_n31796_), .B(new_n31794_), .ZN(new_n31797_));
  INV_X1     g28555(.I(new_n31794_), .ZN(new_n31798_));
  NAND3_X1   g28556(.A1(new_n31798_), .A2(new_n3647_), .A3(new_n31796_), .ZN(new_n31799_));
  NAND4_X1   g28557(.A1(new_n31799_), .A2(pi0491), .A3(new_n31093_), .A4(new_n31797_), .ZN(new_n31800_));
  AOI21_X1   g28558(.A1(new_n31791_), .A2(new_n3647_), .B(pi0529), .ZN(new_n31801_));
  NOR3_X1    g28559(.A1(new_n31784_), .A2(new_n3647_), .A3(new_n31795_), .ZN(new_n31802_));
  NAND3_X1   g28560(.A1(new_n31798_), .A2(pi0238), .A3(new_n31093_), .ZN(new_n31803_));
  OAI21_X1   g28561(.A1(new_n31803_), .A2(new_n31802_), .B(new_n30970_), .ZN(new_n31804_));
  OAI22_X1   g28562(.A1(new_n31792_), .A2(new_n31800_), .B1(new_n31801_), .B2(new_n31804_), .ZN(new_n31805_));
  AOI22_X1   g28563(.A1(new_n31376_), .A2(pi0564), .B1(new_n3828_), .B2(pi0482), .ZN(new_n31806_));
  OAI21_X1   g28564(.A1(new_n3828_), .A2(pi0482), .B(new_n31806_), .ZN(new_n31807_));
  INV_X1     g28565(.I(new_n31807_), .ZN(new_n31808_));
  XOR2_X1    g28566(.A1(pi0241), .A2(pi0562), .Z(new_n31809_));
  NOR2_X1    g28567(.A1(new_n31289_), .A2(pi0234), .ZN(new_n31810_));
  NOR2_X1    g28568(.A1(new_n2440_), .A2(pi0570), .ZN(new_n31811_));
  NOR4_X1    g28569(.A1(new_n31808_), .A2(new_n31809_), .A3(new_n31810_), .A4(new_n31811_), .ZN(new_n31812_));
  NAND2_X1   g28570(.A1(new_n31038_), .A2(new_n31812_), .ZN(new_n31813_));
  NOR2_X1    g28571(.A1(pi0248), .A2(pi0565), .ZN(new_n31814_));
  NOR2_X1    g28572(.A1(new_n31379_), .A2(new_n31201_), .ZN(new_n31815_));
  NOR2_X1    g28573(.A1(new_n31815_), .A2(new_n31814_), .ZN(new_n31816_));
  NOR2_X1    g28574(.A1(new_n31376_), .A2(pi0564), .ZN(new_n31817_));
  NOR4_X1    g28575(.A1(new_n31813_), .A2(new_n31186_), .A3(new_n31816_), .A4(new_n31817_), .ZN(new_n31818_));
  NAND2_X1   g28576(.A1(new_n31186_), .A2(pi0240), .ZN(new_n31819_));
  AOI21_X1   g28577(.A1(new_n31368_), .A2(pi0560), .B(new_n31817_), .ZN(new_n31820_));
  XNOR2_X1   g28578(.A1(pi0248), .A2(pi0565), .ZN(new_n31821_));
  INV_X1     g28579(.I(new_n31821_), .ZN(new_n31822_));
  AOI21_X1   g28580(.A1(new_n31819_), .A2(new_n31820_), .B(new_n31822_), .ZN(new_n31823_));
  NAND3_X1   g28581(.A1(new_n31038_), .A2(new_n31812_), .A3(new_n31823_), .ZN(new_n31824_));
  INV_X1     g28582(.I(new_n31824_), .ZN(new_n31825_));
  MUX2_X1    g28583(.I0(new_n31825_), .I1(new_n31818_), .S(pi0240), .Z(new_n31826_));
  INV_X1     g28584(.I(new_n31826_), .ZN(new_n31827_));
  XNOR2_X1   g28585(.A1(pi0239), .A2(pi0569), .ZN(new_n31828_));
  NOR2_X1    g28586(.A1(new_n31827_), .A2(new_n31828_), .ZN(new_n31829_));
  NOR2_X1    g28587(.A1(new_n31195_), .A2(pi0246), .ZN(new_n31830_));
  NOR2_X1    g28588(.A1(new_n31376_), .A2(pi0563), .ZN(new_n31831_));
  NOR2_X1    g28589(.A1(new_n31379_), .A2(pi0554), .ZN(new_n31832_));
  NOR2_X1    g28590(.A1(new_n31167_), .A2(pi0248), .ZN(new_n31833_));
  NOR4_X1    g28591(.A1(new_n31830_), .A2(new_n31831_), .A3(new_n31832_), .A4(new_n31833_), .ZN(new_n31834_));
  NOR2_X1    g28592(.A1(new_n31164_), .A2(pi0241), .ZN(new_n31835_));
  NOR2_X1    g28593(.A1(new_n31370_), .A2(pi0553), .ZN(new_n31836_));
  NOR2_X1    g28594(.A1(new_n31170_), .A2(pi0249), .ZN(new_n31837_));
  NOR2_X1    g28595(.A1(new_n3828_), .A2(pi0555), .ZN(new_n31838_));
  NOR4_X1    g28596(.A1(new_n31835_), .A2(new_n31836_), .A3(new_n31837_), .A4(new_n31838_), .ZN(new_n31839_));
  NAND2_X1   g28597(.A1(new_n2440_), .A2(pi0485), .ZN(new_n31840_));
  NAND2_X1   g28598(.A1(new_n30953_), .A2(pi0234), .ZN(new_n31841_));
  NAND2_X1   g28599(.A1(new_n31368_), .A2(pi0551), .ZN(new_n31842_));
  NAND2_X1   g28600(.A1(new_n31158_), .A2(pi0240), .ZN(new_n31843_));
  NAND4_X1   g28601(.A1(new_n31840_), .A2(new_n31841_), .A3(new_n31842_), .A4(new_n31843_), .ZN(new_n31844_));
  NOR3_X1    g28602(.A1(new_n31834_), .A2(new_n31839_), .A3(new_n31844_), .ZN(new_n31845_));
  NAND2_X1   g28603(.A1(new_n31016_), .A2(new_n31845_), .ZN(new_n31846_));
  NOR2_X1    g28604(.A1(new_n31846_), .A2(pi0550), .ZN(new_n31847_));
  NOR2_X1    g28605(.A1(new_n31847_), .A2(new_n3409_), .ZN(new_n31848_));
  NOR3_X1    g28606(.A1(new_n31824_), .A2(new_n3409_), .A3(pi0569), .ZN(new_n31849_));
  XNOR2_X1   g28607(.A1(pi0239), .A2(pi0550), .ZN(new_n31850_));
  NOR2_X1    g28608(.A1(new_n31846_), .A2(new_n31850_), .ZN(new_n31851_));
  INV_X1     g28609(.I(new_n31851_), .ZN(new_n31852_));
  NAND2_X1   g28610(.A1(new_n31852_), .A2(pi0569), .ZN(new_n31853_));
  NOR4_X1    g28611(.A1(new_n31853_), .A2(new_n31827_), .A3(new_n31848_), .A4(new_n31849_), .ZN(new_n31854_));
  NAND3_X1   g28612(.A1(new_n31854_), .A2(new_n30964_), .A3(new_n31829_), .ZN(new_n31855_));
  INV_X1     g28613(.I(new_n31829_), .ZN(new_n31856_));
  OAI21_X1   g28614(.A1(new_n31854_), .A2(pi0489), .B(new_n31856_), .ZN(new_n31857_));
  NAND3_X1   g28615(.A1(new_n31851_), .A2(new_n30964_), .A3(pi0556), .ZN(new_n31858_));
  NOR2_X1    g28616(.A1(pi0242), .A2(pi0556), .ZN(new_n31859_));
  NAND4_X1   g28617(.A1(new_n31857_), .A2(new_n31855_), .A3(new_n31858_), .A4(new_n31859_), .ZN(new_n31860_));
  MUX2_X1    g28618(.I0(new_n31854_), .I1(new_n31856_), .S(new_n30964_), .Z(new_n31861_));
  NAND2_X1   g28619(.A1(new_n31859_), .A2(pi0489), .ZN(new_n31862_));
  OAI22_X1   g28620(.A1(new_n31861_), .A2(new_n31173_), .B1(new_n31852_), .B2(new_n31862_), .ZN(new_n31863_));
  AOI21_X1   g28621(.A1(new_n31863_), .A2(new_n31860_), .B(new_n31153_), .ZN(new_n31864_));
  NOR2_X1    g28622(.A1(new_n4929_), .A2(new_n31173_), .ZN(new_n31865_));
  NOR2_X1    g28623(.A1(new_n31865_), .A2(new_n31859_), .ZN(new_n31866_));
  NOR2_X1    g28624(.A1(new_n31856_), .A2(new_n31866_), .ZN(new_n31867_));
  OAI21_X1   g28625(.A1(new_n31867_), .A2(pi0549), .B(new_n3511_), .ZN(new_n31868_));
  XOR2_X1    g28626(.A1(pi0242), .A2(pi0489), .Z(new_n31869_));
  NOR2_X1    g28627(.A1(new_n31852_), .A2(new_n31869_), .ZN(new_n31870_));
  NAND2_X1   g28628(.A1(new_n31870_), .A2(new_n31153_), .ZN(new_n31871_));
  AOI21_X1   g28629(.A1(new_n31871_), .A2(new_n3511_), .B(new_n31099_), .ZN(new_n31872_));
  OAI21_X1   g28630(.A1(new_n31864_), .A2(new_n31868_), .B(new_n31872_), .ZN(new_n31873_));
  NAND2_X1   g28631(.A1(new_n31867_), .A2(pi0549), .ZN(new_n31874_));
  AOI21_X1   g28632(.A1(new_n31870_), .A2(pi0549), .B(pi0235), .ZN(new_n31875_));
  NAND2_X1   g28633(.A1(new_n31874_), .A2(new_n31875_), .ZN(new_n31876_));
  OAI21_X1   g28634(.A1(new_n31864_), .A2(new_n31876_), .B(new_n31099_), .ZN(new_n31877_));
  NAND3_X1   g28635(.A1(new_n31873_), .A2(new_n31877_), .A3(pi0486), .ZN(new_n31878_));
  XNOR2_X1   g28636(.A1(pi0235), .A2(pi0531), .ZN(new_n31879_));
  NAND2_X1   g28637(.A1(new_n31867_), .A2(new_n31879_), .ZN(new_n31880_));
  AOI21_X1   g28638(.A1(new_n31880_), .A2(new_n30956_), .B(pi0244), .ZN(new_n31881_));
  XOR2_X1    g28639(.A1(pi0235), .A2(pi0549), .Z(new_n31882_));
  NOR3_X1    g28640(.A1(new_n31852_), .A2(new_n31869_), .A3(new_n31882_), .ZN(new_n31883_));
  INV_X1     g28641(.I(new_n31883_), .ZN(new_n31884_));
  OAI21_X1   g28642(.A1(new_n31884_), .A2(pi0486), .B(new_n4842_), .ZN(new_n31885_));
  NAND2_X1   g28643(.A1(new_n31885_), .A2(pi0566), .ZN(new_n31886_));
  AOI21_X1   g28644(.A1(new_n31878_), .A2(new_n31881_), .B(new_n31886_), .ZN(new_n31887_));
  NOR2_X1    g28645(.A1(new_n31880_), .A2(new_n30956_), .ZN(new_n31888_));
  OAI21_X1   g28646(.A1(new_n31884_), .A2(new_n30956_), .B(new_n4842_), .ZN(new_n31889_));
  NOR2_X1    g28647(.A1(new_n31888_), .A2(new_n31889_), .ZN(new_n31890_));
  AOI21_X1   g28648(.A1(new_n31878_), .A2(new_n31890_), .B(pi0566), .ZN(new_n31891_));
  NOR3_X1    g28649(.A1(new_n31887_), .A2(new_n31891_), .A3(new_n31284_), .ZN(new_n31892_));
  XOR2_X1    g28650(.A1(pi0244), .A2(pi0486), .Z(new_n31893_));
  NOR2_X1    g28651(.A1(new_n31884_), .A2(new_n31893_), .ZN(new_n31894_));
  OAI21_X1   g28652(.A1(new_n31894_), .A2(pi0568), .B(new_n4693_), .ZN(new_n31895_));
  XOR2_X1    g28653(.A1(pi0244), .A2(pi0566), .Z(new_n31896_));
  NOR2_X1    g28654(.A1(new_n31880_), .A2(new_n31896_), .ZN(new_n31897_));
  NAND2_X1   g28655(.A1(new_n31897_), .A2(new_n31284_), .ZN(new_n31898_));
  AOI21_X1   g28656(.A1(new_n31898_), .A2(new_n4693_), .B(new_n31320_), .ZN(new_n31899_));
  OAI21_X1   g28657(.A1(new_n31892_), .A2(new_n31895_), .B(new_n31899_), .ZN(new_n31900_));
  INV_X1     g28658(.I(new_n31897_), .ZN(new_n31901_));
  NAND2_X1   g28659(.A1(new_n4693_), .A2(pi0568), .ZN(new_n31902_));
  AOI21_X1   g28660(.A1(new_n31894_), .A2(pi0568), .B(pi0245), .ZN(new_n31903_));
  OAI21_X1   g28661(.A1(new_n31901_), .A2(new_n31902_), .B(new_n31903_), .ZN(new_n31904_));
  OAI21_X1   g28662(.A1(new_n31892_), .A2(new_n31904_), .B(new_n31320_), .ZN(new_n31905_));
  NAND3_X1   g28663(.A1(new_n31900_), .A2(new_n31905_), .A3(pi0552), .ZN(new_n31906_));
  XOR2_X1    g28664(.A1(pi0245), .A2(pi0568), .Z(new_n31907_));
  NOR2_X1    g28665(.A1(new_n31901_), .A2(new_n31907_), .ZN(new_n31908_));
  XOR2_X1    g28666(.A1(pi0245), .A2(pi0580), .Z(new_n31909_));
  NOR3_X1    g28667(.A1(new_n31884_), .A2(new_n31893_), .A3(new_n31909_), .ZN(new_n31910_));
  INV_X1     g28668(.I(new_n31910_), .ZN(new_n31911_));
  OAI21_X1   g28669(.A1(new_n31911_), .A2(new_n31161_), .B(new_n4258_), .ZN(new_n31912_));
  AOI21_X1   g28670(.A1(new_n31908_), .A2(pi0552), .B(new_n31912_), .ZN(new_n31913_));
  NAND2_X1   g28671(.A1(new_n31906_), .A2(new_n31913_), .ZN(new_n31914_));
  NAND2_X1   g28672(.A1(new_n31914_), .A2(new_n31102_), .ZN(new_n31915_));
  INV_X1     g28673(.I(new_n31908_), .ZN(new_n31916_));
  AOI21_X1   g28674(.A1(new_n31916_), .A2(new_n31161_), .B(pi0247), .ZN(new_n31917_));
  NAND2_X1   g28675(.A1(new_n31906_), .A2(new_n31917_), .ZN(new_n31918_));
  OAI21_X1   g28676(.A1(new_n31911_), .A2(pi0552), .B(new_n4258_), .ZN(new_n31919_));
  NAND3_X1   g28677(.A1(new_n31918_), .A2(pi0532), .A3(new_n31919_), .ZN(new_n31920_));
  NAND2_X1   g28678(.A1(new_n31920_), .A2(new_n31915_), .ZN(new_n31921_));
  NAND2_X1   g28679(.A1(new_n31921_), .A2(pi0238), .ZN(new_n31922_));
  XOR2_X1    g28680(.A1(pi0247), .A2(pi0532), .Z(new_n31923_));
  NOR2_X1    g28681(.A1(new_n31916_), .A2(new_n31923_), .ZN(new_n31924_));
  XOR2_X1    g28682(.A1(pi0247), .A2(pi0552), .Z(new_n31925_));
  NOR2_X1    g28683(.A1(new_n31911_), .A2(new_n31925_), .ZN(new_n31926_));
  OAI21_X1   g28684(.A1(pi0238), .A2(new_n31926_), .B(new_n31924_), .ZN(new_n31927_));
  INV_X1     g28685(.I(new_n31926_), .ZN(new_n31928_));
  OR3_X2     g28686(.A1(new_n31924_), .A2(pi0238), .A3(new_n31928_), .Z(new_n31929_));
  NAND4_X1   g28687(.A1(new_n31929_), .A2(pi0498), .A3(new_n31311_), .A4(new_n31927_), .ZN(new_n31930_));
  AOI21_X1   g28688(.A1(new_n31922_), .A2(pi0577), .B(new_n31930_), .ZN(new_n31931_));
  NAND2_X1   g28689(.A1(new_n31921_), .A2(new_n3647_), .ZN(new_n31932_));
  NAND3_X1   g28690(.A1(new_n31928_), .A2(pi0238), .A3(new_n31311_), .ZN(new_n31933_));
  OAI21_X1   g28691(.A1(new_n31924_), .A2(new_n31933_), .B(new_n30989_), .ZN(new_n31934_));
  AOI21_X1   g28692(.A1(new_n31932_), .A2(new_n31311_), .B(new_n31934_), .ZN(new_n31935_));
  OAI21_X1   g28693(.A1(new_n31931_), .A2(new_n31935_), .B(new_n24069_), .ZN(new_n31936_));
  NAND2_X1   g28694(.A1(new_n31936_), .A2(new_n24070_), .ZN(new_n31937_));
  AOI21_X1   g28695(.A1(new_n31805_), .A2(pi0233), .B(new_n31937_), .ZN(new_n31938_));
  AOI21_X1   g28696(.A1(new_n31660_), .A2(pi0237), .B(new_n31938_), .ZN(po0750));
  INV_X1     g28697(.I(pi0806), .ZN(new_n31940_));
  NAND3_X1   g28698(.A1(new_n30831_), .A2(new_n31940_), .A3(pi0990), .ZN(new_n31941_));
  INV_X1     g28699(.I(new_n31941_), .ZN(new_n31942_));
  NAND2_X1   g28700(.A1(new_n31940_), .A2(pi0990), .ZN(new_n31943_));
  INV_X1     g28701(.I(new_n31943_), .ZN(new_n31944_));
  NAND3_X1   g28702(.A1(new_n31944_), .A2(new_n2563_), .A3(pi0600), .ZN(new_n31945_));
  NAND2_X1   g28703(.A1(new_n2563_), .A2(pi0594), .ZN(new_n31946_));
  AOI21_X1   g28704(.A1(new_n31945_), .A2(new_n31946_), .B(new_n31942_), .ZN(po0751));
  NAND3_X1   g28705(.A1(new_n30831_), .A2(pi0597), .A3(pi0601), .ZN(new_n31948_));
  NOR3_X1    g28706(.A1(new_n31948_), .A2(new_n30844_), .A3(pi0806), .ZN(new_n31949_));
  XOR2_X1    g28707(.A1(new_n31949_), .A2(new_n30836_), .Z(new_n31950_));
  NOR2_X1    g28708(.A1(new_n31950_), .A2(pi0332), .ZN(po0752));
  INV_X1     g28709(.I(pi0600), .ZN(new_n31952_));
  NAND2_X1   g28710(.A1(pi0595), .A2(pi0597), .ZN(new_n31953_));
  NOR4_X1    g28711(.A1(new_n31943_), .A2(new_n31946_), .A3(new_n31952_), .A4(new_n31953_), .ZN(new_n31954_));
  INV_X1     g28712(.I(pi0596), .ZN(new_n31955_));
  NAND2_X1   g28713(.A1(new_n31954_), .A2(new_n31955_), .ZN(new_n31956_));
  NAND2_X1   g28714(.A1(new_n2563_), .A2(pi0596), .ZN(new_n31957_));
  OAI21_X1   g28715(.A1(new_n31954_), .A2(new_n31957_), .B(new_n31956_), .ZN(po0753));
  XOR2_X1    g28716(.A1(new_n31941_), .A2(pi0597), .Z(new_n31959_));
  NOR2_X1    g28717(.A1(new_n31959_), .A2(pi0332), .ZN(po0754));
  INV_X1     g28718(.I(pi0882), .ZN(new_n31961_));
  NAND2_X1   g28719(.A1(new_n6845_), .A2(new_n31961_), .ZN(new_n31962_));
  NAND2_X1   g28720(.A1(new_n31962_), .A2(new_n5473_), .ZN(new_n31963_));
  NAND2_X1   g28721(.A1(pi0740), .A2(pi0780), .ZN(new_n31964_));
  OAI22_X1   g28722(.A1(new_n31963_), .A2(pi0598), .B1(new_n5427_), .B2(new_n31964_), .ZN(po0755));
  AND4_X2    g28723(.A1(pi0332), .A2(new_n31954_), .A3(pi0596), .A4(pi0599), .Z(po0756));
  NAND2_X1   g28724(.A1(new_n31944_), .A2(new_n31952_), .ZN(new_n31967_));
  NAND2_X1   g28725(.A1(new_n31943_), .A2(pi0600), .ZN(new_n31968_));
  AOI21_X1   g28726(.A1(new_n31967_), .A2(new_n31968_), .B(pi0332), .ZN(po0757));
  NOR2_X1    g28727(.A1(pi0806), .A2(pi0989), .ZN(new_n31970_));
  NOR2_X1    g28728(.A1(new_n31940_), .A2(pi0601), .ZN(new_n31971_));
  NOR3_X1    g28729(.A1(new_n31971_), .A2(pi0332), .A3(new_n31970_), .ZN(po0758));
  NOR3_X1    g28730(.A1(new_n12066_), .A2(new_n11885_), .A3(new_n26307_), .ZN(new_n31973_));
  NOR2_X1    g28731(.A1(new_n12099_), .A2(pi1160), .ZN(new_n31974_));
  OAI21_X1   g28732(.A1(new_n14197_), .A2(new_n31974_), .B(pi0790), .ZN(new_n31975_));
  NAND4_X1   g28733(.A1(new_n31973_), .A2(new_n13637_), .A3(new_n13748_), .A4(new_n31975_), .ZN(new_n31976_));
  OAI22_X1   g28734(.A1(new_n13717_), .A2(new_n31976_), .B1(pi0230), .B2(new_n5394_), .ZN(po0759));
  INV_X1     g28735(.I(pi0966), .ZN(new_n31978_));
  INV_X1     g28736(.I(pi0952), .ZN(new_n31979_));
  INV_X1     g28737(.I(pi1038), .ZN(new_n31980_));
  INV_X1     g28738(.I(pi1060), .ZN(new_n31981_));
  NOR3_X1    g28739(.A1(new_n31980_), .A2(new_n31981_), .A3(pi0980), .ZN(new_n31982_));
  INV_X1     g28740(.I(new_n31982_), .ZN(new_n31983_));
  NOR3_X1    g28741(.A1(new_n31983_), .A2(new_n31979_), .A3(pi1061), .ZN(new_n31984_));
  NOR2_X1    g28742(.A1(new_n13184_), .A2(pi1100), .ZN(new_n31985_));
  AOI21_X1   g28743(.A1(new_n31984_), .A2(new_n31985_), .B(pi0966), .ZN(new_n31986_));
  NAND2_X1   g28744(.A1(new_n31984_), .A2(pi0832), .ZN(new_n31987_));
  NAND2_X1   g28745(.A1(new_n31987_), .A2(new_n5101_), .ZN(new_n31988_));
  NOR2_X1    g28746(.A1(pi0871), .A2(pi0872), .ZN(new_n31989_));
  OAI22_X1   g28747(.A1(new_n31988_), .A2(new_n31986_), .B1(new_n31978_), .B2(new_n31989_), .ZN(po0760));
  INV_X1     g28748(.I(pi0983), .ZN(new_n31991_));
  NOR4_X1    g28749(.A1(new_n15305_), .A2(new_n31991_), .A3(pi0299), .A4(pi0604), .ZN(new_n31992_));
  NOR2_X1    g28750(.A1(new_n12461_), .A2(pi0823), .ZN(new_n31993_));
  MUX2_X1    g28751(.I0(new_n31992_), .I1(pi0779), .S(new_n31993_), .Z(po0761));
  NAND2_X1   g28752(.A1(new_n30844_), .A2(new_n31940_), .ZN(new_n31995_));
  NAND2_X1   g28753(.A1(pi0605), .A2(pi0806), .ZN(new_n31996_));
  AOI21_X1   g28754(.A1(new_n31995_), .A2(new_n31996_), .B(pi0332), .ZN(po0762));
  INV_X1     g28755(.I(pi1104), .ZN(new_n31998_));
  NOR2_X1    g28756(.A1(new_n31987_), .A2(new_n31998_), .ZN(new_n31999_));
  AOI21_X1   g28757(.A1(pi0606), .A2(new_n31987_), .B(new_n31999_), .ZN(new_n32000_));
  NAND2_X1   g28758(.A1(pi0837), .A2(pi0966), .ZN(new_n32001_));
  OAI21_X1   g28759(.A1(new_n32000_), .A2(pi0966), .B(new_n32001_), .ZN(po0763));
  OAI21_X1   g28760(.A1(new_n31987_), .A2(pi1107), .B(new_n31978_), .ZN(new_n32003_));
  AOI21_X1   g28761(.A1(new_n24509_), .A2(new_n31987_), .B(new_n32003_), .ZN(po0764));
  OAI21_X1   g28762(.A1(new_n31987_), .A2(pi1116), .B(new_n31978_), .ZN(new_n32005_));
  AOI21_X1   g28763(.A1(new_n13657_), .A2(new_n31987_), .B(new_n32005_), .ZN(po0765));
  OAI21_X1   g28764(.A1(new_n31987_), .A2(pi1118), .B(new_n31978_), .ZN(new_n32007_));
  AOI21_X1   g28765(.A1(new_n11903_), .A2(new_n31987_), .B(new_n32007_), .ZN(po0766));
  INV_X1     g28766(.I(new_n31987_), .ZN(po0897));
  NOR2_X1    g28767(.A1(po0897), .A2(pi0610), .ZN(new_n32010_));
  OAI21_X1   g28768(.A1(new_n31987_), .A2(pi1113), .B(new_n31978_), .ZN(new_n32011_));
  NOR2_X1    g28769(.A1(new_n32010_), .A2(new_n32011_), .ZN(po0767));
  NOR2_X1    g28770(.A1(po0897), .A2(pi0611), .ZN(new_n32013_));
  OAI21_X1   g28771(.A1(new_n31987_), .A2(pi1114), .B(new_n31978_), .ZN(new_n32014_));
  NOR2_X1    g28772(.A1(new_n32013_), .A2(new_n32014_), .ZN(po0768));
  OAI21_X1   g28773(.A1(new_n31987_), .A2(pi1111), .B(new_n31978_), .ZN(new_n32016_));
  AOI21_X1   g28774(.A1(new_n24919_), .A2(new_n31987_), .B(new_n32016_), .ZN(po0769));
  NOR2_X1    g28775(.A1(po0897), .A2(pi0613), .ZN(new_n32018_));
  OAI21_X1   g28776(.A1(new_n31987_), .A2(pi1115), .B(new_n31978_), .ZN(new_n32019_));
  NOR2_X1    g28777(.A1(new_n32018_), .A2(new_n32019_), .ZN(po0770));
  INV_X1     g28778(.I(pi0871), .ZN(new_n32021_));
  NOR2_X1    g28779(.A1(po0897), .A2(pi0614), .ZN(new_n32022_));
  OAI21_X1   g28780(.A1(new_n31987_), .A2(pi1102), .B(new_n31978_), .ZN(new_n32023_));
  OAI22_X1   g28781(.A1(new_n32022_), .A2(new_n32023_), .B1(new_n32021_), .B2(new_n31978_), .ZN(po0771));
  NAND2_X1   g28782(.A1(new_n31962_), .A2(new_n15305_), .ZN(new_n32025_));
  AND2_X2    g28783(.A1(pi0779), .A2(pi0797), .Z(new_n32026_));
  AOI21_X1   g28784(.A1(new_n5100_), .A2(new_n32026_), .B(pi0615), .ZN(new_n32027_));
  NAND2_X1   g28785(.A1(new_n32025_), .A2(new_n32027_), .ZN(po0772));
  INV_X1     g28786(.I(pi0872), .ZN(new_n32029_));
  NOR2_X1    g28787(.A1(po0897), .A2(pi0616), .ZN(new_n32030_));
  OAI21_X1   g28788(.A1(new_n31987_), .A2(pi1101), .B(new_n31978_), .ZN(new_n32031_));
  OAI22_X1   g28789(.A1(new_n32030_), .A2(new_n32031_), .B1(new_n32029_), .B2(new_n31978_), .ZN(po0773));
  INV_X1     g28790(.I(pi1105), .ZN(new_n32033_));
  NOR2_X1    g28791(.A1(new_n31987_), .A2(new_n32033_), .ZN(new_n32034_));
  AOI21_X1   g28792(.A1(pi0617), .A2(new_n31987_), .B(new_n32034_), .ZN(new_n32035_));
  NAND2_X1   g28793(.A1(pi0850), .A2(pi0966), .ZN(new_n32036_));
  OAI21_X1   g28794(.A1(new_n32035_), .A2(pi0966), .B(new_n32036_), .ZN(po0774));
  OAI21_X1   g28795(.A1(new_n31987_), .A2(pi1117), .B(new_n31978_), .ZN(new_n32038_));
  AOI21_X1   g28796(.A1(new_n11934_), .A2(new_n31987_), .B(new_n32038_), .ZN(po0775));
  OAI21_X1   g28797(.A1(new_n31987_), .A2(pi1122), .B(new_n31978_), .ZN(new_n32040_));
  AOI21_X1   g28798(.A1(new_n11967_), .A2(new_n31987_), .B(new_n32040_), .ZN(po0776));
  NOR2_X1    g28799(.A1(po0897), .A2(pi0620), .ZN(new_n32042_));
  OAI21_X1   g28800(.A1(new_n31987_), .A2(pi1112), .B(new_n31978_), .ZN(new_n32043_));
  NOR2_X1    g28801(.A1(new_n32042_), .A2(new_n32043_), .ZN(po0777));
  OAI21_X1   g28802(.A1(new_n31987_), .A2(pi1108), .B(new_n31978_), .ZN(new_n32045_));
  AOI21_X1   g28803(.A1(new_n11872_), .A2(new_n31987_), .B(new_n32045_), .ZN(po0778));
  OAI21_X1   g28804(.A1(new_n31987_), .A2(pi1109), .B(new_n31978_), .ZN(new_n32047_));
  AOI21_X1   g28805(.A1(new_n24556_), .A2(new_n31987_), .B(new_n32047_), .ZN(po0779));
  OAI21_X1   g28806(.A1(new_n31987_), .A2(pi1106), .B(new_n31978_), .ZN(new_n32049_));
  AOI21_X1   g28807(.A1(new_n24325_), .A2(new_n31987_), .B(new_n32049_), .ZN(po0780));
  NOR4_X1    g28808(.A1(new_n5473_), .A2(new_n31991_), .A3(pi0299), .A4(pi0624), .ZN(new_n32051_));
  NOR2_X1    g28809(.A1(new_n12168_), .A2(pi0831), .ZN(new_n32052_));
  MUX2_X1    g28810(.I0(new_n32051_), .I1(pi0780), .S(new_n32052_), .Z(po0781));
  INV_X1     g28811(.I(pi0953), .ZN(new_n32054_));
  INV_X1     g28812(.I(pi1054), .ZN(new_n32055_));
  NAND3_X1   g28813(.A1(new_n32055_), .A2(pi1066), .A3(pi1088), .ZN(new_n32056_));
  NOR3_X1    g28814(.A1(new_n32056_), .A2(new_n13184_), .A3(pi0973), .ZN(new_n32057_));
  NAND2_X1   g28815(.A1(new_n32057_), .A2(new_n32054_), .ZN(new_n32058_));
  INV_X1     g28816(.I(pi0962), .ZN(new_n32059_));
  OAI21_X1   g28817(.A1(new_n32058_), .A2(pi1116), .B(new_n32059_), .ZN(new_n32060_));
  AOI21_X1   g28818(.A1(new_n12970_), .A2(new_n32058_), .B(new_n32060_), .ZN(po0782));
  OAI21_X1   g28819(.A1(new_n31987_), .A2(pi1121), .B(new_n31978_), .ZN(new_n32062_));
  AOI21_X1   g28820(.A1(new_n11994_), .A2(new_n31987_), .B(new_n32062_), .ZN(po0783));
  OAI21_X1   g28821(.A1(new_n32058_), .A2(pi1117), .B(new_n32059_), .ZN(new_n32064_));
  AOI21_X1   g28822(.A1(new_n11949_), .A2(new_n32058_), .B(new_n32064_), .ZN(po0784));
  OAI21_X1   g28823(.A1(new_n32058_), .A2(pi1119), .B(new_n32059_), .ZN(new_n32066_));
  AOI21_X1   g28824(.A1(new_n12031_), .A2(new_n32058_), .B(new_n32066_), .ZN(po0785));
  OAI21_X1   g28825(.A1(new_n31987_), .A2(pi1119), .B(new_n31978_), .ZN(new_n32068_));
  AOI21_X1   g28826(.A1(new_n12030_), .A2(new_n31987_), .B(new_n32068_), .ZN(po0786));
  OAI21_X1   g28827(.A1(new_n31987_), .A2(pi1120), .B(new_n31978_), .ZN(new_n32070_));
  AOI21_X1   g28828(.A1(new_n12060_), .A2(new_n31987_), .B(new_n32070_), .ZN(po0787));
  NAND3_X1   g28829(.A1(new_n32058_), .A2(pi0631), .A3(pi1113), .ZN(new_n32072_));
  INV_X1     g28830(.I(pi1113), .ZN(new_n32073_));
  INV_X1     g28831(.I(new_n32058_), .ZN(po0954));
  OAI21_X1   g28832(.A1(po0954), .A2(pi0631), .B(new_n32073_), .ZN(new_n32075_));
  NAND3_X1   g28833(.A1(new_n32075_), .A2(new_n32059_), .A3(new_n32072_), .ZN(po0788));
  NAND3_X1   g28834(.A1(new_n32058_), .A2(pi0632), .A3(pi1115), .ZN(new_n32077_));
  INV_X1     g28835(.I(pi1115), .ZN(new_n32078_));
  OAI21_X1   g28836(.A1(po0954), .A2(pi0632), .B(new_n32078_), .ZN(new_n32079_));
  NAND3_X1   g28837(.A1(new_n32079_), .A2(new_n32059_), .A3(new_n32077_), .ZN(po0789));
  OAI21_X1   g28838(.A1(new_n31987_), .A2(pi1110), .B(new_n31978_), .ZN(new_n32081_));
  AOI21_X1   g28839(.A1(new_n23202_), .A2(new_n31987_), .B(new_n32081_), .ZN(po0790));
  OAI21_X1   g28840(.A1(new_n32058_), .A2(pi1110), .B(new_n32059_), .ZN(new_n32083_));
  AOI21_X1   g28841(.A1(new_n23318_), .A2(new_n32058_), .B(new_n32083_), .ZN(po0791));
  NAND3_X1   g28842(.A1(new_n32058_), .A2(pi0635), .A3(pi1112), .ZN(new_n32085_));
  INV_X1     g28843(.I(pi1112), .ZN(new_n32086_));
  OAI21_X1   g28844(.A1(po0954), .A2(pi0635), .B(new_n32086_), .ZN(new_n32087_));
  NAND3_X1   g28845(.A1(new_n32087_), .A2(new_n32059_), .A3(new_n32085_), .ZN(po0792));
  NOR2_X1    g28846(.A1(po0897), .A2(pi0636), .ZN(new_n32089_));
  OAI21_X1   g28847(.A1(new_n31987_), .A2(pi1127), .B(new_n31978_), .ZN(new_n32090_));
  NOR2_X1    g28848(.A1(new_n32089_), .A2(new_n32090_), .ZN(po0793));
  OAI21_X1   g28849(.A1(new_n32058_), .A2(pi1105), .B(new_n32059_), .ZN(new_n32092_));
  AOI21_X1   g28850(.A1(new_n23598_), .A2(new_n32058_), .B(new_n32092_), .ZN(po0794));
  OAI21_X1   g28851(.A1(new_n32058_), .A2(pi1107), .B(new_n32059_), .ZN(new_n32094_));
  AOI21_X1   g28852(.A1(new_n24498_), .A2(new_n32058_), .B(new_n32094_), .ZN(po0795));
  OAI21_X1   g28853(.A1(new_n32058_), .A2(pi1109), .B(new_n32059_), .ZN(new_n32096_));
  AOI21_X1   g28854(.A1(new_n24557_), .A2(new_n32058_), .B(new_n32096_), .ZN(po0796));
  NOR2_X1    g28855(.A1(po0897), .A2(pi0640), .ZN(new_n32098_));
  OAI21_X1   g28856(.A1(new_n31987_), .A2(pi1128), .B(new_n31978_), .ZN(new_n32099_));
  NOR2_X1    g28857(.A1(new_n32098_), .A2(new_n32099_), .ZN(po0797));
  OAI21_X1   g28858(.A1(new_n32058_), .A2(pi1121), .B(new_n32059_), .ZN(new_n32101_));
  AOI21_X1   g28859(.A1(new_n11989_), .A2(new_n32058_), .B(new_n32101_), .ZN(po0798));
  OAI21_X1   g28860(.A1(new_n31987_), .A2(pi1103), .B(new_n31978_), .ZN(new_n32103_));
  AOI21_X1   g28861(.A1(new_n12384_), .A2(new_n31987_), .B(new_n32103_), .ZN(po0799));
  OAI21_X1   g28862(.A1(new_n32058_), .A2(pi1104), .B(new_n32059_), .ZN(new_n32105_));
  AOI21_X1   g28863(.A1(new_n23901_), .A2(new_n32058_), .B(new_n32105_), .ZN(po0800));
  OAI21_X1   g28864(.A1(new_n31987_), .A2(pi1123), .B(new_n31978_), .ZN(new_n32107_));
  AOI21_X1   g28865(.A1(new_n12082_), .A2(new_n31987_), .B(new_n32107_), .ZN(po0801));
  NOR2_X1    g28866(.A1(po0897), .A2(pi0645), .ZN(new_n32109_));
  OAI21_X1   g28867(.A1(new_n31987_), .A2(pi1125), .B(new_n31978_), .ZN(new_n32110_));
  NOR2_X1    g28868(.A1(new_n32109_), .A2(new_n32110_), .ZN(po0802));
  NAND3_X1   g28869(.A1(new_n32058_), .A2(pi0646), .A3(pi1114), .ZN(new_n32112_));
  INV_X1     g28870(.I(pi1114), .ZN(new_n32113_));
  OAI21_X1   g28871(.A1(po0954), .A2(pi0646), .B(new_n32113_), .ZN(new_n32114_));
  NAND3_X1   g28872(.A1(new_n32114_), .A2(new_n32059_), .A3(new_n32112_), .ZN(po0803));
  OAI21_X1   g28873(.A1(new_n32058_), .A2(pi1120), .B(new_n32059_), .ZN(new_n32116_));
  AOI21_X1   g28874(.A1(new_n12061_), .A2(new_n32058_), .B(new_n32116_), .ZN(po0804));
  OAI21_X1   g28875(.A1(new_n32058_), .A2(pi1122), .B(new_n32059_), .ZN(new_n32118_));
  AOI21_X1   g28876(.A1(new_n11966_), .A2(new_n32058_), .B(new_n32118_), .ZN(po0805));
  NAND3_X1   g28877(.A1(new_n32058_), .A2(pi0649), .A3(pi1126), .ZN(new_n32120_));
  INV_X1     g28878(.I(pi1126), .ZN(new_n32121_));
  OAI21_X1   g28879(.A1(po0954), .A2(pi0649), .B(new_n32121_), .ZN(new_n32122_));
  NAND3_X1   g28880(.A1(new_n32122_), .A2(new_n32059_), .A3(new_n32120_), .ZN(po0806));
  NAND3_X1   g28881(.A1(new_n32058_), .A2(pi0650), .A3(pi1127), .ZN(new_n32124_));
  INV_X1     g28882(.I(pi1127), .ZN(new_n32125_));
  OAI21_X1   g28883(.A1(po0954), .A2(pi0650), .B(new_n32125_), .ZN(new_n32126_));
  NAND3_X1   g28884(.A1(new_n32126_), .A2(new_n32059_), .A3(new_n32124_), .ZN(po0807));
  NOR2_X1    g28885(.A1(po0897), .A2(pi0651), .ZN(new_n32128_));
  OAI21_X1   g28886(.A1(new_n31987_), .A2(pi1130), .B(new_n31978_), .ZN(new_n32129_));
  NOR2_X1    g28887(.A1(new_n32128_), .A2(new_n32129_), .ZN(po0808));
  NOR2_X1    g28888(.A1(po0897), .A2(pi0652), .ZN(new_n32131_));
  OAI21_X1   g28889(.A1(new_n31987_), .A2(pi1131), .B(new_n31978_), .ZN(new_n32132_));
  NOR2_X1    g28890(.A1(new_n32131_), .A2(new_n32132_), .ZN(po0809));
  NOR2_X1    g28891(.A1(po0897), .A2(pi0653), .ZN(new_n32134_));
  OAI21_X1   g28892(.A1(new_n31987_), .A2(pi1129), .B(new_n31978_), .ZN(new_n32135_));
  NOR2_X1    g28893(.A1(new_n32134_), .A2(new_n32135_), .ZN(po0810));
  NAND3_X1   g28894(.A1(new_n32058_), .A2(pi0654), .A3(pi1130), .ZN(new_n32137_));
  INV_X1     g28895(.I(pi1130), .ZN(new_n32138_));
  OAI21_X1   g28896(.A1(po0954), .A2(pi0654), .B(new_n32138_), .ZN(new_n32139_));
  NAND3_X1   g28897(.A1(new_n32139_), .A2(new_n32059_), .A3(new_n32137_), .ZN(po0811));
  NAND3_X1   g28898(.A1(new_n32058_), .A2(pi0655), .A3(pi1124), .ZN(new_n32141_));
  INV_X1     g28899(.I(pi1124), .ZN(new_n32142_));
  OAI21_X1   g28900(.A1(po0954), .A2(pi0655), .B(new_n32142_), .ZN(new_n32143_));
  NAND3_X1   g28901(.A1(new_n32143_), .A2(new_n32059_), .A3(new_n32141_), .ZN(po0812));
  NOR2_X1    g28902(.A1(po0897), .A2(pi0656), .ZN(new_n32145_));
  OAI21_X1   g28903(.A1(new_n31987_), .A2(pi1126), .B(new_n31978_), .ZN(new_n32146_));
  NOR2_X1    g28904(.A1(new_n32145_), .A2(new_n32146_), .ZN(po0813));
  NAND3_X1   g28905(.A1(new_n32058_), .A2(pi0657), .A3(pi1131), .ZN(new_n32148_));
  INV_X1     g28906(.I(pi1131), .ZN(new_n32149_));
  OAI21_X1   g28907(.A1(po0954), .A2(pi0657), .B(new_n32149_), .ZN(new_n32150_));
  NAND3_X1   g28908(.A1(new_n32150_), .A2(new_n32059_), .A3(new_n32148_), .ZN(po0814));
  NOR2_X1    g28909(.A1(po0897), .A2(pi0658), .ZN(new_n32152_));
  OAI21_X1   g28910(.A1(new_n31987_), .A2(pi1124), .B(new_n31978_), .ZN(new_n32153_));
  NOR2_X1    g28911(.A1(new_n32152_), .A2(new_n32153_), .ZN(po0815));
  NOR2_X1    g28912(.A1(new_n4559_), .A2(pi0280), .ZN(new_n32155_));
  NAND2_X1   g28913(.A1(new_n32155_), .A2(pi0992), .ZN(new_n32156_));
  NOR3_X1    g28914(.A1(new_n32156_), .A2(pi0269), .A3(pi0281), .ZN(new_n32157_));
  NOR3_X1    g28915(.A1(pi0270), .A2(pi0277), .A3(pi0282), .ZN(new_n32158_));
  NAND2_X1   g28916(.A1(new_n32157_), .A2(new_n32158_), .ZN(new_n32159_));
  NOR3_X1    g28917(.A1(new_n32159_), .A2(pi0264), .A3(pi0265), .ZN(new_n32160_));
  XOR2_X1    g28918(.A1(new_n32160_), .A2(new_n3434_), .Z(po0816));
  OAI21_X1   g28919(.A1(new_n32058_), .A2(pi1118), .B(new_n32059_), .ZN(new_n32162_));
  AOI21_X1   g28920(.A1(new_n11923_), .A2(new_n32058_), .B(new_n32162_), .ZN(po0817));
  OAI21_X1   g28921(.A1(new_n32058_), .A2(pi1101), .B(new_n32059_), .ZN(new_n32164_));
  AOI21_X1   g28922(.A1(new_n24950_), .A2(new_n32058_), .B(new_n32164_), .ZN(po0818));
  OAI21_X1   g28923(.A1(new_n32058_), .A2(pi1102), .B(new_n32059_), .ZN(new_n32166_));
  AOI21_X1   g28924(.A1(new_n24848_), .A2(new_n32058_), .B(new_n32166_), .ZN(po0819));
  NOR2_X1    g28925(.A1(pi1137), .A2(pi1138), .ZN(new_n32168_));
  INV_X1     g28926(.I(new_n32168_), .ZN(new_n32169_));
  NOR2_X1    g28927(.A1(new_n32169_), .A2(pi1134), .ZN(new_n32170_));
  INV_X1     g28928(.I(new_n32170_), .ZN(new_n32171_));
  MUX2_X1    g28929(.I0(pi0784), .I1(pi0634), .S(pi1136), .Z(new_n32172_));
  NAND2_X1   g28930(.A1(new_n32172_), .A2(pi1135), .ZN(new_n32173_));
  AOI21_X1   g28931(.A1(new_n23202_), .A2(pi1136), .B(pi1135), .ZN(new_n32174_));
  OAI21_X1   g28932(.A1(pi0815), .A2(pi1136), .B(new_n32174_), .ZN(new_n32175_));
  AOI21_X1   g28933(.A1(new_n32173_), .A2(new_n32175_), .B(new_n32171_), .ZN(new_n32176_));
  AOI21_X1   g28934(.A1(new_n32168_), .A2(pi1135), .B(new_n4543_), .ZN(new_n32177_));
  INV_X1     g28935(.I(new_n32177_), .ZN(new_n32178_));
  NOR2_X1    g28936(.A1(new_n32178_), .A2(pi0766), .ZN(new_n32179_));
  INV_X1     g28937(.I(pi0855), .ZN(new_n32180_));
  NOR2_X1    g28938(.A1(new_n4696_), .A2(pi1136), .ZN(new_n32181_));
  NOR2_X1    g28939(.A1(new_n32169_), .A2(new_n29634_), .ZN(new_n32182_));
  INV_X1     g28940(.I(new_n32181_), .ZN(new_n32183_));
  NAND2_X1   g28941(.A1(new_n32182_), .A2(new_n32183_), .ZN(new_n32184_));
  INV_X1     g28942(.I(new_n32184_), .ZN(new_n32185_));
  NAND4_X1   g28943(.A1(new_n32185_), .A2(new_n15745_), .A3(new_n32180_), .A4(new_n32181_), .ZN(new_n32186_));
  OAI21_X1   g28944(.A1(new_n32186_), .A2(new_n32179_), .B(new_n10332_), .ZN(new_n32187_));
  NOR2_X1    g28945(.A1(new_n32187_), .A2(new_n32176_), .ZN(new_n32188_));
  XNOR2_X1   g28946(.A1(pi0591), .A2(pi0592), .ZN(new_n32189_));
  INV_X1     g28947(.I(new_n32189_), .ZN(new_n32190_));
  NOR2_X1    g28948(.A1(pi0365), .A2(pi0591), .ZN(new_n32191_));
  AOI21_X1   g28949(.A1(new_n6204_), .A2(pi0591), .B(new_n32191_), .ZN(new_n32192_));
  AOI21_X1   g28950(.A1(new_n32190_), .A2(new_n32192_), .B(pi0590), .ZN(new_n32193_));
  NOR2_X1    g28951(.A1(pi0591), .A2(pi0592), .ZN(new_n32194_));
  NAND2_X1   g28952(.A1(new_n32194_), .A2(pi0590), .ZN(new_n32195_));
  INV_X1     g28953(.I(new_n32195_), .ZN(new_n32196_));
  NAND2_X1   g28954(.A1(new_n32196_), .A2(pi0323), .ZN(new_n32197_));
  INV_X1     g28955(.I(new_n25876_), .ZN(new_n32198_));
  NOR2_X1    g28956(.A1(new_n6798_), .A2(pi0592), .ZN(new_n32199_));
  NAND4_X1   g28957(.A1(new_n32199_), .A2(pi0464), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32200_));
  NAND3_X1   g28958(.A1(new_n32200_), .A2(new_n6711_), .A3(new_n32197_), .ZN(new_n32201_));
  NOR2_X1    g28959(.A1(pi0199), .A2(pi0257), .ZN(new_n32202_));
  OAI21_X1   g28960(.A1(new_n8094_), .A2(pi1065), .B(new_n32198_), .ZN(new_n32203_));
  OAI22_X1   g28961(.A1(new_n32201_), .A2(new_n32193_), .B1(new_n32202_), .B2(new_n32203_), .ZN(new_n32204_));
  NAND2_X1   g28962(.A1(new_n32204_), .A2(new_n6953_), .ZN(new_n32205_));
  XOR2_X1    g28963(.A1(new_n32188_), .A2(new_n32205_), .Z(po0820));
  NOR4_X1    g28964(.A1(new_n32029_), .A2(pi1134), .A3(pi1135), .A4(pi1136), .ZN(new_n32208_));
  OAI21_X1   g28965(.A1(pi0811), .A2(pi1135), .B(pi0785), .ZN(new_n32209_));
  NAND3_X1   g28966(.A1(new_n11870_), .A2(new_n4696_), .A3(pi0811), .ZN(new_n32210_));
  NAND4_X1   g28967(.A1(new_n12443_), .A2(new_n24848_), .A3(new_n4543_), .A4(pi1135), .ZN(new_n32211_));
  NAND4_X1   g28968(.A1(new_n32211_), .A2(new_n4543_), .A3(new_n32210_), .A4(new_n32209_), .ZN(new_n32212_));
  NAND2_X1   g28969(.A1(new_n32212_), .A2(new_n29634_), .ZN(new_n32213_));
  NOR2_X1    g28970(.A1(new_n32169_), .A2(new_n6953_), .ZN(new_n32214_));
  NAND2_X1   g28971(.A1(new_n32213_), .A2(new_n32214_), .ZN(new_n32215_));
  NOR2_X1    g28972(.A1(pi0199), .A2(pi0292), .ZN(new_n32216_));
  NOR2_X1    g28973(.A1(new_n8094_), .A2(pi1084), .ZN(new_n32217_));
  NOR3_X1    g28974(.A1(new_n32217_), .A2(new_n25876_), .A3(new_n32216_), .ZN(new_n32218_));
  NAND2_X1   g28975(.A1(new_n32196_), .A2(pi0355), .ZN(new_n32219_));
  AOI21_X1   g28976(.A1(new_n6203_), .A2(pi0592), .B(pi0588), .ZN(new_n32220_));
  INV_X1     g28977(.I(new_n32220_), .ZN(new_n32221_));
  NOR3_X1    g28978(.A1(new_n9393_), .A2(new_n5940_), .A3(pi0590), .ZN(new_n32222_));
  NOR2_X1    g28979(.A1(new_n30672_), .A2(pi0591), .ZN(new_n32223_));
  AOI22_X1   g28980(.A1(new_n32221_), .A2(new_n32222_), .B1(new_n6084_), .B2(new_n32223_), .ZN(new_n32224_));
  NAND2_X1   g28981(.A1(new_n32224_), .A2(new_n32219_), .ZN(new_n32225_));
  INV_X1     g28982(.I(new_n32199_), .ZN(new_n32226_));
  NOR4_X1    g28983(.A1(new_n32226_), .A2(new_n9301_), .A3(pi0588), .A4(new_n25876_), .ZN(new_n32227_));
  AOI21_X1   g28984(.A1(new_n32225_), .A2(new_n32227_), .B(new_n32218_), .ZN(new_n32228_));
  OAI22_X1   g28985(.A1(new_n32228_), .A2(new_n10332_), .B1(new_n32208_), .B2(new_n32215_), .ZN(po0821));
  OAI21_X1   g28986(.A1(new_n32058_), .A2(pi1108), .B(new_n32059_), .ZN(new_n32230_));
  AOI21_X1   g28987(.A1(new_n11882_), .A2(new_n32058_), .B(new_n32230_), .ZN(po0822));
  NAND3_X1   g28988(.A1(new_n4696_), .A2(pi0790), .A3(pi0799), .ZN(new_n32232_));
  OAI21_X1   g28989(.A1(pi0799), .A2(pi1135), .B(new_n11867_), .ZN(new_n32233_));
  NAND3_X1   g28990(.A1(new_n32233_), .A2(new_n4543_), .A3(new_n32232_), .ZN(new_n32235_));
  NOR2_X1    g28991(.A1(new_n32178_), .A2(pi0764), .ZN(new_n32236_));
  INV_X1     g28992(.I(pi0873), .ZN(new_n32237_));
  NAND4_X1   g28993(.A1(new_n32185_), .A2(new_n16401_), .A3(new_n32237_), .A4(new_n32181_), .ZN(new_n32238_));
  OAI21_X1   g28994(.A1(new_n32238_), .A2(new_n32236_), .B(new_n10332_), .ZN(new_n32239_));
  AOI21_X1   g28995(.A1(new_n32170_), .A2(new_n32235_), .B(new_n32239_), .ZN(new_n32240_));
  NAND4_X1   g28996(.A1(new_n32221_), .A2(pi0456), .A3(new_n6203_), .A4(pi0591), .ZN(new_n32241_));
  NAND3_X1   g28997(.A1(new_n5940_), .A2(new_n6084_), .A3(pi0337), .ZN(new_n32242_));
  NAND2_X1   g28998(.A1(new_n32241_), .A2(new_n32242_), .ZN(new_n32243_));
  AOI21_X1   g28999(.A1(pi0441), .A2(new_n32196_), .B(new_n32243_), .ZN(new_n32244_));
  NAND4_X1   g29000(.A1(new_n32199_), .A2(pi0443), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32245_));
  NOR2_X1    g29001(.A1(pi0199), .A2(pi0297), .ZN(new_n32246_));
  OAI21_X1   g29002(.A1(new_n8094_), .A2(pi1044), .B(new_n32198_), .ZN(new_n32247_));
  OAI22_X1   g29003(.A1(new_n32244_), .A2(new_n32245_), .B1(new_n32246_), .B2(new_n32247_), .ZN(new_n32248_));
  NAND2_X1   g29004(.A1(new_n32248_), .A2(new_n6953_), .ZN(new_n32249_));
  XOR2_X1    g29005(.A1(new_n32249_), .A2(new_n32240_), .Z(po0823));
  NOR4_X1    g29006(.A1(new_n32021_), .A2(pi1134), .A3(pi1135), .A4(pi1136), .ZN(new_n32252_));
  OAI21_X1   g29007(.A1(pi0809), .A2(pi1136), .B(new_n4696_), .ZN(new_n32253_));
  AND3_X2    g29008(.A1(new_n32253_), .A2(pi0642), .A3(pi1136), .Z(new_n32254_));
  OAI21_X1   g29009(.A1(pi0681), .A2(new_n4543_), .B(new_n4696_), .ZN(new_n32255_));
  AOI21_X1   g29010(.A1(new_n11868_), .A2(new_n4543_), .B(new_n32255_), .ZN(new_n32256_));
  OAI21_X1   g29011(.A1(new_n32254_), .A2(new_n32256_), .B(new_n29634_), .ZN(new_n32257_));
  NAND2_X1   g29012(.A1(new_n32257_), .A2(new_n32214_), .ZN(new_n32258_));
  NOR2_X1    g29013(.A1(pi0199), .A2(pi0294), .ZN(new_n32259_));
  NOR2_X1    g29014(.A1(new_n8094_), .A2(pi1072), .ZN(new_n32260_));
  NOR3_X1    g29015(.A1(new_n32260_), .A2(new_n25876_), .A3(new_n32259_), .ZN(new_n32261_));
  NAND2_X1   g29016(.A1(new_n32196_), .A2(pi0458), .ZN(new_n32262_));
  NOR3_X1    g29017(.A1(new_n6212_), .A2(new_n5940_), .A3(pi0590), .ZN(new_n32263_));
  NOR2_X1    g29018(.A1(new_n30571_), .A2(pi0591), .ZN(new_n32264_));
  AOI22_X1   g29019(.A1(new_n32221_), .A2(new_n32263_), .B1(new_n6084_), .B2(new_n32264_), .ZN(new_n32265_));
  NAND2_X1   g29020(.A1(new_n32265_), .A2(new_n32262_), .ZN(new_n32266_));
  NOR4_X1    g29021(.A1(new_n32226_), .A2(new_n6804_), .A3(pi0588), .A4(new_n25876_), .ZN(new_n32267_));
  AOI21_X1   g29022(.A1(new_n32266_), .A2(new_n32267_), .B(new_n32261_), .ZN(new_n32268_));
  OAI22_X1   g29023(.A1(new_n32268_), .A2(new_n10332_), .B1(new_n32258_), .B2(new_n32252_), .ZN(po0824));
  AOI21_X1   g29024(.A1(pi0603), .A2(new_n5095_), .B(new_n4696_), .ZN(new_n32270_));
  NAND2_X1   g29025(.A1(new_n32270_), .A2(pi1136), .ZN(new_n32271_));
  AOI21_X1   g29026(.A1(new_n11891_), .A2(pi1135), .B(pi1136), .ZN(new_n32272_));
  OAI21_X1   g29027(.A1(pi0981), .A2(pi1135), .B(new_n32272_), .ZN(new_n32273_));
  AOI21_X1   g29028(.A1(new_n32273_), .A2(new_n32271_), .B(new_n32171_), .ZN(new_n32274_));
  NOR2_X1    g29029(.A1(new_n32178_), .A2(pi0759), .ZN(new_n32275_));
  INV_X1     g29030(.I(pi0837), .ZN(new_n32276_));
  NAND4_X1   g29031(.A1(new_n32185_), .A2(new_n15674_), .A3(new_n32276_), .A4(new_n32181_), .ZN(new_n32277_));
  OAI21_X1   g29032(.A1(new_n32277_), .A2(new_n32275_), .B(new_n10332_), .ZN(new_n32278_));
  NOR2_X1    g29033(.A1(new_n32278_), .A2(new_n32274_), .ZN(new_n32279_));
  NAND4_X1   g29034(.A1(new_n32221_), .A2(pi0390), .A3(new_n6203_), .A4(pi0591), .ZN(new_n32280_));
  NAND3_X1   g29035(.A1(new_n5940_), .A2(new_n6084_), .A3(pi0363), .ZN(new_n32281_));
  NAND2_X1   g29036(.A1(new_n32280_), .A2(new_n32281_), .ZN(new_n32282_));
  AOI21_X1   g29037(.A1(pi0342), .A2(new_n32196_), .B(new_n32282_), .ZN(new_n32283_));
  NAND4_X1   g29038(.A1(new_n32199_), .A2(pi0414), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32284_));
  NOR2_X1    g29039(.A1(pi0199), .A2(pi0291), .ZN(new_n32285_));
  OAI21_X1   g29040(.A1(new_n8094_), .A2(pi1049), .B(new_n32198_), .ZN(new_n32286_));
  OAI22_X1   g29041(.A1(new_n32283_), .A2(new_n32284_), .B1(new_n32285_), .B2(new_n32286_), .ZN(new_n32287_));
  NAND2_X1   g29042(.A1(new_n32287_), .A2(new_n6953_), .ZN(new_n32288_));
  XOR2_X1    g29043(.A1(new_n32288_), .A2(new_n32279_), .Z(po0825));
  NAND3_X1   g29044(.A1(new_n32058_), .A2(pi0669), .A3(pi1125), .ZN(new_n32290_));
  INV_X1     g29045(.I(pi1125), .ZN(new_n32291_));
  OAI21_X1   g29046(.A1(po0954), .A2(pi0669), .B(new_n32291_), .ZN(new_n32292_));
  NAND3_X1   g29047(.A1(new_n32292_), .A2(new_n32059_), .A3(new_n32290_), .ZN(po0826));
  NAND2_X1   g29048(.A1(new_n32177_), .A2(pi0745), .ZN(new_n32294_));
  NOR4_X1    g29049(.A1(new_n32184_), .A2(new_n15593_), .A3(pi0852), .A4(new_n32183_), .ZN(new_n32295_));
  NOR2_X1    g29050(.A1(new_n32169_), .A2(new_n4543_), .ZN(new_n32296_));
  AOI21_X1   g29051(.A1(new_n24919_), .A2(new_n4696_), .B(pi1134), .ZN(new_n32297_));
  NOR3_X1    g29052(.A1(new_n32297_), .A2(new_n24920_), .A3(new_n4696_), .ZN(new_n32298_));
  AOI22_X1   g29053(.A1(new_n32295_), .A2(new_n32294_), .B1(new_n32296_), .B2(new_n32298_), .ZN(new_n32299_));
  NAND2_X1   g29054(.A1(new_n30637_), .A2(pi0592), .ZN(new_n32300_));
  OAI21_X1   g29055(.A1(pi0391), .A2(pi0592), .B(new_n32300_), .ZN(new_n32301_));
  OAI21_X1   g29056(.A1(new_n32301_), .A2(new_n32189_), .B(new_n6203_), .ZN(new_n32302_));
  NAND4_X1   g29057(.A1(new_n32199_), .A2(pi0415), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32303_));
  NAND2_X1   g29058(.A1(new_n32303_), .A2(new_n6711_), .ZN(new_n32304_));
  AOI21_X1   g29059(.A1(pi0343), .A2(new_n32196_), .B(new_n32304_), .ZN(new_n32305_));
  NOR2_X1    g29060(.A1(pi0199), .A2(pi0258), .ZN(new_n32306_));
  NOR2_X1    g29061(.A1(new_n8094_), .A2(pi1062), .ZN(new_n32307_));
  NOR3_X1    g29062(.A1(new_n32307_), .A2(new_n25876_), .A3(new_n32306_), .ZN(new_n32308_));
  AOI21_X1   g29063(.A1(new_n32305_), .A2(new_n32302_), .B(new_n32308_), .ZN(new_n32309_));
  MUX2_X1    g29064(.I0(new_n32309_), .I1(new_n32299_), .S(new_n10332_), .Z(po0827));
  NAND2_X1   g29065(.A1(new_n32177_), .A2(pi0741), .ZN(new_n32311_));
  NOR4_X1    g29066(.A1(new_n32184_), .A2(new_n15811_), .A3(pi0865), .A4(new_n32183_), .ZN(new_n32312_));
  OAI21_X1   g29067(.A1(pi0611), .A2(pi1135), .B(new_n29634_), .ZN(new_n32313_));
  AND3_X2    g29068(.A1(new_n32296_), .A2(pi0646), .A3(pi1135), .Z(new_n32314_));
  AOI22_X1   g29069(.A1(new_n32312_), .A2(new_n32311_), .B1(new_n32313_), .B2(new_n32314_), .ZN(new_n32315_));
  NAND2_X1   g29070(.A1(new_n6286_), .A2(pi0591), .ZN(new_n32316_));
  OAI21_X1   g29071(.A1(pi0447), .A2(pi0591), .B(new_n32316_), .ZN(new_n32317_));
  OAI21_X1   g29072(.A1(new_n32317_), .A2(new_n32189_), .B(new_n6203_), .ZN(new_n32318_));
  NAND4_X1   g29073(.A1(new_n32199_), .A2(pi0453), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32319_));
  NAND2_X1   g29074(.A1(new_n32319_), .A2(new_n6711_), .ZN(new_n32320_));
  AOI21_X1   g29075(.A1(pi0327), .A2(new_n32196_), .B(new_n32320_), .ZN(new_n32321_));
  NOR2_X1    g29076(.A1(pi0199), .A2(pi0261), .ZN(new_n32322_));
  NOR2_X1    g29077(.A1(new_n8094_), .A2(pi1040), .ZN(new_n32323_));
  NOR3_X1    g29078(.A1(new_n32323_), .A2(new_n25876_), .A3(new_n32322_), .ZN(new_n32324_));
  AOI21_X1   g29079(.A1(new_n32321_), .A2(new_n32318_), .B(new_n32324_), .ZN(new_n32325_));
  MUX2_X1    g29080(.I0(new_n32325_), .I1(new_n32315_), .S(new_n10332_), .Z(po0828));
  AOI21_X1   g29081(.A1(pi0616), .A2(new_n24950_), .B(new_n4696_), .ZN(new_n32327_));
  NAND2_X1   g29082(.A1(new_n32327_), .A2(pi1136), .ZN(new_n32328_));
  AOI21_X1   g29083(.A1(new_n11969_), .A2(pi1135), .B(pi1136), .ZN(new_n32329_));
  OAI21_X1   g29084(.A1(pi0808), .A2(pi1135), .B(new_n32329_), .ZN(new_n32330_));
  AOI21_X1   g29085(.A1(new_n32330_), .A2(new_n32328_), .B(new_n32171_), .ZN(new_n32331_));
  NOR2_X1    g29086(.A1(new_n32178_), .A2(pi0758), .ZN(new_n32332_));
  INV_X1     g29087(.I(pi0850), .ZN(new_n32333_));
  NAND4_X1   g29088(.A1(new_n32185_), .A2(new_n14611_), .A3(new_n32333_), .A4(new_n32181_), .ZN(new_n32334_));
  OAI21_X1   g29089(.A1(new_n32334_), .A2(new_n32332_), .B(new_n10332_), .ZN(new_n32335_));
  NOR2_X1    g29090(.A1(new_n32335_), .A2(new_n32331_), .ZN(new_n32336_));
  NOR2_X1    g29091(.A1(new_n32195_), .A2(new_n6132_), .ZN(new_n32337_));
  NOR4_X1    g29092(.A1(new_n32220_), .A2(new_n6211_), .A3(pi0590), .A4(new_n5940_), .ZN(new_n32338_));
  NOR3_X1    g29093(.A1(new_n6331_), .A2(pi0591), .A3(pi0592), .ZN(new_n32339_));
  NOR3_X1    g29094(.A1(new_n32338_), .A2(new_n32337_), .A3(new_n32339_), .ZN(new_n32340_));
  NAND4_X1   g29095(.A1(new_n32199_), .A2(pi0422), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32341_));
  NOR2_X1    g29096(.A1(pi0199), .A2(pi0290), .ZN(new_n32342_));
  OAI21_X1   g29097(.A1(new_n8094_), .A2(pi1048), .B(new_n32198_), .ZN(new_n32343_));
  OAI22_X1   g29098(.A1(new_n32340_), .A2(new_n32341_), .B1(new_n32342_), .B2(new_n32343_), .ZN(new_n32344_));
  NAND2_X1   g29099(.A1(new_n32344_), .A2(new_n6953_), .ZN(new_n32345_));
  XOR2_X1    g29100(.A1(new_n32336_), .A2(new_n32345_), .Z(po0829));
  NAND3_X1   g29101(.A1(new_n4696_), .A2(pi0788), .A3(pi0814), .ZN(new_n32347_));
  OAI21_X1   g29102(.A1(pi0814), .A2(pi1135), .B(new_n11986_), .ZN(new_n32348_));
  NAND3_X1   g29103(.A1(new_n32348_), .A2(new_n4543_), .A3(new_n32347_), .ZN(new_n32350_));
  NOR2_X1    g29104(.A1(new_n32178_), .A2(pi0749), .ZN(new_n32351_));
  INV_X1     g29105(.I(pi0866), .ZN(new_n32352_));
  NAND4_X1   g29106(.A1(new_n32185_), .A2(new_n13199_), .A3(new_n32352_), .A4(new_n32181_), .ZN(new_n32353_));
  OAI21_X1   g29107(.A1(new_n32353_), .A2(new_n32351_), .B(new_n10332_), .ZN(new_n32354_));
  AOI21_X1   g29108(.A1(new_n32170_), .A2(new_n32350_), .B(new_n32354_), .ZN(new_n32355_));
  NOR2_X1    g29109(.A1(new_n32195_), .A2(new_n6500_), .ZN(new_n32356_));
  NOR4_X1    g29110(.A1(new_n32220_), .A2(new_n6210_), .A3(pi0590), .A4(new_n5940_), .ZN(new_n32357_));
  NOR3_X1    g29111(.A1(new_n6337_), .A2(pi0591), .A3(pi0592), .ZN(new_n32358_));
  NOR3_X1    g29112(.A1(new_n32357_), .A2(new_n32356_), .A3(new_n32358_), .ZN(new_n32359_));
  NAND4_X1   g29113(.A1(new_n32199_), .A2(pi0435), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32360_));
  NOR2_X1    g29114(.A1(pi0199), .A2(pi0295), .ZN(new_n32361_));
  OAI21_X1   g29115(.A1(new_n8094_), .A2(pi1053), .B(new_n32198_), .ZN(new_n32362_));
  OAI22_X1   g29116(.A1(new_n32359_), .A2(new_n32360_), .B1(new_n32361_), .B2(new_n32362_), .ZN(new_n32363_));
  NAND2_X1   g29117(.A1(new_n32363_), .A2(new_n6953_), .ZN(new_n32364_));
  XOR2_X1    g29118(.A1(new_n32355_), .A2(new_n32364_), .Z(po0830));
  INV_X1     g29119(.I(pi0859), .ZN(new_n32366_));
  NOR4_X1    g29120(.A1(new_n32366_), .A2(pi1134), .A3(pi1135), .A4(pi1136), .ZN(new_n32368_));
  OAI21_X1   g29121(.A1(pi0804), .A2(pi1135), .B(pi0783), .ZN(new_n32369_));
  INV_X1     g29122(.I(new_n32369_), .ZN(new_n32370_));
  NOR3_X1    g29123(.A1(new_n30832_), .A2(pi0783), .A3(pi1135), .ZN(new_n32371_));
  NOR4_X1    g29124(.A1(new_n4696_), .A2(pi0622), .A3(pi0639), .A4(pi1136), .ZN(new_n32372_));
  NOR4_X1    g29125(.A1(new_n32370_), .A2(new_n32372_), .A3(new_n32371_), .A4(pi1136), .ZN(new_n32373_));
  OAI21_X1   g29126(.A1(new_n32373_), .A2(pi1134), .B(new_n32214_), .ZN(new_n32374_));
  NOR2_X1    g29127(.A1(pi0199), .A2(pi0256), .ZN(new_n32375_));
  NOR2_X1    g29128(.A1(new_n8094_), .A2(pi1070), .ZN(new_n32376_));
  NOR3_X1    g29129(.A1(new_n32376_), .A2(new_n25876_), .A3(new_n32375_), .ZN(new_n32377_));
  NAND2_X1   g29130(.A1(new_n30565_), .A2(pi0592), .ZN(new_n32378_));
  OAI21_X1   g29131(.A1(pi0463), .A2(pi0592), .B(new_n32378_), .ZN(new_n32379_));
  OAI21_X1   g29132(.A1(new_n32379_), .A2(new_n32189_), .B(new_n6203_), .ZN(new_n32380_));
  NOR2_X1    g29133(.A1(new_n32195_), .A2(new_n6102_), .ZN(new_n32381_));
  NOR4_X1    g29134(.A1(new_n32226_), .A2(new_n6727_), .A3(pi0588), .A4(new_n25876_), .ZN(new_n32382_));
  NOR3_X1    g29135(.A1(new_n32382_), .A2(pi0588), .A3(new_n32381_), .ZN(new_n32383_));
  AOI21_X1   g29136(.A1(new_n32383_), .A2(new_n32380_), .B(new_n32377_), .ZN(new_n32384_));
  OAI22_X1   g29137(.A1(new_n32384_), .A2(new_n10332_), .B1(new_n32368_), .B2(new_n32374_), .ZN(po0831));
  NAND3_X1   g29138(.A1(new_n16315_), .A2(pi0730), .A3(pi1135), .ZN(new_n32386_));
  OAI21_X1   g29139(.A1(new_n4696_), .A2(pi0730), .B(pi0748), .ZN(new_n32387_));
  AOI21_X1   g29140(.A1(new_n32387_), .A2(new_n32386_), .B(new_n4543_), .ZN(new_n32388_));
  NOR2_X1    g29141(.A1(pi1135), .A2(pi1136), .ZN(new_n32389_));
  AND2_X2    g29142(.A1(new_n32389_), .A2(pi0876), .Z(new_n32390_));
  OAI21_X1   g29143(.A1(new_n32388_), .A2(new_n32390_), .B(new_n32182_), .ZN(new_n32391_));
  NOR2_X1    g29144(.A1(pi0803), .A2(pi1135), .ZN(new_n32392_));
  NOR2_X1    g29145(.A1(new_n32392_), .A2(pi1136), .ZN(new_n32393_));
  NAND4_X1   g29146(.A1(new_n4543_), .A2(pi0710), .A3(pi0789), .A4(pi1135), .ZN(new_n32394_));
  OAI21_X1   g29147(.A1(new_n32393_), .A2(new_n32394_), .B(new_n32170_), .ZN(new_n32395_));
  NAND3_X1   g29148(.A1(new_n32395_), .A2(new_n24325_), .A3(new_n32177_), .ZN(new_n32396_));
  NAND3_X1   g29149(.A1(new_n32396_), .A2(new_n10332_), .A3(new_n32391_), .ZN(new_n32397_));
  NOR2_X1    g29150(.A1(new_n32195_), .A2(new_n6503_), .ZN(new_n32398_));
  NOR4_X1    g29151(.A1(new_n32220_), .A2(new_n9405_), .A3(pi0590), .A4(new_n5940_), .ZN(new_n32399_));
  NOR3_X1    g29152(.A1(new_n30689_), .A2(pi0591), .A3(pi0592), .ZN(new_n32400_));
  NOR3_X1    g29153(.A1(new_n32399_), .A2(new_n32398_), .A3(new_n32400_), .ZN(new_n32401_));
  NAND4_X1   g29154(.A1(new_n32199_), .A2(pi0436), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32402_));
  NOR2_X1    g29155(.A1(pi0199), .A2(pi0296), .ZN(new_n32403_));
  OAI21_X1   g29156(.A1(new_n8094_), .A2(pi1037), .B(new_n32198_), .ZN(new_n32404_));
  OAI22_X1   g29157(.A1(new_n32401_), .A2(new_n32402_), .B1(new_n32403_), .B2(new_n32404_), .ZN(new_n32405_));
  NAND2_X1   g29158(.A1(new_n32405_), .A2(new_n6953_), .ZN(new_n32406_));
  XNOR2_X1   g29159(.A1(new_n32406_), .A2(new_n32397_), .ZN(po0832));
  NAND3_X1   g29160(.A1(new_n4696_), .A2(pi0787), .A3(pi0812), .ZN(new_n32408_));
  OAI21_X1   g29161(.A1(pi0812), .A2(pi1135), .B(new_n12048_), .ZN(new_n32409_));
  NAND3_X1   g29162(.A1(new_n32409_), .A2(new_n4543_), .A3(new_n32408_), .ZN(new_n32411_));
  NOR2_X1    g29163(.A1(new_n32178_), .A2(pi0746), .ZN(new_n32412_));
  INV_X1     g29164(.I(pi0881), .ZN(new_n32413_));
  NAND4_X1   g29165(.A1(new_n32185_), .A2(new_n16303_), .A3(new_n32413_), .A4(new_n32181_), .ZN(new_n32414_));
  OAI21_X1   g29166(.A1(new_n32414_), .A2(new_n32412_), .B(new_n10332_), .ZN(new_n32415_));
  AOI21_X1   g29167(.A1(new_n32170_), .A2(new_n32411_), .B(new_n32415_), .ZN(new_n32416_));
  NAND4_X1   g29168(.A1(new_n32221_), .A2(pi0410), .A3(new_n6203_), .A4(pi0591), .ZN(new_n32417_));
  NAND3_X1   g29169(.A1(new_n5940_), .A2(new_n6084_), .A3(pi0386), .ZN(new_n32418_));
  NAND2_X1   g29170(.A1(new_n32417_), .A2(new_n32418_), .ZN(new_n32419_));
  AOI21_X1   g29171(.A1(pi0361), .A2(new_n32196_), .B(new_n32419_), .ZN(new_n32420_));
  NAND4_X1   g29172(.A1(new_n32199_), .A2(pi0434), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32421_));
  NOR2_X1    g29173(.A1(pi0199), .A2(pi0293), .ZN(new_n32422_));
  OAI21_X1   g29174(.A1(new_n8094_), .A2(pi1059), .B(new_n32198_), .ZN(new_n32423_));
  OAI22_X1   g29175(.A1(new_n32420_), .A2(new_n32421_), .B1(new_n32422_), .B2(new_n32423_), .ZN(new_n32424_));
  NAND2_X1   g29176(.A1(new_n32424_), .A2(new_n6953_), .ZN(new_n32425_));
  XOR2_X1    g29177(.A1(new_n32425_), .A2(new_n32416_), .Z(po0833));
  NAND2_X1   g29178(.A1(new_n32177_), .A2(pi0742), .ZN(new_n32427_));
  NOR4_X1    g29179(.A1(new_n32184_), .A2(new_n15756_), .A3(pi0870), .A4(new_n32183_), .ZN(new_n32428_));
  OAI21_X1   g29180(.A1(pi0620), .A2(pi1135), .B(new_n29634_), .ZN(new_n32429_));
  AND3_X2    g29181(.A1(new_n32296_), .A2(pi0635), .A3(pi1135), .Z(new_n32430_));
  AOI22_X1   g29182(.A1(new_n32428_), .A2(new_n32427_), .B1(new_n32429_), .B2(new_n32430_), .ZN(new_n32431_));
  INV_X1     g29183(.I(pi0335), .ZN(new_n32432_));
  NAND2_X1   g29184(.A1(new_n32432_), .A2(pi0591), .ZN(new_n32433_));
  OAI21_X1   g29185(.A1(pi0366), .A2(pi0591), .B(new_n32433_), .ZN(new_n32434_));
  OAI21_X1   g29186(.A1(new_n32434_), .A2(new_n32189_), .B(new_n6203_), .ZN(new_n32435_));
  NAND4_X1   g29187(.A1(new_n32199_), .A2(pi0416), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32436_));
  NAND2_X1   g29188(.A1(new_n32436_), .A2(new_n6711_), .ZN(new_n32437_));
  AOI21_X1   g29189(.A1(pi0344), .A2(new_n32196_), .B(new_n32437_), .ZN(new_n32438_));
  NOR2_X1    g29190(.A1(pi0199), .A2(pi0259), .ZN(new_n32439_));
  NOR2_X1    g29191(.A1(new_n8094_), .A2(pi1069), .ZN(new_n32440_));
  NOR3_X1    g29192(.A1(new_n32440_), .A2(new_n25876_), .A3(new_n32439_), .ZN(new_n32441_));
  AOI21_X1   g29193(.A1(new_n32438_), .A2(new_n32435_), .B(new_n32441_), .ZN(new_n32442_));
  MUX2_X1    g29194(.I0(new_n32431_), .I1(new_n32442_), .S(new_n6953_), .Z(po0834));
  NAND2_X1   g29195(.A1(new_n32177_), .A2(pi0760), .ZN(new_n32444_));
  NOR4_X1    g29196(.A1(new_n32184_), .A2(new_n15830_), .A3(pi0856), .A4(new_n32183_), .ZN(new_n32445_));
  OAI21_X1   g29197(.A1(pi0613), .A2(pi1135), .B(new_n29634_), .ZN(new_n32446_));
  AND3_X2    g29198(.A1(new_n32296_), .A2(pi0632), .A3(pi1135), .Z(new_n32447_));
  AOI22_X1   g29199(.A1(new_n32445_), .A2(new_n32444_), .B1(new_n32446_), .B2(new_n32447_), .ZN(new_n32448_));
  NAND2_X1   g29200(.A1(new_n6321_), .A2(pi0592), .ZN(new_n32449_));
  OAI21_X1   g29201(.A1(pi0393), .A2(pi0592), .B(new_n32449_), .ZN(new_n32450_));
  OAI21_X1   g29202(.A1(new_n32450_), .A2(new_n32189_), .B(new_n6203_), .ZN(new_n32451_));
  NOR2_X1    g29203(.A1(new_n32195_), .A2(new_n6094_), .ZN(new_n32452_));
  NOR4_X1    g29204(.A1(new_n32226_), .A2(new_n6725_), .A3(pi0588), .A4(new_n25876_), .ZN(new_n32453_));
  NOR3_X1    g29205(.A1(new_n32453_), .A2(pi0588), .A3(new_n32452_), .ZN(new_n32454_));
  NOR2_X1    g29206(.A1(pi0199), .A2(pi0260), .ZN(new_n32455_));
  NOR2_X1    g29207(.A1(new_n8094_), .A2(pi1067), .ZN(new_n32456_));
  NOR3_X1    g29208(.A1(new_n32456_), .A2(new_n25876_), .A3(new_n32455_), .ZN(new_n32457_));
  AOI21_X1   g29209(.A1(new_n32454_), .A2(new_n32451_), .B(new_n32457_), .ZN(new_n32458_));
  MUX2_X1    g29210(.I0(new_n32458_), .I1(new_n32448_), .S(new_n10332_), .Z(po0835));
  MUX2_X1    g29211(.I0(pi0791), .I1(pi0665), .S(pi1136), .Z(new_n32460_));
  NAND2_X1   g29212(.A1(new_n32460_), .A2(pi1135), .ZN(new_n32461_));
  AOI21_X1   g29213(.A1(new_n11872_), .A2(pi1136), .B(pi1135), .ZN(new_n32462_));
  OAI21_X1   g29214(.A1(pi0810), .A2(pi1136), .B(new_n32462_), .ZN(new_n32463_));
  AOI21_X1   g29215(.A1(new_n32461_), .A2(new_n32463_), .B(new_n32171_), .ZN(new_n32464_));
  NOR2_X1    g29216(.A1(new_n32178_), .A2(pi0739), .ZN(new_n32465_));
  INV_X1     g29217(.I(pi0874), .ZN(new_n32466_));
  NAND4_X1   g29218(.A1(new_n32185_), .A2(new_n16448_), .A3(new_n32466_), .A4(new_n32181_), .ZN(new_n32467_));
  OAI21_X1   g29219(.A1(new_n32467_), .A2(new_n32465_), .B(new_n10332_), .ZN(new_n32468_));
  NOR2_X1    g29220(.A1(new_n32468_), .A2(new_n32464_), .ZN(new_n32469_));
  NOR2_X1    g29221(.A1(pi0413), .A2(pi0592), .ZN(new_n32470_));
  AOI21_X1   g29222(.A1(new_n6319_), .A2(pi0592), .B(new_n32470_), .ZN(new_n32471_));
  AOI21_X1   g29223(.A1(new_n32190_), .A2(new_n32471_), .B(pi0590), .ZN(new_n32472_));
  NAND2_X1   g29224(.A1(new_n32196_), .A2(pi0450), .ZN(new_n32473_));
  NAND4_X1   g29225(.A1(new_n32199_), .A2(pi0438), .A3(new_n6711_), .A4(new_n32198_), .ZN(new_n32474_));
  NAND3_X1   g29226(.A1(new_n32474_), .A2(new_n6711_), .A3(new_n32473_), .ZN(new_n32475_));
  NOR2_X1    g29227(.A1(pi0199), .A2(pi0255), .ZN(new_n32476_));
  OAI21_X1   g29228(.A1(new_n8094_), .A2(pi1036), .B(new_n32198_), .ZN(new_n32477_));
  OAI22_X1   g29229(.A1(new_n32475_), .A2(new_n32472_), .B1(new_n32476_), .B2(new_n32477_), .ZN(new_n32478_));
  NAND2_X1   g29230(.A1(new_n32478_), .A2(new_n6953_), .ZN(new_n32479_));
  XOR2_X1    g29231(.A1(new_n32469_), .A2(new_n32479_), .Z(po0836));
  OAI21_X1   g29232(.A1(new_n32058_), .A2(pi1100), .B(new_n32059_), .ZN(new_n32481_));
  AOI21_X1   g29233(.A1(new_n5095_), .A2(new_n32058_), .B(new_n32481_), .ZN(po0837));
  OAI21_X1   g29234(.A1(new_n32058_), .A2(pi1103), .B(new_n32059_), .ZN(new_n32483_));
  AOI21_X1   g29235(.A1(new_n12731_), .A2(new_n32058_), .B(new_n32483_), .ZN(po0838));
  NAND2_X1   g29236(.A1(new_n32177_), .A2(pi0757), .ZN(new_n32485_));
  NOR4_X1    g29237(.A1(new_n32184_), .A2(new_n15794_), .A3(pi0848), .A4(new_n32183_), .ZN(new_n32486_));
  OAI21_X1   g29238(.A1(pi0610), .A2(pi1135), .B(new_n29634_), .ZN(new_n32487_));
  AND3_X2    g29239(.A1(new_n32296_), .A2(pi0631), .A3(pi1135), .Z(new_n32488_));
  AOI22_X1   g29240(.A1(new_n32486_), .A2(new_n32485_), .B1(new_n32487_), .B2(new_n32488_), .ZN(new_n32489_));
  NAND2_X1   g29241(.A1(new_n30644_), .A2(pi0592), .ZN(new_n32490_));
  OAI21_X1   g29242(.A1(pi0392), .A2(pi0592), .B(new_n32490_), .ZN(new_n32491_));
  OAI21_X1   g29243(.A1(new_n32491_), .A2(new_n32189_), .B(new_n6203_), .ZN(new_n32492_));
  NOR2_X1    g29244(.A1(new_n32195_), .A2(new_n6093_), .ZN(new_n32493_));
  NOR4_X1    g29245(.A1(new_n32226_), .A2(new_n6724_), .A3(pi0588), .A4(new_n25876_), .ZN(new_n32494_));
  NOR3_X1    g29246(.A1(new_n32494_), .A2(pi0588), .A3(new_n32493_), .ZN(new_n32495_));
  NOR2_X1    g29247(.A1(pi0199), .A2(pi0251), .ZN(new_n32496_));
  NOR2_X1    g29248(.A1(new_n8094_), .A2(pi1039), .ZN(new_n32497_));
  NOR3_X1    g29249(.A1(new_n32497_), .A2(new_n25876_), .A3(new_n32496_), .ZN(new_n32498_));
  AOI21_X1   g29250(.A1(new_n32495_), .A2(new_n32492_), .B(new_n32498_), .ZN(new_n32499_));
  MUX2_X1    g29251(.I0(new_n32499_), .I1(new_n32489_), .S(new_n10332_), .Z(po0839));
  NAND2_X1   g29252(.A1(new_n32057_), .A2(pi0953), .ZN(new_n32501_));
  NAND3_X1   g29253(.A1(new_n32501_), .A2(pi0684), .A3(pi1130), .ZN(new_n32502_));
  INV_X1     g29254(.I(new_n32501_), .ZN(po0980));
  OAI21_X1   g29255(.A1(po0980), .A2(pi0684), .B(new_n32138_), .ZN(new_n32504_));
  NAND3_X1   g29256(.A1(new_n32504_), .A2(new_n32059_), .A3(new_n32502_), .ZN(po0841));
  NAND3_X1   g29257(.A1(new_n32501_), .A2(pi0686), .A3(pi1113), .ZN(new_n32507_));
  OAI21_X1   g29258(.A1(po0980), .A2(pi0686), .B(new_n32073_), .ZN(new_n32508_));
  NAND3_X1   g29259(.A1(new_n32508_), .A2(new_n32059_), .A3(new_n32507_), .ZN(po0843));
  OAI21_X1   g29260(.A1(new_n32501_), .A2(pi1127), .B(new_n32059_), .ZN(new_n32510_));
  AOI21_X1   g29261(.A1(new_n14216_), .A2(new_n32501_), .B(new_n32510_), .ZN(po0844));
  NAND3_X1   g29262(.A1(new_n32501_), .A2(pi0688), .A3(pi1115), .ZN(new_n32512_));
  OAI21_X1   g29263(.A1(po0980), .A2(pi0688), .B(new_n32078_), .ZN(new_n32513_));
  NAND3_X1   g29264(.A1(new_n32513_), .A2(new_n32059_), .A3(new_n32512_), .ZN(po0845));
  OAI21_X1   g29265(.A1(new_n32501_), .A2(pi1108), .B(new_n32059_), .ZN(new_n32516_));
  AOI21_X1   g29266(.A1(new_n16448_), .A2(new_n32501_), .B(new_n32516_), .ZN(po0847));
  OAI21_X1   g29267(.A1(new_n32501_), .A2(pi1107), .B(new_n32059_), .ZN(new_n32518_));
  AOI21_X1   g29268(.A1(new_n16401_), .A2(new_n32501_), .B(new_n32518_), .ZN(po0848));
  NAND4_X1   g29269(.A1(new_n15427_), .A2(new_n4543_), .A3(pi0726), .A4(pi1135), .ZN(new_n32520_));
  NAND4_X1   g29270(.A1(new_n32520_), .A2(pi0844), .A3(new_n29634_), .A4(new_n32389_), .ZN(new_n32521_));
  NAND2_X1   g29271(.A1(new_n32389_), .A2(pi0801), .ZN(new_n32522_));
  NAND4_X1   g29272(.A1(new_n32521_), .A2(new_n10332_), .A3(new_n32170_), .A4(new_n32522_), .ZN(new_n32523_));
  NAND4_X1   g29273(.A1(new_n6203_), .A2(new_n6084_), .A3(pi0402), .A4(pi0591), .ZN(new_n32524_));
  XNOR2_X1   g29274(.A1(pi0590), .A2(pi0592), .ZN(new_n32525_));
  NAND2_X1   g29275(.A1(new_n6356_), .A2(pi0592), .ZN(new_n32526_));
  OAI21_X1   g29276(.A1(pi0352), .A2(pi0592), .B(new_n32526_), .ZN(new_n32527_));
  OAI21_X1   g29277(.A1(new_n32527_), .A2(new_n32525_), .B(new_n5940_), .ZN(new_n32528_));
  NAND3_X1   g29278(.A1(new_n6203_), .A2(new_n5940_), .A3(pi0588), .ZN(new_n32529_));
  NAND2_X1   g29279(.A1(new_n6084_), .A2(pi0427), .ZN(new_n32530_));
  OAI21_X1   g29280(.A1(new_n32529_), .A2(new_n32530_), .B(new_n6711_), .ZN(new_n32531_));
  AOI21_X1   g29281(.A1(new_n32528_), .A2(new_n32524_), .B(new_n32531_), .ZN(new_n32532_));
  NOR3_X1    g29282(.A1(new_n29387_), .A2(pi0199), .A3(new_n30606_), .ZN(new_n32533_));
  AOI21_X1   g29283(.A1(new_n29387_), .A2(new_n8094_), .B(pi1078), .ZN(new_n32534_));
  NOR4_X1    g29284(.A1(new_n32533_), .A2(new_n32534_), .A3(new_n10332_), .A4(new_n25876_), .ZN(new_n32535_));
  OAI21_X1   g29285(.A1(new_n32532_), .A2(new_n32198_), .B(new_n32535_), .ZN(new_n32536_));
  NAND2_X1   g29286(.A1(new_n32536_), .A2(new_n32523_), .ZN(po0849));
  NAND3_X1   g29287(.A1(new_n32058_), .A2(pi0693), .A3(pi1129), .ZN(new_n32538_));
  INV_X1     g29288(.I(pi1129), .ZN(new_n32539_));
  OAI21_X1   g29289(.A1(po0954), .A2(pi0693), .B(new_n32539_), .ZN(new_n32540_));
  NAND3_X1   g29290(.A1(new_n32540_), .A2(new_n32059_), .A3(new_n32538_), .ZN(po0850));
  NAND3_X1   g29291(.A1(new_n32501_), .A2(pi0694), .A3(pi1128), .ZN(new_n32542_));
  INV_X1     g29292(.I(pi1128), .ZN(new_n32543_));
  OAI21_X1   g29293(.A1(po0980), .A2(pi0694), .B(new_n32543_), .ZN(new_n32544_));
  NAND3_X1   g29294(.A1(new_n32544_), .A2(new_n32059_), .A3(new_n32542_), .ZN(po0851));
  NAND3_X1   g29295(.A1(new_n32058_), .A2(pi0695), .A3(pi1111), .ZN(new_n32546_));
  INV_X1     g29296(.I(pi1111), .ZN(new_n32547_));
  OAI21_X1   g29297(.A1(po0954), .A2(pi0695), .B(new_n32547_), .ZN(new_n32548_));
  NAND3_X1   g29298(.A1(new_n32548_), .A2(new_n32059_), .A3(new_n32546_), .ZN(po0852));
  OAI21_X1   g29299(.A1(new_n32501_), .A2(pi1100), .B(new_n32059_), .ZN(new_n32550_));
  AOI21_X1   g29300(.A1(new_n15674_), .A2(new_n32501_), .B(new_n32550_), .ZN(po0853));
  NAND3_X1   g29301(.A1(new_n32501_), .A2(pi0697), .A3(pi1129), .ZN(new_n32552_));
  OAI21_X1   g29302(.A1(po0980), .A2(pi0697), .B(new_n32539_), .ZN(new_n32553_));
  NAND3_X1   g29303(.A1(new_n32553_), .A2(new_n32059_), .A3(new_n32552_), .ZN(po0854));
  NAND3_X1   g29304(.A1(new_n32501_), .A2(pi0698), .A3(pi1116), .ZN(new_n32555_));
  INV_X1     g29305(.I(pi1116), .ZN(new_n32556_));
  OAI21_X1   g29306(.A1(po0980), .A2(pi0698), .B(new_n32556_), .ZN(new_n32557_));
  NAND3_X1   g29307(.A1(new_n32557_), .A2(new_n32059_), .A3(new_n32555_), .ZN(po0855));
  OAI21_X1   g29308(.A1(new_n32501_), .A2(pi1103), .B(new_n32059_), .ZN(new_n32559_));
  AOI21_X1   g29309(.A1(new_n16255_), .A2(new_n32501_), .B(new_n32559_), .ZN(po0856));
  OAI21_X1   g29310(.A1(new_n32501_), .A2(pi1110), .B(new_n32059_), .ZN(new_n32561_));
  AOI21_X1   g29311(.A1(new_n15745_), .A2(new_n32501_), .B(new_n32561_), .ZN(po0857));
  NAND3_X1   g29312(.A1(new_n32501_), .A2(pi0701), .A3(pi1123), .ZN(new_n32563_));
  INV_X1     g29313(.I(pi1123), .ZN(new_n32564_));
  OAI21_X1   g29314(.A1(po0980), .A2(pi0701), .B(new_n32564_), .ZN(new_n32565_));
  NAND3_X1   g29315(.A1(new_n32565_), .A2(new_n32059_), .A3(new_n32563_), .ZN(po0858));
  NAND3_X1   g29316(.A1(new_n32501_), .A2(pi0702), .A3(pi1117), .ZN(new_n32567_));
  INV_X1     g29317(.I(pi1117), .ZN(new_n32568_));
  OAI21_X1   g29318(.A1(po0980), .A2(pi0702), .B(new_n32568_), .ZN(new_n32569_));
  NAND3_X1   g29319(.A1(new_n32569_), .A2(new_n32059_), .A3(new_n32567_), .ZN(po0859));
  OAI21_X1   g29320(.A1(new_n32501_), .A2(pi1124), .B(new_n32059_), .ZN(new_n32571_));
  AOI21_X1   g29321(.A1(new_n16094_), .A2(new_n32501_), .B(new_n32571_), .ZN(po0860));
  NAND3_X1   g29322(.A1(new_n32501_), .A2(pi0704), .A3(pi1112), .ZN(new_n32573_));
  OAI21_X1   g29323(.A1(po0980), .A2(pi0704), .B(new_n32086_), .ZN(new_n32574_));
  NAND3_X1   g29324(.A1(new_n32574_), .A2(new_n32059_), .A3(new_n32573_), .ZN(po0861));
  OAI21_X1   g29325(.A1(new_n32501_), .A2(pi1125), .B(new_n32059_), .ZN(new_n32576_));
  AOI21_X1   g29326(.A1(new_n16198_), .A2(new_n32501_), .B(new_n32576_), .ZN(po0862));
  OAI21_X1   g29327(.A1(new_n32501_), .A2(pi1105), .B(new_n32059_), .ZN(new_n32578_));
  AOI21_X1   g29328(.A1(new_n13199_), .A2(new_n32501_), .B(new_n32578_), .ZN(po0863));
  MUX2_X1    g29329(.I0(new_n11903_), .I1(new_n11923_), .S(pi1135), .Z(new_n32581_));
  NAND2_X1   g29330(.A1(new_n32296_), .A2(new_n29634_), .ZN(new_n32582_));
  OAI21_X1   g29331(.A1(new_n32582_), .A2(new_n32581_), .B(new_n10332_), .ZN(new_n32583_));
  NOR2_X1    g29332(.A1(new_n32169_), .A2(new_n32181_), .ZN(new_n32584_));
  OR2_X2     g29333(.A1(pi0857), .A2(pi1136), .Z(new_n32585_));
  NAND2_X1   g29334(.A1(pi0709), .A2(pi1135), .ZN(new_n32586_));
  NAND4_X1   g29335(.A1(new_n32584_), .A2(pi1134), .A3(new_n32585_), .A4(new_n32586_), .ZN(new_n32587_));
  NAND4_X1   g29336(.A1(new_n32583_), .A2(pi0754), .A3(new_n32177_), .A4(new_n32587_), .ZN(new_n32588_));
  NAND4_X1   g29337(.A1(new_n25876_), .A2(new_n32194_), .A3(pi0588), .A4(new_n6203_), .ZN(new_n32589_));
  NOR3_X1    g29338(.A1(new_n32589_), .A2(new_n6714_), .A3(new_n6953_), .ZN(new_n32590_));
  INV_X1     g29339(.I(pi0305), .ZN(new_n32591_));
  NOR2_X1    g29340(.A1(new_n32591_), .A2(pi0200), .ZN(new_n32592_));
  AOI21_X1   g29341(.A1(pi0200), .A2(pi1084), .B(new_n32592_), .ZN(new_n32593_));
  NAND3_X1   g29342(.A1(new_n32593_), .A2(pi0199), .A3(pi1058), .ZN(new_n32594_));
  INV_X1     g29343(.I(new_n32593_), .ZN(new_n32595_));
  OAI21_X1   g29344(.A1(new_n8094_), .A2(pi1058), .B(new_n32595_), .ZN(new_n32596_));
  AOI21_X1   g29345(.A1(new_n32596_), .A2(new_n32594_), .B(new_n25876_), .ZN(new_n32597_));
  NOR2_X1    g29346(.A1(new_n32195_), .A2(new_n32198_), .ZN(new_n32598_));
  NOR3_X1    g29347(.A1(new_n32198_), .A2(pi0591), .A3(new_n6084_), .ZN(new_n32599_));
  NAND2_X1   g29348(.A1(new_n32599_), .A2(pi0442), .ZN(new_n32600_));
  NOR3_X1    g29349(.A1(new_n32198_), .A2(new_n5940_), .A3(pi0592), .ZN(new_n32601_));
  AOI21_X1   g29350(.A1(new_n32601_), .A2(pi0328), .B(pi0590), .ZN(new_n32602_));
  AOI22_X1   g29351(.A1(new_n32602_), .A2(new_n32600_), .B1(pi0321), .B2(new_n32598_), .ZN(new_n32603_));
  NOR3_X1    g29352(.A1(new_n32597_), .A2(pi0588), .A3(new_n32603_), .ZN(new_n32604_));
  OAI21_X1   g29353(.A1(new_n32604_), .A2(new_n32590_), .B(new_n32588_), .ZN(po0865));
  NAND3_X1   g29354(.A1(new_n32501_), .A2(pi0709), .A3(pi1118), .ZN(new_n32606_));
  INV_X1     g29355(.I(pi1118), .ZN(new_n32607_));
  OAI21_X1   g29356(.A1(po0980), .A2(pi0709), .B(new_n32607_), .ZN(new_n32608_));
  NAND3_X1   g29357(.A1(new_n32608_), .A2(new_n32059_), .A3(new_n32606_), .ZN(po0866));
  OAI21_X1   g29358(.A1(new_n32058_), .A2(pi1106), .B(new_n32059_), .ZN(new_n32610_));
  AOI21_X1   g29359(.A1(new_n24174_), .A2(new_n32058_), .B(new_n32610_), .ZN(po0867));
  INV_X1     g29360(.I(new_n32582_), .ZN(new_n32613_));
  NAND2_X1   g29361(.A1(new_n32177_), .A2(pi0751), .ZN(new_n32614_));
  INV_X1     g29362(.I(new_n32584_), .ZN(new_n32615_));
  NOR2_X1    g29363(.A1(pi0842), .A2(pi1136), .ZN(new_n32616_));
  NOR2_X1    g29364(.A1(new_n15564_), .A2(new_n4696_), .ZN(new_n32617_));
  NOR4_X1    g29365(.A1(new_n32615_), .A2(new_n29634_), .A3(new_n32616_), .A4(new_n32617_), .ZN(new_n32618_));
  MUX2_X1    g29366(.I0(pi0644), .I1(pi0715), .S(pi1135), .Z(new_n32619_));
  AOI22_X1   g29367(.A1(new_n32618_), .A2(new_n32614_), .B1(new_n32613_), .B2(new_n32619_), .ZN(new_n32620_));
  NOR2_X1    g29368(.A1(pi0400), .A2(pi0592), .ZN(new_n32621_));
  AOI21_X1   g29369(.A1(new_n6689_), .A2(pi0592), .B(new_n32621_), .ZN(new_n32622_));
  NAND2_X1   g29370(.A1(new_n32190_), .A2(new_n32622_), .ZN(new_n32623_));
  NOR3_X1    g29371(.A1(new_n32195_), .A2(new_n6108_), .A3(pi0590), .ZN(new_n32624_));
  AOI21_X1   g29372(.A1(new_n32623_), .A2(new_n32624_), .B(pi0588), .ZN(new_n32625_));
  NAND2_X1   g29373(.A1(new_n6084_), .A2(pi0425), .ZN(new_n32626_));
  OAI21_X1   g29374(.A1(new_n32529_), .A2(new_n32626_), .B(new_n25876_), .ZN(new_n32627_));
  INV_X1     g29375(.I(pi0298), .ZN(new_n32628_));
  NOR2_X1    g29376(.A1(new_n26635_), .A2(new_n30408_), .ZN(new_n32629_));
  OAI21_X1   g29377(.A1(new_n8094_), .A2(new_n30600_), .B(new_n32198_), .ZN(new_n32630_));
  OAI22_X1   g29378(.A1(new_n32629_), .A2(new_n32630_), .B1(new_n32628_), .B2(new_n8161_), .ZN(new_n32631_));
  OAI21_X1   g29379(.A1(new_n32625_), .A2(new_n32627_), .B(new_n32631_), .ZN(new_n32632_));
  MUX2_X1    g29380(.I0(new_n32620_), .I1(new_n32632_), .S(new_n6953_), .Z(po0869));
  OAI21_X1   g29381(.A1(new_n32058_), .A2(pi1123), .B(new_n32059_), .ZN(new_n32636_));
  AOI21_X1   g29382(.A1(new_n12099_), .A2(new_n32058_), .B(new_n32636_), .ZN(po0872));
  MUX2_X1    g29383(.I0(new_n11994_), .I1(new_n11989_), .S(pi1135), .Z(new_n32638_));
  OAI21_X1   g29384(.A1(new_n32582_), .A2(new_n32638_), .B(new_n10332_), .ZN(new_n32639_));
  OR2_X2     g29385(.A1(pi0845), .A2(pi1136), .Z(new_n32640_));
  NAND2_X1   g29386(.A1(pi0738), .A2(pi1135), .ZN(new_n32641_));
  NAND4_X1   g29387(.A1(new_n32584_), .A2(pi1134), .A3(new_n32640_), .A4(new_n32641_), .ZN(new_n32642_));
  NAND4_X1   g29388(.A1(new_n32639_), .A2(pi0761), .A3(new_n32177_), .A4(new_n32642_), .ZN(new_n32643_));
  NOR3_X1    g29389(.A1(new_n32589_), .A2(new_n6713_), .A3(new_n6953_), .ZN(new_n32644_));
  INV_X1     g29390(.I(pi0307), .ZN(new_n32645_));
  NOR2_X1    g29391(.A1(new_n32645_), .A2(pi0200), .ZN(new_n32646_));
  AOI21_X1   g29392(.A1(pi0200), .A2(pi1053), .B(new_n32646_), .ZN(new_n32647_));
  NAND3_X1   g29393(.A1(new_n32647_), .A2(pi0199), .A3(pi1043), .ZN(new_n32648_));
  INV_X1     g29394(.I(new_n32647_), .ZN(new_n32649_));
  OAI21_X1   g29395(.A1(new_n8094_), .A2(pi1043), .B(new_n32649_), .ZN(new_n32650_));
  AOI21_X1   g29396(.A1(new_n32650_), .A2(new_n32648_), .B(new_n25876_), .ZN(new_n32651_));
  NAND2_X1   g29397(.A1(new_n32599_), .A2(pi0440), .ZN(new_n32652_));
  AOI21_X1   g29398(.A1(new_n32601_), .A2(pi0329), .B(pi0590), .ZN(new_n32653_));
  AOI22_X1   g29399(.A1(new_n32653_), .A2(new_n32652_), .B1(pi0349), .B2(new_n32598_), .ZN(new_n32654_));
  NOR3_X1    g29400(.A1(new_n32651_), .A2(pi0588), .A3(new_n32654_), .ZN(new_n32655_));
  OAI21_X1   g29401(.A1(new_n32655_), .A2(new_n32644_), .B(new_n32643_), .ZN(po0873));
  NOR2_X1    g29402(.A1(new_n5940_), .A2(pi0318), .ZN(new_n32657_));
  AOI21_X1   g29403(.A1(new_n6354_), .A2(new_n5940_), .B(new_n32657_), .ZN(new_n32658_));
  NAND2_X1   g29404(.A1(new_n32190_), .A2(new_n32658_), .ZN(new_n32659_));
  NOR3_X1    g29405(.A1(new_n32195_), .A2(new_n6193_), .A3(pi0590), .ZN(new_n32660_));
  NAND2_X1   g29406(.A1(new_n25876_), .A2(new_n6711_), .ZN(new_n32661_));
  AOI21_X1   g29407(.A1(new_n32659_), .A2(new_n32660_), .B(new_n32661_), .ZN(new_n32662_));
  NOR3_X1    g29408(.A1(new_n29381_), .A2(pi0199), .A3(new_n30509_), .ZN(new_n32663_));
  AOI21_X1   g29409(.A1(new_n29381_), .A2(new_n8094_), .B(pi1074), .ZN(new_n32664_));
  NOR2_X1    g29410(.A1(pi0223), .A2(pi0224), .ZN(new_n32665_));
  NOR3_X1    g29411(.A1(new_n32663_), .A2(new_n32664_), .A3(new_n32665_), .ZN(new_n32666_));
  NOR2_X1    g29412(.A1(new_n32662_), .A2(new_n32666_), .ZN(new_n32667_));
  INV_X1     g29413(.I(pi0669), .ZN(new_n32668_));
  MUX2_X1    g29414(.I0(pi0645), .I1(new_n32668_), .S(pi1135), .Z(new_n32669_));
  AOI22_X1   g29415(.A1(new_n32669_), .A2(pi1136), .B1(pi0800), .B2(new_n32389_), .ZN(new_n32670_));
  NOR2_X1    g29416(.A1(pi0839), .A2(pi1136), .ZN(new_n32671_));
  NOR2_X1    g29417(.A1(new_n16198_), .A2(pi1135), .ZN(new_n32672_));
  NOR4_X1    g29418(.A1(new_n32615_), .A2(new_n29634_), .A3(new_n32671_), .A4(new_n32672_), .ZN(new_n32673_));
  NAND2_X1   g29419(.A1(new_n32177_), .A2(pi0768), .ZN(new_n32674_));
  OAI22_X1   g29420(.A1(new_n32673_), .A2(new_n32674_), .B1(new_n32171_), .B2(new_n32670_), .ZN(new_n32675_));
  MUX2_X1    g29421(.I0(new_n32675_), .I1(new_n32667_), .S(new_n6953_), .Z(po0874));
  MUX2_X1    g29422(.I0(new_n13657_), .I1(new_n12970_), .S(pi1135), .Z(new_n32677_));
  OAI21_X1   g29423(.A1(new_n32582_), .A2(new_n32677_), .B(new_n10332_), .ZN(new_n32678_));
  OR2_X2     g29424(.A1(pi0853), .A2(pi1136), .Z(new_n32679_));
  NAND2_X1   g29425(.A1(pi0698), .A2(pi1135), .ZN(new_n32680_));
  NAND4_X1   g29426(.A1(new_n32584_), .A2(pi1134), .A3(new_n32679_), .A4(new_n32680_), .ZN(new_n32681_));
  NAND4_X1   g29427(.A1(new_n32678_), .A2(pi0767), .A3(new_n32177_), .A4(new_n32681_), .ZN(new_n32682_));
  NAND2_X1   g29428(.A1(new_n10332_), .A2(pi0419), .ZN(new_n32683_));
  NOR2_X1    g29429(.A1(new_n32683_), .A2(new_n32589_), .ZN(new_n32684_));
  INV_X1     g29430(.I(pi0303), .ZN(new_n32685_));
  NOR2_X1    g29431(.A1(new_n32685_), .A2(pi0200), .ZN(new_n32686_));
  AOI21_X1   g29432(.A1(pi0200), .A2(pi1049), .B(new_n32686_), .ZN(new_n32687_));
  NAND3_X1   g29433(.A1(new_n32687_), .A2(pi0199), .A3(pi1080), .ZN(new_n32688_));
  INV_X1     g29434(.I(new_n32687_), .ZN(new_n32689_));
  OAI21_X1   g29435(.A1(new_n8094_), .A2(pi1080), .B(new_n32689_), .ZN(new_n32690_));
  AOI21_X1   g29436(.A1(new_n32690_), .A2(new_n32688_), .B(new_n25876_), .ZN(new_n32691_));
  NAND2_X1   g29437(.A1(new_n32599_), .A2(pi0369), .ZN(new_n32692_));
  AOI21_X1   g29438(.A1(new_n32601_), .A2(pi0394), .B(pi0590), .ZN(new_n32693_));
  AOI22_X1   g29439(.A1(new_n32693_), .A2(new_n32692_), .B1(pi0315), .B2(new_n32598_), .ZN(new_n32694_));
  NOR3_X1    g29440(.A1(new_n32691_), .A2(pi0588), .A3(new_n32694_), .ZN(new_n32695_));
  OAI21_X1   g29441(.A1(new_n32695_), .A2(new_n32684_), .B(new_n32682_), .ZN(po0875));
  NOR2_X1    g29442(.A1(new_n5940_), .A2(pi0325), .ZN(new_n32697_));
  AOI21_X1   g29443(.A1(new_n6358_), .A2(new_n5940_), .B(new_n32697_), .ZN(new_n32698_));
  NAND2_X1   g29444(.A1(new_n32190_), .A2(new_n32698_), .ZN(new_n32699_));
  AND3_X2    g29445(.A1(new_n32196_), .A2(pi0353), .A3(new_n6203_), .Z(new_n32700_));
  AOI21_X1   g29446(.A1(new_n32700_), .A2(new_n32699_), .B(new_n32661_), .ZN(new_n32701_));
  NOR3_X1    g29447(.A1(new_n29393_), .A2(pi0199), .A3(new_n30529_), .ZN(new_n32702_));
  AOI21_X1   g29448(.A1(new_n29393_), .A2(new_n8094_), .B(pi1063), .ZN(new_n32703_));
  NOR2_X1    g29449(.A1(pi0223), .A2(pi0224), .ZN(new_n32704_));
  NOR3_X1    g29450(.A1(new_n32702_), .A2(new_n32703_), .A3(new_n32704_), .ZN(new_n32705_));
  NOR2_X1    g29451(.A1(new_n32701_), .A2(new_n32705_), .ZN(new_n32706_));
  INV_X1     g29452(.I(pi0650), .ZN(new_n32707_));
  MUX2_X1    g29453(.I0(pi0636), .I1(new_n32707_), .S(pi1135), .Z(new_n32708_));
  AOI22_X1   g29454(.A1(new_n32708_), .A2(pi1136), .B1(pi0807), .B2(new_n32389_), .ZN(new_n32709_));
  NOR2_X1    g29455(.A1(pi0868), .A2(pi1136), .ZN(new_n32710_));
  NOR2_X1    g29456(.A1(new_n14216_), .A2(pi1135), .ZN(new_n32711_));
  NOR4_X1    g29457(.A1(new_n32615_), .A2(new_n29634_), .A3(new_n32710_), .A4(new_n32711_), .ZN(new_n32712_));
  NAND2_X1   g29458(.A1(new_n32177_), .A2(pi0774), .ZN(new_n32713_));
  OAI22_X1   g29459(.A1(new_n32712_), .A2(new_n32713_), .B1(new_n32171_), .B2(new_n32709_), .ZN(new_n32714_));
  MUX2_X1    g29460(.I0(new_n32714_), .I1(new_n32706_), .S(new_n6953_), .Z(po0876));
  INV_X1     g29461(.I(pi0816), .ZN(new_n32717_));
  INV_X1     g29462(.I(pi0721), .ZN(new_n32718_));
  INV_X1     g29463(.I(pi0813), .ZN(new_n32719_));
  XNOR2_X1   g29464(.A1(pi0771), .A2(pi0800), .ZN(new_n32720_));
  INV_X1     g29465(.I(pi0747), .ZN(new_n32721_));
  INV_X1     g29466(.I(pi0807), .ZN(new_n32722_));
  XOR2_X1    g29467(.A1(pi0765), .A2(pi0798), .Z(new_n32723_));
  NOR2_X1    g29468(.A1(new_n32723_), .A2(new_n32722_), .ZN(new_n32724_));
  INV_X1     g29469(.I(new_n32724_), .ZN(new_n32725_));
  INV_X1     g29470(.I(pi0798), .ZN(new_n32726_));
  NOR2_X1    g29471(.A1(new_n32726_), .A2(pi0765), .ZN(new_n32727_));
  INV_X1     g29472(.I(pi0765), .ZN(new_n32728_));
  NOR2_X1    g29473(.A1(new_n32728_), .A2(pi0798), .ZN(new_n32729_));
  NOR4_X1    g29474(.A1(new_n32727_), .A2(new_n32729_), .A3(pi0747), .A4(pi0807), .ZN(new_n32730_));
  OAI21_X1   g29475(.A1(new_n32725_), .A2(new_n32721_), .B(new_n32730_), .ZN(new_n32731_));
  INV_X1     g29476(.I(new_n32731_), .ZN(new_n32732_));
  XOR2_X1    g29477(.A1(pi0769), .A2(pi0794), .Z(new_n32733_));
  NOR2_X1    g29478(.A1(new_n32732_), .A2(new_n32733_), .ZN(new_n32734_));
  NAND2_X1   g29479(.A1(new_n32734_), .A2(new_n32720_), .ZN(new_n32735_));
  XOR2_X1    g29480(.A1(pi0773), .A2(pi0801), .Z(new_n32736_));
  NOR2_X1    g29481(.A1(new_n32735_), .A2(new_n32736_), .ZN(new_n32737_));
  INV_X1     g29482(.I(new_n32737_), .ZN(new_n32738_));
  NOR3_X1    g29483(.A1(new_n32738_), .A2(new_n32718_), .A3(new_n32719_), .ZN(new_n32739_));
  INV_X1     g29484(.I(new_n32720_), .ZN(new_n32740_));
  NOR2_X1    g29485(.A1(new_n32725_), .A2(new_n32740_), .ZN(new_n32741_));
  INV_X1     g29486(.I(pi0794), .ZN(new_n32742_));
  INV_X1     g29487(.I(pi0801), .ZN(new_n32743_));
  NOR4_X1    g29488(.A1(new_n32742_), .A2(new_n32743_), .A3(pi0721), .A4(pi0813), .ZN(new_n32744_));
  AOI21_X1   g29489(.A1(new_n32741_), .A2(new_n32744_), .B(new_n32739_), .ZN(new_n32745_));
  INV_X1     g29490(.I(pi0775), .ZN(new_n32746_));
  INV_X1     g29491(.I(pi0731), .ZN(new_n32747_));
  INV_X1     g29492(.I(pi0945), .ZN(new_n32748_));
  NAND2_X1   g29493(.A1(new_n32748_), .A2(pi0988), .ZN(new_n32749_));
  NOR2_X1    g29494(.A1(new_n32749_), .A2(new_n32747_), .ZN(new_n32750_));
  AND2_X2    g29495(.A1(pi0747), .A2(pi0773), .Z(new_n32751_));
  NAND2_X1   g29496(.A1(new_n32751_), .A2(pi0769), .ZN(new_n32752_));
  XOR2_X1    g29497(.A1(new_n32752_), .A2(pi0721), .Z(new_n32753_));
  NOR2_X1    g29498(.A1(new_n32718_), .A2(pi0775), .ZN(new_n32754_));
  NOR4_X1    g29499(.A1(new_n32753_), .A2(new_n32746_), .A3(pi0795), .A4(new_n32750_), .ZN(new_n32755_));
  OAI21_X1   g29500(.A1(new_n32745_), .A2(new_n32717_), .B(new_n32755_), .ZN(new_n32756_));
  INV_X1     g29501(.I(new_n32750_), .ZN(new_n32757_));
  NOR2_X1    g29502(.A1(pi0775), .A2(pi0816), .ZN(new_n32758_));
  NOR2_X1    g29503(.A1(new_n32746_), .A2(new_n32717_), .ZN(new_n32759_));
  OAI21_X1   g29504(.A1(new_n32758_), .A2(new_n32759_), .B(new_n32739_), .ZN(new_n32760_));
  INV_X1     g29505(.I(new_n32760_), .ZN(new_n32761_));
  XNOR2_X1   g29506(.A1(pi0731), .A2(pi0795), .ZN(new_n32762_));
  NAND4_X1   g29507(.A1(new_n32761_), .A2(new_n32718_), .A3(new_n32757_), .A4(new_n32762_), .ZN(new_n32763_));
  NAND2_X1   g29508(.A1(new_n32760_), .A2(new_n32754_), .ZN(new_n32764_));
  NAND3_X1   g29509(.A1(new_n32763_), .A2(new_n32764_), .A3(new_n32756_), .ZN(po0878));
  INV_X1     g29510(.I(pi0795), .ZN(new_n32766_));
  NAND3_X1   g29511(.A1(new_n32766_), .A2(pi0851), .A3(pi1134), .ZN(new_n32767_));
  OAI21_X1   g29512(.A1(new_n29634_), .A2(pi0851), .B(pi0795), .ZN(new_n32768_));
  AOI21_X1   g29513(.A1(new_n32768_), .A2(new_n32767_), .B(pi1136), .ZN(new_n32769_));
  INV_X1     g29514(.I(pi0776), .ZN(new_n32770_));
  OAI21_X1   g29515(.A1(pi0640), .A2(pi1134), .B(new_n32770_), .ZN(new_n32771_));
  NAND3_X1   g29516(.A1(new_n29634_), .A2(pi0640), .A3(pi0776), .ZN(new_n32772_));
  AOI21_X1   g29517(.A1(new_n32771_), .A2(new_n32772_), .B(new_n4543_), .ZN(new_n32773_));
  OAI21_X1   g29518(.A1(new_n32773_), .A2(new_n32769_), .B(new_n4696_), .ZN(new_n32774_));
  INV_X1     g29519(.I(pi0694), .ZN(new_n32775_));
  AOI22_X1   g29520(.A1(new_n32775_), .A2(pi1134), .B1(pi1135), .B2(pi1136), .ZN(new_n32776_));
  OAI21_X1   g29521(.A1(pi0732), .A2(pi1134), .B(new_n32776_), .ZN(new_n32777_));
  NAND3_X1   g29522(.A1(new_n32774_), .A2(new_n32214_), .A3(new_n32777_), .ZN(new_n32778_));
  NOR3_X1    g29523(.A1(new_n29399_), .A2(pi0199), .A3(new_n30611_), .ZN(new_n32779_));
  AOI21_X1   g29524(.A1(new_n29399_), .A2(new_n8094_), .B(pi1045), .ZN(new_n32780_));
  NOR2_X1    g29525(.A1(pi0403), .A2(pi0592), .ZN(new_n32781_));
  AOI21_X1   g29526(.A1(new_n30669_), .A2(pi0592), .B(new_n32781_), .ZN(new_n32782_));
  NAND2_X1   g29527(.A1(new_n32190_), .A2(new_n32782_), .ZN(new_n32783_));
  NOR3_X1    g29528(.A1(new_n32195_), .A2(new_n6192_), .A3(pi0590), .ZN(new_n32784_));
  AOI21_X1   g29529(.A1(new_n32783_), .A2(new_n32784_), .B(pi0588), .ZN(new_n32785_));
  NOR2_X1    g29530(.A1(pi0223), .A2(pi0224), .ZN(new_n32786_));
  NOR4_X1    g29531(.A1(new_n32785_), .A2(new_n32779_), .A3(new_n32780_), .A4(new_n32786_), .ZN(new_n32787_));
  NOR2_X1    g29532(.A1(new_n32787_), .A2(new_n10332_), .ZN(new_n32788_));
  XNOR2_X1   g29533(.A1(new_n32788_), .A2(new_n32778_), .ZN(po0879));
  NAND3_X1   g29534(.A1(new_n32501_), .A2(pi0723), .A3(pi1111), .ZN(new_n32790_));
  OAI21_X1   g29535(.A1(po0980), .A2(pi0723), .B(new_n32547_), .ZN(new_n32791_));
  NAND3_X1   g29536(.A1(new_n32791_), .A2(new_n32059_), .A3(new_n32790_), .ZN(po0880));
  NAND3_X1   g29537(.A1(new_n32501_), .A2(pi0724), .A3(pi1114), .ZN(new_n32793_));
  OAI21_X1   g29538(.A1(po0980), .A2(pi0724), .B(new_n32113_), .ZN(new_n32794_));
  NAND3_X1   g29539(.A1(new_n32794_), .A2(new_n32059_), .A3(new_n32793_), .ZN(po0881));
  NAND3_X1   g29540(.A1(new_n32501_), .A2(pi0725), .A3(pi1120), .ZN(new_n32796_));
  INV_X1     g29541(.I(pi1120), .ZN(new_n32797_));
  OAI21_X1   g29542(.A1(po0980), .A2(pi0725), .B(new_n32797_), .ZN(new_n32798_));
  NAND3_X1   g29543(.A1(new_n32798_), .A2(new_n32059_), .A3(new_n32796_), .ZN(po0882));
  OAI21_X1   g29544(.A1(new_n32501_), .A2(pi1126), .B(new_n32059_), .ZN(new_n32800_));
  AOI21_X1   g29545(.A1(new_n15463_), .A2(new_n32501_), .B(new_n32800_), .ZN(po0883));
  OAI21_X1   g29546(.A1(new_n32501_), .A2(pi1102), .B(new_n32059_), .ZN(new_n32802_));
  AOI21_X1   g29547(.A1(new_n16128_), .A2(new_n32501_), .B(new_n32802_), .ZN(po0884));
  NAND3_X1   g29548(.A1(new_n32501_), .A2(pi0728), .A3(pi1131), .ZN(new_n32804_));
  OAI21_X1   g29549(.A1(po0980), .A2(pi0728), .B(new_n32149_), .ZN(new_n32805_));
  NAND3_X1   g29550(.A1(new_n32805_), .A2(new_n32059_), .A3(new_n32804_), .ZN(po0885));
  OAI21_X1   g29551(.A1(new_n32501_), .A2(pi1104), .B(new_n32059_), .ZN(new_n32807_));
  AOI21_X1   g29552(.A1(new_n16303_), .A2(new_n32501_), .B(new_n32807_), .ZN(po0886));
  OAI21_X1   g29553(.A1(new_n32501_), .A2(pi1106), .B(new_n32059_), .ZN(new_n32809_));
  AOI21_X1   g29554(.A1(new_n16318_), .A2(new_n32501_), .B(new_n32809_), .ZN(po0887));
  XNOR2_X1   g29555(.A1(pi0721), .A2(pi0813), .ZN(new_n32811_));
  INV_X1     g29556(.I(new_n32811_), .ZN(new_n32812_));
  XNOR2_X1   g29557(.A1(pi0775), .A2(pi0816), .ZN(new_n32813_));
  INV_X1     g29558(.I(new_n32813_), .ZN(new_n32814_));
  NOR2_X1    g29559(.A1(new_n32812_), .A2(new_n32814_), .ZN(new_n32815_));
  XNOR2_X1   g29560(.A1(pi0769), .A2(pi0794), .ZN(new_n32816_));
  NOR2_X1    g29561(.A1(new_n32743_), .A2(pi0795), .ZN(new_n32817_));
  NOR4_X1    g29562(.A1(new_n32815_), .A2(new_n32751_), .A3(new_n32816_), .A4(new_n32817_), .ZN(new_n32818_));
  NAND2_X1   g29563(.A1(new_n32818_), .A2(new_n32741_), .ZN(new_n32819_));
  XOR2_X1    g29564(.A1(pi0721), .A2(pi0813), .Z(new_n32820_));
  NOR2_X1    g29565(.A1(new_n32738_), .A2(new_n32820_), .ZN(new_n32821_));
  NAND3_X1   g29566(.A1(new_n32821_), .A2(pi0795), .A3(new_n32813_), .ZN(new_n32822_));
  NAND2_X1   g29567(.A1(new_n32822_), .A2(pi0731), .ZN(new_n32823_));
  AOI22_X1   g29568(.A1(new_n32823_), .A2(new_n32749_), .B1(new_n32747_), .B2(new_n32819_), .ZN(po0888));
  NAND3_X1   g29569(.A1(new_n32058_), .A2(pi0732), .A3(pi1128), .ZN(new_n32827_));
  OAI21_X1   g29570(.A1(po0954), .A2(pi0732), .B(new_n32543_), .ZN(new_n32828_));
  NAND3_X1   g29571(.A1(new_n32828_), .A2(new_n32059_), .A3(new_n32827_), .ZN(po0889));
  MUX2_X1    g29572(.I0(new_n11967_), .I1(new_n11966_), .S(pi1135), .Z(new_n32830_));
  OAI21_X1   g29573(.A1(new_n32582_), .A2(new_n32830_), .B(new_n10332_), .ZN(new_n32831_));
  OR2_X2     g29574(.A1(pi0838), .A2(pi1136), .Z(new_n32832_));
  NAND2_X1   g29575(.A1(pi0737), .A2(pi1135), .ZN(new_n32833_));
  NAND4_X1   g29576(.A1(new_n32584_), .A2(pi1134), .A3(new_n32832_), .A4(new_n32833_), .ZN(new_n32834_));
  NAND4_X1   g29577(.A1(new_n32831_), .A2(pi0777), .A3(new_n32177_), .A4(new_n32834_), .ZN(new_n32835_));
  NAND2_X1   g29578(.A1(new_n10332_), .A2(pi0424), .ZN(new_n32836_));
  NOR2_X1    g29579(.A1(new_n32836_), .A2(new_n32589_), .ZN(new_n32837_));
  INV_X1     g29580(.I(pi0308), .ZN(new_n32838_));
  NOR2_X1    g29581(.A1(new_n32838_), .A2(pi0200), .ZN(new_n32839_));
  AOI21_X1   g29582(.A1(pi0200), .A2(pi1037), .B(new_n32839_), .ZN(new_n32840_));
  NAND3_X1   g29583(.A1(new_n32840_), .A2(pi0199), .A3(pi1047), .ZN(new_n32841_));
  INV_X1     g29584(.I(new_n32840_), .ZN(new_n32842_));
  OAI21_X1   g29585(.A1(new_n8094_), .A2(pi1047), .B(new_n32842_), .ZN(new_n32843_));
  AOI21_X1   g29586(.A1(new_n32843_), .A2(new_n32841_), .B(new_n25876_), .ZN(new_n32844_));
  NAND2_X1   g29587(.A1(new_n32599_), .A2(pi0375), .ZN(new_n32845_));
  AOI21_X1   g29588(.A1(new_n32601_), .A2(pi0399), .B(pi0590), .ZN(new_n32846_));
  AOI22_X1   g29589(.A1(new_n32846_), .A2(new_n32845_), .B1(pi0316), .B2(new_n32598_), .ZN(new_n32847_));
  NOR3_X1    g29590(.A1(new_n32844_), .A2(pi0588), .A3(new_n32847_), .ZN(new_n32848_));
  OAI21_X1   g29591(.A1(new_n32848_), .A2(new_n32837_), .B(new_n32835_), .ZN(po0890));
  NAND3_X1   g29592(.A1(new_n32501_), .A2(pi0734), .A3(pi1119), .ZN(new_n32850_));
  INV_X1     g29593(.I(pi1119), .ZN(new_n32851_));
  OAI21_X1   g29594(.A1(po0980), .A2(pi0734), .B(new_n32851_), .ZN(new_n32852_));
  NAND3_X1   g29595(.A1(new_n32852_), .A2(new_n32059_), .A3(new_n32850_), .ZN(po0891));
  OAI21_X1   g29596(.A1(new_n32501_), .A2(pi1109), .B(new_n32059_), .ZN(new_n32854_));
  AOI21_X1   g29597(.A1(new_n13638_), .A2(new_n32501_), .B(new_n32854_), .ZN(po0892));
  OAI21_X1   g29598(.A1(new_n32501_), .A2(pi1101), .B(new_n32059_), .ZN(new_n32856_));
  AOI21_X1   g29599(.A1(new_n14611_), .A2(new_n32501_), .B(new_n32856_), .ZN(po0893));
  NAND3_X1   g29600(.A1(new_n32501_), .A2(pi0737), .A3(pi1122), .ZN(new_n32858_));
  INV_X1     g29601(.I(pi1122), .ZN(new_n32859_));
  OAI21_X1   g29602(.A1(po0980), .A2(pi0737), .B(new_n32859_), .ZN(new_n32860_));
  NAND3_X1   g29603(.A1(new_n32860_), .A2(new_n32059_), .A3(new_n32858_), .ZN(po0894));
  NAND3_X1   g29604(.A1(new_n32501_), .A2(pi0738), .A3(pi1121), .ZN(new_n32862_));
  INV_X1     g29605(.I(pi1121), .ZN(new_n32863_));
  OAI21_X1   g29606(.A1(po0980), .A2(pi0738), .B(new_n32863_), .ZN(new_n32864_));
  NAND3_X1   g29607(.A1(new_n32864_), .A2(new_n32059_), .A3(new_n32862_), .ZN(po0895));
  OR3_X2     g29608(.A1(new_n31983_), .A2(pi0952), .A3(pi1061), .Z(new_n32866_));
  NOR2_X1    g29609(.A1(new_n32866_), .A2(new_n13184_), .ZN(po0988));
  OAI21_X1   g29610(.A1(po0988), .A2(pi0739), .B(pi1108), .ZN(new_n32868_));
  INV_X1     g29611(.I(pi1108), .ZN(new_n32869_));
  INV_X1     g29612(.I(po0988), .ZN(new_n32870_));
  NAND3_X1   g29613(.A1(new_n32870_), .A2(pi0739), .A3(new_n32869_), .ZN(new_n32871_));
  NAND3_X1   g29614(.A1(new_n32871_), .A2(new_n31978_), .A3(new_n32868_), .ZN(po0896));
  AOI21_X1   g29615(.A1(new_n32870_), .A2(new_n15815_), .B(pi0966), .ZN(new_n32873_));
  NOR3_X1    g29616(.A1(new_n32873_), .A2(new_n32113_), .A3(new_n32870_), .ZN(po0898));
  AOI21_X1   g29617(.A1(new_n32870_), .A2(new_n15764_), .B(pi0966), .ZN(new_n32875_));
  NOR3_X1    g29618(.A1(new_n32875_), .A2(new_n32086_), .A3(new_n32870_), .ZN(po0899));
  OAI21_X1   g29619(.A1(po0988), .A2(pi0743), .B(pi1109), .ZN(new_n32877_));
  INV_X1     g29620(.I(pi1109), .ZN(new_n32878_));
  NAND3_X1   g29621(.A1(new_n32870_), .A2(pi0743), .A3(new_n32878_), .ZN(new_n32879_));
  NAND3_X1   g29622(.A1(new_n32879_), .A2(new_n31978_), .A3(new_n32877_), .ZN(po0900));
  OR2_X2     g29623(.A1(po0988), .A2(pi0744), .Z(new_n32881_));
  NAND2_X1   g29624(.A1(po0988), .A2(pi1131), .ZN(new_n32882_));
  AOI21_X1   g29625(.A1(new_n32881_), .A2(new_n31978_), .B(new_n32882_), .ZN(po0901));
  AOI21_X1   g29626(.A1(new_n32870_), .A2(new_n15596_), .B(pi0966), .ZN(new_n32884_));
  NOR3_X1    g29627(.A1(new_n32884_), .A2(new_n32547_), .A3(new_n32870_), .ZN(po0902));
  OAI21_X1   g29628(.A1(po0988), .A2(pi0746), .B(pi1104), .ZN(new_n32886_));
  NAND3_X1   g29629(.A1(new_n32870_), .A2(pi0746), .A3(new_n31998_), .ZN(new_n32887_));
  NAND3_X1   g29630(.A1(new_n32887_), .A2(new_n31978_), .A3(new_n32886_), .ZN(po0903));
  INV_X1     g29631(.I(new_n32749_), .ZN(new_n32889_));
  NAND2_X1   g29632(.A1(new_n32889_), .A2(pi0773), .ZN(new_n32890_));
  NOR2_X1    g29633(.A1(new_n32724_), .A2(new_n32890_), .ZN(new_n32891_));
  XNOR2_X1   g29634(.A1(pi0773), .A2(pi0801), .ZN(new_n32892_));
  OAI22_X1   g29635(.A1(new_n32891_), .A2(new_n32892_), .B1(new_n32743_), .B2(new_n32730_), .ZN(new_n32893_));
  INV_X1     g29636(.I(new_n32815_), .ZN(new_n32894_));
  NAND2_X1   g29637(.A1(new_n32894_), .A2(new_n32762_), .ZN(new_n32895_));
  NOR2_X1    g29638(.A1(new_n32895_), .A2(new_n32740_), .ZN(new_n32896_));
  NOR2_X1    g29639(.A1(new_n32896_), .A2(new_n32816_), .ZN(new_n32897_));
  XOR2_X1    g29640(.A1(new_n32890_), .A2(pi0747), .Z(new_n32898_));
  AOI21_X1   g29641(.A1(new_n32897_), .A2(new_n32893_), .B(new_n32898_), .ZN(po0904));
  OAI21_X1   g29642(.A1(po0988), .A2(pi0748), .B(pi1106), .ZN(new_n32900_));
  INV_X1     g29643(.I(pi1106), .ZN(new_n32901_));
  NAND3_X1   g29644(.A1(new_n32870_), .A2(pi0748), .A3(new_n32901_), .ZN(new_n32902_));
  NAND3_X1   g29645(.A1(new_n32902_), .A2(new_n31978_), .A3(new_n32900_), .ZN(po0905));
  OAI21_X1   g29646(.A1(po0988), .A2(pi0749), .B(pi1105), .ZN(new_n32904_));
  NAND3_X1   g29647(.A1(new_n32870_), .A2(pi0749), .A3(new_n32033_), .ZN(new_n32905_));
  NAND3_X1   g29648(.A1(new_n32905_), .A2(new_n31978_), .A3(new_n32904_), .ZN(po0906));
  OR2_X2     g29649(.A1(po0988), .A2(pi0750), .Z(new_n32907_));
  NAND2_X1   g29650(.A1(po0988), .A2(pi1130), .ZN(new_n32908_));
  AOI21_X1   g29651(.A1(new_n32907_), .A2(new_n31978_), .B(new_n32908_), .ZN(po0907));
  AOI21_X1   g29652(.A1(new_n32870_), .A2(new_n15546_), .B(pi0966), .ZN(new_n32910_));
  NOR3_X1    g29653(.A1(new_n32910_), .A2(new_n32564_), .A3(new_n32870_), .ZN(po0908));
  AOI21_X1   g29654(.A1(new_n32870_), .A2(new_n16089_), .B(pi0966), .ZN(new_n32912_));
  NOR3_X1    g29655(.A1(new_n32912_), .A2(new_n32142_), .A3(new_n32870_), .ZN(po0909));
  AOI21_X1   g29656(.A1(new_n32870_), .A2(new_n15866_), .B(pi0966), .ZN(new_n32914_));
  NOR3_X1    g29657(.A1(new_n32914_), .A2(new_n32568_), .A3(new_n32870_), .ZN(po0910));
  AOI21_X1   g29658(.A1(new_n32870_), .A2(new_n15896_), .B(pi0966), .ZN(new_n32916_));
  NOR3_X1    g29659(.A1(new_n32916_), .A2(new_n32607_), .A3(new_n32870_), .ZN(po0911));
  AOI21_X1   g29660(.A1(new_n32870_), .A2(new_n15509_), .B(pi0966), .ZN(new_n32918_));
  NOR3_X1    g29661(.A1(new_n32918_), .A2(new_n32797_), .A3(new_n32870_), .ZN(po0912));
  AOI21_X1   g29662(.A1(new_n32870_), .A2(new_n15926_), .B(pi0966), .ZN(new_n32920_));
  NOR3_X1    g29663(.A1(new_n32920_), .A2(new_n32851_), .A3(new_n32870_), .ZN(po0913));
  AOI21_X1   g29664(.A1(new_n32870_), .A2(new_n15787_), .B(pi0966), .ZN(new_n32922_));
  NOR3_X1    g29665(.A1(new_n32922_), .A2(new_n32073_), .A3(new_n32870_), .ZN(po0914));
  OAI21_X1   g29666(.A1(po0988), .A2(pi0758), .B(pi1101), .ZN(new_n32924_));
  INV_X1     g29667(.I(pi1101), .ZN(new_n32925_));
  NAND3_X1   g29668(.A1(new_n32870_), .A2(pi0758), .A3(new_n32925_), .ZN(new_n32926_));
  NAND3_X1   g29669(.A1(new_n32926_), .A2(new_n31978_), .A3(new_n32924_), .ZN(po0915));
  NOR3_X1    g29670(.A1(new_n32866_), .A2(new_n13184_), .A3(pi1100), .ZN(new_n32928_));
  NOR2_X1    g29671(.A1(po0988), .A2(pi0759), .ZN(new_n32929_));
  OAI21_X1   g29672(.A1(new_n32929_), .A2(new_n32928_), .B(new_n31978_), .ZN(po0916));
  AOI21_X1   g29673(.A1(new_n32870_), .A2(new_n15831_), .B(pi0966), .ZN(new_n32931_));
  NOR3_X1    g29674(.A1(new_n32931_), .A2(new_n32078_), .A3(new_n32870_), .ZN(po0917));
  AOI21_X1   g29675(.A1(new_n32870_), .A2(new_n12116_), .B(pi0966), .ZN(new_n32933_));
  NOR3_X1    g29676(.A1(new_n32933_), .A2(new_n32863_), .A3(new_n32870_), .ZN(po0918));
  OR2_X2     g29677(.A1(po0988), .A2(pi0762), .Z(new_n32935_));
  NAND2_X1   g29678(.A1(po0988), .A2(pi1129), .ZN(new_n32936_));
  AOI21_X1   g29679(.A1(new_n32935_), .A2(new_n31978_), .B(new_n32936_), .ZN(po0919));
  OAI21_X1   g29680(.A1(po0988), .A2(pi0763), .B(pi1103), .ZN(new_n32938_));
  INV_X1     g29681(.I(pi1103), .ZN(new_n32939_));
  NAND3_X1   g29682(.A1(new_n32870_), .A2(pi0763), .A3(new_n32939_), .ZN(new_n32940_));
  NAND3_X1   g29683(.A1(new_n32940_), .A2(new_n31978_), .A3(new_n32938_), .ZN(po0920));
  OAI21_X1   g29684(.A1(po0988), .A2(pi0764), .B(pi1107), .ZN(new_n32942_));
  INV_X1     g29685(.I(pi1107), .ZN(new_n32943_));
  NAND3_X1   g29686(.A1(new_n32870_), .A2(pi0764), .A3(new_n32943_), .ZN(new_n32944_));
  NAND3_X1   g29687(.A1(new_n32944_), .A2(new_n31978_), .A3(new_n32942_), .ZN(po0921));
  NOR2_X1    g29688(.A1(new_n32738_), .A2(new_n32895_), .ZN(po0978));
  NOR3_X1    g29689(.A1(po0978), .A2(new_n32728_), .A3(new_n32748_), .ZN(po0922));
  OAI21_X1   g29690(.A1(po0988), .A2(pi0766), .B(pi1110), .ZN(new_n32948_));
  INV_X1     g29691(.I(pi1110), .ZN(new_n32949_));
  NAND3_X1   g29692(.A1(new_n32870_), .A2(pi0766), .A3(new_n32949_), .ZN(new_n32950_));
  NAND3_X1   g29693(.A1(new_n32950_), .A2(new_n31978_), .A3(new_n32948_), .ZN(po0923));
  AOI21_X1   g29694(.A1(new_n32870_), .A2(new_n15145_), .B(pi0966), .ZN(new_n32952_));
  NOR3_X1    g29695(.A1(new_n32952_), .A2(new_n32556_), .A3(new_n32870_), .ZN(po0924));
  AOI21_X1   g29696(.A1(new_n32870_), .A2(new_n16201_), .B(pi0966), .ZN(new_n32954_));
  NOR3_X1    g29697(.A1(new_n32954_), .A2(new_n32291_), .A3(new_n32870_), .ZN(po0925));
  INV_X1     g29698(.I(pi0769), .ZN(new_n32956_));
  NOR2_X1    g29699(.A1(new_n32740_), .A2(new_n32742_), .ZN(new_n32957_));
  NOR4_X1    g29700(.A1(new_n32732_), .A2(new_n32815_), .A3(new_n32892_), .A4(new_n32957_), .ZN(new_n32958_));
  NAND4_X1   g29701(.A1(new_n32958_), .A2(new_n32956_), .A3(new_n32757_), .A4(new_n32762_), .ZN(new_n32959_));
  INV_X1     g29702(.I(new_n32958_), .ZN(new_n32960_));
  NAND2_X1   g29703(.A1(new_n32821_), .A2(pi0816), .ZN(new_n32961_));
  AOI21_X1   g29704(.A1(new_n32746_), .A2(new_n32960_), .B(new_n32961_), .ZN(new_n32962_));
  NAND3_X1   g29705(.A1(new_n32961_), .A2(new_n32746_), .A3(new_n32958_), .ZN(new_n32963_));
  NAND2_X1   g29706(.A1(new_n32751_), .A2(pi0775), .ZN(new_n32964_));
  XOR2_X1    g29707(.A1(new_n32964_), .A2(new_n32956_), .Z(new_n32965_));
  AOI21_X1   g29708(.A1(new_n32965_), .A2(new_n32750_), .B(new_n32766_), .ZN(new_n32966_));
  NAND2_X1   g29709(.A1(new_n32963_), .A2(new_n32966_), .ZN(new_n32967_));
  OAI21_X1   g29710(.A1(new_n32967_), .A2(new_n32962_), .B(new_n32959_), .ZN(po0926));
  AOI21_X1   g29711(.A1(new_n32870_), .A2(new_n15427_), .B(pi0966), .ZN(new_n32969_));
  NOR3_X1    g29712(.A1(new_n32969_), .A2(new_n32121_), .A3(new_n32870_), .ZN(po0927));
  NAND2_X1   g29713(.A1(pi0771), .A2(pi0945), .ZN(new_n32971_));
  NAND2_X1   g29714(.A1(pi0731), .A2(pi0795), .ZN(new_n32972_));
  INV_X1     g29715(.I(new_n32735_), .ZN(new_n32973_));
  INV_X1     g29716(.I(new_n32892_), .ZN(new_n32974_));
  NOR2_X1    g29717(.A1(new_n32725_), .A2(new_n32721_), .ZN(new_n32975_));
  AOI21_X1   g29718(.A1(pi0771), .A2(pi0800), .B(pi0765), .ZN(new_n32976_));
  OR3_X2     g29719(.A1(new_n32976_), .A2(new_n32956_), .A3(new_n32742_), .Z(new_n32977_));
  OAI21_X1   g29720(.A1(new_n32975_), .A2(new_n32977_), .B(pi0773), .ZN(new_n32978_));
  OAI21_X1   g29721(.A1(new_n32973_), .A2(new_n32978_), .B(new_n32974_), .ZN(new_n32979_));
  NOR2_X1    g29722(.A1(new_n32758_), .A2(pi0721), .ZN(new_n32980_));
  AOI21_X1   g29723(.A1(new_n32979_), .A2(new_n32980_), .B(new_n32759_), .ZN(new_n32981_));
  NAND2_X1   g29724(.A1(new_n32747_), .A2(new_n32766_), .ZN(new_n32982_));
  OAI22_X1   g29725(.A1(new_n32981_), .A2(new_n32982_), .B1(new_n32814_), .B2(new_n32972_), .ZN(new_n32983_));
  AND2_X2    g29726(.A1(new_n32983_), .A2(new_n32821_), .Z(po0963));
  NOR2_X1    g29727(.A1(po0963), .A2(pi0945), .ZN(new_n32985_));
  OAI22_X1   g29728(.A1(new_n32985_), .A2(pi0987), .B1(po0978), .B2(new_n32971_), .ZN(po0928));
  OAI21_X1   g29729(.A1(po0988), .A2(pi0772), .B(pi1102), .ZN(new_n32987_));
  INV_X1     g29730(.I(pi1102), .ZN(new_n32988_));
  NAND3_X1   g29731(.A1(new_n32870_), .A2(pi0772), .A3(new_n32988_), .ZN(new_n32989_));
  NAND3_X1   g29732(.A1(new_n32989_), .A2(new_n31978_), .A3(new_n32987_), .ZN(po0929));
  NAND3_X1   g29733(.A1(po0963), .A2(new_n32743_), .A3(new_n32973_), .ZN(new_n32991_));
  AOI21_X1   g29734(.A1(pi0801), .A2(new_n32895_), .B(new_n32738_), .ZN(new_n32992_));
  XOR2_X1    g29735(.A1(new_n32749_), .A2(pi0773), .Z(new_n32993_));
  OAI21_X1   g29736(.A1(new_n32992_), .A2(new_n32889_), .B(new_n32993_), .ZN(new_n32994_));
  AOI21_X1   g29737(.A1(new_n32991_), .A2(new_n32889_), .B(new_n32994_), .ZN(po0930));
  AOI21_X1   g29738(.A1(new_n32870_), .A2(new_n14348_), .B(pi0966), .ZN(new_n32996_));
  NOR3_X1    g29739(.A1(new_n32996_), .A2(new_n32125_), .A3(new_n32870_), .ZN(po0931));
  NAND3_X1   g29740(.A1(new_n32751_), .A2(pi0765), .A3(pi0771), .ZN(new_n32998_));
  NAND2_X1   g29741(.A1(new_n32822_), .A2(new_n32998_), .ZN(new_n32999_));
  NOR3_X1    g29742(.A1(new_n32747_), .A2(new_n32746_), .A3(pi0945), .ZN(new_n33000_));
  NOR2_X1    g29743(.A1(new_n32747_), .A2(pi0945), .ZN(new_n33001_));
  NAND4_X1   g29744(.A1(new_n32717_), .A2(pi0795), .A3(pi0800), .A4(pi0801), .ZN(new_n33002_));
  NOR2_X1    g29745(.A1(new_n32812_), .A2(new_n33002_), .ZN(new_n33003_));
  AOI21_X1   g29746(.A1(new_n32734_), .A2(new_n33003_), .B(new_n32998_), .ZN(new_n33004_));
  OAI21_X1   g29747(.A1(new_n33004_), .A2(pi0775), .B(new_n33001_), .ZN(new_n33005_));
  OAI21_X1   g29748(.A1(new_n32738_), .A2(new_n32895_), .B(pi0775), .ZN(new_n33006_));
  AOI22_X1   g29749(.A1(new_n32999_), .A2(new_n33000_), .B1(new_n33005_), .B2(new_n33006_), .ZN(po0932));
  AOI21_X1   g29750(.A1(new_n32870_), .A2(new_n32770_), .B(pi0966), .ZN(new_n33008_));
  NOR3_X1    g29751(.A1(new_n33008_), .A2(new_n32543_), .A3(new_n32870_), .ZN(po0933));
  AOI21_X1   g29752(.A1(new_n32870_), .A2(new_n16049_), .B(pi0966), .ZN(new_n33010_));
  NOR3_X1    g29753(.A1(new_n33010_), .A2(new_n32859_), .A3(new_n32870_), .ZN(po0934));
  NOR2_X1    g29754(.A1(pi1046), .A2(pi1083), .ZN(new_n33012_));
  NAND4_X1   g29755(.A1(new_n33012_), .A2(pi0832), .A3(pi0956), .A4(pi1085), .ZN(new_n33013_));
  NOR2_X1    g29756(.A1(new_n33013_), .A2(pi0968), .ZN(new_n33014_));
  NAND2_X1   g29757(.A1(new_n33014_), .A2(pi1100), .ZN(new_n33015_));
  OAI21_X1   g29758(.A1(new_n11891_), .A2(new_n33014_), .B(new_n33015_), .ZN(po0935));
  NOR2_X1    g29759(.A1(new_n32025_), .A2(pi0779), .ZN(po0936));
  NOR2_X1    g29760(.A1(new_n31963_), .A2(pi0780), .ZN(po0937));
  NAND2_X1   g29761(.A1(new_n33014_), .A2(pi1101), .ZN(new_n33019_));
  OAI21_X1   g29762(.A1(new_n11969_), .A2(new_n33014_), .B(new_n33019_), .ZN(po0938));
  NAND4_X1   g29763(.A1(new_n31962_), .A2(new_n2587_), .A3(pi0983), .A4(new_n29015_), .ZN(po0939));
  INV_X1     g29764(.I(pi0783), .ZN(new_n33022_));
  NAND2_X1   g29765(.A1(new_n33014_), .A2(pi1109), .ZN(new_n33023_));
  OAI21_X1   g29766(.A1(new_n33022_), .A2(new_n33014_), .B(new_n33023_), .ZN(po0940));
  INV_X1     g29767(.I(pi0784), .ZN(new_n33025_));
  NAND2_X1   g29768(.A1(new_n33014_), .A2(pi1110), .ZN(new_n33026_));
  OAI21_X1   g29769(.A1(new_n33025_), .A2(new_n33014_), .B(new_n33026_), .ZN(po0941));
  NAND2_X1   g29770(.A1(new_n33014_), .A2(pi1102), .ZN(new_n33028_));
  OAI21_X1   g29771(.A1(new_n11870_), .A2(new_n33014_), .B(new_n33028_), .ZN(po0942));
  NAND2_X1   g29772(.A1(new_n7876_), .A2(pi0954), .ZN(new_n33030_));
  OAI21_X1   g29773(.A1(pi0024), .A2(pi0954), .B(new_n33030_), .ZN(po0943));
  NAND2_X1   g29774(.A1(new_n33014_), .A2(pi1104), .ZN(new_n33032_));
  OAI21_X1   g29775(.A1(new_n12048_), .A2(new_n33014_), .B(new_n33032_), .ZN(po0944));
  NAND2_X1   g29776(.A1(new_n33014_), .A2(pi1105), .ZN(new_n33034_));
  OAI21_X1   g29777(.A1(new_n11986_), .A2(new_n33014_), .B(new_n33034_), .ZN(po0945));
  NAND2_X1   g29778(.A1(new_n33014_), .A2(pi1106), .ZN(new_n33036_));
  OAI21_X1   g29779(.A1(new_n11985_), .A2(new_n33014_), .B(new_n33036_), .ZN(po0946));
  NAND2_X1   g29780(.A1(new_n33014_), .A2(pi1107), .ZN(new_n33038_));
  OAI21_X1   g29781(.A1(new_n11867_), .A2(new_n33014_), .B(new_n33038_), .ZN(po0947));
  INV_X1     g29782(.I(pi0791), .ZN(new_n33040_));
  NAND2_X1   g29783(.A1(new_n33014_), .A2(pi1108), .ZN(new_n33041_));
  OAI21_X1   g29784(.A1(new_n33040_), .A2(new_n33014_), .B(new_n33041_), .ZN(po0948));
  NAND2_X1   g29785(.A1(new_n33014_), .A2(pi1103), .ZN(new_n33043_));
  OAI21_X1   g29786(.A1(new_n11868_), .A2(new_n33014_), .B(new_n33043_), .ZN(po0949));
  INV_X1     g29787(.I(new_n26268_), .ZN(po0950));
  INV_X1     g29788(.I(pi0968), .ZN(new_n33046_));
  NOR2_X1    g29789(.A1(new_n33013_), .A2(new_n33046_), .ZN(new_n33047_));
  NAND2_X1   g29790(.A1(new_n33047_), .A2(pi1130), .ZN(new_n33048_));
  OAI21_X1   g29791(.A1(new_n32742_), .A2(new_n33047_), .B(new_n33048_), .ZN(po0951));
  NAND2_X1   g29792(.A1(new_n33047_), .A2(pi1128), .ZN(new_n33050_));
  OAI21_X1   g29793(.A1(new_n32766_), .A2(new_n33047_), .B(new_n33050_), .ZN(po0952));
  INV_X1     g29794(.I(new_n32155_), .ZN(new_n33052_));
  NOR4_X1    g29795(.A1(new_n33052_), .A2(pi0269), .A3(po1130), .A4(new_n4711_), .ZN(new_n33053_));
  NAND3_X1   g29796(.A1(new_n33053_), .A2(new_n4119_), .A3(new_n32158_), .ZN(new_n33054_));
  XOR2_X1    g29797(.A1(new_n33054_), .A2(new_n29593_), .Z(po0953));
  NAND2_X1   g29798(.A1(new_n33047_), .A2(pi1124), .ZN(new_n33056_));
  OAI21_X1   g29799(.A1(new_n32726_), .A2(new_n33047_), .B(new_n33056_), .ZN(po0955));
  NAND2_X1   g29800(.A1(new_n33047_), .A2(pi1107), .ZN(new_n33058_));
  OAI21_X1   g29801(.A1(pi0799), .A2(new_n33047_), .B(new_n33058_), .ZN(po0956));
  INV_X1     g29802(.I(pi0800), .ZN(new_n33060_));
  NAND2_X1   g29803(.A1(new_n33047_), .A2(pi1125), .ZN(new_n33061_));
  OAI21_X1   g29804(.A1(new_n33060_), .A2(new_n33047_), .B(new_n33061_), .ZN(po0957));
  NAND2_X1   g29805(.A1(new_n33047_), .A2(pi1126), .ZN(new_n33063_));
  OAI21_X1   g29806(.A1(new_n32743_), .A2(new_n33047_), .B(new_n33063_), .ZN(po0958));
  NOR4_X1    g29807(.A1(new_n32159_), .A2(pi0264), .A3(pi0265), .A4(pi0274), .ZN(po0959));
  NAND2_X1   g29808(.A1(new_n33047_), .A2(pi1106), .ZN(new_n33066_));
  OAI21_X1   g29809(.A1(pi0803), .A2(new_n33047_), .B(new_n33066_), .ZN(po0960));
  NAND2_X1   g29810(.A1(new_n33047_), .A2(pi1109), .ZN(new_n33068_));
  OAI21_X1   g29811(.A1(new_n30832_), .A2(new_n33047_), .B(new_n33068_), .ZN(po0961));
  INV_X1     g29812(.I(new_n32157_), .ZN(new_n33070_));
  NOR2_X1    g29813(.A1(new_n33070_), .A2(pi0282), .ZN(new_n33071_));
  INV_X1     g29814(.I(pi0282), .ZN(new_n33072_));
  NAND2_X1   g29815(.A1(new_n33072_), .A2(pi0270), .ZN(new_n33073_));
  OAI22_X1   g29816(.A1(new_n33071_), .A2(pi0270), .B1(new_n33070_), .B2(new_n33073_), .ZN(po0962));
  NAND2_X1   g29817(.A1(new_n33047_), .A2(pi1127), .ZN(new_n33075_));
  OAI21_X1   g29818(.A1(new_n32722_), .A2(new_n33047_), .B(new_n33075_), .ZN(po0964));
  INV_X1     g29819(.I(pi0808), .ZN(new_n33077_));
  NAND2_X1   g29820(.A1(new_n33047_), .A2(pi1101), .ZN(new_n33078_));
  OAI21_X1   g29821(.A1(new_n33077_), .A2(new_n33047_), .B(new_n33078_), .ZN(po0965));
  NAND2_X1   g29822(.A1(new_n33047_), .A2(pi1103), .ZN(new_n33080_));
  OAI21_X1   g29823(.A1(pi0809), .A2(new_n33047_), .B(new_n33080_), .ZN(po0966));
  NAND2_X1   g29824(.A1(new_n33047_), .A2(pi1108), .ZN(new_n33082_));
  OAI21_X1   g29825(.A1(new_n30833_), .A2(new_n33047_), .B(new_n33082_), .ZN(po0967));
  INV_X1     g29826(.I(pi0811), .ZN(new_n33084_));
  NAND2_X1   g29827(.A1(new_n33047_), .A2(pi1102), .ZN(new_n33085_));
  OAI21_X1   g29828(.A1(new_n33084_), .A2(new_n33047_), .B(new_n33085_), .ZN(po0968));
  NAND2_X1   g29829(.A1(new_n33047_), .A2(pi1104), .ZN(new_n33087_));
  OAI21_X1   g29830(.A1(pi0812), .A2(new_n33047_), .B(new_n33087_), .ZN(po0969));
  NAND2_X1   g29831(.A1(new_n33047_), .A2(pi1131), .ZN(new_n33089_));
  OAI21_X1   g29832(.A1(new_n32719_), .A2(new_n33047_), .B(new_n33089_), .ZN(po0970));
  NAND2_X1   g29833(.A1(new_n33047_), .A2(pi1105), .ZN(new_n33091_));
  OAI21_X1   g29834(.A1(pi0814), .A2(new_n33047_), .B(new_n33091_), .ZN(po0971));
  NAND2_X1   g29835(.A1(new_n33047_), .A2(pi1110), .ZN(new_n33093_));
  OAI21_X1   g29836(.A1(new_n30830_), .A2(new_n33047_), .B(new_n33093_), .ZN(po0972));
  NAND2_X1   g29837(.A1(new_n33047_), .A2(pi1129), .ZN(new_n33095_));
  OAI21_X1   g29838(.A1(new_n32717_), .A2(new_n33047_), .B(new_n33095_), .ZN(po0973));
  XOR2_X1    g29839(.A1(new_n32156_), .A2(pi0269), .Z(po0974));
  OAI21_X1   g29840(.A1(new_n10370_), .A2(new_n10332_), .B(new_n10255_), .ZN(po0975));
  NOR2_X1    g29841(.A1(new_n32159_), .A2(pi0264), .ZN(new_n33099_));
  NAND2_X1   g29842(.A1(new_n29593_), .A2(pi0265), .ZN(new_n33100_));
  OAI22_X1   g29843(.A1(new_n33099_), .A2(pi0265), .B1(new_n32159_), .B2(new_n33100_), .ZN(po0976));
  AOI21_X1   g29844(.A1(new_n29936_), .A2(new_n33072_), .B(new_n32157_), .ZN(new_n33102_));
  XOR2_X1    g29845(.A1(new_n33102_), .A2(pi0277), .Z(po0977));
  NOR2_X1    g29846(.A1(pi0811), .A2(pi0893), .ZN(po0979));
  NOR2_X1    g29847(.A1(new_n7757_), .A2(pi0982), .ZN(new_n33105_));
  OAI21_X1   g29848(.A1(new_n9141_), .A2(new_n10332_), .B(new_n2955_), .ZN(new_n33106_));
  NOR2_X1    g29849(.A1(new_n33105_), .A2(new_n33106_), .ZN(po0981));
  INV_X1     g29850(.I(pi0825), .ZN(po1147));
  INV_X1     g29851(.I(pi0123), .ZN(new_n33109_));
  NOR2_X1    g29852(.A1(new_n3590_), .A2(new_n33109_), .ZN(new_n33110_));
  INV_X1     g29853(.I(new_n33110_), .ZN(new_n33111_));
  NOR2_X1    g29854(.A1(new_n33111_), .A2(po1147), .ZN(new_n33112_));
  AOI21_X1   g29855(.A1(new_n32125_), .A2(new_n32149_), .B(new_n33110_), .ZN(new_n33113_));
  OR2_X2     g29856(.A1(new_n33112_), .A2(new_n33113_), .Z(new_n33114_));
  XOR2_X1    g29857(.A1(pi1125), .A2(pi1126), .Z(new_n33115_));
  XOR2_X1    g29858(.A1(new_n33115_), .A2(new_n32539_), .Z(new_n33116_));
  XOR2_X1    g29859(.A1(new_n33116_), .A2(pi1128), .Z(new_n33117_));
  XOR2_X1    g29860(.A1(pi1124), .A2(pi1130), .Z(new_n33118_));
  INV_X1     g29861(.I(new_n33118_), .ZN(new_n33119_));
  XNOR2_X1   g29862(.A1(pi1124), .A2(pi1130), .ZN(new_n33120_));
  NOR2_X1    g29863(.A1(new_n33117_), .A2(new_n33120_), .ZN(new_n33121_));
  AOI21_X1   g29864(.A1(new_n33117_), .A2(new_n33119_), .B(new_n33121_), .ZN(new_n33122_));
  INV_X1     g29865(.I(new_n33122_), .ZN(new_n33123_));
  NAND4_X1   g29866(.A1(new_n33122_), .A2(pi1127), .A3(pi1131), .A4(new_n33111_), .ZN(new_n33124_));
  NAND3_X1   g29867(.A1(new_n33111_), .A2(pi1127), .A3(pi1131), .ZN(new_n33125_));
  NAND4_X1   g29868(.A1(new_n33112_), .A2(new_n32125_), .A3(new_n32149_), .A4(new_n33111_), .ZN(new_n33126_));
  OAI21_X1   g29869(.A1(new_n33125_), .A2(new_n33126_), .B(new_n33123_), .ZN(new_n33127_));
  AOI22_X1   g29870(.A1(new_n33127_), .A2(new_n33124_), .B1(new_n33114_), .B2(new_n33123_), .ZN(po0982));
  INV_X1     g29871(.I(pi0826), .ZN(po1148));
  NOR2_X1    g29872(.A1(new_n33111_), .A2(po1148), .ZN(new_n33130_));
  AOI21_X1   g29873(.A1(new_n32859_), .A2(new_n32564_), .B(new_n33110_), .ZN(new_n33131_));
  OR2_X2     g29874(.A1(new_n33130_), .A2(new_n33131_), .Z(new_n33132_));
  XOR2_X1    g29875(.A1(pi1116), .A2(pi1117), .Z(new_n33133_));
  XOR2_X1    g29876(.A1(new_n33133_), .A2(new_n32863_), .Z(new_n33134_));
  XOR2_X1    g29877(.A1(new_n33134_), .A2(pi1120), .Z(new_n33135_));
  XOR2_X1    g29878(.A1(pi1118), .A2(pi1119), .Z(new_n33136_));
  INV_X1     g29879(.I(new_n33136_), .ZN(new_n33137_));
  XNOR2_X1   g29880(.A1(pi1118), .A2(pi1119), .ZN(new_n33138_));
  NOR2_X1    g29881(.A1(new_n33135_), .A2(new_n33138_), .ZN(new_n33139_));
  AOI21_X1   g29882(.A1(new_n33135_), .A2(new_n33137_), .B(new_n33139_), .ZN(new_n33140_));
  INV_X1     g29883(.I(new_n33140_), .ZN(new_n33141_));
  NAND4_X1   g29884(.A1(new_n33140_), .A2(pi1122), .A3(pi1123), .A4(new_n33111_), .ZN(new_n33142_));
  NAND3_X1   g29885(.A1(new_n33111_), .A2(pi1122), .A3(pi1123), .ZN(new_n33143_));
  NAND4_X1   g29886(.A1(new_n33130_), .A2(new_n32859_), .A3(new_n32564_), .A4(new_n33111_), .ZN(new_n33144_));
  OAI21_X1   g29887(.A1(new_n33143_), .A2(new_n33144_), .B(new_n33141_), .ZN(new_n33145_));
  AOI22_X1   g29888(.A1(new_n33145_), .A2(new_n33142_), .B1(new_n33132_), .B2(new_n33141_), .ZN(po0983));
  INV_X1     g29889(.I(pi0827), .ZN(po1178));
  NOR2_X1    g29890(.A1(new_n33111_), .A2(po1178), .ZN(new_n33148_));
  INV_X1     g29891(.I(pi1100), .ZN(new_n33149_));
  AOI21_X1   g29892(.A1(new_n33149_), .A2(new_n32943_), .B(new_n33110_), .ZN(new_n33150_));
  OR2_X2     g29893(.A1(new_n33148_), .A2(new_n33150_), .Z(new_n33151_));
  XOR2_X1    g29894(.A1(pi1101), .A2(pi1102), .Z(new_n33152_));
  XOR2_X1    g29895(.A1(new_n33152_), .A2(new_n32901_), .Z(new_n33153_));
  XOR2_X1    g29896(.A1(new_n33153_), .A2(pi1104), .Z(new_n33154_));
  XOR2_X1    g29897(.A1(pi1103), .A2(pi1105), .Z(new_n33155_));
  INV_X1     g29898(.I(new_n33155_), .ZN(new_n33156_));
  XNOR2_X1   g29899(.A1(pi1103), .A2(pi1105), .ZN(new_n33157_));
  NOR2_X1    g29900(.A1(new_n33154_), .A2(new_n33157_), .ZN(new_n33158_));
  AOI21_X1   g29901(.A1(new_n33154_), .A2(new_n33156_), .B(new_n33158_), .ZN(new_n33159_));
  INV_X1     g29902(.I(new_n33159_), .ZN(new_n33160_));
  NAND4_X1   g29903(.A1(new_n33159_), .A2(pi1100), .A3(pi1107), .A4(new_n33111_), .ZN(new_n33161_));
  NAND3_X1   g29904(.A1(new_n33111_), .A2(pi1100), .A3(pi1107), .ZN(new_n33162_));
  NAND4_X1   g29905(.A1(new_n33148_), .A2(new_n33149_), .A3(new_n32943_), .A4(new_n33111_), .ZN(new_n33163_));
  OAI21_X1   g29906(.A1(new_n33162_), .A2(new_n33163_), .B(new_n33160_), .ZN(new_n33164_));
  AOI22_X1   g29907(.A1(new_n33164_), .A2(new_n33161_), .B1(new_n33151_), .B2(new_n33160_), .ZN(po0984));
  INV_X1     g29908(.I(pi0828), .ZN(po1182));
  NOR2_X1    g29909(.A1(new_n33111_), .A2(po1182), .ZN(new_n33167_));
  AOI21_X1   g29910(.A1(new_n32113_), .A2(new_n32078_), .B(new_n33110_), .ZN(new_n33168_));
  OR2_X2     g29911(.A1(new_n33167_), .A2(new_n33168_), .Z(new_n33169_));
  XOR2_X1    g29912(.A1(pi1108), .A2(pi1109), .Z(new_n33170_));
  XOR2_X1    g29913(.A1(new_n33170_), .A2(new_n32073_), .Z(new_n33171_));
  XOR2_X1    g29914(.A1(new_n33171_), .A2(pi1112), .Z(new_n33172_));
  XOR2_X1    g29915(.A1(pi1110), .A2(pi1111), .Z(new_n33173_));
  INV_X1     g29916(.I(new_n33173_), .ZN(new_n33174_));
  XNOR2_X1   g29917(.A1(pi1110), .A2(pi1111), .ZN(new_n33175_));
  NOR2_X1    g29918(.A1(new_n33172_), .A2(new_n33175_), .ZN(new_n33176_));
  AOI21_X1   g29919(.A1(new_n33172_), .A2(new_n33174_), .B(new_n33176_), .ZN(new_n33177_));
  INV_X1     g29920(.I(new_n33177_), .ZN(new_n33178_));
  NAND4_X1   g29921(.A1(new_n33177_), .A2(pi1114), .A3(pi1115), .A4(new_n33111_), .ZN(new_n33179_));
  NAND3_X1   g29922(.A1(new_n33111_), .A2(pi1114), .A3(pi1115), .ZN(new_n33180_));
  NAND4_X1   g29923(.A1(new_n33167_), .A2(new_n32113_), .A3(new_n32078_), .A4(new_n33111_), .ZN(new_n33181_));
  OAI21_X1   g29924(.A1(new_n33180_), .A2(new_n33181_), .B(new_n33178_), .ZN(new_n33182_));
  AOI22_X1   g29925(.A1(new_n33182_), .A2(new_n33179_), .B1(new_n33169_), .B2(new_n33178_), .ZN(po0985));
  NOR4_X1    g29926(.A1(new_n7756_), .A2(pi0951), .A3(pi1092), .A4(new_n10332_), .ZN(po0986));
  XOR2_X1    g29927(.A1(new_n33053_), .A2(new_n4119_), .Z(po0987));
  INV_X1     g29928(.I(pi1162), .ZN(new_n33186_));
  NOR4_X1    g29929(.A1(new_n6957_), .A2(pi0832), .A3(new_n2918_), .A4(new_n33186_), .ZN(po0989));
  MUX2_X1    g29930(.I0(pi1091), .I1(new_n2553_), .S(new_n2925_), .Z(po0990));
  AND2_X2    g29931(.A1(new_n2925_), .A2(pi0946), .Z(po0991));
  XOR2_X1    g29932(.A1(new_n32157_), .A2(new_n33072_), .Z(po0992));
  NAND2_X1   g29933(.A1(pi0837), .A2(pi0955), .ZN(new_n33191_));
  OAI21_X1   g29934(.A1(pi0955), .A2(new_n30390_), .B(new_n33191_), .ZN(po0993));
  NAND2_X1   g29935(.A1(pi0838), .A2(pi0955), .ZN(new_n33193_));
  OAI21_X1   g29936(.A1(pi0955), .A2(new_n30502_), .B(new_n33193_), .ZN(po0994));
  NAND2_X1   g29937(.A1(pi0839), .A2(pi0955), .ZN(new_n33195_));
  OAI21_X1   g29938(.A1(pi0955), .A2(new_n30509_), .B(new_n33195_), .ZN(po0995));
  NAND2_X1   g29939(.A1(new_n2926_), .A2(pi0840), .ZN(new_n33197_));
  OAI21_X1   g29940(.A1(new_n6209_), .A2(new_n2926_), .B(new_n33197_), .ZN(po0996));
  NOR2_X1    g29941(.A1(new_n7318_), .A2(pi0033), .ZN(po0997));
  NAND2_X1   g29942(.A1(pi0842), .A2(pi0955), .ZN(new_n33200_));
  OAI21_X1   g29943(.A1(pi0955), .A2(new_n30600_), .B(new_n33200_), .ZN(po0998));
  NAND2_X1   g29944(.A1(pi0843), .A2(pi0955), .ZN(new_n33202_));
  OAI21_X1   g29945(.A1(pi0955), .A2(new_n30603_), .B(new_n33202_), .ZN(po0999));
  NAND2_X1   g29946(.A1(pi0844), .A2(pi0955), .ZN(new_n33204_));
  OAI21_X1   g29947(.A1(pi0955), .A2(new_n30606_), .B(new_n33204_), .ZN(po1000));
  NAND2_X1   g29948(.A1(pi0845), .A2(pi0955), .ZN(new_n33206_));
  OAI21_X1   g29949(.A1(pi0955), .A2(new_n30539_), .B(new_n33206_), .ZN(po1001));
  NAND2_X1   g29950(.A1(new_n29419_), .A2(pi0846), .ZN(new_n33208_));
  OAI21_X1   g29951(.A1(new_n29634_), .A2(new_n29419_), .B(new_n33208_), .ZN(po1002));
  NAND2_X1   g29952(.A1(pi0847), .A2(pi0955), .ZN(new_n33210_));
  OAI21_X1   g29953(.A1(pi0955), .A2(new_n30592_), .B(new_n33210_), .ZN(po1003));
  NAND2_X1   g29954(.A1(pi0848), .A2(pi0955), .ZN(new_n33212_));
  OAI21_X1   g29955(.A1(pi0955), .A2(new_n29011_), .B(new_n33212_), .ZN(po1004));
  NAND2_X1   g29956(.A1(new_n2926_), .A2(pi0849), .ZN(new_n33214_));
  OAI21_X1   g29957(.A1(new_n6156_), .A2(new_n2926_), .B(new_n33214_), .ZN(po1005));
  NAND2_X1   g29958(.A1(pi0850), .A2(pi0955), .ZN(new_n33216_));
  OAI21_X1   g29959(.A1(pi0955), .A2(new_n30387_), .B(new_n33216_), .ZN(po1006));
  NAND2_X1   g29960(.A1(pi0851), .A2(pi0955), .ZN(new_n33218_));
  OAI21_X1   g29961(.A1(pi0955), .A2(new_n30611_), .B(new_n33218_), .ZN(po1007));
  NAND2_X1   g29962(.A1(pi0852), .A2(pi0955), .ZN(new_n33220_));
  OAI21_X1   g29963(.A1(pi0955), .A2(new_n29391_), .B(new_n33220_), .ZN(po1008));
  NAND2_X1   g29964(.A1(pi0853), .A2(pi0955), .ZN(new_n33222_));
  OAI21_X1   g29965(.A1(pi0955), .A2(new_n30497_), .B(new_n33222_), .ZN(po1009));
  NAND2_X1   g29966(.A1(pi0854), .A2(pi0955), .ZN(new_n33224_));
  OAI21_X1   g29967(.A1(pi0955), .A2(new_n30521_), .B(new_n33224_), .ZN(po1010));
  NAND2_X1   g29968(.A1(pi0855), .A2(pi0955), .ZN(new_n33226_));
  OAI21_X1   g29969(.A1(pi0955), .A2(new_n29385_), .B(new_n33226_), .ZN(po1011));
  NAND2_X1   g29970(.A1(pi0856), .A2(pi0955), .ZN(new_n33228_));
  OAI21_X1   g29971(.A1(pi0955), .A2(new_n29404_), .B(new_n33228_), .ZN(po1012));
  NAND2_X1   g29972(.A1(pi0857), .A2(pi0955), .ZN(new_n33230_));
  OAI21_X1   g29973(.A1(pi0955), .A2(new_n30518_), .B(new_n33230_), .ZN(po1013));
  NAND2_X1   g29974(.A1(pi0858), .A2(pi0955), .ZN(new_n33232_));
  OAI21_X1   g29975(.A1(pi0955), .A2(new_n30595_), .B(new_n33232_), .ZN(po1014));
  NAND2_X1   g29976(.A1(pi0859), .A2(pi0955), .ZN(new_n33234_));
  OAI21_X1   g29977(.A1(pi0955), .A2(new_n29379_), .B(new_n33234_), .ZN(po1015));
  NAND2_X1   g29978(.A1(pi0860), .A2(pi0955), .ZN(new_n33236_));
  OAI21_X1   g29979(.A1(pi0955), .A2(new_n30619_), .B(new_n33236_), .ZN(po1016));
  MUX2_X1    g29980(.I0(pi0861), .I1(pi1141), .S(pi1093), .Z(new_n33238_));
  NAND2_X1   g29981(.A1(new_n33238_), .A2(new_n2523_), .ZN(new_n33239_));
  MUX2_X1    g29982(.I0(new_n3831_), .I1(new_n3839_), .S(pi0123), .Z(new_n33240_));
  OAI21_X1   g29983(.A1(new_n2523_), .A2(new_n33240_), .B(new_n33239_), .ZN(po1017));
  NAND2_X1   g29984(.A1(new_n29419_), .A2(pi0862), .ZN(new_n33242_));
  OAI21_X1   g29985(.A1(new_n4115_), .A2(new_n29419_), .B(new_n33242_), .ZN(po1018));
  NAND2_X1   g29986(.A1(new_n2926_), .A2(pi0863), .ZN(new_n33244_));
  OAI21_X1   g29987(.A1(new_n6088_), .A2(new_n2926_), .B(new_n33244_), .ZN(po1019));
  NAND2_X1   g29988(.A1(new_n2926_), .A2(pi0864), .ZN(new_n33246_));
  OAI21_X1   g29989(.A1(new_n6090_), .A2(new_n2926_), .B(new_n33246_), .ZN(po1020));
  NAND2_X1   g29990(.A1(pi0865), .A2(pi0955), .ZN(new_n33248_));
  OAI21_X1   g29991(.A1(pi0955), .A2(new_n29410_), .B(new_n33248_), .ZN(po1021));
  NAND2_X1   g29992(.A1(pi0866), .A2(pi0955), .ZN(new_n33250_));
  OAI21_X1   g29993(.A1(pi0955), .A2(new_n30402_), .B(new_n33250_), .ZN(po1022));
  NAND2_X1   g29994(.A1(pi0867), .A2(pi0955), .ZN(new_n33252_));
  OAI21_X1   g29995(.A1(pi0955), .A2(new_n30532_), .B(new_n33252_), .ZN(po1023));
  NAND2_X1   g29996(.A1(pi0868), .A2(pi0955), .ZN(new_n33254_));
  OAI21_X1   g29997(.A1(pi0955), .A2(new_n30529_), .B(new_n33254_), .ZN(po1024));
  MUX2_X1    g29998(.I0(pi0869), .I1(pi1140), .S(pi1093), .Z(new_n33256_));
  NAND2_X1   g29999(.A1(new_n33256_), .A2(new_n2523_), .ZN(new_n33257_));
  MUX2_X1    g30000(.I0(new_n3973_), .I1(new_n3981_), .S(pi0123), .Z(new_n33258_));
  OAI21_X1   g30001(.A1(new_n2523_), .A2(new_n33258_), .B(new_n33257_), .ZN(po1025));
  NAND2_X1   g30002(.A1(pi0870), .A2(pi0955), .ZN(new_n33260_));
  OAI21_X1   g30003(.A1(pi0955), .A2(new_n29397_), .B(new_n33260_), .ZN(po1026));
  NAND2_X1   g30004(.A1(pi0871), .A2(pi0955), .ZN(new_n33262_));
  OAI21_X1   g30005(.A1(pi0955), .A2(new_n30399_), .B(new_n33262_), .ZN(po1027));
  NAND2_X1   g30006(.A1(pi0872), .A2(pi0955), .ZN(new_n33264_));
  OAI21_X1   g30007(.A1(pi0955), .A2(new_n30393_), .B(new_n33264_), .ZN(po1028));
  NAND2_X1   g30008(.A1(pi0873), .A2(pi0955), .ZN(new_n33266_));
  OAI21_X1   g30009(.A1(pi0955), .A2(new_n30408_), .B(new_n33266_), .ZN(po1029));
  NAND2_X1   g30010(.A1(pi0874), .A2(pi0955), .ZN(new_n33268_));
  OAI21_X1   g30011(.A1(pi0955), .A2(new_n29374_), .B(new_n33268_), .ZN(po1030));
  OAI21_X1   g30012(.A1(new_n33109_), .A2(pi0875), .B(new_n2523_), .ZN(new_n33270_));
  AOI21_X1   g30013(.A1(new_n33109_), .A2(new_n4543_), .B(new_n33270_), .ZN(new_n33271_));
  NOR2_X1    g30014(.A1(new_n2924_), .A2(new_n4543_), .ZN(new_n33272_));
  NOR2_X1    g30015(.A1(new_n2924_), .A2(pi0875), .ZN(new_n33273_));
  NOR4_X1    g30016(.A1(new_n33271_), .A2(pi0228), .A3(new_n33272_), .A4(new_n33273_), .ZN(po1031));
  NAND2_X1   g30017(.A1(pi0876), .A2(pi0955), .ZN(new_n33275_));
  OAI21_X1   g30018(.A1(pi0955), .A2(new_n30405_), .B(new_n33275_), .ZN(po1032));
  MUX2_X1    g30019(.I0(pi0877), .I1(pi1138), .S(pi1093), .Z(new_n33277_));
  NAND2_X1   g30020(.A1(new_n33277_), .A2(new_n2523_), .ZN(new_n33278_));
  MUX2_X1    g30021(.I0(new_n4261_), .I1(new_n4269_), .S(pi0123), .Z(new_n33279_));
  OAI21_X1   g30022(.A1(new_n2523_), .A2(new_n33279_), .B(new_n33278_), .ZN(po1033));
  MUX2_X1    g30023(.I0(pi0878), .I1(pi1137), .S(pi1093), .Z(new_n33281_));
  NAND2_X1   g30024(.A1(new_n33281_), .A2(new_n2523_), .ZN(new_n33282_));
  MUX2_X1    g30025(.I0(new_n4402_), .I1(new_n4410_), .S(pi0123), .Z(new_n33283_));
  OAI21_X1   g30026(.A1(new_n2523_), .A2(new_n33283_), .B(new_n33282_), .ZN(po1034));
  MUX2_X1    g30027(.I0(pi0879), .I1(pi1135), .S(pi1093), .Z(new_n33285_));
  NAND2_X1   g30028(.A1(new_n33285_), .A2(new_n2523_), .ZN(new_n33286_));
  MUX2_X1    g30029(.I0(new_n4696_), .I1(new_n4702_), .S(pi0123), .Z(new_n33287_));
  OAI21_X1   g30030(.A1(new_n2523_), .A2(new_n33287_), .B(new_n33286_), .ZN(po1035));
  NAND2_X1   g30031(.A1(pi0880), .A2(pi0955), .ZN(new_n33289_));
  OAI21_X1   g30032(.A1(pi0955), .A2(new_n30616_), .B(new_n33289_), .ZN(po1036));
  NAND2_X1   g30033(.A1(pi0881), .A2(pi0955), .ZN(new_n33291_));
  OAI21_X1   g30034(.A1(pi0955), .A2(new_n30396_), .B(new_n33291_), .ZN(po1037));
  INV_X1     g30035(.I(pi0883), .ZN(po1163));
  NAND2_X1   g30036(.A1(new_n33110_), .A2(po1163), .ZN(new_n33294_));
  OAI21_X1   g30037(.A1(new_n32943_), .A2(new_n33110_), .B(new_n33294_), .ZN(po1039));
  INV_X1     g30038(.I(pi0884), .ZN(po1180));
  NAND2_X1   g30039(.A1(new_n33110_), .A2(po1180), .ZN(new_n33297_));
  OAI21_X1   g30040(.A1(new_n32142_), .A2(new_n33110_), .B(new_n33297_), .ZN(po1040));
  INV_X1     g30041(.I(pi0885), .ZN(po1172));
  NAND2_X1   g30042(.A1(new_n33110_), .A2(po1172), .ZN(new_n33300_));
  OAI21_X1   g30043(.A1(new_n32291_), .A2(new_n33110_), .B(new_n33300_), .ZN(po1041));
  INV_X1     g30044(.I(pi0886), .ZN(po1166));
  NAND2_X1   g30045(.A1(new_n33110_), .A2(po1166), .ZN(new_n33303_));
  OAI21_X1   g30046(.A1(new_n32878_), .A2(new_n33110_), .B(new_n33303_), .ZN(po1042));
  INV_X1     g30047(.I(pi0887), .ZN(po1179));
  NAND2_X1   g30048(.A1(new_n33110_), .A2(po1179), .ZN(new_n33306_));
  OAI21_X1   g30049(.A1(new_n33149_), .A2(new_n33110_), .B(new_n33306_), .ZN(po1043));
  INV_X1     g30050(.I(pi0888), .ZN(po1164));
  NAND2_X1   g30051(.A1(new_n33110_), .A2(po1164), .ZN(new_n33309_));
  OAI21_X1   g30052(.A1(new_n32797_), .A2(new_n33110_), .B(new_n33309_), .ZN(po1044));
  INV_X1     g30053(.I(pi0889), .ZN(po1170));
  NAND2_X1   g30054(.A1(new_n33110_), .A2(po1170), .ZN(new_n33312_));
  OAI21_X1   g30055(.A1(new_n32939_), .A2(new_n33110_), .B(new_n33312_), .ZN(po1045));
  INV_X1     g30056(.I(pi0890), .ZN(po1153));
  NAND2_X1   g30057(.A1(new_n33110_), .A2(po1153), .ZN(new_n33315_));
  OAI21_X1   g30058(.A1(new_n32121_), .A2(new_n33110_), .B(new_n33315_), .ZN(po1046));
  INV_X1     g30059(.I(pi0891), .ZN(po1160));
  NAND2_X1   g30060(.A1(new_n33110_), .A2(po1160), .ZN(new_n33318_));
  OAI21_X1   g30061(.A1(new_n32556_), .A2(new_n33110_), .B(new_n33318_), .ZN(po1047));
  INV_X1     g30062(.I(pi0892), .ZN(po1183));
  NAND2_X1   g30063(.A1(new_n33110_), .A2(po1183), .ZN(new_n33321_));
  OAI21_X1   g30064(.A1(new_n32925_), .A2(new_n33110_), .B(new_n33321_), .ZN(po1048));
  INV_X1     g30065(.I(pi0894), .ZN(po1150));
  NAND2_X1   g30066(.A1(new_n33110_), .A2(po1150), .ZN(new_n33324_));
  OAI21_X1   g30067(.A1(new_n32851_), .A2(new_n33110_), .B(new_n33324_), .ZN(po1050));
  INV_X1     g30068(.I(pi0895), .ZN(po1168));
  NAND2_X1   g30069(.A1(new_n33110_), .A2(po1168), .ZN(new_n33327_));
  OAI21_X1   g30070(.A1(new_n32073_), .A2(new_n33110_), .B(new_n33327_), .ZN(po1051));
  INV_X1     g30071(.I(pi0896), .ZN(po1156));
  NAND2_X1   g30072(.A1(new_n33110_), .A2(po1156), .ZN(new_n33330_));
  OAI21_X1   g30073(.A1(new_n32607_), .A2(new_n33110_), .B(new_n33330_), .ZN(po1052));
  INV_X1     g30074(.I(pi0898), .ZN(po1176));
  NAND2_X1   g30075(.A1(new_n33110_), .A2(po1176), .ZN(new_n33333_));
  OAI21_X1   g30076(.A1(new_n32539_), .A2(new_n33110_), .B(new_n33333_), .ZN(po1054));
  INV_X1     g30077(.I(pi0899), .ZN(po1174));
  NAND2_X1   g30078(.A1(new_n33110_), .A2(po1174), .ZN(new_n33336_));
  OAI21_X1   g30079(.A1(new_n32078_), .A2(new_n33110_), .B(new_n33336_), .ZN(po1055));
  INV_X1     g30080(.I(pi0900), .ZN(po1171));
  NAND2_X1   g30081(.A1(new_n33110_), .A2(po1171), .ZN(new_n33339_));
  OAI21_X1   g30082(.A1(new_n32949_), .A2(new_n33110_), .B(new_n33339_), .ZN(po1056));
  INV_X1     g30083(.I(pi0902), .ZN(po1161));
  NAND2_X1   g30084(.A1(new_n33110_), .A2(po1161), .ZN(new_n33342_));
  OAI21_X1   g30085(.A1(new_n32547_), .A2(new_n33110_), .B(new_n33342_), .ZN(po1058));
  INV_X1     g30086(.I(pi0903), .ZN(po1162));
  NAND2_X1   g30087(.A1(new_n33110_), .A2(po1162), .ZN(new_n33345_));
  OAI21_X1   g30088(.A1(new_n32863_), .A2(new_n33110_), .B(new_n33345_), .ZN(po1059));
  INV_X1     g30089(.I(pi0904), .ZN(po1173));
  NAND2_X1   g30090(.A1(new_n33110_), .A2(po1173), .ZN(new_n33348_));
  OAI21_X1   g30091(.A1(new_n32125_), .A2(new_n33110_), .B(new_n33348_), .ZN(po1060));
  INV_X1     g30092(.I(pi0905), .ZN(po1151));
  NAND2_X1   g30093(.A1(new_n33110_), .A2(po1151), .ZN(new_n33351_));
  OAI21_X1   g30094(.A1(new_n32149_), .A2(new_n33110_), .B(new_n33351_), .ZN(po1061));
  INV_X1     g30095(.I(pi0906), .ZN(po1155));
  NAND2_X1   g30096(.A1(new_n33110_), .A2(po1155), .ZN(new_n33354_));
  OAI21_X1   g30097(.A1(new_n32543_), .A2(new_n33110_), .B(new_n33354_), .ZN(po1062));
  INV_X1     g30098(.I(pi0782), .ZN(new_n33356_));
  INV_X1     g30099(.I(pi0598), .ZN(new_n33357_));
  INV_X1     g30100(.I(pi0624), .ZN(new_n33358_));
  MUX2_X1    g30101(.I0(new_n33358_), .I1(new_n33357_), .S(pi0979), .Z(new_n33359_));
  NOR2_X1    g30102(.A1(new_n33359_), .A2(new_n33356_), .ZN(new_n33360_));
  NOR2_X1    g30103(.A1(new_n5119_), .A2(pi0615), .ZN(new_n33361_));
  INV_X1     g30104(.I(pi0604), .ZN(new_n33362_));
  OAI21_X1   g30105(.A1(new_n33362_), .A2(pi0979), .B(pi0782), .ZN(new_n33363_));
  OAI22_X1   g30106(.A1(new_n33363_), .A2(new_n33361_), .B1(pi0782), .B2(pi0907), .ZN(new_n33364_));
  NOR2_X1    g30107(.A1(new_n33360_), .A2(new_n33364_), .ZN(po1063));
  INV_X1     g30108(.I(pi0908), .ZN(po1159));
  NAND2_X1   g30109(.A1(new_n33110_), .A2(po1159), .ZN(new_n33367_));
  OAI21_X1   g30110(.A1(new_n32859_), .A2(new_n33110_), .B(new_n33367_), .ZN(po1064));
  INV_X1     g30111(.I(pi0909), .ZN(po1157));
  NAND2_X1   g30112(.A1(new_n33110_), .A2(po1157), .ZN(new_n33370_));
  OAI21_X1   g30113(.A1(new_n32033_), .A2(new_n33110_), .B(new_n33370_), .ZN(po1065));
  INV_X1     g30114(.I(pi0910), .ZN(po1181));
  NAND2_X1   g30115(.A1(new_n33110_), .A2(po1181), .ZN(new_n33373_));
  OAI21_X1   g30116(.A1(new_n32568_), .A2(new_n33110_), .B(new_n33373_), .ZN(po1066));
  INV_X1     g30117(.I(pi0911), .ZN(po1158));
  NAND2_X1   g30118(.A1(new_n33110_), .A2(po1158), .ZN(new_n33376_));
  OAI21_X1   g30119(.A1(new_n32138_), .A2(new_n33110_), .B(new_n33376_), .ZN(po1067));
  INV_X1     g30120(.I(pi0912), .ZN(po1167));
  NAND2_X1   g30121(.A1(new_n33110_), .A2(po1167), .ZN(new_n33379_));
  OAI21_X1   g30122(.A1(new_n32113_), .A2(new_n33110_), .B(new_n33379_), .ZN(po1068));
  INV_X1     g30123(.I(pi0913), .ZN(po1149));
  NAND2_X1   g30124(.A1(new_n33110_), .A2(po1149), .ZN(new_n33382_));
  OAI21_X1   g30125(.A1(new_n32901_), .A2(new_n33110_), .B(new_n33382_), .ZN(po1069));
  NAND2_X1   g30126(.A1(pi0266), .A2(pi0992), .ZN(new_n33384_));
  XOR2_X1    g30127(.A1(new_n33384_), .A2(pi0280), .Z(po1070));
  INV_X1     g30128(.I(pi0915), .ZN(po1146));
  NAND2_X1   g30129(.A1(new_n33110_), .A2(po1146), .ZN(new_n33387_));
  OAI21_X1   g30130(.A1(new_n32869_), .A2(new_n33110_), .B(new_n33387_), .ZN(po1071));
  INV_X1     g30131(.I(pi0916), .ZN(po1169));
  NAND2_X1   g30132(.A1(new_n33110_), .A2(po1169), .ZN(new_n33390_));
  OAI21_X1   g30133(.A1(new_n32564_), .A2(new_n33110_), .B(new_n33390_), .ZN(po1072));
  INV_X1     g30134(.I(pi0917), .ZN(po1177));
  NAND2_X1   g30135(.A1(new_n33110_), .A2(po1177), .ZN(new_n33393_));
  OAI21_X1   g30136(.A1(new_n32086_), .A2(new_n33110_), .B(new_n33393_), .ZN(po1073));
  INV_X1     g30137(.I(pi0918), .ZN(po1175));
  NAND2_X1   g30138(.A1(new_n33110_), .A2(po1175), .ZN(new_n33396_));
  OAI21_X1   g30139(.A1(new_n31998_), .A2(new_n33110_), .B(new_n33396_), .ZN(po1074));
  INV_X1     g30140(.I(pi0919), .ZN(po1165));
  NAND2_X1   g30141(.A1(new_n33110_), .A2(po1165), .ZN(new_n33399_));
  OAI21_X1   g30142(.A1(new_n32988_), .A2(new_n33110_), .B(new_n33399_), .ZN(po1075));
  NAND2_X1   g30143(.A1(new_n2924_), .A2(pi0920), .ZN(new_n33401_));
  OAI21_X1   g30144(.A1(new_n2924_), .A2(new_n4115_), .B(new_n33401_), .ZN(po1076));
  NAND2_X1   g30145(.A1(pi1093), .A2(pi1140), .ZN(new_n33403_));
  OAI21_X1   g30146(.A1(new_n3974_), .A2(pi1093), .B(new_n33403_), .ZN(po1077));
  NAND2_X1   g30147(.A1(pi1093), .A2(pi1152), .ZN(new_n33405_));
  OAI21_X1   g30148(.A1(new_n30910_), .A2(pi1093), .B(new_n33405_), .ZN(po1078));
  NAND2_X1   g30149(.A1(new_n2924_), .A2(pi0923), .ZN(new_n33407_));
  OAI21_X1   g30150(.A1(new_n2924_), .A2(new_n11950_), .B(new_n33407_), .ZN(po1079));
  NOR4_X1    g30151(.A1(new_n30423_), .A2(new_n30478_), .A3(pi0300), .A4(pi0312), .ZN(po1080));
  NAND2_X1   g30152(.A1(new_n2924_), .A2(pi0925), .ZN(new_n33410_));
  OAI21_X1   g30153(.A1(new_n2924_), .A2(new_n11912_), .B(new_n33410_), .ZN(po1081));
  NAND2_X1   g30154(.A1(new_n2924_), .A2(pi0926), .ZN(new_n33412_));
  OAI21_X1   g30155(.A1(new_n2924_), .A2(new_n12049_), .B(new_n33412_), .ZN(po1082));
  NAND2_X1   g30156(.A1(pi1093), .A2(pi1145), .ZN(new_n33414_));
  OAI21_X1   g30157(.A1(new_n3412_), .A2(pi1093), .B(new_n33414_), .ZN(po1083));
  INV_X1     g30158(.I(new_n33272_), .ZN(new_n33416_));
  OAI21_X1   g30159(.A1(new_n4568_), .A2(pi1093), .B(new_n33416_), .ZN(po1084));
  NAND2_X1   g30160(.A1(pi1093), .A2(pi1144), .ZN(new_n33418_));
  OAI21_X1   g30161(.A1(new_n2551_), .A2(pi1093), .B(new_n33418_), .ZN(po1085));
  NAND2_X1   g30162(.A1(new_n2924_), .A2(pi0930), .ZN(new_n33420_));
  OAI21_X1   g30163(.A1(new_n2924_), .A2(new_n29634_), .B(new_n33420_), .ZN(po1086));
  NAND2_X1   g30164(.A1(pi1093), .A2(pi1150), .ZN(new_n33422_));
  OAI21_X1   g30165(.A1(new_n30917_), .A2(pi1093), .B(new_n33422_), .ZN(po1087));
  NAND2_X1   g30166(.A1(pi1093), .A2(pi1142), .ZN(new_n33424_));
  OAI21_X1   g30167(.A1(new_n3701_), .A2(pi1093), .B(new_n33424_), .ZN(po1088));
  NAND2_X1   g30168(.A1(pi1093), .A2(pi1137), .ZN(new_n33426_));
  OAI21_X1   g30169(.A1(new_n4403_), .A2(pi1093), .B(new_n33426_), .ZN(po1089));
  NAND2_X1   g30170(.A1(new_n2924_), .A2(pi0934), .ZN(new_n33428_));
  OAI21_X1   g30171(.A1(new_n2924_), .A2(new_n27494_), .B(new_n33428_), .ZN(po1090));
  NAND2_X1   g30172(.A1(pi1093), .A2(pi1141), .ZN(new_n33430_));
  OAI21_X1   g30173(.A1(new_n3832_), .A2(pi1093), .B(new_n33430_), .ZN(po1091));
  NAND2_X1   g30174(.A1(pi1093), .A2(pi1149), .ZN(new_n33432_));
  OAI21_X1   g30175(.A1(new_n30924_), .A2(pi1093), .B(new_n33432_), .ZN(po1092));
  NAND2_X1   g30176(.A1(pi1093), .A2(pi1148), .ZN(new_n33434_));
  OAI21_X1   g30177(.A1(new_n30440_), .A2(pi1093), .B(new_n33434_), .ZN(po1093));
  NAND2_X1   g30178(.A1(pi1093), .A2(pi1135), .ZN(new_n33436_));
  OAI21_X1   g30179(.A1(new_n4732_), .A2(pi1093), .B(new_n33436_), .ZN(po1094));
  NAND2_X1   g30180(.A1(pi1093), .A2(pi1146), .ZN(new_n33438_));
  OAI21_X1   g30181(.A1(new_n3261_), .A2(pi1093), .B(new_n33438_), .ZN(po1095));
  NAND2_X1   g30182(.A1(pi1093), .A2(pi1138), .ZN(new_n33440_));
  OAI21_X1   g30183(.A1(new_n4262_), .A2(pi1093), .B(new_n33440_), .ZN(po1096));
  NAND2_X1   g30184(.A1(new_n2924_), .A2(pi0941), .ZN(new_n33442_));
  OAI21_X1   g30185(.A1(new_n2924_), .A2(new_n11893_), .B(new_n33442_), .ZN(po1097));
  NAND2_X1   g30186(.A1(new_n2924_), .A2(pi0942), .ZN(new_n33444_));
  OAI21_X1   g30187(.A1(new_n2924_), .A2(new_n12026_), .B(new_n33444_), .ZN(po1098));
  NAND2_X1   g30188(.A1(pi1093), .A2(pi1151), .ZN(new_n33446_));
  OAI21_X1   g30189(.A1(new_n30870_), .A2(pi1093), .B(new_n33446_), .ZN(po1099));
  NAND2_X1   g30190(.A1(pi1093), .A2(pi1143), .ZN(new_n33448_));
  OAI21_X1   g30191(.A1(new_n3549_), .A2(pi1093), .B(new_n33448_), .ZN(po1100));
  NOR2_X1    g30192(.A1(new_n2926_), .A2(new_n26307_), .ZN(po1102));
  INV_X1     g30193(.I(new_n33360_), .ZN(new_n33451_));
  OAI21_X1   g30194(.A1(pi0782), .A2(new_n5473_), .B(new_n33451_), .ZN(po1103));
  XOR2_X1    g30195(.A1(pi0266), .A2(pi0992), .Z(po1104));
  NAND2_X1   g30196(.A1(pi0949), .A2(pi0954), .ZN(new_n33454_));
  OAI21_X1   g30197(.A1(pi0313), .A2(pi0954), .B(new_n33454_), .ZN(po1105));
  NOR3_X1    g30198(.A1(new_n6003_), .A2(new_n2927_), .A3(new_n2923_), .ZN(po1107));
  OAI21_X1   g30199(.A1(new_n2919_), .A2(new_n2923_), .B(new_n6958_), .ZN(po1112));
  NOR2_X1    g30200(.A1(new_n5645_), .A2(pi0782), .ZN(po1115));
  NOR2_X1    g30201(.A1(new_n5600_), .A2(pi0230), .ZN(po1116));
  NOR2_X1    g30202(.A1(new_n5697_), .A2(pi0782), .ZN(po1118));
  NOR2_X1    g30203(.A1(new_n5514_), .A2(pi0230), .ZN(po1122));
  NOR2_X1    g30204(.A1(new_n5704_), .A2(pi0230), .ZN(po1124));
  NOR2_X1    g30205(.A1(new_n5504_), .A2(pi0782), .ZN(po1125));
  NOR2_X1    g30206(.A1(new_n5756_), .A2(pi0230), .ZN(po1126));
  NOR2_X1    g30207(.A1(new_n5593_), .A2(pi0782), .ZN(po1127));
  NOR2_X1    g30208(.A1(new_n5807_), .A2(pi0230), .ZN(po1128));
  NOR2_X1    g30209(.A1(new_n5749_), .A2(pi0782), .ZN(po1129));
  NOR2_X1    g30210(.A1(new_n5652_), .A2(pi0230), .ZN(po1131));
  NOR2_X1    g30211(.A1(new_n5803_), .A2(pi0782), .ZN(po1132));
  NAND2_X1   g30212(.A1(new_n33357_), .A2(pi0615), .ZN(po1133));
  NOR2_X1    g30213(.A1(new_n5366_), .A2(new_n2923_), .ZN(po1135));
  NAND2_X1   g30214(.A1(new_n33362_), .A2(new_n33358_), .ZN(po1137));
  assign     po0166 = 1'b1;
  assign     po0436 = 1'b0;
  assign     po0439 = 1'b0;
  assign     po0441 = 1'b0;
  assign     po0622 = 1'b0;
  assign     po0626 = 1'b0;
  assign     po0627 = 1'b0;
  assign     po0628 = 1'b0;
  assign     po0629 = 1'b0;
  assign     po0842 = 1'b0;
  assign     po0846 = 1'b0;
  assign     po0864 = 1'b0;
  assign     po0868 = 1'b0;
  assign     po0870 = 1'b0;
  assign     po0871 = 1'b0;
  assign     po0877 = 1'b0;
  BUF_X16    g30215(.I(pi0668), .Z(po0000));
  BUF_X16    g30216(.I(pi0672), .Z(po0001));
  BUF_X16    g30217(.I(pi0664), .Z(po0002));
  BUF_X16    g30218(.I(pi0667), .Z(po0003));
  BUF_X16    g30219(.I(pi0676), .Z(po0004));
  BUF_X16    g30220(.I(pi0673), .Z(po0005));
  BUF_X16    g30221(.I(pi0675), .Z(po0006));
  BUF_X16    g30222(.I(pi0666), .Z(po0007));
  BUF_X16    g30223(.I(pi0679), .Z(po0008));
  BUF_X16    g30224(.I(pi0674), .Z(po0009));
  BUF_X16    g30225(.I(pi0663), .Z(po0010));
  BUF_X16    g30226(.I(pi0670), .Z(po0011));
  BUF_X16    g30227(.I(pi0677), .Z(po0012));
  BUF_X16    g30228(.I(pi0682), .Z(po0013));
  BUF_X16    g30229(.I(pi0671), .Z(po0014));
  BUF_X16    g30230(.I(pi0678), .Z(po0015));
  BUF_X16    g30231(.I(pi0718), .Z(po0016));
  BUF_X16    g30232(.I(pi0707), .Z(po0017));
  BUF_X16    g30233(.I(pi0708), .Z(po0018));
  BUF_X16    g30234(.I(pi0713), .Z(po0019));
  BUF_X16    g30235(.I(pi0711), .Z(po0020));
  BUF_X16    g30236(.I(pi0716), .Z(po0021));
  BUF_X16    g30237(.I(pi0733), .Z(po0022));
  BUF_X16    g30238(.I(pi0712), .Z(po0023));
  BUF_X16    g30239(.I(pi0689), .Z(po0024));
  BUF_X16    g30240(.I(pi0717), .Z(po0025));
  BUF_X16    g30241(.I(pi0692), .Z(po0026));
  BUF_X16    g30242(.I(pi0719), .Z(po0027));
  BUF_X16    g30243(.I(pi0722), .Z(po0028));
  BUF_X16    g30244(.I(pi0714), .Z(po0029));
  BUF_X16    g30245(.I(pi0720), .Z(po0030));
  BUF_X16    g30246(.I(pi0685), .Z(po0031));
  BUF_X16    g30247(.I(pi0837), .Z(po0032));
  BUF_X16    g30248(.I(pi0850), .Z(po0033));
  BUF_X16    g30249(.I(pi0872), .Z(po0034));
  BUF_X16    g30250(.I(pi0871), .Z(po0035));
  BUF_X16    g30251(.I(pi0881), .Z(po0036));
  BUF_X16    g30252(.I(pi0866), .Z(po0037));
  BUF_X16    g30253(.I(pi0876), .Z(po0038));
  BUF_X16    g30254(.I(pi0873), .Z(po0039));
  BUF_X16    g30255(.I(pi0874), .Z(po0040));
  BUF_X16    g30256(.I(pi0859), .Z(po0041));
  BUF_X16    g30257(.I(pi0855), .Z(po0042));
  BUF_X16    g30258(.I(pi0852), .Z(po0043));
  BUF_X16    g30259(.I(pi0870), .Z(po0044));
  BUF_X16    g30260(.I(pi0848), .Z(po0045));
  BUF_X16    g30261(.I(pi0865), .Z(po0046));
  BUF_X16    g30262(.I(pi0856), .Z(po0047));
  BUF_X16    g30263(.I(pi0853), .Z(po0048));
  BUF_X16    g30264(.I(pi0847), .Z(po0049));
  BUF_X16    g30265(.I(pi0857), .Z(po0050));
  BUF_X16    g30266(.I(pi0854), .Z(po0051));
  BUF_X16    g30267(.I(pi0858), .Z(po0052));
  BUF_X16    g30268(.I(pi0845), .Z(po0053));
  BUF_X16    g30269(.I(pi0838), .Z(po0054));
  BUF_X16    g30270(.I(pi0842), .Z(po0055));
  BUF_X16    g30271(.I(pi0843), .Z(po0056));
  BUF_X16    g30272(.I(pi0839), .Z(po0057));
  BUF_X16    g30273(.I(pi0844), .Z(po0058));
  BUF_X16    g30274(.I(pi0868), .Z(po0059));
  BUF_X16    g30275(.I(pi0851), .Z(po0060));
  BUF_X16    g30276(.I(pi0867), .Z(po0061));
  BUF_X16    g30277(.I(pi0880), .Z(po0062));
  BUF_X16    g30278(.I(pi0860), .Z(po0063));
  BUF_X16    g30279(.I(pi1030), .Z(po0064));
  BUF_X16    g30280(.I(pi1034), .Z(po0065));
  BUF_X16    g30281(.I(pi1015), .Z(po0066));
  BUF_X16    g30282(.I(pi1020), .Z(po0067));
  BUF_X16    g30283(.I(pi1025), .Z(po0068));
  BUF_X16    g30284(.I(pi1005), .Z(po0069));
  BUF_X16    g30285(.I(pi0996), .Z(po0070));
  BUF_X16    g30286(.I(pi1012), .Z(po0071));
  BUF_X16    g30287(.I(pi0993), .Z(po0072));
  BUF_X16    g30288(.I(pi1016), .Z(po0073));
  BUF_X16    g30289(.I(pi1021), .Z(po0074));
  BUF_X16    g30290(.I(pi1010), .Z(po0075));
  BUF_X16    g30291(.I(pi1027), .Z(po0076));
  BUF_X16    g30292(.I(pi1018), .Z(po0077));
  BUF_X16    g30293(.I(pi1017), .Z(po0078));
  BUF_X16    g30294(.I(pi1024), .Z(po0079));
  BUF_X16    g30295(.I(pi1009), .Z(po0080));
  BUF_X16    g30296(.I(pi1032), .Z(po0081));
  BUF_X16    g30297(.I(pi1003), .Z(po0082));
  BUF_X16    g30298(.I(pi0997), .Z(po0083));
  BUF_X16    g30299(.I(pi1013), .Z(po0084));
  BUF_X16    g30300(.I(pi1011), .Z(po0085));
  BUF_X16    g30301(.I(pi1008), .Z(po0086));
  BUF_X16    g30302(.I(pi1019), .Z(po0087));
  BUF_X16    g30303(.I(pi1031), .Z(po0088));
  BUF_X16    g30304(.I(pi1022), .Z(po0089));
  BUF_X16    g30305(.I(pi1000), .Z(po0090));
  BUF_X16    g30306(.I(pi1023), .Z(po0091));
  BUF_X16    g30307(.I(pi1002), .Z(po0092));
  BUF_X16    g30308(.I(pi1026), .Z(po0093));
  BUF_X16    g30309(.I(pi1006), .Z(po0094));
  BUF_X16    g30310(.I(pi0998), .Z(po0095));
  BUF_X16    g30311(.I(pi0031), .Z(po0096));
  BUF_X16    g30312(.I(pi0080), .Z(po0097));
  BUF_X16    g30313(.I(pi0893), .Z(po0098));
  BUF_X16    g30314(.I(pi0467), .Z(po0099));
  BUF_X16    g30315(.I(pi0078), .Z(po0100));
  BUF_X16    g30316(.I(pi0112), .Z(po0101));
  BUF_X16    g30317(.I(pi0013), .Z(po0102));
  BUF_X16    g30318(.I(pi0025), .Z(po0103));
  BUF_X16    g30319(.I(pi0226), .Z(po0104));
  BUF_X16    g30320(.I(pi0127), .Z(po0105));
  BUF_X16    g30321(.I(pi0822), .Z(po0106));
  BUF_X16    g30322(.I(pi0808), .Z(po0107));
  BUF_X16    g30323(.I(pi0227), .Z(po0108));
  BUF_X16    g30324(.I(pi0477), .Z(po0109));
  BUF_X16    g30325(.I(pi0834), .Z(po0110));
  BUF_X16    g30326(.I(pi0229), .Z(po0111));
  BUF_X16    g30327(.I(pi0012), .Z(po0112));
  BUF_X16    g30328(.I(pi0011), .Z(po0113));
  BUF_X16    g30329(.I(pi0010), .Z(po0114));
  BUF_X16    g30330(.I(pi0009), .Z(po0115));
  BUF_X16    g30331(.I(pi0008), .Z(po0116));
  BUF_X16    g30332(.I(pi0007), .Z(po0117));
  BUF_X16    g30333(.I(pi0006), .Z(po0118));
  BUF_X16    g30334(.I(pi0005), .Z(po0119));
  BUF_X16    g30335(.I(pi0004), .Z(po0120));
  BUF_X16    g30336(.I(pi0003), .Z(po0121));
  BUF_X16    g30337(.I(pi0000), .Z(po0122));
  BUF_X16    g30338(.I(pi0002), .Z(po0123));
  BUF_X16    g30339(.I(pi0001), .Z(po0124));
  BUF_X16    g30340(.I(pi0310), .Z(po0125));
  BUF_X16    g30341(.I(pi0302), .Z(po0126));
  BUF_X16    g30342(.I(pi0475), .Z(po0127));
  BUF_X16    g30343(.I(pi0474), .Z(po0128));
  BUF_X16    g30344(.I(pi0466), .Z(po0129));
  BUF_X16    g30345(.I(pi0473), .Z(po0130));
  BUF_X16    g30346(.I(pi0471), .Z(po0131));
  BUF_X16    g30347(.I(pi0472), .Z(po0132));
  BUF_X16    g30348(.I(pi0470), .Z(po0133));
  BUF_X16    g30349(.I(pi0469), .Z(po0134));
  BUF_X16    g30350(.I(pi0465), .Z(po0135));
  BUF_X16    g30351(.I(pi1028), .Z(po0136));
  BUF_X16    g30352(.I(pi1033), .Z(po0137));
  BUF_X16    g30353(.I(pi0995), .Z(po0138));
  BUF_X16    g30354(.I(pi0994), .Z(po0139));
  BUF_X16    g30355(.I(pi0028), .Z(po0140));
  BUF_X16    g30356(.I(pi0027), .Z(po0141));
  BUF_X16    g30357(.I(pi0026), .Z(po0142));
  BUF_X16    g30358(.I(pi0029), .Z(po0143));
  BUF_X16    g30359(.I(pi0015), .Z(po0144));
  BUF_X16    g30360(.I(pi0014), .Z(po0145));
  BUF_X16    g30361(.I(pi0021), .Z(po0146));
  BUF_X16    g30362(.I(pi0020), .Z(po0147));
  BUF_X16    g30363(.I(pi0019), .Z(po0148));
  BUF_X16    g30364(.I(pi0018), .Z(po0149));
  BUF_X16    g30365(.I(pi0017), .Z(po0150));
  BUF_X16    g30366(.I(pi0016), .Z(po0151));
  BUF_X16    g30367(.I(pi1096), .Z(po0152));
  BUF_X16    g30368(.I(pi0228), .Z(po0168));
  BUF_X16    g30369(.I(pi0022), .Z(po0169));
  BUF_X16    g30370(.I(pi1089), .Z(po0179));
  BUF_X16    g30371(.I(pi0023), .Z(po0180));
  OAI22_X1   g30372(.A1(new_n5202_), .A2(new_n5204_), .B1(new_n5055_), .B2(new_n5209_), .ZN(po0181));
  BUF_X16    g30373(.I(pi0037), .Z(po0188));
  BUF_X16    g30374(.I(pi0117), .Z(po0263));
  BUF_X16    g30375(.I(pi0131), .Z(po0285));
  BUF_X16    g30376(.I(pi0232), .Z(po0386));
  BUF_X16    g30377(.I(pi0236), .Z(po0388));
  BUF_X16    g30378(.I(pi0583), .Z(po0636));
  BUF_X16    g30379(.I(pi0067), .Z(po1053));
  BUF_X16    g30380(.I(pi1134), .Z(po1108));
  BUF_X16    g30381(.I(pi0964), .Z(po1109));
  BUF_X16    g30382(.I(pi0965), .Z(po1111));
  BUF_X16    g30383(.I(pi0991), .Z(po1113));
  BUF_X16    g30384(.I(pi0985), .Z(po1114));
  BUF_X16    g30385(.I(pi1014), .Z(po1117));
  BUF_X16    g30386(.I(pi1029), .Z(po1119));
  BUF_X16    g30387(.I(pi1004), .Z(po1120));
  BUF_X16    g30388(.I(pi1007), .Z(po1121));
  BUF_X16    g30389(.I(pi1135), .Z(po1123));
  BUF_X16    g30390(.I(pi1064), .Z(po1134));
  BUF_X16    g30391(.I(pi0299), .Z(po1136));
  BUF_X16    g30392(.I(pi1075), .Z(po1138));
  BUF_X16    g30393(.I(pi1052), .Z(po1139));
  BUF_X16    g30394(.I(pi0771), .Z(po1140));
  BUF_X16    g30395(.I(pi0765), .Z(po1141));
  BUF_X16    g30396(.I(pi0605), .Z(po1142));
  BUF_X16    g30397(.I(pi0601), .Z(po1143));
  BUF_X16    g30398(.I(pi0278), .Z(po1144));
  BUF_X16    g30399(.I(pi0279), .Z(po1145));
  BUF_X16    g30400(.I(pi1095), .Z(po1152));
  BUF_X16    g30401(.I(pi1094), .Z(po1154));
  BUF_X16    g30402(.I(pi1187), .Z(po1184));
  BUF_X16    g30403(.I(pi1172), .Z(po1185));
  BUF_X16    g30404(.I(pi1170), .Z(po1186));
  BUF_X16    g30405(.I(pi1138), .Z(po1187));
  BUF_X16    g30406(.I(pi1177), .Z(po1188));
  BUF_X16    g30407(.I(pi1178), .Z(po1189));
  BUF_X16    g30408(.I(pi0863), .Z(po1190));
  BUF_X16    g30409(.I(pi1203), .Z(po1191));
  BUF_X16    g30410(.I(pi1185), .Z(po1192));
  BUF_X16    g30411(.I(pi1171), .Z(po1193));
  BUF_X16    g30412(.I(pi1192), .Z(po1194));
  BUF_X16    g30413(.I(pi1137), .Z(po1195));
  BUF_X16    g30414(.I(pi1186), .Z(po1196));
  BUF_X16    g30415(.I(pi1165), .Z(po1197));
  BUF_X16    g30416(.I(pi1164), .Z(po1198));
  BUF_X16    g30417(.I(pi1098), .Z(po1199));
  BUF_X16    g30418(.I(pi1183), .Z(po1200));
  BUF_X16    g30419(.I(pi0230), .Z(po1201));
  BUF_X16    g30420(.I(pi1169), .Z(po1202));
  BUF_X16    g30421(.I(pi1136), .Z(po1203));
  BUF_X16    g30422(.I(pi1181), .Z(po1204));
  BUF_X16    g30423(.I(pi0849), .Z(po1205));
  BUF_X16    g30424(.I(pi1193), .Z(po1206));
  BUF_X16    g30425(.I(pi1182), .Z(po1207));
  BUF_X16    g30426(.I(pi1168), .Z(po1208));
  BUF_X16    g30427(.I(pi1175), .Z(po1209));
  BUF_X16    g30428(.I(pi1191), .Z(po1210));
  BUF_X16    g30429(.I(pi1099), .Z(po1211));
  BUF_X16    g30430(.I(pi1174), .Z(po1212));
  BUF_X16    g30431(.I(pi1179), .Z(po1213));
  BUF_X16    g30432(.I(pi1202), .Z(po1214));
  BUF_X16    g30433(.I(pi1176), .Z(po1215));
  BUF_X16    g30434(.I(pi1173), .Z(po1216));
  BUF_X16    g30435(.I(pi1201), .Z(po1217));
  BUF_X16    g30436(.I(pi1167), .Z(po1218));
  BUF_X16    g30437(.I(pi0840), .Z(po1219));
  BUF_X16    g30438(.I(pi1189), .Z(po1220));
  BUF_X16    g30439(.I(pi1195), .Z(po1221));
  BUF_X16    g30440(.I(pi0864), .Z(po1222));
  BUF_X16    g30441(.I(pi1190), .Z(po1223));
  BUF_X16    g30442(.I(pi1188), .Z(po1224));
  BUF_X16    g30443(.I(pi1180), .Z(po1225));
  BUF_X16    g30444(.I(pi1194), .Z(po1226));
  BUF_X16    g30445(.I(pi1097), .Z(po1227));
  BUF_X16    g30446(.I(pi1166), .Z(po1228));
  BUF_X16    g30447(.I(pi1200), .Z(po1229));
  BUF_X16    g30448(.I(pi1184), .Z(po1230));
endmodule


