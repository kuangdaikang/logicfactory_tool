// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:26 2022

module soar  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43,
    v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57,
    v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71,
    v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82,
    \v83.0 , \v83.1 , \v83.2 , \v83.3 , \v83.4 , \v83.5 , \v83.6 , \v83.7 ,
    \v83.8 , \v83.9 , \v83.10 , \v83.11 , \v83.12 , \v83.13 , \v83.14 ,
    \v83.15 , \v83.16 , \v83.17 , \v83.18 , \v83.19 , \v83.20 , \v83.21 ,
    \v83.22 , \v83.23 , \v83.24 , \v83.25 , \v83.26 , \v83.27 , \v83.28 ,
    \v83.29 , \v83.30 , \v83.31 , \v83.32 , \v83.33 , \v83.34 , \v83.35 ,
    \v83.36 , \v83.37 , \v83.38 , \v83.39 , \v83.40 , \v83.41 , \v83.42 ,
    \v83.43 , \v83.44 , \v83.45 , \v83.46 , \v83.47 , \v83.48 , \v83.49 ,
    \v83.50 , \v83.51 , \v83.52 , \v83.53 , \v83.54 , \v83.55 , \v83.56 ,
    \v83.57 , \v83.58 , \v83.59 , \v83.60 , \v83.61 , \v83.62 , \v83.63 ,
    \v83.64 , \v83.65 , \v83.66 , \v83.67 , \v83.68 , \v83.69 , \v83.70 ,
    \v83.71 , \v83.72 , \v83.73 , \v83.74 , \v83.75 , \v83.76 , \v83.77 ,
    \v83.78 , \v83.79 , \v83.80 , \v83.81 , \v83.82 , \v83.83 , \v83.84 ,
    \v83.85 , \v83.86 , \v83.87 , \v83.88 , \v83.89 , \v83.90 , \v83.91 ,
    \v83.92 , \v83.93   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42,
    v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56,
    v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70,
    v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82;
  output \v83.0 , \v83.1 , \v83.2 , \v83.3 , \v83.4 , \v83.5 , \v83.6 ,
    \v83.7 , \v83.8 , \v83.9 , \v83.10 , \v83.11 , \v83.12 , \v83.13 ,
    \v83.14 , \v83.15 , \v83.16 , \v83.17 , \v83.18 , \v83.19 , \v83.20 ,
    \v83.21 , \v83.22 , \v83.23 , \v83.24 , \v83.25 , \v83.26 , \v83.27 ,
    \v83.28 , \v83.29 , \v83.30 , \v83.31 , \v83.32 , \v83.33 , \v83.34 ,
    \v83.35 , \v83.36 , \v83.37 , \v83.38 , \v83.39 , \v83.40 , \v83.41 ,
    \v83.42 , \v83.43 , \v83.44 , \v83.45 , \v83.46 , \v83.47 , \v83.48 ,
    \v83.49 , \v83.50 , \v83.51 , \v83.52 , \v83.53 , \v83.54 , \v83.55 ,
    \v83.56 , \v83.57 , \v83.58 , \v83.59 , \v83.60 , \v83.61 , \v83.62 ,
    \v83.63 , \v83.64 , \v83.65 , \v83.66 , \v83.67 , \v83.68 , \v83.69 ,
    \v83.70 , \v83.71 , \v83.72 , \v83.73 , \v83.74 , \v83.75 , \v83.76 ,
    \v83.77 , \v83.78 , \v83.79 , \v83.80 , \v83.81 , \v83.82 , \v83.83 ,
    \v83.84 , \v83.85 , \v83.86 , \v83.87 , \v83.88 , \v83.89 , \v83.90 ,
    \v83.91 , \v83.92 , \v83.93 ;
  wire new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n201_, new_n202_, new_n203_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n267_, new_n268_, new_n270_, new_n271_,
    new_n272_, new_n274_, new_n275_, new_n276_, new_n277_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n339_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n358_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n376_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n513_, new_n514_, new_n515_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n553_, new_n554_, new_n555_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n564_, new_n566_, new_n567_,
    new_n569_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n579_, new_n581_, new_n582_, new_n584_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n613_,
    new_n614_, new_n615_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n708_, new_n711_, new_n712_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n750_, new_n752_, new_n754_, new_n755_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n889_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_;
  assign new_n178_ = ~v7 & v8;
  assign new_n179_ = v6 & ~new_n178_;
  assign new_n180_ = v9 & ~new_n179_;
  assign new_n181_ = ~v11 & ~new_n180_;
  assign new_n182_ = ~v6 & ~v7;
  assign new_n183_ = ~v8 & v11;
  assign new_n184_ = new_n182_ & new_n183_;
  assign new_n185_ = v12 & ~new_n184_;
  assign new_n186_ = v10 & new_n185_;
  assign new_n187_ = ~new_n181_ & new_n186_;
  assign new_n188_ = v5 & ~new_n187_;
  assign new_n189_ = ~v4 & new_n188_;
  assign new_n190_ = ~v3 & new_n189_;
  assign new_n191_ = ~v2 & new_n190_;
  assign new_n192_ = ~v1 & new_n191_;
  assign \v83.0  = ~v0 | new_n192_;
  assign new_n194_ = ~v14 & v15;
  assign new_n195_ = v13 & new_n194_;
  assign new_n196_ = ~v16 & ~new_n195_;
  assign new_n197_ = ~v19 & ~new_n196_;
  assign new_n198_ = ~v18 & new_n197_;
  assign new_n199_ = ~v17 & new_n198_;
  assign \v83.2  = v0 & new_n199_;
  assign new_n201_ = v17 & v18;
  assign new_n202_ = v0 & new_n201_;
  assign new_n203_ = ~v20 & ~new_n202_;
  assign \v83.3  = ~v19 & new_n203_;
  assign new_n205_ = ~v16 & v18;
  assign new_n206_ = ~v13 & v15;
  assign new_n207_ = v16 & ~v18;
  assign new_n208_ = new_n206_ & new_n207_;
  assign new_n209_ = ~new_n205_ & ~new_n208_;
  assign new_n210_ = v14 & ~new_n209_;
  assign new_n211_ = ~v13 & ~v15;
  assign new_n212_ = v18 & ~new_n211_;
  assign new_n213_ = ~v16 & new_n212_;
  assign new_n214_ = ~new_n210_ & ~new_n213_;
  assign new_n215_ = ~v19 & ~new_n214_;
  assign new_n216_ = v17 & new_n215_;
  assign \v83.4  = v0 & new_n216_;
  assign new_n218_ = v13 & v17;
  assign new_n219_ = v16 & ~new_n218_;
  assign new_n220_ = ~new_n194_ & ~new_n219_;
  assign new_n221_ = v13 & ~v17;
  assign new_n222_ = ~v16 & ~new_n221_;
  assign new_n223_ = ~new_n220_ & ~new_n222_;
  assign new_n224_ = ~v18 & ~new_n223_;
  assign new_n225_ = ~v14 & ~v15;
  assign new_n226_ = ~v13 & new_n225_;
  assign new_n227_ = v17 & ~new_n226_;
  assign new_n228_ = v18 & ~new_n227_;
  assign new_n229_ = v0 & ~v19;
  assign new_n230_ = ~new_n228_ & new_n229_;
  assign \v83.5  = new_n224_ | ~new_n230_;
  assign new_n232_ = v0 & ~v13;
  assign new_n233_ = ~v14 & new_n232_;
  assign new_n234_ = ~v15 & new_n233_;
  assign new_n235_ = v16 & new_n234_;
  assign new_n236_ = v17 & new_n235_;
  assign new_n237_ = ~v18 & new_n236_;
  assign \v83.6  = ~v19 & new_n237_;
  assign new_n239_ = v14 & ~v15;
  assign new_n240_ = ~v13 & new_n239_;
  assign new_n241_ = ~new_n212_ & ~new_n240_;
  assign new_n242_ = ~v19 & ~new_n241_;
  assign new_n243_ = v17 & new_n242_;
  assign new_n244_ = v16 & new_n243_;
  assign \v83.7  = v0 & new_n244_;
  assign new_n246_ = ~v22 & v23;
  assign new_n247_ = v22 & ~v23;
  assign new_n248_ = ~new_n246_ & ~new_n247_;
  assign new_n249_ = v21 & ~new_n248_;
  assign new_n250_ = v22 & v23;
  assign new_n251_ = ~v22 & ~v23;
  assign new_n252_ = ~new_n250_ & ~new_n251_;
  assign new_n253_ = ~v21 & ~new_n252_;
  assign \v83.9  = new_n249_ | new_n253_;
  assign new_n255_ = v21 & ~v22;
  assign new_n256_ = ~v21 & v22;
  assign new_n257_ = ~new_n255_ & ~new_n256_;
  assign new_n258_ = v24 & ~new_n257_;
  assign new_n259_ = v23 & v24;
  assign new_n260_ = v22 & ~new_n259_;
  assign new_n261_ = v21 & new_n260_;
  assign new_n262_ = ~v23 & v24;
  assign new_n263_ = ~v22 & ~new_n262_;
  assign new_n264_ = ~v21 & new_n263_;
  assign new_n265_ = ~new_n261_ & ~new_n264_;
  assign \v83.10  = new_n258_ | ~new_n265_;
  assign new_n267_ = v21 & v22;
  assign new_n268_ = ~v21 & ~v22;
  assign \v83.11  = new_n267_ | new_n268_;
  assign new_n270_ = v24 & ~new_n268_;
  assign new_n271_ = ~v22 & ~v24;
  assign new_n272_ = ~v21 & new_n271_;
  assign \v83.12  = new_n270_ | new_n272_;
  assign new_n274_ = ~v20 & ~new_n226_;
  assign new_n275_ = v18 & new_n274_;
  assign new_n276_ = v17 & new_n275_;
  assign new_n277_ = ~v16 & new_n276_;
  assign \v83.13  = v0 & new_n277_;
  assign new_n279_ = v13 & ~v14;
  assign new_n280_ = ~v16 & ~v17;
  assign new_n281_ = v15 & new_n280_;
  assign new_n282_ = new_n279_ & new_n281_;
  assign new_n283_ = v0 & ~new_n282_;
  assign new_n284_ = ~v18 & ~new_n283_;
  assign \v83.14  = ~v20 & ~new_n284_;
  assign new_n286_ = ~v9 & v11;
  assign new_n287_ = v8 & new_n286_;
  assign new_n288_ = v9 & ~v11;
  assign new_n289_ = ~new_n287_ & ~new_n288_;
  assign new_n290_ = v7 & ~new_n289_;
  assign new_n291_ = ~v8 & v9;
  assign new_n292_ = ~v7 & new_n291_;
  assign new_n293_ = v6 & ~new_n292_;
  assign new_n294_ = v11 & ~new_n293_;
  assign new_n295_ = ~new_n290_ & ~new_n294_;
  assign new_n296_ = v12 & ~new_n295_;
  assign \v83.15  = ~v10 & new_n296_;
  assign new_n298_ = ~v7 & v9;
  assign new_n299_ = ~v11 & ~new_n298_;
  assign new_n300_ = v10 & ~new_n299_;
  assign new_n301_ = ~v1 & ~v2;
  assign new_n302_ = ~v4 & v5;
  assign new_n303_ = ~v3 & new_n302_;
  assign new_n304_ = new_n301_ & new_n303_;
  assign new_n305_ = v25 & ~new_n304_;
  assign new_n306_ = ~v26 & v27;
  assign new_n307_ = ~new_n305_ & ~new_n306_;
  assign new_n308_ = v11 & ~new_n307_;
  assign new_n309_ = ~v9 & new_n308_;
  assign new_n310_ = v0 & new_n309_;
  assign new_n311_ = ~new_n300_ & ~new_n310_;
  assign new_n312_ = v8 & ~new_n311_;
  assign new_n313_ = ~v9 & ~new_n307_;
  assign new_n314_ = v0 & new_n313_;
  assign new_n315_ = ~v10 & ~new_n314_;
  assign new_n316_ = ~new_n182_ & ~new_n315_;
  assign new_n317_ = ~v10 & ~new_n307_;
  assign new_n318_ = ~v9 & new_n317_;
  assign new_n319_ = v0 & new_n318_;
  assign new_n320_ = ~new_n316_ & ~new_n319_;
  assign new_n321_ = v11 & ~new_n320_;
  assign new_n322_ = v10 & ~new_n288_;
  assign new_n323_ = v7 & ~new_n322_;
  assign new_n324_ = ~v8 & new_n288_;
  assign new_n325_ = ~new_n323_ & ~new_n324_;
  assign new_n326_ = v6 & ~new_n325_;
  assign new_n327_ = v8 & ~v9;
  assign new_n328_ = ~v10 & ~new_n327_;
  assign new_n329_ = ~new_n326_ & ~new_n328_;
  assign new_n330_ = ~new_n307_ & ~new_n329_;
  assign new_n331_ = v0 & new_n330_;
  assign new_n332_ = ~v6 & v9;
  assign new_n333_ = v10 & ~v11;
  assign new_n334_ = new_n332_ & new_n333_;
  assign new_n335_ = ~new_n331_ & ~new_n334_;
  assign new_n336_ = ~new_n321_ & new_n335_;
  assign new_n337_ = ~new_n312_ & new_n336_;
  assign \v83.16  = v12 & ~new_n337_;
  assign new_n339_ = v0 & v17;
  assign \v83.17  = ~v18 | ~new_n339_;
  assign new_n341_ = v12 & new_n305_;
  assign new_n342_ = v11 & new_n341_;
  assign new_n343_ = v10 & new_n342_;
  assign new_n344_ = ~v9 & new_n343_;
  assign new_n345_ = ~v8 & new_n344_;
  assign new_n346_ = ~v7 & new_n345_;
  assign new_n347_ = ~v6 & new_n346_;
  assign \v83.18  = v0 & new_n347_;
  assign new_n349_ = v0 & ~v6;
  assign new_n350_ = ~v7 & new_n349_;
  assign new_n351_ = ~v8 & new_n350_;
  assign new_n352_ = ~v9 & new_n351_;
  assign new_n353_ = v10 & new_n352_;
  assign new_n354_ = v11 & new_n353_;
  assign new_n355_ = v12 & new_n354_;
  assign new_n356_ = ~v26 & new_n355_;
  assign \v83.19  = v27 & new_n356_;
  assign new_n358_ = ~v0 & ~v18;
  assign \v83.20  = ~v20 & new_n358_;
  assign new_n360_ = v17 & ~new_n225_;
  assign new_n361_ = ~v13 & ~new_n360_;
  assign new_n362_ = ~v15 & v16;
  assign new_n363_ = ~v14 & new_n362_;
  assign new_n364_ = v15 & ~v16;
  assign new_n365_ = v14 & new_n364_;
  assign new_n366_ = ~new_n363_ & ~new_n365_;
  assign new_n367_ = ~v17 & ~new_n366_;
  assign new_n368_ = ~new_n361_ & ~new_n367_;
  assign new_n369_ = v18 & ~new_n368_;
  assign new_n370_ = ~v17 & ~new_n206_;
  assign new_n371_ = ~v18 & ~new_n370_;
  assign new_n372_ = ~v16 & new_n371_;
  assign new_n373_ = ~new_n369_ & ~new_n372_;
  assign new_n374_ = ~v20 & ~new_n373_;
  assign \v83.21  = v0 & new_n374_;
  assign new_n376_ = v0 & v16;
  assign \v83.22  = ~new_n201_ | ~new_n376_;
  assign new_n378_ = ~v18 & ~new_n211_;
  assign new_n379_ = v14 & ~new_n378_;
  assign new_n380_ = v15 & v18;
  assign new_n381_ = ~new_n379_ & ~new_n380_;
  assign new_n382_ = ~v20 & ~new_n381_;
  assign new_n383_ = v17 & new_n382_;
  assign new_n384_ = v16 & new_n383_;
  assign \v83.23  = v0 & new_n384_;
  assign new_n386_ = ~v36 & ~v38;
  assign new_n387_ = ~v35 & ~new_n386_;
  assign new_n388_ = v30 & v31;
  assign new_n389_ = ~v28 & ~new_n388_;
  assign new_n390_ = ~v30 & v31;
  assign new_n391_ = ~v29 & new_n390_;
  assign new_n392_ = v30 & ~v31;
  assign new_n393_ = v29 & new_n392_;
  assign new_n394_ = ~new_n391_ & ~new_n393_;
  assign new_n395_ = ~new_n389_ & new_n394_;
  assign new_n396_ = v33 & ~new_n395_;
  assign new_n397_ = ~v32 & new_n396_;
  assign new_n398_ = v32 & ~v33;
  assign new_n399_ = ~v31 & new_n398_;
  assign new_n400_ = ~new_n397_ & ~new_n399_;
  assign new_n401_ = ~new_n387_ & ~new_n400_;
  assign new_n402_ = v31 & new_n387_;
  assign new_n403_ = v35 & new_n386_;
  assign new_n404_ = ~new_n402_ & ~new_n403_;
  assign new_n405_ = v30 & ~new_n404_;
  assign new_n406_ = ~v28 & ~v30;
  assign new_n407_ = v31 & ~v35;
  assign new_n408_ = new_n406_ & new_n407_;
  assign new_n409_ = ~new_n405_ & ~new_n408_;
  assign new_n410_ = ~v33 & ~new_n409_;
  assign new_n411_ = v32 & new_n410_;
  assign new_n412_ = ~v29 & new_n411_;
  assign new_n413_ = ~new_n401_ & ~new_n412_;
  assign new_n414_ = v37 & ~new_n413_;
  assign \v83.24  = v34 & new_n414_;
  assign new_n416_ = ~v36 & ~v48;
  assign new_n417_ = ~v49 & ~v50;
  assign new_n418_ = new_n416_ & new_n417_;
  assign new_n419_ = v47 & ~new_n418_;
  assign new_n420_ = v32 & ~new_n419_;
  assign new_n421_ = ~v30 & new_n420_;
  assign new_n422_ = ~v29 & new_n421_;
  assign new_n423_ = ~v28 & new_n422_;
  assign new_n424_ = ~v32 & v35;
  assign new_n425_ = ~new_n423_ & ~new_n424_;
  assign new_n426_ = v37 & ~new_n425_;
  assign new_n427_ = v34 & new_n426_;
  assign new_n428_ = ~v33 & new_n427_;
  assign new_n429_ = ~v45 & v46;
  assign new_n430_ = ~new_n428_ & ~new_n429_;
  assign new_n431_ = v31 & ~new_n430_;
  assign new_n432_ = ~v29 & ~v30;
  assign new_n433_ = ~v28 & new_n432_;
  assign new_n434_ = v32 & ~new_n433_;
  assign new_n435_ = ~v33 & v34;
  assign new_n436_ = new_n434_ & new_n435_;
  assign new_n437_ = v46 & ~new_n436_;
  assign new_n438_ = ~v45 & new_n437_;
  assign new_n439_ = ~v39 & ~new_n438_;
  assign new_n440_ = ~new_n431_ & new_n439_;
  assign new_n441_ = ~v40 & ~new_n440_;
  assign new_n442_ = ~v41 & ~new_n441_;
  assign new_n443_ = ~v42 & ~new_n442_;
  assign new_n444_ = ~v43 & ~new_n443_;
  assign \v83.25  = ~v44 & ~new_n444_;
  assign new_n446_ = v37 & ~new_n419_;
  assign new_n447_ = v31 & new_n446_;
  assign new_n448_ = ~v30 & new_n447_;
  assign new_n449_ = ~v29 & new_n448_;
  assign new_n450_ = ~v28 & new_n449_;
  assign new_n451_ = ~v31 & ~new_n433_;
  assign new_n452_ = ~new_n450_ & ~new_n451_;
  assign new_n453_ = v32 & ~new_n452_;
  assign new_n454_ = v31 & ~v32;
  assign new_n455_ = v35 & v37;
  assign new_n456_ = new_n454_ & new_n455_;
  assign new_n457_ = ~new_n453_ & ~new_n456_;
  assign new_n458_ = ~v40 & ~new_n457_;
  assign new_n459_ = ~v39 & new_n458_;
  assign new_n460_ = v34 & new_n459_;
  assign new_n461_ = ~v33 & new_n460_;
  assign new_n462_ = ~v41 & ~v42;
  assign new_n463_ = ~new_n461_ & new_n462_;
  assign new_n464_ = ~v44 & ~new_n463_;
  assign \v83.26  = ~v43 & new_n464_;
  assign new_n466_ = v34 & ~new_n457_;
  assign new_n467_ = ~v33 & new_n466_;
  assign new_n468_ = ~v39 & ~v40;
  assign new_n469_ = ~new_n467_ & new_n468_;
  assign new_n470_ = ~v44 & ~new_n469_;
  assign new_n471_ = ~v43 & new_n470_;
  assign new_n472_ = ~v42 & new_n471_;
  assign \v83.27  = ~v41 & new_n472_;
  assign new_n474_ = ~v45 & ~v46;
  assign new_n475_ = v31 & v37;
  assign new_n476_ = ~new_n434_ & ~new_n475_;
  assign new_n477_ = ~new_n418_ & ~new_n451_;
  assign new_n478_ = v47 & new_n477_;
  assign new_n479_ = v31 & ~new_n433_;
  assign new_n480_ = ~new_n478_ & ~new_n479_;
  assign new_n481_ = v32 & ~new_n480_;
  assign new_n482_ = ~v32 & ~v35;
  assign new_n483_ = v31 & ~v37;
  assign new_n484_ = ~new_n482_ & ~new_n483_;
  assign new_n485_ = new_n435_ & new_n484_;
  assign new_n486_ = ~new_n481_ & new_n485_;
  assign new_n487_ = ~new_n476_ & new_n486_;
  assign new_n488_ = ~new_n474_ & ~new_n487_;
  assign new_n489_ = ~v44 & new_n488_;
  assign new_n490_ = ~v43 & new_n489_;
  assign new_n491_ = ~v42 & new_n490_;
  assign new_n492_ = ~v41 & new_n491_;
  assign new_n493_ = ~v40 & new_n492_;
  assign \v83.28  = ~v39 & new_n493_;
  assign new_n495_ = v17 & ~new_n207_;
  assign new_n496_ = v13 & ~new_n495_;
  assign new_n497_ = ~v15 & v18;
  assign new_n498_ = ~v13 & new_n497_;
  assign new_n499_ = ~new_n207_ & ~new_n498_;
  assign new_n500_ = ~v14 & ~new_n499_;
  assign new_n501_ = v16 & v18;
  assign new_n502_ = ~v15 & new_n501_;
  assign new_n503_ = ~v17 & ~new_n502_;
  assign new_n504_ = ~new_n500_ & ~new_n503_;
  assign new_n505_ = ~new_n496_ & new_n504_;
  assign \v83.29  = v0 & ~new_n505_;
  assign new_n507_ = ~v53 & v54;
  assign new_n508_ = ~v52 & new_n507_;
  assign new_n509_ = v53 & ~v54;
  assign new_n510_ = v52 & new_n509_;
  assign new_n511_ = ~new_n508_ & ~new_n510_;
  assign \v83.30  = v51 & ~new_n511_;
  assign new_n513_ = ~v15 & new_n232_;
  assign new_n514_ = ~v16 & new_n513_;
  assign new_n515_ = ~v17 & new_n514_;
  assign \v83.31  = v18 & new_n515_;
  assign new_n517_ = v11 & v12;
  assign new_n518_ = new_n327_ & new_n517_;
  assign new_n519_ = ~new_n288_ & ~new_n518_;
  assign new_n520_ = v7 & ~new_n519_;
  assign new_n521_ = v6 & v8;
  assign new_n522_ = ~v9 & ~v11;
  assign new_n523_ = new_n521_ & new_n522_;
  assign new_n524_ = new_n291_ & new_n517_;
  assign new_n525_ = ~new_n523_ & ~new_n524_;
  assign new_n526_ = ~v7 & ~new_n525_;
  assign new_n527_ = ~v6 & new_n517_;
  assign new_n528_ = ~new_n526_ & ~new_n527_;
  assign new_n529_ = ~new_n520_ & new_n528_;
  assign new_n530_ = ~v10 & ~new_n529_;
  assign new_n531_ = ~v11 & ~v12;
  assign \v83.32  = new_n530_ | new_n531_;
  assign new_n533_ = ~v1 & ~v3;
  assign new_n534_ = ~new_n187_ & ~new_n533_;
  assign new_n535_ = v5 & new_n534_;
  assign new_n536_ = ~v4 & new_n535_;
  assign new_n537_ = ~v2 & new_n536_;
  assign new_n538_ = ~v2 & new_n302_;
  assign new_n539_ = ~v9 & ~new_n286_;
  assign new_n540_ = v8 & new_n539_;
  assign new_n541_ = ~v10 & ~new_n540_;
  assign new_n542_ = ~new_n326_ & ~new_n541_;
  assign new_n543_ = ~new_n538_ & ~new_n542_;
  assign new_n544_ = v25 & new_n543_;
  assign new_n545_ = v12 & new_n544_;
  assign new_n546_ = ~new_n537_ & ~new_n545_;
  assign \v83.33  = v0 & ~new_n546_;
  assign new_n548_ = v0 & v13;
  assign new_n549_ = v16 & new_n548_;
  assign new_n550_ = ~v17 & new_n549_;
  assign new_n551_ = ~v18 & new_n550_;
  assign \v83.36  = ~v20 & new_n551_;
  assign new_n553_ = v0 & v15;
  assign new_n554_ = v16 & new_n553_;
  assign new_n555_ = ~v17 & new_n554_;
  assign \v83.37  = ~v18 & new_n555_;
  assign new_n557_ = v15 & new_n233_;
  assign new_n558_ = v16 & new_n557_;
  assign new_n559_ = ~v17 & new_n558_;
  assign new_n560_ = v18 & new_n559_;
  assign new_n561_ = ~v55 & new_n560_;
  assign new_n562_ = ~v56 & new_n561_;
  assign \v83.38  = v57 & new_n562_;
  assign new_n564_ = v56 & new_n561_;
  assign \v83.39  = v57 & new_n564_;
  assign new_n566_ = v55 & new_n560_;
  assign new_n567_ = ~v56 & new_n566_;
  assign \v83.40  = v57 & new_n567_;
  assign new_n569_ = v56 & new_n566_;
  assign \v83.41  = v57 & new_n569_;
  assign new_n571_ = v14 & new_n232_;
  assign new_n572_ = v15 & new_n571_;
  assign new_n573_ = v16 & new_n572_;
  assign new_n574_ = ~v17 & new_n573_;
  assign new_n575_ = v18 & new_n574_;
  assign new_n576_ = ~v55 & new_n575_;
  assign new_n577_ = ~v56 & new_n576_;
  assign \v83.42  = v57 & new_n577_;
  assign new_n579_ = v56 & new_n576_;
  assign \v83.43  = v57 & new_n579_;
  assign new_n581_ = v55 & new_n575_;
  assign new_n582_ = ~v56 & new_n581_;
  assign \v83.44  = v57 & new_n582_;
  assign new_n584_ = v56 & new_n581_;
  assign \v83.45  = v57 & new_n584_;
  assign new_n586_ = v0 & new_n279_;
  assign new_n587_ = ~v17 & ~v18;
  assign new_n588_ = new_n364_ & new_n587_;
  assign new_n589_ = new_n586_ & new_n588_;
  assign \v83.46  = ~v20 & ~new_n589_;
  assign new_n591_ = v6 & ~v7;
  assign new_n592_ = ~v9 & ~v10;
  assign new_n593_ = v8 & new_n592_;
  assign new_n594_ = new_n591_ & new_n593_;
  assign new_n595_ = v12 & ~new_n594_;
  assign \v83.47  = ~v11 & ~new_n595_;
  assign new_n597_ = v7 & v9;
  assign new_n598_ = ~v10 & new_n597_;
  assign new_n599_ = ~v11 & new_n598_;
  assign \v83.48  = v12 & new_n599_;
  assign new_n601_ = ~v14 & new_n207_;
  assign new_n602_ = ~new_n201_ & ~new_n601_;
  assign new_n603_ = v15 & ~new_n602_;
  assign new_n604_ = ~v18 & ~new_n218_;
  assign new_n605_ = v16 & new_n604_;
  assign new_n606_ = ~v13 & ~v14;
  assign new_n607_ = v18 & ~new_n606_;
  assign new_n608_ = v17 & new_n607_;
  assign new_n609_ = v0 & ~new_n608_;
  assign new_n610_ = ~new_n605_ & new_n609_;
  assign new_n611_ = ~new_n603_ & new_n610_;
  assign \v83.49  = ~v20 & ~new_n611_;
  assign new_n613_ = v16 & new_n587_;
  assign new_n614_ = v0 & ~new_n613_;
  assign new_n615_ = ~v20 & ~new_n614_;
  assign \v83.50  = ~v19 & new_n615_;
  assign new_n617_ = ~v54 & ~v63;
  assign new_n618_ = ~v51 & ~new_n617_;
  assign new_n619_ = v53 & ~v63;
  assign new_n620_ = v51 & new_n619_;
  assign new_n621_ = ~new_n507_ & ~new_n620_;
  assign new_n622_ = v52 & ~new_n621_;
  assign new_n623_ = v53 & v54;
  assign new_n624_ = ~v53 & v63;
  assign new_n625_ = ~new_n623_ & ~new_n624_;
  assign new_n626_ = ~v52 & ~new_n625_;
  assign new_n627_ = v59 & v62;
  assign new_n628_ = ~new_n626_ & ~new_n627_;
  assign new_n629_ = ~new_n622_ & new_n628_;
  assign new_n630_ = ~new_n618_ & new_n629_;
  assign new_n631_ = v61 & ~new_n630_;
  assign new_n632_ = v62 & ~v63;
  assign new_n633_ = v59 & new_n632_;
  assign new_n634_ = ~new_n631_ & ~new_n633_;
  assign new_n635_ = ~v60 & ~new_n634_;
  assign new_n636_ = ~v52 & new_n509_;
  assign new_n637_ = ~v53 & ~v54;
  assign new_n638_ = v53 & v63;
  assign new_n639_ = ~new_n637_ & ~new_n638_;
  assign new_n640_ = v52 & ~new_n639_;
  assign new_n641_ = ~new_n636_ & ~new_n640_;
  assign new_n642_ = v61 & ~new_n641_;
  assign new_n643_ = ~v53 & ~v63;
  assign new_n644_ = ~v52 & new_n643_;
  assign new_n645_ = ~new_n642_ & ~new_n644_;
  assign new_n646_ = v51 & ~new_n645_;
  assign new_n647_ = ~v51 & ~v54;
  assign new_n648_ = v61 & ~new_n647_;
  assign new_n649_ = ~v63 & ~new_n648_;
  assign new_n650_ = ~new_n646_ & ~new_n649_;
  assign new_n651_ = ~new_n627_ & ~new_n650_;
  assign new_n652_ = v60 & new_n651_;
  assign new_n653_ = ~new_n635_ & ~new_n652_;
  assign new_n654_ = ~v64 & ~new_n653_;
  assign new_n655_ = ~v52 & v53;
  assign new_n656_ = v52 & ~v53;
  assign new_n657_ = ~new_n655_ & ~new_n656_;
  assign new_n658_ = ~v59 & v60;
  assign new_n659_ = v51 & ~v54;
  assign new_n660_ = new_n658_ & new_n659_;
  assign new_n661_ = ~v58 & ~v60;
  assign new_n662_ = v54 & new_n661_;
  assign new_n663_ = ~new_n660_ & ~new_n662_;
  assign new_n664_ = ~new_n657_ & ~new_n663_;
  assign new_n665_ = v51 & v52;
  assign new_n666_ = v53 & ~v59;
  assign new_n667_ = new_n665_ & new_n666_;
  assign new_n668_ = ~v58 & ~new_n667_;
  assign new_n669_ = v60 & ~new_n668_;
  assign new_n670_ = ~v52 & ~v53;
  assign new_n671_ = ~v59 & ~new_n670_;
  assign new_n672_ = v51 & new_n671_;
  assign new_n673_ = ~v60 & ~new_n672_;
  assign new_n674_ = ~v58 & new_n673_;
  assign new_n675_ = ~new_n669_ & ~new_n674_;
  assign new_n676_ = v64 & ~new_n675_;
  assign new_n677_ = ~new_n664_ & ~new_n676_;
  assign new_n678_ = ~v63 & ~new_n677_;
  assign new_n679_ = ~v62 & new_n678_;
  assign new_n680_ = v61 & new_n679_;
  assign \v83.51  = new_n654_ | new_n680_;
  assign new_n682_ = new_n497_ & new_n606_;
  assign new_n683_ = v17 & ~new_n682_;
  assign new_n684_ = new_n376_ & new_n683_;
  assign new_n685_ = ~new_n378_ & new_n684_;
  assign \v83.52  = ~v20 & ~new_n685_;
  assign new_n687_ = v27 & ~new_n542_;
  assign new_n688_ = ~v26 & new_n687_;
  assign new_n689_ = v12 & new_n688_;
  assign \v83.53  = v0 & new_n689_;
  assign new_n691_ = v17 & new_n376_;
  assign \v83.54  = v18 & new_n691_;
  assign new_n693_ = ~v9 & v10;
  assign new_n694_ = v11 & new_n693_;
  assign \v83.55  = v12 & new_n694_;
  assign new_n696_ = v13 & v14;
  assign new_n697_ = v15 & ~new_n696_;
  assign new_n698_ = ~v17 & ~new_n697_;
  assign new_n699_ = ~v18 & ~new_n698_;
  assign new_n700_ = ~v16 & new_n699_;
  assign new_n701_ = ~new_n369_ & ~new_n700_;
  assign new_n702_ = ~v20 & ~new_n701_;
  assign new_n703_ = ~v19 & new_n702_;
  assign \v83.56  = v0 & new_n703_;
  assign new_n705_ = v2 & new_n190_;
  assign new_n706_ = v1 & new_n705_;
  assign \v83.57  = v0 & new_n706_;
  assign new_n708_ = ~v1 & new_n705_;
  assign \v83.58  = v0 & new_n708_;
  assign \v83.59  = v18 & new_n236_;
  assign new_n711_ = v16 & new_n201_;
  assign new_n712_ = v65 & ~new_n711_;
  assign \v83.60  = v0 & new_n712_;
  assign \v83.61  = ~v0 | new_n712_;
  assign new_n715_ = v3 & new_n189_;
  assign new_n716_ = v2 & new_n715_;
  assign \v83.63  = v0 & new_n716_;
  assign new_n718_ = ~v17 & v18;
  assign new_n719_ = v14 & new_n718_;
  assign new_n720_ = v17 & ~v18;
  assign new_n721_ = v16 & new_n720_;
  assign new_n722_ = ~new_n719_ & ~new_n721_;
  assign new_n723_ = ~v15 & ~new_n722_;
  assign new_n724_ = v16 & v17;
  assign new_n725_ = ~new_n280_ & ~new_n724_;
  assign new_n726_ = ~v18 & ~new_n725_;
  assign new_n727_ = v14 & new_n726_;
  assign new_n728_ = v15 & v16;
  assign new_n729_ = ~v14 & ~v16;
  assign new_n730_ = ~new_n728_ & ~new_n729_;
  assign new_n731_ = v18 & ~new_n730_;
  assign new_n732_ = ~v17 & new_n731_;
  assign new_n733_ = ~new_n727_ & ~new_n732_;
  assign new_n734_ = ~new_n723_ & new_n733_;
  assign new_n735_ = v13 & ~new_n734_;
  assign new_n736_ = ~v15 & ~v16;
  assign new_n737_ = new_n587_ & new_n736_;
  assign new_n738_ = ~new_n735_ & ~new_n737_;
  assign new_n739_ = v0 & ~new_n738_;
  assign \v83.64  = v66 | new_n739_;
  assign new_n741_ = v28 & v29;
  assign new_n742_ = v37 & ~new_n741_;
  assign new_n743_ = v34 & new_n742_;
  assign new_n744_ = v33 & new_n743_;
  assign new_n745_ = ~v32 & new_n744_;
  assign new_n746_ = v31 & new_n745_;
  assign \v83.65  = ~v30 & new_n746_;
  assign new_n748_ = ~v1 & new_n716_;
  assign \v83.66  = v0 & new_n748_;
  assign new_n750_ = v1 & new_n191_;
  assign \v83.67  = v0 & new_n750_;
  assign new_n752_ = v1 & new_n716_;
  assign \v83.68  = v0 & new_n752_;
  assign new_n754_ = ~v2 & new_n715_;
  assign new_n755_ = ~v1 & new_n754_;
  assign \v83.69  = v0 & new_n755_;
  assign new_n757_ = v1 & new_n754_;
  assign \v83.70  = v0 & new_n757_;
  assign new_n759_ = v13 & ~v15;
  assign new_n760_ = ~v18 & ~new_n759_;
  assign new_n761_ = v17 & new_n760_;
  assign new_n762_ = v16 & new_n761_;
  assign new_n763_ = ~v14 & new_n762_;
  assign \v83.71  = v0 & new_n763_;
  assign new_n765_ = ~v71 & ~v72;
  assign new_n766_ = v71 & v72;
  assign new_n767_ = v73 & v74;
  assign new_n768_ = ~new_n766_ & ~new_n767_;
  assign new_n769_ = ~new_n765_ & ~new_n768_;
  assign new_n770_ = v70 & ~new_n769_;
  assign new_n771_ = v68 & ~v69;
  assign new_n772_ = ~v67 & new_n771_;
  assign \v83.72  = new_n770_ | ~new_n772_;
  assign new_n774_ = ~new_n286_ & ~new_n328_;
  assign new_n775_ = ~new_n326_ & new_n774_;
  assign new_n776_ = v79 & ~new_n775_;
  assign new_n777_ = ~v78 & new_n776_;
  assign new_n778_ = ~v77 & new_n777_;
  assign new_n779_ = ~v76 & new_n778_;
  assign new_n780_ = v75 & new_n779_;
  assign \v83.73  = v12 & new_n780_;
  assign new_n782_ = v77 & new_n777_;
  assign new_n783_ = ~v76 & new_n782_;
  assign new_n784_ = ~v75 & new_n783_;
  assign \v83.74  = v12 & new_n784_;
  assign new_n786_ = v75 & new_n783_;
  assign \v83.75  = v12 & new_n786_;
  assign new_n788_ = v9 & v10;
  assign new_n789_ = v8 & new_n522_;
  assign new_n790_ = ~new_n788_ & ~new_n789_;
  assign new_n791_ = ~v6 & ~new_n790_;
  assign new_n792_ = ~new_n522_ & ~new_n788_;
  assign new_n793_ = ~v7 & ~new_n792_;
  assign new_n794_ = v10 & new_n517_;
  assign new_n795_ = ~new_n793_ & ~new_n794_;
  assign new_n796_ = v8 & ~new_n795_;
  assign new_n797_ = v12 & ~new_n182_;
  assign new_n798_ = ~v9 & ~new_n797_;
  assign new_n799_ = v11 & ~new_n798_;
  assign new_n800_ = ~new_n522_ & ~new_n799_;
  assign new_n801_ = v10 & ~new_n800_;
  assign new_n802_ = v12 & v25;
  assign new_n803_ = ~new_n304_ & new_n802_;
  assign new_n804_ = ~new_n801_ & new_n803_;
  assign new_n805_ = ~new_n796_ & new_n804_;
  assign new_n806_ = ~new_n791_ & new_n805_;
  assign \v83.76  = v0 & ~new_n806_;
  assign new_n808_ = v12 & new_n306_;
  assign new_n809_ = ~new_n801_ & new_n808_;
  assign new_n810_ = ~new_n796_ & new_n809_;
  assign new_n811_ = ~new_n791_ & new_n810_;
  assign \v83.77  = v0 & ~new_n811_;
  assign new_n813_ = v14 & ~new_n503_;
  assign new_n814_ = ~v13 & new_n813_;
  assign new_n815_ = ~v16 & ~v18;
  assign new_n816_ = ~new_n212_ & ~new_n815_;
  assign new_n817_ = v17 & ~new_n816_;
  assign new_n818_ = ~new_n814_ & ~new_n817_;
  assign \v83.78  = v0 & ~new_n818_;
  assign new_n820_ = ~v16 & new_n572_;
  assign new_n821_ = ~v17 & new_n820_;
  assign \v83.79  = v18 & new_n821_;
  assign new_n823_ = v14 & new_n548_;
  assign new_n824_ = v15 & new_n823_;
  assign new_n825_ = ~v16 & new_n824_;
  assign new_n826_ = ~v17 & new_n825_;
  assign \v83.80  = v18 & new_n826_;
  assign new_n828_ = ~v13 & ~v16;
  assign new_n829_ = ~v15 & ~new_n828_;
  assign new_n830_ = v14 & ~v16;
  assign new_n831_ = v13 & ~new_n830_;
  assign new_n832_ = v0 & new_n718_;
  assign new_n833_ = ~new_n831_ & new_n832_;
  assign \v83.81  = new_n829_ | ~new_n833_;
  assign new_n835_ = ~v16 & new_n557_;
  assign new_n836_ = ~v17 & new_n835_;
  assign \v83.82  = v18 & new_n836_;
  assign new_n838_ = ~v80 & v81;
  assign new_n839_ = v80 & v82;
  assign new_n840_ = v14 & new_n839_;
  assign new_n841_ = ~new_n838_ & ~new_n840_;
  assign new_n842_ = v18 & ~new_n841_;
  assign new_n843_ = ~v17 & new_n842_;
  assign new_n844_ = ~v16 & new_n843_;
  assign new_n845_ = ~v15 & new_n844_;
  assign new_n846_ = ~v13 & new_n845_;
  assign \v83.83  = v0 & new_n846_;
  assign new_n848_ = ~v14 & ~v80;
  assign new_n849_ = v81 & ~new_n848_;
  assign new_n850_ = v18 & new_n849_;
  assign new_n851_ = ~v17 & new_n850_;
  assign new_n852_ = ~v16 & new_n851_;
  assign new_n853_ = ~v15 & new_n852_;
  assign new_n854_ = ~v13 & new_n853_;
  assign \v83.84  = v0 & new_n854_;
  assign new_n856_ = ~v28 & ~v29;
  assign new_n857_ = ~v30 & new_n856_;
  assign new_n858_ = ~v31 & new_n857_;
  assign new_n859_ = v32 & new_n858_;
  assign new_n860_ = ~v33 & new_n859_;
  assign \v83.85  = v34 & new_n860_;
  assign new_n862_ = v16 & new_n513_;
  assign new_n863_ = v17 & new_n862_;
  assign \v83.86  = ~v18 & new_n863_;
  assign new_n865_ = ~v14 & new_n548_;
  assign new_n866_ = v15 & new_n865_;
  assign new_n867_ = ~v16 & new_n866_;
  assign new_n868_ = ~v17 & new_n867_;
  assign \v83.87  = ~v18 & new_n868_;
  assign new_n870_ = ~v8 & v10;
  assign new_n871_ = ~v7 & ~new_n870_;
  assign new_n872_ = ~v11 & ~new_n871_;
  assign new_n873_ = v6 & new_n872_;
  assign new_n874_ = ~v10 & v12;
  assign new_n875_ = v7 & new_n874_;
  assign new_n876_ = ~new_n873_ & ~new_n875_;
  assign new_n877_ = v9 & ~new_n876_;
  assign new_n878_ = v11 & ~new_n788_;
  assign new_n879_ = ~v6 & v8;
  assign new_n880_ = ~v10 & ~new_n879_;
  assign new_n881_ = ~v9 & new_n880_;
  assign new_n882_ = ~new_n878_ & ~new_n881_;
  assign new_n883_ = v12 & ~new_n882_;
  assign new_n884_ = ~new_n531_ & ~new_n883_;
  assign \v83.88  = new_n877_ | ~new_n884_;
  assign new_n886_ = v76 & new_n782_;
  assign new_n887_ = ~v75 & new_n886_;
  assign \v83.89  = v12 & new_n887_;
  assign new_n889_ = v75 & new_n886_;
  assign \v83.90  = v12 & new_n889_;
  assign new_n891_ = v76 & new_n778_;
  assign new_n892_ = v75 & new_n891_;
  assign \v83.91  = v12 & new_n892_;
  assign new_n894_ = ~v75 & new_n891_;
  assign \v83.92  = v12 & new_n894_;
  assign new_n896_ = v0 & ~v14;
  assign new_n897_ = v15 & new_n896_;
  assign new_n898_ = v16 & new_n897_;
  assign new_n899_ = v17 & new_n898_;
  assign new_n900_ = ~v18 & new_n899_;
  assign \v83.93  = ~v19 & new_n900_;
  assign \v83.1  = ~v0;
  assign \v83.8  = ~v21;
  assign \v83.34  = \v83.32 ;
  assign \v83.35  = \v83.20 ;
  assign \v83.62  = \v83.17 ;
endmodule


