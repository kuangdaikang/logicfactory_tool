// Benchmark "c499.blif" written by ABC on Fri Feb 25 15:13:01 2022

module c499  ( 
    Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9, Gid10,
    Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19, Gid20,
    Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29, Gid30,
    Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr,
    God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10,
    God11, God12, God13, God14, God15, God16, God17, God18, God19, God20,
    God21, God22, God23, God24, God25, God26, God27, God28, God29, God30,
    God31  );
  input  Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9,
    Gid10, Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19,
    Gid20, Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29,
    Gid30, Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr;
  output God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10,
    God11, God12, God13, God14, God15, God16, God17, God18, God19, God20,
    God21, God22, God23, God24, God25, God26, God27, God28, God29, God30,
    God31;
  wire new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n320_, new_n321_, new_n322_, new_n324_, new_n325_,
    new_n326_, new_n328_, new_n329_, new_n330_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n339_, new_n340_,
    new_n341_, new_n343_, new_n344_, new_n345_, new_n347_, new_n348_,
    new_n349_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n359_, new_n360_, new_n361_, new_n363_,
    new_n364_, new_n365_, new_n367_, new_n368_, new_n369_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n378_,
    new_n379_, new_n380_, new_n382_, new_n383_, new_n384_, new_n386_,
    new_n387_, new_n388_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n407_, new_n408_, new_n409_, new_n411_, new_n412_, new_n413_,
    new_n415_, new_n416_, new_n417_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n425_, new_n426_, new_n427_, new_n429_,
    new_n430_, new_n431_, new_n433_, new_n434_, new_n435_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n444_,
    new_n445_, new_n446_, new_n448_, new_n449_, new_n450_, new_n452_,
    new_n453_, new_n454_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n462_, new_n463_, new_n464_, new_n466_, new_n467_,
    new_n468_, new_n470_, new_n471_, new_n472_;
  assign new_n74_ = ~Gid0 & Gid4;
  assign new_n75_ = Gid0 & ~Gid4;
  assign new_n76_ = ~new_n74_ & ~new_n75_;
  assign new_n77_ = ~Gid8 & Gid12;
  assign new_n78_ = Gid8 & ~Gid12;
  assign new_n79_ = ~new_n77_ & ~new_n78_;
  assign new_n80_ = new_n76_ & ~new_n79_;
  assign new_n81_ = ~new_n76_ & new_n79_;
  assign new_n82_ = ~new_n80_ & ~new_n81_;
  assign new_n83_ = Gic0 & Gr;
  assign new_n84_ = ~Gid16 & Gid17;
  assign new_n85_ = Gid16 & ~Gid17;
  assign new_n86_ = ~new_n84_ & ~new_n85_;
  assign new_n87_ = ~Gid18 & Gid19;
  assign new_n88_ = Gid18 & ~Gid19;
  assign new_n89_ = ~new_n87_ & ~new_n88_;
  assign new_n90_ = new_n86_ & ~new_n89_;
  assign new_n91_ = ~new_n86_ & new_n89_;
  assign new_n92_ = ~new_n90_ & ~new_n91_;
  assign new_n93_ = ~Gid20 & Gid21;
  assign new_n94_ = Gid20 & ~Gid21;
  assign new_n95_ = ~new_n93_ & ~new_n94_;
  assign new_n96_ = ~Gid22 & Gid23;
  assign new_n97_ = Gid22 & ~Gid23;
  assign new_n98_ = ~new_n96_ & ~new_n97_;
  assign new_n99_ = new_n95_ & ~new_n98_;
  assign new_n100_ = ~new_n95_ & new_n98_;
  assign new_n101_ = ~new_n99_ & ~new_n100_;
  assign new_n102_ = new_n92_ & ~new_n101_;
  assign new_n103_ = ~new_n92_ & new_n101_;
  assign new_n104_ = ~new_n102_ & ~new_n103_;
  assign new_n105_ = ~new_n83_ & ~new_n104_;
  assign new_n106_ = new_n83_ & new_n104_;
  assign new_n107_ = ~new_n105_ & ~new_n106_;
  assign new_n108_ = new_n82_ & ~new_n107_;
  assign new_n109_ = ~new_n82_ & new_n107_;
  assign new_n110_ = ~new_n108_ & ~new_n109_;
  assign new_n111_ = ~Gid16 & Gid20;
  assign new_n112_ = Gid16 & ~Gid20;
  assign new_n113_ = ~new_n111_ & ~new_n112_;
  assign new_n114_ = ~Gid24 & Gid28;
  assign new_n115_ = Gid24 & ~Gid28;
  assign new_n116_ = ~new_n114_ & ~new_n115_;
  assign new_n117_ = new_n113_ & ~new_n116_;
  assign new_n118_ = ~new_n113_ & new_n116_;
  assign new_n119_ = ~new_n117_ & ~new_n118_;
  assign new_n120_ = Gic4 & Gr;
  assign new_n121_ = ~Gid0 & Gid1;
  assign new_n122_ = Gid0 & ~Gid1;
  assign new_n123_ = ~new_n121_ & ~new_n122_;
  assign new_n124_ = ~Gid2 & Gid3;
  assign new_n125_ = Gid2 & ~Gid3;
  assign new_n126_ = ~new_n124_ & ~new_n125_;
  assign new_n127_ = new_n123_ & ~new_n126_;
  assign new_n128_ = ~new_n123_ & new_n126_;
  assign new_n129_ = ~new_n127_ & ~new_n128_;
  assign new_n130_ = ~Gid4 & Gid5;
  assign new_n131_ = Gid4 & ~Gid5;
  assign new_n132_ = ~new_n130_ & ~new_n131_;
  assign new_n133_ = ~Gid6 & Gid7;
  assign new_n134_ = Gid6 & ~Gid7;
  assign new_n135_ = ~new_n133_ & ~new_n134_;
  assign new_n136_ = new_n132_ & ~new_n135_;
  assign new_n137_ = ~new_n132_ & new_n135_;
  assign new_n138_ = ~new_n136_ & ~new_n137_;
  assign new_n139_ = new_n129_ & ~new_n138_;
  assign new_n140_ = ~new_n129_ & new_n138_;
  assign new_n141_ = ~new_n139_ & ~new_n140_;
  assign new_n142_ = ~new_n120_ & ~new_n141_;
  assign new_n143_ = new_n120_ & new_n141_;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = new_n119_ & ~new_n144_;
  assign new_n146_ = ~new_n119_ & new_n144_;
  assign new_n147_ = ~new_n145_ & ~new_n146_;
  assign new_n148_ = ~Gid17 & Gid21;
  assign new_n149_ = Gid17 & ~Gid21;
  assign new_n150_ = ~new_n148_ & ~new_n149_;
  assign new_n151_ = ~Gid25 & Gid29;
  assign new_n152_ = Gid25 & ~Gid29;
  assign new_n153_ = ~new_n151_ & ~new_n152_;
  assign new_n154_ = new_n150_ & ~new_n153_;
  assign new_n155_ = ~new_n150_ & new_n153_;
  assign new_n156_ = ~new_n154_ & ~new_n155_;
  assign new_n157_ = Gic5 & Gr;
  assign new_n158_ = ~Gid8 & Gid9;
  assign new_n159_ = Gid8 & ~Gid9;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_ = ~Gid10 & Gid11;
  assign new_n162_ = Gid10 & ~Gid11;
  assign new_n163_ = ~new_n161_ & ~new_n162_;
  assign new_n164_ = new_n160_ & ~new_n163_;
  assign new_n165_ = ~new_n160_ & new_n163_;
  assign new_n166_ = ~new_n164_ & ~new_n165_;
  assign new_n167_ = ~Gid12 & Gid13;
  assign new_n168_ = Gid12 & ~Gid13;
  assign new_n169_ = ~new_n167_ & ~new_n168_;
  assign new_n170_ = ~Gid14 & Gid15;
  assign new_n171_ = Gid14 & ~Gid15;
  assign new_n172_ = ~new_n170_ & ~new_n171_;
  assign new_n173_ = new_n169_ & ~new_n172_;
  assign new_n174_ = ~new_n169_ & new_n172_;
  assign new_n175_ = ~new_n173_ & ~new_n174_;
  assign new_n176_ = new_n166_ & ~new_n175_;
  assign new_n177_ = ~new_n166_ & new_n175_;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = ~new_n157_ & ~new_n178_;
  assign new_n180_ = new_n157_ & new_n178_;
  assign new_n181_ = ~new_n179_ & ~new_n180_;
  assign new_n182_ = new_n156_ & ~new_n181_;
  assign new_n183_ = ~new_n156_ & new_n181_;
  assign new_n184_ = ~new_n182_ & ~new_n183_;
  assign new_n185_ = ~Gid18 & Gid22;
  assign new_n186_ = Gid18 & ~Gid22;
  assign new_n187_ = ~new_n185_ & ~new_n186_;
  assign new_n188_ = ~Gid26 & Gid30;
  assign new_n189_ = Gid26 & ~Gid30;
  assign new_n190_ = ~new_n188_ & ~new_n189_;
  assign new_n191_ = new_n187_ & ~new_n190_;
  assign new_n192_ = ~new_n187_ & new_n190_;
  assign new_n193_ = ~new_n191_ & ~new_n192_;
  assign new_n194_ = Gic6 & Gr;
  assign new_n195_ = new_n129_ & ~new_n166_;
  assign new_n196_ = ~new_n129_ & new_n166_;
  assign new_n197_ = ~new_n195_ & ~new_n196_;
  assign new_n198_ = ~new_n194_ & ~new_n197_;
  assign new_n199_ = new_n194_ & new_n197_;
  assign new_n200_ = ~new_n198_ & ~new_n199_;
  assign new_n201_ = new_n193_ & ~new_n200_;
  assign new_n202_ = ~new_n193_ & new_n200_;
  assign new_n203_ = ~new_n201_ & ~new_n202_;
  assign new_n204_ = ~Gid19 & Gid23;
  assign new_n205_ = Gid19 & ~Gid23;
  assign new_n206_ = ~new_n204_ & ~new_n205_;
  assign new_n207_ = ~Gid27 & Gid31;
  assign new_n208_ = Gid27 & ~Gid31;
  assign new_n209_ = ~new_n207_ & ~new_n208_;
  assign new_n210_ = new_n206_ & ~new_n209_;
  assign new_n211_ = ~new_n206_ & new_n209_;
  assign new_n212_ = ~new_n210_ & ~new_n211_;
  assign new_n213_ = Gic7 & Gr;
  assign new_n214_ = new_n138_ & ~new_n175_;
  assign new_n215_ = ~new_n138_ & new_n175_;
  assign new_n216_ = ~new_n214_ & ~new_n215_;
  assign new_n217_ = ~new_n213_ & ~new_n216_;
  assign new_n218_ = new_n213_ & new_n216_;
  assign new_n219_ = ~new_n217_ & ~new_n218_;
  assign new_n220_ = new_n212_ & ~new_n219_;
  assign new_n221_ = ~new_n212_ & new_n219_;
  assign new_n222_ = ~new_n220_ & ~new_n221_;
  assign new_n223_ = ~Gid1 & Gid5;
  assign new_n224_ = Gid1 & ~Gid5;
  assign new_n225_ = ~new_n223_ & ~new_n224_;
  assign new_n226_ = ~Gid9 & Gid13;
  assign new_n227_ = Gid9 & ~Gid13;
  assign new_n228_ = ~new_n226_ & ~new_n227_;
  assign new_n229_ = new_n225_ & ~new_n228_;
  assign new_n230_ = ~new_n225_ & new_n228_;
  assign new_n231_ = ~new_n229_ & ~new_n230_;
  assign new_n232_ = Gic1 & Gr;
  assign new_n233_ = ~Gid24 & Gid25;
  assign new_n234_ = Gid24 & ~Gid25;
  assign new_n235_ = ~new_n233_ & ~new_n234_;
  assign new_n236_ = ~Gid26 & Gid27;
  assign new_n237_ = Gid26 & ~Gid27;
  assign new_n238_ = ~new_n236_ & ~new_n237_;
  assign new_n239_ = new_n235_ & ~new_n238_;
  assign new_n240_ = ~new_n235_ & new_n238_;
  assign new_n241_ = ~new_n239_ & ~new_n240_;
  assign new_n242_ = ~Gid28 & Gid29;
  assign new_n243_ = Gid28 & ~Gid29;
  assign new_n244_ = ~new_n242_ & ~new_n243_;
  assign new_n245_ = ~Gid30 & Gid31;
  assign new_n246_ = Gid30 & ~Gid31;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign new_n248_ = new_n244_ & ~new_n247_;
  assign new_n249_ = ~new_n244_ & new_n247_;
  assign new_n250_ = ~new_n248_ & ~new_n249_;
  assign new_n251_ = new_n241_ & ~new_n250_;
  assign new_n252_ = ~new_n241_ & new_n250_;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign new_n254_ = ~new_n232_ & ~new_n253_;
  assign new_n255_ = new_n232_ & new_n253_;
  assign new_n256_ = ~new_n254_ & ~new_n255_;
  assign new_n257_ = new_n231_ & ~new_n256_;
  assign new_n258_ = ~new_n231_ & new_n256_;
  assign new_n259_ = ~new_n257_ & ~new_n258_;
  assign new_n260_ = ~Gid2 & Gid6;
  assign new_n261_ = Gid2 & ~Gid6;
  assign new_n262_ = ~new_n260_ & ~new_n261_;
  assign new_n263_ = ~Gid10 & Gid14;
  assign new_n264_ = Gid10 & ~Gid14;
  assign new_n265_ = ~new_n263_ & ~new_n264_;
  assign new_n266_ = new_n262_ & ~new_n265_;
  assign new_n267_ = ~new_n262_ & new_n265_;
  assign new_n268_ = ~new_n266_ & ~new_n267_;
  assign new_n269_ = Gic2 & Gr;
  assign new_n270_ = new_n92_ & ~new_n241_;
  assign new_n271_ = ~new_n92_ & new_n241_;
  assign new_n272_ = ~new_n270_ & ~new_n271_;
  assign new_n273_ = ~new_n269_ & ~new_n272_;
  assign new_n274_ = new_n269_ & new_n272_;
  assign new_n275_ = ~new_n273_ & ~new_n274_;
  assign new_n276_ = new_n268_ & ~new_n275_;
  assign new_n277_ = ~new_n268_ & new_n275_;
  assign new_n278_ = ~new_n276_ & ~new_n277_;
  assign new_n279_ = ~Gid3 & Gid7;
  assign new_n280_ = Gid3 & ~Gid7;
  assign new_n281_ = ~new_n279_ & ~new_n280_;
  assign new_n282_ = ~Gid11 & Gid15;
  assign new_n283_ = Gid11 & ~Gid15;
  assign new_n284_ = ~new_n282_ & ~new_n283_;
  assign new_n285_ = new_n281_ & ~new_n284_;
  assign new_n286_ = ~new_n281_ & new_n284_;
  assign new_n287_ = ~new_n285_ & ~new_n286_;
  assign new_n288_ = Gic3 & Gr;
  assign new_n289_ = new_n101_ & ~new_n250_;
  assign new_n290_ = ~new_n101_ & new_n250_;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = ~new_n288_ & ~new_n291_;
  assign new_n293_ = new_n288_ & new_n291_;
  assign new_n294_ = ~new_n292_ & ~new_n293_;
  assign new_n295_ = new_n287_ & ~new_n294_;
  assign new_n296_ = ~new_n287_ & new_n294_;
  assign new_n297_ = ~new_n295_ & ~new_n296_;
  assign new_n298_ = new_n110_ & new_n259_;
  assign new_n299_ = new_n278_ & new_n298_;
  assign new_n300_ = ~new_n297_ & new_n299_;
  assign new_n301_ = ~new_n278_ & new_n298_;
  assign new_n302_ = new_n297_ & new_n301_;
  assign new_n303_ = new_n110_ & ~new_n259_;
  assign new_n304_ = new_n278_ & new_n303_;
  assign new_n305_ = new_n297_ & new_n304_;
  assign new_n306_ = ~new_n110_ & new_n259_;
  assign new_n307_ = new_n278_ & new_n306_;
  assign new_n308_ = new_n297_ & new_n307_;
  assign new_n309_ = ~new_n305_ & ~new_n308_;
  assign new_n310_ = ~new_n300_ & ~new_n302_;
  assign new_n311_ = new_n309_ & new_n310_;
  assign new_n312_ = ~new_n147_ & new_n184_;
  assign new_n313_ = ~new_n203_ & new_n312_;
  assign new_n314_ = new_n222_ & new_n313_;
  assign new_n315_ = ~new_n311_ & new_n314_;
  assign new_n316_ = ~new_n110_ & new_n315_;
  assign new_n317_ = ~Gid0 & new_n316_;
  assign new_n318_ = Gid0 & ~new_n316_;
  assign God0 = new_n317_ | new_n318_;
  assign new_n320_ = ~new_n259_ & new_n315_;
  assign new_n321_ = ~Gid1 & new_n320_;
  assign new_n322_ = Gid1 & ~new_n320_;
  assign God1 = new_n321_ | new_n322_;
  assign new_n324_ = ~new_n278_ & new_n315_;
  assign new_n325_ = ~Gid2 & new_n324_;
  assign new_n326_ = Gid2 & ~new_n324_;
  assign God2 = new_n325_ | new_n326_;
  assign new_n328_ = ~new_n297_ & new_n315_;
  assign new_n329_ = ~Gid3 & new_n328_;
  assign new_n330_ = Gid3 & ~new_n328_;
  assign God3 = new_n329_ | new_n330_;
  assign new_n332_ = new_n203_ & new_n312_;
  assign new_n333_ = ~new_n222_ & new_n332_;
  assign new_n334_ = ~new_n311_ & new_n333_;
  assign new_n335_ = ~new_n110_ & new_n334_;
  assign new_n336_ = ~Gid4 & new_n335_;
  assign new_n337_ = Gid4 & ~new_n335_;
  assign God4 = new_n336_ | new_n337_;
  assign new_n339_ = ~new_n259_ & new_n334_;
  assign new_n340_ = ~Gid5 & new_n339_;
  assign new_n341_ = Gid5 & ~new_n339_;
  assign God5 = new_n340_ | new_n341_;
  assign new_n343_ = ~new_n278_ & new_n334_;
  assign new_n344_ = ~Gid6 & new_n343_;
  assign new_n345_ = Gid6 & ~new_n343_;
  assign God6 = new_n344_ | new_n345_;
  assign new_n347_ = ~new_n297_ & new_n334_;
  assign new_n348_ = ~Gid7 & new_n347_;
  assign new_n349_ = Gid7 & ~new_n347_;
  assign God7 = new_n348_ | new_n349_;
  assign new_n351_ = new_n147_ & ~new_n184_;
  assign new_n352_ = ~new_n203_ & new_n351_;
  assign new_n353_ = new_n222_ & new_n352_;
  assign new_n354_ = ~new_n311_ & new_n353_;
  assign new_n355_ = ~new_n110_ & new_n354_;
  assign new_n356_ = ~Gid8 & new_n355_;
  assign new_n357_ = Gid8 & ~new_n355_;
  assign God8 = new_n356_ | new_n357_;
  assign new_n359_ = ~new_n259_ & new_n354_;
  assign new_n360_ = ~Gid9 & new_n359_;
  assign new_n361_ = Gid9 & ~new_n359_;
  assign God9 = new_n360_ | new_n361_;
  assign new_n363_ = ~new_n278_ & new_n354_;
  assign new_n364_ = ~Gid10 & new_n363_;
  assign new_n365_ = Gid10 & ~new_n363_;
  assign God10 = new_n364_ | new_n365_;
  assign new_n367_ = ~new_n297_ & new_n354_;
  assign new_n368_ = ~Gid11 & new_n367_;
  assign new_n369_ = Gid11 & ~new_n367_;
  assign God11 = new_n368_ | new_n369_;
  assign new_n371_ = new_n203_ & new_n351_;
  assign new_n372_ = ~new_n222_ & new_n371_;
  assign new_n373_ = ~new_n311_ & new_n372_;
  assign new_n374_ = ~new_n110_ & new_n373_;
  assign new_n375_ = ~Gid12 & new_n374_;
  assign new_n376_ = Gid12 & ~new_n374_;
  assign God12 = new_n375_ | new_n376_;
  assign new_n378_ = ~new_n259_ & new_n373_;
  assign new_n379_ = ~Gid13 & new_n378_;
  assign new_n380_ = Gid13 & ~new_n378_;
  assign God13 = new_n379_ | new_n380_;
  assign new_n382_ = ~new_n278_ & new_n373_;
  assign new_n383_ = ~Gid14 & new_n382_;
  assign new_n384_ = Gid14 & ~new_n382_;
  assign God14 = new_n383_ | new_n384_;
  assign new_n386_ = ~new_n297_ & new_n373_;
  assign new_n387_ = ~Gid15 & new_n386_;
  assign new_n388_ = Gid15 & ~new_n386_;
  assign God15 = new_n387_ | new_n388_;
  assign new_n390_ = new_n147_ & new_n184_;
  assign new_n391_ = new_n203_ & new_n390_;
  assign new_n392_ = ~new_n222_ & new_n391_;
  assign new_n393_ = ~new_n203_ & new_n390_;
  assign new_n394_ = new_n222_ & new_n393_;
  assign new_n395_ = new_n222_ & new_n371_;
  assign new_n396_ = new_n222_ & new_n332_;
  assign new_n397_ = ~new_n395_ & ~new_n396_;
  assign new_n398_ = ~new_n392_ & ~new_n394_;
  assign new_n399_ = new_n397_ & new_n398_;
  assign new_n400_ = ~new_n278_ & new_n306_;
  assign new_n401_ = new_n297_ & new_n400_;
  assign new_n402_ = ~new_n399_ & new_n401_;
  assign new_n403_ = ~new_n147_ & new_n402_;
  assign new_n404_ = ~Gid16 & new_n403_;
  assign new_n405_ = Gid16 & ~new_n403_;
  assign God16 = new_n404_ | new_n405_;
  assign new_n407_ = ~new_n184_ & new_n402_;
  assign new_n408_ = ~Gid17 & new_n407_;
  assign new_n409_ = Gid17 & ~new_n407_;
  assign God17 = new_n408_ | new_n409_;
  assign new_n411_ = ~new_n203_ & new_n402_;
  assign new_n412_ = ~Gid18 & new_n411_;
  assign new_n413_ = Gid18 & ~new_n411_;
  assign God18 = new_n412_ | new_n413_;
  assign new_n415_ = ~new_n222_ & new_n402_;
  assign new_n416_ = ~Gid19 & new_n415_;
  assign new_n417_ = Gid19 & ~new_n415_;
  assign God19 = new_n416_ | new_n417_;
  assign new_n419_ = ~new_n297_ & new_n307_;
  assign new_n420_ = ~new_n399_ & new_n419_;
  assign new_n421_ = ~new_n147_ & new_n420_;
  assign new_n422_ = ~Gid20 & new_n421_;
  assign new_n423_ = Gid20 & ~new_n421_;
  assign God20 = new_n422_ | new_n423_;
  assign new_n425_ = ~new_n184_ & new_n420_;
  assign new_n426_ = ~Gid21 & new_n425_;
  assign new_n427_ = Gid21 & ~new_n425_;
  assign God21 = new_n426_ | new_n427_;
  assign new_n429_ = ~new_n203_ & new_n420_;
  assign new_n430_ = ~Gid22 & new_n429_;
  assign new_n431_ = Gid22 & ~new_n429_;
  assign God22 = new_n430_ | new_n431_;
  assign new_n433_ = ~new_n222_ & new_n420_;
  assign new_n434_ = ~Gid23 & new_n433_;
  assign new_n435_ = Gid23 & ~new_n433_;
  assign God23 = new_n434_ | new_n435_;
  assign new_n437_ = ~new_n278_ & new_n303_;
  assign new_n438_ = new_n297_ & new_n437_;
  assign new_n439_ = ~new_n399_ & new_n438_;
  assign new_n440_ = ~new_n147_ & new_n439_;
  assign new_n441_ = ~Gid24 & new_n440_;
  assign new_n442_ = Gid24 & ~new_n440_;
  assign God24 = new_n441_ | new_n442_;
  assign new_n444_ = ~new_n184_ & new_n439_;
  assign new_n445_ = ~Gid25 & new_n444_;
  assign new_n446_ = Gid25 & ~new_n444_;
  assign God25 = new_n445_ | new_n446_;
  assign new_n448_ = ~new_n203_ & new_n439_;
  assign new_n449_ = ~Gid26 & new_n448_;
  assign new_n450_ = Gid26 & ~new_n448_;
  assign God26 = new_n449_ | new_n450_;
  assign new_n452_ = ~new_n222_ & new_n439_;
  assign new_n453_ = ~Gid27 & new_n452_;
  assign new_n454_ = Gid27 & ~new_n452_;
  assign God27 = new_n453_ | new_n454_;
  assign new_n456_ = ~new_n297_ & new_n304_;
  assign new_n457_ = ~new_n399_ & new_n456_;
  assign new_n458_ = ~new_n147_ & new_n457_;
  assign new_n459_ = ~Gid28 & new_n458_;
  assign new_n460_ = Gid28 & ~new_n458_;
  assign God28 = new_n459_ | new_n460_;
  assign new_n462_ = ~new_n184_ & new_n457_;
  assign new_n463_ = ~Gid29 & new_n462_;
  assign new_n464_ = Gid29 & ~new_n462_;
  assign God29 = new_n463_ | new_n464_;
  assign new_n466_ = ~new_n203_ & new_n457_;
  assign new_n467_ = ~Gid30 & new_n466_;
  assign new_n468_ = Gid30 & ~new_n466_;
  assign God30 = new_n467_ | new_n468_;
  assign new_n470_ = ~new_n222_ & new_n457_;
  assign new_n471_ = ~Gid31 & new_n470_;
  assign new_n472_ = Gid31 & ~new_n470_;
  assign God31 = new_n471_ | new_n472_;
endmodule


