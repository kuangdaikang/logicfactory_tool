// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:54 2022

module bca  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25,
    \v26.0 , \v26.1 , \v26.2 , \v26.3 , \v26.4 , \v26.5 , \v26.6 , \v26.7 ,
    \v26.8 , \v26.9 , \v26.10 , \v26.11 , \v26.12 , \v26.13 , \v26.14 ,
    \v26.15 , \v26.16 , \v26.17 , \v26.18 , \v26.19 , \v26.20 , \v26.21 ,
    \v26.22 , \v26.23 , \v26.24 , \v26.25 , \v26.26 , \v26.27 , \v26.28 ,
    \v26.29 , \v26.30 , \v26.31 , \v26.32 , \v26.33 , \v26.34 , \v26.35 ,
    \v26.36 , \v26.37 , \v26.38 , \v26.39 , \v26.40 , \v26.41 , \v26.42 ,
    \v26.43 , \v26.44 , \v26.45   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25;
  output \v26.0 , \v26.1 , \v26.2 , \v26.3 , \v26.4 , \v26.5 , \v26.6 ,
    \v26.7 , \v26.8 , \v26.9 , \v26.10 , \v26.11 , \v26.12 , \v26.13 ,
    \v26.14 , \v26.15 , \v26.16 , \v26.17 , \v26.18 , \v26.19 , \v26.20 ,
    \v26.21 , \v26.22 , \v26.23 , \v26.24 , \v26.25 , \v26.26 , \v26.27 ,
    \v26.28 , \v26.29 , \v26.30 , \v26.31 , \v26.32 , \v26.33 , \v26.34 ,
    \v26.35 , \v26.36 , \v26.37 , \v26.38 , \v26.39 , \v26.40 , \v26.41 ,
    \v26.42 , \v26.43 , \v26.44 , \v26.45 ;
  wire new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2148_, new_n2149_, new_n2150_, new_n2151_,
    new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_,
    new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_,
    new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_,
    new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_,
    new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_,
    new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_,
    new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_,
    new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_,
    new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_,
    new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_,
    new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_,
    new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_,
    new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_,
    new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_,
    new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_,
    new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_,
    new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_,
    new_n2321_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2564_,
    new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_,
    new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_,
    new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_,
    new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_,
    new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_,
    new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_,
    new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_,
    new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_,
    new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_,
    new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_,
    new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_,
    new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_,
    new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_,
    new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2709_, new_n2710_,
    new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_,
    new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_,
    new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_,
    new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_,
    new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_,
    new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_,
    new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_,
    new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3147_, new_n3148_, new_n3149_, new_n3150_,
    new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_,
    new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_,
    new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_,
    new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_,
    new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_,
    new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_,
    new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_,
    new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_,
    new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_,
    new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_,
    new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_,
    new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_,
    new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_,
    new_n3242_, new_n3243_, new_n3244_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_,
    new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_,
    new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_,
    new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_,
    new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_,
    new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_,
    new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_,
    new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_,
    new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_,
    new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_,
    new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_,
    new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_,
    new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_,
    new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3587_, new_n3588_,
    new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_,
    new_n3595_, new_n3596_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_,
    new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_,
    new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_,
    new_n3621_, new_n3622_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_,
    new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_,
    new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_,
    new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_,
    new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_,
    new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_,
    new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_,
    new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_,
    new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_,
    new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_,
    new_n3739_, new_n3740_;
  assign new_n73_ = v5 & ~v7;
  assign new_n74_ = v5 & ~new_n73_;
  assign new_n75_ = ~v6 & ~new_n74_;
  assign new_n76_ = v7 & v10;
  assign new_n77_ = ~v7 & ~v10;
  assign new_n78_ = ~new_n76_ & ~new_n77_;
  assign new_n79_ = ~v5 & ~new_n78_;
  assign new_n80_ = v5 & new_n77_;
  assign new_n81_ = ~new_n79_ & ~new_n80_;
  assign new_n82_ = v6 & ~new_n81_;
  assign new_n83_ = ~new_n75_ & ~new_n82_;
  assign new_n84_ = ~v25 & ~new_n83_;
  assign new_n85_ = ~v24 & new_n84_;
  assign new_n86_ = ~v23 & new_n85_;
  assign new_n87_ = ~v22 & new_n86_;
  assign new_n88_ = v9 & new_n87_;
  assign new_n89_ = ~v8 & new_n88_;
  assign new_n90_ = v4 & new_n89_;
  assign new_n91_ = v3 & new_n90_;
  assign new_n92_ = v2 & new_n91_;
  assign new_n93_ = v1 & new_n92_;
  assign \v26.0  = ~v0 & new_n93_;
  assign new_n95_ = ~v0 & ~v1;
  assign new_n96_ = ~v2 & new_n95_;
  assign new_n97_ = ~v3 & new_n96_;
  assign new_n98_ = ~v4 & new_n97_;
  assign new_n99_ = ~v5 & new_n98_;
  assign new_n100_ = ~v6 & new_n99_;
  assign new_n101_ = ~v7 & new_n100_;
  assign new_n102_ = ~v8 & new_n101_;
  assign new_n103_ = ~v9 & new_n102_;
  assign new_n104_ = ~v10 & new_n103_;
  assign new_n105_ = ~v22 & new_n104_;
  assign new_n106_ = ~v23 & new_n105_;
  assign new_n107_ = ~v24 & new_n106_;
  assign \v26.1  = ~v25 & new_n107_;
  assign new_n109_ = v9 & ~new_n83_;
  assign new_n110_ = v4 & new_n109_;
  assign new_n111_ = v3 & new_n110_;
  assign new_n112_ = v2 & new_n111_;
  assign new_n113_ = v1 & new_n112_;
  assign new_n114_ = ~v1 & ~v2;
  assign new_n115_ = ~v3 & ~v4;
  assign new_n116_ = new_n114_ & new_n115_;
  assign new_n117_ = ~v5 & ~v6;
  assign new_n118_ = ~v9 & ~v10;
  assign new_n119_ = ~v7 & new_n118_;
  assign new_n120_ = new_n117_ & new_n119_;
  assign new_n121_ = new_n116_ & new_n120_;
  assign new_n122_ = ~new_n113_ & ~new_n121_;
  assign new_n123_ = ~v25 & ~new_n122_;
  assign new_n124_ = ~v24 & new_n123_;
  assign new_n125_ = ~v23 & new_n124_;
  assign new_n126_ = ~v22 & new_n125_;
  assign new_n127_ = ~v8 & new_n126_;
  assign \v26.2  = ~v0 & new_n127_;
  assign new_n129_ = ~v23 & v25;
  assign new_n130_ = v6 & new_n129_;
  assign new_n131_ = ~v5 & new_n130_;
  assign new_n132_ = v3 & new_n131_;
  assign new_n133_ = ~v2 & new_n132_;
  assign new_n134_ = v1 & new_n133_;
  assign new_n135_ = v0 & new_n134_;
  assign new_n136_ = v2 & ~v3;
  assign new_n137_ = new_n95_ & new_n136_;
  assign new_n138_ = v5 & ~v6;
  assign new_n139_ = v23 & ~v25;
  assign new_n140_ = v10 & new_n139_;
  assign new_n141_ = new_n138_ & new_n140_;
  assign new_n142_ = new_n137_ & new_n141_;
  assign new_n143_ = ~new_n135_ & ~new_n142_;
  assign new_n144_ = v7 & ~new_n143_;
  assign new_n145_ = ~v3 & v5;
  assign new_n146_ = v2 & new_n145_;
  assign new_n147_ = new_n95_ & new_n146_;
  assign new_n148_ = ~v6 & ~v7;
  assign new_n149_ = new_n140_ & new_n148_;
  assign new_n150_ = new_n147_ & new_n149_;
  assign new_n151_ = ~new_n144_ & ~new_n150_;
  assign new_n152_ = v9 & ~new_n151_;
  assign new_n153_ = ~v9 & new_n129_;
  assign new_n154_ = v7 & new_n153_;
  assign new_n155_ = v6 & new_n154_;
  assign new_n156_ = ~v5 & new_n155_;
  assign new_n157_ = v3 & new_n156_;
  assign new_n158_ = ~v2 & new_n157_;
  assign new_n159_ = v1 & new_n158_;
  assign new_n160_ = v0 & new_n159_;
  assign new_n161_ = ~new_n152_ & ~new_n160_;
  assign new_n162_ = ~v8 & ~new_n161_;
  assign new_n163_ = v8 & new_n129_;
  assign new_n164_ = v7 & new_n163_;
  assign new_n165_ = v6 & new_n164_;
  assign new_n166_ = ~v5 & new_n165_;
  assign new_n167_ = v3 & new_n166_;
  assign new_n168_ = ~v2 & new_n167_;
  assign new_n169_ = v1 & new_n168_;
  assign new_n170_ = v0 & new_n169_;
  assign new_n171_ = ~new_n162_ & ~new_n170_;
  assign new_n172_ = v4 & ~new_n171_;
  assign new_n173_ = ~v23 & ~v25;
  assign new_n174_ = ~v9 & new_n173_;
  assign new_n175_ = ~v8 & new_n174_;
  assign new_n176_ = v7 & new_n175_;
  assign new_n177_ = v6 & new_n176_;
  assign new_n178_ = v5 & new_n177_;
  assign new_n179_ = ~v4 & new_n178_;
  assign new_n180_ = v3 & new_n179_;
  assign new_n181_ = v2 & new_n180_;
  assign new_n182_ = ~v1 & new_n181_;
  assign new_n183_ = ~v0 & new_n182_;
  assign new_n184_ = ~new_n172_ & ~new_n183_;
  assign new_n185_ = v24 & ~new_n184_;
  assign \v26.3  = ~v22 & new_n185_;
  assign new_n187_ = ~v24 & v25;
  assign new_n188_ = v24 & ~v25;
  assign new_n189_ = ~new_n187_ & ~new_n188_;
  assign new_n190_ = ~v6 & ~new_n189_;
  assign new_n191_ = ~v4 & new_n190_;
  assign new_n192_ = ~v0 & new_n191_;
  assign new_n193_ = v0 & v4;
  assign new_n194_ = ~v24 & ~v25;
  assign new_n195_ = v6 & new_n194_;
  assign new_n196_ = new_n193_ & new_n195_;
  assign new_n197_ = ~new_n192_ & ~new_n196_;
  assign new_n198_ = v2 & ~new_n197_;
  assign new_n199_ = ~v1 & new_n198_;
  assign new_n200_ = v24 & v25;
  assign new_n201_ = ~new_n194_ & ~new_n200_;
  assign new_n202_ = v6 & ~new_n201_;
  assign new_n203_ = v4 & new_n202_;
  assign new_n204_ = ~v2 & new_n203_;
  assign new_n205_ = v1 & new_n204_;
  assign new_n206_ = v0 & new_n205_;
  assign new_n207_ = ~new_n199_ & ~new_n206_;
  assign new_n208_ = v10 & ~new_n207_;
  assign new_n209_ = ~v10 & ~new_n201_;
  assign new_n210_ = v6 & new_n209_;
  assign new_n211_ = v4 & new_n210_;
  assign new_n212_ = ~v2 & new_n211_;
  assign new_n213_ = v1 & new_n212_;
  assign new_n214_ = v0 & new_n213_;
  assign new_n215_ = ~new_n208_ & ~new_n214_;
  assign new_n216_ = ~v8 & ~new_n215_;
  assign new_n217_ = v8 & ~new_n201_;
  assign new_n218_ = v6 & new_n217_;
  assign new_n219_ = v4 & new_n218_;
  assign new_n220_ = ~v2 & new_n219_;
  assign new_n221_ = v1 & new_n220_;
  assign new_n222_ = v0 & new_n221_;
  assign new_n223_ = ~new_n216_ & ~new_n222_;
  assign new_n224_ = v3 & ~new_n223_;
  assign new_n225_ = ~v10 & v24;
  assign new_n226_ = v8 & new_n225_;
  assign new_n227_ = v6 & new_n226_;
  assign new_n228_ = ~v4 & new_n227_;
  assign new_n229_ = ~v3 & new_n228_;
  assign new_n230_ = ~v2 & new_n229_;
  assign new_n231_ = v1 & new_n230_;
  assign new_n232_ = v0 & new_n231_;
  assign new_n233_ = ~new_n224_ & ~new_n232_;
  assign new_n234_ = ~v5 & ~new_n233_;
  assign new_n235_ = ~v0 & new_n114_;
  assign new_n236_ = ~v4 & v5;
  assign new_n237_ = ~v3 & new_n236_;
  assign new_n238_ = new_n235_ & new_n237_;
  assign new_n239_ = v8 & ~v10;
  assign new_n240_ = ~v6 & new_n239_;
  assign new_n241_ = ~v19 & new_n187_;
  assign new_n242_ = new_n240_ & new_n241_;
  assign new_n243_ = new_n238_ & new_n242_;
  assign new_n244_ = ~new_n234_ & ~new_n243_;
  assign new_n245_ = ~v3 & v24;
  assign new_n246_ = v1 & new_n245_;
  assign new_n247_ = v3 & ~v24;
  assign new_n248_ = ~v1 & new_n247_;
  assign new_n249_ = ~new_n246_ & ~new_n248_;
  assign new_n250_ = ~v10 & ~new_n249_;
  assign new_n251_ = ~v9 & new_n250_;
  assign new_n252_ = ~v4 & new_n251_;
  assign new_n253_ = v0 & new_n252_;
  assign new_n254_ = ~v0 & v1;
  assign new_n255_ = v3 & v4;
  assign new_n256_ = new_n254_ & new_n255_;
  assign new_n257_ = ~v8 & v9;
  assign new_n258_ = v10 & v24;
  assign new_n259_ = new_n257_ & new_n258_;
  assign new_n260_ = new_n256_ & new_n259_;
  assign new_n261_ = ~new_n253_ & ~new_n260_;
  assign new_n262_ = v6 & ~new_n261_;
  assign new_n263_ = v9 & v24;
  assign new_n264_ = ~v8 & new_n263_;
  assign new_n265_ = ~v6 & new_n264_;
  assign new_n266_ = v4 & new_n265_;
  assign new_n267_ = v3 & new_n266_;
  assign new_n268_ = v1 & new_n267_;
  assign new_n269_ = ~v0 & new_n268_;
  assign new_n270_ = ~new_n262_ & ~new_n269_;
  assign new_n271_ = v2 & ~new_n270_;
  assign new_n272_ = v3 & v8;
  assign new_n273_ = ~v3 & ~v8;
  assign new_n274_ = ~new_n272_ & ~new_n273_;
  assign new_n275_ = ~v24 & ~new_n274_;
  assign new_n276_ = ~v1 & new_n275_;
  assign new_n277_ = v1 & ~v3;
  assign new_n278_ = ~v8 & v24;
  assign new_n279_ = new_n277_ & new_n278_;
  assign new_n280_ = ~new_n276_ & ~new_n279_;
  assign new_n281_ = ~v10 & ~new_n280_;
  assign new_n282_ = ~v9 & new_n281_;
  assign new_n283_ = v6 & new_n282_;
  assign new_n284_ = ~v4 & new_n283_;
  assign new_n285_ = ~v2 & new_n284_;
  assign new_n286_ = v0 & new_n285_;
  assign new_n287_ = ~new_n271_ & ~new_n286_;
  assign new_n288_ = ~v5 & ~new_n287_;
  assign new_n289_ = v0 & v1;
  assign new_n290_ = v2 & new_n115_;
  assign new_n291_ = new_n289_ & new_n290_;
  assign new_n292_ = v6 & v8;
  assign new_n293_ = v5 & new_n292_;
  assign new_n294_ = v9 & new_n225_;
  assign new_n295_ = new_n293_ & new_n294_;
  assign new_n296_ = new_n291_ & new_n295_;
  assign new_n297_ = ~new_n288_ & ~new_n296_;
  assign new_n298_ = ~v9 & v10;
  assign new_n299_ = v8 & new_n298_;
  assign new_n300_ = v9 & ~v10;
  assign new_n301_ = ~v8 & new_n300_;
  assign new_n302_ = ~new_n299_ & ~new_n301_;
  assign new_n303_ = v1 & ~new_n302_;
  assign new_n304_ = ~v1 & ~v8;
  assign new_n305_ = new_n298_ & new_n304_;
  assign new_n306_ = ~new_n303_ & ~new_n305_;
  assign new_n307_ = v25 & ~new_n306_;
  assign new_n308_ = ~v2 & new_n307_;
  assign new_n309_ = ~v0 & new_n308_;
  assign new_n310_ = v8 & v9;
  assign new_n311_ = ~v8 & new_n118_;
  assign new_n312_ = ~new_n310_ & ~new_n311_;
  assign new_n313_ = ~v25 & ~new_n312_;
  assign new_n314_ = v2 & new_n313_;
  assign new_n315_ = ~v1 & new_n314_;
  assign new_n316_ = v0 & new_n315_;
  assign new_n317_ = ~new_n309_ & ~new_n316_;
  assign new_n318_ = v4 & ~new_n317_;
  assign new_n319_ = ~v2 & ~v4;
  assign new_n320_ = new_n95_ & new_n319_;
  assign new_n321_ = v8 & ~v9;
  assign new_n322_ = ~v10 & ~v25;
  assign new_n323_ = new_n321_ & new_n322_;
  assign new_n324_ = new_n320_ & new_n323_;
  assign new_n325_ = ~new_n318_ & ~new_n324_;
  assign new_n326_ = ~v24 & ~new_n325_;
  assign new_n327_ = ~v8 & v25;
  assign new_n328_ = v8 & ~v25;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign new_n330_ = v2 & ~new_n329_;
  assign new_n331_ = ~v2 & new_n328_;
  assign new_n332_ = ~new_n330_ & ~new_n331_;
  assign new_n333_ = ~v1 & ~new_n332_;
  assign new_n334_ = v1 & v2;
  assign new_n335_ = new_n327_ & new_n334_;
  assign new_n336_ = ~new_n333_ & ~new_n335_;
  assign new_n337_ = v24 & ~new_n336_;
  assign new_n338_ = ~v10 & new_n337_;
  assign new_n339_ = ~v9 & new_n338_;
  assign new_n340_ = ~v4 & new_n339_;
  assign new_n341_ = v0 & new_n340_;
  assign new_n342_ = ~new_n326_ & ~new_n341_;
  assign new_n343_ = v6 & ~new_n342_;
  assign new_n344_ = ~v4 & v8;
  assign new_n345_ = v2 & new_n344_;
  assign new_n346_ = ~v2 & v4;
  assign new_n347_ = ~v8 & ~v10;
  assign new_n348_ = new_n346_ & new_n347_;
  assign new_n349_ = ~new_n345_ & ~new_n348_;
  assign new_n350_ = ~v25 & ~new_n349_;
  assign new_n351_ = ~v24 & new_n350_;
  assign new_n352_ = ~v9 & new_n351_;
  assign new_n353_ = ~v6 & new_n352_;
  assign new_n354_ = ~v1 & new_n353_;
  assign new_n355_ = ~v0 & new_n354_;
  assign new_n356_ = ~new_n343_ & ~new_n355_;
  assign new_n357_ = v3 & ~new_n356_;
  assign new_n358_ = v2 & ~v6;
  assign new_n359_ = ~v8 & v10;
  assign new_n360_ = new_n358_ & new_n359_;
  assign new_n361_ = ~v2 & v6;
  assign new_n362_ = new_n239_ & new_n361_;
  assign new_n363_ = ~new_n360_ & ~new_n362_;
  assign new_n364_ = ~v24 & ~new_n363_;
  assign new_n365_ = v9 & new_n364_;
  assign new_n366_ = ~v0 & new_n365_;
  assign new_n367_ = v0 & new_n361_;
  assign new_n368_ = ~v8 & ~v9;
  assign new_n369_ = new_n225_ & new_n368_;
  assign new_n370_ = new_n367_ & new_n369_;
  assign new_n371_ = ~new_n366_ & ~new_n370_;
  assign new_n372_ = v25 & ~new_n371_;
  assign new_n373_ = ~v4 & new_n372_;
  assign new_n374_ = ~v3 & new_n373_;
  assign new_n375_ = ~v1 & new_n374_;
  assign new_n376_ = ~new_n357_ & ~new_n375_;
  assign new_n377_ = ~v5 & ~new_n376_;
  assign new_n378_ = ~v9 & ~new_n189_;
  assign new_n379_ = v8 & new_n378_;
  assign new_n380_ = v6 & new_n379_;
  assign new_n381_ = v3 & new_n380_;
  assign new_n382_ = ~v6 & ~v8;
  assign new_n383_ = ~v3 & new_n382_;
  assign new_n384_ = v9 & new_n200_;
  assign new_n385_ = new_n383_ & new_n384_;
  assign new_n386_ = ~new_n381_ & ~new_n385_;
  assign new_n387_ = v10 & ~new_n386_;
  assign new_n388_ = v5 & new_n387_;
  assign new_n389_ = v4 & new_n388_;
  assign new_n390_ = v2 & new_n389_;
  assign new_n391_ = ~v1 & new_n390_;
  assign new_n392_ = ~v0 & new_n391_;
  assign new_n393_ = ~new_n377_ & ~new_n392_;
  assign new_n394_ = new_n297_ & new_n393_;
  assign new_n395_ = new_n244_ & new_n394_;
  assign new_n396_ = v7 & ~new_n395_;
  assign new_n397_ = v2 & v4;
  assign new_n398_ = v9 & v10;
  assign new_n399_ = v5 & new_n398_;
  assign new_n400_ = new_n397_ & new_n399_;
  assign new_n401_ = ~v5 & new_n118_;
  assign new_n402_ = new_n319_ & new_n401_;
  assign new_n403_ = ~new_n400_ & ~new_n402_;
  assign new_n404_ = ~v3 & ~new_n403_;
  assign new_n405_ = ~v1 & new_n404_;
  assign new_n406_ = v4 & v9;
  assign new_n407_ = v3 & new_n406_;
  assign new_n408_ = v2 & new_n407_;
  assign new_n409_ = v1 & new_n408_;
  assign new_n410_ = ~new_n405_ & ~new_n409_;
  assign new_n411_ = ~v6 & ~new_n410_;
  assign new_n412_ = v6 & new_n300_;
  assign new_n413_ = v4 & new_n412_;
  assign new_n414_ = v3 & new_n413_;
  assign new_n415_ = v2 & new_n414_;
  assign new_n416_ = v1 & new_n415_;
  assign new_n417_ = ~new_n411_ & ~new_n416_;
  assign new_n418_ = ~v1 & v2;
  assign new_n419_ = v4 & v5;
  assign new_n420_ = ~v3 & new_n419_;
  assign new_n421_ = new_n418_ & new_n420_;
  assign new_n422_ = v6 & ~v9;
  assign new_n423_ = ~v19 & ~v25;
  assign new_n424_ = ~v10 & new_n423_;
  assign new_n425_ = new_n422_ & new_n424_;
  assign new_n426_ = new_n421_ & new_n425_;
  assign new_n427_ = new_n417_ & ~new_n426_;
  assign new_n428_ = v24 & ~new_n427_;
  assign new_n429_ = ~v3 & v9;
  assign new_n430_ = ~v10 & v25;
  assign new_n431_ = new_n429_ & new_n430_;
  assign new_n432_ = v3 & ~v9;
  assign new_n433_ = v10 & ~v25;
  assign new_n434_ = new_n432_ & new_n433_;
  assign new_n435_ = ~new_n431_ & ~new_n434_;
  assign new_n436_ = v6 & ~new_n435_;
  assign new_n437_ = v4 & new_n436_;
  assign new_n438_ = v1 & new_n437_;
  assign new_n439_ = v3 & ~v4;
  assign new_n440_ = ~v1 & new_n439_;
  assign new_n441_ = ~v6 & v9;
  assign new_n442_ = new_n322_ & new_n441_;
  assign new_n443_ = new_n440_ & new_n442_;
  assign new_n444_ = ~new_n438_ & ~new_n443_;
  assign new_n445_ = ~v24 & ~new_n444_;
  assign new_n446_ = v5 & new_n445_;
  assign new_n447_ = ~v2 & new_n446_;
  assign new_n448_ = ~new_n428_ & ~new_n447_;
  assign new_n449_ = ~v8 & ~new_n448_;
  assign new_n450_ = v4 & ~v5;
  assign new_n451_ = v3 & new_n450_;
  assign new_n452_ = new_n114_ & new_n451_;
  assign new_n453_ = v6 & new_n321_;
  assign new_n454_ = ~v10 & new_n194_;
  assign new_n455_ = new_n453_ & new_n454_;
  assign new_n456_ = new_n452_ & new_n455_;
  assign new_n457_ = ~new_n449_ & ~new_n456_;
  assign new_n458_ = ~v0 & ~new_n457_;
  assign new_n459_ = v3 & new_n188_;
  assign new_n460_ = ~v1 & new_n459_;
  assign new_n461_ = new_n249_ & ~new_n460_;
  assign new_n462_ = ~v10 & ~new_n461_;
  assign new_n463_ = v9 & new_n462_;
  assign new_n464_ = v8 & new_n463_;
  assign new_n465_ = v6 & new_n464_;
  assign new_n466_ = ~v5 & new_n465_;
  assign new_n467_ = ~v4 & new_n466_;
  assign new_n468_ = v0 & new_n467_;
  assign new_n469_ = ~new_n458_ & ~new_n468_;
  assign new_n470_ = ~v7 & ~new_n469_;
  assign new_n471_ = ~new_n396_ & ~new_n470_;
  assign new_n472_ = ~v23 & ~new_n471_;
  assign new_n473_ = ~v6 & new_n398_;
  assign new_n474_ = v5 & new_n473_;
  assign new_n475_ = v4 & new_n474_;
  assign new_n476_ = v2 & new_n475_;
  assign new_n477_ = ~v0 & new_n476_;
  assign new_n478_ = v0 & ~v2;
  assign new_n479_ = ~v4 & ~v5;
  assign new_n480_ = new_n478_ & new_n479_;
  assign new_n481_ = new_n225_ & new_n422_;
  assign new_n482_ = new_n480_ & new_n481_;
  assign new_n483_ = ~new_n477_ & ~new_n482_;
  assign new_n484_ = ~v1 & ~new_n483_;
  assign new_n485_ = ~v9 & new_n225_;
  assign new_n486_ = v6 & new_n485_;
  assign new_n487_ = ~v5 & new_n486_;
  assign new_n488_ = ~v4 & new_n487_;
  assign new_n489_ = v1 & new_n488_;
  assign new_n490_ = v0 & new_n489_;
  assign new_n491_ = ~new_n484_ & ~new_n490_;
  assign new_n492_ = v7 & ~new_n491_;
  assign new_n493_ = v4 & new_n399_;
  assign new_n494_ = v2 & new_n493_;
  assign new_n495_ = ~v2 & new_n479_;
  assign new_n496_ = ~v10 & ~v24;
  assign new_n497_ = ~v9 & new_n496_;
  assign new_n498_ = new_n495_ & new_n497_;
  assign new_n499_ = ~new_n494_ & ~new_n498_;
  assign new_n500_ = ~v7 & ~new_n499_;
  assign new_n501_ = ~v6 & new_n500_;
  assign new_n502_ = ~v1 & new_n501_;
  assign new_n503_ = ~v0 & new_n502_;
  assign new_n504_ = ~new_n492_ & ~new_n503_;
  assign new_n505_ = ~v25 & ~new_n504_;
  assign new_n506_ = ~v1 & ~new_n114_;
  assign new_n507_ = v25 & ~new_n506_;
  assign new_n508_ = ~v24 & new_n507_;
  assign new_n509_ = ~v10 & new_n508_;
  assign new_n510_ = ~v9 & new_n509_;
  assign new_n511_ = v7 & new_n510_;
  assign new_n512_ = v6 & new_n511_;
  assign new_n513_ = ~v5 & new_n512_;
  assign new_n514_ = ~v4 & new_n513_;
  assign new_n515_ = v0 & new_n514_;
  assign new_n516_ = ~new_n505_ & ~new_n515_;
  assign new_n517_ = ~v3 & ~new_n516_;
  assign new_n518_ = ~v10 & ~new_n189_;
  assign new_n519_ = ~v9 & new_n518_;
  assign new_n520_ = v7 & new_n519_;
  assign new_n521_ = v6 & new_n520_;
  assign new_n522_ = ~v5 & new_n521_;
  assign new_n523_ = ~v4 & new_n522_;
  assign new_n524_ = v3 & new_n523_;
  assign new_n525_ = v2 & new_n524_;
  assign new_n526_ = v0 & new_n525_;
  assign new_n527_ = ~new_n517_ & ~new_n526_;
  assign new_n528_ = v23 & ~new_n527_;
  assign new_n529_ = ~v8 & new_n528_;
  assign new_n530_ = ~new_n472_ & ~new_n529_;
  assign \v26.4  = ~v22 & ~new_n530_;
  assign new_n532_ = ~v0 & new_n358_;
  assign new_n533_ = v6 & v7;
  assign new_n534_ = new_n478_ & new_n533_;
  assign new_n535_ = ~new_n532_ & ~new_n534_;
  assign new_n536_ = ~v5 & ~new_n535_;
  assign new_n537_ = ~v0 & v2;
  assign new_n538_ = v5 & new_n148_;
  assign new_n539_ = new_n537_ & new_n538_;
  assign new_n540_ = ~new_n536_ & ~new_n539_;
  assign new_n541_ = v2 & new_n82_;
  assign new_n542_ = ~v0 & new_n541_;
  assign new_n543_ = new_n540_ & ~new_n542_;
  assign new_n544_ = v1 & ~new_n543_;
  assign new_n545_ = ~v0 & new_n418_;
  assign new_n546_ = v5 & v6;
  assign new_n547_ = ~v7 & v10;
  assign new_n548_ = new_n546_ & new_n547_;
  assign new_n549_ = new_n545_ & new_n548_;
  assign new_n550_ = ~new_n544_ & ~new_n549_;
  assign new_n551_ = v3 & ~new_n550_;
  assign new_n552_ = ~v6 & v10;
  assign new_n553_ = v5 & new_n552_;
  assign new_n554_ = ~v3 & new_n553_;
  assign new_n555_ = v2 & new_n554_;
  assign new_n556_ = ~v1 & new_n555_;
  assign new_n557_ = ~v0 & new_n556_;
  assign new_n558_ = ~new_n551_ & ~new_n557_;
  assign new_n559_ = ~v24 & ~new_n558_;
  assign new_n560_ = ~v23 & new_n559_;
  assign new_n561_ = v23 & v24;
  assign new_n562_ = v10 & new_n561_;
  assign new_n563_ = ~v6 & new_n562_;
  assign new_n564_ = v5 & new_n563_;
  assign new_n565_ = ~v3 & new_n564_;
  assign new_n566_ = v2 & new_n565_;
  assign new_n567_ = ~v1 & new_n566_;
  assign new_n568_ = ~v0 & new_n567_;
  assign new_n569_ = ~new_n560_ & ~new_n568_;
  assign new_n570_ = ~v25 & ~new_n569_;
  assign new_n571_ = ~v5 & v7;
  assign new_n572_ = v3 & new_n571_;
  assign new_n573_ = v0 & new_n572_;
  assign new_n574_ = ~v0 & new_n145_;
  assign new_n575_ = ~v7 & new_n496_;
  assign new_n576_ = new_n574_ & new_n575_;
  assign new_n577_ = ~new_n573_ & ~new_n576_;
  assign new_n578_ = v25 & ~new_n577_;
  assign new_n579_ = ~v23 & new_n578_;
  assign new_n580_ = v6 & new_n579_;
  assign new_n581_ = ~v2 & new_n580_;
  assign new_n582_ = v1 & new_n581_;
  assign new_n583_ = ~new_n570_ & ~new_n582_;
  assign new_n584_ = v9 & ~new_n583_;
  assign new_n585_ = ~v5 & v6;
  assign new_n586_ = v3 & new_n585_;
  assign new_n587_ = v1 & new_n586_;
  assign new_n588_ = v0 & new_n587_;
  assign new_n589_ = ~v1 & ~v3;
  assign new_n590_ = ~v0 & new_n589_;
  assign new_n591_ = new_n553_ & new_n590_;
  assign new_n592_ = ~new_n588_ & ~new_n591_;
  assign new_n593_ = ~v1 & v3;
  assign new_n594_ = ~v0 & new_n593_;
  assign new_n595_ = new_n117_ & new_n322_;
  assign new_n596_ = new_n594_ & new_n595_;
  assign new_n597_ = new_n592_ & ~new_n596_;
  assign new_n598_ = ~v24 & ~new_n597_;
  assign new_n599_ = v6 & new_n200_;
  assign new_n600_ = ~v5 & new_n599_;
  assign new_n601_ = v3 & new_n600_;
  assign new_n602_ = v1 & new_n601_;
  assign new_n603_ = v0 & new_n602_;
  assign new_n604_ = ~new_n598_ & ~new_n603_;
  assign new_n605_ = ~v23 & ~new_n604_;
  assign new_n606_ = ~v9 & new_n605_;
  assign new_n607_ = v7 & new_n606_;
  assign new_n608_ = ~v2 & new_n607_;
  assign new_n609_ = ~new_n584_ & ~new_n608_;
  assign new_n610_ = ~v8 & ~new_n609_;
  assign new_n611_ = v3 & new_n546_;
  assign new_n612_ = ~v9 & v25;
  assign new_n613_ = v7 & new_n612_;
  assign new_n614_ = new_n611_ & new_n613_;
  assign new_n615_ = ~v3 & new_n117_;
  assign new_n616_ = v9 & ~v25;
  assign new_n617_ = ~v7 & new_n616_;
  assign new_n618_ = new_n615_ & new_n617_;
  assign new_n619_ = ~new_n614_ & ~new_n618_;
  assign new_n620_ = v2 & ~new_n619_;
  assign new_n621_ = ~v1 & new_n620_;
  assign new_n622_ = ~v0 & new_n621_;
  assign new_n623_ = ~v5 & new_n533_;
  assign new_n624_ = v3 & new_n623_;
  assign new_n625_ = ~v2 & new_n624_;
  assign new_n626_ = v1 & new_n625_;
  assign new_n627_ = v0 & new_n626_;
  assign new_n628_ = ~new_n622_ & ~new_n627_;
  assign new_n629_ = v10 & ~new_n628_;
  assign new_n630_ = v1 & v7;
  assign new_n631_ = v0 & new_n630_;
  assign new_n632_ = ~v9 & ~v25;
  assign new_n633_ = ~v7 & new_n632_;
  assign new_n634_ = new_n95_ & new_n633_;
  assign new_n635_ = ~new_n631_ & ~new_n634_;
  assign new_n636_ = ~v10 & ~new_n635_;
  assign new_n637_ = v6 & new_n636_;
  assign new_n638_ = ~v5 & new_n637_;
  assign new_n639_ = v3 & new_n638_;
  assign new_n640_ = ~v2 & new_n639_;
  assign new_n641_ = ~new_n629_ & ~new_n640_;
  assign new_n642_ = ~v24 & ~new_n641_;
  assign new_n643_ = v7 & new_n200_;
  assign new_n644_ = v6 & new_n643_;
  assign new_n645_ = ~v5 & new_n644_;
  assign new_n646_ = v3 & new_n645_;
  assign new_n647_ = ~v2 & new_n646_;
  assign new_n648_ = v1 & new_n647_;
  assign new_n649_ = v0 & new_n648_;
  assign new_n650_ = ~new_n642_ & ~new_n649_;
  assign new_n651_ = ~v23 & ~new_n650_;
  assign new_n652_ = v8 & new_n651_;
  assign new_n653_ = ~new_n610_ & ~new_n652_;
  assign new_n654_ = v4 & ~new_n653_;
  assign new_n655_ = ~v0 & ~new_n363_;
  assign new_n656_ = ~v2 & v8;
  assign new_n657_ = ~v2 & ~new_n656_;
  assign new_n658_ = ~v10 & ~new_n657_;
  assign new_n659_ = v6 & new_n658_;
  assign new_n660_ = v0 & new_n659_;
  assign new_n661_ = ~new_n655_ & ~new_n660_;
  assign new_n662_ = ~v25 & ~new_n661_;
  assign new_n663_ = ~v24 & new_n662_;
  assign new_n664_ = new_n200_ & new_n359_;
  assign new_n665_ = new_n532_ & new_n664_;
  assign new_n666_ = ~new_n663_ & ~new_n665_;
  assign new_n667_ = ~v9 & ~new_n666_;
  assign new_n668_ = v10 & ~new_n201_;
  assign new_n669_ = v9 & new_n668_;
  assign new_n670_ = ~v8 & new_n669_;
  assign new_n671_ = ~v6 & new_n670_;
  assign new_n672_ = v2 & new_n671_;
  assign new_n673_ = ~v0 & new_n672_;
  assign new_n674_ = ~new_n667_ & ~new_n673_;
  assign new_n675_ = ~v5 & ~new_n674_;
  assign new_n676_ = ~v9 & new_n188_;
  assign new_n677_ = ~v8 & new_n676_;
  assign new_n678_ = v6 & new_n677_;
  assign new_n679_ = v5 & new_n678_;
  assign new_n680_ = v2 & new_n679_;
  assign new_n681_ = ~v0 & new_n680_;
  assign new_n682_ = ~new_n675_ & ~new_n681_;
  assign new_n683_ = v7 & ~new_n682_;
  assign new_n684_ = v9 & new_n454_;
  assign new_n685_ = v8 & new_n684_;
  assign new_n686_ = ~v7 & new_n685_;
  assign new_n687_ = v6 & new_n686_;
  assign new_n688_ = ~v5 & new_n687_;
  assign new_n689_ = v0 & new_n688_;
  assign new_n690_ = ~new_n683_ & ~new_n689_;
  assign new_n691_ = v3 & ~new_n690_;
  assign new_n692_ = new_n148_ & new_n430_;
  assign new_n693_ = new_n433_ & new_n533_;
  assign new_n694_ = ~new_n692_ & ~new_n693_;
  assign new_n695_ = ~v0 & ~new_n694_;
  assign new_n696_ = v0 & v6;
  assign new_n697_ = v7 & new_n322_;
  assign new_n698_ = new_n696_ & new_n697_;
  assign new_n699_ = ~new_n695_ & ~new_n698_;
  assign new_n700_ = ~v24 & ~new_n699_;
  assign new_n701_ = ~v9 & new_n700_;
  assign new_n702_ = ~v8 & new_n701_;
  assign new_n703_ = ~v5 & new_n702_;
  assign new_n704_ = ~v3 & new_n703_;
  assign new_n705_ = ~v2 & new_n704_;
  assign new_n706_ = ~new_n691_ & ~new_n705_;
  assign new_n707_ = ~v23 & ~new_n706_;
  assign new_n708_ = ~v4 & new_n707_;
  assign new_n709_ = ~v1 & new_n708_;
  assign new_n710_ = ~new_n654_ & ~new_n709_;
  assign \v26.5  = ~v22 & ~new_n710_;
  assign new_n712_ = v2 & v3;
  assign new_n713_ = ~v2 & ~v3;
  assign new_n714_ = ~new_n712_ & ~new_n713_;
  assign new_n715_ = v1 & new_n136_;
  assign new_n716_ = new_n714_ & ~new_n715_;
  assign new_n717_ = ~v24 & ~new_n716_;
  assign new_n718_ = v23 & new_n717_;
  assign new_n719_ = ~v10 & new_n718_;
  assign new_n720_ = ~v9 & new_n719_;
  assign new_n721_ = v6 & new_n720_;
  assign new_n722_ = ~v5 & new_n721_;
  assign new_n723_ = ~v4 & new_n722_;
  assign new_n724_ = v0 & new_n723_;
  assign new_n725_ = ~v3 & v4;
  assign new_n726_ = v2 & new_n725_;
  assign new_n727_ = new_n95_ & new_n726_;
  assign new_n728_ = v5 & new_n441_;
  assign new_n729_ = ~v23 & v24;
  assign new_n730_ = v10 & new_n729_;
  assign new_n731_ = new_n728_ & new_n730_;
  assign new_n732_ = new_n727_ & new_n731_;
  assign new_n733_ = ~new_n724_ & ~new_n732_;
  assign new_n734_ = ~v25 & ~new_n733_;
  assign new_n735_ = ~v22 & new_n734_;
  assign new_n736_ = ~v8 & new_n735_;
  assign \v26.6  = v7 & new_n736_;
  assign new_n738_ = v23 & ~v24;
  assign new_n739_ = ~v5 & new_n738_;
  assign new_n740_ = v0 & new_n739_;
  assign new_n741_ = v5 & new_n729_;
  assign new_n742_ = new_n95_ & new_n741_;
  assign new_n743_ = ~new_n740_ & ~new_n742_;
  assign new_n744_ = ~v10 & ~new_n743_;
  assign new_n745_ = ~v1 & v5;
  assign new_n746_ = ~v0 & new_n745_;
  assign new_n747_ = new_n730_ & new_n746_;
  assign new_n748_ = ~new_n744_ & ~new_n747_;
  assign new_n749_ = v3 & ~new_n748_;
  assign new_n750_ = v0 & new_n277_;
  assign new_n751_ = ~v5 & ~v10;
  assign new_n752_ = new_n738_ & new_n751_;
  assign new_n753_ = new_n750_ & new_n752_;
  assign new_n754_ = ~new_n749_ & ~new_n753_;
  assign new_n755_ = v2 & ~new_n754_;
  assign new_n756_ = ~v10 & new_n738_;
  assign new_n757_ = ~v5 & new_n756_;
  assign new_n758_ = ~v3 & new_n757_;
  assign new_n759_ = ~v2 & new_n758_;
  assign new_n760_ = v0 & new_n759_;
  assign new_n761_ = ~new_n755_ & ~new_n760_;
  assign new_n762_ = ~v25 & ~new_n761_;
  assign new_n763_ = ~v8 & new_n762_;
  assign new_n764_ = ~v4 & new_n763_;
  assign new_n765_ = ~v2 & new_n255_;
  assign new_n766_ = new_n289_ & new_n765_;
  assign new_n767_ = v8 & v10;
  assign new_n768_ = ~v5 & new_n767_;
  assign new_n769_ = ~v23 & new_n187_;
  assign new_n770_ = new_n768_ & new_n769_;
  assign new_n771_ = new_n766_ & new_n770_;
  assign new_n772_ = ~new_n764_ & ~new_n771_;
  assign new_n773_ = ~v22 & ~new_n772_;
  assign new_n774_ = ~v9 & new_n773_;
  assign new_n775_ = v7 & new_n774_;
  assign \v26.7  = v6 & new_n775_;
  assign new_n777_ = v3 & new_n292_;
  assign new_n778_ = ~v9 & new_n187_;
  assign new_n779_ = new_n777_ & new_n778_;
  assign new_n780_ = v9 & new_n188_;
  assign new_n781_ = new_n383_ & new_n780_;
  assign new_n782_ = ~new_n779_ & ~new_n781_;
  assign new_n783_ = ~v23 & ~new_n782_;
  assign new_n784_ = v10 & new_n783_;
  assign new_n785_ = v5 & new_n784_;
  assign new_n786_ = v4 & new_n785_;
  assign new_n787_ = ~v0 & new_n786_;
  assign new_n788_ = v0 & v3;
  assign new_n789_ = ~v4 & new_n585_;
  assign new_n790_ = new_n788_ & new_n789_;
  assign new_n791_ = v23 & new_n194_;
  assign new_n792_ = new_n311_ & new_n791_;
  assign new_n793_ = new_n790_ & new_n792_;
  assign new_n794_ = ~new_n787_ & ~new_n793_;
  assign new_n795_ = ~v1 & ~new_n794_;
  assign new_n796_ = ~v10 & new_n791_;
  assign new_n797_ = ~v9 & new_n796_;
  assign new_n798_ = ~v8 & new_n797_;
  assign new_n799_ = v6 & new_n798_;
  assign new_n800_ = ~v5 & new_n799_;
  assign new_n801_ = ~v4 & new_n800_;
  assign new_n802_ = v1 & new_n801_;
  assign new_n803_ = v0 & new_n802_;
  assign new_n804_ = ~new_n795_ & ~new_n803_;
  assign new_n805_ = v2 & ~new_n804_;
  assign new_n806_ = new_n163_ & new_n255_;
  assign new_n807_ = ~v8 & new_n139_;
  assign new_n808_ = new_n115_ & new_n807_;
  assign new_n809_ = ~new_n806_ & ~new_n808_;
  assign new_n810_ = v1 & ~new_n809_;
  assign new_n811_ = ~v1 & new_n115_;
  assign new_n812_ = new_n807_ & new_n811_;
  assign new_n813_ = ~new_n810_ & ~new_n812_;
  assign new_n814_ = ~v24 & ~new_n813_;
  assign new_n815_ = ~v10 & new_n814_;
  assign new_n816_ = ~v9 & new_n815_;
  assign new_n817_ = v6 & new_n816_;
  assign new_n818_ = ~v5 & new_n817_;
  assign new_n819_ = ~v2 & new_n818_;
  assign new_n820_ = v0 & new_n819_;
  assign new_n821_ = ~new_n805_ & ~new_n820_;
  assign new_n822_ = ~v22 & ~new_n821_;
  assign \v26.8  = v7 & new_n822_;
  assign new_n824_ = v1 & v4;
  assign new_n825_ = ~v4 & ~v9;
  assign new_n826_ = ~v1 & new_n825_;
  assign new_n827_ = ~new_n824_ & ~new_n826_;
  assign new_n828_ = v7 & ~new_n827_;
  assign new_n829_ = ~v1 & ~v4;
  assign new_n830_ = ~v7 & v9;
  assign new_n831_ = new_n829_ & new_n830_;
  assign new_n832_ = ~new_n828_ & ~new_n831_;
  assign new_n833_ = ~v2 & ~new_n832_;
  assign new_n834_ = v7 & ~v9;
  assign new_n835_ = ~new_n830_ & ~new_n834_;
  assign new_n836_ = ~v4 & ~new_n835_;
  assign new_n837_ = v2 & new_n836_;
  assign new_n838_ = ~v1 & new_n837_;
  assign new_n839_ = ~new_n833_ & ~new_n838_;
  assign new_n840_ = v8 & ~new_n839_;
  assign new_n841_ = v1 & new_n346_;
  assign new_n842_ = new_n418_ & new_n825_;
  assign new_n843_ = ~new_n841_ & ~new_n842_;
  assign new_n844_ = ~v8 & ~new_n843_;
  assign new_n845_ = v7 & new_n844_;
  assign new_n846_ = ~new_n840_ & ~new_n845_;
  assign new_n847_ = ~v10 & ~new_n846_;
  assign new_n848_ = v4 & new_n76_;
  assign new_n849_ = ~v2 & new_n848_;
  assign new_n850_ = v1 & new_n849_;
  assign new_n851_ = ~new_n847_ & ~new_n850_;
  assign new_n852_ = ~v25 & ~new_n851_;
  assign new_n853_ = v1 & ~v2;
  assign new_n854_ = v4 & v7;
  assign new_n855_ = new_n853_ & new_n854_;
  assign new_n856_ = v10 & v25;
  assign new_n857_ = new_n310_ & new_n856_;
  assign new_n858_ = new_n855_ & new_n857_;
  assign new_n859_ = ~new_n852_ & ~new_n858_;
  assign new_n860_ = ~v24 & ~new_n859_;
  assign new_n861_ = v4 & new_n643_;
  assign new_n862_ = ~v2 & new_n861_;
  assign new_n863_ = v1 & new_n862_;
  assign new_n864_ = ~new_n860_ & ~new_n863_;
  assign new_n865_ = ~v23 & ~new_n864_;
  assign new_n866_ = v7 & new_n798_;
  assign new_n867_ = ~v4 & new_n866_;
  assign new_n868_ = v2 & new_n867_;
  assign new_n869_ = ~new_n865_ & ~new_n868_;
  assign new_n870_ = v0 & ~new_n869_;
  assign new_n871_ = v9 & ~new_n78_;
  assign new_n872_ = ~v8 & new_n871_;
  assign new_n873_ = v2 & new_n872_;
  assign new_n874_ = v1 & new_n873_;
  assign new_n875_ = ~v2 & ~v7;
  assign new_n876_ = ~v1 & new_n875_;
  assign new_n877_ = v8 & new_n118_;
  assign new_n878_ = new_n876_ & new_n877_;
  assign new_n879_ = ~new_n874_ & ~new_n878_;
  assign new_n880_ = v4 & ~new_n879_;
  assign new_n881_ = ~v1 & new_n319_;
  assign new_n882_ = v7 & v8;
  assign new_n883_ = new_n118_ & new_n882_;
  assign new_n884_ = new_n881_ & new_n883_;
  assign new_n885_ = ~new_n880_ & ~new_n884_;
  assign new_n886_ = ~v25 & ~new_n885_;
  assign new_n887_ = ~v24 & new_n886_;
  assign new_n888_ = ~v23 & new_n887_;
  assign new_n889_ = ~v0 & new_n888_;
  assign new_n890_ = ~new_n870_ & ~new_n889_;
  assign new_n891_ = v3 & ~new_n890_;
  assign new_n892_ = v23 & ~new_n506_;
  assign new_n893_ = ~v2 & ~v23;
  assign new_n894_ = ~v1 & new_n893_;
  assign new_n895_ = ~new_n892_ & ~new_n894_;
  assign new_n896_ = ~v25 & ~new_n895_;
  assign new_n897_ = ~v24 & new_n896_;
  assign new_n898_ = ~v10 & new_n897_;
  assign new_n899_ = ~v9 & new_n898_;
  assign new_n900_ = ~v8 & new_n899_;
  assign new_n901_ = v7 & new_n900_;
  assign new_n902_ = ~v4 & new_n901_;
  assign new_n903_ = ~v3 & new_n902_;
  assign new_n904_ = v0 & new_n903_;
  assign new_n905_ = ~new_n891_ & ~new_n904_;
  assign new_n906_ = v6 & ~new_n905_;
  assign new_n907_ = v2 & v9;
  assign new_n908_ = v1 & new_n907_;
  assign new_n909_ = v7 & new_n118_;
  assign new_n910_ = new_n114_ & new_n909_;
  assign new_n911_ = ~new_n908_ & ~new_n910_;
  assign new_n912_ = ~v25 & ~new_n911_;
  assign new_n913_ = ~v24 & new_n912_;
  assign new_n914_ = ~v23 & new_n913_;
  assign new_n915_ = ~v8 & new_n914_;
  assign new_n916_ = ~v6 & new_n915_;
  assign new_n917_ = v4 & new_n916_;
  assign new_n918_ = v3 & new_n917_;
  assign new_n919_ = ~v0 & new_n918_;
  assign new_n920_ = ~new_n906_ & ~new_n919_;
  assign new_n921_ = ~v5 & ~new_n920_;
  assign new_n922_ = v1 & new_n361_;
  assign new_n923_ = new_n77_ & new_n187_;
  assign new_n924_ = new_n922_ & new_n923_;
  assign new_n925_ = ~v1 & new_n358_;
  assign new_n926_ = new_n76_ & new_n188_;
  assign new_n927_ = new_n925_ & new_n926_;
  assign new_n928_ = ~new_n924_ & ~new_n927_;
  assign new_n929_ = ~v3 & ~new_n928_;
  assign new_n930_ = v6 & ~v10;
  assign new_n931_ = v6 & ~new_n930_;
  assign new_n932_ = ~v25 & ~new_n931_;
  assign new_n933_ = ~v24 & new_n932_;
  assign new_n934_ = ~v7 & new_n933_;
  assign new_n935_ = v3 & new_n934_;
  assign new_n936_ = v2 & new_n935_;
  assign new_n937_ = v1 & new_n936_;
  assign new_n938_ = ~new_n929_ & ~new_n937_;
  assign new_n939_ = v9 & ~new_n938_;
  assign new_n940_ = v4 & new_n939_;
  assign new_n941_ = v7 & new_n676_;
  assign new_n942_ = v6 & new_n941_;
  assign new_n943_ = ~v4 & new_n942_;
  assign new_n944_ = v3 & new_n943_;
  assign new_n945_ = v2 & new_n944_;
  assign new_n946_ = ~v1 & new_n945_;
  assign new_n947_ = ~new_n940_ & ~new_n946_;
  assign new_n948_ = ~v8 & ~new_n947_;
  assign new_n949_ = v4 & v6;
  assign new_n950_ = v3 & new_n949_;
  assign new_n951_ = new_n418_ & new_n950_;
  assign new_n952_ = v7 & new_n321_;
  assign new_n953_ = v10 & new_n187_;
  assign new_n954_ = new_n952_ & new_n953_;
  assign new_n955_ = new_n951_ & new_n954_;
  assign new_n956_ = ~new_n948_ & ~new_n955_;
  assign new_n957_ = ~v23 & ~new_n956_;
  assign new_n958_ = v5 & new_n957_;
  assign new_n959_ = ~v0 & new_n958_;
  assign new_n960_ = ~new_n921_ & ~new_n959_;
  assign \v26.9  = ~v22 & ~new_n960_;
  assign new_n962_ = ~v2 & new_n949_;
  assign new_n963_ = v1 & new_n962_;
  assign new_n964_ = v0 & new_n963_;
  assign new_n965_ = ~v4 & new_n552_;
  assign new_n966_ = new_n545_ & new_n965_;
  assign new_n967_ = ~new_n964_ & ~new_n966_;
  assign new_n968_ = ~v25 & ~new_n967_;
  assign new_n969_ = ~v24 & new_n968_;
  assign new_n970_ = v2 & ~v4;
  assign new_n971_ = new_n95_ & new_n970_;
  assign new_n972_ = new_n200_ & new_n552_;
  assign new_n973_ = new_n971_ & new_n972_;
  assign new_n974_ = ~new_n969_ & ~new_n973_;
  assign new_n975_ = ~v8 & ~new_n974_;
  assign new_n976_ = v8 & new_n194_;
  assign new_n977_ = v6 & new_n976_;
  assign new_n978_ = v4 & new_n977_;
  assign new_n979_ = ~v2 & new_n978_;
  assign new_n980_ = v1 & new_n979_;
  assign new_n981_ = v0 & new_n980_;
  assign new_n982_ = ~new_n975_ & ~new_n981_;
  assign new_n983_ = ~v4 & new_n292_;
  assign new_n984_ = v4 & new_n382_;
  assign new_n985_ = ~new_n983_ & ~new_n984_;
  assign new_n986_ = ~v0 & ~new_n985_;
  assign new_n987_ = v0 & ~v4;
  assign new_n988_ = new_n292_ & new_n987_;
  assign new_n989_ = ~new_n986_ & ~new_n988_;
  assign new_n990_ = ~v2 & ~new_n989_;
  assign new_n991_ = ~v4 & v6;
  assign new_n992_ = v2 & new_n991_;
  assign new_n993_ = v0 & new_n992_;
  assign new_n994_ = ~new_n990_ & ~new_n993_;
  assign new_n995_ = ~v25 & ~new_n994_;
  assign new_n996_ = ~v9 & new_n995_;
  assign new_n997_ = ~v1 & new_n996_;
  assign new_n998_ = new_n289_ & new_n346_;
  assign new_n999_ = v9 & v25;
  assign new_n1000_ = new_n292_ & new_n999_;
  assign new_n1001_ = new_n998_ & new_n1000_;
  assign new_n1002_ = ~new_n997_ & ~new_n1001_;
  assign new_n1003_ = ~v24 & ~new_n1002_;
  assign new_n1004_ = ~v10 & new_n1003_;
  assign new_n1005_ = new_n982_ & ~new_n1004_;
  assign new_n1006_ = v7 & ~new_n1005_;
  assign new_n1007_ = ~v4 & v9;
  assign new_n1008_ = v0 & new_n1007_;
  assign new_n1009_ = ~v0 & ~v2;
  assign new_n1010_ = v4 & ~v9;
  assign new_n1011_ = new_n1009_ & new_n1010_;
  assign new_n1012_ = ~new_n1008_ & ~new_n1011_;
  assign new_n1013_ = ~v25 & ~new_n1012_;
  assign new_n1014_ = ~v24 & new_n1013_;
  assign new_n1015_ = ~v10 & new_n1014_;
  assign new_n1016_ = v8 & new_n1015_;
  assign new_n1017_ = ~v7 & new_n1016_;
  assign new_n1018_ = v6 & new_n1017_;
  assign new_n1019_ = ~v1 & new_n1018_;
  assign new_n1020_ = ~new_n1006_ & ~new_n1019_;
  assign new_n1021_ = v3 & ~new_n1020_;
  assign new_n1022_ = ~v9 & ~new_n699_;
  assign new_n1023_ = ~v8 & new_n1022_;
  assign new_n1024_ = ~v4 & new_n1023_;
  assign new_n1025_ = ~v2 & new_n1024_;
  assign new_n1026_ = v4 & ~v6;
  assign new_n1027_ = new_n537_ & new_n1026_;
  assign new_n1028_ = ~v7 & v8;
  assign new_n1029_ = v9 & new_n433_;
  assign new_n1030_ = new_n1028_ & new_n1029_;
  assign new_n1031_ = new_n1027_ & new_n1030_;
  assign new_n1032_ = ~new_n1025_ & ~new_n1031_;
  assign new_n1033_ = ~v24 & ~new_n1032_;
  assign new_n1034_ = ~v3 & new_n1033_;
  assign new_n1035_ = ~v1 & new_n1034_;
  assign new_n1036_ = ~new_n1021_ & ~new_n1035_;
  assign new_n1037_ = ~v5 & ~new_n1036_;
  assign new_n1038_ = v2 & ~new_n782_;
  assign new_n1039_ = ~v9 & ~v24;
  assign new_n1040_ = ~v8 & new_n1039_;
  assign new_n1041_ = ~v6 & new_n1040_;
  assign new_n1042_ = ~v3 & new_n1041_;
  assign new_n1043_ = ~v2 & new_n1042_;
  assign new_n1044_ = ~new_n1038_ & ~new_n1043_;
  assign new_n1045_ = v7 & ~new_n1044_;
  assign new_n1046_ = v6 & ~v7;
  assign new_n1047_ = new_n712_ & new_n1046_;
  assign new_n1048_ = new_n194_ & new_n257_;
  assign new_n1049_ = new_n1047_ & new_n1048_;
  assign new_n1050_ = ~new_n1045_ & ~new_n1049_;
  assign new_n1051_ = v10 & ~new_n1050_;
  assign new_n1052_ = ~v1 & new_n1051_;
  assign new_n1053_ = ~v3 & new_n1046_;
  assign new_n1054_ = new_n853_ & new_n1053_;
  assign new_n1055_ = ~v10 & new_n187_;
  assign new_n1056_ = new_n257_ & new_n1055_;
  assign new_n1057_ = new_n1054_ & new_n1056_;
  assign new_n1058_ = ~new_n1052_ & ~new_n1057_;
  assign new_n1059_ = v5 & ~new_n1058_;
  assign new_n1060_ = v4 & new_n1059_;
  assign new_n1061_ = ~v0 & new_n1060_;
  assign new_n1062_ = ~new_n1037_ & ~new_n1061_;
  assign new_n1063_ = ~v23 & ~new_n1062_;
  assign new_n1064_ = ~v25 & ~new_n716_;
  assign new_n1065_ = ~v24 & new_n1064_;
  assign new_n1066_ = v23 & new_n1065_;
  assign new_n1067_ = ~v10 & new_n1066_;
  assign new_n1068_ = ~v9 & new_n1067_;
  assign new_n1069_ = ~v8 & new_n1068_;
  assign new_n1070_ = v7 & new_n1069_;
  assign new_n1071_ = v6 & new_n1070_;
  assign new_n1072_ = ~v5 & new_n1071_;
  assign new_n1073_ = ~v4 & new_n1072_;
  assign new_n1074_ = v0 & new_n1073_;
  assign new_n1075_ = ~new_n1063_ & ~new_n1074_;
  assign \v26.10  = ~v22 & ~new_n1075_;
  assign new_n1077_ = v1 & new_n255_;
  assign new_n1078_ = new_n589_ & new_n825_;
  assign new_n1079_ = ~new_n1077_ & ~new_n1078_;
  assign new_n1080_ = ~v25 & ~new_n1079_;
  assign new_n1081_ = v7 & new_n1080_;
  assign new_n1082_ = ~v5 & new_n1081_;
  assign new_n1083_ = v0 & new_n1082_;
  assign new_n1084_ = new_n254_ & new_n725_;
  assign new_n1085_ = new_n73_ & new_n999_;
  assign new_n1086_ = new_n1084_ & new_n1085_;
  assign new_n1087_ = ~new_n1083_ & ~new_n1086_;
  assign new_n1088_ = ~v8 & ~new_n1087_;
  assign new_n1089_ = v0 & ~new_n835_;
  assign new_n1090_ = ~v0 & new_n834_;
  assign new_n1091_ = ~new_n1089_ & ~new_n1090_;
  assign new_n1092_ = ~v4 & ~new_n1091_;
  assign new_n1093_ = ~v0 & v4;
  assign new_n1094_ = ~v7 & ~v9;
  assign new_n1095_ = new_n1093_ & new_n1094_;
  assign new_n1096_ = ~new_n1092_ & ~new_n1095_;
  assign new_n1097_ = ~v1 & ~new_n1096_;
  assign new_n1098_ = v1 & new_n854_;
  assign new_n1099_ = v0 & new_n1098_;
  assign new_n1100_ = ~new_n1097_ & ~new_n1099_;
  assign new_n1101_ = ~v25 & ~new_n1100_;
  assign new_n1102_ = v8 & new_n1101_;
  assign new_n1103_ = ~v5 & new_n1102_;
  assign new_n1104_ = v3 & new_n1103_;
  assign new_n1105_ = ~new_n1088_ & ~new_n1104_;
  assign new_n1106_ = ~v10 & ~new_n1105_;
  assign new_n1107_ = ~v8 & new_n612_;
  assign new_n1108_ = v25 & ~new_n1107_;
  assign new_n1109_ = v10 & ~new_n1108_;
  assign new_n1110_ = v7 & new_n1109_;
  assign new_n1111_ = ~v5 & new_n1110_;
  assign new_n1112_ = v4 & new_n1111_;
  assign new_n1113_ = v3 & new_n1112_;
  assign new_n1114_ = v1 & new_n1113_;
  assign new_n1115_ = v0 & new_n1114_;
  assign new_n1116_ = ~new_n1106_ & ~new_n1115_;
  assign new_n1117_ = ~v2 & ~new_n1116_;
  assign new_n1118_ = ~v7 & new_n310_;
  assign new_n1119_ = ~new_n834_ & ~new_n1118_;
  assign new_n1120_ = ~v10 & ~new_n1119_;
  assign new_n1121_ = ~v5 & new_n1120_;
  assign new_n1122_ = ~v4 & new_n1121_;
  assign new_n1123_ = v0 & new_n1122_;
  assign new_n1124_ = ~v0 & new_n419_;
  assign new_n1125_ = ~v7 & ~v8;
  assign new_n1126_ = new_n398_ & new_n1125_;
  assign new_n1127_ = new_n1124_ & new_n1126_;
  assign new_n1128_ = ~new_n1123_ & ~new_n1127_;
  assign new_n1129_ = ~v25 & ~new_n1128_;
  assign new_n1130_ = v3 & new_n1129_;
  assign new_n1131_ = v2 & new_n1130_;
  assign new_n1132_ = ~v1 & new_n1131_;
  assign new_n1133_ = ~new_n1117_ & ~new_n1132_;
  assign new_n1134_ = ~v23 & ~new_n1133_;
  assign new_n1135_ = v23 & new_n1064_;
  assign new_n1136_ = ~v10 & new_n1135_;
  assign new_n1137_ = ~v9 & new_n1136_;
  assign new_n1138_ = ~v8 & new_n1137_;
  assign new_n1139_ = v7 & new_n1138_;
  assign new_n1140_ = ~v5 & new_n1139_;
  assign new_n1141_ = ~v4 & new_n1140_;
  assign new_n1142_ = v0 & new_n1141_;
  assign new_n1143_ = ~new_n1134_ & ~new_n1142_;
  assign new_n1144_ = v6 & ~new_n1143_;
  assign new_n1145_ = ~v3 & new_n399_;
  assign new_n1146_ = v2 & new_n1145_;
  assign new_n1147_ = v3 & ~v5;
  assign new_n1148_ = ~v2 & new_n1147_;
  assign new_n1149_ = new_n909_ & new_n1148_;
  assign new_n1150_ = ~new_n1146_ & ~new_n1149_;
  assign new_n1151_ = ~v25 & ~new_n1150_;
  assign new_n1152_ = ~v23 & new_n1151_;
  assign new_n1153_ = ~v8 & new_n1152_;
  assign new_n1154_ = ~v6 & new_n1153_;
  assign new_n1155_ = v4 & new_n1154_;
  assign new_n1156_ = ~v1 & new_n1155_;
  assign new_n1157_ = ~v0 & new_n1156_;
  assign new_n1158_ = ~new_n1144_ & ~new_n1157_;
  assign new_n1159_ = ~v24 & ~new_n1158_;
  assign new_n1160_ = new_n138_ & new_n725_;
  assign new_n1161_ = new_n545_ & new_n1160_;
  assign new_n1162_ = v7 & new_n257_;
  assign new_n1163_ = v10 & ~v23;
  assign new_n1164_ = new_n188_ & new_n1163_;
  assign new_n1165_ = new_n1162_ & new_n1164_;
  assign new_n1166_ = new_n1161_ & new_n1165_;
  assign new_n1167_ = ~new_n1159_ & ~new_n1166_;
  assign \v26.11  = ~v22 & ~new_n1167_;
  assign new_n1169_ = ~v9 & new_n430_;
  assign new_n1170_ = ~v4 & ~v8;
  assign new_n1171_ = ~v2 & new_n1170_;
  assign new_n1172_ = new_n1169_ & new_n1171_;
  assign new_n1173_ = v4 & v8;
  assign new_n1174_ = v2 & new_n1173_;
  assign new_n1175_ = new_n1029_ & new_n1174_;
  assign new_n1176_ = ~new_n1172_ & ~new_n1175_;
  assign new_n1177_ = ~v23 & ~new_n1176_;
  assign new_n1178_ = ~v7 & new_n1177_;
  assign new_n1179_ = ~v6 & new_n1178_;
  assign new_n1180_ = ~v0 & new_n1179_;
  assign new_n1181_ = ~v4 & new_n533_;
  assign new_n1182_ = new_n478_ & new_n1181_;
  assign new_n1183_ = ~v10 & new_n139_;
  assign new_n1184_ = new_n368_ & new_n1183_;
  assign new_n1185_ = new_n1182_ & new_n1184_;
  assign new_n1186_ = ~new_n1180_ & ~new_n1185_;
  assign new_n1187_ = ~v1 & ~new_n1186_;
  assign new_n1188_ = ~v9 & new_n1183_;
  assign new_n1189_ = ~v8 & new_n1188_;
  assign new_n1190_ = v7 & new_n1189_;
  assign new_n1191_ = v6 & new_n1190_;
  assign new_n1192_ = ~v4 & new_n1191_;
  assign new_n1193_ = v1 & new_n1192_;
  assign new_n1194_ = v0 & new_n1193_;
  assign new_n1195_ = ~new_n1187_ & ~new_n1194_;
  assign new_n1196_ = ~v3 & ~new_n1195_;
  assign new_n1197_ = new_n129_ & new_n346_;
  assign new_n1198_ = new_n139_ & new_n970_;
  assign new_n1199_ = ~new_n1197_ & ~new_n1198_;
  assign new_n1200_ = v1 & ~new_n1199_;
  assign new_n1201_ = ~v4 & new_n139_;
  assign new_n1202_ = new_n418_ & new_n1201_;
  assign new_n1203_ = ~new_n1200_ & ~new_n1202_;
  assign new_n1204_ = ~v10 & ~new_n1203_;
  assign new_n1205_ = ~v9 & new_n1204_;
  assign new_n1206_ = ~v8 & new_n1205_;
  assign new_n1207_ = v7 & new_n1206_;
  assign new_n1208_ = v6 & new_n1207_;
  assign new_n1209_ = v3 & new_n1208_;
  assign new_n1210_ = v0 & new_n1209_;
  assign new_n1211_ = ~new_n1196_ & ~new_n1210_;
  assign new_n1212_ = ~v24 & ~new_n1211_;
  assign new_n1213_ = ~v23 & new_n200_;
  assign new_n1214_ = v10 & new_n1213_;
  assign new_n1215_ = ~v8 & new_n1214_;
  assign new_n1216_ = v7 & new_n1215_;
  assign new_n1217_ = ~v6 & new_n1216_;
  assign new_n1218_ = ~v4 & new_n1217_;
  assign new_n1219_ = v3 & new_n1218_;
  assign new_n1220_ = v2 & new_n1219_;
  assign new_n1221_ = ~v1 & new_n1220_;
  assign new_n1222_ = ~v0 & new_n1221_;
  assign new_n1223_ = ~new_n1212_ & ~new_n1222_;
  assign new_n1224_ = ~v5 & ~new_n1223_;
  assign new_n1225_ = ~v4 & new_n422_;
  assign new_n1226_ = v3 & new_n1225_;
  assign new_n1227_ = new_n473_ & new_n725_;
  assign new_n1228_ = ~new_n1226_ & ~new_n1227_;
  assign new_n1229_ = ~v25 & ~new_n1228_;
  assign new_n1230_ = v24 & new_n1229_;
  assign new_n1231_ = ~v23 & new_n1230_;
  assign new_n1232_ = ~v8 & new_n1231_;
  assign new_n1233_ = v7 & new_n1232_;
  assign new_n1234_ = v5 & new_n1233_;
  assign new_n1235_ = v2 & new_n1234_;
  assign new_n1236_ = ~v1 & new_n1235_;
  assign new_n1237_ = ~v0 & new_n1236_;
  assign new_n1238_ = ~new_n1224_ & ~new_n1237_;
  assign \v26.12  = ~v22 & ~new_n1238_;
  assign new_n1240_ = ~v2 & new_n1039_;
  assign new_n1241_ = ~new_n907_ & ~new_n1240_;
  assign new_n1242_ = ~v25 & ~new_n1241_;
  assign new_n1243_ = ~v2 & ~v9;
  assign new_n1244_ = new_n187_ & new_n1243_;
  assign new_n1245_ = ~new_n1242_ & ~new_n1244_;
  assign new_n1246_ = ~v6 & ~new_n1245_;
  assign new_n1247_ = v5 & new_n1246_;
  assign new_n1248_ = v4 & new_n1247_;
  assign new_n1249_ = new_n194_ & new_n422_;
  assign new_n1250_ = new_n495_ & new_n1249_;
  assign new_n1251_ = ~new_n1248_ & ~new_n1250_;
  assign new_n1252_ = ~v3 & ~new_n1251_;
  assign new_n1253_ = ~v1 & new_n1252_;
  assign new_n1254_ = ~v0 & new_n1253_;
  assign new_n1255_ = v9 & new_n187_;
  assign new_n1256_ = new_n585_ & new_n1255_;
  assign new_n1257_ = new_n766_ & new_n1256_;
  assign new_n1258_ = ~new_n1254_ & ~new_n1257_;
  assign new_n1259_ = v7 & ~new_n1258_;
  assign new_n1260_ = v9 & new_n194_;
  assign new_n1261_ = new_n538_ & new_n1260_;
  assign new_n1262_ = new_n727_ & new_n1261_;
  assign new_n1263_ = ~new_n1259_ & ~new_n1262_;
  assign new_n1264_ = ~v23 & ~new_n1263_;
  assign new_n1265_ = ~v22 & new_n1264_;
  assign new_n1266_ = v10 & new_n1265_;
  assign \v26.13  = ~v8 & new_n1266_;
  assign new_n1268_ = v2 & new_n616_;
  assign new_n1269_ = ~new_n1244_ & ~new_n1268_;
  assign new_n1270_ = v10 & ~new_n1269_;
  assign new_n1271_ = ~v6 & new_n1270_;
  assign new_n1272_ = v5 & new_n1271_;
  assign new_n1273_ = ~v3 & new_n1272_;
  assign new_n1274_ = ~v1 & new_n1273_;
  assign new_n1275_ = ~v0 & new_n1274_;
  assign new_n1276_ = new_n289_ & new_n1148_;
  assign new_n1277_ = v6 & v9;
  assign new_n1278_ = new_n1055_ & new_n1277_;
  assign new_n1279_ = new_n1276_ & new_n1278_;
  assign new_n1280_ = ~new_n1275_ & ~new_n1279_;
  assign new_n1281_ = ~v23 & ~new_n1280_;
  assign new_n1282_ = v23 & new_n188_;
  assign new_n1283_ = new_n473_ & new_n1282_;
  assign new_n1284_ = new_n147_ & new_n1283_;
  assign new_n1285_ = ~new_n1281_ & ~new_n1284_;
  assign new_n1286_ = v7 & ~new_n1285_;
  assign new_n1287_ = ~v23 & ~v24;
  assign new_n1288_ = ~new_n561_ & ~new_n1287_;
  assign new_n1289_ = ~v25 & ~new_n1288_;
  assign new_n1290_ = v10 & new_n1289_;
  assign new_n1291_ = v9 & new_n1290_;
  assign new_n1292_ = ~v7 & new_n1291_;
  assign new_n1293_ = ~v6 & new_n1292_;
  assign new_n1294_ = v5 & new_n1293_;
  assign new_n1295_ = ~v3 & new_n1294_;
  assign new_n1296_ = v2 & new_n1295_;
  assign new_n1297_ = ~v1 & new_n1296_;
  assign new_n1298_ = ~v0 & new_n1297_;
  assign new_n1299_ = ~new_n1286_ & ~new_n1298_;
  assign new_n1300_ = ~v22 & ~new_n1299_;
  assign new_n1301_ = ~v8 & new_n1300_;
  assign \v26.14  = v4 & new_n1301_;
  assign new_n1303_ = v23 & ~new_n714_;
  assign new_n1304_ = ~v10 & new_n1303_;
  assign new_n1305_ = v6 & new_n1304_;
  assign new_n1306_ = v0 & new_n1305_;
  assign new_n1307_ = ~v0 & new_n712_;
  assign new_n1308_ = ~v6 & new_n1163_;
  assign new_n1309_ = new_n1307_ & new_n1308_;
  assign new_n1310_ = ~new_n1306_ & ~new_n1309_;
  assign new_n1311_ = v25 & ~new_n1310_;
  assign new_n1312_ = ~v8 & new_n1311_;
  assign new_n1313_ = v8 & new_n173_;
  assign new_n1314_ = ~v6 & new_n1313_;
  assign new_n1315_ = v3 & new_n1314_;
  assign new_n1316_ = v2 & new_n1315_;
  assign new_n1317_ = ~v0 & new_n1316_;
  assign new_n1318_ = ~new_n1312_ & ~new_n1317_;
  assign new_n1319_ = ~v24 & ~new_n1318_;
  assign new_n1320_ = v7 & new_n1319_;
  assign new_n1321_ = ~v10 & new_n729_;
  assign new_n1322_ = ~v8 & new_n1321_;
  assign new_n1323_ = ~v7 & new_n1322_;
  assign new_n1324_ = ~v6 & new_n1323_;
  assign new_n1325_ = ~v3 & new_n1324_;
  assign new_n1326_ = ~v2 & new_n1325_;
  assign new_n1327_ = ~v0 & new_n1326_;
  assign new_n1328_ = ~new_n1320_ & ~new_n1327_;
  assign new_n1329_ = ~v4 & ~new_n1328_;
  assign new_n1330_ = v6 & new_n1028_;
  assign new_n1331_ = v7 & ~v8;
  assign new_n1332_ = ~v6 & new_n1331_;
  assign new_n1333_ = ~new_n1330_ & ~new_n1332_;
  assign new_n1334_ = ~v25 & ~new_n1333_;
  assign new_n1335_ = ~v24 & new_n1334_;
  assign new_n1336_ = ~v23 & new_n1335_;
  assign new_n1337_ = ~v10 & new_n1336_;
  assign new_n1338_ = v4 & new_n1337_;
  assign new_n1339_ = v3 & new_n1338_;
  assign new_n1340_ = ~v2 & new_n1339_;
  assign new_n1341_ = ~v0 & new_n1340_;
  assign new_n1342_ = ~new_n1329_ & ~new_n1341_;
  assign new_n1343_ = ~v5 & ~new_n1342_;
  assign new_n1344_ = v3 & new_n882_;
  assign new_n1345_ = new_n953_ & new_n1344_;
  assign new_n1346_ = ~v3 & new_n1125_;
  assign new_n1347_ = ~v10 & ~v19;
  assign new_n1348_ = new_n188_ & new_n1347_;
  assign new_n1349_ = new_n1346_ & new_n1348_;
  assign new_n1350_ = ~new_n1345_ & ~new_n1349_;
  assign new_n1351_ = ~v23 & ~new_n1350_;
  assign new_n1352_ = v6 & new_n1351_;
  assign new_n1353_ = v5 & new_n1352_;
  assign new_n1354_ = v4 & new_n1353_;
  assign new_n1355_ = v2 & new_n1354_;
  assign new_n1356_ = ~v0 & new_n1355_;
  assign new_n1357_ = ~new_n1343_ & ~new_n1356_;
  assign new_n1358_ = ~v1 & ~new_n1357_;
  assign new_n1359_ = ~v2 & ~new_n713_;
  assign new_n1360_ = v25 & ~new_n1359_;
  assign new_n1361_ = ~v24 & new_n1360_;
  assign new_n1362_ = v23 & new_n1361_;
  assign new_n1363_ = ~v10 & new_n1362_;
  assign new_n1364_ = ~v8 & new_n1363_;
  assign new_n1365_ = v7 & new_n1364_;
  assign new_n1366_ = v6 & new_n1365_;
  assign new_n1367_ = ~v5 & new_n1366_;
  assign new_n1368_ = ~v4 & new_n1367_;
  assign new_n1369_ = v1 & new_n1368_;
  assign new_n1370_ = v0 & new_n1369_;
  assign new_n1371_ = ~new_n1358_ & ~new_n1370_;
  assign new_n1372_ = ~v9 & ~new_n1371_;
  assign new_n1373_ = new_n418_ & new_n439_;
  assign new_n1374_ = new_n76_ & new_n117_;
  assign new_n1375_ = new_n1373_ & new_n1374_;
  assign new_n1376_ = new_n725_ & new_n853_;
  assign new_n1377_ = new_n77_ & new_n546_;
  assign new_n1378_ = new_n1376_ & new_n1377_;
  assign new_n1379_ = ~new_n1375_ & ~new_n1378_;
  assign new_n1380_ = v25 & ~new_n1379_;
  assign new_n1381_ = ~v0 & new_n1380_;
  assign new_n1382_ = v0 & ~v1;
  assign new_n1383_ = v2 & new_n255_;
  assign new_n1384_ = new_n1382_ & new_n1383_;
  assign new_n1385_ = v7 & new_n433_;
  assign new_n1386_ = new_n585_ & new_n1385_;
  assign new_n1387_ = new_n1384_ & new_n1386_;
  assign new_n1388_ = ~new_n1381_ & ~new_n1387_;
  assign new_n1389_ = ~v24 & ~new_n1388_;
  assign new_n1390_ = ~v23 & new_n1389_;
  assign new_n1391_ = v9 & new_n1390_;
  assign new_n1392_ = ~v8 & new_n1391_;
  assign new_n1393_ = ~new_n1372_ & ~new_n1392_;
  assign \v26.15  = ~v22 & ~new_n1393_;
  assign new_n1395_ = v5 & v8;
  assign new_n1396_ = new_n713_ & new_n1395_;
  assign new_n1397_ = new_n187_ & new_n1347_;
  assign new_n1398_ = new_n1396_ & new_n1397_;
  assign new_n1399_ = v2 & new_n1147_;
  assign new_n1400_ = new_n188_ & new_n359_;
  assign new_n1401_ = new_n1399_ & new_n1400_;
  assign new_n1402_ = ~new_n1398_ & ~new_n1401_;
  assign new_n1403_ = ~v6 & ~new_n1402_;
  assign new_n1404_ = ~v1 & new_n1403_;
  assign new_n1405_ = ~v0 & new_n1404_;
  assign new_n1406_ = ~v3 & ~v5;
  assign new_n1407_ = ~v2 & new_n1406_;
  assign new_n1408_ = new_n289_ & new_n1407_;
  assign new_n1409_ = ~v10 & new_n200_;
  assign new_n1410_ = new_n292_ & new_n1409_;
  assign new_n1411_ = new_n1408_ & new_n1410_;
  assign new_n1412_ = ~new_n1405_ & ~new_n1411_;
  assign new_n1413_ = ~v4 & ~new_n1412_;
  assign new_n1414_ = ~v5 & new_n195_;
  assign new_n1415_ = v4 & new_n1414_;
  assign new_n1416_ = v3 & new_n1415_;
  assign new_n1417_ = ~v2 & new_n1416_;
  assign new_n1418_ = v1 & new_n1417_;
  assign new_n1419_ = v0 & new_n1418_;
  assign new_n1420_ = ~new_n1413_ & ~new_n1419_;
  assign new_n1421_ = ~new_n310_ & ~new_n368_;
  assign new_n1422_ = ~v10 & ~new_n1421_;
  assign new_n1423_ = ~v5 & new_n1422_;
  assign new_n1424_ = v0 & new_n1423_;
  assign new_n1425_ = ~v0 & v5;
  assign new_n1426_ = new_n299_ & new_n1425_;
  assign new_n1427_ = ~new_n1424_ & ~new_n1426_;
  assign new_n1428_ = ~v24 & ~new_n1427_;
  assign new_n1429_ = v6 & new_n1428_;
  assign new_n1430_ = v3 & new_n1429_;
  assign new_n1431_ = ~v0 & ~v3;
  assign new_n1432_ = new_n138_ & new_n1431_;
  assign new_n1433_ = new_n259_ & new_n1432_;
  assign new_n1434_ = ~new_n1430_ & ~new_n1433_;
  assign new_n1435_ = v4 & ~new_n1434_;
  assign new_n1436_ = new_n479_ & new_n788_;
  assign new_n1437_ = v6 & ~v8;
  assign new_n1438_ = new_n485_ & new_n1437_;
  assign new_n1439_ = new_n1436_ & new_n1438_;
  assign new_n1440_ = ~new_n1435_ & ~new_n1439_;
  assign new_n1441_ = ~v1 & ~new_n1440_;
  assign new_n1442_ = ~v5 & ~v9;
  assign new_n1443_ = v5 & new_n310_;
  assign new_n1444_ = ~new_n1442_ & ~new_n1443_;
  assign new_n1445_ = ~v3 & ~new_n1444_;
  assign new_n1446_ = new_n368_ & new_n1147_;
  assign new_n1447_ = ~new_n1445_ & ~new_n1446_;
  assign new_n1448_ = v24 & ~new_n1447_;
  assign new_n1449_ = ~v10 & new_n1448_;
  assign new_n1450_ = v6 & new_n1449_;
  assign new_n1451_ = ~v4 & new_n1450_;
  assign new_n1452_ = v1 & new_n1451_;
  assign new_n1453_ = v0 & new_n1452_;
  assign new_n1454_ = ~new_n1441_ & ~new_n1453_;
  assign new_n1455_ = v25 & ~new_n1454_;
  assign new_n1456_ = ~v0 & new_n824_;
  assign new_n1457_ = v9 & new_n258_;
  assign new_n1458_ = new_n1456_ & new_n1457_;
  assign new_n1459_ = v0 & new_n829_;
  assign new_n1460_ = new_n497_ & new_n1459_;
  assign new_n1461_ = ~new_n1458_ & ~new_n1460_;
  assign new_n1462_ = v6 & ~new_n1461_;
  assign new_n1463_ = ~v6 & new_n263_;
  assign new_n1464_ = v4 & new_n1463_;
  assign new_n1465_ = v1 & new_n1464_;
  assign new_n1466_ = ~v0 & new_n1465_;
  assign new_n1467_ = ~new_n1462_ & ~new_n1466_;
  assign new_n1468_ = ~v8 & ~new_n1467_;
  assign new_n1469_ = v6 & new_n877_;
  assign new_n1470_ = ~v4 & new_n1469_;
  assign new_n1471_ = ~v1 & new_n1470_;
  assign new_n1472_ = v0 & new_n1471_;
  assign new_n1473_ = ~new_n1468_ & ~new_n1472_;
  assign new_n1474_ = ~v25 & ~new_n1473_;
  assign new_n1475_ = ~v5 & new_n1474_;
  assign new_n1476_ = v3 & new_n1475_;
  assign new_n1477_ = ~new_n1455_ & ~new_n1476_;
  assign new_n1478_ = v2 & ~new_n1477_;
  assign new_n1479_ = ~v0 & ~v24;
  assign new_n1480_ = ~v0 & ~new_n1479_;
  assign new_n1481_ = ~v25 & ~new_n1480_;
  assign new_n1482_ = ~v9 & new_n1481_;
  assign new_n1483_ = v3 & new_n1482_;
  assign new_n1484_ = new_n1255_ & new_n1431_;
  assign new_n1485_ = ~new_n1483_ & ~new_n1484_;
  assign new_n1486_ = v8 & ~new_n1485_;
  assign new_n1487_ = ~v9 & ~new_n201_;
  assign new_n1488_ = ~v8 & new_n1487_;
  assign new_n1489_ = ~v3 & new_n1488_;
  assign new_n1490_ = v0 & new_n1489_;
  assign new_n1491_ = ~new_n1486_ & ~new_n1490_;
  assign new_n1492_ = ~v1 & ~new_n1491_;
  assign new_n1493_ = new_n200_ & new_n368_;
  assign new_n1494_ = new_n750_ & new_n1493_;
  assign new_n1495_ = ~new_n1492_ & ~new_n1494_;
  assign new_n1496_ = ~v10 & ~new_n1495_;
  assign new_n1497_ = v6 & new_n1496_;
  assign new_n1498_ = ~v5 & new_n1497_;
  assign new_n1499_ = ~v4 & new_n1498_;
  assign new_n1500_ = ~v2 & new_n1499_;
  assign new_n1501_ = ~new_n1478_ & ~new_n1500_;
  assign new_n1502_ = new_n1420_ & new_n1501_;
  assign new_n1503_ = v7 & ~new_n1502_;
  assign new_n1504_ = ~v1 & new_n344_;
  assign new_n1505_ = v0 & new_n1504_;
  assign new_n1506_ = v4 & new_n278_;
  assign new_n1507_ = new_n254_ & new_n1506_;
  assign new_n1508_ = ~new_n1505_ & ~new_n1507_;
  assign new_n1509_ = v6 & ~new_n1508_;
  assign new_n1510_ = ~v6 & new_n278_;
  assign new_n1511_ = new_n1456_ & new_n1510_;
  assign new_n1512_ = ~new_n1509_ & ~new_n1511_;
  assign new_n1513_ = v2 & ~new_n1512_;
  assign new_n1514_ = ~v2 & new_n983_;
  assign new_n1515_ = ~v1 & new_n1514_;
  assign new_n1516_ = v0 & new_n1515_;
  assign new_n1517_ = ~new_n1513_ & ~new_n1516_;
  assign new_n1518_ = ~v25 & ~new_n1517_;
  assign new_n1519_ = v3 & new_n1518_;
  assign new_n1520_ = v8 & new_n200_;
  assign new_n1521_ = v6 & new_n1520_;
  assign new_n1522_ = ~v4 & new_n1521_;
  assign new_n1523_ = ~v3 & new_n1522_;
  assign new_n1524_ = v1 & new_n1523_;
  assign new_n1525_ = v0 & new_n1524_;
  assign new_n1526_ = ~new_n1519_ & ~new_n1525_;
  assign new_n1527_ = ~v5 & ~new_n1526_;
  assign new_n1528_ = ~v8 & new_n200_;
  assign new_n1529_ = v5 & new_n1528_;
  assign new_n1530_ = v4 & new_n1529_;
  assign new_n1531_ = v3 & new_n1530_;
  assign new_n1532_ = v2 & new_n1531_;
  assign new_n1533_ = v1 & new_n1532_;
  assign new_n1534_ = ~v0 & new_n1533_;
  assign new_n1535_ = ~new_n1527_ & ~new_n1534_;
  assign new_n1536_ = ~v10 & ~new_n1535_;
  assign new_n1537_ = v5 & v25;
  assign new_n1538_ = ~v5 & ~v25;
  assign new_n1539_ = ~new_n1537_ & ~new_n1538_;
  assign new_n1540_ = v3 & ~new_n1539_;
  assign new_n1541_ = v1 & new_n1540_;
  assign new_n1542_ = new_n589_ & new_n1537_;
  assign new_n1543_ = ~new_n1541_ & ~new_n1542_;
  assign new_n1544_ = v24 & ~new_n1543_;
  assign new_n1545_ = v10 & new_n1544_;
  assign new_n1546_ = ~v8 & new_n1545_;
  assign new_n1547_ = ~v6 & new_n1546_;
  assign new_n1548_ = v4 & new_n1547_;
  assign new_n1549_ = v2 & new_n1548_;
  assign new_n1550_ = ~v0 & new_n1549_;
  assign new_n1551_ = ~new_n1536_ & ~new_n1550_;
  assign new_n1552_ = v9 & ~new_n1551_;
  assign new_n1553_ = new_n117_ & new_n319_;
  assign new_n1554_ = v6 & ~v19;
  assign new_n1555_ = v5 & new_n1554_;
  assign new_n1556_ = new_n397_ & new_n1555_;
  assign new_n1557_ = ~new_n1553_ & ~new_n1556_;
  assign new_n1558_ = v24 & ~new_n1557_;
  assign new_n1559_ = ~v10 & new_n1558_;
  assign new_n1560_ = ~v3 & new_n1559_;
  assign new_n1561_ = ~v1 & new_n1560_;
  assign new_n1562_ = new_n255_ & new_n853_;
  assign new_n1563_ = v10 & ~v24;
  assign new_n1564_ = new_n546_ & new_n1563_;
  assign new_n1565_ = new_n1562_ & new_n1564_;
  assign new_n1566_ = ~new_n1561_ & ~new_n1565_;
  assign new_n1567_ = ~v25 & ~new_n1566_;
  assign new_n1568_ = new_n117_ & new_n1409_;
  assign new_n1569_ = new_n116_ & new_n1568_;
  assign new_n1570_ = ~new_n1567_ & ~new_n1569_;
  assign new_n1571_ = ~v9 & ~new_n1570_;
  assign new_n1572_ = ~v8 & new_n1571_;
  assign new_n1573_ = ~v0 & new_n1572_;
  assign new_n1574_ = ~new_n1552_ & ~new_n1573_;
  assign new_n1575_ = ~v7 & ~new_n1574_;
  assign new_n1576_ = ~new_n1503_ & ~new_n1575_;
  assign new_n1577_ = ~v23 & ~new_n1576_;
  assign new_n1578_ = ~v3 & new_n475_;
  assign new_n1579_ = ~v0 & new_n1578_;
  assign new_n1580_ = new_n481_ & new_n1436_;
  assign new_n1581_ = ~new_n1579_ & ~new_n1580_;
  assign new_n1582_ = ~v1 & ~new_n1581_;
  assign new_n1583_ = ~new_n490_ & ~new_n1582_;
  assign new_n1584_ = v2 & ~new_n1583_;
  assign new_n1585_ = ~v3 & new_n488_;
  assign new_n1586_ = ~v2 & new_n1585_;
  assign new_n1587_ = v0 & new_n1586_;
  assign new_n1588_ = ~new_n1584_ & ~new_n1587_;
  assign new_n1589_ = v7 & ~new_n1588_;
  assign new_n1590_ = ~v3 & new_n501_;
  assign new_n1591_ = ~v1 & new_n1590_;
  assign new_n1592_ = ~v0 & new_n1591_;
  assign new_n1593_ = ~new_n1589_ & ~new_n1592_;
  assign new_n1594_ = ~v25 & ~new_n1593_;
  assign new_n1595_ = v23 & new_n1594_;
  assign new_n1596_ = ~v8 & new_n1595_;
  assign new_n1597_ = ~new_n1577_ & ~new_n1596_;
  assign \v26.16  = ~v22 & ~new_n1597_;
  assign new_n1599_ = ~v10 & v23;
  assign new_n1600_ = v6 & new_n1599_;
  assign new_n1601_ = v0 & new_n1600_;
  assign new_n1602_ = new_n95_ & new_n1308_;
  assign new_n1603_ = ~new_n1601_ & ~new_n1602_;
  assign new_n1604_ = ~v9 & ~new_n1603_;
  assign new_n1605_ = ~v1 & ~v6;
  assign new_n1606_ = ~v0 & new_n1605_;
  assign new_n1607_ = v9 & new_n1163_;
  assign new_n1608_ = new_n1606_ & new_n1607_;
  assign new_n1609_ = ~new_n1604_ & ~new_n1608_;
  assign new_n1610_ = ~v24 & ~new_n1609_;
  assign new_n1611_ = ~v4 & new_n1610_;
  assign new_n1612_ = v6 & v10;
  assign new_n1613_ = v6 & ~new_n1612_;
  assign new_n1614_ = v24 & ~new_n1613_;
  assign new_n1615_ = ~v23 & new_n1614_;
  assign new_n1616_ = v9 & new_n1615_;
  assign new_n1617_ = v4 & new_n1616_;
  assign new_n1618_ = v1 & new_n1617_;
  assign new_n1619_ = ~v0 & new_n1618_;
  assign new_n1620_ = ~new_n1611_ & ~new_n1619_;
  assign new_n1621_ = v2 & ~new_n1620_;
  assign new_n1622_ = v6 & new_n729_;
  assign new_n1623_ = v4 & new_n1622_;
  assign new_n1624_ = ~v2 & new_n1623_;
  assign new_n1625_ = v1 & new_n1624_;
  assign new_n1626_ = v0 & new_n1625_;
  assign new_n1627_ = ~new_n1621_ & ~new_n1626_;
  assign new_n1628_ = v25 & ~new_n1627_;
  assign new_n1629_ = v0 & v2;
  assign new_n1630_ = v6 & new_n398_;
  assign new_n1631_ = new_n1629_ & new_n1630_;
  assign new_n1632_ = ~v6 & new_n118_;
  assign new_n1633_ = new_n1009_ & new_n1632_;
  assign new_n1634_ = ~new_n1631_ & ~new_n1633_;
  assign new_n1635_ = ~v24 & ~new_n1634_;
  assign new_n1636_ = v4 & new_n1635_;
  assign new_n1637_ = ~v6 & new_n258_;
  assign new_n1638_ = ~v4 & new_n1637_;
  assign new_n1639_ = v2 & new_n1638_;
  assign new_n1640_ = ~v0 & new_n1639_;
  assign new_n1641_ = ~new_n1636_ & ~new_n1640_;
  assign new_n1642_ = ~v25 & ~new_n1641_;
  assign new_n1643_ = ~v23 & new_n1642_;
  assign new_n1644_ = ~v1 & new_n1643_;
  assign new_n1645_ = ~new_n1628_ & ~new_n1644_;
  assign new_n1646_ = ~v8 & ~new_n1645_;
  assign new_n1647_ = v8 & new_n1213_;
  assign new_n1648_ = v6 & new_n1647_;
  assign new_n1649_ = v4 & new_n1648_;
  assign new_n1650_ = ~v2 & new_n1649_;
  assign new_n1651_ = v1 & new_n1650_;
  assign new_n1652_ = v0 & new_n1651_;
  assign new_n1653_ = ~new_n1646_ & ~new_n1652_;
  assign new_n1654_ = v7 & ~new_n1653_;
  assign new_n1655_ = ~v8 & new_n384_;
  assign new_n1656_ = v2 & new_n1655_;
  assign new_n1657_ = v1 & new_n1656_;
  assign new_n1658_ = ~v1 & new_n361_;
  assign new_n1659_ = new_n194_ & new_n321_;
  assign new_n1660_ = new_n1658_ & new_n1659_;
  assign new_n1661_ = ~new_n1657_ & ~new_n1660_;
  assign new_n1662_ = ~v10 & ~new_n1661_;
  assign new_n1663_ = new_n334_ & new_n382_;
  assign new_n1664_ = new_n200_ & new_n398_;
  assign new_n1665_ = new_n1663_ & new_n1664_;
  assign new_n1666_ = ~new_n1662_ & ~new_n1665_;
  assign new_n1667_ = ~v23 & ~new_n1666_;
  assign new_n1668_ = ~v7 & new_n1667_;
  assign new_n1669_ = v4 & new_n1668_;
  assign new_n1670_ = ~v0 & new_n1669_;
  assign new_n1671_ = ~new_n1654_ & ~new_n1670_;
  assign new_n1672_ = v3 & ~new_n1671_;
  assign new_n1673_ = ~v23 & ~new_n363_;
  assign new_n1674_ = v9 & new_n1673_;
  assign new_n1675_ = ~v0 & new_n1674_;
  assign new_n1676_ = new_n368_ & new_n1599_;
  assign new_n1677_ = new_n367_ & new_n1676_;
  assign new_n1678_ = ~new_n1675_ & ~new_n1677_;
  assign new_n1679_ = ~v1 & ~new_n1678_;
  assign new_n1680_ = ~v9 & new_n1599_;
  assign new_n1681_ = ~v8 & new_n1680_;
  assign new_n1682_ = v6 & new_n1681_;
  assign new_n1683_ = v1 & new_n1682_;
  assign new_n1684_ = v0 & new_n1683_;
  assign new_n1685_ = ~new_n1679_ & ~new_n1684_;
  assign new_n1686_ = v25 & ~new_n1685_;
  assign new_n1687_ = ~v24 & new_n1686_;
  assign new_n1688_ = v7 & new_n1687_;
  assign new_n1689_ = ~v4 & new_n1688_;
  assign new_n1690_ = ~v3 & new_n1689_;
  assign new_n1691_ = ~new_n1672_ & ~new_n1690_;
  assign new_n1692_ = ~v5 & ~new_n1691_;
  assign new_n1693_ = v3 & ~v25;
  assign new_n1694_ = v1 & new_n1693_;
  assign new_n1695_ = new_n589_ & new_n856_;
  assign new_n1696_ = ~new_n1694_ & ~new_n1695_;
  assign new_n1697_ = ~v7 & ~new_n1696_;
  assign new_n1698_ = v7 & new_n856_;
  assign new_n1699_ = new_n589_ & new_n1698_;
  assign new_n1700_ = ~new_n1697_ & ~new_n1699_;
  assign new_n1701_ = ~v6 & ~new_n1700_;
  assign new_n1702_ = v3 & v6;
  assign new_n1703_ = v1 & new_n1702_;
  assign new_n1704_ = ~v7 & new_n322_;
  assign new_n1705_ = new_n1703_ & new_n1704_;
  assign new_n1706_ = ~new_n1701_ & ~new_n1705_;
  assign new_n1707_ = v24 & ~new_n1706_;
  assign new_n1708_ = v2 & new_n1707_;
  assign new_n1709_ = ~v3 & v6;
  assign new_n1710_ = new_n853_ & new_n1709_;
  assign new_n1711_ = new_n923_ & new_n1710_;
  assign new_n1712_ = ~new_n1708_ & ~new_n1711_;
  assign new_n1713_ = ~v23 & ~new_n1712_;
  assign new_n1714_ = v9 & new_n1713_;
  assign new_n1715_ = ~v8 & new_n1714_;
  assign new_n1716_ = v5 & new_n1715_;
  assign new_n1717_ = v4 & new_n1716_;
  assign new_n1718_ = ~v0 & new_n1717_;
  assign new_n1719_ = ~new_n1692_ & ~new_n1718_;
  assign \v26.17  = ~v22 & ~new_n1719_;
  assign new_n1721_ = v3 & ~v6;
  assign new_n1722_ = new_n359_ & new_n1721_;
  assign new_n1723_ = new_n545_ & new_n1722_;
  assign new_n1724_ = v0 & new_n853_;
  assign new_n1725_ = new_n239_ & new_n1709_;
  assign new_n1726_ = new_n1724_ & new_n1725_;
  assign new_n1727_ = ~new_n1723_ & ~new_n1726_;
  assign new_n1728_ = ~v25 & ~new_n1727_;
  assign new_n1729_ = ~v4 & new_n1728_;
  assign new_n1730_ = v6 & v25;
  assign new_n1731_ = v4 & new_n1730_;
  assign new_n1732_ = v3 & new_n1731_;
  assign new_n1733_ = ~v2 & new_n1732_;
  assign new_n1734_ = v1 & new_n1733_;
  assign new_n1735_ = v0 & new_n1734_;
  assign new_n1736_ = ~new_n1729_ & ~new_n1735_;
  assign new_n1737_ = ~v2 & ~v8;
  assign new_n1738_ = ~v2 & ~new_n1737_;
  assign new_n1739_ = ~v25 & ~new_n1738_;
  assign new_n1740_ = ~v10 & new_n1739_;
  assign new_n1741_ = ~v9 & new_n1740_;
  assign new_n1742_ = v6 & new_n1741_;
  assign new_n1743_ = ~v4 & new_n1742_;
  assign new_n1744_ = ~v3 & new_n1743_;
  assign new_n1745_ = v1 & new_n1744_;
  assign new_n1746_ = v0 & new_n1745_;
  assign new_n1747_ = new_n1736_ & ~new_n1746_;
  assign new_n1748_ = v24 & ~new_n1747_;
  assign new_n1749_ = v2 & new_n1422_;
  assign new_n1750_ = v0 & new_n1749_;
  assign new_n1751_ = ~v8 & new_n298_;
  assign new_n1752_ = new_n1009_ & new_n1751_;
  assign new_n1753_ = ~new_n1750_ & ~new_n1752_;
  assign new_n1754_ = ~v1 & ~new_n1753_;
  assign new_n1755_ = ~v2 & ~new_n302_;
  assign new_n1756_ = v1 & new_n1755_;
  assign new_n1757_ = ~v0 & new_n1756_;
  assign new_n1758_ = ~new_n1754_ & ~new_n1757_;
  assign new_n1759_ = v4 & ~new_n1758_;
  assign new_n1760_ = ~v9 & new_n658_;
  assign new_n1761_ = ~v4 & new_n1760_;
  assign new_n1762_ = ~v1 & new_n1761_;
  assign new_n1763_ = v0 & new_n1762_;
  assign new_n1764_ = ~new_n1759_ & ~new_n1763_;
  assign new_n1765_ = v3 & ~new_n1764_;
  assign new_n1766_ = ~v0 & new_n310_;
  assign new_n1767_ = v0 & new_n368_;
  assign new_n1768_ = ~new_n1766_ & ~new_n1767_;
  assign new_n1769_ = ~v10 & ~new_n1768_;
  assign new_n1770_ = ~v4 & new_n1769_;
  assign new_n1771_ = ~v3 & new_n1770_;
  assign new_n1772_ = ~v2 & new_n1771_;
  assign new_n1773_ = ~v1 & new_n1772_;
  assign new_n1774_ = ~new_n1765_ & ~new_n1773_;
  assign new_n1775_ = v25 & ~new_n1774_;
  assign new_n1776_ = ~v24 & new_n1775_;
  assign new_n1777_ = v6 & new_n1776_;
  assign new_n1778_ = ~new_n1748_ & ~new_n1777_;
  assign new_n1779_ = v7 & ~new_n1778_;
  assign new_n1780_ = new_n187_ & new_n593_;
  assign new_n1781_ = new_n188_ & new_n277_;
  assign new_n1782_ = ~new_n1780_ & ~new_n1781_;
  assign new_n1783_ = v9 & ~new_n1782_;
  assign new_n1784_ = v8 & new_n1783_;
  assign new_n1785_ = v6 & new_n1784_;
  assign new_n1786_ = v0 & new_n1785_;
  assign new_n1787_ = new_n95_ & new_n713_;
  assign new_n1788_ = ~v9 & new_n200_;
  assign new_n1789_ = new_n382_ & new_n1788_;
  assign new_n1790_ = new_n1787_ & new_n1789_;
  assign new_n1791_ = ~new_n1786_ & ~new_n1790_;
  assign new_n1792_ = ~v10 & ~new_n1791_;
  assign new_n1793_ = ~v7 & new_n1792_;
  assign new_n1794_ = ~v4 & new_n1793_;
  assign new_n1795_ = ~new_n1779_ & ~new_n1794_;
  assign new_n1796_ = ~v5 & ~new_n1795_;
  assign new_n1797_ = v7 & ~new_n386_;
  assign new_n1798_ = ~v3 & new_n148_;
  assign new_n1799_ = new_n200_ & new_n257_;
  assign new_n1800_ = new_n1798_ & new_n1799_;
  assign new_n1801_ = ~new_n1797_ & ~new_n1800_;
  assign new_n1802_ = v10 & ~new_n1801_;
  assign new_n1803_ = new_n1125_ & new_n1709_;
  assign new_n1804_ = ~v19 & new_n188_;
  assign new_n1805_ = new_n118_ & new_n1804_;
  assign new_n1806_ = new_n1803_ & new_n1805_;
  assign new_n1807_ = ~new_n1802_ & ~new_n1806_;
  assign new_n1808_ = v4 & ~new_n1807_;
  assign new_n1809_ = ~v1 & new_n1808_;
  assign new_n1810_ = ~v0 & new_n1809_;
  assign new_n1811_ = ~v3 & new_n991_;
  assign new_n1812_ = new_n289_ & new_n1811_;
  assign new_n1813_ = v7 & new_n310_;
  assign new_n1814_ = ~v10 & new_n188_;
  assign new_n1815_ = new_n1813_ & new_n1814_;
  assign new_n1816_ = new_n1812_ & new_n1815_;
  assign new_n1817_ = ~new_n1810_ & ~new_n1816_;
  assign new_n1818_ = v5 & ~new_n1817_;
  assign new_n1819_ = v2 & new_n1818_;
  assign new_n1820_ = ~new_n1796_ & ~new_n1819_;
  assign new_n1821_ = ~v23 & ~new_n1820_;
  assign new_n1822_ = new_n115_ & new_n117_;
  assign new_n1823_ = new_n235_ & new_n1822_;
  assign new_n1824_ = ~v7 & new_n368_;
  assign new_n1825_ = new_n194_ & new_n1599_;
  assign new_n1826_ = new_n1824_ & new_n1825_;
  assign new_n1827_ = new_n1823_ & new_n1826_;
  assign new_n1828_ = ~new_n1821_ & ~new_n1827_;
  assign \v26.18  = ~v22 & ~new_n1828_;
  assign new_n1830_ = v4 & new_n194_;
  assign new_n1831_ = v3 & new_n1830_;
  assign new_n1832_ = new_n115_ & new_n1409_;
  assign new_n1833_ = ~new_n1831_ & ~new_n1832_;
  assign new_n1834_ = v6 & ~new_n1833_;
  assign new_n1835_ = ~v5 & new_n1834_;
  assign new_n1836_ = v1 & new_n1835_;
  assign new_n1837_ = v0 & new_n1836_;
  assign new_n1838_ = new_n95_ & new_n237_;
  assign new_n1839_ = ~v6 & ~v10;
  assign new_n1840_ = new_n241_ & new_n1839_;
  assign new_n1841_ = new_n1838_ & new_n1840_;
  assign new_n1842_ = ~new_n1837_ & ~new_n1841_;
  assign new_n1843_ = v8 & ~new_n1842_;
  assign new_n1844_ = ~v8 & new_n194_;
  assign new_n1845_ = v6 & new_n1844_;
  assign new_n1846_ = ~v5 & new_n1845_;
  assign new_n1847_ = v4 & new_n1846_;
  assign new_n1848_ = v3 & new_n1847_;
  assign new_n1849_ = v1 & new_n1848_;
  assign new_n1850_ = v0 & new_n1849_;
  assign new_n1851_ = ~new_n1843_ & ~new_n1850_;
  assign new_n1852_ = ~v3 & new_n327_;
  assign new_n1853_ = v3 & new_n328_;
  assign new_n1854_ = ~new_n1852_ & ~new_n1853_;
  assign new_n1855_ = v24 & ~new_n1854_;
  assign new_n1856_ = v0 & new_n1855_;
  assign new_n1857_ = ~v0 & v3;
  assign new_n1858_ = new_n976_ & new_n1857_;
  assign new_n1859_ = ~new_n1856_ & ~new_n1858_;
  assign new_n1860_ = v6 & ~new_n1859_;
  assign new_n1861_ = ~v4 & new_n1860_;
  assign new_n1862_ = ~v0 & new_n255_;
  assign new_n1863_ = new_n194_ & new_n382_;
  assign new_n1864_ = new_n1862_ & new_n1863_;
  assign new_n1865_ = ~new_n1861_ & ~new_n1864_;
  assign new_n1866_ = ~v1 & ~new_n1865_;
  assign new_n1867_ = new_n115_ & new_n289_;
  assign new_n1868_ = new_n200_ & new_n1437_;
  assign new_n1869_ = new_n1867_ & new_n1868_;
  assign new_n1870_ = ~new_n1866_ & ~new_n1869_;
  assign new_n1871_ = ~v10 & ~new_n1870_;
  assign new_n1872_ = ~v9 & new_n1871_;
  assign new_n1873_ = ~v5 & new_n1872_;
  assign new_n1874_ = new_n1851_ & ~new_n1873_;
  assign new_n1875_ = ~v2 & ~new_n1874_;
  assign new_n1876_ = new_n236_ & new_n277_;
  assign new_n1877_ = new_n200_ & new_n239_;
  assign new_n1878_ = new_n1876_ & new_n1877_;
  assign new_n1879_ = new_n450_ & new_n593_;
  assign new_n1880_ = new_n194_ & new_n359_;
  assign new_n1881_ = new_n1879_ & new_n1880_;
  assign new_n1882_ = ~new_n1878_ & ~new_n1881_;
  assign new_n1883_ = v9 & ~new_n1882_;
  assign new_n1884_ = ~v1 & ~new_n329_;
  assign new_n1885_ = v1 & new_n327_;
  assign new_n1886_ = ~new_n1884_ & ~new_n1885_;
  assign new_n1887_ = v3 & ~new_n1886_;
  assign new_n1888_ = ~v3 & v25;
  assign new_n1889_ = v1 & new_n1888_;
  assign new_n1890_ = ~new_n1887_ & ~new_n1889_;
  assign new_n1891_ = v24 & ~new_n1890_;
  assign new_n1892_ = ~v10 & new_n1891_;
  assign new_n1893_ = ~v9 & new_n1892_;
  assign new_n1894_ = ~v5 & new_n1893_;
  assign new_n1895_ = ~v4 & new_n1894_;
  assign new_n1896_ = ~new_n1883_ & ~new_n1895_;
  assign new_n1897_ = v6 & ~new_n1896_;
  assign new_n1898_ = v2 & new_n1897_;
  assign new_n1899_ = v0 & new_n1898_;
  assign new_n1900_ = ~new_n1875_ & ~new_n1899_;
  assign new_n1901_ = v7 & ~new_n1900_;
  assign new_n1902_ = ~v4 & new_n263_;
  assign new_n1903_ = v0 & new_n1902_;
  assign new_n1904_ = v4 & new_n1039_;
  assign new_n1905_ = new_n1009_ & new_n1904_;
  assign new_n1906_ = ~new_n1903_ & ~new_n1905_;
  assign new_n1907_ = v8 & ~new_n1906_;
  assign new_n1908_ = v6 & new_n1907_;
  assign new_n1909_ = v3 & new_n1908_;
  assign new_n1910_ = new_n115_ & new_n1009_;
  assign new_n1911_ = new_n382_ & new_n1039_;
  assign new_n1912_ = new_n1910_ & new_n1911_;
  assign new_n1913_ = ~new_n1909_ & ~new_n1912_;
  assign new_n1914_ = ~v25 & ~new_n1913_;
  assign new_n1915_ = ~v1 & new_n1914_;
  assign new_n1916_ = v8 & new_n384_;
  assign new_n1917_ = v6 & new_n1916_;
  assign new_n1918_ = ~v4 & new_n1917_;
  assign new_n1919_ = ~v3 & new_n1918_;
  assign new_n1920_ = v1 & new_n1919_;
  assign new_n1921_ = v0 & new_n1920_;
  assign new_n1922_ = ~new_n1915_ & ~new_n1921_;
  assign new_n1923_ = ~v5 & ~new_n1922_;
  assign new_n1924_ = ~v2 & new_n725_;
  assign new_n1925_ = new_n254_ & new_n1924_;
  assign new_n1926_ = v5 & new_n1437_;
  assign new_n1927_ = new_n1255_ & new_n1926_;
  assign new_n1928_ = new_n1925_ & new_n1927_;
  assign new_n1929_ = ~new_n1923_ & ~new_n1928_;
  assign new_n1930_ = ~v10 & ~new_n1929_;
  assign new_n1931_ = ~v7 & new_n1930_;
  assign new_n1932_ = ~new_n1901_ & ~new_n1931_;
  assign new_n1933_ = ~v23 & ~new_n1932_;
  assign \v26.19  = ~v22 & new_n1933_;
  assign new_n1935_ = v6 & new_n359_;
  assign new_n1936_ = new_n451_ & new_n1935_;
  assign new_n1937_ = ~v6 & v8;
  assign new_n1938_ = new_n1347_ & new_n1937_;
  assign new_n1939_ = new_n237_ & new_n1938_;
  assign new_n1940_ = ~new_n1936_ & ~new_n1939_;
  assign new_n1941_ = ~v9 & ~new_n1940_;
  assign new_n1942_ = ~v1 & new_n1941_;
  assign new_n1943_ = v1 & v3;
  assign new_n1944_ = new_n450_ & new_n1943_;
  assign new_n1945_ = new_n300_ & new_n1437_;
  assign new_n1946_ = new_n1944_ & new_n1945_;
  assign new_n1947_ = ~new_n1942_ & ~new_n1946_;
  assign new_n1948_ = ~v24 & ~new_n1947_;
  assign new_n1949_ = ~v2 & new_n1948_;
  assign new_n1950_ = v9 & new_n1614_;
  assign new_n1951_ = ~v8 & new_n1950_;
  assign new_n1952_ = ~v5 & new_n1951_;
  assign new_n1953_ = v4 & new_n1952_;
  assign new_n1954_ = v3 & new_n1953_;
  assign new_n1955_ = v2 & new_n1954_;
  assign new_n1956_ = v1 & new_n1955_;
  assign new_n1957_ = ~new_n1949_ & ~new_n1956_;
  assign new_n1958_ = v7 & ~new_n1957_;
  assign new_n1959_ = v24 & ~new_n931_;
  assign new_n1960_ = v9 & new_n1959_;
  assign new_n1961_ = ~v8 & new_n1960_;
  assign new_n1962_ = ~v7 & new_n1961_;
  assign new_n1963_ = v4 & new_n1962_;
  assign new_n1964_ = v3 & new_n1963_;
  assign new_n1965_ = v2 & new_n1964_;
  assign new_n1966_ = v1 & new_n1965_;
  assign new_n1967_ = ~new_n1958_ & ~new_n1966_;
  assign new_n1968_ = v25 & ~new_n1967_;
  assign new_n1969_ = v24 & new_n84_;
  assign new_n1970_ = v9 & new_n1969_;
  assign new_n1971_ = ~v8 & new_n1970_;
  assign new_n1972_ = v4 & new_n1971_;
  assign new_n1973_ = v3 & new_n1972_;
  assign new_n1974_ = v2 & new_n1973_;
  assign new_n1975_ = v1 & new_n1974_;
  assign new_n1976_ = ~new_n1968_ & ~new_n1975_;
  assign new_n1977_ = ~v0 & ~new_n1976_;
  assign new_n1978_ = ~new_n249_ & ~new_n835_;
  assign new_n1979_ = v8 & new_n1978_;
  assign new_n1980_ = ~v9 & v24;
  assign new_n1981_ = ~v8 & new_n1980_;
  assign new_n1982_ = ~v3 & v7;
  assign new_n1983_ = v1 & new_n1982_;
  assign new_n1984_ = new_n1981_ & new_n1983_;
  assign new_n1985_ = ~new_n1979_ & ~new_n1984_;
  assign new_n1986_ = ~v24 & ~new_n714_;
  assign new_n1987_ = ~v9 & new_n1986_;
  assign new_n1988_ = ~v8 & new_n1987_;
  assign new_n1989_ = ~v1 & new_n1988_;
  assign new_n1990_ = v1 & new_n713_;
  assign new_n1991_ = v8 & new_n263_;
  assign new_n1992_ = new_n1990_ & new_n1991_;
  assign new_n1993_ = ~new_n1989_ & ~new_n1992_;
  assign new_n1994_ = v7 & ~new_n1993_;
  assign new_n1995_ = new_n1985_ & ~new_n1994_;
  assign new_n1996_ = ~v5 & ~new_n1995_;
  assign new_n1997_ = new_n145_ & new_n334_;
  assign new_n1998_ = new_n263_ & new_n882_;
  assign new_n1999_ = new_n1997_ & new_n1998_;
  assign new_n2000_ = ~new_n1996_ & ~new_n1999_;
  assign new_n2001_ = ~v25 & ~new_n2000_;
  assign new_n2002_ = ~v10 & new_n2001_;
  assign new_n2003_ = v6 & new_n2002_;
  assign new_n2004_ = ~v4 & new_n2003_;
  assign new_n2005_ = v0 & new_n2004_;
  assign new_n2006_ = ~new_n1977_ & ~new_n2005_;
  assign new_n2007_ = ~v23 & ~new_n2006_;
  assign new_n2008_ = ~new_n1827_ & ~new_n2007_;
  assign \v26.20  = ~v22 & ~new_n2008_;
  assign new_n2010_ = v4 & new_n1334_;
  assign new_n2011_ = ~v0 & new_n2010_;
  assign new_n2012_ = v0 & new_n991_;
  assign new_n2013_ = v8 & v25;
  assign new_n2014_ = v7 & new_n2013_;
  assign new_n2015_ = new_n2012_ & new_n2014_;
  assign new_n2016_ = ~new_n2011_ & ~new_n2015_;
  assign new_n2017_ = ~v2 & ~new_n2016_;
  assign new_n2018_ = v7 & v25;
  assign new_n2019_ = v6 & new_n2018_;
  assign new_n2020_ = ~v4 & new_n2019_;
  assign new_n2021_ = v2 & new_n2020_;
  assign new_n2022_ = v0 & new_n2021_;
  assign new_n2023_ = ~new_n2017_ & ~new_n2022_;
  assign new_n2024_ = ~v23 & ~new_n2023_;
  assign new_n2025_ = ~v8 & v23;
  assign new_n2026_ = v7 & new_n2025_;
  assign new_n2027_ = v6 & new_n2026_;
  assign new_n2028_ = ~v4 & new_n2027_;
  assign new_n2029_ = v2 & new_n2028_;
  assign new_n2030_ = v0 & new_n2029_;
  assign new_n2031_ = ~new_n2024_ & ~new_n2030_;
  assign new_n2032_ = v3 & ~new_n2031_;
  assign new_n2033_ = ~v23 & ~new_n129_;
  assign new_n2034_ = ~v8 & ~new_n2033_;
  assign new_n2035_ = v7 & new_n2034_;
  assign new_n2036_ = v6 & new_n2035_;
  assign new_n2037_ = ~v4 & new_n2036_;
  assign new_n2038_ = ~v3 & new_n2037_;
  assign new_n2039_ = ~v2 & new_n2038_;
  assign new_n2040_ = v0 & new_n2039_;
  assign new_n2041_ = ~new_n2032_ & ~new_n2040_;
  assign new_n2042_ = ~v1 & ~new_n2041_;
  assign new_n2043_ = v23 & ~new_n1359_;
  assign new_n2044_ = ~v8 & new_n2043_;
  assign new_n2045_ = v7 & new_n2044_;
  assign new_n2046_ = v6 & new_n2045_;
  assign new_n2047_ = ~v4 & new_n2046_;
  assign new_n2048_ = v1 & new_n2047_;
  assign new_n2049_ = v0 & new_n2048_;
  assign new_n2050_ = ~new_n2042_ & ~new_n2049_;
  assign new_n2051_ = ~v9 & ~new_n2050_;
  assign new_n2052_ = v9 & new_n129_;
  assign new_n2053_ = v8 & new_n2052_;
  assign new_n2054_ = ~v7 & new_n2053_;
  assign new_n2055_ = v6 & new_n2054_;
  assign new_n2056_ = ~v4 & new_n2055_;
  assign new_n2057_ = v3 & new_n2056_;
  assign new_n2058_ = ~v1 & new_n2057_;
  assign new_n2059_ = v0 & new_n2058_;
  assign new_n2060_ = ~new_n2051_ & ~new_n2059_;
  assign new_n2061_ = ~v10 & ~new_n2060_;
  assign new_n2062_ = v10 & new_n129_;
  assign new_n2063_ = ~v8 & new_n2062_;
  assign new_n2064_ = v7 & new_n2063_;
  assign new_n2065_ = ~v6 & new_n2064_;
  assign new_n2066_ = ~v4 & new_n2065_;
  assign new_n2067_ = v3 & new_n2066_;
  assign new_n2068_ = v2 & new_n2067_;
  assign new_n2069_ = ~v1 & new_n2068_;
  assign new_n2070_ = ~v0 & new_n2069_;
  assign new_n2071_ = ~new_n2061_ & ~new_n2070_;
  assign new_n2072_ = ~v24 & ~new_n2071_;
  assign new_n2073_ = ~v22 & new_n2072_;
  assign \v26.21  = ~v5 & new_n2073_;
  assign new_n2075_ = v7 & new_n658_;
  assign new_n2076_ = ~v5 & new_n2075_;
  assign new_n2077_ = ~v4 & new_n2076_;
  assign new_n2078_ = ~v1 & new_n2077_;
  assign new_n2079_ = v0 & new_n2078_;
  assign new_n2080_ = new_n254_ & new_n346_;
  assign new_n2081_ = new_n73_ & new_n359_;
  assign new_n2082_ = new_n2080_ & new_n2081_;
  assign new_n2083_ = ~new_n2079_ & ~new_n2082_;
  assign new_n2084_ = ~v24 & ~new_n2083_;
  assign new_n2085_ = v4 & new_n767_;
  assign new_n2086_ = ~new_n1170_ & ~new_n2085_;
  assign new_n2087_ = v24 & ~new_n2086_;
  assign new_n2088_ = v7 & new_n2087_;
  assign new_n2089_ = v5 & new_n2088_;
  assign new_n2090_ = v2 & new_n2089_;
  assign new_n2091_ = ~v1 & new_n2090_;
  assign new_n2092_ = ~v0 & new_n2091_;
  assign new_n2093_ = ~new_n2084_ & ~new_n2092_;
  assign new_n2094_ = v3 & ~new_n2093_;
  assign new_n2095_ = v1 & v24;
  assign new_n2096_ = ~v8 & ~v24;
  assign new_n2097_ = new_n114_ & new_n2096_;
  assign new_n2098_ = ~new_n2095_ & ~new_n2097_;
  assign new_n2099_ = ~v10 & ~new_n2098_;
  assign new_n2100_ = v7 & new_n2099_;
  assign new_n2101_ = ~v5 & new_n2100_;
  assign new_n2102_ = ~v4 & new_n2101_;
  assign new_n2103_ = ~v3 & new_n2102_;
  assign new_n2104_ = v0 & new_n2103_;
  assign new_n2105_ = ~new_n2094_ & ~new_n2104_;
  assign new_n2106_ = ~v9 & ~new_n2105_;
  assign new_n2107_ = ~v7 & ~new_n249_;
  assign new_n2108_ = v7 & v24;
  assign new_n2109_ = ~v3 & new_n2108_;
  assign new_n2110_ = new_n853_ & new_n2109_;
  assign new_n2111_ = ~new_n2107_ & ~new_n2110_;
  assign new_n2112_ = ~v5 & ~new_n2111_;
  assign new_n2113_ = v5 & new_n2108_;
  assign new_n2114_ = new_n715_ & new_n2113_;
  assign new_n2115_ = ~new_n2112_ & ~new_n2114_;
  assign new_n2116_ = ~v10 & ~new_n2115_;
  assign new_n2117_ = v9 & new_n2116_;
  assign new_n2118_ = v8 & new_n2117_;
  assign new_n2119_ = ~v4 & new_n2118_;
  assign new_n2120_ = v0 & new_n2119_;
  assign new_n2121_ = ~new_n2106_ & ~new_n2120_;
  assign new_n2122_ = ~v25 & ~new_n2121_;
  assign new_n2123_ = v6 & new_n2122_;
  assign new_n2124_ = ~v10 & new_n241_;
  assign new_n2125_ = v8 & new_n2124_;
  assign new_n2126_ = v7 & new_n2125_;
  assign new_n2127_ = ~v6 & new_n2126_;
  assign new_n2128_ = v5 & new_n2127_;
  assign new_n2129_ = ~v4 & new_n2128_;
  assign new_n2130_ = ~v3 & new_n2129_;
  assign new_n2131_ = ~v2 & new_n2130_;
  assign new_n2132_ = ~v1 & new_n2131_;
  assign new_n2133_ = ~v0 & new_n2132_;
  assign new_n2134_ = ~new_n2123_ & ~new_n2133_;
  assign new_n2135_ = ~v23 & ~new_n2134_;
  assign new_n2136_ = v10 & new_n1282_;
  assign new_n2137_ = v9 & new_n2136_;
  assign new_n2138_ = ~v8 & new_n2137_;
  assign new_n2139_ = ~v6 & new_n2138_;
  assign new_n2140_ = v5 & new_n2139_;
  assign new_n2141_ = v4 & new_n2140_;
  assign new_n2142_ = ~v3 & new_n2141_;
  assign new_n2143_ = v2 & new_n2142_;
  assign new_n2144_ = ~v1 & new_n2143_;
  assign new_n2145_ = ~v0 & new_n2144_;
  assign new_n2146_ = ~new_n2135_ & ~new_n2145_;
  assign \v26.22  = ~v22 & ~new_n2146_;
  assign new_n2148_ = v3 & v25;
  assign new_n2149_ = v1 & new_n2148_;
  assign new_n2150_ = v5 & ~v25;
  assign new_n2151_ = new_n589_ & new_n2150_;
  assign new_n2152_ = ~new_n2149_ & ~new_n2151_;
  assign new_n2153_ = ~v7 & ~new_n2152_;
  assign new_n2154_ = v7 & ~v25;
  assign new_n2155_ = v5 & new_n2154_;
  assign new_n2156_ = new_n589_ & new_n2155_;
  assign new_n2157_ = ~new_n2153_ & ~new_n2156_;
  assign new_n2158_ = v4 & ~new_n2157_;
  assign new_n2159_ = ~new_n1693_ & ~new_n1888_;
  assign new_n2160_ = v7 & ~new_n2159_;
  assign new_n2161_ = ~v5 & new_n2160_;
  assign new_n2162_ = ~v4 & new_n2161_;
  assign new_n2163_ = ~v1 & new_n2162_;
  assign new_n2164_ = ~new_n2158_ & ~new_n2163_;
  assign new_n2165_ = ~v24 & ~new_n2164_;
  assign new_n2166_ = new_n200_ & new_n571_;
  assign new_n2167_ = new_n440_ & new_n2166_;
  assign new_n2168_ = ~new_n2165_ & ~new_n2167_;
  assign new_n2169_ = v9 & ~new_n2168_;
  assign new_n2170_ = v7 & new_n1487_;
  assign new_n2171_ = ~v5 & new_n2170_;
  assign new_n2172_ = ~v4 & new_n2171_;
  assign new_n2173_ = v3 & new_n2172_;
  assign new_n2174_ = ~v1 & new_n2173_;
  assign new_n2175_ = ~new_n2169_ & ~new_n2174_;
  assign new_n2176_ = v2 & ~new_n2175_;
  assign new_n2177_ = v7 & new_n1039_;
  assign new_n2178_ = v5 & new_n2177_;
  assign new_n2179_ = v4 & new_n2178_;
  assign new_n2180_ = ~v3 & new_n2179_;
  assign new_n2181_ = ~v2 & new_n2180_;
  assign new_n2182_ = ~v1 & new_n2181_;
  assign new_n2183_ = ~new_n2176_ & ~new_n2182_;
  assign new_n2184_ = v10 & ~new_n2183_;
  assign new_n2185_ = new_n612_ & new_n1406_;
  assign new_n2186_ = v3 & v5;
  assign new_n2187_ = new_n616_ & new_n2186_;
  assign new_n2188_ = ~new_n2185_ & ~new_n2187_;
  assign new_n2189_ = ~v24 & ~new_n2188_;
  assign new_n2190_ = ~v10 & new_n2189_;
  assign new_n2191_ = ~v7 & new_n2190_;
  assign new_n2192_ = ~v4 & new_n2191_;
  assign new_n2193_ = ~v2 & new_n2192_;
  assign new_n2194_ = ~v1 & new_n2193_;
  assign new_n2195_ = ~new_n2184_ & ~new_n2194_;
  assign new_n2196_ = ~v6 & ~new_n2195_;
  assign new_n2197_ = v5 & new_n830_;
  assign new_n2198_ = new_n1383_ & new_n2197_;
  assign new_n2199_ = ~v2 & new_n115_;
  assign new_n2200_ = ~v5 & new_n834_;
  assign new_n2201_ = new_n2199_ & new_n2200_;
  assign new_n2202_ = ~new_n2198_ & ~new_n2201_;
  assign new_n2203_ = ~v25 & ~new_n2202_;
  assign new_n2204_ = ~v24 & new_n2203_;
  assign new_n2205_ = v10 & new_n2204_;
  assign new_n2206_ = v6 & new_n2205_;
  assign new_n2207_ = ~v1 & new_n2206_;
  assign new_n2208_ = ~new_n2196_ & ~new_n2207_;
  assign new_n2209_ = ~v8 & ~new_n2208_;
  assign new_n2210_ = ~v1 & new_n136_;
  assign new_n2211_ = v4 & new_n117_;
  assign new_n2212_ = new_n2210_ & new_n2211_;
  assign new_n2213_ = v10 & new_n194_;
  assign new_n2214_ = new_n1118_ & new_n2213_;
  assign new_n2215_ = new_n2212_ & new_n2214_;
  assign new_n2216_ = ~new_n2209_ & ~new_n2215_;
  assign new_n2217_ = ~v23 & ~new_n2216_;
  assign new_n2218_ = ~v22 & new_n2217_;
  assign \v26.23  = ~v0 & new_n2218_;
  assign new_n2220_ = v4 & new_n187_;
  assign new_n2221_ = v3 & new_n2220_;
  assign new_n2222_ = new_n115_ & new_n1814_;
  assign new_n2223_ = ~new_n2221_ & ~new_n2222_;
  assign new_n2224_ = v6 & ~new_n2223_;
  assign new_n2225_ = ~v5 & new_n2224_;
  assign new_n2226_ = v1 & new_n2225_;
  assign new_n2227_ = v0 & new_n2226_;
  assign new_n2228_ = ~new_n1841_ & ~new_n2227_;
  assign new_n2229_ = v8 & ~new_n2228_;
  assign new_n2230_ = ~v8 & new_n187_;
  assign new_n2231_ = v6 & new_n2230_;
  assign new_n2232_ = ~v5 & new_n2231_;
  assign new_n2233_ = v4 & new_n2232_;
  assign new_n2234_ = v3 & new_n2233_;
  assign new_n2235_ = v1 & new_n2234_;
  assign new_n2236_ = v0 & new_n2235_;
  assign new_n2237_ = ~new_n2229_ & ~new_n2236_;
  assign new_n2238_ = new_n187_ & new_n767_;
  assign new_n2239_ = new_n1862_ & new_n2238_;
  assign new_n2240_ = v0 & new_n115_;
  assign new_n2241_ = new_n188_ & new_n347_;
  assign new_n2242_ = new_n2240_ & new_n2241_;
  assign new_n2243_ = ~new_n2239_ & ~new_n2242_;
  assign new_n2244_ = v1 & ~new_n2243_;
  assign new_n2245_ = ~v25 & ~new_n274_;
  assign new_n2246_ = ~v24 & new_n2245_;
  assign new_n2247_ = ~v10 & new_n2246_;
  assign new_n2248_ = ~v4 & new_n2247_;
  assign new_n2249_ = ~v1 & new_n2248_;
  assign new_n2250_ = v0 & new_n2249_;
  assign new_n2251_ = ~new_n2244_ & ~new_n2250_;
  assign new_n2252_ = ~v9 & ~new_n2251_;
  assign new_n2253_ = v6 & new_n2252_;
  assign new_n2254_ = ~v5 & new_n2253_;
  assign new_n2255_ = new_n2237_ & ~new_n2254_;
  assign new_n2256_ = ~v2 & ~new_n2255_;
  assign new_n2257_ = ~v25 & ~new_n249_;
  assign new_n2258_ = ~v4 & new_n2257_;
  assign new_n2259_ = ~v1 & new_n255_;
  assign new_n2260_ = new_n2230_ & new_n2259_;
  assign new_n2261_ = ~new_n2258_ & ~new_n2260_;
  assign new_n2262_ = ~v9 & ~new_n2261_;
  assign new_n2263_ = new_n187_ & new_n310_;
  assign new_n2264_ = new_n2259_ & new_n2263_;
  assign new_n2265_ = ~new_n2262_ & ~new_n2264_;
  assign new_n2266_ = ~v5 & ~new_n2265_;
  assign new_n2267_ = new_n188_ & new_n310_;
  assign new_n2268_ = new_n1876_ & new_n2267_;
  assign new_n2269_ = ~new_n2266_ & ~new_n2268_;
  assign new_n2270_ = ~v10 & ~new_n2269_;
  assign new_n2271_ = v6 & new_n2270_;
  assign new_n2272_ = v0 & new_n2271_;
  assign new_n2273_ = ~v3 & new_n479_;
  assign new_n2274_ = new_n95_ & new_n2273_;
  assign new_n2275_ = ~v6 & new_n257_;
  assign new_n2276_ = new_n953_ & new_n2275_;
  assign new_n2277_ = new_n2274_ & new_n2276_;
  assign new_n2278_ = ~new_n2272_ & ~new_n2277_;
  assign new_n2279_ = v2 & ~new_n2278_;
  assign new_n2280_ = ~new_n2256_ & ~new_n2279_;
  assign new_n2281_ = v7 & ~new_n2280_;
  assign new_n2282_ = v8 & ~new_n249_;
  assign new_n2283_ = v6 & new_n2282_;
  assign new_n2284_ = ~v5 & new_n2283_;
  assign new_n2285_ = v0 & new_n2284_;
  assign new_n2286_ = new_n138_ & new_n2096_;
  assign new_n2287_ = new_n594_ & new_n2286_;
  assign new_n2288_ = ~new_n2285_ & ~new_n2287_;
  assign new_n2289_ = ~v10 & ~new_n2288_;
  assign new_n2290_ = v9 & new_n2289_;
  assign new_n2291_ = ~v4 & new_n2290_;
  assign new_n2292_ = v3 & new_n419_;
  assign new_n2293_ = new_n254_ & new_n2292_;
  assign new_n2294_ = ~v9 & new_n1563_;
  assign new_n2295_ = new_n1437_ & new_n2294_;
  assign new_n2296_ = new_n2293_ & new_n2295_;
  assign new_n2297_ = ~new_n2291_ & ~new_n2296_;
  assign new_n2298_ = ~v2 & ~new_n2297_;
  assign new_n2299_ = v9 & new_n250_;
  assign new_n2300_ = v8 & new_n2299_;
  assign new_n2301_ = v6 & new_n2300_;
  assign new_n2302_ = ~v5 & new_n2301_;
  assign new_n2303_ = ~v4 & new_n2302_;
  assign new_n2304_ = v2 & new_n2303_;
  assign new_n2305_ = v0 & new_n2304_;
  assign new_n2306_ = ~new_n2298_ & ~new_n2305_;
  assign new_n2307_ = ~v25 & ~new_n2306_;
  assign new_n2308_ = ~v7 & new_n2307_;
  assign new_n2309_ = ~new_n2281_ & ~new_n2308_;
  assign new_n2310_ = ~v23 & ~new_n2309_;
  assign new_n2311_ = v10 & new_n791_;
  assign new_n2312_ = v9 & new_n2311_;
  assign new_n2313_ = ~v8 & new_n2312_;
  assign new_n2314_ = ~v6 & new_n2313_;
  assign new_n2315_ = v5 & new_n2314_;
  assign new_n2316_ = v4 & new_n2315_;
  assign new_n2317_ = ~v3 & new_n2316_;
  assign new_n2318_ = v2 & new_n2317_;
  assign new_n2319_ = ~v1 & new_n2318_;
  assign new_n2320_ = ~v0 & new_n2319_;
  assign new_n2321_ = ~new_n2310_ & ~new_n2320_;
  assign \v26.24  = ~v22 & ~new_n2321_;
  assign new_n2323_ = ~v2 & new_n533_;
  assign new_n2324_ = v0 & new_n2323_;
  assign new_n2325_ = ~v6 & new_n547_;
  assign new_n2326_ = new_n537_ & new_n2325_;
  assign new_n2327_ = ~new_n2324_ & ~new_n2326_;
  assign new_n2328_ = ~v5 & ~new_n2327_;
  assign new_n2329_ = v2 & v5;
  assign new_n2330_ = ~v0 & new_n2329_;
  assign new_n2331_ = new_n2325_ & new_n2330_;
  assign new_n2332_ = ~new_n2328_ & ~new_n2331_;
  assign new_n2333_ = v25 & ~new_n2332_;
  assign new_n2334_ = ~v23 & new_n2333_;
  assign new_n2335_ = v3 & new_n2334_;
  assign new_n2336_ = v1 & new_n2335_;
  assign new_n2337_ = ~v6 & new_n140_;
  assign new_n2338_ = v5 & new_n2337_;
  assign new_n2339_ = ~v3 & new_n2338_;
  assign new_n2340_ = v2 & new_n2339_;
  assign new_n2341_ = ~v1 & new_n2340_;
  assign new_n2342_ = ~v0 & new_n2341_;
  assign new_n2343_ = ~new_n2336_ & ~new_n2342_;
  assign new_n2344_ = v9 & ~new_n2343_;
  assign new_n2345_ = ~new_n160_ & ~new_n2344_;
  assign new_n2346_ = ~v24 & ~new_n2345_;
  assign new_n2347_ = ~v6 & new_n2137_;
  assign new_n2348_ = v5 & new_n2347_;
  assign new_n2349_ = ~v3 & new_n2348_;
  assign new_n2350_ = v2 & new_n2349_;
  assign new_n2351_ = ~v1 & new_n2350_;
  assign new_n2352_ = ~v0 & new_n2351_;
  assign new_n2353_ = ~new_n2346_ & ~new_n2352_;
  assign new_n2354_ = ~v8 & ~new_n2353_;
  assign new_n2355_ = v8 & new_n769_;
  assign new_n2356_ = v7 & new_n2355_;
  assign new_n2357_ = v6 & new_n2356_;
  assign new_n2358_ = ~v5 & new_n2357_;
  assign new_n2359_ = v3 & new_n2358_;
  assign new_n2360_ = ~v2 & new_n2359_;
  assign new_n2361_ = v1 & new_n2360_;
  assign new_n2362_ = v0 & new_n2361_;
  assign new_n2363_ = ~new_n2354_ & ~new_n2362_;
  assign new_n2364_ = v4 & ~new_n2363_;
  assign new_n2365_ = ~v5 & ~v24;
  assign new_n2366_ = v0 & new_n2365_;
  assign new_n2367_ = new_n278_ & new_n1425_;
  assign new_n2368_ = ~new_n2366_ & ~new_n2367_;
  assign new_n2369_ = ~v10 & ~new_n2368_;
  assign new_n2370_ = ~v8 & new_n258_;
  assign new_n2371_ = new_n1425_ & new_n2370_;
  assign new_n2372_ = ~new_n2369_ & ~new_n2371_;
  assign new_n2373_ = ~v9 & ~new_n2372_;
  assign new_n2374_ = v7 & new_n2373_;
  assign new_n2375_ = ~v5 & ~v7;
  assign new_n2376_ = v0 & new_n2375_;
  assign new_n2377_ = new_n310_ & new_n496_;
  assign new_n2378_ = new_n2376_ & new_n2377_;
  assign new_n2379_ = ~new_n2374_ & ~new_n2378_;
  assign new_n2380_ = v2 & ~new_n2379_;
  assign new_n2381_ = ~v24 & ~new_n835_;
  assign new_n2382_ = ~v10 & new_n2381_;
  assign new_n2383_ = v8 & new_n2382_;
  assign new_n2384_ = ~v5 & new_n2383_;
  assign new_n2385_ = ~v2 & new_n2384_;
  assign new_n2386_ = v0 & new_n2385_;
  assign new_n2387_ = ~new_n2380_ & ~new_n2386_;
  assign new_n2388_ = v3 & ~new_n2387_;
  assign new_n2389_ = new_n478_ & new_n1406_;
  assign new_n2390_ = new_n497_ & new_n1331_;
  assign new_n2391_ = new_n2389_ & new_n2390_;
  assign new_n2392_ = ~new_n2388_ & ~new_n2391_;
  assign new_n2393_ = ~v25 & ~new_n2392_;
  assign new_n2394_ = ~v23 & new_n2393_;
  assign new_n2395_ = v6 & new_n2394_;
  assign new_n2396_ = ~v4 & new_n2395_;
  assign new_n2397_ = ~v1 & new_n2396_;
  assign new_n2398_ = ~new_n2364_ & ~new_n2397_;
  assign \v26.25  = ~v22 & ~new_n2398_;
  assign new_n2400_ = new_n263_ & new_n1709_;
  assign new_n2401_ = new_n1039_ & new_n1721_;
  assign new_n2402_ = ~new_n2400_ & ~new_n2401_;
  assign new_n2403_ = ~v10 & ~new_n2402_;
  assign new_n2404_ = ~v7 & new_n2403_;
  assign new_n2405_ = v1 & new_n2404_;
  assign new_n2406_ = ~v3 & ~v6;
  assign new_n2407_ = ~v1 & new_n2406_;
  assign new_n2408_ = new_n834_ & new_n1563_;
  assign new_n2409_ = new_n2407_ & new_n2408_;
  assign new_n2410_ = ~new_n2405_ & ~new_n2409_;
  assign new_n2411_ = ~v25 & ~new_n2410_;
  assign new_n2412_ = ~v6 & v7;
  assign new_n2413_ = new_n589_ & new_n2412_;
  assign new_n2414_ = new_n187_ & new_n298_;
  assign new_n2415_ = new_n2413_ & new_n2414_;
  assign new_n2416_ = ~new_n2411_ & ~new_n2415_;
  assign new_n2417_ = v4 & ~new_n2416_;
  assign new_n2418_ = ~v4 & ~v6;
  assign new_n2419_ = new_n593_ & new_n2418_;
  assign new_n2420_ = new_n454_ & new_n834_;
  assign new_n2421_ = new_n2419_ & new_n2420_;
  assign new_n2422_ = ~new_n2417_ & ~new_n2421_;
  assign new_n2423_ = v5 & ~new_n2422_;
  assign new_n2424_ = v6 & new_n76_;
  assign new_n2425_ = ~new_n692_ & ~new_n2424_;
  assign new_n2426_ = ~v24 & ~new_n2425_;
  assign new_n2427_ = ~v9 & new_n2426_;
  assign new_n2428_ = ~v5 & new_n2427_;
  assign new_n2429_ = ~v4 & new_n2428_;
  assign new_n2430_ = ~v3 & new_n2429_;
  assign new_n2431_ = ~v1 & new_n2430_;
  assign new_n2432_ = ~new_n2423_ & ~new_n2431_;
  assign new_n2433_ = ~v2 & ~new_n2432_;
  assign new_n2434_ = v6 & ~v25;
  assign new_n2435_ = v5 & new_n2434_;
  assign new_n2436_ = new_n117_ & new_n856_;
  assign new_n2437_ = ~new_n2435_ & ~new_n2436_;
  assign new_n2438_ = ~v9 & ~new_n2437_;
  assign new_n2439_ = v9 & new_n856_;
  assign new_n2440_ = new_n117_ & new_n2439_;
  assign new_n2441_ = ~new_n2438_ & ~new_n2440_;
  assign new_n2442_ = v24 & ~new_n2441_;
  assign new_n2443_ = v7 & new_n2442_;
  assign new_n2444_ = ~v4 & new_n2443_;
  assign new_n2445_ = v3 & new_n2444_;
  assign new_n2446_ = v2 & new_n2445_;
  assign new_n2447_ = ~v1 & new_n2446_;
  assign new_n2448_ = ~new_n2433_ & ~new_n2447_;
  assign new_n2449_ = ~v0 & ~new_n2448_;
  assign new_n2450_ = v0 & new_n334_;
  assign new_n2451_ = v3 & new_n479_;
  assign new_n2452_ = new_n2450_ & new_n2451_;
  assign new_n2453_ = v6 & new_n834_;
  assign new_n2454_ = new_n1055_ & new_n2453_;
  assign new_n2455_ = new_n2452_ & new_n2454_;
  assign new_n2456_ = ~new_n2449_ & ~new_n2455_;
  assign new_n2457_ = ~v23 & ~new_n2456_;
  assign new_n2458_ = v24 & new_n1064_;
  assign new_n2459_ = v23 & new_n2458_;
  assign new_n2460_ = ~v10 & new_n2459_;
  assign new_n2461_ = ~v9 & new_n2460_;
  assign new_n2462_ = v7 & new_n2461_;
  assign new_n2463_ = v6 & new_n2462_;
  assign new_n2464_ = ~v5 & new_n2463_;
  assign new_n2465_ = ~v4 & new_n2464_;
  assign new_n2466_ = v0 & new_n2465_;
  assign new_n2467_ = ~new_n2457_ & ~new_n2466_;
  assign new_n2468_ = ~v8 & ~new_n2467_;
  assign new_n2469_ = v25 & ~new_n835_;
  assign new_n2470_ = v6 & new_n2469_;
  assign new_n2471_ = ~v5 & new_n2470_;
  assign new_n2472_ = v2 & new_n2471_;
  assign new_n2473_ = v1 & new_n2472_;
  assign new_n2474_ = v0 & new_n2473_;
  assign new_n2475_ = ~v2 & v5;
  assign new_n2476_ = new_n95_ & new_n2475_;
  assign new_n2477_ = new_n148_ & new_n632_;
  assign new_n2478_ = new_n2476_ & new_n2477_;
  assign new_n2479_ = ~new_n2474_ & ~new_n2478_;
  assign new_n2480_ = v3 & ~new_n2479_;
  assign new_n2481_ = v7 & new_n616_;
  assign new_n2482_ = new_n585_ & new_n2481_;
  assign new_n2483_ = new_n1787_ & new_n2482_;
  assign new_n2484_ = ~new_n2480_ & ~new_n2483_;
  assign new_n2485_ = ~v10 & ~new_n2484_;
  assign new_n2486_ = ~v4 & new_n2485_;
  assign new_n2487_ = ~v5 & new_n148_;
  assign new_n2488_ = new_n1029_ & new_n2487_;
  assign new_n2489_ = new_n727_ & new_n2488_;
  assign new_n2490_ = ~new_n2486_ & ~new_n2489_;
  assign new_n2491_ = ~v24 & ~new_n2490_;
  assign new_n2492_ = ~v23 & new_n2491_;
  assign new_n2493_ = v8 & new_n2492_;
  assign new_n2494_ = ~new_n2468_ & ~new_n2493_;
  assign \v26.26  = ~v22 & ~new_n2494_;
  assign new_n2496_ = ~v0 & new_n1308_;
  assign new_n2497_ = new_n696_ & new_n1680_;
  assign new_n2498_ = ~new_n2496_ & ~new_n2497_;
  assign new_n2499_ = ~new_n189_ & ~new_n2498_;
  assign new_n2500_ = v3 & new_n2499_;
  assign new_n2501_ = new_n441_ & new_n1431_;
  assign new_n2502_ = new_n187_ & new_n1163_;
  assign new_n2503_ = new_n2501_ & new_n2502_;
  assign new_n2504_ = ~new_n2500_ & ~new_n2503_;
  assign new_n2505_ = ~v5 & ~new_n2504_;
  assign new_n2506_ = ~v4 & new_n2505_;
  assign new_n2507_ = v10 & new_n188_;
  assign new_n2508_ = v9 & new_n2507_;
  assign new_n2509_ = ~v6 & new_n2508_;
  assign new_n2510_ = v5 & new_n2509_;
  assign new_n2511_ = v4 & new_n2510_;
  assign new_n2512_ = ~v3 & new_n2511_;
  assign new_n2513_ = ~v0 & new_n2512_;
  assign new_n2514_ = ~new_n2506_ & ~new_n2513_;
  assign new_n2515_ = ~v1 & ~new_n2514_;
  assign new_n2516_ = v23 & ~new_n189_;
  assign new_n2517_ = ~v10 & new_n2516_;
  assign new_n2518_ = ~v9 & new_n2517_;
  assign new_n2519_ = v6 & new_n2518_;
  assign new_n2520_ = ~v5 & new_n2519_;
  assign new_n2521_ = ~v4 & new_n2520_;
  assign new_n2522_ = v1 & new_n2521_;
  assign new_n2523_ = v0 & new_n2522_;
  assign new_n2524_ = ~new_n2515_ & ~new_n2523_;
  assign new_n2525_ = v2 & ~new_n2524_;
  assign new_n2526_ = ~v3 & new_n2521_;
  assign new_n2527_ = ~v2 & new_n2526_;
  assign new_n2528_ = v0 & new_n2527_;
  assign new_n2529_ = ~new_n2525_ & ~new_n2528_;
  assign new_n2530_ = ~v8 & ~new_n2529_;
  assign new_n2531_ = ~v23 & new_n194_;
  assign new_n2532_ = ~v10 & new_n2531_;
  assign new_n2533_ = v8 & new_n2532_;
  assign new_n2534_ = ~v6 & new_n2533_;
  assign new_n2535_ = v5 & new_n2534_;
  assign new_n2536_ = ~v4 & new_n2535_;
  assign new_n2537_ = ~v3 & new_n2536_;
  assign new_n2538_ = ~v2 & new_n2537_;
  assign new_n2539_ = ~v1 & new_n2538_;
  assign new_n2540_ = ~v0 & new_n2539_;
  assign new_n2541_ = ~new_n2530_ & ~new_n2540_;
  assign new_n2542_ = v7 & ~new_n2541_;
  assign new_n2543_ = new_n422_ & new_n1347_;
  assign new_n2544_ = ~new_n473_ & ~new_n2543_;
  assign new_n2545_ = v24 & ~new_n2544_;
  assign new_n2546_ = v2 & new_n2545_;
  assign new_n2547_ = ~v1 & new_n2546_;
  assign new_n2548_ = v9 & new_n496_;
  assign new_n2549_ = new_n922_ & new_n2548_;
  assign new_n2550_ = ~new_n2547_ & ~new_n2549_;
  assign new_n2551_ = ~v23 & ~new_n2550_;
  assign new_n2552_ = new_n398_ & new_n561_;
  assign new_n2553_ = new_n925_ & new_n2552_;
  assign new_n2554_ = ~new_n2551_ & ~new_n2553_;
  assign new_n2555_ = ~v25 & ~new_n2554_;
  assign new_n2556_ = ~v8 & new_n2555_;
  assign new_n2557_ = ~v7 & new_n2556_;
  assign new_n2558_ = v5 & new_n2557_;
  assign new_n2559_ = v4 & new_n2558_;
  assign new_n2560_ = ~v3 & new_n2559_;
  assign new_n2561_ = ~v0 & new_n2560_;
  assign new_n2562_ = ~new_n2542_ & ~new_n2561_;
  assign \v26.27  = ~v22 & ~new_n2562_;
  assign new_n2564_ = ~v24 & new_n1311_;
  assign new_n2565_ = new_n537_ & new_n1721_;
  assign new_n2566_ = new_n1164_ & new_n2565_;
  assign new_n2567_ = ~new_n2564_ & ~new_n2566_;
  assign new_n2568_ = ~v9 & ~new_n2567_;
  assign new_n2569_ = ~v23 & ~new_n189_;
  assign new_n2570_ = v10 & new_n2569_;
  assign new_n2571_ = v9 & new_n2570_;
  assign new_n2572_ = ~v6 & new_n2571_;
  assign new_n2573_ = v3 & new_n2572_;
  assign new_n2574_ = v2 & new_n2573_;
  assign new_n2575_ = ~v0 & new_n2574_;
  assign new_n2576_ = ~new_n2568_ & ~new_n2575_;
  assign new_n2577_ = ~v4 & ~new_n2576_;
  assign new_n2578_ = v3 & new_n1026_;
  assign new_n2579_ = new_n1009_ & new_n2578_;
  assign new_n2580_ = new_n118_ & new_n2531_;
  assign new_n2581_ = new_n2579_ & new_n2580_;
  assign new_n2582_ = ~new_n2577_ & ~new_n2581_;
  assign new_n2583_ = ~v5 & ~new_n2582_;
  assign new_n2584_ = new_n420_ & new_n537_;
  assign new_n2585_ = ~v23 & new_n188_;
  assign new_n2586_ = new_n473_ & new_n2585_;
  assign new_n2587_ = new_n2584_ & new_n2586_;
  assign new_n2588_ = ~new_n2583_ & ~new_n2587_;
  assign new_n2589_ = v7 & ~new_n2588_;
  assign new_n2590_ = v4 & new_n258_;
  assign new_n2591_ = new_n136_ & new_n2590_;
  assign new_n2592_ = ~v2 & v3;
  assign new_n2593_ = ~v4 & new_n496_;
  assign new_n2594_ = new_n2592_ & new_n2593_;
  assign new_n2595_ = ~new_n2591_ & ~new_n2594_;
  assign new_n2596_ = ~v25 & ~new_n2595_;
  assign new_n2597_ = ~v23 & new_n2596_;
  assign new_n2598_ = v9 & new_n2597_;
  assign new_n2599_ = ~v7 & new_n2598_;
  assign new_n2600_ = ~v6 & new_n2599_;
  assign new_n2601_ = v5 & new_n2600_;
  assign new_n2602_ = ~v0 & new_n2601_;
  assign new_n2603_ = ~new_n2589_ & ~new_n2602_;
  assign new_n2604_ = ~v8 & ~new_n2603_;
  assign new_n2605_ = new_n136_ & new_n473_;
  assign new_n2606_ = v6 & new_n118_;
  assign new_n2607_ = new_n2592_ & new_n2606_;
  assign new_n2608_ = ~new_n2605_ & ~new_n2607_;
  assign new_n2609_ = ~v25 & ~new_n2608_;
  assign new_n2610_ = ~v24 & new_n2609_;
  assign new_n2611_ = ~v23 & new_n2610_;
  assign new_n2612_ = v8 & new_n2611_;
  assign new_n2613_ = ~v7 & new_n2612_;
  assign new_n2614_ = ~v5 & new_n2613_;
  assign new_n2615_ = v4 & new_n2614_;
  assign new_n2616_ = ~v0 & new_n2615_;
  assign new_n2617_ = ~new_n2604_ & ~new_n2616_;
  assign new_n2618_ = ~v1 & ~new_n2617_;
  assign new_n2619_ = ~v9 & new_n2043_;
  assign new_n2620_ = v7 & new_n2619_;
  assign new_n2621_ = ~v5 & new_n2620_;
  assign new_n2622_ = ~v4 & new_n2621_;
  assign new_n2623_ = v0 & new_n2622_;
  assign new_n2624_ = new_n725_ & new_n1009_;
  assign new_n2625_ = v9 & ~v23;
  assign new_n2626_ = new_n73_ & new_n2625_;
  assign new_n2627_ = new_n2624_ & new_n2626_;
  assign new_n2628_ = ~new_n2623_ & ~new_n2627_;
  assign new_n2629_ = v25 & ~new_n2628_;
  assign new_n2630_ = ~v24 & new_n2629_;
  assign new_n2631_ = ~v10 & new_n2630_;
  assign new_n2632_ = ~v8 & new_n2631_;
  assign new_n2633_ = v6 & new_n2632_;
  assign new_n2634_ = v1 & new_n2633_;
  assign new_n2635_ = ~new_n2618_ & ~new_n2634_;
  assign \v26.28  = ~v22 & ~new_n2635_;
  assign new_n2637_ = v9 & ~new_n189_;
  assign new_n2638_ = ~v2 & new_n2637_;
  assign new_n2639_ = v1 & new_n2638_;
  assign new_n2640_ = v2 & ~v9;
  assign new_n2641_ = ~v1 & new_n2640_;
  assign new_n2642_ = new_n1804_ & new_n2641_;
  assign new_n2643_ = ~new_n2639_ & ~new_n2642_;
  assign new_n2644_ = ~v10 & ~new_n2643_;
  assign new_n2645_ = v6 & new_n2644_;
  assign new_n2646_ = new_n188_ & new_n398_;
  assign new_n2647_ = new_n925_ & new_n2646_;
  assign new_n2648_ = ~new_n2645_ & ~new_n2647_;
  assign new_n2649_ = ~v7 & ~new_n2648_;
  assign new_n2650_ = new_n418_ & new_n2412_;
  assign new_n2651_ = new_n2646_ & new_n2650_;
  assign new_n2652_ = ~new_n2649_ & ~new_n2651_;
  assign new_n2653_ = v5 & ~new_n2652_;
  assign new_n2654_ = v4 & new_n2653_;
  assign new_n2655_ = ~v6 & new_n77_;
  assign new_n2656_ = ~new_n2424_ & ~new_n2655_;
  assign new_n2657_ = ~v9 & ~new_n2656_;
  assign new_n2658_ = ~v2 & new_n2657_;
  assign new_n2659_ = v7 & new_n398_;
  assign new_n2660_ = new_n358_ & new_n2659_;
  assign new_n2661_ = ~new_n2658_ & ~new_n2660_;
  assign new_n2662_ = v25 & ~new_n2661_;
  assign new_n2663_ = ~v24 & new_n2662_;
  assign new_n2664_ = ~v5 & new_n2663_;
  assign new_n2665_ = ~v4 & new_n2664_;
  assign new_n2666_ = ~v1 & new_n2665_;
  assign new_n2667_ = ~new_n2654_ & ~new_n2666_;
  assign new_n2668_ = ~v3 & ~new_n2667_;
  assign new_n2669_ = v7 & new_n258_;
  assign new_n2670_ = ~v5 & new_n2669_;
  assign new_n2671_ = v2 & new_n2670_;
  assign new_n2672_ = ~v2 & new_n73_;
  assign new_n2673_ = new_n2548_ & new_n2672_;
  assign new_n2674_ = ~new_n2671_ & ~new_n2673_;
  assign new_n2675_ = ~v4 & ~new_n2674_;
  assign new_n2676_ = ~v2 & new_n450_;
  assign new_n2677_ = new_n496_ & new_n834_;
  assign new_n2678_ = new_n2676_ & new_n2677_;
  assign new_n2679_ = ~new_n2675_ & ~new_n2678_;
  assign new_n2680_ = ~v25 & ~new_n2679_;
  assign new_n2681_ = v10 & new_n200_;
  assign new_n2682_ = v7 & new_n2681_;
  assign new_n2683_ = ~v5 & new_n2682_;
  assign new_n2684_ = ~v4 & new_n2683_;
  assign new_n2685_ = v2 & new_n2684_;
  assign new_n2686_ = ~new_n2680_ & ~new_n2685_;
  assign new_n2687_ = ~v6 & ~new_n2686_;
  assign new_n2688_ = v3 & new_n2687_;
  assign new_n2689_ = ~v1 & new_n2688_;
  assign new_n2690_ = ~new_n2668_ & ~new_n2689_;
  assign new_n2691_ = ~v23 & ~new_n2690_;
  assign new_n2692_ = v4 & new_n2348_;
  assign new_n2693_ = ~v3 & new_n2692_;
  assign new_n2694_ = v2 & new_n2693_;
  assign new_n2695_ = ~v1 & new_n2694_;
  assign new_n2696_ = ~new_n2691_ & ~new_n2695_;
  assign new_n2697_ = ~v8 & ~new_n2696_;
  assign new_n2698_ = ~v1 & new_n2615_;
  assign new_n2699_ = ~new_n2697_ & ~new_n2698_;
  assign new_n2700_ = ~v0 & ~new_n2699_;
  assign new_n2701_ = ~v8 & new_n2461_;
  assign new_n2702_ = v7 & new_n2701_;
  assign new_n2703_ = v6 & new_n2702_;
  assign new_n2704_ = ~v5 & new_n2703_;
  assign new_n2705_ = ~v4 & new_n2704_;
  assign new_n2706_ = v0 & new_n2705_;
  assign new_n2707_ = ~new_n2700_ & ~new_n2706_;
  assign \v26.29  = ~v22 & ~new_n2707_;
  assign new_n2709_ = ~v4 & ~new_n1727_;
  assign new_n2710_ = ~v2 & new_n950_;
  assign new_n2711_ = v1 & new_n2710_;
  assign new_n2712_ = v0 & new_n2711_;
  assign new_n2713_ = ~new_n2709_ & ~new_n2712_;
  assign new_n2714_ = new_n712_ & new_n1382_;
  assign new_n2715_ = ~v8 & new_n1563_;
  assign new_n2716_ = new_n949_ & new_n2715_;
  assign new_n2717_ = new_n2714_ & new_n2716_;
  assign new_n2718_ = new_n2713_ & ~new_n2717_;
  assign new_n2719_ = v7 & ~new_n2718_;
  assign new_n2720_ = new_n95_ & new_n290_;
  assign new_n2721_ = ~v8 & new_n496_;
  assign new_n2722_ = new_n1046_ & new_n2721_;
  assign new_n2723_ = new_n2720_ & new_n2722_;
  assign new_n2724_ = ~new_n2719_ & ~new_n2723_;
  assign new_n2725_ = ~v23 & ~new_n2724_;
  assign new_n2726_ = v7 & new_n791_;
  assign new_n2727_ = v6 & new_n2726_;
  assign new_n2728_ = v4 & new_n2727_;
  assign new_n2729_ = v3 & new_n2728_;
  assign new_n2730_ = ~v2 & new_n2729_;
  assign new_n2731_ = v1 & new_n2730_;
  assign new_n2732_ = v0 & new_n2731_;
  assign new_n2733_ = ~new_n2725_ & ~new_n2732_;
  assign new_n2734_ = ~v5 & ~new_n2733_;
  assign new_n2735_ = v24 & ~new_n188_;
  assign new_n2736_ = ~v23 & ~new_n2735_;
  assign new_n2737_ = ~v10 & new_n2736_;
  assign new_n2738_ = v8 & new_n2737_;
  assign new_n2739_ = v7 & new_n2738_;
  assign new_n2740_ = ~v6 & new_n2739_;
  assign new_n2741_ = v5 & new_n2740_;
  assign new_n2742_ = ~v4 & new_n2741_;
  assign new_n2743_ = ~v3 & new_n2742_;
  assign new_n2744_ = ~v2 & new_n2743_;
  assign new_n2745_ = ~v1 & new_n2744_;
  assign new_n2746_ = ~v0 & new_n2745_;
  assign new_n2747_ = ~new_n2734_ & ~new_n2746_;
  assign new_n2748_ = v23 & ~new_n738_;
  assign new_n2749_ = v1 & new_n1147_;
  assign new_n2750_ = v5 & v10;
  assign new_n2751_ = new_n589_ & new_n2750_;
  assign new_n2752_ = ~new_n2749_ & ~new_n2751_;
  assign new_n2753_ = ~new_n2748_ & ~new_n2752_;
  assign new_n2754_ = v5 & new_n562_;
  assign new_n2755_ = ~v3 & new_n2754_;
  assign new_n2756_ = ~v1 & new_n2755_;
  assign new_n2757_ = ~new_n2753_ & ~new_n2756_;
  assign new_n2758_ = ~v7 & ~new_n2748_;
  assign new_n2759_ = v5 & new_n2758_;
  assign new_n2760_ = v3 & new_n2759_;
  assign new_n2761_ = v1 & new_n2760_;
  assign new_n2762_ = new_n2757_ & ~new_n2761_;
  assign new_n2763_ = ~v6 & ~new_n2762_;
  assign new_n2764_ = ~new_n81_ & ~new_n2748_;
  assign new_n2765_ = v1 & new_n2764_;
  assign new_n2766_ = v10 & new_n1287_;
  assign new_n2767_ = ~v1 & new_n73_;
  assign new_n2768_ = new_n2766_ & new_n2767_;
  assign new_n2769_ = ~new_n2765_ & ~new_n2768_;
  assign new_n2770_ = v6 & ~new_n2769_;
  assign new_n2771_ = v3 & new_n2770_;
  assign new_n2772_ = ~new_n2763_ & ~new_n2771_;
  assign new_n2773_ = v9 & ~new_n2772_;
  assign new_n2774_ = v3 & new_n552_;
  assign new_n2775_ = ~v3 & new_n930_;
  assign new_n2776_ = ~new_n2774_ & ~new_n2775_;
  assign new_n2777_ = ~v24 & ~new_n2776_;
  assign new_n2778_ = v6 & new_n225_;
  assign new_n2779_ = ~v3 & new_n2778_;
  assign new_n2780_ = ~new_n2777_ & ~new_n2779_;
  assign new_n2781_ = ~v23 & ~new_n2780_;
  assign new_n2782_ = ~v9 & new_n2781_;
  assign new_n2783_ = ~v7 & new_n2782_;
  assign new_n2784_ = v5 & new_n2783_;
  assign new_n2785_ = ~v1 & new_n2784_;
  assign new_n2786_ = ~new_n2773_ & ~new_n2785_;
  assign new_n2787_ = v2 & ~new_n2786_;
  assign new_n2788_ = ~v3 & new_n73_;
  assign new_n2789_ = ~new_n572_ & ~new_n2788_;
  assign new_n2790_ = ~v10 & ~new_n2789_;
  assign new_n2791_ = v9 & new_n2790_;
  assign new_n2792_ = v1 & new_n2791_;
  assign new_n2793_ = ~v1 & new_n1147_;
  assign new_n2794_ = v7 & new_n298_;
  assign new_n2795_ = new_n2793_ & new_n2794_;
  assign new_n2796_ = ~new_n2792_ & ~new_n2795_;
  assign new_n2797_ = ~new_n2735_ & ~new_n2796_;
  assign new_n2798_ = new_n73_ & new_n1943_;
  assign new_n2799_ = new_n194_ & new_n298_;
  assign new_n2800_ = new_n2798_ & new_n2799_;
  assign new_n2801_ = ~new_n2797_ & ~new_n2800_;
  assign new_n2802_ = v6 & ~new_n2801_;
  assign new_n2803_ = ~v3 & new_n2750_;
  assign new_n2804_ = v3 & new_n751_;
  assign new_n2805_ = ~new_n2803_ & ~new_n2804_;
  assign new_n2806_ = v7 & ~new_n2805_;
  assign new_n2807_ = ~v1 & new_n2806_;
  assign new_n2808_ = new_n80_ & new_n1943_;
  assign new_n2809_ = ~new_n2807_ & ~new_n2808_;
  assign new_n2810_ = ~v24 & ~new_n2809_;
  assign new_n2811_ = ~v9 & new_n2810_;
  assign new_n2812_ = ~v6 & new_n2811_;
  assign new_n2813_ = ~new_n2802_ & ~new_n2812_;
  assign new_n2814_ = ~v23 & ~new_n2813_;
  assign new_n2815_ = ~v2 & new_n2814_;
  assign new_n2816_ = ~new_n2787_ & ~new_n2815_;
  assign new_n2817_ = v4 & ~new_n2816_;
  assign new_n2818_ = v5 & ~new_n835_;
  assign new_n2819_ = v3 & new_n2818_;
  assign new_n2820_ = new_n1094_ & new_n1406_;
  assign new_n2821_ = ~new_n2819_ & ~new_n2820_;
  assign new_n2822_ = ~v10 & ~new_n2821_;
  assign new_n2823_ = ~v6 & new_n2822_;
  assign new_n2824_ = ~v3 & new_n585_;
  assign new_n2825_ = new_n2794_ & new_n2824_;
  assign new_n2826_ = ~new_n2823_ & ~new_n2825_;
  assign new_n2827_ = ~v2 & ~new_n2826_;
  assign new_n2828_ = v5 & new_n422_;
  assign new_n2829_ = v3 & new_n2828_;
  assign new_n2830_ = new_n473_ & new_n1406_;
  assign new_n2831_ = ~new_n2829_ & ~new_n2830_;
  assign new_n2832_ = v7 & ~new_n2831_;
  assign new_n2833_ = v2 & new_n2832_;
  assign new_n2834_ = ~new_n2827_ & ~new_n2833_;
  assign new_n2835_ = ~v24 & ~new_n2834_;
  assign new_n2836_ = v5 & new_n533_;
  assign new_n2837_ = v3 & new_n2836_;
  assign new_n2838_ = v2 & new_n2837_;
  assign new_n2839_ = new_n1407_ & new_n2655_;
  assign new_n2840_ = ~new_n2838_ & ~new_n2839_;
  assign new_n2841_ = v24 & ~new_n2840_;
  assign new_n2842_ = ~v9 & new_n2841_;
  assign new_n2843_ = ~new_n2835_ & ~new_n2842_;
  assign new_n2844_ = ~v1 & ~new_n2843_;
  assign new_n2845_ = new_n853_ & new_n1147_;
  assign new_n2846_ = new_n1046_ & new_n2548_;
  assign new_n2847_ = new_n2845_ & new_n2846_;
  assign new_n2848_ = ~new_n2844_ & ~new_n2847_;
  assign new_n2849_ = v3 & new_n117_;
  assign new_n2850_ = new_n114_ & new_n2849_;
  assign new_n2851_ = v7 & v9;
  assign new_n2852_ = new_n454_ & new_n2851_;
  assign new_n2853_ = new_n2850_ & new_n2852_;
  assign new_n2854_ = new_n2848_ & ~new_n2853_;
  assign new_n2855_ = ~v23 & ~new_n2854_;
  assign new_n2856_ = ~v25 & ~new_n2840_;
  assign new_n2857_ = ~v24 & new_n2856_;
  assign new_n2858_ = v23 & new_n2857_;
  assign new_n2859_ = ~v9 & new_n2858_;
  assign new_n2860_ = ~v1 & new_n2859_;
  assign new_n2861_ = ~new_n2855_ & ~new_n2860_;
  assign new_n2862_ = ~v4 & ~new_n2861_;
  assign new_n2863_ = ~new_n2817_ & ~new_n2862_;
  assign new_n2864_ = ~v0 & ~new_n2863_;
  assign new_n2865_ = ~new_n714_ & ~new_n2748_;
  assign new_n2866_ = ~v3 & ~new_n2748_;
  assign new_n2867_ = v2 & new_n2866_;
  assign new_n2868_ = v1 & new_n2867_;
  assign new_n2869_ = ~new_n2865_ & ~new_n2868_;
  assign new_n2870_ = ~v4 & ~new_n2869_;
  assign new_n2871_ = ~v1 & new_n712_;
  assign new_n2872_ = v4 & new_n1287_;
  assign new_n2873_ = new_n2871_ & new_n2872_;
  assign new_n2874_ = ~new_n2870_ & ~new_n2873_;
  assign new_n2875_ = ~v4 & new_n2459_;
  assign new_n2876_ = new_n2874_ & ~new_n2875_;
  assign new_n2877_ = ~v10 & ~new_n2876_;
  assign new_n2878_ = ~v9 & new_n2877_;
  assign new_n2879_ = v7 & new_n2878_;
  assign new_n2880_ = v6 & new_n2879_;
  assign new_n2881_ = ~v5 & new_n2880_;
  assign new_n2882_ = v0 & new_n2881_;
  assign new_n2883_ = ~new_n2864_ & ~new_n2882_;
  assign new_n2884_ = ~v8 & ~new_n2883_;
  assign new_n2885_ = v3 & ~new_n1091_;
  assign new_n2886_ = new_n1431_ & new_n2851_;
  assign new_n2887_ = ~new_n2885_ & ~new_n2886_;
  assign new_n2888_ = ~v2 & ~new_n2887_;
  assign new_n2889_ = v3 & ~new_n835_;
  assign new_n2890_ = v2 & new_n2889_;
  assign new_n2891_ = v0 & new_n2890_;
  assign new_n2892_ = ~new_n2888_ & ~new_n2891_;
  assign new_n2893_ = ~v10 & ~new_n2892_;
  assign new_n2894_ = ~v0 & new_n713_;
  assign new_n2895_ = ~v7 & new_n398_;
  assign new_n2896_ = new_n2894_ & new_n2895_;
  assign new_n2897_ = ~new_n2893_ & ~new_n2896_;
  assign new_n2898_ = v6 & ~new_n2897_;
  assign new_n2899_ = ~v6 & new_n834_;
  assign new_n2900_ = v3 & new_n2899_;
  assign new_n2901_ = v2 & new_n2900_;
  assign new_n2902_ = ~v0 & new_n2901_;
  assign new_n2903_ = ~new_n2898_ & ~new_n2902_;
  assign new_n2904_ = ~v1 & ~new_n2903_;
  assign new_n2905_ = v2 & ~new_n835_;
  assign new_n2906_ = new_n713_ & new_n830_;
  assign new_n2907_ = ~new_n2905_ & ~new_n2906_;
  assign new_n2908_ = ~v10 & ~new_n2907_;
  assign new_n2909_ = v6 & new_n2908_;
  assign new_n2910_ = v1 & new_n2909_;
  assign new_n2911_ = v0 & new_n2910_;
  assign new_n2912_ = ~new_n2904_ & ~new_n2911_;
  assign new_n2913_ = ~v5 & ~new_n2912_;
  assign new_n2914_ = ~new_n1046_ & ~new_n2412_;
  assign new_n2915_ = v3 & ~new_n2914_;
  assign new_n2916_ = ~new_n1053_ & ~new_n2915_;
  assign new_n2917_ = v10 & ~new_n2916_;
  assign new_n2918_ = ~v2 & new_n2917_;
  assign new_n2919_ = ~v1 & new_n2918_;
  assign new_n2920_ = ~v0 & new_n2919_;
  assign new_n2921_ = v7 & ~v10;
  assign new_n2922_ = new_n1709_ & new_n2921_;
  assign new_n2923_ = new_n2450_ & new_n2922_;
  assign new_n2924_ = ~new_n2920_ & ~new_n2923_;
  assign new_n2925_ = v9 & ~new_n2924_;
  assign new_n2926_ = new_n95_ & new_n2592_;
  assign new_n2927_ = new_n118_ & new_n148_;
  assign new_n2928_ = new_n2926_ & new_n2927_;
  assign new_n2929_ = ~new_n2925_ & ~new_n2928_;
  assign new_n2930_ = v5 & ~new_n2929_;
  assign new_n2931_ = ~new_n2913_ & ~new_n2930_;
  assign new_n2932_ = ~v4 & ~new_n2931_;
  assign new_n2933_ = ~v5 & v9;
  assign new_n2934_ = v0 & new_n2933_;
  assign new_n2935_ = new_n298_ & new_n1425_;
  assign new_n2936_ = ~new_n2934_ & ~new_n2935_;
  assign new_n2937_ = v7 & ~new_n2936_;
  assign new_n2938_ = v6 & new_n2937_;
  assign new_n2939_ = ~v0 & new_n138_;
  assign new_n2940_ = ~v7 & new_n298_;
  assign new_n2941_ = new_n2939_ & new_n2940_;
  assign new_n2942_ = ~new_n2938_ & ~new_n2941_;
  assign new_n2943_ = v2 & ~new_n2942_;
  assign new_n2944_ = ~v2 & ~v5;
  assign new_n2945_ = ~v0 & new_n2944_;
  assign new_n2946_ = new_n118_ & new_n1046_;
  assign new_n2947_ = new_n2945_ & new_n2946_;
  assign new_n2948_ = ~new_n2943_ & ~new_n2947_;
  assign new_n2949_ = ~v1 & ~new_n2948_;
  assign new_n2950_ = new_n254_ & new_n2944_;
  assign new_n2951_ = new_n298_ & new_n533_;
  assign new_n2952_ = new_n2950_ & new_n2951_;
  assign new_n2953_ = ~new_n2949_ & ~new_n2952_;
  assign new_n2954_ = v4 & ~new_n2953_;
  assign new_n2955_ = v3 & new_n2954_;
  assign new_n2956_ = ~new_n2932_ & ~new_n2955_;
  assign new_n2957_ = ~v24 & ~new_n2956_;
  assign new_n2958_ = v5 & v9;
  assign new_n2959_ = ~new_n1442_ & ~new_n2958_;
  assign new_n2960_ = ~v10 & ~new_n2959_;
  assign new_n2961_ = ~v4 & new_n2960_;
  assign new_n2962_ = ~v3 & new_n2961_;
  assign new_n2963_ = v1 & new_n2962_;
  assign new_n2964_ = v0 & new_n2963_;
  assign new_n2965_ = new_n298_ & new_n419_;
  assign new_n2966_ = new_n594_ & new_n2965_;
  assign new_n2967_ = ~new_n2964_ & ~new_n2966_;
  assign new_n2968_ = v7 & ~new_n2967_;
  assign new_n2969_ = new_n300_ & new_n2375_;
  assign new_n2970_ = new_n1867_ & new_n2969_;
  assign new_n2971_ = ~new_n2968_ & ~new_n2970_;
  assign new_n2972_ = v2 & ~new_n2971_;
  assign new_n2973_ = new_n289_ & new_n713_;
  assign new_n2974_ = ~v7 & new_n300_;
  assign new_n2975_ = new_n479_ & new_n2974_;
  assign new_n2976_ = new_n2973_ & new_n2975_;
  assign new_n2977_ = ~new_n2972_ & ~new_n2976_;
  assign new_n2978_ = v24 & ~new_n2977_;
  assign new_n2979_ = v6 & new_n2978_;
  assign new_n2980_ = ~new_n2957_ & ~new_n2979_;
  assign new_n2981_ = v0 & new_n2889_;
  assign new_n2982_ = ~new_n2886_ & ~new_n2981_;
  assign new_n2983_ = ~v10 & ~new_n2982_;
  assign new_n2984_ = new_n1431_ & new_n2895_;
  assign new_n2985_ = ~new_n2983_ & ~new_n2984_;
  assign new_n2986_ = ~v2 & ~new_n2985_;
  assign new_n2987_ = ~v10 & ~new_n835_;
  assign new_n2988_ = v3 & new_n2987_;
  assign new_n2989_ = v2 & new_n2988_;
  assign new_n2990_ = v0 & new_n2989_;
  assign new_n2991_ = ~new_n2986_ & ~new_n2990_;
  assign new_n2992_ = ~v5 & ~new_n2991_;
  assign new_n2993_ = v5 & new_n2895_;
  assign new_n2994_ = ~v2 & new_n2993_;
  assign new_n2995_ = ~v0 & new_n2994_;
  assign new_n2996_ = ~new_n2992_ & ~new_n2995_;
  assign new_n2997_ = v24 & ~new_n2996_;
  assign new_n2998_ = v6 & new_n2997_;
  assign new_n2999_ = ~v4 & new_n2998_;
  assign new_n3000_ = ~v3 & new_n450_;
  assign new_n3001_ = new_n537_ & new_n3000_;
  assign new_n3002_ = v9 & new_n1563_;
  assign new_n3003_ = new_n148_ & new_n3002_;
  assign new_n3004_ = new_n3001_ & new_n3003_;
  assign new_n3005_ = ~new_n2999_ & ~new_n3004_;
  assign new_n3006_ = ~v25 & ~new_n3005_;
  assign new_n3007_ = ~v1 & new_n3006_;
  assign new_n3008_ = new_n2980_ & ~new_n3007_;
  assign new_n3009_ = ~v23 & ~new_n3008_;
  assign new_n3010_ = v8 & new_n3009_;
  assign new_n3011_ = ~new_n2884_ & ~new_n3010_;
  assign new_n3012_ = new_n2747_ & new_n3011_;
  assign \v26.30  = ~v22 & ~new_n3012_;
  assign new_n3014_ = v10 & v23;
  assign new_n3015_ = ~v8 & new_n3014_;
  assign new_n3016_ = ~v6 & new_n3015_;
  assign new_n3017_ = v5 & new_n3016_;
  assign new_n3018_ = v4 & new_n3017_;
  assign new_n3019_ = v2 & new_n3018_;
  assign new_n3020_ = ~v1 & new_n3019_;
  assign new_n3021_ = ~v0 & new_n3020_;
  assign new_n3022_ = new_n289_ & new_n319_;
  assign new_n3023_ = ~v10 & ~v23;
  assign new_n3024_ = v8 & new_n3023_;
  assign new_n3025_ = new_n585_ & new_n3024_;
  assign new_n3026_ = new_n3022_ & new_n3025_;
  assign new_n3027_ = ~new_n3021_ & ~new_n3026_;
  assign new_n3028_ = v5 & v7;
  assign new_n3029_ = ~new_n2375_ & ~new_n3028_;
  assign new_n3030_ = ~v23 & ~new_n3029_;
  assign new_n3031_ = ~v10 & new_n3030_;
  assign new_n3032_ = v8 & new_n3031_;
  assign new_n3033_ = v6 & new_n3032_;
  assign new_n3034_ = ~v4 & new_n3033_;
  assign new_n3035_ = v2 & new_n3034_;
  assign new_n3036_ = v1 & new_n3035_;
  assign new_n3037_ = v0 & new_n3036_;
  assign new_n3038_ = new_n3027_ & ~new_n3037_;
  assign new_n3039_ = v25 & ~new_n3038_;
  assign new_n3040_ = ~v2 & new_n419_;
  assign new_n3041_ = new_n254_ & new_n3040_;
  assign new_n3042_ = v6 & new_n1125_;
  assign new_n3043_ = ~v10 & new_n173_;
  assign new_n3044_ = new_n3042_ & new_n3043_;
  assign new_n3045_ = new_n3041_ & new_n3044_;
  assign new_n3046_ = ~new_n3039_ & ~new_n3045_;
  assign new_n3047_ = ~v3 & ~new_n3046_;
  assign new_n3048_ = v8 & new_n322_;
  assign new_n3049_ = ~v7 & new_n3048_;
  assign new_n3050_ = v6 & new_n3049_;
  assign new_n3051_ = v0 & new_n3050_;
  assign new_n3052_ = new_n856_ & new_n1331_;
  assign new_n3053_ = new_n532_ & new_n3052_;
  assign new_n3054_ = ~new_n3051_ & ~new_n3053_;
  assign new_n3055_ = ~v4 & ~new_n3054_;
  assign new_n3056_ = ~v1 & new_n3055_;
  assign new_n3057_ = ~v8 & new_n322_;
  assign new_n3058_ = new_n533_ & new_n3057_;
  assign new_n3059_ = new_n2080_ & new_n3058_;
  assign new_n3060_ = ~new_n3056_ & ~new_n3059_;
  assign new_n3061_ = ~v23 & ~new_n3060_;
  assign new_n3062_ = ~v5 & new_n3061_;
  assign new_n3063_ = v3 & new_n3062_;
  assign new_n3064_ = ~new_n3047_ & ~new_n3063_;
  assign new_n3065_ = v9 & ~new_n3064_;
  assign new_n3066_ = v6 & new_n3048_;
  assign new_n3067_ = v0 & new_n3066_;
  assign new_n3068_ = ~v8 & new_n856_;
  assign new_n3069_ = new_n532_ & new_n3068_;
  assign new_n3070_ = ~new_n3067_ & ~new_n3069_;
  assign new_n3071_ = ~v4 & ~new_n3070_;
  assign new_n3072_ = ~v0 & new_n346_;
  assign new_n3073_ = new_n433_ & new_n1437_;
  assign new_n3074_ = new_n3072_ & new_n3073_;
  assign new_n3075_ = ~new_n3071_ & ~new_n3074_;
  assign new_n3076_ = v3 & ~new_n3075_;
  assign new_n3077_ = ~v1 & new_n3076_;
  assign new_n3078_ = v8 & new_n430_;
  assign new_n3079_ = v6 & new_n3078_;
  assign new_n3080_ = ~v4 & new_n3079_;
  assign new_n3081_ = ~v3 & new_n3080_;
  assign new_n3082_ = v1 & new_n3081_;
  assign new_n3083_ = v0 & new_n3082_;
  assign new_n3084_ = ~new_n3077_ & ~new_n3083_;
  assign new_n3085_ = v7 & ~new_n3084_;
  assign new_n3086_ = ~v5 & new_n3085_;
  assign new_n3087_ = new_n420_ & new_n545_;
  assign new_n3088_ = new_n424_ & new_n3042_;
  assign new_n3089_ = new_n3087_ & new_n3088_;
  assign new_n3090_ = ~new_n3086_ & ~new_n3089_;
  assign new_n3091_ = ~v23 & ~new_n3090_;
  assign new_n3092_ = ~v9 & new_n3091_;
  assign new_n3093_ = ~new_n3065_ & ~new_n3092_;
  assign new_n3094_ = v24 & ~new_n3093_;
  assign new_n3095_ = ~v4 & v7;
  assign new_n3096_ = new_n327_ & new_n3095_;
  assign new_n3097_ = v4 & ~v7;
  assign new_n3098_ = new_n328_ & new_n3097_;
  assign new_n3099_ = ~new_n3096_ & ~new_n3098_;
  assign new_n3100_ = v10 & ~new_n3099_;
  assign new_n3101_ = v9 & new_n3100_;
  assign new_n3102_ = ~v3 & new_n3101_;
  assign new_n3103_ = v2 & new_n3102_;
  assign new_n3104_ = new_n854_ & new_n2592_;
  assign new_n3105_ = new_n368_ & new_n430_;
  assign new_n3106_ = new_n3104_ & new_n3105_;
  assign new_n3107_ = ~new_n3103_ & ~new_n3106_;
  assign new_n3108_ = ~v6 & ~new_n3107_;
  assign new_n3109_ = ~new_n3095_ & ~new_n3097_;
  assign new_n3110_ = v25 & ~new_n3109_;
  assign new_n3111_ = ~v10 & new_n3110_;
  assign new_n3112_ = ~v9 & new_n3111_;
  assign new_n3113_ = v8 & new_n3112_;
  assign new_n3114_ = v6 & new_n3113_;
  assign new_n3115_ = v3 & new_n3114_;
  assign new_n3116_ = ~v2 & new_n3115_;
  assign new_n3117_ = ~new_n3108_ & ~new_n3116_;
  assign new_n3118_ = ~v5 & ~new_n3117_;
  assign new_n3119_ = ~v19 & v25;
  assign new_n3120_ = ~v10 & new_n3119_;
  assign new_n3121_ = v8 & new_n3120_;
  assign new_n3122_ = v7 & new_n3121_;
  assign new_n3123_ = ~v6 & new_n3122_;
  assign new_n3124_ = v5 & new_n3123_;
  assign new_n3125_ = ~v4 & new_n3124_;
  assign new_n3126_ = ~v3 & new_n3125_;
  assign new_n3127_ = ~v2 & new_n3126_;
  assign new_n3128_ = ~new_n3118_ & ~new_n3127_;
  assign new_n3129_ = ~v23 & ~new_n3128_;
  assign new_n3130_ = ~v4 & new_n117_;
  assign new_n3131_ = new_n713_ & new_n3130_;
  assign new_n3132_ = new_n1183_ & new_n1824_;
  assign new_n3133_ = new_n3131_ & new_n3132_;
  assign new_n3134_ = ~new_n3129_ & ~new_n3133_;
  assign new_n3135_ = ~v1 & ~new_n3134_;
  assign new_n3136_ = v1 & new_n2592_;
  assign new_n3137_ = v4 & new_n546_;
  assign new_n3138_ = new_n3136_ & new_n3137_;
  assign new_n3139_ = v10 & new_n173_;
  assign new_n3140_ = new_n1824_ & new_n3139_;
  assign new_n3141_ = new_n3138_ & new_n3140_;
  assign new_n3142_ = ~new_n3135_ & ~new_n3141_;
  assign new_n3143_ = ~v24 & ~new_n3142_;
  assign new_n3144_ = ~v0 & new_n3143_;
  assign new_n3145_ = ~new_n3094_ & ~new_n3144_;
  assign \v26.31  = ~v22 & ~new_n3145_;
  assign new_n3147_ = ~v3 & new_n344_;
  assign new_n3148_ = v0 & new_n3147_;
  assign new_n3149_ = v4 & ~v8;
  assign new_n3150_ = v3 & new_n3149_;
  assign new_n3151_ = new_n537_ & new_n3150_;
  assign new_n3152_ = ~new_n3148_ & ~new_n3151_;
  assign new_n3153_ = ~v25 & ~new_n3152_;
  assign new_n3154_ = v4 & new_n327_;
  assign new_n3155_ = new_n1307_ & new_n3154_;
  assign new_n3156_ = ~new_n3153_ & ~new_n3155_;
  assign new_n3157_ = v24 & ~new_n3156_;
  assign new_n3158_ = v1 & new_n3157_;
  assign new_n3159_ = ~v4 & new_n976_;
  assign new_n3160_ = v3 & new_n3159_;
  assign new_n3161_ = ~v1 & new_n3160_;
  assign new_n3162_ = v0 & new_n3161_;
  assign new_n3163_ = ~new_n3158_ & ~new_n3162_;
  assign new_n3164_ = v6 & ~new_n3163_;
  assign new_n3165_ = v4 & new_n1510_;
  assign new_n3166_ = v3 & new_n3165_;
  assign new_n3167_ = v2 & new_n3166_;
  assign new_n3168_ = v1 & new_n3167_;
  assign new_n3169_ = ~v0 & new_n3168_;
  assign new_n3170_ = ~new_n3164_ & ~new_n3169_;
  assign new_n3171_ = ~v7 & ~new_n3170_;
  assign new_n3172_ = ~v6 & v24;
  assign new_n3173_ = v2 & new_n3172_;
  assign new_n3174_ = new_n187_ & new_n361_;
  assign new_n3175_ = ~new_n3173_ & ~new_n3174_;
  assign new_n3176_ = ~v8 & ~new_n3175_;
  assign new_n3177_ = v7 & new_n3176_;
  assign new_n3178_ = v4 & new_n3177_;
  assign new_n3179_ = v3 & new_n3178_;
  assign new_n3180_ = v1 & new_n3179_;
  assign new_n3181_ = ~v0 & new_n3180_;
  assign new_n3182_ = ~new_n3171_ & ~new_n3181_;
  assign new_n3183_ = ~v10 & ~new_n3182_;
  assign new_n3184_ = v6 & ~new_n533_;
  assign new_n3185_ = v24 & ~new_n3184_;
  assign new_n3186_ = v10 & new_n3185_;
  assign new_n3187_ = ~v8 & new_n3186_;
  assign new_n3188_ = v4 & new_n3187_;
  assign new_n3189_ = v3 & new_n3188_;
  assign new_n3190_ = v2 & new_n3189_;
  assign new_n3191_ = v1 & new_n3190_;
  assign new_n3192_ = ~v0 & new_n3191_;
  assign new_n3193_ = ~new_n3183_ & ~new_n3192_;
  assign new_n3194_ = ~v5 & ~new_n3193_;
  assign new_n3195_ = ~v8 & new_n1959_;
  assign new_n3196_ = ~v7 & new_n3195_;
  assign new_n3197_ = v5 & new_n3196_;
  assign new_n3198_ = v4 & new_n3197_;
  assign new_n3199_ = v3 & new_n3198_;
  assign new_n3200_ = v2 & new_n3199_;
  assign new_n3201_ = v1 & new_n3200_;
  assign new_n3202_ = ~v0 & new_n3201_;
  assign new_n3203_ = ~new_n3194_ & ~new_n3202_;
  assign new_n3204_ = v9 & ~new_n3203_;
  assign new_n3205_ = new_n235_ & new_n451_;
  assign new_n3206_ = v6 & new_n1331_;
  assign new_n3207_ = new_n2414_ & new_n3206_;
  assign new_n3208_ = new_n3205_ & new_n3207_;
  assign new_n3209_ = ~new_n3204_ & ~new_n3208_;
  assign new_n3210_ = ~v23 & ~new_n3209_;
  assign \v26.32  = ~v22 & new_n3210_;
  assign new_n3212_ = new_n1147_ & new_n2018_;
  assign new_n3213_ = ~v7 & ~v25;
  assign new_n3214_ = new_n145_ & new_n3213_;
  assign new_n3215_ = ~new_n3212_ & ~new_n3214_;
  assign new_n3216_ = ~v8 & ~new_n3215_;
  assign new_n3217_ = v6 & new_n3216_;
  assign new_n3218_ = v4 & new_n3217_;
  assign new_n3219_ = v1 & new_n3218_;
  assign new_n3220_ = new_n236_ & new_n589_;
  assign new_n3221_ = new_n328_ & new_n2412_;
  assign new_n3222_ = new_n3220_ & new_n3221_;
  assign new_n3223_ = ~new_n3219_ & ~new_n3222_;
  assign new_n3224_ = v9 & ~new_n3223_;
  assign new_n3225_ = v8 & new_n632_;
  assign new_n3226_ = new_n2412_ & new_n3225_;
  assign new_n3227_ = new_n3220_ & new_n3226_;
  assign new_n3228_ = ~new_n3224_ & ~new_n3227_;
  assign new_n3229_ = ~v10 & ~new_n3228_;
  assign new_n3230_ = v4 & new_n585_;
  assign new_n3231_ = new_n593_ & new_n3230_;
  assign new_n3232_ = ~v9 & new_n856_;
  assign new_n3233_ = new_n1331_ & new_n3232_;
  assign new_n3234_ = new_n3231_ & new_n3233_;
  assign new_n3235_ = ~new_n3229_ & ~new_n3234_;
  assign new_n3236_ = ~v24 & ~new_n3235_;
  assign new_n3237_ = ~v2 & new_n3236_;
  assign new_n3238_ = v1 & new_n712_;
  assign new_n3239_ = new_n2211_ & new_n3238_;
  assign new_n3240_ = new_n1162_ & new_n1814_;
  assign new_n3241_ = new_n3239_ & new_n3240_;
  assign new_n3242_ = ~new_n3237_ & ~new_n3241_;
  assign new_n3243_ = ~v23 & ~new_n3242_;
  assign new_n3244_ = ~v22 & new_n3243_;
  assign \v26.33  = ~v0 & new_n3244_;
  assign new_n3246_ = ~v3 & new_n882_;
  assign new_n3247_ = v3 & new_n1125_;
  assign new_n3248_ = ~new_n3246_ & ~new_n3247_;
  assign new_n3249_ = ~v24 & ~new_n3248_;
  assign new_n3250_ = ~v4 & new_n3249_;
  assign new_n3251_ = ~v2 & new_n3250_;
  assign new_n3252_ = ~v1 & new_n3251_;
  assign new_n3253_ = new_n278_ & new_n3097_;
  assign new_n3254_ = new_n3238_ & new_n3253_;
  assign new_n3255_ = ~new_n3252_ & ~new_n3254_;
  assign new_n3256_ = v9 & ~new_n3255_;
  assign new_n3257_ = new_n882_ & new_n1039_;
  assign new_n3258_ = new_n116_ & new_n3257_;
  assign new_n3259_ = ~new_n3256_ & ~new_n3258_;
  assign new_n3260_ = v5 & ~new_n3259_;
  assign new_n3261_ = ~v5 & new_n264_;
  assign new_n3262_ = v4 & new_n3261_;
  assign new_n3263_ = v3 & new_n3262_;
  assign new_n3264_ = v2 & new_n3263_;
  assign new_n3265_ = v1 & new_n3264_;
  assign new_n3266_ = ~new_n3260_ & ~new_n3265_;
  assign new_n3267_ = ~v25 & ~new_n3266_;
  assign new_n3268_ = v25 & ~new_n74_;
  assign new_n3269_ = v24 & new_n3268_;
  assign new_n3270_ = v9 & new_n3269_;
  assign new_n3271_ = ~v8 & new_n3270_;
  assign new_n3272_ = v4 & new_n3271_;
  assign new_n3273_ = v3 & new_n3272_;
  assign new_n3274_ = v2 & new_n3273_;
  assign new_n3275_ = v1 & new_n3274_;
  assign new_n3276_ = ~new_n3267_ & ~new_n3275_;
  assign new_n3277_ = ~v10 & ~new_n3276_;
  assign new_n3278_ = ~v5 & new_n2018_;
  assign new_n3279_ = v7 & ~new_n3278_;
  assign new_n3280_ = v24 & ~new_n3279_;
  assign new_n3281_ = v4 & new_n3280_;
  assign new_n3282_ = v3 & new_n3281_;
  assign new_n3283_ = v1 & new_n3282_;
  assign new_n3284_ = new_n187_ & new_n571_;
  assign new_n3285_ = new_n811_ & new_n3284_;
  assign new_n3286_ = ~new_n3283_ & ~new_n3285_;
  assign new_n3287_ = v10 & ~new_n3286_;
  assign new_n3288_ = v9 & new_n3287_;
  assign new_n3289_ = ~v8 & new_n3288_;
  assign new_n3290_ = v2 & new_n3289_;
  assign new_n3291_ = ~new_n3277_ & ~new_n3290_;
  assign new_n3292_ = ~v6 & ~new_n3291_;
  assign new_n3293_ = v9 & new_n430_;
  assign new_n3294_ = new_n571_ & new_n3293_;
  assign new_n3295_ = ~v9 & new_n433_;
  assign new_n3296_ = new_n73_ & new_n3295_;
  assign new_n3297_ = ~new_n3294_ & ~new_n3296_;
  assign new_n3298_ = v1 & ~new_n3297_;
  assign new_n3299_ = ~v1 & new_n571_;
  assign new_n3300_ = new_n3232_ & new_n3299_;
  assign new_n3301_ = ~new_n3298_ & ~new_n3300_;
  assign new_n3302_ = ~v24 & ~new_n3301_;
  assign new_n3303_ = ~v2 & new_n3302_;
  assign new_n3304_ = new_n571_ & new_n856_;
  assign new_n3305_ = ~new_n77_ & ~new_n3304_;
  assign new_n3306_ = v24 & ~new_n3305_;
  assign new_n3307_ = v9 & new_n3306_;
  assign new_n3308_ = v2 & new_n3307_;
  assign new_n3309_ = v1 & new_n3308_;
  assign new_n3310_ = ~new_n3303_ & ~new_n3309_;
  assign new_n3311_ = v3 & ~new_n3310_;
  assign new_n3312_ = new_n145_ & new_n853_;
  assign new_n3313_ = new_n454_ & new_n830_;
  assign new_n3314_ = new_n3312_ & new_n3313_;
  assign new_n3315_ = ~new_n3311_ & ~new_n3314_;
  assign new_n3316_ = ~v8 & ~new_n3315_;
  assign new_n3317_ = v6 & new_n3316_;
  assign new_n3318_ = v4 & new_n3317_;
  assign new_n3319_ = ~new_n3292_ & ~new_n3318_;
  assign new_n3320_ = ~v0 & ~new_n3319_;
  assign new_n3321_ = ~v10 & new_n2257_;
  assign new_n3322_ = v9 & new_n3321_;
  assign new_n3323_ = v8 & new_n3322_;
  assign new_n3324_ = ~v7 & new_n3323_;
  assign new_n3325_ = v6 & new_n3324_;
  assign new_n3326_ = ~v5 & new_n3325_;
  assign new_n3327_ = ~v4 & new_n3326_;
  assign new_n3328_ = v0 & new_n3327_;
  assign new_n3329_ = ~new_n3320_ & ~new_n3328_;
  assign new_n3330_ = ~v23 & ~new_n3329_;
  assign \v26.34  = ~v22 & new_n3330_;
  assign new_n3332_ = ~v2 & new_n138_;
  assign new_n3333_ = v19 & v25;
  assign new_n3334_ = new_n882_ & new_n3333_;
  assign new_n3335_ = new_n3332_ & new_n3334_;
  assign new_n3336_ = v2 & new_n585_;
  assign new_n3337_ = ~v8 & ~v25;
  assign new_n3338_ = ~v7 & new_n3337_;
  assign new_n3339_ = new_n3336_ & new_n3338_;
  assign new_n3340_ = ~new_n3335_ & ~new_n3339_;
  assign new_n3341_ = ~v10 & ~new_n3340_;
  assign new_n3342_ = v7 & new_n368_;
  assign new_n3343_ = ~new_n1118_ & ~new_n3342_;
  assign new_n3344_ = v6 & ~new_n3343_;
  assign new_n3345_ = ~v2 & new_n3344_;
  assign new_n3346_ = new_n358_ & new_n1162_;
  assign new_n3347_ = ~new_n3345_ & ~new_n3346_;
  assign new_n3348_ = ~v5 & ~new_n3347_;
  assign new_n3349_ = ~v2 & new_n546_;
  assign new_n3350_ = new_n1118_ & new_n3349_;
  assign new_n3351_ = ~new_n3348_ & ~new_n3350_;
  assign new_n3352_ = ~v25 & ~new_n3351_;
  assign new_n3353_ = v10 & new_n3352_;
  assign new_n3354_ = ~new_n3341_ & ~new_n3353_;
  assign new_n3355_ = ~v3 & ~new_n3354_;
  assign new_n3356_ = v2 & new_n3342_;
  assign new_n3357_ = v8 & new_n398_;
  assign new_n3358_ = new_n875_ & new_n3357_;
  assign new_n3359_ = ~new_n3356_ & ~new_n3358_;
  assign new_n3360_ = v6 & ~new_n3359_;
  assign new_n3361_ = ~v2 & new_n2412_;
  assign new_n3362_ = new_n3357_ & new_n3361_;
  assign new_n3363_ = ~new_n3360_ & ~new_n3362_;
  assign new_n3364_ = ~v25 & ~new_n3363_;
  assign new_n3365_ = v5 & new_n3364_;
  assign new_n3366_ = new_n533_ & new_n2944_;
  assign new_n3367_ = new_n321_ & new_n430_;
  assign new_n3368_ = new_n3366_ & new_n3367_;
  assign new_n3369_ = ~new_n3365_ & ~new_n3368_;
  assign new_n3370_ = v3 & ~new_n3369_;
  assign new_n3371_ = ~new_n3355_ & ~new_n3370_;
  assign new_n3372_ = ~v4 & ~new_n3371_;
  assign new_n3373_ = v25 & ~new_n1333_;
  assign new_n3374_ = ~v10 & new_n3373_;
  assign new_n3375_ = ~v5 & new_n3374_;
  assign new_n3376_ = ~v2 & new_n3375_;
  assign new_n3377_ = v6 & new_n882_;
  assign new_n3378_ = ~new_n148_ & ~new_n3377_;
  assign new_n3379_ = ~v25 & ~new_n3378_;
  assign new_n3380_ = v10 & new_n3379_;
  assign new_n3381_ = v5 & new_n3380_;
  assign new_n3382_ = v2 & new_n3381_;
  assign new_n3383_ = ~new_n3376_ & ~new_n3382_;
  assign new_n3384_ = ~v9 & ~new_n3383_;
  assign new_n3385_ = new_n1046_ & new_n2329_;
  assign new_n3386_ = new_n257_ & new_n433_;
  assign new_n3387_ = new_n3385_ & new_n3386_;
  assign new_n3388_ = ~new_n3384_ & ~new_n3387_;
  assign new_n3389_ = v3 & ~new_n3388_;
  assign new_n3390_ = new_n138_ & new_n713_;
  assign new_n3391_ = new_n1331_ & new_n3295_;
  assign new_n3392_ = new_n3390_ & new_n3391_;
  assign new_n3393_ = ~new_n3389_ & ~new_n3392_;
  assign new_n3394_ = v4 & ~new_n3393_;
  assign new_n3395_ = ~new_n3372_ & ~new_n3394_;
  assign new_n3396_ = ~v1 & ~new_n3395_;
  assign new_n3397_ = new_n853_ & new_n2451_;
  assign new_n3398_ = v9 & new_n322_;
  assign new_n3399_ = new_n3042_ & new_n3398_;
  assign new_n3400_ = new_n3397_ & new_n3399_;
  assign new_n3401_ = ~new_n3396_ & ~new_n3400_;
  assign new_n3402_ = ~v23 & ~new_n3401_;
  assign new_n3403_ = v23 & new_n84_;
  assign new_n3404_ = v9 & new_n3403_;
  assign new_n3405_ = ~v8 & new_n3404_;
  assign new_n3406_ = v4 & new_n3405_;
  assign new_n3407_ = v3 & new_n3406_;
  assign new_n3408_ = v2 & new_n3407_;
  assign new_n3409_ = v1 & new_n3408_;
  assign new_n3410_ = ~new_n3402_ & ~new_n3409_;
  assign new_n3411_ = ~v24 & ~new_n3410_;
  assign new_n3412_ = ~v2 & ~new_n2796_;
  assign new_n3413_ = new_n145_ & new_n418_;
  assign new_n3414_ = ~v10 & v19;
  assign new_n3415_ = new_n1094_ & new_n3414_;
  assign new_n3416_ = new_n3413_ & new_n3415_;
  assign new_n3417_ = ~new_n3412_ & ~new_n3416_;
  assign new_n3418_ = ~v25 & ~new_n3417_;
  assign new_n3419_ = ~v23 & new_n3418_;
  assign new_n3420_ = v6 & new_n3419_;
  assign new_n3421_ = v23 & v25;
  assign new_n3422_ = v19 & new_n3421_;
  assign new_n3423_ = v10 & new_n3422_;
  assign new_n3424_ = v9 & new_n3423_;
  assign new_n3425_ = ~v6 & new_n3424_;
  assign new_n3426_ = v5 & new_n3425_;
  assign new_n3427_ = ~v3 & new_n3426_;
  assign new_n3428_ = v2 & new_n3427_;
  assign new_n3429_ = ~v1 & new_n3428_;
  assign new_n3430_ = ~new_n3420_ & ~new_n3429_;
  assign new_n3431_ = v24 & ~new_n3430_;
  assign new_n3432_ = ~v8 & new_n3431_;
  assign new_n3433_ = v4 & new_n3432_;
  assign new_n3434_ = ~new_n3411_ & ~new_n3433_;
  assign new_n3435_ = ~v22 & ~new_n3434_;
  assign \v26.35  = ~v0 & new_n3435_;
  assign new_n3437_ = v25 & ~new_n1421_;
  assign new_n3438_ = ~v10 & new_n3437_;
  assign new_n3439_ = ~v1 & new_n3438_;
  assign new_n3440_ = v0 & new_n3439_;
  assign new_n3441_ = v1 & ~v8;
  assign new_n3442_ = ~v0 & new_n3441_;
  assign new_n3443_ = new_n1029_ & new_n3442_;
  assign new_n3444_ = ~new_n3440_ & ~new_n3443_;
  assign new_n3445_ = v6 & ~new_n3444_;
  assign new_n3446_ = ~v8 & new_n616_;
  assign new_n3447_ = ~v6 & new_n3446_;
  assign new_n3448_ = v1 & new_n3447_;
  assign new_n3449_ = ~v0 & new_n3448_;
  assign new_n3450_ = ~new_n3445_ & ~new_n3449_;
  assign new_n3451_ = v7 & ~new_n3450_;
  assign new_n3452_ = v9 & new_n932_;
  assign new_n3453_ = ~v8 & new_n3452_;
  assign new_n3454_ = ~v7 & new_n3453_;
  assign new_n3455_ = v1 & new_n3454_;
  assign new_n3456_ = ~v0 & new_n3455_;
  assign new_n3457_ = ~new_n3451_ & ~new_n3456_;
  assign new_n3458_ = ~v5 & ~new_n3457_;
  assign new_n3459_ = ~v7 & new_n257_;
  assign new_n3460_ = ~new_n952_ & ~new_n3459_;
  assign new_n3461_ = v6 & ~new_n3460_;
  assign new_n3462_ = ~v6 & new_n1094_;
  assign new_n3463_ = ~new_n3461_ & ~new_n3462_;
  assign new_n3464_ = ~v1 & ~new_n3463_;
  assign new_n3465_ = v1 & ~v6;
  assign new_n3466_ = new_n3459_ & new_n3465_;
  assign new_n3467_ = ~new_n3464_ & ~new_n3466_;
  assign new_n3468_ = v10 & ~new_n3467_;
  assign new_n3469_ = ~v7 & new_n301_;
  assign new_n3470_ = v1 & new_n3469_;
  assign new_n3471_ = ~new_n3468_ & ~new_n3470_;
  assign new_n3472_ = ~v25 & ~new_n3471_;
  assign new_n3473_ = v5 & new_n3472_;
  assign new_n3474_ = ~v0 & new_n3473_;
  assign new_n3475_ = ~new_n3458_ & ~new_n3474_;
  assign new_n3476_ = v2 & ~new_n3475_;
  assign new_n3477_ = ~v10 & ~new_n1333_;
  assign new_n3478_ = ~v1 & new_n3477_;
  assign new_n3479_ = v1 & v6;
  assign new_n3480_ = v7 & new_n767_;
  assign new_n3481_ = new_n3479_ & new_n3480_;
  assign new_n3482_ = ~new_n3478_ & ~new_n3481_;
  assign new_n3483_ = v25 & ~new_n3482_;
  assign new_n3484_ = ~v9 & new_n3483_;
  assign new_n3485_ = ~v5 & new_n3484_;
  assign new_n3486_ = ~v2 & new_n3485_;
  assign new_n3487_ = ~v0 & new_n3486_;
  assign new_n3488_ = ~new_n3476_ & ~new_n3487_;
  assign new_n3489_ = v4 & ~new_n3488_;
  assign new_n3490_ = ~v1 & ~new_n3369_;
  assign new_n3491_ = new_n585_ & new_n853_;
  assign new_n3492_ = new_n1125_ & new_n3398_;
  assign new_n3493_ = new_n3491_ & new_n3492_;
  assign new_n3494_ = ~new_n3490_ & ~new_n3493_;
  assign new_n3495_ = ~v4 & ~new_n3494_;
  assign new_n3496_ = ~v0 & new_n3495_;
  assign new_n3497_ = ~new_n3489_ & ~new_n3496_;
  assign new_n3498_ = v3 & ~new_n3497_;
  assign new_n3499_ = ~v2 & new_n117_;
  assign new_n3500_ = new_n632_ & new_n1125_;
  assign new_n3501_ = new_n3499_ & new_n3500_;
  assign new_n3502_ = new_n3340_ & ~new_n3501_;
  assign new_n3503_ = ~v10 & ~new_n3502_;
  assign new_n3504_ = ~new_n3353_ & ~new_n3503_;
  assign new_n3505_ = ~v4 & ~new_n3504_;
  assign new_n3506_ = new_n138_ & new_n346_;
  assign new_n3507_ = new_n3391_ & new_n3506_;
  assign new_n3508_ = ~new_n3505_ & ~new_n3507_;
  assign new_n3509_ = ~v3 & ~new_n3508_;
  assign new_n3510_ = ~v1 & new_n3509_;
  assign new_n3511_ = ~v0 & new_n3510_;
  assign new_n3512_ = ~new_n3498_ & ~new_n3511_;
  assign new_n3513_ = ~v23 & ~new_n3512_;
  assign new_n3514_ = ~v0 & new_n3409_;
  assign new_n3515_ = ~new_n3513_ & ~new_n3514_;
  assign new_n3516_ = ~v24 & ~new_n3515_;
  assign new_n3517_ = ~v0 & new_n3433_;
  assign new_n3518_ = ~new_n3516_ & ~new_n3517_;
  assign \v26.36  = ~v22 & ~new_n3518_;
  assign new_n3520_ = ~v23 & ~new_n3475_;
  assign new_n3521_ = v1 & new_n3405_;
  assign new_n3522_ = ~v0 & new_n3521_;
  assign new_n3523_ = ~new_n3520_ & ~new_n3522_;
  assign new_n3524_ = v4 & ~new_n3523_;
  assign new_n3525_ = ~v1 & new_n179_;
  assign new_n3526_ = ~v0 & new_n3525_;
  assign new_n3527_ = ~new_n3524_ & ~new_n3526_;
  assign new_n3528_ = v2 & ~new_n3527_;
  assign new_n3529_ = v4 & new_n882_;
  assign new_n3530_ = new_n3232_ & new_n3529_;
  assign new_n3531_ = ~v4 & new_n1125_;
  assign new_n3532_ = new_n3398_ & new_n3531_;
  assign new_n3533_ = ~new_n3530_ & ~new_n3532_;
  assign new_n3534_ = ~v5 & ~new_n3533_;
  assign new_n3535_ = v1 & new_n3534_;
  assign new_n3536_ = new_n73_ & new_n829_;
  assign new_n3537_ = new_n310_ & new_n433_;
  assign new_n3538_ = new_n3536_ & new_n3537_;
  assign new_n3539_ = ~new_n3535_ & ~new_n3538_;
  assign new_n3540_ = v6 & ~new_n3539_;
  assign new_n3541_ = new_n138_ & new_n829_;
  assign new_n3542_ = new_n882_ & new_n1029_;
  assign new_n3543_ = new_n3541_ & new_n3542_;
  assign new_n3544_ = ~new_n3540_ & ~new_n3543_;
  assign new_n3545_ = ~v23 & ~new_n3544_;
  assign new_n3546_ = ~v2 & new_n3545_;
  assign new_n3547_ = ~v0 & new_n3546_;
  assign new_n3548_ = ~new_n3528_ & ~new_n3547_;
  assign new_n3549_ = v3 & ~new_n3548_;
  assign new_n3550_ = v2 & new_n347_;
  assign new_n3551_ = new_n398_ & new_n656_;
  assign new_n3552_ = ~new_n3550_ & ~new_n3551_;
  assign new_n3553_ = ~v5 & ~new_n3552_;
  assign new_n3554_ = new_n2475_ & new_n3357_;
  assign new_n3555_ = ~new_n3553_ & ~new_n3554_;
  assign new_n3556_ = ~v7 & ~new_n3555_;
  assign new_n3557_ = v6 & new_n3556_;
  assign new_n3558_ = v2 & new_n117_;
  assign new_n3559_ = new_n398_ & new_n1331_;
  assign new_n3560_ = new_n3558_ & new_n3559_;
  assign new_n3561_ = ~new_n3557_ & ~new_n3560_;
  assign new_n3562_ = ~v25 & ~new_n3561_;
  assign new_n3563_ = ~v23 & new_n3562_;
  assign new_n3564_ = ~v4 & new_n3563_;
  assign new_n3565_ = ~v3 & new_n3564_;
  assign new_n3566_ = ~v1 & new_n3565_;
  assign new_n3567_ = ~v0 & new_n3566_;
  assign new_n3568_ = ~new_n3549_ & ~new_n3567_;
  assign new_n3569_ = ~v24 & ~new_n3568_;
  assign new_n3570_ = v10 & new_n3421_;
  assign new_n3571_ = v9 & new_n3570_;
  assign new_n3572_ = ~v6 & new_n3571_;
  assign new_n3573_ = v6 & new_n1094_;
  assign new_n3574_ = new_n3043_ & new_n3573_;
  assign new_n3575_ = ~new_n3572_ & ~new_n3574_;
  assign new_n3576_ = v24 & ~new_n3575_;
  assign new_n3577_ = v19 & new_n3576_;
  assign new_n3578_ = ~v8 & new_n3577_;
  assign new_n3579_ = v5 & new_n3578_;
  assign new_n3580_ = v4 & new_n3579_;
  assign new_n3581_ = ~v3 & new_n3580_;
  assign new_n3582_ = v2 & new_n3581_;
  assign new_n3583_ = ~v1 & new_n3582_;
  assign new_n3584_ = ~v0 & new_n3583_;
  assign new_n3585_ = ~new_n3569_ & ~new_n3584_;
  assign \v26.37  = ~v22 & ~new_n3585_;
  assign new_n3587_ = v25 & ~new_n83_;
  assign new_n3588_ = v24 & new_n3587_;
  assign new_n3589_ = ~v23 & new_n3588_;
  assign new_n3590_ = ~v22 & new_n3589_;
  assign new_n3591_ = v9 & new_n3590_;
  assign new_n3592_ = ~v8 & new_n3591_;
  assign new_n3593_ = v4 & new_n3592_;
  assign new_n3594_ = v3 & new_n3593_;
  assign new_n3595_ = v2 & new_n3594_;
  assign new_n3596_ = v1 & new_n3595_;
  assign \v26.39  = ~v0 & new_n3596_;
  assign new_n3598_ = v24 & ~new_n716_;
  assign new_n3599_ = v23 & new_n3598_;
  assign new_n3600_ = ~v10 & new_n3599_;
  assign new_n3601_ = ~v9 & new_n3600_;
  assign new_n3602_ = ~v8 & new_n3601_;
  assign new_n3603_ = v7 & new_n3602_;
  assign new_n3604_ = v6 & new_n3603_;
  assign new_n3605_ = ~v4 & new_n3604_;
  assign new_n3606_ = v0 & new_n3605_;
  assign new_n3607_ = ~v3 & new_n1026_;
  assign new_n3608_ = new_n545_ & new_n3607_;
  assign new_n3609_ = new_n1118_ & new_n2766_;
  assign new_n3610_ = new_n3608_ & new_n3609_;
  assign new_n3611_ = ~new_n3606_ & ~new_n3610_;
  assign new_n3612_ = ~v25 & ~new_n3611_;
  assign new_n3613_ = ~v22 & new_n3612_;
  assign \v26.40  = ~v5 & new_n3613_;
  assign new_n3615_ = ~v22 & new_n2459_;
  assign new_n3616_ = ~v10 & new_n3615_;
  assign new_n3617_ = ~v9 & new_n3616_;
  assign new_n3618_ = ~v8 & new_n3617_;
  assign new_n3619_ = v7 & new_n3618_;
  assign new_n3620_ = v6 & new_n3619_;
  assign new_n3621_ = ~v5 & new_n3620_;
  assign new_n3622_ = ~v4 & new_n3621_;
  assign \v26.41  = v0 & new_n3622_;
  assign new_n3624_ = v24 & ~new_n81_;
  assign new_n3625_ = ~v23 & new_n3624_;
  assign new_n3626_ = ~v22 & new_n3625_;
  assign new_n3627_ = v9 & new_n3626_;
  assign new_n3628_ = ~v8 & new_n3627_;
  assign new_n3629_ = v6 & new_n3628_;
  assign new_n3630_ = v4 & new_n3629_;
  assign new_n3631_ = v3 & new_n3630_;
  assign new_n3632_ = v2 & new_n3631_;
  assign new_n3633_ = v1 & new_n3632_;
  assign \v26.42  = ~v0 & new_n3633_;
  assign new_n3635_ = ~v23 & new_n2257_;
  assign new_n3636_ = ~v22 & new_n3635_;
  assign new_n3637_ = ~v10 & new_n3636_;
  assign new_n3638_ = v9 & new_n3637_;
  assign new_n3639_ = v8 & new_n3638_;
  assign new_n3640_ = ~v7 & new_n3639_;
  assign new_n3641_ = v6 & new_n3640_;
  assign new_n3642_ = ~v5 & new_n3641_;
  assign new_n3643_ = ~v4 & new_n3642_;
  assign \v26.43  = v0 & new_n3643_;
  assign new_n3645_ = v4 & new_n645_;
  assign new_n3646_ = v1 & new_n3645_;
  assign new_n3647_ = v0 & new_n3646_;
  assign new_n3648_ = new_n95_ & new_n236_;
  assign new_n3649_ = new_n148_ & new_n454_;
  assign new_n3650_ = new_n3648_ & new_n3649_;
  assign new_n3651_ = ~new_n3647_ & ~new_n3650_;
  assign new_n3652_ = v3 & ~new_n3651_;
  assign new_n3653_ = ~v2 & new_n3652_;
  assign new_n3654_ = ~v5 & new_n2412_;
  assign new_n3655_ = new_n953_ & new_n3654_;
  assign new_n3656_ = new_n2720_ & new_n3655_;
  assign new_n3657_ = ~new_n3653_ & ~new_n3656_;
  assign new_n3658_ = v9 & ~new_n3657_;
  assign new_n3659_ = v7 & new_n1788_;
  assign new_n3660_ = v6 & new_n3659_;
  assign new_n3661_ = ~v5 & new_n3660_;
  assign new_n3662_ = v4 & new_n3661_;
  assign new_n3663_ = v3 & new_n3662_;
  assign new_n3664_ = ~v2 & new_n3663_;
  assign new_n3665_ = v1 & new_n3664_;
  assign new_n3666_ = v0 & new_n3665_;
  assign new_n3667_ = ~new_n3658_ & ~new_n3666_;
  assign new_n3668_ = ~v8 & ~new_n3667_;
  assign new_n3669_ = v7 & new_n1520_;
  assign new_n3670_ = v6 & new_n3669_;
  assign new_n3671_ = ~v5 & new_n3670_;
  assign new_n3672_ = v4 & new_n3671_;
  assign new_n3673_ = v3 & new_n3672_;
  assign new_n3674_ = ~v2 & new_n3673_;
  assign new_n3675_ = v1 & new_n3674_;
  assign new_n3676_ = v0 & new_n3675_;
  assign new_n3677_ = ~new_n3668_ & ~new_n3676_;
  assign new_n3678_ = ~v23 & ~new_n3677_;
  assign \v26.44  = ~v22 & new_n3678_;
  assign new_n3680_ = new_n292_ & new_n430_;
  assign new_n3681_ = new_n2973_ & new_n3680_;
  assign new_n3682_ = new_n95_ & new_n712_;
  assign new_n3683_ = new_n382_ & new_n433_;
  assign new_n3684_ = new_n3682_ & new_n3683_;
  assign new_n3685_ = ~new_n3681_ & ~new_n3684_;
  assign new_n3686_ = ~v2 & new_n273_;
  assign new_n3687_ = ~v2 & ~new_n3686_;
  assign new_n3688_ = v25 & ~new_n3687_;
  assign new_n3689_ = ~v10 & new_n3688_;
  assign new_n3690_ = ~v9 & new_n3689_;
  assign new_n3691_ = v6 & new_n3690_;
  assign new_n3692_ = v1 & new_n3691_;
  assign new_n3693_ = v0 & new_n3692_;
  assign new_n3694_ = new_n3685_ & ~new_n3693_;
  assign new_n3695_ = v7 & ~new_n3694_;
  assign new_n3696_ = ~v10 & new_n1360_;
  assign new_n3697_ = v9 & new_n3696_;
  assign new_n3698_ = v8 & new_n3697_;
  assign new_n3699_ = ~v7 & new_n3698_;
  assign new_n3700_ = v6 & new_n3699_;
  assign new_n3701_ = v1 & new_n3700_;
  assign new_n3702_ = v0 & new_n3701_;
  assign new_n3703_ = ~new_n3695_ & ~new_n3702_;
  assign new_n3704_ = ~v4 & ~new_n3703_;
  assign new_n3705_ = ~new_n547_ & ~new_n2921_;
  assign new_n3706_ = ~v6 & ~new_n3705_;
  assign new_n3707_ = new_n78_ & ~new_n3706_;
  assign new_n3708_ = v25 & ~new_n3707_;
  assign new_n3709_ = v9 & new_n3708_;
  assign new_n3710_ = ~v8 & new_n3709_;
  assign new_n3711_ = v4 & new_n3710_;
  assign new_n3712_ = v3 & new_n3711_;
  assign new_n3713_ = v2 & new_n3712_;
  assign new_n3714_ = v1 & new_n3713_;
  assign new_n3715_ = ~v0 & new_n3714_;
  assign new_n3716_ = ~new_n3704_ & ~new_n3715_;
  assign new_n3717_ = ~v5 & ~new_n3716_;
  assign new_n3718_ = ~v3 & v10;
  assign new_n3719_ = ~v1 & new_n3718_;
  assign new_n3720_ = ~new_n1943_ & ~new_n3719_;
  assign new_n3721_ = ~v7 & ~new_n3720_;
  assign new_n3722_ = new_n76_ & new_n589_;
  assign new_n3723_ = ~new_n3721_ & ~new_n3722_;
  assign new_n3724_ = ~v6 & ~new_n3723_;
  assign new_n3725_ = v6 & new_n77_;
  assign new_n3726_ = new_n1943_ & new_n3725_;
  assign new_n3727_ = ~new_n3724_ & ~new_n3726_;
  assign new_n3728_ = ~v8 & ~new_n3727_;
  assign new_n3729_ = v4 & new_n3728_;
  assign new_n3730_ = ~v0 & new_n3729_;
  assign new_n3731_ = new_n239_ & new_n533_;
  assign new_n3732_ = new_n1867_ & new_n3731_;
  assign new_n3733_ = ~new_n3730_ & ~new_n3732_;
  assign new_n3734_ = v25 & ~new_n3733_;
  assign new_n3735_ = v9 & new_n3734_;
  assign new_n3736_ = v5 & new_n3735_;
  assign new_n3737_ = v2 & new_n3736_;
  assign new_n3738_ = ~new_n3717_ & ~new_n3737_;
  assign new_n3739_ = ~v24 & ~new_n3738_;
  assign new_n3740_ = ~v23 & new_n3739_;
  assign \v26.45  = ~v22 & new_n3740_;
  assign \v26.38  = \v26.32 ;
endmodule


