// Benchmark "ttt2" written by ABC on Fri Feb 25 15:12:27 2022

module ttt2 ( 
    a, b, c, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0,
    r0, s0, t0  );
  input  a, b, c, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v,
    w, x, y;
  output z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0,
    q0, r0, s0, t0;
  wire new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_,
    new_n53_, new_n54_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_,
    new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_,
    new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_,
    new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_,
    new_n98_, new_n99_, new_n100_, new_n101_, new_n102_, new_n103_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_, new_n142_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n252_, new_n253_, new_n254_, new_n256_, new_n257_,
    new_n258_, new_n260_, new_n261_, new_n262_;
  assign new_n46_ = s & ~t;
  assign new_n47_ = ~e & ~new_n46_;
  assign new_n48_ = ~t & ~u;
  assign new_n49_ = ~s & new_n48_;
  assign new_n50_ = ~new_n47_ & ~new_n49_;
  assign new_n51_ = v & ~new_n50_;
  assign new_n52_ = e & v;
  assign new_n53_ = u & ~new_n52_;
  assign new_n54_ = ~new_n51_ & ~new_n53_;
  assign z = ~w & new_n54_;
  assign new_n56_ = ~v & ~y;
  assign new_n57_ = ~u & v;
  assign new_n58_ = ~v & y;
  assign new_n59_ = u & new_n58_;
  assign new_n60_ = ~new_n57_ & ~new_n59_;
  assign new_n61_ = ~s & ~new_n60_;
  assign new_n62_ = ~t & new_n61_;
  assign new_n63_ = f & ~new_n48_;
  assign new_n64_ = v & new_n63_;
  assign new_n65_ = ~new_n62_ & ~new_n64_;
  assign new_n66_ = v & ~w;
  assign new_n67_ = q & ~new_n66_;
  assign new_n68_ = ~w & new_n65_;
  assign new_n69_ = ~t & u;
  assign new_n70_ = s & new_n56_;
  assign new_n71_ = new_n69_ & new_n70_;
  assign new_n72_ = ~new_n68_ & ~new_n71_;
  assign a0 = ~new_n67_ & new_n72_;
  assign new_n74_ = new_n46_ & new_n56_;
  assign new_n75_ = ~s & new_n58_;
  assign new_n76_ = u & ~new_n75_;
  assign new_n77_ = ~t & ~new_n76_;
  assign new_n78_ = ~u & ~v;
  assign new_n79_ = ~g & v;
  assign new_n80_ = ~new_n78_ & ~new_n79_;
  assign new_n81_ = ~new_n77_ & new_n80_;
  assign new_n82_ = w & ~new_n74_;
  assign b0 = new_n81_ & ~new_n82_;
  assign new_n84_ = ~q & w;
  assign new_n85_ = u & v;
  assign new_n86_ = u & ~v;
  assign new_n87_ = t & ~new_n86_;
  assign new_n88_ = ~new_n85_ & ~new_n87_;
  assign new_n89_ = ~w & new_n78_;
  assign new_n90_ = ~s & ~t;
  assign new_n91_ = q & new_n58_;
  assign new_n92_ = new_n90_ & new_n91_;
  assign new_n93_ = ~new_n89_ & ~new_n92_;
  assign new_n94_ = q & ~new_n74_;
  assign new_n95_ = ~h & ~new_n88_;
  assign new_n96_ = ~w & new_n95_;
  assign new_n97_ = ~u & ~new_n84_;
  assign new_n98_ = new_n46_ & new_n97_;
  assign new_n99_ = ~new_n96_ & ~new_n98_;
  assign new_n100_ = ~new_n94_ & new_n99_;
  assign new_n101_ = ~new_n95_ & ~new_n98_;
  assign new_n102_ = ~w & new_n101_;
  assign new_n103_ = ~new_n100_ & ~new_n102_;
  assign c0 = new_n93_ & ~new_n103_;
  assign new_n105_ = s & ~u;
  assign new_n106_ = ~v & ~new_n105_;
  assign new_n107_ = ~i & v;
  assign new_n108_ = ~new_n48_ & ~new_n107_;
  assign new_n109_ = ~new_n106_ & new_n108_;
  assign d0 = ~w & new_n109_;
  assign new_n111_ = t & v;
  assign new_n112_ = ~u & ~new_n111_;
  assign new_n113_ = ~j & ~new_n112_;
  assign new_n114_ = new_n57_ & new_n90_;
  assign new_n115_ = t & ~v;
  assign new_n116_ = s & new_n115_;
  assign new_n117_ = ~new_n114_ & ~new_n116_;
  assign new_n118_ = ~new_n113_ & new_n117_;
  assign new_n119_ = ~new_n86_ & new_n118_;
  assign e0 = ~w & new_n119_;
  assign f0 = ~a & ~k;
  assign new_n122_ = ~m & n;
  assign new_n123_ = ~l & ~new_n122_;
  assign new_n124_ = k & new_n123_;
  assign new_n125_ = ~k & l;
  assign new_n126_ = ~new_n124_ & ~new_n125_;
  assign g0 = ~a & ~new_n126_;
  assign new_n128_ = k & l;
  assign new_n129_ = m & ~new_n128_;
  assign new_n130_ = l & ~m;
  assign new_n131_ = k & new_n130_;
  assign new_n132_ = ~new_n129_ & ~new_n131_;
  assign h0 = ~a & ~new_n132_;
  assign new_n134_ = l & m;
  assign new_n135_ = k & new_n134_;
  assign new_n136_ = ~l & ~m;
  assign new_n137_ = m & n;
  assign new_n138_ = l & new_n137_;
  assign new_n139_ = ~new_n136_ & ~new_n138_;
  assign new_n140_ = k & ~new_n139_;
  assign new_n141_ = ~a & ~new_n140_;
  assign new_n142_ = ~n & ~new_n135_;
  assign i0 = new_n141_ & ~new_n142_;
  assign new_n144_ = n & o;
  assign new_n145_ = k & ~l;
  assign new_n146_ = new_n122_ & new_n145_;
  assign new_n147_ = ~x & ~new_n146_;
  assign new_n148_ = ~o & ~new_n147_;
  assign new_n149_ = ~o & ~new_n146_;
  assign new_n150_ = ~x & ~new_n149_;
  assign new_n151_ = ~new_n148_ & ~new_n150_;
  assign new_n152_ = ~m & new_n144_;
  assign new_n153_ = new_n145_ & new_n152_;
  assign new_n154_ = ~new_n151_ & ~new_n153_;
  assign j0 = ~a & new_n154_;
  assign new_n156_ = ~q & r;
  assign new_n157_ = ~p & ~new_n156_;
  assign new_n158_ = x & ~new_n157_;
  assign new_n159_ = o & new_n158_;
  assign new_n160_ = ~o & ~p;
  assign new_n161_ = ~a & ~new_n160_;
  assign new_n162_ = ~new_n159_ & new_n161_;
  assign new_n163_ = ~p & ~new_n146_;
  assign new_n164_ = ~x & new_n163_;
  assign new_n165_ = new_n152_ & ~new_n157_;
  assign new_n166_ = new_n145_ & new_n165_;
  assign new_n167_ = ~new_n164_ & ~new_n166_;
  assign k0 = new_n162_ & new_n167_;
  assign new_n169_ = o & p;
  assign new_n170_ = ~q & ~new_n169_;
  assign new_n171_ = ~a & ~new_n170_;
  assign new_n172_ = q & ~new_n147_;
  assign new_n173_ = new_n169_ & new_n172_;
  assign new_n174_ = ~new_n147_ & ~new_n173_;
  assign new_n175_ = p & ~new_n147_;
  assign new_n176_ = o & new_n175_;
  assign new_n177_ = q & ~new_n176_;
  assign new_n178_ = ~new_n174_ & ~new_n177_;
  assign l0 = new_n171_ & ~new_n178_;
  assign new_n180_ = ~p & ~q;
  assign new_n181_ = q & r;
  assign new_n182_ = p & new_n181_;
  assign new_n183_ = ~new_n180_ & ~new_n182_;
  assign new_n184_ = p & q;
  assign new_n185_ = o & new_n184_;
  assign new_n186_ = ~r & ~new_n185_;
  assign new_n187_ = ~a & ~new_n186_;
  assign new_n188_ = ~r & ~new_n146_;
  assign new_n189_ = ~x & new_n188_;
  assign new_n190_ = ~l & new_n152_;
  assign new_n191_ = k & new_n190_;
  assign new_n192_ = ~o & ~new_n191_;
  assign new_n193_ = ~new_n183_ & ~new_n192_;
  assign new_n194_ = ~new_n189_ & ~new_n193_;
  assign new_n195_ = ~new_n188_ & ~new_n191_;
  assign new_n196_ = ~x & new_n195_;
  assign new_n197_ = ~new_n194_ & ~new_n196_;
  assign m0 = new_n187_ & ~new_n197_;
  assign new_n199_ = r & s;
  assign new_n200_ = ~q & new_n199_;
  assign new_n201_ = ~new_n147_ & new_n156_;
  assign new_n202_ = o & ~p;
  assign new_n203_ = new_n201_ & new_n202_;
  assign new_n204_ = ~s & ~new_n203_;
  assign new_n205_ = ~new_n147_ & new_n200_;
  assign new_n206_ = new_n202_ & new_n205_;
  assign new_n207_ = ~new_n204_ & ~new_n206_;
  assign n0 = ~a & new_n207_;
  assign new_n209_ = new_n46_ & new_n156_;
  assign new_n210_ = ~l & new_n122_;
  assign new_n211_ = k & new_n210_;
  assign new_n212_ = ~x & ~new_n211_;
  assign new_n213_ = ~new_n57_ & ~new_n212_;
  assign new_n214_ = o & ~q;
  assign new_n215_ = new_n199_ & new_n214_;
  assign new_n216_ = ~new_n147_ & new_n215_;
  assign new_n217_ = ~p & new_n216_;
  assign new_n218_ = new_n209_ & new_n213_;
  assign new_n219_ = new_n202_ & new_n218_;
  assign new_n220_ = t & ~new_n217_;
  assign new_n221_ = ~new_n219_ & ~new_n220_;
  assign o0 = ~a & ~new_n221_;
  assign new_n223_ = o & new_n180_;
  assign new_n224_ = t & ~u;
  assign new_n225_ = new_n199_ & new_n224_;
  assign new_n226_ = o & r;
  assign new_n227_ = s & t;
  assign new_n228_ = new_n226_ & new_n227_;
  assign new_n229_ = ~new_n147_ & new_n228_;
  assign new_n230_ = ~q & new_n229_;
  assign new_n231_ = ~p & new_n230_;
  assign new_n232_ = ~new_n147_ & new_n225_;
  assign new_n233_ = new_n223_ & new_n232_;
  assign new_n234_ = u & ~new_n231_;
  assign new_n235_ = ~new_n233_ & ~new_n234_;
  assign p0 = ~a & ~new_n235_;
  assign new_n237_ = new_n156_ & new_n202_;
  assign new_n238_ = new_n86_ & new_n227_;
  assign new_n239_ = t & u;
  assign new_n240_ = ~new_n48_ & ~new_n239_;
  assign new_n241_ = r & ~new_n240_;
  assign new_n242_ = s & new_n241_;
  assign new_n243_ = o & new_n242_;
  assign new_n244_ = ~new_n147_ & new_n243_;
  assign new_n245_ = ~q & new_n244_;
  assign new_n246_ = ~p & new_n245_;
  assign new_n247_ = new_n237_ & new_n238_;
  assign new_n248_ = ~new_n147_ & new_n247_;
  assign new_n249_ = v & ~new_n246_;
  assign new_n250_ = ~new_n248_ & ~new_n249_;
  assign q0 = ~a & ~new_n250_;
  assign new_n252_ = new_n69_ & new_n75_;
  assign new_n253_ = ~w & ~new_n252_;
  assign new_n254_ = ~new_n71_ & ~new_n253_;
  assign r0 = ~a & new_n254_;
  assign new_n256_ = b & ~x;
  assign new_n257_ = ~b & x;
  assign new_n258_ = ~new_n256_ & ~new_n257_;
  assign s0 = ~a & ~new_n258_;
  assign new_n260_ = c & ~y;
  assign new_n261_ = ~c & y;
  assign new_n262_ = ~new_n260_ & ~new_n261_;
  assign t0 = ~a & ~new_n262_;
endmodule


