// Benchmark "max" written by ABC on Tue Sep  5 18:12:16 2023

module max ( 
    \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] , \in0[6] ,
    \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] , \in0[12] ,
    \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] , \in0[18] ,
    \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] , \in0[24] ,
    \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] , \in0[30] ,
    \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] , \in0[36] ,
    \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] , \in0[42] ,
    \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] , \in0[48] ,
    \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] , \in0[54] ,
    \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] ,
    \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] ,
    \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72] ,
    \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] , \in0[78] ,
    \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] , \in0[84] ,
    \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] , \in0[90] ,
    \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] , \in0[96] ,
    \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] , \in0[102] ,
    \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] , \in0[108] ,
    \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] ,
    \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] , \in0[120] ,
    \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] ,
    \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] ,
    \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] ,
    \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] ,
    \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] , \in1[23] ,
    \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] ,
    \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] , \in1[35] ,
    \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] ,
    \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] ,
    \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53] ,
    \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] , \in1[59] ,
    \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] , \in1[65] ,
    \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] , \in1[71] ,
    \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] , \in1[77] ,
    \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] , \in1[83] ,
    \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] , \in1[89] ,
    \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] , \in1[95] ,
    \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] , \in1[101] ,
    \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] ,
    \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] , \in1[113] ,
    \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] , \in1[119] ,
    \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] ,
    \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] ,
    \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] ,
    \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] ,
    \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] ,
    \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] ,
    \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] , \in2[34] ,
    \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] , \in2[40] ,
    \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] , \in2[46] ,
    \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] , \in2[52] ,
    \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] , \in2[58] ,
    \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] , \in2[64] ,
    \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] , \in2[70] ,
    \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] , \in2[76] ,
    \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] ,
    \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] ,
    \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94] ,
    \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] , \in2[100] ,
    \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] , \in2[106] ,
    \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] , \in2[112] ,
    \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] , \in2[118] ,
    \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
    \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] ,
    \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] , \in3[9] ,
    \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] , \in3[15] ,
    \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] , \in3[21] ,
    \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] , \in3[27] ,
    \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] , \in3[33] ,
    \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] , \in3[39] ,
    \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] , \in3[45] ,
    \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] , \in3[51] ,
    \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] , \in3[57] ,
    \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] ,
    \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] ,
    \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75] ,
    \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] , \in3[81] ,
    \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] , \in3[87] ,
    \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] , \in3[93] ,
    \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] , \in3[99] ,
    \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] , \in3[105] ,
    \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] , \in3[111] ,
    \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] ,
    \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] ,
    \in3[124] , \in3[125] , \in3[126] , \in3[127] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1]   );
  input  \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
    \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
    \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] ,
    \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] ,
    \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] ,
    \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] ,
    \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] ,
    \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] ,
    \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] ,
    \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] ,
    \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] ,
    \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] ,
    \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
    \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] ,
    \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] ,
    \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] ,
    \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] ,
    \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] ,
    \in0[108] , \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] ,
    \in0[114] , \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] ,
    \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] ,
    \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] ,
    \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] ,
    \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] ,
    \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] ,
    \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] ,
    \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] ,
    \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] ,
    \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] ,
    \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] ,
    \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
    \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] ,
    \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] ,
    \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] ,
    \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] ,
    \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] ,
    \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] ,
    \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] ,
    \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] ,
    \in1[107] , \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] ,
    \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] ,
    \in1[119] , \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] ,
    \in1[125] , \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] ,
    \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] ,
    \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] ,
    \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] ,
    \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] ,
    \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
    \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] ,
    \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] ,
    \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] ,
    \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] ,
    \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] ,
    \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] ,
    \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] ,
    \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] ,
    \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] ,
    \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] ,
    \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
    \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] ,
    \in2[106] , \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] ,
    \in2[112] , \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] ,
    \in2[118] , \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] ,
    \in2[124] , \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] ,
    \in3[2] , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
    \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
    \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] ,
    \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] ,
    \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] ,
    \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] ,
    \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] ,
    \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] ,
    \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] ,
    \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] ,
    \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] ,
    \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] ,
    \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
    \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] ,
    \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] ,
    \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] ,
    \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] ,
    \in3[105] , \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] ,
    \in3[111] , \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] ,
    \in3[117] , \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] ,
    \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1] ;
  wire new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_,
    new_n2721_, new_n2722_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2774_,
    new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_,
    new_n2781_, new_n2782_, new_n2784_, new_n2785_, new_n2787_, new_n2788_,
    new_n2790_, new_n2791_, new_n2793_, new_n2794_, new_n2796_, new_n2797_,
    new_n2799_, new_n2800_, new_n2802_, new_n2803_, new_n2805_, new_n2806_,
    new_n2807_, new_n2809_, new_n2810_, new_n2812_, new_n2813_, new_n2815_,
    new_n2816_, new_n2818_, new_n2819_, new_n2821_, new_n2822_, new_n2824_,
    new_n2825_, new_n2827_, new_n2828_, new_n2830_, new_n2831_, new_n2832_,
    new_n2834_, new_n2835_, new_n2837_, new_n2838_, new_n2840_, new_n2841_,
    new_n2843_, new_n2844_, new_n2846_, new_n2847_, new_n2849_, new_n2850_,
    new_n2852_, new_n2853_, new_n2855_, new_n2856_, new_n2858_, new_n2859_,
    new_n2860_, new_n2862_, new_n2863_, new_n2865_, new_n2866_, new_n2867_,
    new_n2869_, new_n2870_, new_n2872_, new_n2873_, new_n2875_, new_n2876_,
    new_n2878_, new_n2879_, new_n2881_, new_n2882_, new_n2884_, new_n2885_,
    new_n2887_, new_n2888_, new_n2889_, new_n2891_, new_n2892_, new_n2894_,
    new_n2895_, new_n2897_, new_n2898_, new_n2900_, new_n2901_, new_n2903_,
    new_n2904_, new_n2906_, new_n2907_, new_n2909_, new_n2910_, new_n2912_,
    new_n2913_, new_n2915_, new_n2916_, new_n2918_, new_n2919_, new_n2921_,
    new_n2922_, new_n2924_, new_n2925_, new_n2927_, new_n2928_, new_n2929_,
    new_n2931_, new_n2932_, new_n2934_, new_n2935_, new_n2937_, new_n2938_,
    new_n2939_, new_n2941_, new_n2942_, new_n2943_, new_n2945_, new_n2946_,
    new_n2948_, new_n2949_, new_n2951_, new_n2952_, new_n2954_, new_n2955_,
    new_n2957_, new_n2958_, new_n2960_, new_n2961_, new_n2963_, new_n2964_,
    new_n2966_, new_n2967_, new_n2969_, new_n2970_, new_n2972_, new_n2973_,
    new_n2975_, new_n2976_, new_n2978_, new_n2979_, new_n2981_, new_n2982_,
    new_n2984_, new_n2985_, new_n2987_, new_n2988_, new_n2990_, new_n2991_,
    new_n2993_, new_n2994_, new_n2996_, new_n2997_, new_n2999_, new_n3000_,
    new_n3002_, new_n3003_, new_n3005_, new_n3006_, new_n3008_, new_n3009_,
    new_n3011_, new_n3012_, new_n3014_, new_n3015_, new_n3016_, new_n3018_,
    new_n3019_, new_n3021_, new_n3022_, new_n3024_, new_n3025_, new_n3027_,
    new_n3028_, new_n3030_, new_n3031_, new_n3033_, new_n3034_, new_n3036_,
    new_n3037_, new_n3039_, new_n3040_, new_n3042_, new_n3043_, new_n3045_,
    new_n3046_, new_n3048_, new_n3049_, new_n3051_, new_n3052_, new_n3054_,
    new_n3055_, new_n3057_, new_n3058_, new_n3060_, new_n3061_, new_n3063_,
    new_n3064_, new_n3066_, new_n3067_, new_n3069_, new_n3070_, new_n3072_,
    new_n3073_, new_n3075_, new_n3076_, new_n3078_, new_n3079_, new_n3081_,
    new_n3082_, new_n3084_, new_n3085_, new_n3087_, new_n3088_, new_n3089_,
    new_n3091_, new_n3092_, new_n3094_, new_n3095_, new_n3097_, new_n3098_,
    new_n3100_, new_n3101_, new_n3103_, new_n3104_, new_n3106_, new_n3107_,
    new_n3109_, new_n3110_, new_n3112_, new_n3113_, new_n3115_, new_n3116_,
    new_n3118_, new_n3119_, new_n3121_, new_n3122_, new_n3124_, new_n3125_,
    new_n3127_, new_n3128_, new_n3130_, new_n3131_, new_n3133_, new_n3134_,
    new_n3135_, new_n3137_, new_n3138_, new_n3139_, new_n3141_, new_n3142_,
    new_n3144_, new_n3145_, new_n3147_, new_n3148_, new_n3150_, new_n3152_,
    new_n3153_;
  INV_X1     g0000(.I(\in3[0] ), .ZN(new_n643_));
  INV_X1     g0001(.I(\in3[127] ), .ZN(new_n644_));
  NOR2_X1    g0002(.A1(new_n644_), .A2(\in2[127] ), .ZN(new_n645_));
  INV_X1     g0003(.I(new_n645_), .ZN(new_n646_));
  INV_X1     g0004(.I(\in2[125] ), .ZN(new_n647_));
  INV_X1     g0005(.I(\in2[126] ), .ZN(new_n648_));
  AOI22_X1   g0006(.A1(new_n647_), .A2(\in3[125] ), .B1(new_n648_), .B2(\in3[126] ), .ZN(new_n649_));
  INV_X1     g0007(.I(new_n649_), .ZN(new_n650_));
  INV_X1     g0008(.I(\in3[124] ), .ZN(new_n651_));
  INV_X1     g0009(.I(\in3[125] ), .ZN(new_n652_));
  AOI22_X1   g0010(.A1(\in2[124] ), .A2(new_n651_), .B1(new_n652_), .B2(\in2[125] ), .ZN(new_n653_));
  NAND2_X1   g0011(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1     g0012(.I(\in3[126] ), .ZN(new_n655_));
  AOI22_X1   g0013(.A1(\in2[126] ), .A2(new_n655_), .B1(new_n644_), .B2(\in2[127] ), .ZN(new_n656_));
  AND2_X2    g0014(.A1(new_n654_), .A2(new_n656_), .Z(new_n657_));
  INV_X1     g0015(.I(new_n657_), .ZN(new_n658_));
  INV_X1     g0016(.I(\in2[47] ), .ZN(new_n659_));
  NAND2_X1   g0017(.A1(new_n659_), .A2(\in3[47] ), .ZN(new_n660_));
  INV_X1     g0018(.I(\in2[46] ), .ZN(new_n661_));
  NAND2_X1   g0019(.A1(new_n661_), .A2(\in3[46] ), .ZN(new_n662_));
  INV_X1     g0020(.I(\in2[45] ), .ZN(new_n663_));
  NAND2_X1   g0021(.A1(new_n663_), .A2(\in3[45] ), .ZN(new_n664_));
  INV_X1     g0022(.I(\in2[44] ), .ZN(new_n665_));
  NAND2_X1   g0023(.A1(new_n665_), .A2(\in3[44] ), .ZN(new_n666_));
  AOI22_X1   g0024(.A1(new_n660_), .A2(new_n662_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1     g0025(.I(\in2[43] ), .ZN(new_n668_));
  INV_X1     g0026(.I(\in2[42] ), .ZN(new_n669_));
  AOI22_X1   g0027(.A1(new_n669_), .A2(\in3[42] ), .B1(new_n668_), .B2(\in3[43] ), .ZN(new_n670_));
  INV_X1     g0028(.I(\in3[41] ), .ZN(new_n671_));
  INV_X1     g0029(.I(\in3[42] ), .ZN(new_n672_));
  AOI22_X1   g0030(.A1(\in2[41] ), .A2(new_n671_), .B1(new_n672_), .B2(\in2[42] ), .ZN(new_n673_));
  INV_X1     g0031(.I(\in2[41] ), .ZN(new_n674_));
  NOR4_X1    g0032(.A1(new_n674_), .A2(\in2[40] ), .A3(\in3[40] ), .A4(\in3[41] ), .ZN(new_n675_));
  NOR2_X1    g0033(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  OAI22_X1   g0034(.A1(new_n676_), .A2(new_n670_), .B1(new_n668_), .B2(\in3[43] ), .ZN(new_n677_));
  INV_X1     g0035(.I(\in3[47] ), .ZN(new_n678_));
  NOR2_X1    g0036(.A1(new_n678_), .A2(\in2[47] ), .ZN(new_n679_));
  INV_X1     g0037(.I(\in3[45] ), .ZN(new_n680_));
  NOR2_X1    g0038(.A1(new_n680_), .A2(\in2[45] ), .ZN(new_n681_));
  NOR3_X1    g0039(.A1(new_n679_), .A2(new_n681_), .A3(new_n662_), .ZN(new_n682_));
  NOR3_X1    g0040(.A1(new_n679_), .A2(new_n661_), .A3(\in3[46] ), .ZN(new_n683_));
  NOR3_X1    g0041(.A1(new_n681_), .A2(new_n665_), .A3(\in3[44] ), .ZN(new_n684_));
  NOR2_X1    g0042(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1   g0043(.A1(new_n685_), .A2(new_n682_), .ZN(new_n686_));
  AOI21_X1   g0044(.A1(new_n677_), .A2(new_n667_), .B(new_n686_), .ZN(new_n687_));
  INV_X1     g0045(.I(\in2[39] ), .ZN(new_n688_));
  NAND2_X1   g0046(.A1(new_n688_), .A2(\in3[39] ), .ZN(new_n689_));
  INV_X1     g0047(.I(\in2[38] ), .ZN(new_n690_));
  NAND2_X1   g0048(.A1(new_n690_), .A2(\in3[38] ), .ZN(new_n691_));
  INV_X1     g0049(.I(\in2[37] ), .ZN(new_n692_));
  NAND2_X1   g0050(.A1(new_n692_), .A2(\in3[37] ), .ZN(new_n693_));
  INV_X1     g0051(.I(\in2[36] ), .ZN(new_n694_));
  NAND2_X1   g0052(.A1(new_n694_), .A2(\in3[36] ), .ZN(new_n695_));
  AOI22_X1   g0053(.A1(new_n689_), .A2(new_n691_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1     g0054(.I(\in2[35] ), .ZN(new_n697_));
  NAND2_X1   g0055(.A1(new_n697_), .A2(\in3[35] ), .ZN(new_n698_));
  INV_X1     g0056(.I(\in2[34] ), .ZN(new_n699_));
  NAND2_X1   g0057(.A1(new_n699_), .A2(\in3[34] ), .ZN(new_n700_));
  INV_X1     g0058(.I(\in2[33] ), .ZN(new_n701_));
  OAI22_X1   g0059(.A1(new_n701_), .A2(\in3[33] ), .B1(new_n699_), .B2(\in3[34] ), .ZN(new_n702_));
  INV_X1     g0060(.I(\in2[32] ), .ZN(new_n703_));
  INV_X1     g0061(.I(\in3[32] ), .ZN(new_n704_));
  INV_X1     g0062(.I(\in3[33] ), .ZN(new_n705_));
  NAND4_X1   g0063(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .A4(\in2[33] ), .ZN(new_n706_));
  AOI22_X1   g0064(.A1(new_n702_), .A2(new_n706_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n707_));
  NOR2_X1    g0065(.A1(new_n697_), .A2(\in3[35] ), .ZN(new_n708_));
  OAI21_X1   g0066(.A1(new_n707_), .A2(new_n708_), .B(new_n696_), .ZN(new_n709_));
  INV_X1     g0067(.I(\in2[40] ), .ZN(new_n710_));
  AOI22_X1   g0068(.A1(new_n710_), .A2(\in3[40] ), .B1(new_n674_), .B2(\in3[41] ), .ZN(new_n711_));
  NOR2_X1    g0069(.A1(new_n670_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1   g0070(.A1(new_n712_), .A2(new_n667_), .ZN(new_n713_));
  INV_X1     g0071(.I(\in2[31] ), .ZN(new_n714_));
  NAND2_X1   g0072(.A1(new_n714_), .A2(\in3[31] ), .ZN(new_n715_));
  INV_X1     g0073(.I(\in3[39] ), .ZN(new_n716_));
  NOR2_X1    g0074(.A1(new_n716_), .A2(\in2[39] ), .ZN(new_n717_));
  INV_X1     g0075(.I(\in3[37] ), .ZN(new_n718_));
  NOR2_X1    g0076(.A1(new_n718_), .A2(\in2[37] ), .ZN(new_n719_));
  NOR2_X1    g0077(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  AND2_X2    g0078(.A1(new_n720_), .A2(new_n715_), .Z(new_n721_));
  NOR2_X1    g0079(.A1(new_n694_), .A2(\in3[36] ), .ZN(new_n722_));
  AOI21_X1   g0080(.A1(new_n690_), .A2(\in3[38] ), .B(new_n717_), .ZN(new_n723_));
  AOI21_X1   g0081(.A1(new_n693_), .A2(new_n722_), .B(new_n723_), .ZN(new_n724_));
  NAND4_X1   g0082(.A1(new_n709_), .A2(new_n713_), .A3(new_n721_), .A4(new_n724_), .ZN(new_n725_));
  INV_X1     g0083(.I(\in2[54] ), .ZN(new_n726_));
  INV_X1     g0084(.I(\in2[55] ), .ZN(new_n727_));
  AOI22_X1   g0085(.A1(new_n726_), .A2(\in3[54] ), .B1(new_n727_), .B2(\in3[55] ), .ZN(new_n728_));
  INV_X1     g0086(.I(\in2[53] ), .ZN(new_n729_));
  NAND2_X1   g0087(.A1(new_n729_), .A2(\in3[53] ), .ZN(new_n730_));
  INV_X1     g0088(.I(\in2[52] ), .ZN(new_n731_));
  NOR2_X1    g0089(.A1(new_n731_), .A2(\in3[52] ), .ZN(new_n732_));
  NAND3_X1   g0090(.A1(new_n728_), .A2(new_n730_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1     g0091(.I(\in3[51] ), .ZN(new_n734_));
  NOR2_X1    g0092(.A1(new_n734_), .A2(\in2[51] ), .ZN(new_n735_));
  INV_X1     g0093(.I(\in3[50] ), .ZN(new_n736_));
  NOR2_X1    g0094(.A1(new_n736_), .A2(\in2[50] ), .ZN(new_n737_));
  INV_X1     g0095(.I(\in3[49] ), .ZN(new_n738_));
  AOI22_X1   g0096(.A1(\in2[49] ), .A2(new_n738_), .B1(new_n736_), .B2(\in2[50] ), .ZN(new_n739_));
  INV_X1     g0097(.I(\in2[49] ), .ZN(new_n740_));
  NOR4_X1    g0098(.A1(new_n740_), .A2(\in2[48] ), .A3(\in3[48] ), .A4(\in3[49] ), .ZN(new_n741_));
  OAI22_X1   g0099(.A1(new_n739_), .A2(new_n741_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n742_));
  INV_X1     g0100(.I(\in2[51] ), .ZN(new_n743_));
  NOR2_X1    g0101(.A1(new_n743_), .A2(\in3[51] ), .ZN(new_n744_));
  INV_X1     g0102(.I(new_n744_), .ZN(new_n745_));
  AOI21_X1   g0103(.A1(new_n742_), .A2(new_n745_), .B(new_n733_), .ZN(new_n746_));
  INV_X1     g0104(.I(\in3[54] ), .ZN(new_n747_));
  INV_X1     g0105(.I(\in3[55] ), .ZN(new_n748_));
  OAI22_X1   g0106(.A1(\in2[54] ), .A2(new_n747_), .B1(new_n748_), .B2(\in2[55] ), .ZN(new_n749_));
  INV_X1     g0107(.I(\in3[53] ), .ZN(new_n750_));
  NOR2_X1    g0108(.A1(new_n750_), .A2(\in2[53] ), .ZN(new_n751_));
  INV_X1     g0109(.I(\in3[52] ), .ZN(new_n752_));
  NAND2_X1   g0110(.A1(new_n752_), .A2(\in2[52] ), .ZN(new_n753_));
  NOR3_X1    g0111(.A1(new_n749_), .A2(new_n751_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1     g0112(.I(\in2[50] ), .ZN(new_n755_));
  AOI22_X1   g0113(.A1(new_n755_), .A2(\in3[50] ), .B1(new_n743_), .B2(\in3[51] ), .ZN(new_n756_));
  INV_X1     g0114(.I(\in2[48] ), .ZN(new_n757_));
  AOI22_X1   g0115(.A1(new_n757_), .A2(\in3[48] ), .B1(new_n740_), .B2(\in3[49] ), .ZN(new_n758_));
  NOR2_X1    g0116(.A1(new_n727_), .A2(\in3[55] ), .ZN(new_n759_));
  NOR3_X1    g0117(.A1(new_n756_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1   g0118(.A1(new_n760_), .A2(new_n754_), .ZN(new_n761_));
  INV_X1     g0119(.I(\in3[63] ), .ZN(new_n762_));
  NOR2_X1    g0120(.A1(new_n762_), .A2(\in2[63] ), .ZN(new_n763_));
  INV_X1     g0121(.I(\in3[62] ), .ZN(new_n764_));
  NOR2_X1    g0122(.A1(new_n764_), .A2(\in2[62] ), .ZN(new_n765_));
  INV_X1     g0123(.I(\in3[61] ), .ZN(new_n766_));
  NOR2_X1    g0124(.A1(new_n766_), .A2(\in2[61] ), .ZN(new_n767_));
  INV_X1     g0125(.I(\in3[60] ), .ZN(new_n768_));
  NOR2_X1    g0126(.A1(new_n768_), .A2(\in2[60] ), .ZN(new_n769_));
  OAI22_X1   g0127(.A1(new_n763_), .A2(new_n765_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1     g0128(.I(\in3[56] ), .ZN(new_n771_));
  INV_X1     g0129(.I(\in3[57] ), .ZN(new_n772_));
  OAI22_X1   g0130(.A1(\in2[56] ), .A2(new_n771_), .B1(new_n772_), .B2(\in2[57] ), .ZN(new_n773_));
  INV_X1     g0131(.I(\in3[58] ), .ZN(new_n774_));
  INV_X1     g0132(.I(\in3[59] ), .ZN(new_n775_));
  OAI22_X1   g0133(.A1(\in2[58] ), .A2(new_n774_), .B1(new_n775_), .B2(\in2[59] ), .ZN(new_n776_));
  NAND2_X1   g0134(.A1(new_n773_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1   g0135(.A1(new_n747_), .A2(\in2[54] ), .ZN(new_n778_));
  NAND2_X1   g0136(.A1(new_n750_), .A2(\in2[53] ), .ZN(new_n779_));
  AOI22_X1   g0137(.A1(new_n730_), .A2(new_n732_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  OAI22_X1   g0138(.A1(new_n770_), .A2(new_n777_), .B1(new_n780_), .B2(new_n728_), .ZN(new_n781_));
  NOR3_X1    g0139(.A1(new_n781_), .A2(new_n746_), .A3(new_n761_), .ZN(new_n782_));
  OAI21_X1   g0140(.A1(new_n687_), .A2(new_n725_), .B(new_n782_), .ZN(new_n783_));
  INV_X1     g0141(.I(\in2[63] ), .ZN(new_n784_));
  NAND2_X1   g0142(.A1(new_n784_), .A2(\in3[63] ), .ZN(new_n785_));
  INV_X1     g0143(.I(\in2[62] ), .ZN(new_n786_));
  NAND2_X1   g0144(.A1(new_n786_), .A2(\in3[62] ), .ZN(new_n787_));
  INV_X1     g0145(.I(\in2[61] ), .ZN(new_n788_));
  NAND2_X1   g0146(.A1(new_n788_), .A2(\in3[61] ), .ZN(new_n789_));
  INV_X1     g0147(.I(\in2[60] ), .ZN(new_n790_));
  NAND2_X1   g0148(.A1(new_n790_), .A2(\in3[60] ), .ZN(new_n791_));
  AOI22_X1   g0149(.A1(new_n785_), .A2(new_n787_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1     g0150(.I(\in2[58] ), .ZN(new_n793_));
  INV_X1     g0151(.I(\in2[59] ), .ZN(new_n794_));
  AOI22_X1   g0152(.A1(new_n793_), .A2(\in3[58] ), .B1(new_n794_), .B2(\in3[59] ), .ZN(new_n795_));
  INV_X1     g0153(.I(\in2[57] ), .ZN(new_n796_));
  OAI22_X1   g0154(.A1(new_n796_), .A2(\in3[57] ), .B1(new_n793_), .B2(\in3[58] ), .ZN(new_n797_));
  INV_X1     g0155(.I(\in2[56] ), .ZN(new_n798_));
  NAND4_X1   g0156(.A1(new_n798_), .A2(new_n771_), .A3(new_n772_), .A4(\in2[57] ), .ZN(new_n799_));
  AOI21_X1   g0157(.A1(new_n797_), .A2(new_n799_), .B(new_n795_), .ZN(new_n800_));
  NOR2_X1    g0158(.A1(new_n794_), .A2(\in3[59] ), .ZN(new_n801_));
  OAI21_X1   g0159(.A1(new_n800_), .A2(new_n801_), .B(new_n792_), .ZN(new_n802_));
  INV_X1     g0160(.I(\in3[65] ), .ZN(new_n803_));
  NOR2_X1    g0161(.A1(new_n803_), .A2(\in2[65] ), .ZN(new_n804_));
  NOR2_X1    g0162(.A1(new_n804_), .A2(\in3[64] ), .ZN(new_n805_));
  NAND2_X1   g0163(.A1(new_n803_), .A2(\in2[65] ), .ZN(new_n806_));
  INV_X1     g0164(.I(\in3[66] ), .ZN(new_n807_));
  AOI21_X1   g0165(.A1(new_n807_), .A2(\in2[66] ), .B(\in2[64] ), .ZN(new_n808_));
  NAND2_X1   g0166(.A1(new_n808_), .A2(new_n806_), .ZN(new_n809_));
  INV_X1     g0167(.I(\in3[67] ), .ZN(new_n810_));
  OAI22_X1   g0168(.A1(\in2[66] ), .A2(new_n807_), .B1(new_n810_), .B2(\in2[67] ), .ZN(new_n811_));
  OAI21_X1   g0169(.A1(new_n809_), .A2(new_n805_), .B(new_n811_), .ZN(new_n812_));
  NOR3_X1    g0170(.A1(new_n767_), .A2(new_n790_), .A3(\in3[60] ), .ZN(new_n813_));
  AOI21_X1   g0171(.A1(new_n786_), .A2(\in3[62] ), .B(new_n763_), .ZN(new_n814_));
  INV_X1     g0172(.I(\in2[64] ), .ZN(new_n815_));
  NOR4_X1    g0173(.A1(new_n811_), .A2(new_n815_), .A3(\in3[64] ), .A4(new_n804_), .ZN(new_n816_));
  NAND2_X1   g0174(.A1(new_n810_), .A2(\in2[67] ), .ZN(new_n817_));
  NAND3_X1   g0175(.A1(new_n785_), .A2(new_n789_), .A3(new_n817_), .ZN(new_n818_));
  NOR4_X1    g0176(.A1(new_n816_), .A2(new_n813_), .A3(new_n814_), .A4(new_n818_), .ZN(new_n819_));
  NAND3_X1   g0177(.A1(new_n819_), .A2(new_n802_), .A3(new_n812_), .ZN(new_n820_));
  INV_X1     g0178(.I(new_n820_), .ZN(new_n821_));
  INV_X1     g0179(.I(\in3[70] ), .ZN(new_n822_));
  INV_X1     g0180(.I(\in3[71] ), .ZN(new_n823_));
  OAI22_X1   g0181(.A1(\in2[70] ), .A2(new_n822_), .B1(new_n823_), .B2(\in2[71] ), .ZN(new_n824_));
  INV_X1     g0182(.I(new_n824_), .ZN(new_n825_));
  INV_X1     g0183(.I(\in2[71] ), .ZN(new_n826_));
  AOI22_X1   g0184(.A1(\in2[70] ), .A2(new_n822_), .B1(new_n826_), .B2(\in3[71] ), .ZN(new_n827_));
  INV_X1     g0185(.I(\in2[69] ), .ZN(new_n828_));
  INV_X1     g0186(.I(\in3[68] ), .ZN(new_n829_));
  AOI22_X1   g0187(.A1(\in2[68] ), .A2(new_n829_), .B1(new_n828_), .B2(\in3[69] ), .ZN(new_n830_));
  AOI21_X1   g0188(.A1(new_n824_), .A2(new_n830_), .B(new_n827_), .ZN(new_n831_));
  INV_X1     g0189(.I(\in2[72] ), .ZN(new_n832_));
  INV_X1     g0190(.I(\in3[74] ), .ZN(new_n833_));
  INV_X1     g0191(.I(\in3[75] ), .ZN(new_n834_));
  OAI22_X1   g0192(.A1(\in2[74] ), .A2(new_n833_), .B1(new_n834_), .B2(\in2[75] ), .ZN(new_n835_));
  INV_X1     g0193(.I(\in3[73] ), .ZN(new_n836_));
  NOR2_X1    g0194(.A1(new_n836_), .A2(\in2[73] ), .ZN(new_n837_));
  NOR4_X1    g0195(.A1(new_n835_), .A2(new_n832_), .A3(\in3[72] ), .A4(new_n837_), .ZN(new_n838_));
  INV_X1     g0196(.I(\in3[69] ), .ZN(new_n839_));
  OAI22_X1   g0197(.A1(\in2[68] ), .A2(new_n829_), .B1(new_n839_), .B2(\in2[69] ), .ZN(new_n840_));
  INV_X1     g0198(.I(new_n840_), .ZN(new_n841_));
  NOR4_X1    g0199(.A1(new_n831_), .A2(new_n838_), .A3(new_n825_), .A4(new_n841_), .ZN(new_n842_));
  INV_X1     g0200(.I(new_n842_), .ZN(new_n843_));
  AOI21_X1   g0201(.A1(new_n783_), .A2(new_n821_), .B(new_n843_), .ZN(new_n844_));
  NOR2_X1    g0202(.A1(new_n837_), .A2(\in3[72] ), .ZN(new_n845_));
  INV_X1     g0203(.I(\in2[73] ), .ZN(new_n846_));
  AOI21_X1   g0204(.A1(new_n833_), .A2(\in2[74] ), .B(\in2[72] ), .ZN(new_n847_));
  OAI21_X1   g0205(.A1(new_n846_), .A2(\in3[73] ), .B(new_n847_), .ZN(new_n848_));
  OR2_X2     g0206(.A1(new_n848_), .A2(new_n845_), .Z(new_n849_));
  AOI22_X1   g0207(.A1(new_n849_), .A2(new_n835_), .B1(\in2[75] ), .B2(new_n834_), .ZN(new_n850_));
  INV_X1     g0208(.I(\in2[79] ), .ZN(new_n851_));
  INV_X1     g0209(.I(\in3[78] ), .ZN(new_n852_));
  AOI22_X1   g0210(.A1(\in2[78] ), .A2(new_n852_), .B1(new_n851_), .B2(\in3[79] ), .ZN(new_n853_));
  INV_X1     g0211(.I(\in3[79] ), .ZN(new_n854_));
  OAI22_X1   g0212(.A1(\in2[78] ), .A2(new_n852_), .B1(new_n854_), .B2(\in2[79] ), .ZN(new_n855_));
  INV_X1     g0213(.I(\in3[76] ), .ZN(new_n856_));
  INV_X1     g0214(.I(\in3[77] ), .ZN(new_n857_));
  NOR2_X1    g0215(.A1(new_n857_), .A2(\in2[77] ), .ZN(new_n858_));
  AOI21_X1   g0216(.A1(\in2[76] ), .A2(new_n856_), .B(new_n858_), .ZN(new_n859_));
  AOI21_X1   g0217(.A1(new_n859_), .A2(new_n855_), .B(new_n853_), .ZN(new_n860_));
  NOR2_X1    g0218(.A1(new_n856_), .A2(\in2[76] ), .ZN(new_n861_));
  OAI21_X1   g0219(.A1(new_n858_), .A2(new_n861_), .B(new_n855_), .ZN(new_n862_));
  INV_X1     g0220(.I(new_n862_), .ZN(new_n863_));
  NOR3_X1    g0221(.A1(new_n850_), .A2(new_n860_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1     g0222(.I(new_n864_), .ZN(new_n865_));
  INV_X1     g0223(.I(\in3[81] ), .ZN(new_n866_));
  NOR2_X1    g0224(.A1(new_n866_), .A2(\in2[81] ), .ZN(new_n867_));
  NOR2_X1    g0225(.A1(new_n867_), .A2(\in3[80] ), .ZN(new_n868_));
  NAND2_X1   g0226(.A1(new_n866_), .A2(\in2[81] ), .ZN(new_n869_));
  INV_X1     g0227(.I(\in3[82] ), .ZN(new_n870_));
  AOI21_X1   g0228(.A1(new_n870_), .A2(\in2[82] ), .B(\in2[80] ), .ZN(new_n871_));
  NAND2_X1   g0229(.A1(new_n871_), .A2(new_n869_), .ZN(new_n872_));
  INV_X1     g0230(.I(\in3[83] ), .ZN(new_n873_));
  OAI22_X1   g0231(.A1(\in2[82] ), .A2(new_n870_), .B1(new_n873_), .B2(\in2[83] ), .ZN(new_n874_));
  OAI21_X1   g0232(.A1(new_n872_), .A2(new_n868_), .B(new_n874_), .ZN(new_n875_));
  INV_X1     g0233(.I(\in3[86] ), .ZN(new_n876_));
  INV_X1     g0234(.I(\in3[87] ), .ZN(new_n877_));
  OAI22_X1   g0235(.A1(\in2[86] ), .A2(new_n876_), .B1(new_n877_), .B2(\in2[87] ), .ZN(new_n878_));
  INV_X1     g0236(.I(\in3[85] ), .ZN(new_n879_));
  NOR2_X1    g0237(.A1(new_n879_), .A2(\in2[85] ), .ZN(new_n880_));
  INV_X1     g0238(.I(\in3[84] ), .ZN(new_n881_));
  NOR2_X1    g0239(.A1(new_n881_), .A2(\in2[84] ), .ZN(new_n882_));
  OAI21_X1   g0240(.A1(new_n880_), .A2(new_n882_), .B(new_n878_), .ZN(new_n883_));
  INV_X1     g0241(.I(\in2[83] ), .ZN(new_n884_));
  NOR2_X1    g0242(.A1(new_n884_), .A2(\in3[83] ), .ZN(new_n885_));
  INV_X1     g0243(.I(\in3[80] ), .ZN(new_n886_));
  NAND2_X1   g0244(.A1(new_n886_), .A2(\in2[80] ), .ZN(new_n887_));
  NOR4_X1    g0245(.A1(new_n874_), .A2(new_n867_), .A3(new_n885_), .A4(new_n887_), .ZN(new_n888_));
  NAND3_X1   g0246(.A1(new_n875_), .A2(new_n883_), .A3(new_n888_), .ZN(new_n889_));
  INV_X1     g0247(.I(new_n889_), .ZN(new_n890_));
  OAI21_X1   g0248(.A1(new_n844_), .A2(new_n865_), .B(new_n890_), .ZN(new_n891_));
  INV_X1     g0249(.I(\in3[89] ), .ZN(new_n892_));
  NOR2_X1    g0250(.A1(new_n892_), .A2(\in2[89] ), .ZN(new_n893_));
  NOR2_X1    g0251(.A1(new_n893_), .A2(\in3[88] ), .ZN(new_n894_));
  INV_X1     g0252(.I(new_n894_), .ZN(new_n895_));
  INV_X1     g0253(.I(\in3[90] ), .ZN(new_n896_));
  AOI21_X1   g0254(.A1(new_n896_), .A2(\in2[90] ), .B(\in2[88] ), .ZN(new_n897_));
  INV_X1     g0255(.I(new_n897_), .ZN(new_n898_));
  AOI21_X1   g0256(.A1(\in2[89] ), .A2(new_n892_), .B(new_n898_), .ZN(new_n899_));
  INV_X1     g0257(.I(\in3[91] ), .ZN(new_n900_));
  OAI22_X1   g0258(.A1(\in2[90] ), .A2(new_n896_), .B1(new_n900_), .B2(\in2[91] ), .ZN(new_n901_));
  INV_X1     g0259(.I(new_n901_), .ZN(new_n902_));
  AOI21_X1   g0260(.A1(new_n899_), .A2(new_n895_), .B(new_n902_), .ZN(new_n903_));
  INV_X1     g0261(.I(new_n880_), .ZN(new_n904_));
  NAND2_X1   g0262(.A1(new_n881_), .A2(\in2[84] ), .ZN(new_n905_));
  AND3_X2    g0263(.A1(new_n904_), .A2(new_n878_), .A3(new_n905_), .Z(new_n906_));
  INV_X1     g0264(.I(\in2[87] ), .ZN(new_n907_));
  AOI22_X1   g0265(.A1(\in2[86] ), .A2(new_n876_), .B1(new_n907_), .B2(\in3[87] ), .ZN(new_n908_));
  INV_X1     g0266(.I(\in2[88] ), .ZN(new_n909_));
  NOR3_X1    g0267(.A1(new_n893_), .A2(new_n909_), .A3(\in3[88] ), .ZN(new_n910_));
  AOI22_X1   g0268(.A1(new_n902_), .A2(new_n910_), .B1(\in2[91] ), .B2(new_n900_), .ZN(new_n911_));
  INV_X1     g0269(.I(new_n911_), .ZN(new_n912_));
  NOR4_X1    g0270(.A1(new_n912_), .A2(new_n903_), .A3(new_n906_), .A4(new_n908_), .ZN(new_n913_));
  INV_X1     g0271(.I(\in3[94] ), .ZN(new_n914_));
  INV_X1     g0272(.I(\in3[95] ), .ZN(new_n915_));
  OAI22_X1   g0273(.A1(\in2[94] ), .A2(new_n914_), .B1(new_n915_), .B2(\in2[95] ), .ZN(new_n916_));
  INV_X1     g0274(.I(new_n916_), .ZN(new_n917_));
  INV_X1     g0275(.I(\in2[95] ), .ZN(new_n918_));
  AOI22_X1   g0276(.A1(\in2[94] ), .A2(new_n914_), .B1(new_n918_), .B2(\in3[95] ), .ZN(new_n919_));
  INV_X1     g0277(.I(\in2[93] ), .ZN(new_n920_));
  INV_X1     g0278(.I(\in3[92] ), .ZN(new_n921_));
  AOI22_X1   g0279(.A1(\in2[92] ), .A2(new_n921_), .B1(new_n920_), .B2(\in3[93] ), .ZN(new_n922_));
  AOI21_X1   g0280(.A1(new_n916_), .A2(new_n922_), .B(new_n919_), .ZN(new_n923_));
  INV_X1     g0281(.I(\in2[96] ), .ZN(new_n924_));
  INV_X1     g0282(.I(\in2[98] ), .ZN(new_n925_));
  INV_X1     g0283(.I(\in2[99] ), .ZN(new_n926_));
  AOI22_X1   g0284(.A1(new_n925_), .A2(\in3[98] ), .B1(new_n926_), .B2(\in3[99] ), .ZN(new_n927_));
  INV_X1     g0285(.I(new_n927_), .ZN(new_n928_));
  INV_X1     g0286(.I(\in3[97] ), .ZN(new_n929_));
  NOR2_X1    g0287(.A1(new_n929_), .A2(\in2[97] ), .ZN(new_n930_));
  NOR4_X1    g0288(.A1(new_n928_), .A2(new_n924_), .A3(\in3[96] ), .A4(new_n930_), .ZN(new_n931_));
  INV_X1     g0289(.I(\in3[93] ), .ZN(new_n932_));
  OAI22_X1   g0290(.A1(\in2[92] ), .A2(new_n921_), .B1(new_n932_), .B2(\in2[93] ), .ZN(new_n933_));
  INV_X1     g0291(.I(new_n933_), .ZN(new_n934_));
  NOR4_X1    g0292(.A1(new_n931_), .A2(new_n917_), .A3(new_n923_), .A4(new_n934_), .ZN(new_n935_));
  INV_X1     g0293(.I(new_n935_), .ZN(new_n936_));
  AOI21_X1   g0294(.A1(new_n891_), .A2(new_n913_), .B(new_n936_), .ZN(new_n937_));
  NOR2_X1    g0295(.A1(new_n930_), .A2(\in3[96] ), .ZN(new_n938_));
  NAND2_X1   g0296(.A1(new_n929_), .A2(\in2[97] ), .ZN(new_n939_));
  INV_X1     g0297(.I(new_n939_), .ZN(new_n940_));
  NOR2_X1    g0298(.A1(new_n925_), .A2(\in3[98] ), .ZN(new_n941_));
  NOR4_X1    g0299(.A1(new_n938_), .A2(new_n940_), .A3(\in2[96] ), .A4(new_n941_), .ZN(new_n942_));
  OAI22_X1   g0300(.A1(new_n942_), .A2(new_n927_), .B1(new_n926_), .B2(\in3[99] ), .ZN(new_n943_));
  INV_X1     g0301(.I(new_n943_), .ZN(new_n944_));
  INV_X1     g0302(.I(\in2[103] ), .ZN(new_n945_));
  INV_X1     g0303(.I(\in3[102] ), .ZN(new_n946_));
  AOI22_X1   g0304(.A1(\in2[102] ), .A2(new_n946_), .B1(new_n945_), .B2(\in3[103] ), .ZN(new_n947_));
  INV_X1     g0305(.I(\in3[103] ), .ZN(new_n948_));
  OAI22_X1   g0306(.A1(\in2[102] ), .A2(new_n946_), .B1(new_n948_), .B2(\in2[103] ), .ZN(new_n949_));
  INV_X1     g0307(.I(\in3[100] ), .ZN(new_n950_));
  INV_X1     g0308(.I(\in3[101] ), .ZN(new_n951_));
  NOR2_X1    g0309(.A1(new_n951_), .A2(\in2[101] ), .ZN(new_n952_));
  AOI21_X1   g0310(.A1(\in2[100] ), .A2(new_n950_), .B(new_n952_), .ZN(new_n953_));
  AOI21_X1   g0311(.A1(new_n953_), .A2(new_n949_), .B(new_n947_), .ZN(new_n954_));
  NOR2_X1    g0312(.A1(new_n950_), .A2(\in2[100] ), .ZN(new_n955_));
  OAI21_X1   g0313(.A1(new_n952_), .A2(new_n955_), .B(new_n949_), .ZN(new_n956_));
  INV_X1     g0314(.I(new_n956_), .ZN(new_n957_));
  NOR3_X1    g0315(.A1(new_n944_), .A2(new_n954_), .A3(new_n957_), .ZN(new_n958_));
  INV_X1     g0316(.I(new_n958_), .ZN(new_n959_));
  INV_X1     g0317(.I(\in3[105] ), .ZN(new_n960_));
  NOR2_X1    g0318(.A1(new_n960_), .A2(\in2[105] ), .ZN(new_n961_));
  NOR2_X1    g0319(.A1(new_n961_), .A2(\in3[104] ), .ZN(new_n962_));
  NAND2_X1   g0320(.A1(new_n960_), .A2(\in2[105] ), .ZN(new_n963_));
  INV_X1     g0321(.I(\in3[106] ), .ZN(new_n964_));
  AOI21_X1   g0322(.A1(new_n964_), .A2(\in2[106] ), .B(\in2[104] ), .ZN(new_n965_));
  NAND2_X1   g0323(.A1(new_n965_), .A2(new_n963_), .ZN(new_n966_));
  INV_X1     g0324(.I(\in3[107] ), .ZN(new_n967_));
  OAI22_X1   g0325(.A1(\in2[106] ), .A2(new_n964_), .B1(new_n967_), .B2(\in2[107] ), .ZN(new_n968_));
  OAI21_X1   g0326(.A1(new_n966_), .A2(new_n962_), .B(new_n968_), .ZN(new_n969_));
  INV_X1     g0327(.I(\in2[110] ), .ZN(new_n970_));
  INV_X1     g0328(.I(\in2[111] ), .ZN(new_n971_));
  AOI22_X1   g0329(.A1(new_n970_), .A2(\in3[110] ), .B1(new_n971_), .B2(\in3[111] ), .ZN(new_n972_));
  INV_X1     g0330(.I(new_n972_), .ZN(new_n973_));
  INV_X1     g0331(.I(\in3[109] ), .ZN(new_n974_));
  NOR2_X1    g0332(.A1(new_n974_), .A2(\in2[109] ), .ZN(new_n975_));
  INV_X1     g0333(.I(\in3[108] ), .ZN(new_n976_));
  NOR2_X1    g0334(.A1(new_n976_), .A2(\in2[108] ), .ZN(new_n977_));
  OAI21_X1   g0335(.A1(new_n975_), .A2(new_n977_), .B(new_n973_), .ZN(new_n978_));
  INV_X1     g0336(.I(\in2[107] ), .ZN(new_n979_));
  NOR2_X1    g0337(.A1(new_n979_), .A2(\in3[107] ), .ZN(new_n980_));
  INV_X1     g0338(.I(\in3[104] ), .ZN(new_n981_));
  NAND2_X1   g0339(.A1(new_n981_), .A2(\in2[104] ), .ZN(new_n982_));
  NOR4_X1    g0340(.A1(new_n968_), .A2(new_n961_), .A3(new_n980_), .A4(new_n982_), .ZN(new_n983_));
  NAND3_X1   g0341(.A1(new_n978_), .A2(new_n969_), .A3(new_n983_), .ZN(new_n984_));
  INV_X1     g0342(.I(new_n984_), .ZN(new_n985_));
  OAI21_X1   g0343(.A1(new_n937_), .A2(new_n959_), .B(new_n985_), .ZN(new_n986_));
  INV_X1     g0344(.I(\in3[113] ), .ZN(new_n987_));
  NOR2_X1    g0345(.A1(new_n987_), .A2(\in2[113] ), .ZN(new_n988_));
  NOR2_X1    g0346(.A1(new_n988_), .A2(\in3[112] ), .ZN(new_n989_));
  INV_X1     g0347(.I(new_n989_), .ZN(new_n990_));
  INV_X1     g0348(.I(\in3[114] ), .ZN(new_n991_));
  AOI21_X1   g0349(.A1(new_n991_), .A2(\in2[114] ), .B(\in2[112] ), .ZN(new_n992_));
  INV_X1     g0350(.I(new_n992_), .ZN(new_n993_));
  AOI21_X1   g0351(.A1(\in2[113] ), .A2(new_n987_), .B(new_n993_), .ZN(new_n994_));
  INV_X1     g0352(.I(\in3[115] ), .ZN(new_n995_));
  OAI22_X1   g0353(.A1(\in2[114] ), .A2(new_n991_), .B1(new_n995_), .B2(\in2[115] ), .ZN(new_n996_));
  INV_X1     g0354(.I(new_n996_), .ZN(new_n997_));
  AOI21_X1   g0355(.A1(new_n994_), .A2(new_n990_), .B(new_n997_), .ZN(new_n998_));
  NAND2_X1   g0356(.A1(new_n976_), .A2(\in2[108] ), .ZN(new_n999_));
  INV_X1     g0357(.I(new_n999_), .ZN(new_n1000_));
  NOR3_X1    g0358(.A1(new_n1000_), .A2(new_n972_), .A3(new_n975_), .ZN(new_n1001_));
  INV_X1     g0359(.I(\in3[110] ), .ZN(new_n1002_));
  AOI22_X1   g0360(.A1(\in2[110] ), .A2(new_n1002_), .B1(new_n971_), .B2(\in3[111] ), .ZN(new_n1003_));
  INV_X1     g0361(.I(\in2[112] ), .ZN(new_n1004_));
  NOR3_X1    g0362(.A1(new_n988_), .A2(new_n1004_), .A3(\in3[112] ), .ZN(new_n1005_));
  AOI22_X1   g0363(.A1(new_n997_), .A2(new_n1005_), .B1(\in2[115] ), .B2(new_n995_), .ZN(new_n1006_));
  INV_X1     g0364(.I(new_n1006_), .ZN(new_n1007_));
  NOR4_X1    g0365(.A1(new_n1007_), .A2(new_n998_), .A3(new_n1001_), .A4(new_n1003_), .ZN(new_n1008_));
  INV_X1     g0366(.I(\in3[118] ), .ZN(new_n1009_));
  INV_X1     g0367(.I(\in3[119] ), .ZN(new_n1010_));
  OAI22_X1   g0368(.A1(\in2[118] ), .A2(new_n1009_), .B1(new_n1010_), .B2(\in2[119] ), .ZN(new_n1011_));
  INV_X1     g0369(.I(new_n1011_), .ZN(new_n1012_));
  INV_X1     g0370(.I(\in2[119] ), .ZN(new_n1013_));
  AOI22_X1   g0371(.A1(\in2[118] ), .A2(new_n1009_), .B1(new_n1013_), .B2(\in3[119] ), .ZN(new_n1014_));
  INV_X1     g0372(.I(\in2[117] ), .ZN(new_n1015_));
  INV_X1     g0373(.I(\in3[116] ), .ZN(new_n1016_));
  AOI22_X1   g0374(.A1(\in2[116] ), .A2(new_n1016_), .B1(new_n1015_), .B2(\in3[117] ), .ZN(new_n1017_));
  AOI21_X1   g0375(.A1(new_n1011_), .A2(new_n1017_), .B(new_n1014_), .ZN(new_n1018_));
  INV_X1     g0376(.I(\in2[120] ), .ZN(new_n1019_));
  INV_X1     g0377(.I(\in2[122] ), .ZN(new_n1020_));
  INV_X1     g0378(.I(\in2[123] ), .ZN(new_n1021_));
  AOI22_X1   g0379(.A1(new_n1020_), .A2(\in3[122] ), .B1(new_n1021_), .B2(\in3[123] ), .ZN(new_n1022_));
  INV_X1     g0380(.I(new_n1022_), .ZN(new_n1023_));
  INV_X1     g0381(.I(\in3[121] ), .ZN(new_n1024_));
  NOR2_X1    g0382(.A1(new_n1024_), .A2(\in2[121] ), .ZN(new_n1025_));
  NOR4_X1    g0383(.A1(new_n1023_), .A2(new_n1019_), .A3(\in3[120] ), .A4(new_n1025_), .ZN(new_n1026_));
  INV_X1     g0384(.I(\in3[117] ), .ZN(new_n1027_));
  OAI22_X1   g0385(.A1(\in2[116] ), .A2(new_n1016_), .B1(new_n1027_), .B2(\in2[117] ), .ZN(new_n1028_));
  INV_X1     g0386(.I(new_n1028_), .ZN(new_n1029_));
  NOR4_X1    g0387(.A1(new_n1026_), .A2(new_n1012_), .A3(new_n1018_), .A4(new_n1029_), .ZN(new_n1030_));
  INV_X1     g0388(.I(new_n1030_), .ZN(new_n1031_));
  AOI21_X1   g0389(.A1(new_n986_), .A2(new_n1008_), .B(new_n1031_), .ZN(new_n1032_));
  INV_X1     g0390(.I(\in2[127] ), .ZN(new_n1033_));
  OAI22_X1   g0391(.A1(\in2[124] ), .A2(new_n651_), .B1(new_n1033_), .B2(\in3[127] ), .ZN(new_n1034_));
  INV_X1     g0392(.I(new_n1034_), .ZN(new_n1035_));
  NOR2_X1    g0393(.A1(new_n1021_), .A2(\in3[123] ), .ZN(new_n1036_));
  NOR2_X1    g0394(.A1(new_n1025_), .A2(\in3[120] ), .ZN(new_n1037_));
  INV_X1     g0395(.I(new_n1037_), .ZN(new_n1038_));
  NOR2_X1    g0396(.A1(new_n1020_), .A2(\in3[122] ), .ZN(new_n1039_));
  NOR2_X1    g0397(.A1(new_n1039_), .A2(\in2[120] ), .ZN(new_n1040_));
  INV_X1     g0398(.I(new_n1040_), .ZN(new_n1041_));
  AOI21_X1   g0399(.A1(\in2[121] ), .A2(new_n1024_), .B(new_n1041_), .ZN(new_n1042_));
  AOI21_X1   g0400(.A1(new_n1042_), .A2(new_n1038_), .B(new_n1022_), .ZN(new_n1043_));
  OAI22_X1   g0401(.A1(new_n1043_), .A2(new_n1036_), .B1(new_n649_), .B2(new_n1035_), .ZN(new_n1044_));
  OAI21_X1   g0402(.A1(new_n1032_), .A2(new_n1044_), .B(new_n658_), .ZN(new_n1045_));
  NAND2_X1   g0403(.A1(new_n1045_), .A2(new_n646_), .ZN(new_n1046_));
  MUX2_X1    g0404(.I0(\in2[0] ), .I1(new_n643_), .S(new_n1046_), .Z(new_n1047_));
  INV_X1     g0405(.I(\in0[127] ), .ZN(new_n1048_));
  INV_X1     g0406(.I(\in1[127] ), .ZN(new_n1049_));
  INV_X1     g0407(.I(\in0[125] ), .ZN(new_n1050_));
  INV_X1     g0408(.I(\in0[126] ), .ZN(new_n1051_));
  AOI22_X1   g0409(.A1(new_n1050_), .A2(\in1[125] ), .B1(new_n1051_), .B2(\in1[126] ), .ZN(new_n1052_));
  INV_X1     g0410(.I(new_n1052_), .ZN(new_n1053_));
  INV_X1     g0411(.I(\in1[124] ), .ZN(new_n1054_));
  INV_X1     g0412(.I(\in1[125] ), .ZN(new_n1055_));
  AOI22_X1   g0413(.A1(\in0[124] ), .A2(new_n1054_), .B1(new_n1055_), .B2(\in0[125] ), .ZN(new_n1056_));
  NAND2_X1   g0414(.A1(new_n1053_), .A2(new_n1056_), .ZN(new_n1057_));
  INV_X1     g0415(.I(\in1[126] ), .ZN(new_n1058_));
  AOI22_X1   g0416(.A1(\in0[126] ), .A2(new_n1058_), .B1(new_n1049_), .B2(\in0[127] ), .ZN(new_n1059_));
  AND2_X2    g0417(.A1(new_n1057_), .A2(new_n1059_), .Z(new_n1060_));
  INV_X1     g0418(.I(new_n1060_), .ZN(new_n1061_));
  INV_X1     g0419(.I(\in0[47] ), .ZN(new_n1062_));
  NAND2_X1   g0420(.A1(new_n1062_), .A2(\in1[47] ), .ZN(new_n1063_));
  INV_X1     g0421(.I(\in0[46] ), .ZN(new_n1064_));
  NAND2_X1   g0422(.A1(new_n1064_), .A2(\in1[46] ), .ZN(new_n1065_));
  NAND2_X1   g0423(.A1(new_n1063_), .A2(new_n1065_), .ZN(new_n1066_));
  INV_X1     g0424(.I(\in0[45] ), .ZN(new_n1067_));
  NAND2_X1   g0425(.A1(new_n1067_), .A2(\in1[45] ), .ZN(new_n1068_));
  INV_X1     g0426(.I(\in0[44] ), .ZN(new_n1069_));
  NAND2_X1   g0427(.A1(new_n1069_), .A2(\in1[44] ), .ZN(new_n1070_));
  NAND2_X1   g0428(.A1(new_n1068_), .A2(new_n1070_), .ZN(new_n1071_));
  NAND2_X1   g0429(.A1(new_n1066_), .A2(new_n1071_), .ZN(new_n1072_));
  INV_X1     g0430(.I(\in1[43] ), .ZN(new_n1073_));
  INV_X1     g0431(.I(\in1[42] ), .ZN(new_n1074_));
  OAI22_X1   g0432(.A1(\in0[42] ), .A2(new_n1074_), .B1(new_n1073_), .B2(\in0[43] ), .ZN(new_n1075_));
  INV_X1     g0433(.I(\in0[41] ), .ZN(new_n1076_));
  INV_X1     g0434(.I(\in0[42] ), .ZN(new_n1077_));
  OAI22_X1   g0435(.A1(new_n1076_), .A2(\in1[41] ), .B1(new_n1077_), .B2(\in1[42] ), .ZN(new_n1078_));
  INV_X1     g0436(.I(\in0[40] ), .ZN(new_n1079_));
  INV_X1     g0437(.I(\in1[40] ), .ZN(new_n1080_));
  INV_X1     g0438(.I(\in1[41] ), .ZN(new_n1081_));
  NAND4_X1   g0439(.A1(new_n1079_), .A2(new_n1080_), .A3(new_n1081_), .A4(\in0[41] ), .ZN(new_n1082_));
  NAND2_X1   g0440(.A1(new_n1078_), .A2(new_n1082_), .ZN(new_n1083_));
  AOI22_X1   g0441(.A1(new_n1083_), .A2(new_n1075_), .B1(\in0[43] ), .B2(new_n1073_), .ZN(new_n1084_));
  NAND4_X1   g0442(.A1(new_n1063_), .A2(new_n1068_), .A3(new_n1064_), .A4(\in1[46] ), .ZN(new_n1085_));
  INV_X1     g0443(.I(\in1[47] ), .ZN(new_n1086_));
  NOR2_X1    g0444(.A1(new_n1086_), .A2(\in0[47] ), .ZN(new_n1087_));
  NOR3_X1    g0445(.A1(new_n1087_), .A2(new_n1064_), .A3(\in1[46] ), .ZN(new_n1088_));
  INV_X1     g0446(.I(\in1[45] ), .ZN(new_n1089_));
  NOR2_X1    g0447(.A1(new_n1089_), .A2(\in0[45] ), .ZN(new_n1090_));
  NOR3_X1    g0448(.A1(new_n1090_), .A2(new_n1069_), .A3(\in1[44] ), .ZN(new_n1091_));
  NOR3_X1    g0449(.A1(new_n1085_), .A2(new_n1088_), .A3(new_n1091_), .ZN(new_n1092_));
  OAI21_X1   g0450(.A1(new_n1084_), .A2(new_n1072_), .B(new_n1092_), .ZN(new_n1093_));
  INV_X1     g0451(.I(new_n1093_), .ZN(new_n1094_));
  INV_X1     g0452(.I(\in0[39] ), .ZN(new_n1095_));
  NAND2_X1   g0453(.A1(new_n1095_), .A2(\in1[39] ), .ZN(new_n1096_));
  INV_X1     g0454(.I(\in0[38] ), .ZN(new_n1097_));
  NAND2_X1   g0455(.A1(new_n1097_), .A2(\in1[38] ), .ZN(new_n1098_));
  INV_X1     g0456(.I(\in0[37] ), .ZN(new_n1099_));
  NAND2_X1   g0457(.A1(new_n1099_), .A2(\in1[37] ), .ZN(new_n1100_));
  INV_X1     g0458(.I(\in0[36] ), .ZN(new_n1101_));
  NAND2_X1   g0459(.A1(new_n1101_), .A2(\in1[36] ), .ZN(new_n1102_));
  AOI22_X1   g0460(.A1(new_n1096_), .A2(new_n1098_), .B1(new_n1100_), .B2(new_n1102_), .ZN(new_n1103_));
  INV_X1     g0461(.I(\in0[35] ), .ZN(new_n1104_));
  NAND2_X1   g0462(.A1(new_n1104_), .A2(\in1[35] ), .ZN(new_n1105_));
  INV_X1     g0463(.I(\in0[34] ), .ZN(new_n1106_));
  NAND2_X1   g0464(.A1(new_n1106_), .A2(\in1[34] ), .ZN(new_n1107_));
  INV_X1     g0465(.I(\in0[33] ), .ZN(new_n1108_));
  OAI22_X1   g0466(.A1(new_n1108_), .A2(\in1[33] ), .B1(new_n1106_), .B2(\in1[34] ), .ZN(new_n1109_));
  INV_X1     g0467(.I(\in0[32] ), .ZN(new_n1110_));
  INV_X1     g0468(.I(\in1[32] ), .ZN(new_n1111_));
  INV_X1     g0469(.I(\in1[33] ), .ZN(new_n1112_));
  NAND4_X1   g0470(.A1(new_n1110_), .A2(new_n1111_), .A3(new_n1112_), .A4(\in0[33] ), .ZN(new_n1113_));
  AOI22_X1   g0471(.A1(new_n1109_), .A2(new_n1113_), .B1(new_n1105_), .B2(new_n1107_), .ZN(new_n1114_));
  NOR2_X1    g0472(.A1(new_n1104_), .A2(\in1[35] ), .ZN(new_n1115_));
  OAI21_X1   g0473(.A1(new_n1114_), .A2(new_n1115_), .B(new_n1103_), .ZN(new_n1116_));
  OAI22_X1   g0474(.A1(\in0[40] ), .A2(new_n1080_), .B1(new_n1081_), .B2(\in0[41] ), .ZN(new_n1117_));
  NAND4_X1   g0475(.A1(new_n1066_), .A2(new_n1071_), .A3(new_n1075_), .A4(new_n1117_), .ZN(new_n1118_));
  INV_X1     g0476(.I(\in1[39] ), .ZN(new_n1119_));
  NOR2_X1    g0477(.A1(new_n1119_), .A2(\in0[39] ), .ZN(new_n1120_));
  INV_X1     g0478(.I(\in1[37] ), .ZN(new_n1121_));
  NOR2_X1    g0479(.A1(new_n1121_), .A2(\in0[37] ), .ZN(new_n1122_));
  INV_X1     g0480(.I(\in1[31] ), .ZN(new_n1123_));
  NOR2_X1    g0481(.A1(new_n1123_), .A2(\in0[31] ), .ZN(new_n1124_));
  NOR3_X1    g0482(.A1(new_n1120_), .A2(new_n1122_), .A3(new_n1124_), .ZN(new_n1125_));
  NOR3_X1    g0483(.A1(new_n1122_), .A2(new_n1101_), .A3(\in1[36] ), .ZN(new_n1126_));
  AOI21_X1   g0484(.A1(new_n1097_), .A2(\in1[38] ), .B(new_n1120_), .ZN(new_n1127_));
  NOR2_X1    g0485(.A1(new_n1127_), .A2(new_n1126_), .ZN(new_n1128_));
  NAND4_X1   g0486(.A1(new_n1116_), .A2(new_n1118_), .A3(new_n1125_), .A4(new_n1128_), .ZN(new_n1129_));
  INV_X1     g0487(.I(\in0[54] ), .ZN(new_n1130_));
  INV_X1     g0488(.I(\in0[55] ), .ZN(new_n1131_));
  AOI22_X1   g0489(.A1(new_n1130_), .A2(\in1[54] ), .B1(new_n1131_), .B2(\in1[55] ), .ZN(new_n1132_));
  INV_X1     g0490(.I(\in0[53] ), .ZN(new_n1133_));
  NAND2_X1   g0491(.A1(new_n1133_), .A2(\in1[53] ), .ZN(new_n1134_));
  INV_X1     g0492(.I(\in0[52] ), .ZN(new_n1135_));
  NOR2_X1    g0493(.A1(new_n1135_), .A2(\in1[52] ), .ZN(new_n1136_));
  NAND3_X1   g0494(.A1(new_n1132_), .A2(new_n1134_), .A3(new_n1136_), .ZN(new_n1137_));
  INV_X1     g0495(.I(\in1[50] ), .ZN(new_n1138_));
  INV_X1     g0496(.I(\in1[51] ), .ZN(new_n1139_));
  OAI22_X1   g0497(.A1(\in0[50] ), .A2(new_n1138_), .B1(new_n1139_), .B2(\in0[51] ), .ZN(new_n1140_));
  INV_X1     g0498(.I(\in1[49] ), .ZN(new_n1141_));
  AOI22_X1   g0499(.A1(\in0[49] ), .A2(new_n1141_), .B1(new_n1138_), .B2(\in0[50] ), .ZN(new_n1142_));
  INV_X1     g0500(.I(\in0[49] ), .ZN(new_n1143_));
  NOR4_X1    g0501(.A1(new_n1143_), .A2(\in0[48] ), .A3(\in1[48] ), .A4(\in1[49] ), .ZN(new_n1144_));
  OAI21_X1   g0502(.A1(new_n1142_), .A2(new_n1144_), .B(new_n1140_), .ZN(new_n1145_));
  INV_X1     g0503(.I(\in0[51] ), .ZN(new_n1146_));
  NOR2_X1    g0504(.A1(new_n1146_), .A2(\in1[51] ), .ZN(new_n1147_));
  INV_X1     g0505(.I(new_n1147_), .ZN(new_n1148_));
  AOI21_X1   g0506(.A1(new_n1145_), .A2(new_n1148_), .B(new_n1137_), .ZN(new_n1149_));
  INV_X1     g0507(.I(\in1[54] ), .ZN(new_n1150_));
  INV_X1     g0508(.I(\in1[55] ), .ZN(new_n1151_));
  OAI22_X1   g0509(.A1(\in0[54] ), .A2(new_n1150_), .B1(new_n1151_), .B2(\in0[55] ), .ZN(new_n1152_));
  INV_X1     g0510(.I(\in1[53] ), .ZN(new_n1153_));
  NOR2_X1    g0511(.A1(new_n1153_), .A2(\in0[53] ), .ZN(new_n1154_));
  INV_X1     g0512(.I(\in1[52] ), .ZN(new_n1155_));
  NAND2_X1   g0513(.A1(new_n1155_), .A2(\in0[52] ), .ZN(new_n1156_));
  NOR3_X1    g0514(.A1(new_n1152_), .A2(new_n1154_), .A3(new_n1156_), .ZN(new_n1157_));
  INV_X1     g0515(.I(\in0[50] ), .ZN(new_n1158_));
  AOI22_X1   g0516(.A1(new_n1158_), .A2(\in1[50] ), .B1(new_n1146_), .B2(\in1[51] ), .ZN(new_n1159_));
  INV_X1     g0517(.I(\in0[48] ), .ZN(new_n1160_));
  AOI22_X1   g0518(.A1(new_n1160_), .A2(\in1[48] ), .B1(new_n1143_), .B2(\in1[49] ), .ZN(new_n1161_));
  NOR2_X1    g0519(.A1(new_n1131_), .A2(\in1[55] ), .ZN(new_n1162_));
  NOR3_X1    g0520(.A1(new_n1159_), .A2(new_n1161_), .A3(new_n1162_), .ZN(new_n1163_));
  NAND2_X1   g0521(.A1(new_n1163_), .A2(new_n1157_), .ZN(new_n1164_));
  INV_X1     g0522(.I(\in0[63] ), .ZN(new_n1165_));
  NAND2_X1   g0523(.A1(new_n1165_), .A2(\in1[63] ), .ZN(new_n1166_));
  INV_X1     g0524(.I(\in0[62] ), .ZN(new_n1167_));
  NAND2_X1   g0525(.A1(new_n1167_), .A2(\in1[62] ), .ZN(new_n1168_));
  NAND2_X1   g0526(.A1(new_n1166_), .A2(new_n1168_), .ZN(new_n1169_));
  INV_X1     g0527(.I(\in0[61] ), .ZN(new_n1170_));
  NAND2_X1   g0528(.A1(new_n1170_), .A2(\in1[61] ), .ZN(new_n1171_));
  INV_X1     g0529(.I(\in0[60] ), .ZN(new_n1172_));
  NAND2_X1   g0530(.A1(new_n1172_), .A2(\in1[60] ), .ZN(new_n1173_));
  NAND2_X1   g0531(.A1(new_n1171_), .A2(new_n1173_), .ZN(new_n1174_));
  NAND2_X1   g0532(.A1(new_n1169_), .A2(new_n1174_), .ZN(new_n1175_));
  INV_X1     g0533(.I(\in1[56] ), .ZN(new_n1176_));
  INV_X1     g0534(.I(\in1[57] ), .ZN(new_n1177_));
  OAI22_X1   g0535(.A1(\in0[56] ), .A2(new_n1176_), .B1(new_n1177_), .B2(\in0[57] ), .ZN(new_n1178_));
  INV_X1     g0536(.I(\in1[58] ), .ZN(new_n1179_));
  INV_X1     g0537(.I(\in1[59] ), .ZN(new_n1180_));
  OAI22_X1   g0538(.A1(\in0[58] ), .A2(new_n1179_), .B1(new_n1180_), .B2(\in0[59] ), .ZN(new_n1181_));
  NAND2_X1   g0539(.A1(new_n1178_), .A2(new_n1181_), .ZN(new_n1182_));
  NAND2_X1   g0540(.A1(new_n1150_), .A2(\in0[54] ), .ZN(new_n1183_));
  NAND2_X1   g0541(.A1(new_n1153_), .A2(\in0[53] ), .ZN(new_n1184_));
  AOI22_X1   g0542(.A1(new_n1134_), .A2(new_n1136_), .B1(new_n1183_), .B2(new_n1184_), .ZN(new_n1185_));
  OAI22_X1   g0543(.A1(new_n1175_), .A2(new_n1182_), .B1(new_n1185_), .B2(new_n1132_), .ZN(new_n1186_));
  NOR3_X1    g0544(.A1(new_n1186_), .A2(new_n1149_), .A3(new_n1164_), .ZN(new_n1187_));
  OAI21_X1   g0545(.A1(new_n1094_), .A2(new_n1129_), .B(new_n1187_), .ZN(new_n1188_));
  AOI22_X1   g0546(.A1(new_n1166_), .A2(new_n1168_), .B1(new_n1171_), .B2(new_n1173_), .ZN(new_n1189_));
  INV_X1     g0547(.I(\in0[59] ), .ZN(new_n1190_));
  AOI22_X1   g0548(.A1(\in0[57] ), .A2(new_n1177_), .B1(new_n1179_), .B2(\in0[58] ), .ZN(new_n1191_));
  INV_X1     g0549(.I(\in0[57] ), .ZN(new_n1192_));
  NOR4_X1    g0550(.A1(new_n1192_), .A2(\in0[56] ), .A3(\in1[56] ), .A4(\in1[57] ), .ZN(new_n1193_));
  OAI21_X1   g0551(.A1(new_n1191_), .A2(new_n1193_), .B(new_n1181_), .ZN(new_n1194_));
  OAI21_X1   g0552(.A1(new_n1190_), .A2(\in1[59] ), .B(new_n1194_), .ZN(new_n1195_));
  INV_X1     g0553(.I(\in1[64] ), .ZN(new_n1196_));
  INV_X1     g0554(.I(\in0[65] ), .ZN(new_n1197_));
  NAND2_X1   g0555(.A1(new_n1197_), .A2(\in1[65] ), .ZN(new_n1198_));
  NAND2_X1   g0556(.A1(new_n1198_), .A2(new_n1196_), .ZN(new_n1199_));
  NOR2_X1    g0557(.A1(new_n1197_), .A2(\in1[65] ), .ZN(new_n1200_));
  INV_X1     g0558(.I(\in0[66] ), .ZN(new_n1201_));
  NOR2_X1    g0559(.A1(new_n1201_), .A2(\in1[66] ), .ZN(new_n1202_));
  NOR3_X1    g0560(.A1(new_n1200_), .A2(new_n1202_), .A3(\in0[64] ), .ZN(new_n1203_));
  NAND2_X1   g0561(.A1(new_n1203_), .A2(new_n1199_), .ZN(new_n1204_));
  INV_X1     g0562(.I(\in1[66] ), .ZN(new_n1205_));
  INV_X1     g0563(.I(\in1[67] ), .ZN(new_n1206_));
  OAI22_X1   g0564(.A1(\in0[66] ), .A2(new_n1205_), .B1(new_n1206_), .B2(\in0[67] ), .ZN(new_n1207_));
  NAND2_X1   g0565(.A1(new_n1204_), .A2(new_n1207_), .ZN(new_n1208_));
  INV_X1     g0566(.I(\in1[61] ), .ZN(new_n1209_));
  NOR2_X1    g0567(.A1(new_n1209_), .A2(\in0[61] ), .ZN(new_n1210_));
  NOR3_X1    g0568(.A1(new_n1210_), .A2(new_n1172_), .A3(\in1[60] ), .ZN(new_n1211_));
  INV_X1     g0569(.I(\in1[63] ), .ZN(new_n1212_));
  NOR2_X1    g0570(.A1(new_n1212_), .A2(\in0[63] ), .ZN(new_n1213_));
  AOI21_X1   g0571(.A1(new_n1167_), .A2(\in1[62] ), .B(new_n1213_), .ZN(new_n1214_));
  NAND3_X1   g0572(.A1(new_n1198_), .A2(\in0[64] ), .A3(new_n1196_), .ZN(new_n1215_));
  NOR2_X1    g0573(.A1(new_n1215_), .A2(new_n1207_), .ZN(new_n1216_));
  NAND2_X1   g0574(.A1(new_n1206_), .A2(\in0[67] ), .ZN(new_n1217_));
  NAND3_X1   g0575(.A1(new_n1166_), .A2(new_n1171_), .A3(new_n1217_), .ZN(new_n1218_));
  NOR4_X1    g0576(.A1(new_n1216_), .A2(new_n1218_), .A3(new_n1211_), .A4(new_n1214_), .ZN(new_n1219_));
  NAND2_X1   g0577(.A1(new_n1219_), .A2(new_n1208_), .ZN(new_n1220_));
  AOI21_X1   g0578(.A1(new_n1189_), .A2(new_n1195_), .B(new_n1220_), .ZN(new_n1221_));
  INV_X1     g0579(.I(\in1[70] ), .ZN(new_n1222_));
  INV_X1     g0580(.I(\in1[71] ), .ZN(new_n1223_));
  OAI22_X1   g0581(.A1(\in0[70] ), .A2(new_n1222_), .B1(new_n1223_), .B2(\in0[71] ), .ZN(new_n1224_));
  INV_X1     g0582(.I(new_n1224_), .ZN(new_n1225_));
  INV_X1     g0583(.I(\in0[71] ), .ZN(new_n1226_));
  AOI22_X1   g0584(.A1(\in0[70] ), .A2(new_n1222_), .B1(new_n1226_), .B2(\in1[71] ), .ZN(new_n1227_));
  INV_X1     g0585(.I(\in0[69] ), .ZN(new_n1228_));
  INV_X1     g0586(.I(\in1[68] ), .ZN(new_n1229_));
  AOI22_X1   g0587(.A1(\in0[68] ), .A2(new_n1229_), .B1(new_n1228_), .B2(\in1[69] ), .ZN(new_n1230_));
  AOI21_X1   g0588(.A1(new_n1224_), .A2(new_n1230_), .B(new_n1227_), .ZN(new_n1231_));
  INV_X1     g0589(.I(\in0[72] ), .ZN(new_n1232_));
  INV_X1     g0590(.I(\in1[74] ), .ZN(new_n1233_));
  INV_X1     g0591(.I(\in1[75] ), .ZN(new_n1234_));
  OAI22_X1   g0592(.A1(\in0[74] ), .A2(new_n1233_), .B1(new_n1234_), .B2(\in0[75] ), .ZN(new_n1235_));
  INV_X1     g0593(.I(\in1[73] ), .ZN(new_n1236_));
  NOR2_X1    g0594(.A1(new_n1236_), .A2(\in0[73] ), .ZN(new_n1237_));
  NOR4_X1    g0595(.A1(new_n1235_), .A2(new_n1232_), .A3(\in1[72] ), .A4(new_n1237_), .ZN(new_n1238_));
  INV_X1     g0596(.I(\in1[69] ), .ZN(new_n1239_));
  OAI22_X1   g0597(.A1(\in0[68] ), .A2(new_n1229_), .B1(new_n1239_), .B2(\in0[69] ), .ZN(new_n1240_));
  INV_X1     g0598(.I(new_n1240_), .ZN(new_n1241_));
  NOR4_X1    g0599(.A1(new_n1231_), .A2(new_n1238_), .A3(new_n1225_), .A4(new_n1241_), .ZN(new_n1242_));
  INV_X1     g0600(.I(new_n1242_), .ZN(new_n1243_));
  AOI21_X1   g0601(.A1(new_n1188_), .A2(new_n1221_), .B(new_n1243_), .ZN(new_n1244_));
  INV_X1     g0602(.I(\in1[72] ), .ZN(new_n1245_));
  OAI21_X1   g0603(.A1(\in0[73] ), .A2(new_n1236_), .B(new_n1245_), .ZN(new_n1246_));
  NAND2_X1   g0604(.A1(new_n1236_), .A2(\in0[73] ), .ZN(new_n1247_));
  AOI21_X1   g0605(.A1(new_n1233_), .A2(\in0[74] ), .B(\in0[72] ), .ZN(new_n1248_));
  NAND3_X1   g0606(.A1(new_n1246_), .A2(new_n1248_), .A3(new_n1247_), .ZN(new_n1249_));
  AOI22_X1   g0607(.A1(new_n1249_), .A2(new_n1235_), .B1(\in0[75] ), .B2(new_n1234_), .ZN(new_n1250_));
  INV_X1     g0608(.I(\in0[79] ), .ZN(new_n1251_));
  INV_X1     g0609(.I(\in1[78] ), .ZN(new_n1252_));
  AOI22_X1   g0610(.A1(\in0[78] ), .A2(new_n1252_), .B1(new_n1251_), .B2(\in1[79] ), .ZN(new_n1253_));
  INV_X1     g0611(.I(\in1[79] ), .ZN(new_n1254_));
  OAI22_X1   g0612(.A1(\in0[78] ), .A2(new_n1252_), .B1(new_n1254_), .B2(\in0[79] ), .ZN(new_n1255_));
  INV_X1     g0613(.I(\in1[76] ), .ZN(new_n1256_));
  INV_X1     g0614(.I(\in1[77] ), .ZN(new_n1257_));
  NOR2_X1    g0615(.A1(new_n1257_), .A2(\in0[77] ), .ZN(new_n1258_));
  AOI21_X1   g0616(.A1(\in0[76] ), .A2(new_n1256_), .B(new_n1258_), .ZN(new_n1259_));
  AOI21_X1   g0617(.A1(new_n1259_), .A2(new_n1255_), .B(new_n1253_), .ZN(new_n1260_));
  NOR2_X1    g0618(.A1(new_n1256_), .A2(\in0[76] ), .ZN(new_n1261_));
  OAI21_X1   g0619(.A1(new_n1258_), .A2(new_n1261_), .B(new_n1255_), .ZN(new_n1262_));
  INV_X1     g0620(.I(new_n1262_), .ZN(new_n1263_));
  NOR3_X1    g0621(.A1(new_n1250_), .A2(new_n1263_), .A3(new_n1260_), .ZN(new_n1264_));
  INV_X1     g0622(.I(new_n1264_), .ZN(new_n1265_));
  INV_X1     g0623(.I(\in1[81] ), .ZN(new_n1266_));
  NOR2_X1    g0624(.A1(new_n1266_), .A2(\in0[81] ), .ZN(new_n1267_));
  NOR2_X1    g0625(.A1(new_n1267_), .A2(\in1[80] ), .ZN(new_n1268_));
  NAND2_X1   g0626(.A1(new_n1266_), .A2(\in0[81] ), .ZN(new_n1269_));
  INV_X1     g0627(.I(\in1[82] ), .ZN(new_n1270_));
  AOI21_X1   g0628(.A1(new_n1270_), .A2(\in0[82] ), .B(\in0[80] ), .ZN(new_n1271_));
  NAND2_X1   g0629(.A1(new_n1271_), .A2(new_n1269_), .ZN(new_n1272_));
  INV_X1     g0630(.I(\in1[83] ), .ZN(new_n1273_));
  OAI22_X1   g0631(.A1(\in0[82] ), .A2(new_n1270_), .B1(new_n1273_), .B2(\in0[83] ), .ZN(new_n1274_));
  OAI21_X1   g0632(.A1(new_n1272_), .A2(new_n1268_), .B(new_n1274_), .ZN(new_n1275_));
  INV_X1     g0633(.I(\in0[86] ), .ZN(new_n1276_));
  INV_X1     g0634(.I(\in0[87] ), .ZN(new_n1277_));
  AOI22_X1   g0635(.A1(new_n1276_), .A2(\in1[86] ), .B1(new_n1277_), .B2(\in1[87] ), .ZN(new_n1278_));
  INV_X1     g0636(.I(new_n1278_), .ZN(new_n1279_));
  INV_X1     g0637(.I(\in1[85] ), .ZN(new_n1280_));
  NOR2_X1    g0638(.A1(new_n1280_), .A2(\in0[85] ), .ZN(new_n1281_));
  INV_X1     g0639(.I(\in1[84] ), .ZN(new_n1282_));
  NOR2_X1    g0640(.A1(new_n1282_), .A2(\in0[84] ), .ZN(new_n1283_));
  OAI21_X1   g0641(.A1(new_n1281_), .A2(new_n1283_), .B(new_n1279_), .ZN(new_n1284_));
  INV_X1     g0642(.I(\in0[83] ), .ZN(new_n1285_));
  NOR2_X1    g0643(.A1(new_n1285_), .A2(\in1[83] ), .ZN(new_n1286_));
  INV_X1     g0644(.I(\in1[80] ), .ZN(new_n1287_));
  NAND2_X1   g0645(.A1(new_n1287_), .A2(\in0[80] ), .ZN(new_n1288_));
  NOR4_X1    g0646(.A1(new_n1274_), .A2(new_n1267_), .A3(new_n1286_), .A4(new_n1288_), .ZN(new_n1289_));
  NAND3_X1   g0647(.A1(new_n1284_), .A2(new_n1275_), .A3(new_n1289_), .ZN(new_n1290_));
  INV_X1     g0648(.I(new_n1290_), .ZN(new_n1291_));
  OAI21_X1   g0649(.A1(new_n1244_), .A2(new_n1265_), .B(new_n1291_), .ZN(new_n1292_));
  INV_X1     g0650(.I(\in1[89] ), .ZN(new_n1293_));
  NOR2_X1    g0651(.A1(new_n1293_), .A2(\in0[89] ), .ZN(new_n1294_));
  NOR2_X1    g0652(.A1(new_n1294_), .A2(\in1[88] ), .ZN(new_n1295_));
  INV_X1     g0653(.I(new_n1295_), .ZN(new_n1296_));
  INV_X1     g0654(.I(\in1[90] ), .ZN(new_n1297_));
  AOI21_X1   g0655(.A1(new_n1297_), .A2(\in0[90] ), .B(\in0[88] ), .ZN(new_n1298_));
  INV_X1     g0656(.I(new_n1298_), .ZN(new_n1299_));
  AOI21_X1   g0657(.A1(\in0[89] ), .A2(new_n1293_), .B(new_n1299_), .ZN(new_n1300_));
  INV_X1     g0658(.I(\in1[91] ), .ZN(new_n1301_));
  OAI22_X1   g0659(.A1(\in0[90] ), .A2(new_n1297_), .B1(new_n1301_), .B2(\in0[91] ), .ZN(new_n1302_));
  INV_X1     g0660(.I(new_n1302_), .ZN(new_n1303_));
  AOI21_X1   g0661(.A1(new_n1300_), .A2(new_n1296_), .B(new_n1303_), .ZN(new_n1304_));
  NAND2_X1   g0662(.A1(new_n1282_), .A2(\in0[84] ), .ZN(new_n1305_));
  INV_X1     g0663(.I(new_n1305_), .ZN(new_n1306_));
  NOR3_X1    g0664(.A1(new_n1306_), .A2(new_n1278_), .A3(new_n1281_), .ZN(new_n1307_));
  INV_X1     g0665(.I(\in1[86] ), .ZN(new_n1308_));
  AOI22_X1   g0666(.A1(\in0[86] ), .A2(new_n1308_), .B1(new_n1277_), .B2(\in1[87] ), .ZN(new_n1309_));
  INV_X1     g0667(.I(\in1[88] ), .ZN(new_n1310_));
  NAND2_X1   g0668(.A1(new_n1310_), .A2(\in0[88] ), .ZN(new_n1311_));
  NOR2_X1    g0669(.A1(new_n1294_), .A2(new_n1311_), .ZN(new_n1312_));
  AOI22_X1   g0670(.A1(new_n1303_), .A2(new_n1312_), .B1(\in0[91] ), .B2(new_n1301_), .ZN(new_n1313_));
  INV_X1     g0671(.I(new_n1313_), .ZN(new_n1314_));
  NOR4_X1    g0672(.A1(new_n1314_), .A2(new_n1304_), .A3(new_n1307_), .A4(new_n1309_), .ZN(new_n1315_));
  INV_X1     g0673(.I(\in1[94] ), .ZN(new_n1316_));
  INV_X1     g0674(.I(\in1[95] ), .ZN(new_n1317_));
  OAI22_X1   g0675(.A1(\in0[94] ), .A2(new_n1316_), .B1(new_n1317_), .B2(\in0[95] ), .ZN(new_n1318_));
  INV_X1     g0676(.I(new_n1318_), .ZN(new_n1319_));
  INV_X1     g0677(.I(\in0[95] ), .ZN(new_n1320_));
  AOI22_X1   g0678(.A1(\in0[94] ), .A2(new_n1316_), .B1(new_n1320_), .B2(\in1[95] ), .ZN(new_n1321_));
  INV_X1     g0679(.I(\in0[93] ), .ZN(new_n1322_));
  INV_X1     g0680(.I(\in1[92] ), .ZN(new_n1323_));
  AOI22_X1   g0681(.A1(\in0[92] ), .A2(new_n1323_), .B1(new_n1322_), .B2(\in1[93] ), .ZN(new_n1324_));
  AOI21_X1   g0682(.A1(new_n1318_), .A2(new_n1324_), .B(new_n1321_), .ZN(new_n1325_));
  INV_X1     g0683(.I(\in0[96] ), .ZN(new_n1326_));
  INV_X1     g0684(.I(\in0[98] ), .ZN(new_n1327_));
  INV_X1     g0685(.I(\in0[99] ), .ZN(new_n1328_));
  AOI22_X1   g0686(.A1(new_n1327_), .A2(\in1[98] ), .B1(new_n1328_), .B2(\in1[99] ), .ZN(new_n1329_));
  INV_X1     g0687(.I(new_n1329_), .ZN(new_n1330_));
  INV_X1     g0688(.I(\in1[97] ), .ZN(new_n1331_));
  NOR2_X1    g0689(.A1(new_n1331_), .A2(\in0[97] ), .ZN(new_n1332_));
  NOR4_X1    g0690(.A1(new_n1330_), .A2(new_n1326_), .A3(\in1[96] ), .A4(new_n1332_), .ZN(new_n1333_));
  INV_X1     g0691(.I(\in1[93] ), .ZN(new_n1334_));
  OAI22_X1   g0692(.A1(\in0[92] ), .A2(new_n1323_), .B1(new_n1334_), .B2(\in0[93] ), .ZN(new_n1335_));
  INV_X1     g0693(.I(new_n1335_), .ZN(new_n1336_));
  NOR4_X1    g0694(.A1(new_n1333_), .A2(new_n1319_), .A3(new_n1325_), .A4(new_n1336_), .ZN(new_n1337_));
  INV_X1     g0695(.I(new_n1337_), .ZN(new_n1338_));
  AOI21_X1   g0696(.A1(new_n1292_), .A2(new_n1315_), .B(new_n1338_), .ZN(new_n1339_));
  NOR2_X1    g0697(.A1(new_n1332_), .A2(\in1[96] ), .ZN(new_n1340_));
  NAND2_X1   g0698(.A1(new_n1331_), .A2(\in0[97] ), .ZN(new_n1341_));
  INV_X1     g0699(.I(new_n1341_), .ZN(new_n1342_));
  NOR2_X1    g0700(.A1(new_n1327_), .A2(\in1[98] ), .ZN(new_n1343_));
  NOR4_X1    g0701(.A1(new_n1340_), .A2(new_n1342_), .A3(\in0[96] ), .A4(new_n1343_), .ZN(new_n1344_));
  OAI22_X1   g0702(.A1(new_n1344_), .A2(new_n1329_), .B1(new_n1328_), .B2(\in1[99] ), .ZN(new_n1345_));
  INV_X1     g0703(.I(new_n1345_), .ZN(new_n1346_));
  INV_X1     g0704(.I(\in0[103] ), .ZN(new_n1347_));
  INV_X1     g0705(.I(\in1[102] ), .ZN(new_n1348_));
  AOI22_X1   g0706(.A1(\in0[102] ), .A2(new_n1348_), .B1(new_n1347_), .B2(\in1[103] ), .ZN(new_n1349_));
  INV_X1     g0707(.I(\in1[103] ), .ZN(new_n1350_));
  OAI22_X1   g0708(.A1(\in0[102] ), .A2(new_n1348_), .B1(new_n1350_), .B2(\in0[103] ), .ZN(new_n1351_));
  INV_X1     g0709(.I(\in1[100] ), .ZN(new_n1352_));
  INV_X1     g0710(.I(\in1[101] ), .ZN(new_n1353_));
  NOR2_X1    g0711(.A1(new_n1353_), .A2(\in0[101] ), .ZN(new_n1354_));
  AOI21_X1   g0712(.A1(\in0[100] ), .A2(new_n1352_), .B(new_n1354_), .ZN(new_n1355_));
  AOI21_X1   g0713(.A1(new_n1355_), .A2(new_n1351_), .B(new_n1349_), .ZN(new_n1356_));
  NOR2_X1    g0714(.A1(new_n1352_), .A2(\in0[100] ), .ZN(new_n1357_));
  OAI21_X1   g0715(.A1(new_n1354_), .A2(new_n1357_), .B(new_n1351_), .ZN(new_n1358_));
  INV_X1     g0716(.I(new_n1358_), .ZN(new_n1359_));
  NOR3_X1    g0717(.A1(new_n1346_), .A2(new_n1356_), .A3(new_n1359_), .ZN(new_n1360_));
  INV_X1     g0718(.I(new_n1360_), .ZN(new_n1361_));
  INV_X1     g0719(.I(\in1[105] ), .ZN(new_n1362_));
  NOR2_X1    g0720(.A1(new_n1362_), .A2(\in0[105] ), .ZN(new_n1363_));
  NOR2_X1    g0721(.A1(new_n1363_), .A2(\in1[104] ), .ZN(new_n1364_));
  NAND2_X1   g0722(.A1(new_n1362_), .A2(\in0[105] ), .ZN(new_n1365_));
  INV_X1     g0723(.I(\in1[106] ), .ZN(new_n1366_));
  AOI21_X1   g0724(.A1(new_n1366_), .A2(\in0[106] ), .B(\in0[104] ), .ZN(new_n1367_));
  NAND2_X1   g0725(.A1(new_n1367_), .A2(new_n1365_), .ZN(new_n1368_));
  INV_X1     g0726(.I(\in1[107] ), .ZN(new_n1369_));
  OAI22_X1   g0727(.A1(\in0[106] ), .A2(new_n1366_), .B1(new_n1369_), .B2(\in0[107] ), .ZN(new_n1370_));
  OAI21_X1   g0728(.A1(new_n1368_), .A2(new_n1364_), .B(new_n1370_), .ZN(new_n1371_));
  INV_X1     g0729(.I(\in0[110] ), .ZN(new_n1372_));
  INV_X1     g0730(.I(\in0[111] ), .ZN(new_n1373_));
  AOI22_X1   g0731(.A1(new_n1372_), .A2(\in1[110] ), .B1(new_n1373_), .B2(\in1[111] ), .ZN(new_n1374_));
  INV_X1     g0732(.I(new_n1374_), .ZN(new_n1375_));
  INV_X1     g0733(.I(\in1[109] ), .ZN(new_n1376_));
  NOR2_X1    g0734(.A1(new_n1376_), .A2(\in0[109] ), .ZN(new_n1377_));
  INV_X1     g0735(.I(\in1[108] ), .ZN(new_n1378_));
  NOR2_X1    g0736(.A1(new_n1378_), .A2(\in0[108] ), .ZN(new_n1379_));
  OAI21_X1   g0737(.A1(new_n1377_), .A2(new_n1379_), .B(new_n1375_), .ZN(new_n1380_));
  INV_X1     g0738(.I(\in0[107] ), .ZN(new_n1381_));
  NOR2_X1    g0739(.A1(new_n1381_), .A2(\in1[107] ), .ZN(new_n1382_));
  INV_X1     g0740(.I(\in1[104] ), .ZN(new_n1383_));
  NAND2_X1   g0741(.A1(new_n1383_), .A2(\in0[104] ), .ZN(new_n1384_));
  NOR4_X1    g0742(.A1(new_n1370_), .A2(new_n1363_), .A3(new_n1382_), .A4(new_n1384_), .ZN(new_n1385_));
  NAND3_X1   g0743(.A1(new_n1380_), .A2(new_n1371_), .A3(new_n1385_), .ZN(new_n1386_));
  INV_X1     g0744(.I(new_n1386_), .ZN(new_n1387_));
  OAI21_X1   g0745(.A1(new_n1339_), .A2(new_n1361_), .B(new_n1387_), .ZN(new_n1388_));
  INV_X1     g0746(.I(\in1[113] ), .ZN(new_n1389_));
  NOR2_X1    g0747(.A1(new_n1389_), .A2(\in0[113] ), .ZN(new_n1390_));
  NOR2_X1    g0748(.A1(new_n1390_), .A2(\in1[112] ), .ZN(new_n1391_));
  INV_X1     g0749(.I(new_n1391_), .ZN(new_n1392_));
  INV_X1     g0750(.I(\in1[114] ), .ZN(new_n1393_));
  AOI21_X1   g0751(.A1(new_n1393_), .A2(\in0[114] ), .B(\in0[112] ), .ZN(new_n1394_));
  INV_X1     g0752(.I(new_n1394_), .ZN(new_n1395_));
  AOI21_X1   g0753(.A1(\in0[113] ), .A2(new_n1389_), .B(new_n1395_), .ZN(new_n1396_));
  INV_X1     g0754(.I(\in1[115] ), .ZN(new_n1397_));
  OAI22_X1   g0755(.A1(\in0[114] ), .A2(new_n1393_), .B1(new_n1397_), .B2(\in0[115] ), .ZN(new_n1398_));
  INV_X1     g0756(.I(new_n1398_), .ZN(new_n1399_));
  AOI21_X1   g0757(.A1(new_n1396_), .A2(new_n1392_), .B(new_n1399_), .ZN(new_n1400_));
  NAND2_X1   g0758(.A1(new_n1378_), .A2(\in0[108] ), .ZN(new_n1401_));
  INV_X1     g0759(.I(new_n1401_), .ZN(new_n1402_));
  NOR3_X1    g0760(.A1(new_n1402_), .A2(new_n1374_), .A3(new_n1377_), .ZN(new_n1403_));
  INV_X1     g0761(.I(\in1[110] ), .ZN(new_n1404_));
  AOI22_X1   g0762(.A1(\in0[110] ), .A2(new_n1404_), .B1(new_n1373_), .B2(\in1[111] ), .ZN(new_n1405_));
  INV_X1     g0763(.I(\in1[112] ), .ZN(new_n1406_));
  NAND2_X1   g0764(.A1(new_n1406_), .A2(\in0[112] ), .ZN(new_n1407_));
  NOR2_X1    g0765(.A1(new_n1390_), .A2(new_n1407_), .ZN(new_n1408_));
  AOI22_X1   g0766(.A1(new_n1399_), .A2(new_n1408_), .B1(\in0[115] ), .B2(new_n1397_), .ZN(new_n1409_));
  INV_X1     g0767(.I(new_n1409_), .ZN(new_n1410_));
  NOR4_X1    g0768(.A1(new_n1410_), .A2(new_n1400_), .A3(new_n1403_), .A4(new_n1405_), .ZN(new_n1411_));
  INV_X1     g0769(.I(\in1[118] ), .ZN(new_n1412_));
  INV_X1     g0770(.I(\in1[119] ), .ZN(new_n1413_));
  OAI22_X1   g0771(.A1(\in0[118] ), .A2(new_n1412_), .B1(new_n1413_), .B2(\in0[119] ), .ZN(new_n1414_));
  INV_X1     g0772(.I(new_n1414_), .ZN(new_n1415_));
  INV_X1     g0773(.I(\in0[119] ), .ZN(new_n1416_));
  AOI22_X1   g0774(.A1(\in0[118] ), .A2(new_n1412_), .B1(new_n1416_), .B2(\in1[119] ), .ZN(new_n1417_));
  INV_X1     g0775(.I(\in0[117] ), .ZN(new_n1418_));
  INV_X1     g0776(.I(\in1[116] ), .ZN(new_n1419_));
  AOI22_X1   g0777(.A1(\in0[116] ), .A2(new_n1419_), .B1(new_n1418_), .B2(\in1[117] ), .ZN(new_n1420_));
  AOI21_X1   g0778(.A1(new_n1414_), .A2(new_n1420_), .B(new_n1417_), .ZN(new_n1421_));
  INV_X1     g0779(.I(\in0[120] ), .ZN(new_n1422_));
  INV_X1     g0780(.I(\in0[122] ), .ZN(new_n1423_));
  INV_X1     g0781(.I(\in0[123] ), .ZN(new_n1424_));
  AOI22_X1   g0782(.A1(new_n1423_), .A2(\in1[122] ), .B1(new_n1424_), .B2(\in1[123] ), .ZN(new_n1425_));
  INV_X1     g0783(.I(new_n1425_), .ZN(new_n1426_));
  INV_X1     g0784(.I(\in1[121] ), .ZN(new_n1427_));
  NOR2_X1    g0785(.A1(new_n1427_), .A2(\in0[121] ), .ZN(new_n1428_));
  NOR4_X1    g0786(.A1(new_n1426_), .A2(new_n1422_), .A3(\in1[120] ), .A4(new_n1428_), .ZN(new_n1429_));
  INV_X1     g0787(.I(\in1[117] ), .ZN(new_n1430_));
  OAI22_X1   g0788(.A1(\in0[116] ), .A2(new_n1419_), .B1(new_n1430_), .B2(\in0[117] ), .ZN(new_n1431_));
  INV_X1     g0789(.I(new_n1431_), .ZN(new_n1432_));
  NOR4_X1    g0790(.A1(new_n1429_), .A2(new_n1415_), .A3(new_n1421_), .A4(new_n1432_), .ZN(new_n1433_));
  INV_X1     g0791(.I(new_n1433_), .ZN(new_n1434_));
  AOI21_X1   g0792(.A1(new_n1388_), .A2(new_n1411_), .B(new_n1434_), .ZN(new_n1435_));
  OAI22_X1   g0793(.A1(\in0[124] ), .A2(new_n1054_), .B1(new_n1048_), .B2(\in1[127] ), .ZN(new_n1436_));
  INV_X1     g0794(.I(new_n1436_), .ZN(new_n1437_));
  NOR2_X1    g0795(.A1(new_n1424_), .A2(\in1[123] ), .ZN(new_n1438_));
  NOR2_X1    g0796(.A1(new_n1428_), .A2(\in1[120] ), .ZN(new_n1439_));
  INV_X1     g0797(.I(new_n1439_), .ZN(new_n1440_));
  INV_X1     g0798(.I(\in1[122] ), .ZN(new_n1441_));
  AOI21_X1   g0799(.A1(new_n1441_), .A2(\in0[122] ), .B(\in0[120] ), .ZN(new_n1442_));
  INV_X1     g0800(.I(new_n1442_), .ZN(new_n1443_));
  AOI21_X1   g0801(.A1(\in0[121] ), .A2(new_n1427_), .B(new_n1443_), .ZN(new_n1444_));
  AOI21_X1   g0802(.A1(new_n1444_), .A2(new_n1440_), .B(new_n1425_), .ZN(new_n1445_));
  OAI22_X1   g0803(.A1(new_n1445_), .A2(new_n1438_), .B1(new_n1052_), .B2(new_n1437_), .ZN(new_n1446_));
  OAI21_X1   g0804(.A1(new_n1435_), .A2(new_n1446_), .B(new_n1061_), .ZN(new_n1447_));
  AOI21_X1   g0805(.A1(new_n1447_), .A2(new_n1049_), .B(new_n1048_), .ZN(new_n1448_));
  INV_X1     g0806(.I(new_n1448_), .ZN(new_n1449_));
  AOI21_X1   g0807(.A1(new_n1045_), .A2(new_n644_), .B(new_n1033_), .ZN(new_n1450_));
  NAND2_X1   g0808(.A1(new_n1449_), .A2(new_n1450_), .ZN(new_n1451_));
  NOR2_X1    g0809(.A1(new_n1449_), .A2(new_n1450_), .ZN(new_n1452_));
  NAND2_X1   g0810(.A1(new_n1096_), .A2(new_n1098_), .ZN(new_n1453_));
  NAND2_X1   g0811(.A1(new_n1100_), .A2(new_n1102_), .ZN(new_n1454_));
  NAND2_X1   g0812(.A1(new_n1453_), .A2(new_n1454_), .ZN(new_n1455_));
  NAND2_X1   g0813(.A1(new_n1105_), .A2(new_n1107_), .ZN(new_n1456_));
  INV_X1     g0814(.I(\in1[34] ), .ZN(new_n1457_));
  AOI22_X1   g0815(.A1(\in0[33] ), .A2(new_n1112_), .B1(new_n1457_), .B2(\in0[34] ), .ZN(new_n1458_));
  NOR4_X1    g0816(.A1(new_n1108_), .A2(\in0[32] ), .A3(\in1[32] ), .A4(\in1[33] ), .ZN(new_n1459_));
  OAI21_X1   g0817(.A1(new_n1458_), .A2(new_n1459_), .B(new_n1456_), .ZN(new_n1460_));
  INV_X1     g0818(.I(new_n1115_), .ZN(new_n1461_));
  AOI21_X1   g0819(.A1(new_n1460_), .A2(new_n1461_), .B(new_n1455_), .ZN(new_n1462_));
  NAND3_X1   g0820(.A1(new_n1118_), .A2(new_n1128_), .A3(new_n1125_), .ZN(new_n1463_));
  NOR2_X1    g0821(.A1(new_n1462_), .A2(new_n1463_), .ZN(new_n1464_));
  OAI22_X1   g0822(.A1(new_n1143_), .A2(\in1[49] ), .B1(new_n1158_), .B2(\in1[50] ), .ZN(new_n1465_));
  INV_X1     g0823(.I(\in1[48] ), .ZN(new_n1466_));
  NAND4_X1   g0824(.A1(new_n1160_), .A2(new_n1466_), .A3(new_n1141_), .A4(\in0[49] ), .ZN(new_n1467_));
  AOI21_X1   g0825(.A1(new_n1465_), .A2(new_n1467_), .B(new_n1159_), .ZN(new_n1468_));
  OAI21_X1   g0826(.A1(new_n1468_), .A2(new_n1147_), .B(new_n1157_), .ZN(new_n1469_));
  NOR4_X1    g0827(.A1(new_n1137_), .A2(new_n1159_), .A3(new_n1161_), .A4(new_n1162_), .ZN(new_n1470_));
  INV_X1     g0828(.I(\in0[56] ), .ZN(new_n1471_));
  AOI22_X1   g0829(.A1(new_n1471_), .A2(\in1[56] ), .B1(new_n1192_), .B2(\in1[57] ), .ZN(new_n1472_));
  INV_X1     g0830(.I(\in0[58] ), .ZN(new_n1473_));
  AOI22_X1   g0831(.A1(new_n1473_), .A2(\in1[58] ), .B1(new_n1190_), .B2(\in1[59] ), .ZN(new_n1474_));
  NOR2_X1    g0832(.A1(new_n1472_), .A2(new_n1474_), .ZN(new_n1475_));
  NOR2_X1    g0833(.A1(new_n1130_), .A2(\in1[54] ), .ZN(new_n1476_));
  NOR2_X1    g0834(.A1(new_n1133_), .A2(\in1[53] ), .ZN(new_n1477_));
  OAI22_X1   g0835(.A1(new_n1476_), .A2(new_n1477_), .B1(new_n1154_), .B2(new_n1156_), .ZN(new_n1478_));
  AOI22_X1   g0836(.A1(new_n1189_), .A2(new_n1475_), .B1(new_n1478_), .B2(new_n1152_), .ZN(new_n1479_));
  NAND3_X1   g0837(.A1(new_n1479_), .A2(new_n1469_), .A3(new_n1470_), .ZN(new_n1480_));
  AOI21_X1   g0838(.A1(new_n1464_), .A2(new_n1093_), .B(new_n1480_), .ZN(new_n1481_));
  NAND2_X1   g0839(.A1(new_n1195_), .A2(new_n1189_), .ZN(new_n1482_));
  NAND3_X1   g0840(.A1(new_n1482_), .A2(new_n1208_), .A3(new_n1219_), .ZN(new_n1483_));
  OAI21_X1   g0841(.A1(new_n1481_), .A2(new_n1483_), .B(new_n1242_), .ZN(new_n1484_));
  AOI21_X1   g0842(.A1(new_n1484_), .A2(new_n1264_), .B(new_n1290_), .ZN(new_n1485_));
  INV_X1     g0843(.I(new_n1315_), .ZN(new_n1486_));
  OAI21_X1   g0844(.A1(new_n1485_), .A2(new_n1486_), .B(new_n1337_), .ZN(new_n1487_));
  AOI21_X1   g0845(.A1(new_n1487_), .A2(new_n1360_), .B(new_n1386_), .ZN(new_n1488_));
  INV_X1     g0846(.I(new_n1411_), .ZN(new_n1489_));
  OAI21_X1   g0847(.A1(new_n1488_), .A2(new_n1489_), .B(new_n1433_), .ZN(new_n1490_));
  INV_X1     g0848(.I(new_n1446_), .ZN(new_n1491_));
  AOI21_X1   g0849(.A1(new_n1490_), .A2(new_n1491_), .B(new_n1060_), .ZN(new_n1492_));
  NOR2_X1    g0850(.A1(new_n1049_), .A2(\in0[127] ), .ZN(new_n1493_));
  NOR2_X1    g0851(.A1(new_n1492_), .A2(new_n1493_), .ZN(new_n1494_));
  NOR2_X1    g0852(.A1(new_n1494_), .A2(\in0[126] ), .ZN(new_n1495_));
  AOI21_X1   g0853(.A1(new_n1058_), .A2(new_n1494_), .B(new_n1495_), .ZN(new_n1496_));
  NOR2_X1    g0854(.A1(new_n1046_), .A2(\in3[126] ), .ZN(new_n1497_));
  AOI21_X1   g0855(.A1(new_n648_), .A2(new_n1046_), .B(new_n1497_), .ZN(new_n1498_));
  INV_X1     g0856(.I(new_n1498_), .ZN(new_n1499_));
  NAND2_X1   g0857(.A1(new_n1499_), .A2(new_n1496_), .ZN(new_n1500_));
  NOR2_X1    g0858(.A1(new_n1494_), .A2(\in0[125] ), .ZN(new_n1501_));
  AOI21_X1   g0859(.A1(new_n1055_), .A2(new_n1494_), .B(new_n1501_), .ZN(new_n1502_));
  NOR2_X1    g0860(.A1(new_n1046_), .A2(\in3[125] ), .ZN(new_n1503_));
  AOI21_X1   g0861(.A1(new_n647_), .A2(new_n1046_), .B(new_n1503_), .ZN(new_n1504_));
  INV_X1     g0862(.I(new_n1504_), .ZN(new_n1505_));
  OAI22_X1   g0863(.A1(new_n1496_), .A2(new_n1499_), .B1(new_n1505_), .B2(new_n1502_), .ZN(new_n1506_));
  NOR2_X1    g0864(.A1(new_n1494_), .A2(\in0[124] ), .ZN(new_n1507_));
  AOI21_X1   g0865(.A1(new_n1054_), .A2(new_n1494_), .B(new_n1507_), .ZN(new_n1508_));
  NAND2_X1   g0866(.A1(new_n677_), .A2(new_n667_), .ZN(new_n1509_));
  INV_X1     g0867(.I(new_n682_), .ZN(new_n1510_));
  NOR3_X1    g0868(.A1(new_n1510_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n1511_));
  NAND2_X1   g0869(.A1(new_n1509_), .A2(new_n1511_), .ZN(new_n1512_));
  INV_X1     g0870(.I(\in3[38] ), .ZN(new_n1513_));
  NOR2_X1    g0871(.A1(new_n1513_), .A2(\in2[38] ), .ZN(new_n1514_));
  INV_X1     g0872(.I(\in3[36] ), .ZN(new_n1515_));
  NOR2_X1    g0873(.A1(new_n1515_), .A2(\in2[36] ), .ZN(new_n1516_));
  OAI22_X1   g0874(.A1(new_n717_), .A2(new_n1514_), .B1(new_n719_), .B2(new_n1516_), .ZN(new_n1517_));
  INV_X1     g0875(.I(\in3[35] ), .ZN(new_n1518_));
  NOR2_X1    g0876(.A1(new_n1518_), .A2(\in2[35] ), .ZN(new_n1519_));
  INV_X1     g0877(.I(\in3[34] ), .ZN(new_n1520_));
  NOR2_X1    g0878(.A1(new_n1520_), .A2(\in2[34] ), .ZN(new_n1521_));
  AOI22_X1   g0879(.A1(\in2[33] ), .A2(new_n705_), .B1(new_n1520_), .B2(\in2[34] ), .ZN(new_n1522_));
  NOR4_X1    g0880(.A1(new_n701_), .A2(\in2[32] ), .A3(\in3[32] ), .A4(\in3[33] ), .ZN(new_n1523_));
  OAI22_X1   g0881(.A1(new_n1522_), .A2(new_n1523_), .B1(new_n1519_), .B2(new_n1521_), .ZN(new_n1524_));
  INV_X1     g0882(.I(new_n708_), .ZN(new_n1525_));
  AOI21_X1   g0883(.A1(new_n1524_), .A2(new_n1525_), .B(new_n1517_), .ZN(new_n1526_));
  AND2_X2    g0884(.A1(new_n712_), .A2(new_n667_), .Z(new_n1527_));
  NAND2_X1   g0885(.A1(new_n722_), .A2(new_n693_), .ZN(new_n1528_));
  OAI21_X1   g0886(.A1(\in2[38] ), .A2(new_n1513_), .B(new_n689_), .ZN(new_n1529_));
  NAND4_X1   g0887(.A1(new_n1529_), .A2(new_n720_), .A3(new_n1528_), .A4(new_n715_), .ZN(new_n1530_));
  NOR3_X1    g0888(.A1(new_n1527_), .A2(new_n1526_), .A3(new_n1530_), .ZN(new_n1531_));
  OAI22_X1   g0889(.A1(new_n740_), .A2(\in3[49] ), .B1(new_n755_), .B2(\in3[50] ), .ZN(new_n1532_));
  INV_X1     g0890(.I(\in3[48] ), .ZN(new_n1533_));
  NAND4_X1   g0891(.A1(new_n757_), .A2(new_n1533_), .A3(new_n738_), .A4(\in2[49] ), .ZN(new_n1534_));
  AOI21_X1   g0892(.A1(new_n1532_), .A2(new_n1534_), .B(new_n756_), .ZN(new_n1535_));
  NOR2_X1    g0893(.A1(new_n1535_), .A2(new_n744_), .ZN(new_n1536_));
  AOI22_X1   g0894(.A1(new_n798_), .A2(\in3[56] ), .B1(new_n796_), .B2(\in3[57] ), .ZN(new_n1537_));
  NOR2_X1    g0895(.A1(new_n1537_), .A2(new_n795_), .ZN(new_n1538_));
  NOR2_X1    g0896(.A1(new_n726_), .A2(\in3[54] ), .ZN(new_n1539_));
  NOR2_X1    g0897(.A1(new_n729_), .A2(\in3[53] ), .ZN(new_n1540_));
  OAI22_X1   g0898(.A1(new_n1539_), .A2(new_n1540_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n1541_));
  AOI22_X1   g0899(.A1(new_n792_), .A2(new_n1538_), .B1(new_n1541_), .B2(new_n749_), .ZN(new_n1542_));
  NAND4_X1   g0900(.A1(new_n1542_), .A2(new_n754_), .A3(new_n1536_), .A4(new_n760_), .ZN(new_n1543_));
  AOI21_X1   g0901(.A1(new_n1512_), .A2(new_n1531_), .B(new_n1543_), .ZN(new_n1544_));
  OAI21_X1   g0902(.A1(new_n1544_), .A2(new_n820_), .B(new_n842_), .ZN(new_n1545_));
  AOI21_X1   g0903(.A1(new_n1545_), .A2(new_n864_), .B(new_n889_), .ZN(new_n1546_));
  INV_X1     g0904(.I(new_n913_), .ZN(new_n1547_));
  OAI21_X1   g0905(.A1(new_n1546_), .A2(new_n1547_), .B(new_n935_), .ZN(new_n1548_));
  AOI21_X1   g0906(.A1(new_n1548_), .A2(new_n958_), .B(new_n984_), .ZN(new_n1549_));
  INV_X1     g0907(.I(new_n1008_), .ZN(new_n1550_));
  OAI21_X1   g0908(.A1(new_n1549_), .A2(new_n1550_), .B(new_n1030_), .ZN(new_n1551_));
  INV_X1     g0909(.I(new_n1044_), .ZN(new_n1552_));
  AOI21_X1   g0910(.A1(new_n1551_), .A2(new_n1552_), .B(new_n657_), .ZN(new_n1553_));
  NOR2_X1    g0911(.A1(new_n1553_), .A2(new_n645_), .ZN(new_n1554_));
  NOR2_X1    g0912(.A1(new_n1554_), .A2(\in2[124] ), .ZN(new_n1555_));
  AOI21_X1   g0913(.A1(new_n651_), .A2(new_n1554_), .B(new_n1555_), .ZN(new_n1556_));
  INV_X1     g0914(.I(new_n1556_), .ZN(new_n1557_));
  NAND2_X1   g0915(.A1(new_n1557_), .A2(new_n1508_), .ZN(new_n1558_));
  NAND2_X1   g0916(.A1(new_n1505_), .A2(new_n1502_), .ZN(new_n1559_));
  NAND3_X1   g0917(.A1(new_n1506_), .A2(new_n1558_), .A3(new_n1559_), .ZN(new_n1560_));
  AOI21_X1   g0918(.A1(new_n1560_), .A2(new_n1500_), .B(new_n1452_), .ZN(new_n1561_));
  INV_X1     g0919(.I(new_n1561_), .ZN(new_n1562_));
  INV_X1     g0920(.I(\in3[23] ), .ZN(new_n1563_));
  NOR2_X1    g0921(.A1(new_n1554_), .A2(\in2[23] ), .ZN(new_n1564_));
  AOI21_X1   g0922(.A1(new_n1563_), .A2(new_n1554_), .B(new_n1564_), .ZN(new_n1565_));
  INV_X1     g0923(.I(new_n1565_), .ZN(new_n1566_));
  NOR2_X1    g0924(.A1(new_n1494_), .A2(\in0[23] ), .ZN(new_n1567_));
  INV_X1     g0925(.I(new_n1494_), .ZN(new_n1568_));
  NOR2_X1    g0926(.A1(new_n1568_), .A2(\in1[23] ), .ZN(new_n1569_));
  NOR2_X1    g0927(.A1(new_n1569_), .A2(new_n1567_), .ZN(new_n1570_));
  NOR2_X1    g0928(.A1(new_n1566_), .A2(new_n1570_), .ZN(new_n1571_));
  INV_X1     g0929(.I(\in3[15] ), .ZN(new_n1572_));
  NOR2_X1    g0930(.A1(new_n1554_), .A2(\in2[15] ), .ZN(new_n1573_));
  AOI21_X1   g0931(.A1(new_n1572_), .A2(new_n1554_), .B(new_n1573_), .ZN(new_n1574_));
  INV_X1     g0932(.I(new_n1574_), .ZN(new_n1575_));
  NOR2_X1    g0933(.A1(new_n1494_), .A2(\in0[15] ), .ZN(new_n1576_));
  NOR2_X1    g0934(.A1(new_n1568_), .A2(\in1[15] ), .ZN(new_n1577_));
  NOR2_X1    g0935(.A1(new_n1577_), .A2(new_n1576_), .ZN(new_n1578_));
  NOR2_X1    g0936(.A1(new_n1575_), .A2(new_n1578_), .ZN(new_n1579_));
  INV_X1     g0937(.I(new_n1579_), .ZN(new_n1580_));
  INV_X1     g0938(.I(\in2[10] ), .ZN(new_n1581_));
  OAI21_X1   g0939(.A1(new_n1553_), .A2(new_n645_), .B(new_n1581_), .ZN(new_n1582_));
  INV_X1     g0940(.I(\in3[10] ), .ZN(new_n1583_));
  NAND3_X1   g0941(.A1(new_n1045_), .A2(new_n1583_), .A3(new_n646_), .ZN(new_n1584_));
  NAND2_X1   g0942(.A1(new_n1582_), .A2(new_n1584_), .ZN(new_n1585_));
  INV_X1     g0943(.I(new_n1493_), .ZN(new_n1586_));
  AOI21_X1   g0944(.A1(new_n1447_), .A2(new_n1586_), .B(\in0[10] ), .ZN(new_n1587_));
  NOR3_X1    g0945(.A1(new_n1492_), .A2(\in1[10] ), .A3(new_n1493_), .ZN(new_n1588_));
  NOR2_X1    g0946(.A1(new_n1587_), .A2(new_n1588_), .ZN(new_n1589_));
  NAND2_X1   g0947(.A1(new_n1589_), .A2(new_n1585_), .ZN(new_n1590_));
  AOI21_X1   g0948(.A1(new_n1045_), .A2(new_n646_), .B(\in2[10] ), .ZN(new_n1591_));
  AOI21_X1   g0949(.A1(new_n1583_), .A2(new_n1554_), .B(new_n1591_), .ZN(new_n1592_));
  INV_X1     g0950(.I(\in0[10] ), .ZN(new_n1593_));
  OAI21_X1   g0951(.A1(new_n1492_), .A2(new_n1493_), .B(new_n1593_), .ZN(new_n1594_));
  INV_X1     g0952(.I(\in1[10] ), .ZN(new_n1595_));
  NAND3_X1   g0953(.A1(new_n1447_), .A2(new_n1595_), .A3(new_n1586_), .ZN(new_n1596_));
  NAND2_X1   g0954(.A1(new_n1596_), .A2(new_n1594_), .ZN(new_n1597_));
  AOI21_X1   g0955(.A1(new_n1447_), .A2(new_n1586_), .B(\in0[9] ), .ZN(new_n1598_));
  NOR3_X1    g0956(.A1(new_n1492_), .A2(\in1[9] ), .A3(new_n1493_), .ZN(new_n1599_));
  NOR2_X1    g0957(.A1(new_n1598_), .A2(new_n1599_), .ZN(new_n1600_));
  INV_X1     g0958(.I(\in2[9] ), .ZN(new_n1601_));
  OAI21_X1   g0959(.A1(new_n1553_), .A2(new_n645_), .B(new_n1601_), .ZN(new_n1602_));
  INV_X1     g0960(.I(\in3[9] ), .ZN(new_n1603_));
  NAND3_X1   g0961(.A1(new_n1045_), .A2(new_n1603_), .A3(new_n646_), .ZN(new_n1604_));
  NAND2_X1   g0962(.A1(new_n1602_), .A2(new_n1604_), .ZN(new_n1605_));
  AOI22_X1   g0963(.A1(new_n1592_), .A2(new_n1597_), .B1(new_n1600_), .B2(new_n1605_), .ZN(new_n1606_));
  INV_X1     g0964(.I(\in2[11] ), .ZN(new_n1607_));
  NAND2_X1   g0965(.A1(new_n1046_), .A2(new_n1607_), .ZN(new_n1608_));
  OAI21_X1   g0966(.A1(\in3[11] ), .A2(new_n1046_), .B(new_n1608_), .ZN(new_n1609_));
  AOI21_X1   g0967(.A1(new_n1606_), .A2(new_n1590_), .B(new_n1609_), .ZN(new_n1610_));
  NOR2_X1    g0968(.A1(new_n1592_), .A2(new_n1597_), .ZN(new_n1611_));
  INV_X1     g0969(.I(\in0[9] ), .ZN(new_n1612_));
  OAI21_X1   g0970(.A1(new_n1492_), .A2(new_n1493_), .B(new_n1612_), .ZN(new_n1613_));
  INV_X1     g0971(.I(\in1[9] ), .ZN(new_n1614_));
  NAND3_X1   g0972(.A1(new_n1447_), .A2(new_n1614_), .A3(new_n1586_), .ZN(new_n1615_));
  NAND2_X1   g0973(.A1(new_n1615_), .A2(new_n1613_), .ZN(new_n1616_));
  AOI21_X1   g0974(.A1(new_n1045_), .A2(new_n646_), .B(\in2[9] ), .ZN(new_n1617_));
  NOR3_X1    g0975(.A1(new_n1553_), .A2(\in3[9] ), .A3(new_n645_), .ZN(new_n1618_));
  NOR2_X1    g0976(.A1(new_n1618_), .A2(new_n1617_), .ZN(new_n1619_));
  NOR2_X1    g0977(.A1(new_n1616_), .A2(new_n1619_), .ZN(new_n1620_));
  NOR2_X1    g0978(.A1(new_n1589_), .A2(new_n1585_), .ZN(new_n1621_));
  NOR2_X1    g0979(.A1(new_n1554_), .A2(\in2[11] ), .ZN(new_n1622_));
  NOR2_X1    g0980(.A1(new_n1046_), .A2(\in3[11] ), .ZN(new_n1623_));
  NOR2_X1    g0981(.A1(new_n1622_), .A2(new_n1623_), .ZN(new_n1624_));
  NOR4_X1    g0982(.A1(new_n1611_), .A2(new_n1620_), .A3(new_n1621_), .A4(new_n1624_), .ZN(new_n1625_));
  INV_X1     g0983(.I(\in1[11] ), .ZN(new_n1626_));
  NOR2_X1    g0984(.A1(new_n1494_), .A2(\in0[11] ), .ZN(new_n1627_));
  AOI21_X1   g0985(.A1(new_n1626_), .A2(new_n1494_), .B(new_n1627_), .ZN(new_n1628_));
  OAI21_X1   g0986(.A1(new_n1610_), .A2(new_n1625_), .B(new_n1628_), .ZN(new_n1629_));
  OAI22_X1   g0987(.A1(new_n1616_), .A2(new_n1619_), .B1(new_n1589_), .B2(new_n1585_), .ZN(new_n1630_));
  NOR2_X1    g0988(.A1(new_n1630_), .A2(new_n1611_), .ZN(new_n1631_));
  INV_X1     g0989(.I(\in1[12] ), .ZN(new_n1632_));
  NOR2_X1    g0990(.A1(new_n1494_), .A2(\in0[12] ), .ZN(new_n1633_));
  AOI21_X1   g0991(.A1(new_n1632_), .A2(new_n1494_), .B(new_n1633_), .ZN(new_n1634_));
  INV_X1     g0992(.I(\in3[12] ), .ZN(new_n1635_));
  NAND2_X1   g0993(.A1(new_n1554_), .A2(new_n1635_), .ZN(new_n1636_));
  OAI21_X1   g0994(.A1(\in2[12] ), .A2(new_n1554_), .B(new_n1636_), .ZN(new_n1637_));
  NAND2_X1   g0995(.A1(new_n1637_), .A2(new_n1634_), .ZN(new_n1638_));
  AOI21_X1   g0996(.A1(new_n1631_), .A2(new_n1609_), .B(new_n1638_), .ZN(new_n1639_));
  INV_X1     g0997(.I(\in3[13] ), .ZN(new_n1640_));
  NAND2_X1   g0998(.A1(new_n1554_), .A2(new_n1640_), .ZN(new_n1641_));
  OAI21_X1   g0999(.A1(\in2[13] ), .A2(new_n1554_), .B(new_n1641_), .ZN(new_n1642_));
  INV_X1     g1000(.I(\in1[13] ), .ZN(new_n1643_));
  NOR2_X1    g1001(.A1(new_n1494_), .A2(\in0[13] ), .ZN(new_n1644_));
  AOI21_X1   g1002(.A1(new_n1643_), .A2(new_n1494_), .B(new_n1644_), .ZN(new_n1645_));
  NAND2_X1   g1003(.A1(new_n1642_), .A2(new_n1645_), .ZN(new_n1646_));
  NOR2_X1    g1004(.A1(new_n1554_), .A2(\in2[13] ), .ZN(new_n1647_));
  AOI21_X1   g1005(.A1(new_n1640_), .A2(new_n1554_), .B(new_n1647_), .ZN(new_n1648_));
  NAND2_X1   g1006(.A1(new_n1494_), .A2(new_n1643_), .ZN(new_n1649_));
  OAI21_X1   g1007(.A1(\in0[13] ), .A2(new_n1494_), .B(new_n1649_), .ZN(new_n1650_));
  NAND2_X1   g1008(.A1(new_n1648_), .A2(new_n1650_), .ZN(new_n1651_));
  NAND3_X1   g1009(.A1(new_n1638_), .A2(new_n1646_), .A3(new_n1651_), .ZN(new_n1652_));
  AOI21_X1   g1010(.A1(new_n1629_), .A2(new_n1639_), .B(new_n1652_), .ZN(new_n1653_));
  INV_X1     g1011(.I(\in3[14] ), .ZN(new_n1654_));
  NOR2_X1    g1012(.A1(new_n1554_), .A2(\in2[14] ), .ZN(new_n1655_));
  AOI21_X1   g1013(.A1(new_n1654_), .A2(new_n1554_), .B(new_n1655_), .ZN(new_n1656_));
  INV_X1     g1014(.I(new_n1656_), .ZN(new_n1657_));
  NOR2_X1    g1015(.A1(new_n1653_), .A2(new_n1657_), .ZN(new_n1658_));
  OAI21_X1   g1016(.A1(new_n1630_), .A2(new_n1611_), .B(new_n1624_), .ZN(new_n1659_));
  NAND3_X1   g1017(.A1(new_n1606_), .A2(new_n1590_), .A3(new_n1609_), .ZN(new_n1660_));
  INV_X1     g1018(.I(new_n1628_), .ZN(new_n1661_));
  AOI21_X1   g1019(.A1(new_n1659_), .A2(new_n1660_), .B(new_n1661_), .ZN(new_n1662_));
  NAND2_X1   g1020(.A1(new_n1606_), .A2(new_n1590_), .ZN(new_n1663_));
  NOR2_X1    g1021(.A1(new_n1568_), .A2(\in1[12] ), .ZN(new_n1664_));
  NOR2_X1    g1022(.A1(new_n1554_), .A2(\in2[12] ), .ZN(new_n1665_));
  AOI21_X1   g1023(.A1(new_n1635_), .A2(new_n1554_), .B(new_n1665_), .ZN(new_n1666_));
  NOR3_X1    g1024(.A1(new_n1666_), .A2(new_n1633_), .A3(new_n1664_), .ZN(new_n1667_));
  OAI21_X1   g1025(.A1(new_n1663_), .A2(new_n1624_), .B(new_n1667_), .ZN(new_n1668_));
  NOR2_X1    g1026(.A1(new_n1648_), .A2(new_n1650_), .ZN(new_n1669_));
  NOR2_X1    g1027(.A1(new_n1642_), .A2(new_n1645_), .ZN(new_n1670_));
  NOR3_X1    g1028(.A1(new_n1667_), .A2(new_n1670_), .A3(new_n1669_), .ZN(new_n1671_));
  OAI21_X1   g1029(.A1(new_n1662_), .A2(new_n1668_), .B(new_n1671_), .ZN(new_n1672_));
  NOR2_X1    g1030(.A1(new_n1672_), .A2(new_n1656_), .ZN(new_n1673_));
  INV_X1     g1031(.I(\in1[14] ), .ZN(new_n1674_));
  NOR2_X1    g1032(.A1(new_n1494_), .A2(\in0[14] ), .ZN(new_n1675_));
  AOI21_X1   g1033(.A1(new_n1674_), .A2(new_n1494_), .B(new_n1675_), .ZN(new_n1676_));
  OAI22_X1   g1034(.A1(new_n1673_), .A2(new_n1658_), .B1(new_n1653_), .B2(new_n1676_), .ZN(new_n1677_));
  NAND2_X1   g1035(.A1(new_n1575_), .A2(new_n1578_), .ZN(new_n1678_));
  INV_X1     g1036(.I(new_n1678_), .ZN(new_n1679_));
  OAI21_X1   g1037(.A1(new_n1677_), .A2(new_n1679_), .B(new_n1580_), .ZN(new_n1680_));
  INV_X1     g1038(.I(\in3[16] ), .ZN(new_n1681_));
  NOR2_X1    g1039(.A1(new_n1554_), .A2(\in2[16] ), .ZN(new_n1682_));
  AOI21_X1   g1040(.A1(new_n1681_), .A2(new_n1554_), .B(new_n1682_), .ZN(new_n1683_));
  INV_X1     g1041(.I(\in1[16] ), .ZN(new_n1684_));
  NOR2_X1    g1042(.A1(new_n1494_), .A2(\in0[16] ), .ZN(new_n1685_));
  AOI21_X1   g1043(.A1(new_n1684_), .A2(new_n1494_), .B(new_n1685_), .ZN(new_n1686_));
  INV_X1     g1044(.I(new_n1686_), .ZN(new_n1687_));
  NOR2_X1    g1045(.A1(new_n1687_), .A2(new_n1683_), .ZN(new_n1688_));
  INV_X1     g1046(.I(new_n1688_), .ZN(new_n1689_));
  NOR2_X1    g1047(.A1(new_n1494_), .A2(\in0[17] ), .ZN(new_n1690_));
  NOR2_X1    g1048(.A1(new_n1568_), .A2(\in1[17] ), .ZN(new_n1691_));
  NOR2_X1    g1049(.A1(new_n1691_), .A2(new_n1690_), .ZN(new_n1692_));
  INV_X1     g1050(.I(\in3[17] ), .ZN(new_n1693_));
  NOR2_X1    g1051(.A1(new_n1554_), .A2(\in2[17] ), .ZN(new_n1694_));
  AOI21_X1   g1052(.A1(new_n1693_), .A2(new_n1554_), .B(new_n1694_), .ZN(new_n1695_));
  INV_X1     g1053(.I(new_n1695_), .ZN(new_n1696_));
  NAND2_X1   g1054(.A1(new_n1696_), .A2(new_n1692_), .ZN(new_n1697_));
  AOI21_X1   g1055(.A1(new_n1683_), .A2(new_n1687_), .B(new_n1697_), .ZN(new_n1698_));
  INV_X1     g1056(.I(new_n1698_), .ZN(new_n1699_));
  AOI21_X1   g1057(.A1(new_n1680_), .A2(new_n1689_), .B(new_n1699_), .ZN(new_n1700_));
  INV_X1     g1058(.I(new_n1697_), .ZN(new_n1701_));
  INV_X1     g1059(.I(\in3[18] ), .ZN(new_n1702_));
  NOR2_X1    g1060(.A1(new_n1554_), .A2(\in2[18] ), .ZN(new_n1703_));
  AOI21_X1   g1061(.A1(new_n1702_), .A2(new_n1554_), .B(new_n1703_), .ZN(new_n1704_));
  INV_X1     g1062(.I(\in1[18] ), .ZN(new_n1705_));
  NOR2_X1    g1063(.A1(new_n1494_), .A2(\in0[18] ), .ZN(new_n1706_));
  AOI21_X1   g1064(.A1(new_n1705_), .A2(new_n1494_), .B(new_n1706_), .ZN(new_n1707_));
  INV_X1     g1065(.I(new_n1707_), .ZN(new_n1708_));
  NOR2_X1    g1066(.A1(new_n1708_), .A2(new_n1704_), .ZN(new_n1709_));
  INV_X1     g1067(.I(new_n1704_), .ZN(new_n1710_));
  NOR2_X1    g1068(.A1(new_n1710_), .A2(new_n1707_), .ZN(new_n1711_));
  NOR3_X1    g1069(.A1(new_n1701_), .A2(new_n1711_), .A3(new_n1709_), .ZN(new_n1712_));
  INV_X1     g1070(.I(new_n1712_), .ZN(new_n1713_));
  INV_X1     g1071(.I(\in3[19] ), .ZN(new_n1714_));
  NOR2_X1    g1072(.A1(new_n1554_), .A2(\in2[19] ), .ZN(new_n1715_));
  AOI21_X1   g1073(.A1(new_n1714_), .A2(new_n1554_), .B(new_n1715_), .ZN(new_n1716_));
  OAI21_X1   g1074(.A1(new_n1700_), .A2(new_n1713_), .B(new_n1716_), .ZN(new_n1717_));
  NAND2_X1   g1075(.A1(new_n1672_), .A2(new_n1656_), .ZN(new_n1718_));
  NAND2_X1   g1076(.A1(new_n1629_), .A2(new_n1639_), .ZN(new_n1719_));
  NAND3_X1   g1077(.A1(new_n1719_), .A2(new_n1671_), .A3(new_n1657_), .ZN(new_n1720_));
  INV_X1     g1078(.I(new_n1676_), .ZN(new_n1721_));
  AOI22_X1   g1079(.A1(new_n1718_), .A2(new_n1720_), .B1(new_n1672_), .B2(new_n1721_), .ZN(new_n1722_));
  AOI21_X1   g1080(.A1(new_n1722_), .A2(new_n1678_), .B(new_n1579_), .ZN(new_n1723_));
  OAI21_X1   g1081(.A1(new_n1723_), .A2(new_n1688_), .B(new_n1698_), .ZN(new_n1724_));
  INV_X1     g1082(.I(new_n1716_), .ZN(new_n1725_));
  NAND3_X1   g1083(.A1(new_n1724_), .A2(new_n1712_), .A3(new_n1725_), .ZN(new_n1726_));
  INV_X1     g1084(.I(\in1[19] ), .ZN(new_n1727_));
  NOR2_X1    g1085(.A1(new_n1494_), .A2(\in0[19] ), .ZN(new_n1728_));
  AOI21_X1   g1086(.A1(new_n1727_), .A2(new_n1494_), .B(new_n1728_), .ZN(new_n1729_));
  INV_X1     g1087(.I(new_n1729_), .ZN(new_n1730_));
  AOI21_X1   g1088(.A1(new_n1717_), .A2(new_n1726_), .B(new_n1730_), .ZN(new_n1731_));
  NOR2_X1    g1089(.A1(new_n1494_), .A2(\in0[20] ), .ZN(new_n1732_));
  NOR2_X1    g1090(.A1(new_n1568_), .A2(\in1[20] ), .ZN(new_n1733_));
  NOR2_X1    g1091(.A1(new_n1733_), .A2(new_n1732_), .ZN(new_n1734_));
  INV_X1     g1092(.I(\in3[20] ), .ZN(new_n1735_));
  NOR2_X1    g1093(.A1(new_n1554_), .A2(\in2[20] ), .ZN(new_n1736_));
  AOI21_X1   g1094(.A1(new_n1735_), .A2(new_n1554_), .B(new_n1736_), .ZN(new_n1737_));
  INV_X1     g1095(.I(new_n1737_), .ZN(new_n1738_));
  NAND2_X1   g1096(.A1(new_n1738_), .A2(new_n1734_), .ZN(new_n1739_));
  INV_X1     g1097(.I(new_n1739_), .ZN(new_n1740_));
  NAND3_X1   g1098(.A1(new_n1724_), .A2(new_n1712_), .A3(new_n1725_), .ZN(new_n1741_));
  NAND2_X1   g1099(.A1(new_n1741_), .A2(new_n1740_), .ZN(new_n1742_));
  INV_X1     g1100(.I(\in3[21] ), .ZN(new_n1743_));
  NOR2_X1    g1101(.A1(new_n1554_), .A2(\in2[21] ), .ZN(new_n1744_));
  AOI21_X1   g1102(.A1(new_n1743_), .A2(new_n1554_), .B(new_n1744_), .ZN(new_n1745_));
  INV_X1     g1103(.I(\in1[21] ), .ZN(new_n1746_));
  NOR2_X1    g1104(.A1(new_n1494_), .A2(\in0[21] ), .ZN(new_n1747_));
  AOI21_X1   g1105(.A1(new_n1746_), .A2(new_n1494_), .B(new_n1747_), .ZN(new_n1748_));
  INV_X1     g1106(.I(new_n1748_), .ZN(new_n1749_));
  NOR2_X1    g1107(.A1(new_n1749_), .A2(new_n1745_), .ZN(new_n1750_));
  INV_X1     g1108(.I(new_n1745_), .ZN(new_n1751_));
  NOR2_X1    g1109(.A1(new_n1751_), .A2(new_n1748_), .ZN(new_n1752_));
  NOR3_X1    g1110(.A1(new_n1740_), .A2(new_n1752_), .A3(new_n1750_), .ZN(new_n1753_));
  OAI21_X1   g1111(.A1(new_n1731_), .A2(new_n1742_), .B(new_n1753_), .ZN(new_n1754_));
  INV_X1     g1112(.I(\in3[22] ), .ZN(new_n1755_));
  NOR2_X1    g1113(.A1(new_n1554_), .A2(\in2[22] ), .ZN(new_n1756_));
  AOI21_X1   g1114(.A1(new_n1755_), .A2(new_n1554_), .B(new_n1756_), .ZN(new_n1757_));
  NAND2_X1   g1115(.A1(new_n1754_), .A2(new_n1757_), .ZN(new_n1758_));
  AOI21_X1   g1116(.A1(new_n1724_), .A2(new_n1712_), .B(new_n1725_), .ZN(new_n1759_));
  NOR3_X1    g1117(.A1(new_n1700_), .A2(new_n1713_), .A3(new_n1716_), .ZN(new_n1760_));
  OAI21_X1   g1118(.A1(new_n1760_), .A2(new_n1759_), .B(new_n1729_), .ZN(new_n1761_));
  NOR2_X1    g1119(.A1(new_n1700_), .A2(new_n1713_), .ZN(new_n1762_));
  AOI21_X1   g1120(.A1(new_n1762_), .A2(new_n1725_), .B(new_n1739_), .ZN(new_n1763_));
  NAND2_X1   g1121(.A1(new_n1761_), .A2(new_n1763_), .ZN(new_n1764_));
  INV_X1     g1122(.I(new_n1757_), .ZN(new_n1765_));
  NAND3_X1   g1123(.A1(new_n1764_), .A2(new_n1753_), .A3(new_n1765_), .ZN(new_n1766_));
  INV_X1     g1124(.I(\in1[22] ), .ZN(new_n1767_));
  NOR2_X1    g1125(.A1(new_n1494_), .A2(\in0[22] ), .ZN(new_n1768_));
  AOI21_X1   g1126(.A1(new_n1767_), .A2(new_n1494_), .B(new_n1768_), .ZN(new_n1769_));
  INV_X1     g1127(.I(new_n1769_), .ZN(new_n1770_));
  AOI22_X1   g1128(.A1(new_n1758_), .A2(new_n1766_), .B1(new_n1754_), .B2(new_n1770_), .ZN(new_n1771_));
  NAND2_X1   g1129(.A1(new_n1566_), .A2(new_n1570_), .ZN(new_n1772_));
  AOI21_X1   g1130(.A1(new_n1771_), .A2(new_n1772_), .B(new_n1571_), .ZN(new_n1773_));
  INV_X1     g1131(.I(\in3[24] ), .ZN(new_n1774_));
  NOR2_X1    g1132(.A1(new_n1554_), .A2(\in2[24] ), .ZN(new_n1775_));
  AOI21_X1   g1133(.A1(new_n1774_), .A2(new_n1554_), .B(new_n1775_), .ZN(new_n1776_));
  INV_X1     g1134(.I(\in1[24] ), .ZN(new_n1777_));
  NOR2_X1    g1135(.A1(new_n1494_), .A2(\in0[24] ), .ZN(new_n1778_));
  AOI21_X1   g1136(.A1(new_n1777_), .A2(new_n1494_), .B(new_n1778_), .ZN(new_n1779_));
  INV_X1     g1137(.I(new_n1779_), .ZN(new_n1780_));
  NOR2_X1    g1138(.A1(new_n1780_), .A2(new_n1776_), .ZN(new_n1781_));
  NOR2_X1    g1139(.A1(new_n1494_), .A2(\in0[25] ), .ZN(new_n1782_));
  NOR2_X1    g1140(.A1(new_n1568_), .A2(\in1[25] ), .ZN(new_n1783_));
  NOR2_X1    g1141(.A1(new_n1783_), .A2(new_n1782_), .ZN(new_n1784_));
  INV_X1     g1142(.I(\in3[25] ), .ZN(new_n1785_));
  NOR2_X1    g1143(.A1(new_n1554_), .A2(\in2[25] ), .ZN(new_n1786_));
  AOI21_X1   g1144(.A1(new_n1785_), .A2(new_n1554_), .B(new_n1786_), .ZN(new_n1787_));
  INV_X1     g1145(.I(new_n1787_), .ZN(new_n1788_));
  NAND2_X1   g1146(.A1(new_n1788_), .A2(new_n1784_), .ZN(new_n1789_));
  AOI21_X1   g1147(.A1(new_n1776_), .A2(new_n1780_), .B(new_n1789_), .ZN(new_n1790_));
  OAI21_X1   g1148(.A1(new_n1773_), .A2(new_n1781_), .B(new_n1790_), .ZN(new_n1791_));
  INV_X1     g1149(.I(new_n1789_), .ZN(new_n1792_));
  INV_X1     g1150(.I(\in3[26] ), .ZN(new_n1793_));
  NOR2_X1    g1151(.A1(new_n1554_), .A2(\in2[26] ), .ZN(new_n1794_));
  AOI21_X1   g1152(.A1(new_n1793_), .A2(new_n1554_), .B(new_n1794_), .ZN(new_n1795_));
  INV_X1     g1153(.I(\in1[26] ), .ZN(new_n1796_));
  NOR2_X1    g1154(.A1(new_n1494_), .A2(\in0[26] ), .ZN(new_n1797_));
  AOI21_X1   g1155(.A1(new_n1796_), .A2(new_n1494_), .B(new_n1797_), .ZN(new_n1798_));
  INV_X1     g1156(.I(new_n1798_), .ZN(new_n1799_));
  NOR2_X1    g1157(.A1(new_n1799_), .A2(new_n1795_), .ZN(new_n1800_));
  INV_X1     g1158(.I(new_n1795_), .ZN(new_n1801_));
  NOR2_X1    g1159(.A1(new_n1801_), .A2(new_n1798_), .ZN(new_n1802_));
  NOR3_X1    g1160(.A1(new_n1792_), .A2(new_n1802_), .A3(new_n1800_), .ZN(new_n1803_));
  INV_X1     g1161(.I(\in3[27] ), .ZN(new_n1804_));
  NOR2_X1    g1162(.A1(new_n1554_), .A2(\in2[27] ), .ZN(new_n1805_));
  AOI21_X1   g1163(.A1(new_n1804_), .A2(new_n1554_), .B(new_n1805_), .ZN(new_n1806_));
  INV_X1     g1164(.I(new_n1806_), .ZN(new_n1807_));
  AOI21_X1   g1165(.A1(new_n1791_), .A2(new_n1803_), .B(new_n1807_), .ZN(new_n1808_));
  INV_X1     g1166(.I(new_n1571_), .ZN(new_n1809_));
  INV_X1     g1167(.I(new_n1753_), .ZN(new_n1810_));
  AOI21_X1   g1168(.A1(new_n1761_), .A2(new_n1763_), .B(new_n1810_), .ZN(new_n1811_));
  NOR2_X1    g1169(.A1(new_n1811_), .A2(new_n1765_), .ZN(new_n1812_));
  NOR2_X1    g1170(.A1(new_n1754_), .A2(new_n1757_), .ZN(new_n1813_));
  OAI22_X1   g1171(.A1(new_n1812_), .A2(new_n1813_), .B1(new_n1811_), .B2(new_n1769_), .ZN(new_n1814_));
  INV_X1     g1172(.I(new_n1772_), .ZN(new_n1815_));
  OAI21_X1   g1173(.A1(new_n1814_), .A2(new_n1815_), .B(new_n1809_), .ZN(new_n1816_));
  INV_X1     g1174(.I(new_n1781_), .ZN(new_n1817_));
  INV_X1     g1175(.I(new_n1790_), .ZN(new_n1818_));
  AOI21_X1   g1176(.A1(new_n1816_), .A2(new_n1817_), .B(new_n1818_), .ZN(new_n1819_));
  INV_X1     g1177(.I(new_n1803_), .ZN(new_n1820_));
  NOR3_X1    g1178(.A1(new_n1819_), .A2(new_n1820_), .A3(new_n1806_), .ZN(new_n1821_));
  INV_X1     g1179(.I(\in1[27] ), .ZN(new_n1822_));
  NOR2_X1    g1180(.A1(new_n1494_), .A2(\in0[27] ), .ZN(new_n1823_));
  AOI21_X1   g1181(.A1(new_n1822_), .A2(new_n1494_), .B(new_n1823_), .ZN(new_n1824_));
  OAI21_X1   g1182(.A1(new_n1821_), .A2(new_n1808_), .B(new_n1824_), .ZN(new_n1825_));
  NOR2_X1    g1183(.A1(new_n1819_), .A2(new_n1820_), .ZN(new_n1826_));
  NOR2_X1    g1184(.A1(new_n1494_), .A2(\in0[28] ), .ZN(new_n1827_));
  NOR2_X1    g1185(.A1(new_n1568_), .A2(\in1[28] ), .ZN(new_n1828_));
  NOR2_X1    g1186(.A1(new_n1828_), .A2(new_n1827_), .ZN(new_n1829_));
  INV_X1     g1187(.I(\in3[28] ), .ZN(new_n1830_));
  NOR2_X1    g1188(.A1(new_n1554_), .A2(\in2[28] ), .ZN(new_n1831_));
  AOI21_X1   g1189(.A1(new_n1830_), .A2(new_n1554_), .B(new_n1831_), .ZN(new_n1832_));
  INV_X1     g1190(.I(new_n1832_), .ZN(new_n1833_));
  NAND2_X1   g1191(.A1(new_n1833_), .A2(new_n1829_), .ZN(new_n1834_));
  AOI21_X1   g1192(.A1(new_n1826_), .A2(new_n1807_), .B(new_n1834_), .ZN(new_n1835_));
  INV_X1     g1193(.I(new_n1834_), .ZN(new_n1836_));
  INV_X1     g1194(.I(\in3[29] ), .ZN(new_n1837_));
  NOR2_X1    g1195(.A1(new_n1554_), .A2(\in2[29] ), .ZN(new_n1838_));
  AOI21_X1   g1196(.A1(new_n1837_), .A2(new_n1554_), .B(new_n1838_), .ZN(new_n1839_));
  INV_X1     g1197(.I(\in1[29] ), .ZN(new_n1840_));
  NOR2_X1    g1198(.A1(new_n1494_), .A2(\in0[29] ), .ZN(new_n1841_));
  AOI21_X1   g1199(.A1(new_n1840_), .A2(new_n1494_), .B(new_n1841_), .ZN(new_n1842_));
  INV_X1     g1200(.I(new_n1842_), .ZN(new_n1843_));
  NOR2_X1    g1201(.A1(new_n1843_), .A2(new_n1839_), .ZN(new_n1844_));
  INV_X1     g1202(.I(new_n1839_), .ZN(new_n1845_));
  NOR2_X1    g1203(.A1(new_n1845_), .A2(new_n1842_), .ZN(new_n1846_));
  NOR3_X1    g1204(.A1(new_n1836_), .A2(new_n1846_), .A3(new_n1844_), .ZN(new_n1847_));
  INV_X1     g1205(.I(new_n1847_), .ZN(new_n1848_));
  AOI21_X1   g1206(.A1(new_n1825_), .A2(new_n1835_), .B(new_n1848_), .ZN(new_n1849_));
  INV_X1     g1207(.I(\in3[30] ), .ZN(new_n1850_));
  NOR2_X1    g1208(.A1(new_n1554_), .A2(\in2[30] ), .ZN(new_n1851_));
  AOI21_X1   g1209(.A1(new_n1850_), .A2(new_n1554_), .B(new_n1851_), .ZN(new_n1852_));
  INV_X1     g1210(.I(new_n1852_), .ZN(new_n1853_));
  NAND2_X1   g1211(.A1(new_n1849_), .A2(new_n1853_), .ZN(new_n1854_));
  NOR2_X1    g1212(.A1(new_n1849_), .A2(new_n1853_), .ZN(new_n1855_));
  OAI21_X1   g1213(.A1(new_n1819_), .A2(new_n1820_), .B(new_n1806_), .ZN(new_n1856_));
  NAND3_X1   g1214(.A1(new_n1791_), .A2(new_n1803_), .A3(new_n1807_), .ZN(new_n1857_));
  INV_X1     g1215(.I(new_n1824_), .ZN(new_n1858_));
  AOI21_X1   g1216(.A1(new_n1856_), .A2(new_n1857_), .B(new_n1858_), .ZN(new_n1859_));
  NAND3_X1   g1217(.A1(new_n1791_), .A2(new_n1803_), .A3(new_n1807_), .ZN(new_n1860_));
  NAND2_X1   g1218(.A1(new_n1860_), .A2(new_n1836_), .ZN(new_n1861_));
  OAI21_X1   g1219(.A1(new_n1859_), .A2(new_n1861_), .B(new_n1847_), .ZN(new_n1862_));
  NOR2_X1    g1220(.A1(new_n1862_), .A2(new_n1852_), .ZN(new_n1863_));
  INV_X1     g1221(.I(\in1[30] ), .ZN(new_n1864_));
  NOR2_X1    g1222(.A1(new_n1494_), .A2(\in0[30] ), .ZN(new_n1865_));
  AOI21_X1   g1223(.A1(new_n1864_), .A2(new_n1494_), .B(new_n1865_), .ZN(new_n1866_));
  OAI21_X1   g1224(.A1(new_n1855_), .A2(new_n1863_), .B(new_n1866_), .ZN(new_n1867_));
  NOR2_X1    g1225(.A1(new_n1494_), .A2(\in0[31] ), .ZN(new_n1868_));
  AOI21_X1   g1226(.A1(new_n1123_), .A2(new_n1494_), .B(new_n1868_), .ZN(new_n1869_));
  INV_X1     g1227(.I(new_n1869_), .ZN(new_n1870_));
  NAND3_X1   g1228(.A1(new_n1867_), .A2(new_n1854_), .A3(new_n1870_), .ZN(new_n1871_));
  NAND2_X1   g1229(.A1(new_n1862_), .A2(new_n1852_), .ZN(new_n1872_));
  NAND2_X1   g1230(.A1(new_n1849_), .A2(new_n1853_), .ZN(new_n1873_));
  INV_X1     g1231(.I(new_n1866_), .ZN(new_n1874_));
  AOI22_X1   g1232(.A1(new_n1873_), .A2(new_n1872_), .B1(new_n1862_), .B2(new_n1874_), .ZN(new_n1875_));
  NAND2_X1   g1233(.A1(new_n1875_), .A2(new_n1869_), .ZN(new_n1876_));
  OAI22_X1   g1234(.A1(new_n1855_), .A2(new_n1863_), .B1(new_n1849_), .B2(new_n1866_), .ZN(new_n1877_));
  NOR2_X1    g1235(.A1(new_n1046_), .A2(\in3[38] ), .ZN(new_n1878_));
  AOI21_X1   g1236(.A1(new_n690_), .A2(new_n1046_), .B(new_n1878_), .ZN(new_n1879_));
  INV_X1     g1237(.I(new_n1879_), .ZN(new_n1880_));
  NOR2_X1    g1238(.A1(new_n1568_), .A2(\in1[38] ), .ZN(new_n1881_));
  AOI21_X1   g1239(.A1(new_n1097_), .A2(new_n1568_), .B(new_n1881_), .ZN(new_n1882_));
  NOR2_X1    g1240(.A1(new_n1046_), .A2(\in3[39] ), .ZN(new_n1883_));
  AOI21_X1   g1241(.A1(new_n688_), .A2(new_n1046_), .B(new_n1883_), .ZN(new_n1884_));
  INV_X1     g1242(.I(new_n1884_), .ZN(new_n1885_));
  NOR2_X1    g1243(.A1(new_n1494_), .A2(\in0[39] ), .ZN(new_n1886_));
  AOI21_X1   g1244(.A1(new_n1119_), .A2(new_n1494_), .B(new_n1886_), .ZN(new_n1887_));
  OAI22_X1   g1245(.A1(new_n1880_), .A2(new_n1882_), .B1(new_n1885_), .B2(new_n1887_), .ZN(new_n1888_));
  NOR2_X1    g1246(.A1(new_n1046_), .A2(\in3[37] ), .ZN(new_n1889_));
  AOI21_X1   g1247(.A1(new_n692_), .A2(new_n1046_), .B(new_n1889_), .ZN(new_n1890_));
  INV_X1     g1248(.I(new_n1890_), .ZN(new_n1891_));
  NOR2_X1    g1249(.A1(new_n1494_), .A2(\in0[37] ), .ZN(new_n1892_));
  AOI21_X1   g1250(.A1(new_n1121_), .A2(new_n1494_), .B(new_n1892_), .ZN(new_n1893_));
  NOR2_X1    g1251(.A1(new_n1891_), .A2(new_n1893_), .ZN(new_n1894_));
  NOR2_X1    g1252(.A1(new_n1046_), .A2(\in3[36] ), .ZN(new_n1895_));
  AOI21_X1   g1253(.A1(new_n694_), .A2(new_n1046_), .B(new_n1895_), .ZN(new_n1896_));
  INV_X1     g1254(.I(new_n1896_), .ZN(new_n1897_));
  INV_X1     g1255(.I(\in1[36] ), .ZN(new_n1898_));
  NOR2_X1    g1256(.A1(new_n1494_), .A2(\in0[36] ), .ZN(new_n1899_));
  AOI21_X1   g1257(.A1(new_n1898_), .A2(new_n1494_), .B(new_n1899_), .ZN(new_n1900_));
  NOR4_X1    g1258(.A1(new_n1888_), .A2(new_n1894_), .A3(new_n1897_), .A4(new_n1900_), .ZN(new_n1901_));
  NOR2_X1    g1259(.A1(new_n1494_), .A2(\in0[32] ), .ZN(new_n1902_));
  AOI21_X1   g1260(.A1(new_n1111_), .A2(new_n1494_), .B(new_n1902_), .ZN(new_n1903_));
  NOR2_X1    g1261(.A1(new_n1046_), .A2(\in3[32] ), .ZN(new_n1904_));
  AOI21_X1   g1262(.A1(new_n703_), .A2(new_n1046_), .B(new_n1904_), .ZN(new_n1905_));
  INV_X1     g1263(.I(new_n1905_), .ZN(new_n1906_));
  NOR2_X1    g1264(.A1(new_n1046_), .A2(\in3[35] ), .ZN(new_n1907_));
  AOI21_X1   g1265(.A1(new_n697_), .A2(new_n1046_), .B(new_n1907_), .ZN(new_n1908_));
  INV_X1     g1266(.I(\in1[35] ), .ZN(new_n1909_));
  NOR2_X1    g1267(.A1(new_n1494_), .A2(\in0[35] ), .ZN(new_n1910_));
  AOI21_X1   g1268(.A1(new_n1909_), .A2(new_n1494_), .B(new_n1910_), .ZN(new_n1911_));
  INV_X1     g1269(.I(new_n1911_), .ZN(new_n1912_));
  NOR2_X1    g1270(.A1(new_n1046_), .A2(\in3[33] ), .ZN(new_n1913_));
  AOI21_X1   g1271(.A1(new_n701_), .A2(new_n1046_), .B(new_n1913_), .ZN(new_n1914_));
  NOR2_X1    g1272(.A1(new_n1494_), .A2(\in0[33] ), .ZN(new_n1915_));
  AOI21_X1   g1273(.A1(new_n1112_), .A2(new_n1494_), .B(new_n1915_), .ZN(new_n1916_));
  INV_X1     g1274(.I(new_n1916_), .ZN(new_n1917_));
  AOI22_X1   g1275(.A1(new_n1908_), .A2(new_n1912_), .B1(new_n1917_), .B2(new_n1914_), .ZN(new_n1918_));
  NOR2_X1    g1276(.A1(new_n1494_), .A2(\in0[34] ), .ZN(new_n1919_));
  AOI21_X1   g1277(.A1(new_n1457_), .A2(new_n1494_), .B(new_n1919_), .ZN(new_n1920_));
  NOR2_X1    g1278(.A1(new_n1046_), .A2(\in3[34] ), .ZN(new_n1921_));
  AOI21_X1   g1279(.A1(new_n699_), .A2(new_n1046_), .B(new_n1921_), .ZN(new_n1922_));
  INV_X1     g1280(.I(new_n1922_), .ZN(new_n1923_));
  NOR2_X1    g1281(.A1(new_n1923_), .A2(new_n1920_), .ZN(new_n1924_));
  NOR2_X1    g1282(.A1(new_n1918_), .A2(new_n1924_), .ZN(new_n1925_));
  INV_X1     g1283(.I(new_n1925_), .ZN(new_n1926_));
  AOI21_X1   g1284(.A1(new_n1903_), .A2(new_n1906_), .B(new_n1926_), .ZN(new_n1927_));
  AOI21_X1   g1285(.A1(new_n1927_), .A2(new_n1901_), .B(new_n1869_), .ZN(new_n1928_));
  INV_X1     g1286(.I(new_n1928_), .ZN(new_n1929_));
  NOR2_X1    g1287(.A1(new_n1046_), .A2(\in3[31] ), .ZN(new_n1930_));
  AOI21_X1   g1288(.A1(new_n714_), .A2(new_n1046_), .B(new_n1930_), .ZN(new_n1931_));
  OAI21_X1   g1289(.A1(new_n1877_), .A2(new_n1929_), .B(new_n1931_), .ZN(new_n1932_));
  AOI21_X1   g1290(.A1(new_n1871_), .A2(new_n1876_), .B(new_n1932_), .ZN(new_n1933_));
  NOR2_X1    g1291(.A1(new_n1046_), .A2(\in3[46] ), .ZN(new_n1934_));
  AOI21_X1   g1292(.A1(new_n661_), .A2(new_n1046_), .B(new_n1934_), .ZN(new_n1935_));
  INV_X1     g1293(.I(new_n1935_), .ZN(new_n1936_));
  NOR2_X1    g1294(.A1(new_n1568_), .A2(\in1[46] ), .ZN(new_n1937_));
  AOI21_X1   g1295(.A1(new_n1064_), .A2(new_n1568_), .B(new_n1937_), .ZN(new_n1938_));
  NOR2_X1    g1296(.A1(new_n1046_), .A2(\in3[47] ), .ZN(new_n1939_));
  AOI21_X1   g1297(.A1(new_n659_), .A2(new_n1046_), .B(new_n1939_), .ZN(new_n1940_));
  INV_X1     g1298(.I(new_n1940_), .ZN(new_n1941_));
  NOR2_X1    g1299(.A1(new_n1494_), .A2(\in0[47] ), .ZN(new_n1942_));
  AOI21_X1   g1300(.A1(new_n1086_), .A2(new_n1494_), .B(new_n1942_), .ZN(new_n1943_));
  OAI22_X1   g1301(.A1(new_n1936_), .A2(new_n1938_), .B1(new_n1941_), .B2(new_n1943_), .ZN(new_n1944_));
  INV_X1     g1302(.I(\in1[44] ), .ZN(new_n1945_));
  NOR2_X1    g1303(.A1(new_n1494_), .A2(\in0[44] ), .ZN(new_n1946_));
  AOI21_X1   g1304(.A1(new_n1945_), .A2(new_n1494_), .B(new_n1946_), .ZN(new_n1947_));
  INV_X1     g1305(.I(new_n1947_), .ZN(new_n1948_));
  NOR2_X1    g1306(.A1(new_n1046_), .A2(\in3[44] ), .ZN(new_n1949_));
  AOI21_X1   g1307(.A1(new_n665_), .A2(new_n1046_), .B(new_n1949_), .ZN(new_n1950_));
  NOR2_X1    g1308(.A1(new_n1948_), .A2(new_n1950_), .ZN(new_n1951_));
  NOR2_X1    g1309(.A1(new_n1046_), .A2(\in3[45] ), .ZN(new_n1952_));
  AOI21_X1   g1310(.A1(new_n663_), .A2(new_n1046_), .B(new_n1952_), .ZN(new_n1953_));
  NOR2_X1    g1311(.A1(new_n1494_), .A2(\in0[45] ), .ZN(new_n1954_));
  AOI21_X1   g1312(.A1(new_n1089_), .A2(new_n1494_), .B(new_n1954_), .ZN(new_n1955_));
  INV_X1     g1313(.I(new_n1953_), .ZN(new_n1956_));
  NAND2_X1   g1314(.A1(new_n1956_), .A2(new_n1955_), .ZN(new_n1957_));
  NOR2_X1    g1315(.A1(new_n1956_), .A2(new_n1955_), .ZN(new_n1958_));
  INV_X1     g1316(.I(new_n1958_), .ZN(new_n1959_));
  AOI22_X1   g1317(.A1(new_n1959_), .A2(new_n1957_), .B1(new_n1951_), .B2(new_n1953_), .ZN(new_n1960_));
  NAND2_X1   g1318(.A1(new_n1960_), .A2(new_n1944_), .ZN(new_n1961_));
  INV_X1     g1319(.I(new_n1950_), .ZN(new_n1962_));
  NOR4_X1    g1320(.A1(new_n1944_), .A2(new_n1947_), .A3(new_n1962_), .A4(new_n1958_), .ZN(new_n1963_));
  INV_X1     g1321(.I(new_n1963_), .ZN(new_n1964_));
  NOR2_X1    g1322(.A1(new_n1494_), .A2(\in0[43] ), .ZN(new_n1965_));
  AOI21_X1   g1323(.A1(new_n1073_), .A2(new_n1494_), .B(new_n1965_), .ZN(new_n1966_));
  NOR2_X1    g1324(.A1(new_n1046_), .A2(\in3[43] ), .ZN(new_n1967_));
  AOI21_X1   g1325(.A1(new_n668_), .A2(new_n1046_), .B(new_n1967_), .ZN(new_n1968_));
  INV_X1     g1326(.I(new_n1968_), .ZN(new_n1969_));
  NAND2_X1   g1327(.A1(new_n1969_), .A2(new_n1966_), .ZN(new_n1970_));
  NOR2_X1    g1328(.A1(new_n1494_), .A2(\in0[42] ), .ZN(new_n1971_));
  AOI21_X1   g1329(.A1(new_n1074_), .A2(new_n1494_), .B(new_n1971_), .ZN(new_n1972_));
  INV_X1     g1330(.I(new_n1972_), .ZN(new_n1973_));
  NOR2_X1    g1331(.A1(new_n1046_), .A2(\in3[42] ), .ZN(new_n1974_));
  AOI21_X1   g1332(.A1(new_n669_), .A2(new_n1046_), .B(new_n1974_), .ZN(new_n1975_));
  NOR2_X1    g1333(.A1(new_n1969_), .A2(new_n1966_), .ZN(new_n1976_));
  AOI21_X1   g1334(.A1(new_n1973_), .A2(new_n1975_), .B(new_n1976_), .ZN(new_n1977_));
  NOR2_X1    g1335(.A1(new_n1046_), .A2(\in3[41] ), .ZN(new_n1978_));
  AOI21_X1   g1336(.A1(new_n674_), .A2(new_n1046_), .B(new_n1978_), .ZN(new_n1979_));
  INV_X1     g1337(.I(new_n1979_), .ZN(new_n1980_));
  NOR2_X1    g1338(.A1(new_n1494_), .A2(\in0[41] ), .ZN(new_n1981_));
  AOI21_X1   g1339(.A1(new_n1081_), .A2(new_n1494_), .B(new_n1981_), .ZN(new_n1982_));
  NOR2_X1    g1340(.A1(new_n1980_), .A2(new_n1982_), .ZN(new_n1983_));
  INV_X1     g1341(.I(new_n1983_), .ZN(new_n1984_));
  NOR2_X1    g1342(.A1(new_n1494_), .A2(\in0[40] ), .ZN(new_n1985_));
  AOI21_X1   g1343(.A1(new_n1080_), .A2(new_n1494_), .B(new_n1985_), .ZN(new_n1986_));
  NOR2_X1    g1344(.A1(new_n1046_), .A2(\in3[40] ), .ZN(new_n1987_));
  AOI21_X1   g1345(.A1(new_n710_), .A2(new_n1046_), .B(new_n1987_), .ZN(new_n1988_));
  OAI21_X1   g1346(.A1(new_n1973_), .A2(new_n1975_), .B(new_n1984_), .ZN(new_n1989_));
  OAI21_X1   g1347(.A1(new_n1989_), .A2(new_n1977_), .B(new_n1970_), .ZN(new_n1990_));
  XNOR2_X1   g1348(.A1(new_n1943_), .A2(new_n1940_), .ZN(new_n1991_));
  AOI21_X1   g1349(.A1(new_n1991_), .A2(new_n1938_), .B(new_n1936_), .ZN(new_n1992_));
  NAND2_X1   g1350(.A1(new_n1941_), .A2(new_n1943_), .ZN(new_n1993_));
  XOR2_X1    g1351(.A1(new_n1992_), .A2(new_n1993_), .Z(new_n1994_));
  NAND4_X1   g1352(.A1(new_n1994_), .A2(new_n1961_), .A3(new_n1964_), .A4(new_n1990_), .ZN(new_n1995_));
  XNOR2_X1   g1353(.A1(new_n1911_), .A2(new_n1908_), .ZN(new_n1996_));
  AOI21_X1   g1354(.A1(new_n1996_), .A2(new_n1920_), .B(new_n1923_), .ZN(new_n1997_));
  OAI21_X1   g1355(.A1(new_n1912_), .A2(new_n1996_), .B(new_n1997_), .ZN(new_n1998_));
  OR3_X2     g1356(.A1(new_n1997_), .A2(new_n1912_), .A3(new_n1996_), .Z(new_n1999_));
  INV_X1     g1357(.I(new_n1903_), .ZN(new_n2000_));
  OAI22_X1   g1358(.A1(new_n2000_), .A2(new_n1905_), .B1(new_n1917_), .B2(new_n1914_), .ZN(new_n2001_));
  NOR3_X1    g1359(.A1(new_n1926_), .A2(new_n1901_), .A3(new_n2001_), .ZN(new_n2002_));
  NAND3_X1   g1360(.A1(new_n1999_), .A2(new_n1998_), .A3(new_n2002_), .ZN(new_n2003_));
  INV_X1     g1361(.I(new_n1888_), .ZN(new_n2004_));
  XNOR2_X1   g1362(.A1(new_n1887_), .A2(new_n1884_), .ZN(new_n2005_));
  AOI21_X1   g1363(.A1(new_n2005_), .A2(new_n1882_), .B(new_n1880_), .ZN(new_n2006_));
  NAND2_X1   g1364(.A1(new_n1885_), .A2(new_n1887_), .ZN(new_n2007_));
  NOR2_X1    g1365(.A1(new_n2006_), .A2(new_n2007_), .ZN(new_n2008_));
  INV_X1     g1366(.I(new_n1988_), .ZN(new_n2009_));
  NOR2_X1    g1367(.A1(new_n2009_), .A2(new_n1986_), .ZN(new_n2010_));
  NOR2_X1    g1368(.A1(new_n1983_), .A2(new_n2010_), .ZN(new_n2011_));
  NOR3_X1    g1369(.A1(new_n1964_), .A2(new_n1977_), .A3(new_n2011_), .ZN(new_n2012_));
  NOR3_X1    g1370(.A1(new_n2012_), .A2(new_n2004_), .A3(new_n2008_), .ZN(new_n2013_));
  XOR2_X1    g1371(.A1(new_n1893_), .A2(new_n1890_), .Z(new_n2014_));
  INV_X1     g1372(.I(new_n1900_), .ZN(new_n2015_));
  OAI21_X1   g1373(.A1(new_n2014_), .A2(new_n2015_), .B(new_n1896_), .ZN(new_n2016_));
  AOI21_X1   g1374(.A1(new_n1893_), .A2(new_n2014_), .B(new_n2016_), .ZN(new_n2017_));
  AND2_X2    g1375(.A1(new_n2006_), .A2(new_n2007_), .Z(new_n2018_));
  AND3_X2    g1376(.A1(new_n1891_), .A2(new_n1897_), .A3(new_n1893_), .Z(new_n2019_));
  NOR3_X1    g1377(.A1(new_n2018_), .A2(new_n2017_), .A3(new_n2019_), .ZN(new_n2020_));
  NAND4_X1   g1378(.A1(new_n1995_), .A2(new_n2003_), .A3(new_n2013_), .A4(new_n2020_), .ZN(new_n2021_));
  NOR2_X1    g1379(.A1(new_n1046_), .A2(\in3[50] ), .ZN(new_n2022_));
  AOI21_X1   g1380(.A1(new_n755_), .A2(new_n1046_), .B(new_n2022_), .ZN(new_n2023_));
  NOR2_X1    g1381(.A1(new_n1494_), .A2(\in0[50] ), .ZN(new_n2024_));
  AOI21_X1   g1382(.A1(new_n1138_), .A2(new_n1494_), .B(new_n2024_), .ZN(new_n2025_));
  NOR2_X1    g1383(.A1(new_n1046_), .A2(\in3[51] ), .ZN(new_n2026_));
  AOI21_X1   g1384(.A1(new_n743_), .A2(new_n1046_), .B(new_n2026_), .ZN(new_n2027_));
  INV_X1     g1385(.I(new_n2027_), .ZN(new_n2028_));
  NOR2_X1    g1386(.A1(new_n1494_), .A2(\in0[51] ), .ZN(new_n2029_));
  AOI21_X1   g1387(.A1(new_n1139_), .A2(new_n1494_), .B(new_n2029_), .ZN(new_n2030_));
  NOR2_X1    g1388(.A1(new_n2028_), .A2(new_n2030_), .ZN(new_n2031_));
  INV_X1     g1389(.I(new_n2031_), .ZN(new_n2032_));
  NAND2_X1   g1390(.A1(new_n2028_), .A2(new_n2030_), .ZN(new_n2033_));
  NAND3_X1   g1391(.A1(new_n2032_), .A2(new_n2025_), .A3(new_n2033_), .ZN(new_n2034_));
  NAND2_X1   g1392(.A1(new_n2034_), .A2(new_n2023_), .ZN(new_n2035_));
  NAND2_X1   g1393(.A1(new_n2028_), .A2(new_n2030_), .ZN(new_n2036_));
  XNOR2_X1   g1394(.A1(new_n2035_), .A2(new_n2036_), .ZN(new_n2037_));
  INV_X1     g1395(.I(new_n2037_), .ZN(new_n2038_));
  INV_X1     g1396(.I(new_n2023_), .ZN(new_n2039_));
  NOR2_X1    g1397(.A1(new_n1046_), .A2(\in3[49] ), .ZN(new_n2040_));
  AOI21_X1   g1398(.A1(new_n740_), .A2(new_n1046_), .B(new_n2040_), .ZN(new_n2041_));
  INV_X1     g1399(.I(new_n2041_), .ZN(new_n2042_));
  NOR2_X1    g1400(.A1(new_n1494_), .A2(\in0[49] ), .ZN(new_n2043_));
  AOI21_X1   g1401(.A1(new_n1141_), .A2(new_n1494_), .B(new_n2043_), .ZN(new_n2044_));
  NOR2_X1    g1402(.A1(new_n2042_), .A2(new_n2044_), .ZN(new_n2045_));
  OAI22_X1   g1403(.A1(new_n2031_), .A2(new_n2045_), .B1(new_n2039_), .B2(new_n2025_), .ZN(new_n2046_));
  NAND2_X1   g1404(.A1(new_n2042_), .A2(new_n2044_), .ZN(new_n2047_));
  NOR2_X1    g1405(.A1(new_n1494_), .A2(\in0[48] ), .ZN(new_n2048_));
  AOI21_X1   g1406(.A1(new_n1466_), .A2(new_n1494_), .B(new_n2048_), .ZN(new_n2049_));
  NOR2_X1    g1407(.A1(new_n1046_), .A2(\in3[48] ), .ZN(new_n2050_));
  AOI21_X1   g1408(.A1(new_n757_), .A2(new_n1046_), .B(new_n2050_), .ZN(new_n2051_));
  INV_X1     g1409(.I(new_n2051_), .ZN(new_n2052_));
  NAND2_X1   g1410(.A1(new_n2052_), .A2(new_n2049_), .ZN(new_n2053_));
  AOI21_X1   g1411(.A1(new_n2047_), .A2(new_n2053_), .B(new_n2046_), .ZN(new_n2054_));
  NOR2_X1    g1412(.A1(new_n1494_), .A2(\in0[54] ), .ZN(new_n2055_));
  AOI21_X1   g1413(.A1(new_n1150_), .A2(new_n1494_), .B(new_n2055_), .ZN(new_n2056_));
  INV_X1     g1414(.I(new_n2056_), .ZN(new_n2057_));
  NOR2_X1    g1415(.A1(new_n1046_), .A2(\in3[54] ), .ZN(new_n2058_));
  AOI21_X1   g1416(.A1(new_n726_), .A2(new_n1046_), .B(new_n2058_), .ZN(new_n2059_));
  NOR2_X1    g1417(.A1(new_n1494_), .A2(\in0[55] ), .ZN(new_n2060_));
  AOI21_X1   g1418(.A1(new_n1151_), .A2(new_n1494_), .B(new_n2060_), .ZN(new_n2061_));
  INV_X1     g1419(.I(new_n2061_), .ZN(new_n2062_));
  NOR2_X1    g1420(.A1(new_n1046_), .A2(\in3[55] ), .ZN(new_n2063_));
  AOI21_X1   g1421(.A1(new_n727_), .A2(new_n1046_), .B(new_n2063_), .ZN(new_n2064_));
  AOI22_X1   g1422(.A1(new_n2057_), .A2(new_n2059_), .B1(new_n2062_), .B2(new_n2064_), .ZN(new_n2065_));
  INV_X1     g1423(.I(new_n2065_), .ZN(new_n2066_));
  INV_X1     g1424(.I(new_n2059_), .ZN(new_n2067_));
  NOR2_X1    g1425(.A1(new_n1046_), .A2(\in3[53] ), .ZN(new_n2068_));
  AOI21_X1   g1426(.A1(new_n729_), .A2(new_n1046_), .B(new_n2068_), .ZN(new_n2069_));
  INV_X1     g1427(.I(new_n2069_), .ZN(new_n2070_));
  NOR2_X1    g1428(.A1(new_n1494_), .A2(\in0[53] ), .ZN(new_n2071_));
  AOI21_X1   g1429(.A1(new_n1153_), .A2(new_n1494_), .B(new_n2071_), .ZN(new_n2072_));
  NOR2_X1    g1430(.A1(new_n2070_), .A2(new_n2072_), .ZN(new_n2073_));
  NOR2_X1    g1431(.A1(new_n1494_), .A2(\in0[52] ), .ZN(new_n2074_));
  AOI21_X1   g1432(.A1(new_n1155_), .A2(new_n1494_), .B(new_n2074_), .ZN(new_n2075_));
  NOR2_X1    g1433(.A1(new_n1046_), .A2(\in3[52] ), .ZN(new_n2076_));
  AOI21_X1   g1434(.A1(new_n731_), .A2(new_n1046_), .B(new_n2076_), .ZN(new_n2077_));
  AOI21_X1   g1435(.A1(new_n2056_), .A2(new_n2067_), .B(new_n2073_), .ZN(new_n2078_));
  NAND2_X1   g1436(.A1(new_n2066_), .A2(new_n2078_), .ZN(new_n2079_));
  INV_X1     g1437(.I(new_n2079_), .ZN(new_n2080_));
  NOR2_X1    g1438(.A1(new_n2062_), .A2(new_n2064_), .ZN(new_n2081_));
  INV_X1     g1439(.I(new_n2073_), .ZN(new_n2082_));
  INV_X1     g1440(.I(new_n2077_), .ZN(new_n2083_));
  NOR2_X1    g1441(.A1(new_n2083_), .A2(new_n2075_), .ZN(new_n2084_));
  NOR3_X1    g1442(.A1(new_n2066_), .A2(new_n2082_), .A3(new_n2084_), .ZN(new_n2085_));
  NOR4_X1    g1443(.A1(new_n2080_), .A2(new_n2054_), .A3(new_n2081_), .A4(new_n2085_), .ZN(new_n2086_));
  NAND2_X1   g1444(.A1(new_n2038_), .A2(new_n2086_), .ZN(new_n2087_));
  NOR2_X1    g1445(.A1(new_n1046_), .A2(\in3[62] ), .ZN(new_n2088_));
  AOI21_X1   g1446(.A1(new_n786_), .A2(new_n1046_), .B(new_n2088_), .ZN(new_n2089_));
  INV_X1     g1447(.I(new_n2089_), .ZN(new_n2090_));
  NOR2_X1    g1448(.A1(new_n1568_), .A2(\in1[62] ), .ZN(new_n2091_));
  AOI21_X1   g1449(.A1(new_n1167_), .A2(new_n1568_), .B(new_n2091_), .ZN(new_n2092_));
  NOR2_X1    g1450(.A1(new_n1046_), .A2(\in3[63] ), .ZN(new_n2093_));
  AOI21_X1   g1451(.A1(new_n784_), .A2(new_n1046_), .B(new_n2093_), .ZN(new_n2094_));
  INV_X1     g1452(.I(new_n2094_), .ZN(new_n2095_));
  NOR2_X1    g1453(.A1(new_n1494_), .A2(\in0[63] ), .ZN(new_n2096_));
  AOI21_X1   g1454(.A1(new_n1212_), .A2(new_n1494_), .B(new_n2096_), .ZN(new_n2097_));
  OAI22_X1   g1455(.A1(new_n2090_), .A2(new_n2092_), .B1(new_n2095_), .B2(new_n2097_), .ZN(new_n2098_));
  NOR2_X1    g1456(.A1(new_n1046_), .A2(\in3[61] ), .ZN(new_n2099_));
  AOI21_X1   g1457(.A1(new_n788_), .A2(new_n1046_), .B(new_n2099_), .ZN(new_n2100_));
  INV_X1     g1458(.I(new_n2100_), .ZN(new_n2101_));
  NOR2_X1    g1459(.A1(new_n1494_), .A2(\in0[61] ), .ZN(new_n2102_));
  AOI21_X1   g1460(.A1(new_n1209_), .A2(new_n1494_), .B(new_n2102_), .ZN(new_n2103_));
  NOR2_X1    g1461(.A1(new_n2101_), .A2(new_n2103_), .ZN(new_n2104_));
  NOR2_X1    g1462(.A1(new_n1046_), .A2(\in3[60] ), .ZN(new_n2105_));
  AOI21_X1   g1463(.A1(new_n790_), .A2(new_n1046_), .B(new_n2105_), .ZN(new_n2106_));
  INV_X1     g1464(.I(new_n2106_), .ZN(new_n2107_));
  NOR2_X1    g1465(.A1(new_n1568_), .A2(\in1[60] ), .ZN(new_n2108_));
  AOI21_X1   g1466(.A1(new_n1172_), .A2(new_n1568_), .B(new_n2108_), .ZN(new_n2109_));
  NOR4_X1    g1467(.A1(new_n2098_), .A2(new_n2104_), .A3(new_n2107_), .A4(new_n2109_), .ZN(new_n2110_));
  INV_X1     g1468(.I(new_n2110_), .ZN(new_n2111_));
  NOR2_X1    g1469(.A1(new_n1046_), .A2(\in3[56] ), .ZN(new_n2112_));
  AOI21_X1   g1470(.A1(new_n798_), .A2(new_n1046_), .B(new_n2112_), .ZN(new_n2113_));
  INV_X1     g1471(.I(new_n2113_), .ZN(new_n2114_));
  NOR2_X1    g1472(.A1(new_n1494_), .A2(\in0[56] ), .ZN(new_n2115_));
  AOI21_X1   g1473(.A1(new_n1176_), .A2(new_n1494_), .B(new_n2115_), .ZN(new_n2116_));
  NOR2_X1    g1474(.A1(new_n2114_), .A2(new_n2116_), .ZN(new_n2117_));
  NOR2_X1    g1475(.A1(new_n1046_), .A2(\in3[57] ), .ZN(new_n2118_));
  AOI21_X1   g1476(.A1(new_n796_), .A2(new_n1046_), .B(new_n2118_), .ZN(new_n2119_));
  INV_X1     g1477(.I(new_n2119_), .ZN(new_n2120_));
  NOR2_X1    g1478(.A1(new_n1494_), .A2(\in0[57] ), .ZN(new_n2121_));
  AOI21_X1   g1479(.A1(new_n1177_), .A2(new_n1494_), .B(new_n2121_), .ZN(new_n2122_));
  NOR2_X1    g1480(.A1(new_n2120_), .A2(new_n2122_), .ZN(new_n2123_));
  NOR2_X1    g1481(.A1(new_n2117_), .A2(new_n2123_), .ZN(new_n2124_));
  NOR2_X1    g1482(.A1(new_n1046_), .A2(\in3[58] ), .ZN(new_n2125_));
  AOI21_X1   g1483(.A1(new_n793_), .A2(new_n1046_), .B(new_n2125_), .ZN(new_n2126_));
  NOR2_X1    g1484(.A1(new_n1494_), .A2(\in0[58] ), .ZN(new_n2127_));
  AOI21_X1   g1485(.A1(new_n1179_), .A2(new_n1494_), .B(new_n2127_), .ZN(new_n2128_));
  INV_X1     g1486(.I(new_n2128_), .ZN(new_n2129_));
  NOR2_X1    g1487(.A1(new_n1046_), .A2(\in3[59] ), .ZN(new_n2130_));
  AOI21_X1   g1488(.A1(new_n794_), .A2(new_n1046_), .B(new_n2130_), .ZN(new_n2131_));
  NOR2_X1    g1489(.A1(new_n1494_), .A2(\in0[59] ), .ZN(new_n2132_));
  AOI21_X1   g1490(.A1(new_n1180_), .A2(new_n1494_), .B(new_n2132_), .ZN(new_n2133_));
  INV_X1     g1491(.I(new_n2133_), .ZN(new_n2134_));
  AOI22_X1   g1492(.A1(new_n2126_), .A2(new_n2129_), .B1(new_n2134_), .B2(new_n2131_), .ZN(new_n2135_));
  NOR3_X1    g1493(.A1(new_n2111_), .A2(new_n2124_), .A3(new_n2135_), .ZN(new_n2136_));
  NAND2_X1   g1494(.A1(new_n2085_), .A2(new_n2053_), .ZN(new_n2137_));
  NOR3_X1    g1495(.A1(new_n2136_), .A2(new_n2046_), .A3(new_n2137_), .ZN(new_n2138_));
  AND2_X2    g1496(.A1(new_n2087_), .A2(new_n2138_), .Z(new_n2139_));
  OAI21_X1   g1497(.A1(new_n1933_), .A2(new_n2021_), .B(new_n2139_), .ZN(new_n2140_));
  NOR2_X1    g1498(.A1(new_n1494_), .A2(\in0[66] ), .ZN(new_n2141_));
  AOI21_X1   g1499(.A1(new_n1205_), .A2(new_n1494_), .B(new_n2141_), .ZN(new_n2142_));
  NOR2_X1    g1500(.A1(new_n1554_), .A2(\in2[66] ), .ZN(new_n2143_));
  AOI21_X1   g1501(.A1(new_n807_), .A2(new_n1554_), .B(new_n2143_), .ZN(new_n2144_));
  INV_X1     g1502(.I(new_n2144_), .ZN(new_n2145_));
  NOR2_X1    g1503(.A1(new_n1494_), .A2(\in0[67] ), .ZN(new_n2146_));
  AOI21_X1   g1504(.A1(new_n1206_), .A2(new_n1494_), .B(new_n2146_), .ZN(new_n2147_));
  NOR2_X1    g1505(.A1(new_n1554_), .A2(\in2[67] ), .ZN(new_n2148_));
  AOI21_X1   g1506(.A1(new_n810_), .A2(new_n1554_), .B(new_n2148_), .ZN(new_n2149_));
  INV_X1     g1507(.I(new_n2149_), .ZN(new_n2150_));
  OAI22_X1   g1508(.A1(new_n2142_), .A2(new_n2145_), .B1(new_n2150_), .B2(new_n2147_), .ZN(new_n2151_));
  NOR2_X1    g1509(.A1(new_n1554_), .A2(\in2[65] ), .ZN(new_n2152_));
  AOI21_X1   g1510(.A1(new_n803_), .A2(new_n1554_), .B(new_n2152_), .ZN(new_n2153_));
  INV_X1     g1511(.I(new_n2153_), .ZN(new_n2154_));
  NOR2_X1    g1512(.A1(new_n1568_), .A2(\in1[65] ), .ZN(new_n2155_));
  AOI21_X1   g1513(.A1(new_n1197_), .A2(new_n1568_), .B(new_n2155_), .ZN(new_n2156_));
  NOR2_X1    g1514(.A1(new_n2154_), .A2(new_n2156_), .ZN(new_n2157_));
  NOR2_X1    g1515(.A1(new_n1494_), .A2(\in0[64] ), .ZN(new_n2158_));
  AOI21_X1   g1516(.A1(new_n1196_), .A2(new_n1494_), .B(new_n2158_), .ZN(new_n2159_));
  NOR2_X1    g1517(.A1(new_n1046_), .A2(\in3[64] ), .ZN(new_n2160_));
  AOI21_X1   g1518(.A1(new_n815_), .A2(new_n1046_), .B(new_n2160_), .ZN(new_n2161_));
  AOI21_X1   g1519(.A1(new_n2142_), .A2(new_n2145_), .B(new_n2157_), .ZN(new_n2162_));
  NAND2_X1   g1520(.A1(new_n2162_), .A2(new_n2151_), .ZN(new_n2163_));
  NAND2_X1   g1521(.A1(new_n2150_), .A2(new_n2147_), .ZN(new_n2164_));
  INV_X1     g1522(.I(new_n2161_), .ZN(new_n2165_));
  OAI21_X1   g1523(.A1(new_n2159_), .A2(new_n2165_), .B(new_n2157_), .ZN(new_n2166_));
  OR2_X2     g1524(.A1(new_n2166_), .A2(new_n2151_), .Z(new_n2167_));
  NAND4_X1   g1525(.A1(new_n2167_), .A2(new_n2111_), .A3(new_n2163_), .A4(new_n2164_), .ZN(new_n2168_));
  INV_X1     g1526(.I(new_n2098_), .ZN(new_n2169_));
  NAND2_X1   g1527(.A1(new_n2109_), .A2(new_n2107_), .ZN(new_n2170_));
  INV_X1     g1528(.I(new_n2103_), .ZN(new_n2171_));
  NOR2_X1    g1529(.A1(new_n2171_), .A2(new_n2100_), .ZN(new_n2172_));
  OAI22_X1   g1530(.A1(new_n2101_), .A2(new_n2170_), .B1(new_n2172_), .B2(new_n2104_), .ZN(new_n2173_));
  XNOR2_X1   g1531(.A1(new_n2097_), .A2(new_n2094_), .ZN(new_n2174_));
  AOI21_X1   g1532(.A1(new_n2174_), .A2(new_n2092_), .B(new_n2090_), .ZN(new_n2175_));
  NAND2_X1   g1533(.A1(new_n2095_), .A2(new_n2097_), .ZN(new_n2176_));
  OAI22_X1   g1534(.A1(new_n2175_), .A2(new_n2176_), .B1(new_n2173_), .B2(new_n2169_), .ZN(new_n2177_));
  NAND2_X1   g1535(.A1(new_n2175_), .A2(new_n2176_), .ZN(new_n2178_));
  NOR2_X1    g1536(.A1(new_n2134_), .A2(new_n2131_), .ZN(new_n2179_));
  INV_X1     g1537(.I(new_n2123_), .ZN(new_n2180_));
  AOI21_X1   g1538(.A1(new_n2114_), .A2(new_n2116_), .B(new_n2180_), .ZN(new_n2181_));
  NOR2_X1    g1539(.A1(new_n2129_), .A2(new_n2126_), .ZN(new_n2182_));
  NOR4_X1    g1540(.A1(new_n2181_), .A2(new_n2123_), .A3(new_n2135_), .A4(new_n2182_), .ZN(new_n2183_));
  OAI21_X1   g1541(.A1(new_n2183_), .A2(new_n2179_), .B(new_n2178_), .ZN(new_n2184_));
  NOR3_X1    g1542(.A1(new_n2184_), .A2(new_n2168_), .A3(new_n2177_), .ZN(new_n2185_));
  INV_X1     g1543(.I(\in2[70] ), .ZN(new_n2186_));
  NOR2_X1    g1544(.A1(new_n1046_), .A2(\in3[70] ), .ZN(new_n2187_));
  AOI21_X1   g1545(.A1(new_n2186_), .A2(new_n1046_), .B(new_n2187_), .ZN(new_n2188_));
  NOR2_X1    g1546(.A1(new_n1494_), .A2(\in0[70] ), .ZN(new_n2189_));
  AOI21_X1   g1547(.A1(new_n1222_), .A2(new_n1494_), .B(new_n2189_), .ZN(new_n2190_));
  NOR2_X1    g1548(.A1(new_n1046_), .A2(\in3[71] ), .ZN(new_n2191_));
  AOI21_X1   g1549(.A1(new_n826_), .A2(new_n1046_), .B(new_n2191_), .ZN(new_n2192_));
  INV_X1     g1550(.I(new_n2192_), .ZN(new_n2193_));
  NOR2_X1    g1551(.A1(new_n1494_), .A2(\in0[71] ), .ZN(new_n2194_));
  AOI21_X1   g1552(.A1(new_n1223_), .A2(new_n1494_), .B(new_n2194_), .ZN(new_n2195_));
  NOR2_X1    g1553(.A1(new_n2193_), .A2(new_n2195_), .ZN(new_n2196_));
  INV_X1     g1554(.I(new_n2196_), .ZN(new_n2197_));
  NAND2_X1   g1555(.A1(new_n2193_), .A2(new_n2195_), .ZN(new_n2198_));
  NAND3_X1   g1556(.A1(new_n2197_), .A2(new_n2190_), .A3(new_n2198_), .ZN(new_n2199_));
  NAND2_X1   g1557(.A1(new_n2199_), .A2(new_n2188_), .ZN(new_n2200_));
  NAND2_X1   g1558(.A1(new_n2193_), .A2(new_n2195_), .ZN(new_n2201_));
  XNOR2_X1   g1559(.A1(new_n2200_), .A2(new_n2201_), .ZN(new_n2202_));
  NOR2_X1    g1560(.A1(new_n1554_), .A2(\in2[68] ), .ZN(new_n2203_));
  AOI21_X1   g1561(.A1(new_n829_), .A2(new_n1554_), .B(new_n2203_), .ZN(new_n2204_));
  INV_X1     g1562(.I(new_n2204_), .ZN(new_n2205_));
  NOR2_X1    g1563(.A1(new_n1494_), .A2(\in0[68] ), .ZN(new_n2206_));
  AOI21_X1   g1564(.A1(new_n1229_), .A2(new_n1494_), .B(new_n2206_), .ZN(new_n2207_));
  NOR2_X1    g1565(.A1(new_n1494_), .A2(\in0[69] ), .ZN(new_n2208_));
  AOI21_X1   g1566(.A1(new_n1239_), .A2(new_n1494_), .B(new_n2208_), .ZN(new_n2209_));
  INV_X1     g1567(.I(new_n2209_), .ZN(new_n2210_));
  NOR2_X1    g1568(.A1(new_n1046_), .A2(\in3[69] ), .ZN(new_n2211_));
  AOI21_X1   g1569(.A1(new_n828_), .A2(new_n1046_), .B(new_n2211_), .ZN(new_n2212_));
  NOR2_X1    g1570(.A1(new_n2210_), .A2(new_n2212_), .ZN(new_n2213_));
  INV_X1     g1571(.I(new_n2212_), .ZN(new_n2214_));
  NOR2_X1    g1572(.A1(new_n2214_), .A2(new_n2209_), .ZN(new_n2215_));
  NOR2_X1    g1573(.A1(new_n2213_), .A2(new_n2215_), .ZN(new_n2216_));
  AOI21_X1   g1574(.A1(new_n2216_), .A2(new_n2207_), .B(new_n2205_), .ZN(new_n2217_));
  INV_X1     g1575(.I(new_n2217_), .ZN(new_n2218_));
  NOR2_X1    g1576(.A1(new_n2210_), .A2(new_n2212_), .ZN(new_n2219_));
  NOR2_X1    g1577(.A1(new_n2218_), .A2(new_n2219_), .ZN(new_n2220_));
  NAND2_X1   g1578(.A1(new_n2218_), .A2(new_n2219_), .ZN(new_n2221_));
  INV_X1     g1579(.I(new_n2188_), .ZN(new_n2222_));
  OAI21_X1   g1580(.A1(new_n2222_), .A2(new_n2190_), .B(new_n2197_), .ZN(new_n2223_));
  NAND2_X1   g1581(.A1(new_n2221_), .A2(new_n2223_), .ZN(new_n2224_));
  NOR2_X1    g1582(.A1(new_n2224_), .A2(new_n2220_), .ZN(new_n2225_));
  NOR2_X1    g1583(.A1(new_n1554_), .A2(\in2[74] ), .ZN(new_n2226_));
  AOI21_X1   g1584(.A1(new_n833_), .A2(new_n1554_), .B(new_n2226_), .ZN(new_n2227_));
  INV_X1     g1585(.I(new_n2227_), .ZN(new_n2228_));
  NOR2_X1    g1586(.A1(new_n1494_), .A2(\in0[74] ), .ZN(new_n2229_));
  AOI21_X1   g1587(.A1(new_n1233_), .A2(new_n1494_), .B(new_n2229_), .ZN(new_n2230_));
  NOR2_X1    g1588(.A1(new_n1554_), .A2(\in2[75] ), .ZN(new_n2231_));
  AOI21_X1   g1589(.A1(new_n834_), .A2(new_n1554_), .B(new_n2231_), .ZN(new_n2232_));
  INV_X1     g1590(.I(new_n2232_), .ZN(new_n2233_));
  NOR2_X1    g1591(.A1(new_n1494_), .A2(\in0[75] ), .ZN(new_n2234_));
  AOI21_X1   g1592(.A1(new_n1234_), .A2(new_n1494_), .B(new_n2234_), .ZN(new_n2235_));
  OAI22_X1   g1593(.A1(new_n2228_), .A2(new_n2230_), .B1(new_n2233_), .B2(new_n2235_), .ZN(new_n2236_));
  NOR2_X1    g1594(.A1(new_n1046_), .A2(\in3[72] ), .ZN(new_n2237_));
  AOI21_X1   g1595(.A1(new_n832_), .A2(new_n1046_), .B(new_n2237_), .ZN(new_n2238_));
  INV_X1     g1596(.I(new_n2238_), .ZN(new_n2239_));
  NOR2_X1    g1597(.A1(new_n1494_), .A2(\in0[72] ), .ZN(new_n2240_));
  AOI21_X1   g1598(.A1(new_n1245_), .A2(new_n1494_), .B(new_n2240_), .ZN(new_n2241_));
  NOR2_X1    g1599(.A1(new_n2239_), .A2(new_n2241_), .ZN(new_n2242_));
  NOR2_X1    g1600(.A1(new_n1046_), .A2(\in3[73] ), .ZN(new_n2243_));
  AOI21_X1   g1601(.A1(new_n846_), .A2(new_n1046_), .B(new_n2243_), .ZN(new_n2244_));
  INV_X1     g1602(.I(new_n2244_), .ZN(new_n2245_));
  NOR2_X1    g1603(.A1(new_n1494_), .A2(\in0[73] ), .ZN(new_n2246_));
  AOI21_X1   g1604(.A1(new_n1236_), .A2(new_n1494_), .B(new_n2246_), .ZN(new_n2247_));
  NOR2_X1    g1605(.A1(new_n2245_), .A2(new_n2247_), .ZN(new_n2248_));
  INV_X1     g1606(.I(new_n2248_), .ZN(new_n2249_));
  NOR3_X1    g1607(.A1(new_n2236_), .A2(new_n2249_), .A3(new_n2242_), .ZN(new_n2250_));
  NOR2_X1    g1608(.A1(new_n2205_), .A2(new_n2207_), .ZN(new_n2251_));
  INV_X1     g1609(.I(new_n2251_), .ZN(new_n2252_));
  NOR4_X1    g1610(.A1(new_n2223_), .A2(new_n2250_), .A3(new_n2215_), .A4(new_n2252_), .ZN(new_n2253_));
  OAI21_X1   g1611(.A1(new_n2225_), .A2(new_n2202_), .B(new_n2253_), .ZN(new_n2254_));
  AOI21_X1   g1612(.A1(new_n2140_), .A2(new_n2185_), .B(new_n2254_), .ZN(new_n2255_));
  NOR2_X1    g1613(.A1(new_n1554_), .A2(\in2[78] ), .ZN(new_n2256_));
  AOI21_X1   g1614(.A1(new_n852_), .A2(new_n1554_), .B(new_n2256_), .ZN(new_n2257_));
  NOR2_X1    g1615(.A1(new_n1494_), .A2(\in0[78] ), .ZN(new_n2258_));
  AOI21_X1   g1616(.A1(new_n1252_), .A2(new_n1494_), .B(new_n2258_), .ZN(new_n2259_));
  NOR2_X1    g1617(.A1(new_n1046_), .A2(\in3[79] ), .ZN(new_n2260_));
  AOI21_X1   g1618(.A1(new_n851_), .A2(new_n1046_), .B(new_n2260_), .ZN(new_n2261_));
  INV_X1     g1619(.I(new_n2261_), .ZN(new_n2262_));
  NOR2_X1    g1620(.A1(new_n1494_), .A2(\in0[79] ), .ZN(new_n2263_));
  AOI21_X1   g1621(.A1(new_n1254_), .A2(new_n1494_), .B(new_n2263_), .ZN(new_n2264_));
  NOR2_X1    g1622(.A1(new_n2262_), .A2(new_n2264_), .ZN(new_n2265_));
  INV_X1     g1623(.I(new_n2265_), .ZN(new_n2266_));
  NAND2_X1   g1624(.A1(new_n2262_), .A2(new_n2264_), .ZN(new_n2267_));
  NAND3_X1   g1625(.A1(new_n2266_), .A2(new_n2259_), .A3(new_n2267_), .ZN(new_n2268_));
  NAND2_X1   g1626(.A1(new_n2268_), .A2(new_n2257_), .ZN(new_n2269_));
  NAND2_X1   g1627(.A1(new_n2262_), .A2(new_n2264_), .ZN(new_n2270_));
  XNOR2_X1   g1628(.A1(new_n2269_), .A2(new_n2270_), .ZN(new_n2271_));
  NOR2_X1    g1629(.A1(new_n1554_), .A2(\in2[76] ), .ZN(new_n2272_));
  AOI21_X1   g1630(.A1(new_n856_), .A2(new_n1554_), .B(new_n2272_), .ZN(new_n2273_));
  INV_X1     g1631(.I(new_n2273_), .ZN(new_n2274_));
  NOR2_X1    g1632(.A1(new_n1494_), .A2(\in0[76] ), .ZN(new_n2275_));
  AOI21_X1   g1633(.A1(new_n1256_), .A2(new_n1494_), .B(new_n2275_), .ZN(new_n2276_));
  NOR2_X1    g1634(.A1(new_n1494_), .A2(\in0[77] ), .ZN(new_n2277_));
  AOI21_X1   g1635(.A1(new_n1257_), .A2(new_n1494_), .B(new_n2277_), .ZN(new_n2278_));
  INV_X1     g1636(.I(new_n2278_), .ZN(new_n2279_));
  NOR2_X1    g1637(.A1(new_n1554_), .A2(\in2[77] ), .ZN(new_n2280_));
  AOI21_X1   g1638(.A1(new_n857_), .A2(new_n1554_), .B(new_n2280_), .ZN(new_n2281_));
  NOR2_X1    g1639(.A1(new_n2279_), .A2(new_n2281_), .ZN(new_n2282_));
  INV_X1     g1640(.I(new_n2281_), .ZN(new_n2283_));
  NOR2_X1    g1641(.A1(new_n2283_), .A2(new_n2278_), .ZN(new_n2284_));
  NOR2_X1    g1642(.A1(new_n2284_), .A2(new_n2282_), .ZN(new_n2285_));
  AOI21_X1   g1643(.A1(new_n2285_), .A2(new_n2276_), .B(new_n2274_), .ZN(new_n2286_));
  NOR2_X1    g1644(.A1(new_n2279_), .A2(new_n2281_), .ZN(new_n2287_));
  INV_X1     g1645(.I(new_n2287_), .ZN(new_n2288_));
  INV_X1     g1646(.I(new_n2257_), .ZN(new_n2289_));
  OAI21_X1   g1647(.A1(new_n2289_), .A2(new_n2259_), .B(new_n2266_), .ZN(new_n2290_));
  OAI21_X1   g1648(.A1(new_n2286_), .A2(new_n2288_), .B(new_n2290_), .ZN(new_n2291_));
  AOI21_X1   g1649(.A1(new_n2286_), .A2(new_n2288_), .B(new_n2291_), .ZN(new_n2292_));
  NOR4_X1    g1650(.A1(new_n2290_), .A2(new_n2274_), .A3(new_n2276_), .A4(new_n2284_), .ZN(new_n2293_));
  NAND2_X1   g1651(.A1(new_n2233_), .A2(new_n2235_), .ZN(new_n2294_));
  NAND2_X1   g1652(.A1(new_n2239_), .A2(new_n2241_), .ZN(new_n2295_));
  NAND2_X1   g1653(.A1(new_n2248_), .A2(new_n2295_), .ZN(new_n2296_));
  NAND2_X1   g1654(.A1(new_n2228_), .A2(new_n2230_), .ZN(new_n2297_));
  NAND4_X1   g1655(.A1(new_n2296_), .A2(new_n2236_), .A3(new_n2249_), .A4(new_n2297_), .ZN(new_n2298_));
  AOI21_X1   g1656(.A1(new_n2298_), .A2(new_n2294_), .B(new_n2293_), .ZN(new_n2299_));
  OAI21_X1   g1657(.A1(new_n2271_), .A2(new_n2292_), .B(new_n2299_), .ZN(new_n2300_));
  NOR2_X1    g1658(.A1(new_n1494_), .A2(\in0[82] ), .ZN(new_n2301_));
  AOI21_X1   g1659(.A1(new_n1270_), .A2(new_n1494_), .B(new_n2301_), .ZN(new_n2302_));
  INV_X1     g1660(.I(new_n2302_), .ZN(new_n2303_));
  NOR2_X1    g1661(.A1(new_n1554_), .A2(\in2[82] ), .ZN(new_n2304_));
  AOI21_X1   g1662(.A1(new_n870_), .A2(new_n1554_), .B(new_n2304_), .ZN(new_n2305_));
  NOR2_X1    g1663(.A1(new_n1494_), .A2(\in0[83] ), .ZN(new_n2306_));
  AOI21_X1   g1664(.A1(new_n1273_), .A2(new_n1494_), .B(new_n2306_), .ZN(new_n2307_));
  INV_X1     g1665(.I(new_n2307_), .ZN(new_n2308_));
  NOR2_X1    g1666(.A1(new_n1046_), .A2(\in3[83] ), .ZN(new_n2309_));
  AOI21_X1   g1667(.A1(new_n884_), .A2(new_n1046_), .B(new_n2309_), .ZN(new_n2310_));
  AOI22_X1   g1668(.A1(new_n2303_), .A2(new_n2305_), .B1(new_n2308_), .B2(new_n2310_), .ZN(new_n2311_));
  INV_X1     g1669(.I(new_n2311_), .ZN(new_n2312_));
  INV_X1     g1670(.I(new_n2305_), .ZN(new_n2313_));
  NOR2_X1    g1671(.A1(new_n1554_), .A2(\in2[81] ), .ZN(new_n2314_));
  AOI21_X1   g1672(.A1(new_n866_), .A2(new_n1554_), .B(new_n2314_), .ZN(new_n2315_));
  INV_X1     g1673(.I(new_n2315_), .ZN(new_n2316_));
  NOR2_X1    g1674(.A1(new_n1494_), .A2(\in0[81] ), .ZN(new_n2317_));
  AOI21_X1   g1675(.A1(new_n1266_), .A2(new_n1494_), .B(new_n2317_), .ZN(new_n2318_));
  NOR2_X1    g1676(.A1(new_n2316_), .A2(new_n2318_), .ZN(new_n2319_));
  NOR2_X1    g1677(.A1(new_n1494_), .A2(\in0[80] ), .ZN(new_n2320_));
  AOI21_X1   g1678(.A1(new_n1287_), .A2(new_n1494_), .B(new_n2320_), .ZN(new_n2321_));
  NOR2_X1    g1679(.A1(new_n1554_), .A2(\in2[80] ), .ZN(new_n2322_));
  AOI21_X1   g1680(.A1(new_n886_), .A2(new_n1554_), .B(new_n2322_), .ZN(new_n2323_));
  AOI21_X1   g1681(.A1(new_n2302_), .A2(new_n2313_), .B(new_n2319_), .ZN(new_n2324_));
  NAND2_X1   g1682(.A1(new_n2324_), .A2(new_n2312_), .ZN(new_n2325_));
  INV_X1     g1683(.I(new_n2325_), .ZN(new_n2326_));
  NOR2_X1    g1684(.A1(new_n1554_), .A2(\in2[86] ), .ZN(new_n2327_));
  AOI21_X1   g1685(.A1(new_n876_), .A2(new_n1554_), .B(new_n2327_), .ZN(new_n2328_));
  INV_X1     g1686(.I(new_n2328_), .ZN(new_n2329_));
  NOR2_X1    g1687(.A1(new_n1494_), .A2(\in0[86] ), .ZN(new_n2330_));
  AOI21_X1   g1688(.A1(new_n1308_), .A2(new_n1494_), .B(new_n2330_), .ZN(new_n2331_));
  NOR2_X1    g1689(.A1(new_n1046_), .A2(\in3[87] ), .ZN(new_n2332_));
  AOI21_X1   g1690(.A1(new_n907_), .A2(new_n1046_), .B(new_n2332_), .ZN(new_n2333_));
  INV_X1     g1691(.I(new_n2333_), .ZN(new_n2334_));
  NOR2_X1    g1692(.A1(new_n1568_), .A2(\in1[87] ), .ZN(new_n2335_));
  AOI21_X1   g1693(.A1(new_n1277_), .A2(new_n1568_), .B(new_n2335_), .ZN(new_n2336_));
  OAI22_X1   g1694(.A1(new_n2329_), .A2(new_n2331_), .B1(new_n2336_), .B2(new_n2334_), .ZN(new_n2337_));
  NOR2_X1    g1695(.A1(new_n1554_), .A2(\in2[85] ), .ZN(new_n2338_));
  AOI21_X1   g1696(.A1(new_n879_), .A2(new_n1554_), .B(new_n2338_), .ZN(new_n2339_));
  INV_X1     g1697(.I(new_n2339_), .ZN(new_n2340_));
  NOR2_X1    g1698(.A1(new_n1494_), .A2(\in0[85] ), .ZN(new_n2341_));
  AOI21_X1   g1699(.A1(new_n1280_), .A2(new_n1494_), .B(new_n2341_), .ZN(new_n2342_));
  NOR2_X1    g1700(.A1(new_n2340_), .A2(new_n2342_), .ZN(new_n2343_));
  NOR2_X1    g1701(.A1(new_n1554_), .A2(\in2[84] ), .ZN(new_n2344_));
  AOI21_X1   g1702(.A1(new_n881_), .A2(new_n1554_), .B(new_n2344_), .ZN(new_n2345_));
  INV_X1     g1703(.I(new_n2345_), .ZN(new_n2346_));
  NOR2_X1    g1704(.A1(new_n1494_), .A2(\in0[84] ), .ZN(new_n2347_));
  AOI21_X1   g1705(.A1(new_n1282_), .A2(new_n1494_), .B(new_n2347_), .ZN(new_n2348_));
  NOR4_X1    g1706(.A1(new_n2337_), .A2(new_n2343_), .A3(new_n2346_), .A4(new_n2348_), .ZN(new_n2349_));
  INV_X1     g1707(.I(new_n2323_), .ZN(new_n2350_));
  NOR2_X1    g1708(.A1(new_n2350_), .A2(new_n2321_), .ZN(new_n2351_));
  OAI21_X1   g1709(.A1(new_n2308_), .A2(new_n2310_), .B(new_n2319_), .ZN(new_n2352_));
  NOR3_X1    g1710(.A1(new_n2352_), .A2(new_n2312_), .A3(new_n2351_), .ZN(new_n2353_));
  INV_X1     g1711(.I(new_n2353_), .ZN(new_n2354_));
  NOR3_X1    g1712(.A1(new_n2354_), .A2(new_n2326_), .A3(new_n2349_), .ZN(new_n2355_));
  OAI21_X1   g1713(.A1(new_n2255_), .A2(new_n2300_), .B(new_n2355_), .ZN(new_n2356_));
  XNOR2_X1   g1714(.A1(new_n2339_), .A2(new_n2342_), .ZN(new_n2357_));
  AOI21_X1   g1715(.A1(new_n2357_), .A2(new_n2348_), .B(new_n2346_), .ZN(new_n2358_));
  NAND2_X1   g1716(.A1(new_n2340_), .A2(new_n2342_), .ZN(new_n2359_));
  OAI21_X1   g1717(.A1(new_n2358_), .A2(new_n2359_), .B(new_n2337_), .ZN(new_n2360_));
  AOI21_X1   g1718(.A1(new_n2358_), .A2(new_n2359_), .B(new_n2360_), .ZN(new_n2361_));
  XOR2_X1    g1719(.A1(new_n2336_), .A2(new_n2334_), .Z(new_n2362_));
  AOI21_X1   g1720(.A1(new_n2362_), .A2(new_n2331_), .B(new_n2329_), .ZN(new_n2363_));
  NAND2_X1   g1721(.A1(new_n2336_), .A2(new_n2334_), .ZN(new_n2364_));
  XOR2_X1    g1722(.A1(new_n2363_), .A2(new_n2364_), .Z(new_n2365_));
  NOR2_X1    g1723(.A1(new_n1494_), .A2(\in0[90] ), .ZN(new_n2366_));
  AOI21_X1   g1724(.A1(new_n1297_), .A2(new_n1494_), .B(new_n2366_), .ZN(new_n2367_));
  NOR2_X1    g1725(.A1(new_n1554_), .A2(\in2[90] ), .ZN(new_n2368_));
  AOI21_X1   g1726(.A1(new_n896_), .A2(new_n1554_), .B(new_n2368_), .ZN(new_n2369_));
  INV_X1     g1727(.I(new_n2369_), .ZN(new_n2370_));
  NOR2_X1    g1728(.A1(new_n1494_), .A2(\in0[91] ), .ZN(new_n2371_));
  AOI21_X1   g1729(.A1(new_n1301_), .A2(new_n1494_), .B(new_n2371_), .ZN(new_n2372_));
  NOR2_X1    g1730(.A1(new_n1554_), .A2(\in2[91] ), .ZN(new_n2373_));
  AOI21_X1   g1731(.A1(new_n900_), .A2(new_n1554_), .B(new_n2373_), .ZN(new_n2374_));
  INV_X1     g1732(.I(new_n2374_), .ZN(new_n2375_));
  OAI22_X1   g1733(.A1(new_n2367_), .A2(new_n2370_), .B1(new_n2375_), .B2(new_n2372_), .ZN(new_n2376_));
  NOR2_X1    g1734(.A1(new_n1554_), .A2(\in2[89] ), .ZN(new_n2377_));
  AOI21_X1   g1735(.A1(new_n892_), .A2(new_n1554_), .B(new_n2377_), .ZN(new_n2378_));
  INV_X1     g1736(.I(new_n2378_), .ZN(new_n2379_));
  NOR2_X1    g1737(.A1(new_n1494_), .A2(\in0[89] ), .ZN(new_n2380_));
  AOI21_X1   g1738(.A1(new_n1293_), .A2(new_n1494_), .B(new_n2380_), .ZN(new_n2381_));
  NOR2_X1    g1739(.A1(new_n2379_), .A2(new_n2381_), .ZN(new_n2382_));
  NOR2_X1    g1740(.A1(new_n1494_), .A2(\in0[88] ), .ZN(new_n2383_));
  AOI21_X1   g1741(.A1(new_n1310_), .A2(new_n1494_), .B(new_n2383_), .ZN(new_n2384_));
  NOR2_X1    g1742(.A1(new_n1046_), .A2(\in3[88] ), .ZN(new_n2385_));
  AOI21_X1   g1743(.A1(new_n909_), .A2(new_n1046_), .B(new_n2385_), .ZN(new_n2386_));
  AOI21_X1   g1744(.A1(new_n2367_), .A2(new_n2370_), .B(new_n2382_), .ZN(new_n2387_));
  NAND2_X1   g1745(.A1(new_n2387_), .A2(new_n2376_), .ZN(new_n2388_));
  NAND2_X1   g1746(.A1(new_n2375_), .A2(new_n2372_), .ZN(new_n2389_));
  INV_X1     g1747(.I(new_n2386_), .ZN(new_n2390_));
  OAI21_X1   g1748(.A1(new_n2384_), .A2(new_n2390_), .B(new_n2382_), .ZN(new_n2391_));
  OR2_X2     g1749(.A1(new_n2391_), .A2(new_n2376_), .Z(new_n2392_));
  NAND3_X1   g1750(.A1(new_n2392_), .A2(new_n2388_), .A3(new_n2389_), .ZN(new_n2393_));
  NOR3_X1    g1751(.A1(new_n2365_), .A2(new_n2361_), .A3(new_n2393_), .ZN(new_n2394_));
  NOR2_X1    g1752(.A1(new_n1554_), .A2(\in2[94] ), .ZN(new_n2395_));
  AOI21_X1   g1753(.A1(new_n914_), .A2(new_n1554_), .B(new_n2395_), .ZN(new_n2396_));
  NOR2_X1    g1754(.A1(new_n1494_), .A2(\in0[94] ), .ZN(new_n2397_));
  AOI21_X1   g1755(.A1(new_n1316_), .A2(new_n1494_), .B(new_n2397_), .ZN(new_n2398_));
  NOR2_X1    g1756(.A1(new_n1046_), .A2(\in3[95] ), .ZN(new_n2399_));
  AOI21_X1   g1757(.A1(new_n918_), .A2(new_n1046_), .B(new_n2399_), .ZN(new_n2400_));
  INV_X1     g1758(.I(new_n2400_), .ZN(new_n2401_));
  NOR2_X1    g1759(.A1(new_n1494_), .A2(\in0[95] ), .ZN(new_n2402_));
  AOI21_X1   g1760(.A1(new_n1317_), .A2(new_n1494_), .B(new_n2402_), .ZN(new_n2403_));
  NOR2_X1    g1761(.A1(new_n2401_), .A2(new_n2403_), .ZN(new_n2404_));
  INV_X1     g1762(.I(new_n2404_), .ZN(new_n2405_));
  NAND2_X1   g1763(.A1(new_n2401_), .A2(new_n2403_), .ZN(new_n2406_));
  NAND3_X1   g1764(.A1(new_n2405_), .A2(new_n2398_), .A3(new_n2406_), .ZN(new_n2407_));
  NAND2_X1   g1765(.A1(new_n2407_), .A2(new_n2396_), .ZN(new_n2408_));
  NAND2_X1   g1766(.A1(new_n2401_), .A2(new_n2403_), .ZN(new_n2409_));
  XNOR2_X1   g1767(.A1(new_n2408_), .A2(new_n2409_), .ZN(new_n2410_));
  NOR2_X1    g1768(.A1(new_n1554_), .A2(\in2[92] ), .ZN(new_n2411_));
  AOI21_X1   g1769(.A1(new_n921_), .A2(new_n1554_), .B(new_n2411_), .ZN(new_n2412_));
  INV_X1     g1770(.I(new_n2412_), .ZN(new_n2413_));
  NOR2_X1    g1771(.A1(new_n1494_), .A2(\in0[92] ), .ZN(new_n2414_));
  AOI21_X1   g1772(.A1(new_n1323_), .A2(new_n1494_), .B(new_n2414_), .ZN(new_n2415_));
  NOR2_X1    g1773(.A1(new_n1494_), .A2(\in0[93] ), .ZN(new_n2416_));
  AOI21_X1   g1774(.A1(new_n1334_), .A2(new_n1494_), .B(new_n2416_), .ZN(new_n2417_));
  INV_X1     g1775(.I(new_n2417_), .ZN(new_n2418_));
  NOR2_X1    g1776(.A1(new_n1046_), .A2(\in3[93] ), .ZN(new_n2419_));
  AOI21_X1   g1777(.A1(new_n920_), .A2(new_n1046_), .B(new_n2419_), .ZN(new_n2420_));
  NOR2_X1    g1778(.A1(new_n2418_), .A2(new_n2420_), .ZN(new_n2421_));
  INV_X1     g1779(.I(new_n2420_), .ZN(new_n2422_));
  NOR2_X1    g1780(.A1(new_n2422_), .A2(new_n2417_), .ZN(new_n2423_));
  NOR2_X1    g1781(.A1(new_n2421_), .A2(new_n2423_), .ZN(new_n2424_));
  AOI21_X1   g1782(.A1(new_n2424_), .A2(new_n2415_), .B(new_n2413_), .ZN(new_n2425_));
  INV_X1     g1783(.I(new_n2425_), .ZN(new_n2426_));
  NOR2_X1    g1784(.A1(new_n2418_), .A2(new_n2420_), .ZN(new_n2427_));
  NOR2_X1    g1785(.A1(new_n2426_), .A2(new_n2427_), .ZN(new_n2428_));
  NAND2_X1   g1786(.A1(new_n2426_), .A2(new_n2427_), .ZN(new_n2429_));
  INV_X1     g1787(.I(new_n2396_), .ZN(new_n2430_));
  OAI21_X1   g1788(.A1(new_n2430_), .A2(new_n2398_), .B(new_n2405_), .ZN(new_n2431_));
  NAND2_X1   g1789(.A1(new_n2429_), .A2(new_n2431_), .ZN(new_n2432_));
  NOR2_X1    g1790(.A1(new_n2432_), .A2(new_n2428_), .ZN(new_n2433_));
  NOR2_X1    g1791(.A1(new_n1046_), .A2(\in3[98] ), .ZN(new_n2434_));
  AOI21_X1   g1792(.A1(new_n925_), .A2(new_n1046_), .B(new_n2434_), .ZN(new_n2435_));
  INV_X1     g1793(.I(new_n2435_), .ZN(new_n2436_));
  NOR2_X1    g1794(.A1(new_n1568_), .A2(\in1[98] ), .ZN(new_n2437_));
  AOI21_X1   g1795(.A1(new_n1327_), .A2(new_n1568_), .B(new_n2437_), .ZN(new_n2438_));
  NOR2_X1    g1796(.A1(new_n1046_), .A2(\in3[99] ), .ZN(new_n2439_));
  AOI21_X1   g1797(.A1(new_n926_), .A2(new_n1046_), .B(new_n2439_), .ZN(new_n2440_));
  INV_X1     g1798(.I(new_n2440_), .ZN(new_n2441_));
  NOR2_X1    g1799(.A1(new_n1568_), .A2(\in1[99] ), .ZN(new_n2442_));
  AOI21_X1   g1800(.A1(new_n1328_), .A2(new_n1568_), .B(new_n2442_), .ZN(new_n2443_));
  OAI22_X1   g1801(.A1(new_n2436_), .A2(new_n2438_), .B1(new_n2443_), .B2(new_n2441_), .ZN(new_n2444_));
  NOR2_X1    g1802(.A1(new_n1046_), .A2(\in3[96] ), .ZN(new_n2445_));
  AOI21_X1   g1803(.A1(new_n924_), .A2(new_n1046_), .B(new_n2445_), .ZN(new_n2446_));
  INV_X1     g1804(.I(new_n2446_), .ZN(new_n2447_));
  NOR2_X1    g1805(.A1(new_n1568_), .A2(\in1[96] ), .ZN(new_n2448_));
  AOI21_X1   g1806(.A1(new_n1326_), .A2(new_n1568_), .B(new_n2448_), .ZN(new_n2449_));
  NOR2_X1    g1807(.A1(new_n2449_), .A2(new_n2447_), .ZN(new_n2450_));
  NOR2_X1    g1808(.A1(new_n1554_), .A2(\in2[97] ), .ZN(new_n2451_));
  AOI21_X1   g1809(.A1(new_n929_), .A2(new_n1554_), .B(new_n2451_), .ZN(new_n2452_));
  INV_X1     g1810(.I(new_n2452_), .ZN(new_n2453_));
  NOR2_X1    g1811(.A1(new_n1494_), .A2(\in0[97] ), .ZN(new_n2454_));
  AOI21_X1   g1812(.A1(new_n1331_), .A2(new_n1494_), .B(new_n2454_), .ZN(new_n2455_));
  NOR2_X1    g1813(.A1(new_n2453_), .A2(new_n2455_), .ZN(new_n2456_));
  INV_X1     g1814(.I(new_n2456_), .ZN(new_n2457_));
  NOR3_X1    g1815(.A1(new_n2457_), .A2(new_n2444_), .A3(new_n2450_), .ZN(new_n2458_));
  NOR2_X1    g1816(.A1(new_n2413_), .A2(new_n2415_), .ZN(new_n2459_));
  INV_X1     g1817(.I(new_n2459_), .ZN(new_n2460_));
  NOR4_X1    g1818(.A1(new_n2431_), .A2(new_n2458_), .A3(new_n2423_), .A4(new_n2460_), .ZN(new_n2461_));
  OAI21_X1   g1819(.A1(new_n2433_), .A2(new_n2410_), .B(new_n2461_), .ZN(new_n2462_));
  AOI21_X1   g1820(.A1(new_n2356_), .A2(new_n2394_), .B(new_n2462_), .ZN(new_n2463_));
  NOR2_X1    g1821(.A1(new_n1554_), .A2(\in2[102] ), .ZN(new_n2464_));
  AOI21_X1   g1822(.A1(new_n946_), .A2(new_n1554_), .B(new_n2464_), .ZN(new_n2465_));
  NOR2_X1    g1823(.A1(new_n1494_), .A2(\in0[102] ), .ZN(new_n2466_));
  AOI21_X1   g1824(.A1(new_n1348_), .A2(new_n1494_), .B(new_n2466_), .ZN(new_n2467_));
  NOR2_X1    g1825(.A1(new_n1046_), .A2(\in3[103] ), .ZN(new_n2468_));
  AOI21_X1   g1826(.A1(new_n945_), .A2(new_n1046_), .B(new_n2468_), .ZN(new_n2469_));
  INV_X1     g1827(.I(new_n2469_), .ZN(new_n2470_));
  NOR2_X1    g1828(.A1(new_n1494_), .A2(\in0[103] ), .ZN(new_n2471_));
  AOI21_X1   g1829(.A1(new_n1350_), .A2(new_n1494_), .B(new_n2471_), .ZN(new_n2472_));
  NOR2_X1    g1830(.A1(new_n2470_), .A2(new_n2472_), .ZN(new_n2473_));
  INV_X1     g1831(.I(new_n2473_), .ZN(new_n2474_));
  NAND2_X1   g1832(.A1(new_n2470_), .A2(new_n2472_), .ZN(new_n2475_));
  NAND3_X1   g1833(.A1(new_n2474_), .A2(new_n2467_), .A3(new_n2475_), .ZN(new_n2476_));
  NAND2_X1   g1834(.A1(new_n2476_), .A2(new_n2465_), .ZN(new_n2477_));
  NAND2_X1   g1835(.A1(new_n2470_), .A2(new_n2472_), .ZN(new_n2478_));
  XNOR2_X1   g1836(.A1(new_n2477_), .A2(new_n2478_), .ZN(new_n2479_));
  NOR2_X1    g1837(.A1(new_n1554_), .A2(\in2[100] ), .ZN(new_n2480_));
  AOI21_X1   g1838(.A1(new_n950_), .A2(new_n1554_), .B(new_n2480_), .ZN(new_n2481_));
  INV_X1     g1839(.I(new_n2481_), .ZN(new_n2482_));
  NOR2_X1    g1840(.A1(new_n1494_), .A2(\in0[100] ), .ZN(new_n2483_));
  AOI21_X1   g1841(.A1(new_n1352_), .A2(new_n1494_), .B(new_n2483_), .ZN(new_n2484_));
  NOR2_X1    g1842(.A1(new_n1494_), .A2(\in0[101] ), .ZN(new_n2485_));
  AOI21_X1   g1843(.A1(new_n1353_), .A2(new_n1494_), .B(new_n2485_), .ZN(new_n2486_));
  INV_X1     g1844(.I(new_n2486_), .ZN(new_n2487_));
  NOR2_X1    g1845(.A1(new_n1554_), .A2(\in2[101] ), .ZN(new_n2488_));
  AOI21_X1   g1846(.A1(new_n951_), .A2(new_n1554_), .B(new_n2488_), .ZN(new_n2489_));
  NOR2_X1    g1847(.A1(new_n2487_), .A2(new_n2489_), .ZN(new_n2490_));
  INV_X1     g1848(.I(new_n2489_), .ZN(new_n2491_));
  NOR2_X1    g1849(.A1(new_n2491_), .A2(new_n2486_), .ZN(new_n2492_));
  NOR2_X1    g1850(.A1(new_n2492_), .A2(new_n2490_), .ZN(new_n2493_));
  AOI21_X1   g1851(.A1(new_n2493_), .A2(new_n2484_), .B(new_n2482_), .ZN(new_n2494_));
  NOR2_X1    g1852(.A1(new_n2487_), .A2(new_n2489_), .ZN(new_n2495_));
  INV_X1     g1853(.I(new_n2495_), .ZN(new_n2496_));
  INV_X1     g1854(.I(new_n2465_), .ZN(new_n2497_));
  OAI21_X1   g1855(.A1(new_n2497_), .A2(new_n2467_), .B(new_n2474_), .ZN(new_n2498_));
  OAI21_X1   g1856(.A1(new_n2494_), .A2(new_n2496_), .B(new_n2498_), .ZN(new_n2499_));
  AOI21_X1   g1857(.A1(new_n2494_), .A2(new_n2496_), .B(new_n2499_), .ZN(new_n2500_));
  NOR4_X1    g1858(.A1(new_n2498_), .A2(new_n2482_), .A3(new_n2484_), .A4(new_n2492_), .ZN(new_n2501_));
  NAND2_X1   g1859(.A1(new_n2443_), .A2(new_n2441_), .ZN(new_n2502_));
  NAND2_X1   g1860(.A1(new_n2449_), .A2(new_n2447_), .ZN(new_n2503_));
  NAND2_X1   g1861(.A1(new_n2456_), .A2(new_n2503_), .ZN(new_n2504_));
  NAND2_X1   g1862(.A1(new_n2438_), .A2(new_n2436_), .ZN(new_n2505_));
  NAND4_X1   g1863(.A1(new_n2504_), .A2(new_n2457_), .A3(new_n2444_), .A4(new_n2505_), .ZN(new_n2506_));
  AOI21_X1   g1864(.A1(new_n2506_), .A2(new_n2502_), .B(new_n2501_), .ZN(new_n2507_));
  OAI21_X1   g1865(.A1(new_n2479_), .A2(new_n2500_), .B(new_n2507_), .ZN(new_n2508_));
  NOR2_X1    g1866(.A1(new_n1494_), .A2(\in0[106] ), .ZN(new_n2509_));
  AOI21_X1   g1867(.A1(new_n1366_), .A2(new_n1494_), .B(new_n2509_), .ZN(new_n2510_));
  INV_X1     g1868(.I(new_n2510_), .ZN(new_n2511_));
  NOR2_X1    g1869(.A1(new_n1554_), .A2(\in2[106] ), .ZN(new_n2512_));
  AOI21_X1   g1870(.A1(new_n964_), .A2(new_n1554_), .B(new_n2512_), .ZN(new_n2513_));
  NOR2_X1    g1871(.A1(new_n1494_), .A2(\in0[107] ), .ZN(new_n2514_));
  AOI21_X1   g1872(.A1(new_n1369_), .A2(new_n1494_), .B(new_n2514_), .ZN(new_n2515_));
  INV_X1     g1873(.I(new_n2515_), .ZN(new_n2516_));
  NOR2_X1    g1874(.A1(new_n1046_), .A2(\in3[107] ), .ZN(new_n2517_));
  AOI21_X1   g1875(.A1(new_n979_), .A2(new_n1046_), .B(new_n2517_), .ZN(new_n2518_));
  AOI22_X1   g1876(.A1(new_n2511_), .A2(new_n2513_), .B1(new_n2516_), .B2(new_n2518_), .ZN(new_n2519_));
  INV_X1     g1877(.I(new_n2519_), .ZN(new_n2520_));
  INV_X1     g1878(.I(new_n2513_), .ZN(new_n2521_));
  NOR2_X1    g1879(.A1(new_n1554_), .A2(\in2[105] ), .ZN(new_n2522_));
  AOI21_X1   g1880(.A1(new_n960_), .A2(new_n1554_), .B(new_n2522_), .ZN(new_n2523_));
  INV_X1     g1881(.I(new_n2523_), .ZN(new_n2524_));
  NOR2_X1    g1882(.A1(new_n1494_), .A2(\in0[105] ), .ZN(new_n2525_));
  AOI21_X1   g1883(.A1(new_n1362_), .A2(new_n1494_), .B(new_n2525_), .ZN(new_n2526_));
  NOR2_X1    g1884(.A1(new_n2524_), .A2(new_n2526_), .ZN(new_n2527_));
  NOR2_X1    g1885(.A1(new_n1494_), .A2(\in0[104] ), .ZN(new_n2528_));
  AOI21_X1   g1886(.A1(new_n1383_), .A2(new_n1494_), .B(new_n2528_), .ZN(new_n2529_));
  NOR2_X1    g1887(.A1(new_n1554_), .A2(\in2[104] ), .ZN(new_n2530_));
  AOI21_X1   g1888(.A1(new_n981_), .A2(new_n1554_), .B(new_n2530_), .ZN(new_n2531_));
  AOI21_X1   g1889(.A1(new_n2510_), .A2(new_n2521_), .B(new_n2527_), .ZN(new_n2532_));
  NAND2_X1   g1890(.A1(new_n2532_), .A2(new_n2520_), .ZN(new_n2533_));
  INV_X1     g1891(.I(new_n2533_), .ZN(new_n2534_));
  NOR2_X1    g1892(.A1(new_n1046_), .A2(\in3[110] ), .ZN(new_n2535_));
  AOI21_X1   g1893(.A1(new_n970_), .A2(new_n1046_), .B(new_n2535_), .ZN(new_n2536_));
  INV_X1     g1894(.I(new_n2536_), .ZN(new_n2537_));
  NOR2_X1    g1895(.A1(new_n1494_), .A2(\in0[110] ), .ZN(new_n2538_));
  AOI21_X1   g1896(.A1(new_n1404_), .A2(new_n1494_), .B(new_n2538_), .ZN(new_n2539_));
  NOR2_X1    g1897(.A1(new_n1046_), .A2(\in3[111] ), .ZN(new_n2540_));
  AOI21_X1   g1898(.A1(new_n971_), .A2(new_n1046_), .B(new_n2540_), .ZN(new_n2541_));
  INV_X1     g1899(.I(new_n2541_), .ZN(new_n2542_));
  NOR2_X1    g1900(.A1(new_n1568_), .A2(\in1[111] ), .ZN(new_n2543_));
  AOI21_X1   g1901(.A1(new_n1373_), .A2(new_n1568_), .B(new_n2543_), .ZN(new_n2544_));
  OAI22_X1   g1902(.A1(new_n2542_), .A2(new_n2544_), .B1(new_n2537_), .B2(new_n2539_), .ZN(new_n2545_));
  NOR2_X1    g1903(.A1(new_n1554_), .A2(\in2[109] ), .ZN(new_n2546_));
  AOI21_X1   g1904(.A1(new_n974_), .A2(new_n1554_), .B(new_n2546_), .ZN(new_n2547_));
  INV_X1     g1905(.I(new_n2547_), .ZN(new_n2548_));
  NOR2_X1    g1906(.A1(new_n1494_), .A2(\in0[109] ), .ZN(new_n2549_));
  AOI21_X1   g1907(.A1(new_n1376_), .A2(new_n1494_), .B(new_n2549_), .ZN(new_n2550_));
  NOR2_X1    g1908(.A1(new_n2548_), .A2(new_n2550_), .ZN(new_n2551_));
  NOR2_X1    g1909(.A1(new_n1554_), .A2(\in2[108] ), .ZN(new_n2552_));
  AOI21_X1   g1910(.A1(new_n976_), .A2(new_n1554_), .B(new_n2552_), .ZN(new_n2553_));
  INV_X1     g1911(.I(new_n2553_), .ZN(new_n2554_));
  NOR2_X1    g1912(.A1(new_n1494_), .A2(\in0[108] ), .ZN(new_n2555_));
  AOI21_X1   g1913(.A1(new_n1378_), .A2(new_n1494_), .B(new_n2555_), .ZN(new_n2556_));
  NOR4_X1    g1914(.A1(new_n2545_), .A2(new_n2551_), .A3(new_n2554_), .A4(new_n2556_), .ZN(new_n2557_));
  INV_X1     g1915(.I(new_n2531_), .ZN(new_n2558_));
  NOR2_X1    g1916(.A1(new_n2558_), .A2(new_n2529_), .ZN(new_n2559_));
  OAI21_X1   g1917(.A1(new_n2516_), .A2(new_n2518_), .B(new_n2527_), .ZN(new_n2560_));
  NOR3_X1    g1918(.A1(new_n2560_), .A2(new_n2520_), .A3(new_n2559_), .ZN(new_n2561_));
  INV_X1     g1919(.I(new_n2561_), .ZN(new_n2562_));
  NOR3_X1    g1920(.A1(new_n2562_), .A2(new_n2534_), .A3(new_n2557_), .ZN(new_n2563_));
  OAI21_X1   g1921(.A1(new_n2463_), .A2(new_n2508_), .B(new_n2563_), .ZN(new_n2564_));
  XNOR2_X1   g1922(.A1(new_n2547_), .A2(new_n2550_), .ZN(new_n2565_));
  AOI21_X1   g1923(.A1(new_n2565_), .A2(new_n2556_), .B(new_n2554_), .ZN(new_n2566_));
  NAND2_X1   g1924(.A1(new_n2548_), .A2(new_n2550_), .ZN(new_n2567_));
  OAI21_X1   g1925(.A1(new_n2566_), .A2(new_n2567_), .B(new_n2545_), .ZN(new_n2568_));
  AOI21_X1   g1926(.A1(new_n2566_), .A2(new_n2567_), .B(new_n2568_), .ZN(new_n2569_));
  XOR2_X1    g1927(.A1(new_n2544_), .A2(new_n2542_), .Z(new_n2570_));
  AOI21_X1   g1928(.A1(new_n2570_), .A2(new_n2539_), .B(new_n2537_), .ZN(new_n2571_));
  NAND2_X1   g1929(.A1(new_n2544_), .A2(new_n2542_), .ZN(new_n2572_));
  XOR2_X1    g1930(.A1(new_n2571_), .A2(new_n2572_), .Z(new_n2573_));
  NOR2_X1    g1931(.A1(new_n1494_), .A2(\in0[114] ), .ZN(new_n2574_));
  AOI21_X1   g1932(.A1(new_n1393_), .A2(new_n1494_), .B(new_n2574_), .ZN(new_n2575_));
  NOR2_X1    g1933(.A1(new_n1554_), .A2(\in2[114] ), .ZN(new_n2576_));
  AOI21_X1   g1934(.A1(new_n991_), .A2(new_n1554_), .B(new_n2576_), .ZN(new_n2577_));
  INV_X1     g1935(.I(new_n2577_), .ZN(new_n2578_));
  NOR2_X1    g1936(.A1(new_n1494_), .A2(\in0[115] ), .ZN(new_n2579_));
  AOI21_X1   g1937(.A1(new_n1397_), .A2(new_n1494_), .B(new_n2579_), .ZN(new_n2580_));
  NOR2_X1    g1938(.A1(new_n1554_), .A2(\in2[115] ), .ZN(new_n2581_));
  AOI21_X1   g1939(.A1(new_n995_), .A2(new_n1554_), .B(new_n2581_), .ZN(new_n2582_));
  INV_X1     g1940(.I(new_n2582_), .ZN(new_n2583_));
  OAI22_X1   g1941(.A1(new_n2575_), .A2(new_n2578_), .B1(new_n2583_), .B2(new_n2580_), .ZN(new_n2584_));
  NOR2_X1    g1942(.A1(new_n1554_), .A2(\in2[113] ), .ZN(new_n2585_));
  AOI21_X1   g1943(.A1(new_n987_), .A2(new_n1554_), .B(new_n2585_), .ZN(new_n2586_));
  INV_X1     g1944(.I(new_n2586_), .ZN(new_n2587_));
  NOR2_X1    g1945(.A1(new_n1494_), .A2(\in0[113] ), .ZN(new_n2588_));
  AOI21_X1   g1946(.A1(new_n1389_), .A2(new_n1494_), .B(new_n2588_), .ZN(new_n2589_));
  NOR2_X1    g1947(.A1(new_n2587_), .A2(new_n2589_), .ZN(new_n2590_));
  NOR2_X1    g1948(.A1(new_n1494_), .A2(\in0[112] ), .ZN(new_n2591_));
  AOI21_X1   g1949(.A1(new_n1406_), .A2(new_n1494_), .B(new_n2591_), .ZN(new_n2592_));
  NOR2_X1    g1950(.A1(new_n1046_), .A2(\in3[112] ), .ZN(new_n2593_));
  AOI21_X1   g1951(.A1(new_n1004_), .A2(new_n1046_), .B(new_n2593_), .ZN(new_n2594_));
  AOI21_X1   g1952(.A1(new_n2575_), .A2(new_n2578_), .B(new_n2590_), .ZN(new_n2595_));
  NAND2_X1   g1953(.A1(new_n2595_), .A2(new_n2584_), .ZN(new_n2596_));
  NAND2_X1   g1954(.A1(new_n2583_), .A2(new_n2580_), .ZN(new_n2597_));
  INV_X1     g1955(.I(new_n2594_), .ZN(new_n2598_));
  OAI21_X1   g1956(.A1(new_n2592_), .A2(new_n2598_), .B(new_n2590_), .ZN(new_n2599_));
  OR2_X2     g1957(.A1(new_n2599_), .A2(new_n2584_), .Z(new_n2600_));
  NAND3_X1   g1958(.A1(new_n2600_), .A2(new_n2596_), .A3(new_n2597_), .ZN(new_n2601_));
  NOR3_X1    g1959(.A1(new_n2573_), .A2(new_n2569_), .A3(new_n2601_), .ZN(new_n2602_));
  NOR2_X1    g1960(.A1(new_n1554_), .A2(\in2[118] ), .ZN(new_n2603_));
  AOI21_X1   g1961(.A1(new_n1009_), .A2(new_n1554_), .B(new_n2603_), .ZN(new_n2604_));
  NOR2_X1    g1962(.A1(new_n1494_), .A2(\in0[118] ), .ZN(new_n2605_));
  AOI21_X1   g1963(.A1(new_n1412_), .A2(new_n1494_), .B(new_n2605_), .ZN(new_n2606_));
  NOR2_X1    g1964(.A1(new_n1046_), .A2(\in3[119] ), .ZN(new_n2607_));
  AOI21_X1   g1965(.A1(new_n1013_), .A2(new_n1046_), .B(new_n2607_), .ZN(new_n2608_));
  INV_X1     g1966(.I(new_n2608_), .ZN(new_n2609_));
  NOR2_X1    g1967(.A1(new_n1494_), .A2(\in0[119] ), .ZN(new_n2610_));
  AOI21_X1   g1968(.A1(new_n1413_), .A2(new_n1494_), .B(new_n2610_), .ZN(new_n2611_));
  NOR2_X1    g1969(.A1(new_n2609_), .A2(new_n2611_), .ZN(new_n2612_));
  INV_X1     g1970(.I(new_n2612_), .ZN(new_n2613_));
  NAND2_X1   g1971(.A1(new_n2609_), .A2(new_n2611_), .ZN(new_n2614_));
  NAND3_X1   g1972(.A1(new_n2613_), .A2(new_n2606_), .A3(new_n2614_), .ZN(new_n2615_));
  NAND2_X1   g1973(.A1(new_n2615_), .A2(new_n2604_), .ZN(new_n2616_));
  NAND2_X1   g1974(.A1(new_n2609_), .A2(new_n2611_), .ZN(new_n2617_));
  XNOR2_X1   g1975(.A1(new_n2616_), .A2(new_n2617_), .ZN(new_n2618_));
  NOR2_X1    g1976(.A1(new_n1554_), .A2(\in2[116] ), .ZN(new_n2619_));
  AOI21_X1   g1977(.A1(new_n1016_), .A2(new_n1554_), .B(new_n2619_), .ZN(new_n2620_));
  INV_X1     g1978(.I(new_n2620_), .ZN(new_n2621_));
  NOR2_X1    g1979(.A1(new_n1494_), .A2(\in0[116] ), .ZN(new_n2622_));
  AOI21_X1   g1980(.A1(new_n1419_), .A2(new_n1494_), .B(new_n2622_), .ZN(new_n2623_));
  NOR2_X1    g1981(.A1(new_n1494_), .A2(\in0[117] ), .ZN(new_n2624_));
  AOI21_X1   g1982(.A1(new_n1430_), .A2(new_n1494_), .B(new_n2624_), .ZN(new_n2625_));
  INV_X1     g1983(.I(new_n2625_), .ZN(new_n2626_));
  NOR2_X1    g1984(.A1(new_n1046_), .A2(\in3[117] ), .ZN(new_n2627_));
  AOI21_X1   g1985(.A1(new_n1015_), .A2(new_n1046_), .B(new_n2627_), .ZN(new_n2628_));
  NOR2_X1    g1986(.A1(new_n2626_), .A2(new_n2628_), .ZN(new_n2629_));
  INV_X1     g1987(.I(new_n2628_), .ZN(new_n2630_));
  NOR2_X1    g1988(.A1(new_n2630_), .A2(new_n2625_), .ZN(new_n2631_));
  NOR2_X1    g1989(.A1(new_n2629_), .A2(new_n2631_), .ZN(new_n2632_));
  AOI21_X1   g1990(.A1(new_n2632_), .A2(new_n2623_), .B(new_n2621_), .ZN(new_n2633_));
  INV_X1     g1991(.I(new_n2633_), .ZN(new_n2634_));
  NOR2_X1    g1992(.A1(new_n2626_), .A2(new_n2628_), .ZN(new_n2635_));
  NOR2_X1    g1993(.A1(new_n2634_), .A2(new_n2635_), .ZN(new_n2636_));
  NAND2_X1   g1994(.A1(new_n2634_), .A2(new_n2635_), .ZN(new_n2637_));
  INV_X1     g1995(.I(new_n2604_), .ZN(new_n2638_));
  OAI21_X1   g1996(.A1(new_n2638_), .A2(new_n2606_), .B(new_n2613_), .ZN(new_n2639_));
  NAND2_X1   g1997(.A1(new_n2637_), .A2(new_n2639_), .ZN(new_n2640_));
  NOR2_X1    g1998(.A1(new_n2640_), .A2(new_n2636_), .ZN(new_n2641_));
  NOR2_X1    g1999(.A1(new_n1046_), .A2(\in3[122] ), .ZN(new_n2642_));
  AOI21_X1   g2000(.A1(new_n1020_), .A2(new_n1046_), .B(new_n2642_), .ZN(new_n2643_));
  NOR2_X1    g2001(.A1(new_n1494_), .A2(\in0[122] ), .ZN(new_n2644_));
  AOI21_X1   g2002(.A1(new_n1441_), .A2(new_n1494_), .B(new_n2644_), .ZN(new_n2645_));
  INV_X1     g2003(.I(new_n2645_), .ZN(new_n2646_));
  NOR2_X1    g2004(.A1(new_n1046_), .A2(\in3[123] ), .ZN(new_n2647_));
  AOI21_X1   g2005(.A1(new_n1021_), .A2(new_n1046_), .B(new_n2647_), .ZN(new_n2648_));
  INV_X1     g2006(.I(\in1[123] ), .ZN(new_n2649_));
  NOR2_X1    g2007(.A1(new_n1494_), .A2(\in0[123] ), .ZN(new_n2650_));
  AOI21_X1   g2008(.A1(new_n2649_), .A2(new_n1494_), .B(new_n2650_), .ZN(new_n2651_));
  INV_X1     g2009(.I(new_n2651_), .ZN(new_n2652_));
  AOI22_X1   g2010(.A1(new_n2643_), .A2(new_n2646_), .B1(new_n2652_), .B2(new_n2648_), .ZN(new_n2653_));
  INV_X1     g2011(.I(new_n2653_), .ZN(new_n2654_));
  NOR2_X1    g2012(.A1(new_n1046_), .A2(\in3[120] ), .ZN(new_n2655_));
  AOI21_X1   g2013(.A1(new_n1019_), .A2(new_n1046_), .B(new_n2655_), .ZN(new_n2656_));
  INV_X1     g2014(.I(new_n2656_), .ZN(new_n2657_));
  NOR2_X1    g2015(.A1(new_n1568_), .A2(\in1[120] ), .ZN(new_n2658_));
  AOI21_X1   g2016(.A1(new_n1422_), .A2(new_n1568_), .B(new_n2658_), .ZN(new_n2659_));
  NOR2_X1    g2017(.A1(new_n1554_), .A2(\in2[121] ), .ZN(new_n2660_));
  AOI21_X1   g2018(.A1(new_n1024_), .A2(new_n1554_), .B(new_n2660_), .ZN(new_n2661_));
  INV_X1     g2019(.I(new_n2661_), .ZN(new_n2662_));
  NOR2_X1    g2020(.A1(new_n1494_), .A2(\in0[121] ), .ZN(new_n2663_));
  AOI21_X1   g2021(.A1(new_n1427_), .A2(new_n1494_), .B(new_n2663_), .ZN(new_n2664_));
  NOR2_X1    g2022(.A1(new_n2662_), .A2(new_n2664_), .ZN(new_n2665_));
  OAI21_X1   g2023(.A1(new_n2657_), .A2(new_n2659_), .B(new_n2665_), .ZN(new_n2666_));
  NOR2_X1    g2024(.A1(new_n2666_), .A2(new_n2654_), .ZN(new_n2667_));
  NOR2_X1    g2025(.A1(new_n2621_), .A2(new_n2623_), .ZN(new_n2668_));
  INV_X1     g2026(.I(new_n2668_), .ZN(new_n2669_));
  NOR4_X1    g2027(.A1(new_n2667_), .A2(new_n2631_), .A3(new_n2639_), .A4(new_n2669_), .ZN(new_n2670_));
  OAI21_X1   g2028(.A1(new_n2641_), .A2(new_n2618_), .B(new_n2670_), .ZN(new_n2671_));
  AOI21_X1   g2029(.A1(new_n2564_), .A2(new_n2602_), .B(new_n2671_), .ZN(new_n2672_));
  OR3_X2     g2030(.A1(new_n1557_), .A2(new_n1452_), .A3(new_n1508_), .Z(new_n2673_));
  NOR2_X1    g2031(.A1(new_n2652_), .A2(new_n2648_), .ZN(new_n2674_));
  INV_X1     g2032(.I(new_n2665_), .ZN(new_n2675_));
  AOI21_X1   g2033(.A1(new_n2657_), .A2(new_n2659_), .B(new_n2675_), .ZN(new_n2676_));
  NOR2_X1    g2034(.A1(new_n2646_), .A2(new_n2643_), .ZN(new_n2677_));
  NOR4_X1    g2035(.A1(new_n2676_), .A2(new_n2653_), .A3(new_n2665_), .A4(new_n2677_), .ZN(new_n2678_));
  OAI22_X1   g2036(.A1(new_n2678_), .A2(new_n2674_), .B1(new_n1506_), .B2(new_n2673_), .ZN(new_n2679_));
  OAI21_X1   g2037(.A1(new_n2672_), .A2(new_n2679_), .B(new_n1562_), .ZN(new_n2680_));
  NOR2_X1    g2038(.A1(new_n1494_), .A2(\in0[0] ), .ZN(new_n2681_));
  NOR2_X1    g2039(.A1(new_n1568_), .A2(\in1[0] ), .ZN(new_n2682_));
  NOR2_X1    g2040(.A1(new_n2682_), .A2(new_n2681_), .ZN(new_n2683_));
  NAND4_X1   g2041(.A1(new_n2680_), .A2(new_n1047_), .A3(new_n1451_), .A4(new_n2683_), .ZN(new_n2684_));
  INV_X1     g2042(.I(new_n1047_), .ZN(new_n2685_));
  NAND2_X1   g2043(.A1(new_n1876_), .A2(new_n1871_), .ZN(new_n2686_));
  INV_X1     g2044(.I(new_n1931_), .ZN(new_n2687_));
  AOI21_X1   g2045(.A1(new_n1875_), .A2(new_n1928_), .B(new_n2687_), .ZN(new_n2688_));
  AOI21_X1   g2046(.A1(new_n2686_), .A2(new_n2688_), .B(new_n2021_), .ZN(new_n2689_));
  INV_X1     g2047(.I(new_n2139_), .ZN(new_n2690_));
  OAI21_X1   g2048(.A1(new_n2689_), .A2(new_n2690_), .B(new_n2185_), .ZN(new_n2691_));
  INV_X1     g2049(.I(new_n2254_), .ZN(new_n2692_));
  AOI21_X1   g2050(.A1(new_n2691_), .A2(new_n2692_), .B(new_n2300_), .ZN(new_n2693_));
  INV_X1     g2051(.I(new_n2355_), .ZN(new_n2694_));
  OAI21_X1   g2052(.A1(new_n2693_), .A2(new_n2694_), .B(new_n2394_), .ZN(new_n2695_));
  INV_X1     g2053(.I(new_n2462_), .ZN(new_n2696_));
  AOI21_X1   g2054(.A1(new_n2695_), .A2(new_n2696_), .B(new_n2508_), .ZN(new_n2697_));
  INV_X1     g2055(.I(new_n2563_), .ZN(new_n2698_));
  OAI21_X1   g2056(.A1(new_n2697_), .A2(new_n2698_), .B(new_n2602_), .ZN(new_n2699_));
  INV_X1     g2057(.I(new_n2671_), .ZN(new_n2700_));
  AOI21_X1   g2058(.A1(new_n2699_), .A2(new_n2700_), .B(new_n2679_), .ZN(new_n2701_));
  OAI21_X1   g2059(.A1(new_n2701_), .A2(new_n1561_), .B(new_n1451_), .ZN(new_n2702_));
  OAI21_X1   g2060(.A1(new_n2702_), .A2(new_n2683_), .B(new_n2685_), .ZN(new_n2703_));
  NAND2_X1   g2061(.A1(new_n2703_), .A2(new_n2684_), .ZN(\result[0] ));
  INV_X1     g2062(.I(\in3[1] ), .ZN(new_n2705_));
  NOR2_X1    g2063(.A1(new_n1554_), .A2(\in2[1] ), .ZN(new_n2706_));
  AOI21_X1   g2064(.A1(new_n2705_), .A2(new_n1554_), .B(new_n2706_), .ZN(new_n2707_));
  NOR2_X1    g2065(.A1(new_n1494_), .A2(\in0[1] ), .ZN(new_n2708_));
  NOR2_X1    g2066(.A1(new_n1568_), .A2(\in1[1] ), .ZN(new_n2709_));
  NOR2_X1    g2067(.A1(new_n2709_), .A2(new_n2708_), .ZN(new_n2710_));
  NAND4_X1   g2068(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2707_), .A4(new_n2710_), .ZN(new_n2711_));
  INV_X1     g2069(.I(new_n2707_), .ZN(new_n2712_));
  OAI21_X1   g2070(.A1(new_n2702_), .A2(new_n2710_), .B(new_n2712_), .ZN(new_n2713_));
  NAND2_X1   g2071(.A1(new_n2713_), .A2(new_n2711_), .ZN(\result[1] ));
  INV_X1     g2072(.I(\in3[2] ), .ZN(new_n2715_));
  MUX2_X1    g2073(.I0(\in2[2] ), .I1(new_n2715_), .S(new_n1046_), .Z(new_n2716_));
  NOR2_X1    g2074(.A1(new_n1494_), .A2(\in0[2] ), .ZN(new_n2717_));
  NOR2_X1    g2075(.A1(new_n1568_), .A2(\in1[2] ), .ZN(new_n2718_));
  NOR2_X1    g2076(.A1(new_n2718_), .A2(new_n2717_), .ZN(new_n2719_));
  NAND4_X1   g2077(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2716_), .A4(new_n2719_), .ZN(new_n2720_));
  INV_X1     g2078(.I(new_n2716_), .ZN(new_n2721_));
  OAI21_X1   g2079(.A1(new_n2702_), .A2(new_n2719_), .B(new_n2721_), .ZN(new_n2722_));
  NAND2_X1   g2080(.A1(new_n2722_), .A2(new_n2720_), .ZN(\result[2] ));
  INV_X1     g2081(.I(\in3[3] ), .ZN(new_n2724_));
  NOR2_X1    g2082(.A1(new_n1554_), .A2(\in2[3] ), .ZN(new_n2725_));
  AOI21_X1   g2083(.A1(new_n2724_), .A2(new_n1554_), .B(new_n2725_), .ZN(new_n2726_));
  NOR2_X1    g2084(.A1(new_n1494_), .A2(\in0[3] ), .ZN(new_n2727_));
  NOR2_X1    g2085(.A1(new_n1568_), .A2(\in1[3] ), .ZN(new_n2728_));
  NOR2_X1    g2086(.A1(new_n2728_), .A2(new_n2727_), .ZN(new_n2729_));
  NAND4_X1   g2087(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2726_), .A4(new_n2729_), .ZN(new_n2730_));
  INV_X1     g2088(.I(new_n2726_), .ZN(new_n2731_));
  OAI21_X1   g2089(.A1(new_n2702_), .A2(new_n2729_), .B(new_n2731_), .ZN(new_n2732_));
  NAND2_X1   g2090(.A1(new_n2732_), .A2(new_n2730_), .ZN(\result[3] ));
  INV_X1     g2091(.I(\in3[4] ), .ZN(new_n2734_));
  NOR2_X1    g2092(.A1(new_n1554_), .A2(\in2[4] ), .ZN(new_n2735_));
  AOI21_X1   g2093(.A1(new_n2734_), .A2(new_n1554_), .B(new_n2735_), .ZN(new_n2736_));
  NOR2_X1    g2094(.A1(new_n1494_), .A2(\in0[4] ), .ZN(new_n2737_));
  NOR2_X1    g2095(.A1(new_n1568_), .A2(\in1[4] ), .ZN(new_n2738_));
  NOR2_X1    g2096(.A1(new_n2738_), .A2(new_n2737_), .ZN(new_n2739_));
  NAND4_X1   g2097(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2736_), .A4(new_n2739_), .ZN(new_n2740_));
  INV_X1     g2098(.I(new_n2736_), .ZN(new_n2741_));
  OAI21_X1   g2099(.A1(new_n2702_), .A2(new_n2739_), .B(new_n2741_), .ZN(new_n2742_));
  NAND2_X1   g2100(.A1(new_n2742_), .A2(new_n2740_), .ZN(\result[4] ));
  INV_X1     g2101(.I(\in3[5] ), .ZN(new_n2744_));
  NOR2_X1    g2102(.A1(new_n1554_), .A2(\in2[5] ), .ZN(new_n2745_));
  AOI21_X1   g2103(.A1(new_n2744_), .A2(new_n1554_), .B(new_n2745_), .ZN(new_n2746_));
  NOR2_X1    g2104(.A1(new_n1494_), .A2(\in0[5] ), .ZN(new_n2747_));
  NOR2_X1    g2105(.A1(new_n1568_), .A2(\in1[5] ), .ZN(new_n2748_));
  NOR2_X1    g2106(.A1(new_n2748_), .A2(new_n2747_), .ZN(new_n2749_));
  NAND4_X1   g2107(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2746_), .A4(new_n2749_), .ZN(new_n2750_));
  INV_X1     g2108(.I(new_n2746_), .ZN(new_n2751_));
  OAI21_X1   g2109(.A1(new_n2702_), .A2(new_n2749_), .B(new_n2751_), .ZN(new_n2752_));
  NAND2_X1   g2110(.A1(new_n2752_), .A2(new_n2750_), .ZN(\result[5] ));
  INV_X1     g2111(.I(\in3[6] ), .ZN(new_n2754_));
  NOR2_X1    g2112(.A1(new_n1554_), .A2(\in2[6] ), .ZN(new_n2755_));
  AOI21_X1   g2113(.A1(new_n2754_), .A2(new_n1554_), .B(new_n2755_), .ZN(new_n2756_));
  NOR2_X1    g2114(.A1(new_n1494_), .A2(\in0[6] ), .ZN(new_n2757_));
  NOR2_X1    g2115(.A1(new_n1568_), .A2(\in1[6] ), .ZN(new_n2758_));
  NOR2_X1    g2116(.A1(new_n2758_), .A2(new_n2757_), .ZN(new_n2759_));
  NAND4_X1   g2117(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2756_), .A4(new_n2759_), .ZN(new_n2760_));
  INV_X1     g2118(.I(new_n2756_), .ZN(new_n2761_));
  OAI21_X1   g2119(.A1(new_n2702_), .A2(new_n2759_), .B(new_n2761_), .ZN(new_n2762_));
  NAND2_X1   g2120(.A1(new_n2762_), .A2(new_n2760_), .ZN(\result[6] ));
  INV_X1     g2121(.I(\in3[7] ), .ZN(new_n2764_));
  NOR2_X1    g2122(.A1(new_n1554_), .A2(\in2[7] ), .ZN(new_n2765_));
  AOI21_X1   g2123(.A1(new_n2764_), .A2(new_n1554_), .B(new_n2765_), .ZN(new_n2766_));
  NOR2_X1    g2124(.A1(new_n1494_), .A2(\in0[7] ), .ZN(new_n2767_));
  NOR2_X1    g2125(.A1(new_n1568_), .A2(\in1[7] ), .ZN(new_n2768_));
  NOR2_X1    g2126(.A1(new_n2768_), .A2(new_n2767_), .ZN(new_n2769_));
  NAND4_X1   g2127(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2766_), .A4(new_n2769_), .ZN(new_n2770_));
  INV_X1     g2128(.I(new_n2766_), .ZN(new_n2771_));
  OAI21_X1   g2129(.A1(new_n2702_), .A2(new_n2769_), .B(new_n2771_), .ZN(new_n2772_));
  NAND2_X1   g2130(.A1(new_n2772_), .A2(new_n2770_), .ZN(\result[7] ));
  INV_X1     g2131(.I(\in3[8] ), .ZN(new_n2774_));
  NOR2_X1    g2132(.A1(new_n1554_), .A2(\in2[8] ), .ZN(new_n2775_));
  AOI21_X1   g2133(.A1(new_n2774_), .A2(new_n1554_), .B(new_n2775_), .ZN(new_n2776_));
  NOR2_X1    g2134(.A1(new_n1494_), .A2(\in0[8] ), .ZN(new_n2777_));
  NOR2_X1    g2135(.A1(new_n1568_), .A2(\in1[8] ), .ZN(new_n2778_));
  NOR2_X1    g2136(.A1(new_n2778_), .A2(new_n2777_), .ZN(new_n2779_));
  NAND4_X1   g2137(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2776_), .A4(new_n2779_), .ZN(new_n2780_));
  INV_X1     g2138(.I(new_n2776_), .ZN(new_n2781_));
  OAI21_X1   g2139(.A1(new_n2702_), .A2(new_n2779_), .B(new_n2781_), .ZN(new_n2782_));
  NAND2_X1   g2140(.A1(new_n2782_), .A2(new_n2780_), .ZN(\result[8] ));
  NAND4_X1   g2141(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1600_), .A4(new_n1619_), .ZN(new_n2784_));
  OAI21_X1   g2142(.A1(new_n2702_), .A2(new_n1600_), .B(new_n1605_), .ZN(new_n2785_));
  NAND2_X1   g2143(.A1(new_n2785_), .A2(new_n2784_), .ZN(\result[9] ));
  NAND4_X1   g2144(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1592_), .A4(new_n1589_), .ZN(new_n2787_));
  OAI21_X1   g2145(.A1(new_n2702_), .A2(new_n1589_), .B(new_n1585_), .ZN(new_n2788_));
  NAND2_X1   g2146(.A1(new_n2788_), .A2(new_n2787_), .ZN(\result[10] ));
  NAND4_X1   g2147(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1624_), .A4(new_n1628_), .ZN(new_n2790_));
  OAI21_X1   g2148(.A1(new_n2702_), .A2(new_n1628_), .B(new_n1609_), .ZN(new_n2791_));
  NAND2_X1   g2149(.A1(new_n2791_), .A2(new_n2790_), .ZN(\result[11] ));
  NAND4_X1   g2150(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1634_), .A4(new_n1666_), .ZN(new_n2793_));
  OAI21_X1   g2151(.A1(new_n2702_), .A2(new_n1634_), .B(new_n1637_), .ZN(new_n2794_));
  NAND2_X1   g2152(.A1(new_n2794_), .A2(new_n2793_), .ZN(\result[12] ));
  NAND4_X1   g2153(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1648_), .A4(new_n1645_), .ZN(new_n2796_));
  OAI21_X1   g2154(.A1(new_n2702_), .A2(new_n1645_), .B(new_n1642_), .ZN(new_n2797_));
  NAND2_X1   g2155(.A1(new_n2797_), .A2(new_n2796_), .ZN(\result[13] ));
  NAND4_X1   g2156(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1656_), .A4(new_n1676_), .ZN(new_n2799_));
  OAI21_X1   g2157(.A1(new_n2702_), .A2(new_n1676_), .B(new_n1657_), .ZN(new_n2800_));
  NAND2_X1   g2158(.A1(new_n2800_), .A2(new_n2799_), .ZN(\result[14] ));
  NAND4_X1   g2159(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1574_), .A4(new_n1578_), .ZN(new_n2802_));
  OAI21_X1   g2160(.A1(new_n2702_), .A2(new_n1578_), .B(new_n1575_), .ZN(new_n2803_));
  NAND2_X1   g2161(.A1(new_n2803_), .A2(new_n2802_), .ZN(\result[15] ));
  NAND4_X1   g2162(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1683_), .A4(new_n1686_), .ZN(new_n2805_));
  INV_X1     g2163(.I(new_n1683_), .ZN(new_n2806_));
  OAI21_X1   g2164(.A1(new_n2702_), .A2(new_n1686_), .B(new_n2806_), .ZN(new_n2807_));
  NAND2_X1   g2165(.A1(new_n2807_), .A2(new_n2805_), .ZN(\result[16] ));
  NAND4_X1   g2166(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1692_), .A4(new_n1695_), .ZN(new_n2809_));
  OAI21_X1   g2167(.A1(new_n2702_), .A2(new_n1692_), .B(new_n1696_), .ZN(new_n2810_));
  NAND2_X1   g2168(.A1(new_n2810_), .A2(new_n2809_), .ZN(\result[17] ));
  NAND4_X1   g2169(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1704_), .A4(new_n1707_), .ZN(new_n2812_));
  OAI21_X1   g2170(.A1(new_n2702_), .A2(new_n1707_), .B(new_n1710_), .ZN(new_n2813_));
  NAND2_X1   g2171(.A1(new_n2813_), .A2(new_n2812_), .ZN(\result[18] ));
  NAND4_X1   g2172(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1716_), .A4(new_n1729_), .ZN(new_n2815_));
  OAI21_X1   g2173(.A1(new_n2702_), .A2(new_n1729_), .B(new_n1725_), .ZN(new_n2816_));
  NAND2_X1   g2174(.A1(new_n2816_), .A2(new_n2815_), .ZN(\result[19] ));
  NAND4_X1   g2175(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1734_), .A4(new_n1737_), .ZN(new_n2818_));
  OAI21_X1   g2176(.A1(new_n2702_), .A2(new_n1734_), .B(new_n1738_), .ZN(new_n2819_));
  NAND2_X1   g2177(.A1(new_n2819_), .A2(new_n2818_), .ZN(\result[20] ));
  NAND4_X1   g2178(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1745_), .A4(new_n1748_), .ZN(new_n2821_));
  OAI21_X1   g2179(.A1(new_n2702_), .A2(new_n1748_), .B(new_n1751_), .ZN(new_n2822_));
  NAND2_X1   g2180(.A1(new_n2822_), .A2(new_n2821_), .ZN(\result[21] ));
  NAND4_X1   g2181(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1757_), .A4(new_n1769_), .ZN(new_n2824_));
  OAI21_X1   g2182(.A1(new_n2702_), .A2(new_n1769_), .B(new_n1765_), .ZN(new_n2825_));
  NAND2_X1   g2183(.A1(new_n2825_), .A2(new_n2824_), .ZN(\result[22] ));
  NAND4_X1   g2184(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1565_), .A4(new_n1570_), .ZN(new_n2827_));
  OAI21_X1   g2185(.A1(new_n2702_), .A2(new_n1570_), .B(new_n1566_), .ZN(new_n2828_));
  NAND2_X1   g2186(.A1(new_n2828_), .A2(new_n2827_), .ZN(\result[23] ));
  NAND4_X1   g2187(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1776_), .A4(new_n1779_), .ZN(new_n2830_));
  INV_X1     g2188(.I(new_n1776_), .ZN(new_n2831_));
  OAI21_X1   g2189(.A1(new_n2702_), .A2(new_n1779_), .B(new_n2831_), .ZN(new_n2832_));
  NAND2_X1   g2190(.A1(new_n2832_), .A2(new_n2830_), .ZN(\result[24] ));
  NAND4_X1   g2191(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1784_), .A4(new_n1787_), .ZN(new_n2834_));
  OAI21_X1   g2192(.A1(new_n2702_), .A2(new_n1784_), .B(new_n1788_), .ZN(new_n2835_));
  NAND2_X1   g2193(.A1(new_n2835_), .A2(new_n2834_), .ZN(\result[25] ));
  NAND4_X1   g2194(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1795_), .A4(new_n1798_), .ZN(new_n2837_));
  OAI21_X1   g2195(.A1(new_n2702_), .A2(new_n1798_), .B(new_n1801_), .ZN(new_n2838_));
  NAND2_X1   g2196(.A1(new_n2838_), .A2(new_n2837_), .ZN(\result[26] ));
  NAND4_X1   g2197(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1806_), .A4(new_n1824_), .ZN(new_n2840_));
  OAI21_X1   g2198(.A1(new_n2702_), .A2(new_n1824_), .B(new_n1807_), .ZN(new_n2841_));
  NAND2_X1   g2199(.A1(new_n2841_), .A2(new_n2840_), .ZN(\result[27] ));
  NAND4_X1   g2200(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1829_), .A4(new_n1832_), .ZN(new_n2843_));
  OAI21_X1   g2201(.A1(new_n2702_), .A2(new_n1829_), .B(new_n1833_), .ZN(new_n2844_));
  NAND2_X1   g2202(.A1(new_n2844_), .A2(new_n2843_), .ZN(\result[28] ));
  NAND4_X1   g2203(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1839_), .A4(new_n1842_), .ZN(new_n2846_));
  OAI21_X1   g2204(.A1(new_n2702_), .A2(new_n1842_), .B(new_n1845_), .ZN(new_n2847_));
  NAND2_X1   g2205(.A1(new_n2847_), .A2(new_n2846_), .ZN(\result[29] ));
  NAND4_X1   g2206(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1852_), .A4(new_n1866_), .ZN(new_n2849_));
  OAI21_X1   g2207(.A1(new_n2702_), .A2(new_n1866_), .B(new_n1853_), .ZN(new_n2850_));
  NAND2_X1   g2208(.A1(new_n2850_), .A2(new_n2849_), .ZN(\result[30] ));
  NAND4_X1   g2209(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1869_), .A4(new_n1931_), .ZN(new_n2852_));
  OAI21_X1   g2210(.A1(new_n2702_), .A2(new_n1869_), .B(new_n2687_), .ZN(new_n2853_));
  NAND2_X1   g2211(.A1(new_n2853_), .A2(new_n2852_), .ZN(\result[31] ));
  NAND4_X1   g2212(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1903_), .A4(new_n1905_), .ZN(new_n2855_));
  OAI21_X1   g2213(.A1(new_n2702_), .A2(new_n1903_), .B(new_n1906_), .ZN(new_n2856_));
  NAND2_X1   g2214(.A1(new_n2856_), .A2(new_n2855_), .ZN(\result[32] ));
  NAND4_X1   g2215(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1914_), .A4(new_n1916_), .ZN(new_n2858_));
  INV_X1     g2216(.I(new_n1914_), .ZN(new_n2859_));
  OAI21_X1   g2217(.A1(new_n2702_), .A2(new_n1916_), .B(new_n2859_), .ZN(new_n2860_));
  NAND2_X1   g2218(.A1(new_n2860_), .A2(new_n2858_), .ZN(\result[33] ));
  NAND4_X1   g2219(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1920_), .A4(new_n1922_), .ZN(new_n2862_));
  OAI21_X1   g2220(.A1(new_n2702_), .A2(new_n1920_), .B(new_n1923_), .ZN(new_n2863_));
  NAND2_X1   g2221(.A1(new_n2863_), .A2(new_n2862_), .ZN(\result[34] ));
  NAND4_X1   g2222(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1908_), .A4(new_n1911_), .ZN(new_n2865_));
  INV_X1     g2223(.I(new_n1908_), .ZN(new_n2866_));
  OAI21_X1   g2224(.A1(new_n2702_), .A2(new_n1911_), .B(new_n2866_), .ZN(new_n2867_));
  NAND2_X1   g2225(.A1(new_n2867_), .A2(new_n2865_), .ZN(\result[35] ));
  NAND4_X1   g2226(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1896_), .A4(new_n1900_), .ZN(new_n2869_));
  OAI21_X1   g2227(.A1(new_n2702_), .A2(new_n1900_), .B(new_n1897_), .ZN(new_n2870_));
  NAND2_X1   g2228(.A1(new_n2870_), .A2(new_n2869_), .ZN(\result[36] ));
  NAND4_X1   g2229(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1890_), .A4(new_n1893_), .ZN(new_n2872_));
  OAI21_X1   g2230(.A1(new_n2702_), .A2(new_n1893_), .B(new_n1891_), .ZN(new_n2873_));
  NAND2_X1   g2231(.A1(new_n2873_), .A2(new_n2872_), .ZN(\result[37] ));
  NAND4_X1   g2232(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1879_), .A4(new_n1882_), .ZN(new_n2875_));
  OAI21_X1   g2233(.A1(new_n2702_), .A2(new_n1882_), .B(new_n1880_), .ZN(new_n2876_));
  NAND2_X1   g2234(.A1(new_n2876_), .A2(new_n2875_), .ZN(\result[38] ));
  NAND4_X1   g2235(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1884_), .A4(new_n1887_), .ZN(new_n2878_));
  OAI21_X1   g2236(.A1(new_n2702_), .A2(new_n1887_), .B(new_n1885_), .ZN(new_n2879_));
  NAND2_X1   g2237(.A1(new_n2879_), .A2(new_n2878_), .ZN(\result[39] ));
  NAND4_X1   g2238(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1986_), .A4(new_n1988_), .ZN(new_n2881_));
  OAI21_X1   g2239(.A1(new_n2702_), .A2(new_n1986_), .B(new_n2009_), .ZN(new_n2882_));
  NAND2_X1   g2240(.A1(new_n2882_), .A2(new_n2881_), .ZN(\result[40] ));
  NAND4_X1   g2241(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1979_), .A4(new_n1982_), .ZN(new_n2884_));
  OAI21_X1   g2242(.A1(new_n2702_), .A2(new_n1982_), .B(new_n1980_), .ZN(new_n2885_));
  NAND2_X1   g2243(.A1(new_n2885_), .A2(new_n2884_), .ZN(\result[41] ));
  NAND4_X1   g2244(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1972_), .A4(new_n1975_), .ZN(new_n2887_));
  INV_X1     g2245(.I(new_n1975_), .ZN(new_n2888_));
  OAI21_X1   g2246(.A1(new_n2702_), .A2(new_n1972_), .B(new_n2888_), .ZN(new_n2889_));
  NAND2_X1   g2247(.A1(new_n2889_), .A2(new_n2887_), .ZN(\result[42] ));
  NAND4_X1   g2248(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1966_), .A4(new_n1968_), .ZN(new_n2891_));
  OAI21_X1   g2249(.A1(new_n2702_), .A2(new_n1966_), .B(new_n1969_), .ZN(new_n2892_));
  NAND2_X1   g2250(.A1(new_n2892_), .A2(new_n2891_), .ZN(\result[43] ));
  NAND4_X1   g2251(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1947_), .A4(new_n1950_), .ZN(new_n2894_));
  OAI21_X1   g2252(.A1(new_n2702_), .A2(new_n1947_), .B(new_n1962_), .ZN(new_n2895_));
  NAND2_X1   g2253(.A1(new_n2895_), .A2(new_n2894_), .ZN(\result[44] ));
  NAND4_X1   g2254(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1955_), .A4(new_n1953_), .ZN(new_n2897_));
  OAI21_X1   g2255(.A1(new_n2702_), .A2(new_n1955_), .B(new_n1956_), .ZN(new_n2898_));
  NAND2_X1   g2256(.A1(new_n2898_), .A2(new_n2897_), .ZN(\result[45] ));
  NAND4_X1   g2257(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1935_), .A4(new_n1938_), .ZN(new_n2900_));
  OAI21_X1   g2258(.A1(new_n2702_), .A2(new_n1938_), .B(new_n1936_), .ZN(new_n2901_));
  NAND2_X1   g2259(.A1(new_n2901_), .A2(new_n2900_), .ZN(\result[46] ));
  NAND4_X1   g2260(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1940_), .A4(new_n1943_), .ZN(new_n2903_));
  OAI21_X1   g2261(.A1(new_n2702_), .A2(new_n1943_), .B(new_n1941_), .ZN(new_n2904_));
  NAND2_X1   g2262(.A1(new_n2904_), .A2(new_n2903_), .ZN(\result[47] ));
  NAND4_X1   g2263(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2049_), .A4(new_n2051_), .ZN(new_n2906_));
  OAI21_X1   g2264(.A1(new_n2702_), .A2(new_n2049_), .B(new_n2052_), .ZN(new_n2907_));
  NAND2_X1   g2265(.A1(new_n2907_), .A2(new_n2906_), .ZN(\result[48] ));
  NAND4_X1   g2266(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2041_), .A4(new_n2044_), .ZN(new_n2909_));
  OAI21_X1   g2267(.A1(new_n2702_), .A2(new_n2044_), .B(new_n2042_), .ZN(new_n2910_));
  NAND2_X1   g2268(.A1(new_n2910_), .A2(new_n2909_), .ZN(\result[49] ));
  NAND4_X1   g2269(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2023_), .A4(new_n2025_), .ZN(new_n2912_));
  OAI21_X1   g2270(.A1(new_n2702_), .A2(new_n2025_), .B(new_n2039_), .ZN(new_n2913_));
  NAND2_X1   g2271(.A1(new_n2913_), .A2(new_n2912_), .ZN(\result[50] ));
  NAND4_X1   g2272(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2027_), .A4(new_n2030_), .ZN(new_n2915_));
  OAI21_X1   g2273(.A1(new_n2702_), .A2(new_n2030_), .B(new_n2028_), .ZN(new_n2916_));
  NAND2_X1   g2274(.A1(new_n2916_), .A2(new_n2915_), .ZN(\result[51] ));
  NAND4_X1   g2275(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2075_), .A4(new_n2077_), .ZN(new_n2918_));
  OAI21_X1   g2276(.A1(new_n2702_), .A2(new_n2075_), .B(new_n2083_), .ZN(new_n2919_));
  NAND2_X1   g2277(.A1(new_n2919_), .A2(new_n2918_), .ZN(\result[52] ));
  NAND4_X1   g2278(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2069_), .A4(new_n2072_), .ZN(new_n2921_));
  OAI21_X1   g2279(.A1(new_n2702_), .A2(new_n2072_), .B(new_n2070_), .ZN(new_n2922_));
  NAND2_X1   g2280(.A1(new_n2922_), .A2(new_n2921_), .ZN(\result[53] ));
  NAND4_X1   g2281(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2056_), .A4(new_n2059_), .ZN(new_n2924_));
  OAI21_X1   g2282(.A1(new_n2702_), .A2(new_n2056_), .B(new_n2067_), .ZN(new_n2925_));
  NAND2_X1   g2283(.A1(new_n2925_), .A2(new_n2924_), .ZN(\result[54] ));
  NAND4_X1   g2284(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2061_), .A4(new_n2064_), .ZN(new_n2927_));
  INV_X1     g2285(.I(new_n2064_), .ZN(new_n2928_));
  OAI21_X1   g2286(.A1(new_n2702_), .A2(new_n2061_), .B(new_n2928_), .ZN(new_n2929_));
  NAND2_X1   g2287(.A1(new_n2929_), .A2(new_n2927_), .ZN(\result[55] ));
  NAND4_X1   g2288(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2113_), .A4(new_n2116_), .ZN(new_n2931_));
  OAI21_X1   g2289(.A1(new_n2702_), .A2(new_n2116_), .B(new_n2114_), .ZN(new_n2932_));
  NAND2_X1   g2290(.A1(new_n2932_), .A2(new_n2931_), .ZN(\result[56] ));
  NAND4_X1   g2291(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2119_), .A4(new_n2122_), .ZN(new_n2934_));
  OAI21_X1   g2292(.A1(new_n2702_), .A2(new_n2122_), .B(new_n2120_), .ZN(new_n2935_));
  NAND2_X1   g2293(.A1(new_n2935_), .A2(new_n2934_), .ZN(\result[57] ));
  NAND4_X1   g2294(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2126_), .A4(new_n2128_), .ZN(new_n2937_));
  INV_X1     g2295(.I(new_n2126_), .ZN(new_n2938_));
  OAI21_X1   g2296(.A1(new_n2702_), .A2(new_n2128_), .B(new_n2938_), .ZN(new_n2939_));
  NAND2_X1   g2297(.A1(new_n2939_), .A2(new_n2937_), .ZN(\result[58] ));
  NAND4_X1   g2298(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2131_), .A4(new_n2133_), .ZN(new_n2941_));
  INV_X1     g2299(.I(new_n2131_), .ZN(new_n2942_));
  OAI21_X1   g2300(.A1(new_n2702_), .A2(new_n2133_), .B(new_n2942_), .ZN(new_n2943_));
  NAND2_X1   g2301(.A1(new_n2943_), .A2(new_n2941_), .ZN(\result[59] ));
  NAND4_X1   g2302(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2106_), .A4(new_n2109_), .ZN(new_n2945_));
  OAI21_X1   g2303(.A1(new_n2702_), .A2(new_n2109_), .B(new_n2107_), .ZN(new_n2946_));
  NAND2_X1   g2304(.A1(new_n2946_), .A2(new_n2945_), .ZN(\result[60] ));
  NAND4_X1   g2305(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2100_), .A4(new_n2103_), .ZN(new_n2948_));
  OAI21_X1   g2306(.A1(new_n2702_), .A2(new_n2103_), .B(new_n2101_), .ZN(new_n2949_));
  NAND2_X1   g2307(.A1(new_n2949_), .A2(new_n2948_), .ZN(\result[61] ));
  NAND4_X1   g2308(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2089_), .A4(new_n2092_), .ZN(new_n2951_));
  OAI21_X1   g2309(.A1(new_n2702_), .A2(new_n2092_), .B(new_n2090_), .ZN(new_n2952_));
  NAND2_X1   g2310(.A1(new_n2952_), .A2(new_n2951_), .ZN(\result[62] ));
  NAND4_X1   g2311(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2094_), .A4(new_n2097_), .ZN(new_n2954_));
  OAI21_X1   g2312(.A1(new_n2702_), .A2(new_n2097_), .B(new_n2095_), .ZN(new_n2955_));
  NAND2_X1   g2313(.A1(new_n2955_), .A2(new_n2954_), .ZN(\result[63] ));
  NAND4_X1   g2314(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2159_), .A4(new_n2161_), .ZN(new_n2957_));
  OAI21_X1   g2315(.A1(new_n2702_), .A2(new_n2159_), .B(new_n2165_), .ZN(new_n2958_));
  NAND2_X1   g2316(.A1(new_n2958_), .A2(new_n2957_), .ZN(\result[64] ));
  NAND4_X1   g2317(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2153_), .A4(new_n2156_), .ZN(new_n2960_));
  OAI21_X1   g2318(.A1(new_n2702_), .A2(new_n2156_), .B(new_n2154_), .ZN(new_n2961_));
  NAND2_X1   g2319(.A1(new_n2961_), .A2(new_n2960_), .ZN(\result[65] ));
  NAND4_X1   g2320(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2142_), .A4(new_n2144_), .ZN(new_n2963_));
  OAI21_X1   g2321(.A1(new_n2702_), .A2(new_n2142_), .B(new_n2145_), .ZN(new_n2964_));
  NAND2_X1   g2322(.A1(new_n2964_), .A2(new_n2963_), .ZN(\result[66] ));
  NAND4_X1   g2323(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2147_), .A4(new_n2149_), .ZN(new_n2966_));
  OAI21_X1   g2324(.A1(new_n2702_), .A2(new_n2147_), .B(new_n2150_), .ZN(new_n2967_));
  NAND2_X1   g2325(.A1(new_n2967_), .A2(new_n2966_), .ZN(\result[67] ));
  NAND4_X1   g2326(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2204_), .A4(new_n2207_), .ZN(new_n2969_));
  OAI21_X1   g2327(.A1(new_n2702_), .A2(new_n2207_), .B(new_n2205_), .ZN(new_n2970_));
  NAND2_X1   g2328(.A1(new_n2970_), .A2(new_n2969_), .ZN(\result[68] ));
  NAND4_X1   g2329(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2209_), .A4(new_n2212_), .ZN(new_n2972_));
  OAI21_X1   g2330(.A1(new_n2702_), .A2(new_n2209_), .B(new_n2214_), .ZN(new_n2973_));
  NAND2_X1   g2331(.A1(new_n2973_), .A2(new_n2972_), .ZN(\result[69] ));
  NAND4_X1   g2332(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2188_), .A4(new_n2190_), .ZN(new_n2975_));
  OAI21_X1   g2333(.A1(new_n2702_), .A2(new_n2190_), .B(new_n2222_), .ZN(new_n2976_));
  NAND2_X1   g2334(.A1(new_n2976_), .A2(new_n2975_), .ZN(\result[70] ));
  NAND4_X1   g2335(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2192_), .A4(new_n2195_), .ZN(new_n2978_));
  OAI21_X1   g2336(.A1(new_n2702_), .A2(new_n2195_), .B(new_n2193_), .ZN(new_n2979_));
  NAND2_X1   g2337(.A1(new_n2979_), .A2(new_n2978_), .ZN(\result[71] ));
  NAND4_X1   g2338(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2238_), .A4(new_n2241_), .ZN(new_n2981_));
  OAI21_X1   g2339(.A1(new_n2702_), .A2(new_n2241_), .B(new_n2239_), .ZN(new_n2982_));
  NAND2_X1   g2340(.A1(new_n2982_), .A2(new_n2981_), .ZN(\result[72] ));
  NAND4_X1   g2341(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2244_), .A4(new_n2247_), .ZN(new_n2984_));
  OAI21_X1   g2342(.A1(new_n2702_), .A2(new_n2247_), .B(new_n2245_), .ZN(new_n2985_));
  NAND2_X1   g2343(.A1(new_n2985_), .A2(new_n2984_), .ZN(\result[73] ));
  NAND4_X1   g2344(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2227_), .A4(new_n2230_), .ZN(new_n2987_));
  OAI21_X1   g2345(.A1(new_n2702_), .A2(new_n2230_), .B(new_n2228_), .ZN(new_n2988_));
  NAND2_X1   g2346(.A1(new_n2988_), .A2(new_n2987_), .ZN(\result[74] ));
  NAND4_X1   g2347(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2232_), .A4(new_n2235_), .ZN(new_n2990_));
  OAI21_X1   g2348(.A1(new_n2702_), .A2(new_n2235_), .B(new_n2233_), .ZN(new_n2991_));
  NAND2_X1   g2349(.A1(new_n2991_), .A2(new_n2990_), .ZN(\result[75] ));
  NAND4_X1   g2350(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2273_), .A4(new_n2276_), .ZN(new_n2993_));
  OAI21_X1   g2351(.A1(new_n2702_), .A2(new_n2276_), .B(new_n2274_), .ZN(new_n2994_));
  NAND2_X1   g2352(.A1(new_n2994_), .A2(new_n2993_), .ZN(\result[76] ));
  NAND4_X1   g2353(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2278_), .A4(new_n2281_), .ZN(new_n2996_));
  OAI21_X1   g2354(.A1(new_n2702_), .A2(new_n2278_), .B(new_n2283_), .ZN(new_n2997_));
  NAND2_X1   g2355(.A1(new_n2997_), .A2(new_n2996_), .ZN(\result[77] ));
  NAND4_X1   g2356(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2257_), .A4(new_n2259_), .ZN(new_n2999_));
  OAI21_X1   g2357(.A1(new_n2702_), .A2(new_n2259_), .B(new_n2289_), .ZN(new_n3000_));
  NAND2_X1   g2358(.A1(new_n3000_), .A2(new_n2999_), .ZN(\result[78] ));
  NAND4_X1   g2359(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2261_), .A4(new_n2264_), .ZN(new_n3002_));
  OAI21_X1   g2360(.A1(new_n2702_), .A2(new_n2264_), .B(new_n2262_), .ZN(new_n3003_));
  NAND2_X1   g2361(.A1(new_n3003_), .A2(new_n3002_), .ZN(\result[79] ));
  NAND4_X1   g2362(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2321_), .A4(new_n2323_), .ZN(new_n3005_));
  OAI21_X1   g2363(.A1(new_n2702_), .A2(new_n2321_), .B(new_n2350_), .ZN(new_n3006_));
  NAND2_X1   g2364(.A1(new_n3006_), .A2(new_n3005_), .ZN(\result[80] ));
  NAND4_X1   g2365(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2315_), .A4(new_n2318_), .ZN(new_n3008_));
  OAI21_X1   g2366(.A1(new_n2702_), .A2(new_n2318_), .B(new_n2316_), .ZN(new_n3009_));
  NAND2_X1   g2367(.A1(new_n3009_), .A2(new_n3008_), .ZN(\result[81] ));
  NAND4_X1   g2368(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2302_), .A4(new_n2305_), .ZN(new_n3011_));
  OAI21_X1   g2369(.A1(new_n2702_), .A2(new_n2302_), .B(new_n2313_), .ZN(new_n3012_));
  NAND2_X1   g2370(.A1(new_n3012_), .A2(new_n3011_), .ZN(\result[82] ));
  NAND4_X1   g2371(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2307_), .A4(new_n2310_), .ZN(new_n3014_));
  INV_X1     g2372(.I(new_n2310_), .ZN(new_n3015_));
  OAI21_X1   g2373(.A1(new_n2702_), .A2(new_n2307_), .B(new_n3015_), .ZN(new_n3016_));
  NAND2_X1   g2374(.A1(new_n3016_), .A2(new_n3014_), .ZN(\result[83] ));
  NAND4_X1   g2375(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2345_), .A4(new_n2348_), .ZN(new_n3018_));
  OAI21_X1   g2376(.A1(new_n2702_), .A2(new_n2348_), .B(new_n2346_), .ZN(new_n3019_));
  NAND2_X1   g2377(.A1(new_n3019_), .A2(new_n3018_), .ZN(\result[84] ));
  NAND4_X1   g2378(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2339_), .A4(new_n2342_), .ZN(new_n3021_));
  OAI21_X1   g2379(.A1(new_n2702_), .A2(new_n2342_), .B(new_n2340_), .ZN(new_n3022_));
  NAND2_X1   g2380(.A1(new_n3022_), .A2(new_n3021_), .ZN(\result[85] ));
  NAND4_X1   g2381(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2328_), .A4(new_n2331_), .ZN(new_n3024_));
  OAI21_X1   g2382(.A1(new_n2702_), .A2(new_n2331_), .B(new_n2329_), .ZN(new_n3025_));
  NAND2_X1   g2383(.A1(new_n3025_), .A2(new_n3024_), .ZN(\result[86] ));
  NAND4_X1   g2384(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2333_), .A4(new_n2336_), .ZN(new_n3027_));
  OAI21_X1   g2385(.A1(new_n2702_), .A2(new_n2336_), .B(new_n2334_), .ZN(new_n3028_));
  NAND2_X1   g2386(.A1(new_n3028_), .A2(new_n3027_), .ZN(\result[87] ));
  NAND4_X1   g2387(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2384_), .A4(new_n2386_), .ZN(new_n3030_));
  OAI21_X1   g2388(.A1(new_n2702_), .A2(new_n2384_), .B(new_n2390_), .ZN(new_n3031_));
  NAND2_X1   g2389(.A1(new_n3031_), .A2(new_n3030_), .ZN(\result[88] ));
  NAND4_X1   g2390(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2378_), .A4(new_n2381_), .ZN(new_n3033_));
  OAI21_X1   g2391(.A1(new_n2702_), .A2(new_n2381_), .B(new_n2379_), .ZN(new_n3034_));
  NAND2_X1   g2392(.A1(new_n3034_), .A2(new_n3033_), .ZN(\result[89] ));
  NAND4_X1   g2393(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2367_), .A4(new_n2369_), .ZN(new_n3036_));
  OAI21_X1   g2394(.A1(new_n2702_), .A2(new_n2367_), .B(new_n2370_), .ZN(new_n3037_));
  NAND2_X1   g2395(.A1(new_n3037_), .A2(new_n3036_), .ZN(\result[90] ));
  NAND4_X1   g2396(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2372_), .A4(new_n2374_), .ZN(new_n3039_));
  OAI21_X1   g2397(.A1(new_n2702_), .A2(new_n2372_), .B(new_n2375_), .ZN(new_n3040_));
  NAND2_X1   g2398(.A1(new_n3040_), .A2(new_n3039_), .ZN(\result[91] ));
  NAND4_X1   g2399(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2412_), .A4(new_n2415_), .ZN(new_n3042_));
  OAI21_X1   g2400(.A1(new_n2702_), .A2(new_n2415_), .B(new_n2413_), .ZN(new_n3043_));
  NAND2_X1   g2401(.A1(new_n3043_), .A2(new_n3042_), .ZN(\result[92] ));
  NAND4_X1   g2402(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2417_), .A4(new_n2420_), .ZN(new_n3045_));
  OAI21_X1   g2403(.A1(new_n2702_), .A2(new_n2417_), .B(new_n2422_), .ZN(new_n3046_));
  NAND2_X1   g2404(.A1(new_n3046_), .A2(new_n3045_), .ZN(\result[93] ));
  NAND4_X1   g2405(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2396_), .A4(new_n2398_), .ZN(new_n3048_));
  OAI21_X1   g2406(.A1(new_n2702_), .A2(new_n2398_), .B(new_n2430_), .ZN(new_n3049_));
  NAND2_X1   g2407(.A1(new_n3049_), .A2(new_n3048_), .ZN(\result[94] ));
  NAND4_X1   g2408(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2400_), .A4(new_n2403_), .ZN(new_n3051_));
  OAI21_X1   g2409(.A1(new_n2702_), .A2(new_n2403_), .B(new_n2401_), .ZN(new_n3052_));
  NAND2_X1   g2410(.A1(new_n3052_), .A2(new_n3051_), .ZN(\result[95] ));
  NAND4_X1   g2411(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2446_), .A4(new_n2449_), .ZN(new_n3054_));
  OAI21_X1   g2412(.A1(new_n2702_), .A2(new_n2449_), .B(new_n2447_), .ZN(new_n3055_));
  NAND2_X1   g2413(.A1(new_n3055_), .A2(new_n3054_), .ZN(\result[96] ));
  NAND4_X1   g2414(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2452_), .A4(new_n2455_), .ZN(new_n3057_));
  OAI21_X1   g2415(.A1(new_n2702_), .A2(new_n2455_), .B(new_n2453_), .ZN(new_n3058_));
  NAND2_X1   g2416(.A1(new_n3058_), .A2(new_n3057_), .ZN(\result[97] ));
  NAND4_X1   g2417(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2435_), .A4(new_n2438_), .ZN(new_n3060_));
  OAI21_X1   g2418(.A1(new_n2702_), .A2(new_n2438_), .B(new_n2436_), .ZN(new_n3061_));
  NAND2_X1   g2419(.A1(new_n3061_), .A2(new_n3060_), .ZN(\result[98] ));
  NAND4_X1   g2420(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2440_), .A4(new_n2443_), .ZN(new_n3063_));
  OAI21_X1   g2421(.A1(new_n2702_), .A2(new_n2443_), .B(new_n2441_), .ZN(new_n3064_));
  NAND2_X1   g2422(.A1(new_n3064_), .A2(new_n3063_), .ZN(\result[99] ));
  NAND4_X1   g2423(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2481_), .A4(new_n2484_), .ZN(new_n3066_));
  OAI21_X1   g2424(.A1(new_n2702_), .A2(new_n2484_), .B(new_n2482_), .ZN(new_n3067_));
  NAND2_X1   g2425(.A1(new_n3067_), .A2(new_n3066_), .ZN(\result[100] ));
  NAND4_X1   g2426(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2486_), .A4(new_n2489_), .ZN(new_n3069_));
  OAI21_X1   g2427(.A1(new_n2702_), .A2(new_n2486_), .B(new_n2491_), .ZN(new_n3070_));
  NAND2_X1   g2428(.A1(new_n3070_), .A2(new_n3069_), .ZN(\result[101] ));
  NAND4_X1   g2429(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2465_), .A4(new_n2467_), .ZN(new_n3072_));
  OAI21_X1   g2430(.A1(new_n2702_), .A2(new_n2467_), .B(new_n2497_), .ZN(new_n3073_));
  NAND2_X1   g2431(.A1(new_n3073_), .A2(new_n3072_), .ZN(\result[102] ));
  NAND4_X1   g2432(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2469_), .A4(new_n2472_), .ZN(new_n3075_));
  OAI21_X1   g2433(.A1(new_n2702_), .A2(new_n2472_), .B(new_n2470_), .ZN(new_n3076_));
  NAND2_X1   g2434(.A1(new_n3076_), .A2(new_n3075_), .ZN(\result[103] ));
  NAND4_X1   g2435(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2529_), .A4(new_n2531_), .ZN(new_n3078_));
  OAI21_X1   g2436(.A1(new_n2702_), .A2(new_n2529_), .B(new_n2558_), .ZN(new_n3079_));
  NAND2_X1   g2437(.A1(new_n3079_), .A2(new_n3078_), .ZN(\result[104] ));
  NAND4_X1   g2438(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2523_), .A4(new_n2526_), .ZN(new_n3081_));
  OAI21_X1   g2439(.A1(new_n2702_), .A2(new_n2526_), .B(new_n2524_), .ZN(new_n3082_));
  NAND2_X1   g2440(.A1(new_n3082_), .A2(new_n3081_), .ZN(\result[105] ));
  NAND4_X1   g2441(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2510_), .A4(new_n2513_), .ZN(new_n3084_));
  OAI21_X1   g2442(.A1(new_n2702_), .A2(new_n2510_), .B(new_n2521_), .ZN(new_n3085_));
  NAND2_X1   g2443(.A1(new_n3085_), .A2(new_n3084_), .ZN(\result[106] ));
  NAND4_X1   g2444(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2515_), .A4(new_n2518_), .ZN(new_n3087_));
  INV_X1     g2445(.I(new_n2518_), .ZN(new_n3088_));
  OAI21_X1   g2446(.A1(new_n2702_), .A2(new_n2515_), .B(new_n3088_), .ZN(new_n3089_));
  NAND2_X1   g2447(.A1(new_n3089_), .A2(new_n3087_), .ZN(\result[107] ));
  NAND4_X1   g2448(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2553_), .A4(new_n2556_), .ZN(new_n3091_));
  OAI21_X1   g2449(.A1(new_n2702_), .A2(new_n2556_), .B(new_n2554_), .ZN(new_n3092_));
  NAND2_X1   g2450(.A1(new_n3092_), .A2(new_n3091_), .ZN(\result[108] ));
  NAND4_X1   g2451(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2547_), .A4(new_n2550_), .ZN(new_n3094_));
  OAI21_X1   g2452(.A1(new_n2702_), .A2(new_n2550_), .B(new_n2548_), .ZN(new_n3095_));
  NAND2_X1   g2453(.A1(new_n3095_), .A2(new_n3094_), .ZN(\result[109] ));
  NAND4_X1   g2454(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2536_), .A4(new_n2539_), .ZN(new_n3097_));
  OAI21_X1   g2455(.A1(new_n2702_), .A2(new_n2539_), .B(new_n2537_), .ZN(new_n3098_));
  NAND2_X1   g2456(.A1(new_n3098_), .A2(new_n3097_), .ZN(\result[110] ));
  NAND4_X1   g2457(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2541_), .A4(new_n2544_), .ZN(new_n3100_));
  OAI21_X1   g2458(.A1(new_n2702_), .A2(new_n2544_), .B(new_n2542_), .ZN(new_n3101_));
  NAND2_X1   g2459(.A1(new_n3101_), .A2(new_n3100_), .ZN(\result[111] ));
  NAND4_X1   g2460(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2592_), .A4(new_n2594_), .ZN(new_n3103_));
  OAI21_X1   g2461(.A1(new_n2702_), .A2(new_n2592_), .B(new_n2598_), .ZN(new_n3104_));
  NAND2_X1   g2462(.A1(new_n3104_), .A2(new_n3103_), .ZN(\result[112] ));
  NAND4_X1   g2463(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2586_), .A4(new_n2589_), .ZN(new_n3106_));
  OAI21_X1   g2464(.A1(new_n2702_), .A2(new_n2589_), .B(new_n2587_), .ZN(new_n3107_));
  NAND2_X1   g2465(.A1(new_n3107_), .A2(new_n3106_), .ZN(\result[113] ));
  NAND4_X1   g2466(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2575_), .A4(new_n2577_), .ZN(new_n3109_));
  OAI21_X1   g2467(.A1(new_n2702_), .A2(new_n2575_), .B(new_n2578_), .ZN(new_n3110_));
  NAND2_X1   g2468(.A1(new_n3110_), .A2(new_n3109_), .ZN(\result[114] ));
  NAND4_X1   g2469(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2580_), .A4(new_n2582_), .ZN(new_n3112_));
  OAI21_X1   g2470(.A1(new_n2702_), .A2(new_n2580_), .B(new_n2583_), .ZN(new_n3113_));
  NAND2_X1   g2471(.A1(new_n3113_), .A2(new_n3112_), .ZN(\result[115] ));
  NAND4_X1   g2472(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2620_), .A4(new_n2623_), .ZN(new_n3115_));
  OAI21_X1   g2473(.A1(new_n2702_), .A2(new_n2623_), .B(new_n2621_), .ZN(new_n3116_));
  NAND2_X1   g2474(.A1(new_n3116_), .A2(new_n3115_), .ZN(\result[116] ));
  NAND4_X1   g2475(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2625_), .A4(new_n2628_), .ZN(new_n3118_));
  OAI21_X1   g2476(.A1(new_n2702_), .A2(new_n2625_), .B(new_n2630_), .ZN(new_n3119_));
  NAND2_X1   g2477(.A1(new_n3119_), .A2(new_n3118_), .ZN(\result[117] ));
  NAND4_X1   g2478(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2604_), .A4(new_n2606_), .ZN(new_n3121_));
  OAI21_X1   g2479(.A1(new_n2702_), .A2(new_n2606_), .B(new_n2638_), .ZN(new_n3122_));
  NAND2_X1   g2480(.A1(new_n3122_), .A2(new_n3121_), .ZN(\result[118] ));
  NAND4_X1   g2481(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2608_), .A4(new_n2611_), .ZN(new_n3124_));
  OAI21_X1   g2482(.A1(new_n2702_), .A2(new_n2611_), .B(new_n2609_), .ZN(new_n3125_));
  NAND2_X1   g2483(.A1(new_n3125_), .A2(new_n3124_), .ZN(\result[119] ));
  NAND4_X1   g2484(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2656_), .A4(new_n2659_), .ZN(new_n3127_));
  OAI21_X1   g2485(.A1(new_n2702_), .A2(new_n2659_), .B(new_n2657_), .ZN(new_n3128_));
  NAND2_X1   g2486(.A1(new_n3128_), .A2(new_n3127_), .ZN(\result[120] ));
  NAND4_X1   g2487(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2661_), .A4(new_n2664_), .ZN(new_n3130_));
  OAI21_X1   g2488(.A1(new_n2702_), .A2(new_n2664_), .B(new_n2662_), .ZN(new_n3131_));
  NAND2_X1   g2489(.A1(new_n3131_), .A2(new_n3130_), .ZN(\result[121] ));
  NAND4_X1   g2490(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2643_), .A4(new_n2645_), .ZN(new_n3133_));
  INV_X1     g2491(.I(new_n2643_), .ZN(new_n3134_));
  OAI21_X1   g2492(.A1(new_n2702_), .A2(new_n2645_), .B(new_n3134_), .ZN(new_n3135_));
  NAND2_X1   g2493(.A1(new_n3135_), .A2(new_n3133_), .ZN(\result[122] ));
  NAND4_X1   g2494(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n2648_), .A4(new_n2651_), .ZN(new_n3137_));
  INV_X1     g2495(.I(new_n2648_), .ZN(new_n3138_));
  OAI21_X1   g2496(.A1(new_n2702_), .A2(new_n2651_), .B(new_n3138_), .ZN(new_n3139_));
  NAND2_X1   g2497(.A1(new_n3139_), .A2(new_n3137_), .ZN(\result[123] ));
  NAND4_X1   g2498(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1508_), .A4(new_n1556_), .ZN(new_n3141_));
  OAI21_X1   g2499(.A1(new_n2702_), .A2(new_n1508_), .B(new_n1557_), .ZN(new_n3142_));
  NAND2_X1   g2500(.A1(new_n3142_), .A2(new_n3141_), .ZN(\result[124] ));
  NAND4_X1   g2501(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1502_), .A4(new_n1504_), .ZN(new_n3144_));
  OAI21_X1   g2502(.A1(new_n2702_), .A2(new_n1502_), .B(new_n1505_), .ZN(new_n3145_));
  NAND2_X1   g2503(.A1(new_n3145_), .A2(new_n3144_), .ZN(\result[125] ));
  NAND4_X1   g2504(.A1(new_n2680_), .A2(new_n1451_), .A3(new_n1496_), .A4(new_n1498_), .ZN(new_n3147_));
  OAI21_X1   g2505(.A1(new_n2702_), .A2(new_n1496_), .B(new_n1499_), .ZN(new_n3148_));
  NAND2_X1   g2506(.A1(new_n3148_), .A2(new_n3147_), .ZN(\result[126] ));
  INV_X1     g2507(.I(new_n1450_), .ZN(new_n3150_));
  AOI21_X1   g2508(.A1(new_n2680_), .A2(new_n3150_), .B(new_n1449_), .ZN(\result[127] ));
  NAND4_X1   g2509(.A1(new_n2680_), .A2(new_n1046_), .A3(new_n1451_), .A4(new_n1568_), .ZN(new_n3152_));
  OAI21_X1   g2510(.A1(new_n2702_), .A2(new_n1568_), .B(new_n1554_), .ZN(new_n3153_));
  NAND2_X1   g2511(.A1(new_n3153_), .A2(new_n3152_), .ZN(\address[0] ));
  INV_X1     g2512(.I(new_n2702_), .ZN(\address[1] ));
endmodule


