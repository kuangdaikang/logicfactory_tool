// Benchmark "i4" written by ABC on Fri Feb 25 15:13:00 2022

module i4 ( 
    \V56(0) , \V28(0) , \V56(1) , \V28(1) , \V56(2) , \V28(2) , \V56(6) ,
    \V28(6) , \V56(10) , \V28(10) , \V56(14) , \V28(14) , \V56(18) ,
    \V28(18) , \V56(22) , \V28(22) , \V56(26) , \V28(26) , \V120(2) ,
    \V88(2) , \V120(6) , \V88(6) , \V120(10) , \V88(10) , \V120(14) ,
    \V88(14) , \V120(18) , \V88(18) , \V120(22) , \V88(22) , \V120(26) ,
    \V88(26) , \V120(30) , \V88(30) , \V132(2) , \V126(2) , \V144(0) ,
    \V28(3) , \V56(3) , \V144(1) , \V56(4) , \V28(4) , \V144(2) , \V28(5) ,
    \V56(5) , \V144(4) , \V28(7) , \V56(7) , \V144(5) , \V56(8) , \V28(8) ,
    \V144(6) , \V28(9) , \V56(9) , \V144(8) , \V28(11) , \V56(11) ,
    \V144(9) , \V56(12) , \V28(12) , \V144(10) , \V28(13) , \V56(13) ,
    \V144(12) , \V28(15) , \V56(15) , \V144(13) , \V56(16) , \V28(16) ,
    \V144(14) , \V28(17) , \V56(17) , \V156(0) , \V28(19) , \V56(19) ,
    \V156(1) , \V56(20) , \V28(20) , \V156(2) , \V28(21) , \V56(21) ,
    \V156(4) , \V28(23) , \V56(23) , \V156(5) , \V56(24) , \V28(24) ,
    \V156(6) , \V28(25) , \V56(25) , \V156(8) , \V28(27) , \V56(27) ,
    \V156(9) , \V120(0) , \V88(0) , \V156(10) , \V88(1) , \V120(1) ,
    \V156(12) , \V88(3) , \V120(3) , \V156(13) , \V120(4) , \V88(4) ,
    \V156(14) , \V88(5) , \V120(5) , \V168(0) , \V88(7) , \V120(7) ,
    \V168(1) , \V120(8) , \V88(8) , \V168(2) , \V88(9) , \V120(9) ,
    \V168(4) , \V88(11) , \V120(11) , \V168(5) , \V120(12) , \V88(12) ,
    \V168(6) , \V88(13) , \V120(13) , \V168(8) , \V88(15) , \V120(15) ,
    \V168(9) , \V120(16) , \V88(16) , \V168(10) , \V88(17) , \V120(17) ,
    \V168(12) , \V88(19) , \V120(19) , \V168(13) , \V120(20) , \V88(20) ,
    \V168(14) , \V88(21) , \V120(21) , \V180(0) , \V88(23) , \V120(23) ,
    \V180(1) , \V120(24) , \V88(24) , \V180(2) , \V88(25) , \V120(25) ,
    \V180(4) , \V88(27) , \V120(27) , \V180(5) , \V120(28) , \V88(28) ,
    \V180(6) , \V88(29) , \V120(29) , \V180(8) , \V88(31) , \V120(31) ,
    \V180(9) , \V132(0) , \V126(0) , \V180(10) , \V126(1) , \V132(1) ,
    \V180(12) , \V126(3) , \V132(3) , \V180(13) , \V132(4) , \V126(4) ,
    \V180(14) , \V126(5) , \V132(5) , \V183(0) , \V183(1) , \V183(2) ,
    \V186(0) , \V186(1) , \V186(2) , \V189(0) , \V189(1) , \V189(2) ,
    \V192(0) , \V192(1) , \V192(2) ,
    \V194(0) , \V194(1) , \V198(0) , \V198(1) , \V198(2) , \V198(3)   );
  input  \V56(0) , \V28(0) , \V56(1) , \V28(1) , \V56(2) , \V28(2) ,
    \V56(6) , \V28(6) , \V56(10) , \V28(10) , \V56(14) , \V28(14) ,
    \V56(18) , \V28(18) , \V56(22) , \V28(22) , \V56(26) , \V28(26) ,
    \V120(2) , \V88(2) , \V120(6) , \V88(6) , \V120(10) , \V88(10) ,
    \V120(14) , \V88(14) , \V120(18) , \V88(18) , \V120(22) , \V88(22) ,
    \V120(26) , \V88(26) , \V120(30) , \V88(30) , \V132(2) , \V126(2) ,
    \V144(0) , \V28(3) , \V56(3) , \V144(1) , \V56(4) , \V28(4) ,
    \V144(2) , \V28(5) , \V56(5) , \V144(4) , \V28(7) , \V56(7) ,
    \V144(5) , \V56(8) , \V28(8) , \V144(6) , \V28(9) , \V56(9) ,
    \V144(8) , \V28(11) , \V56(11) , \V144(9) , \V56(12) , \V28(12) ,
    \V144(10) , \V28(13) , \V56(13) , \V144(12) , \V28(15) , \V56(15) ,
    \V144(13) , \V56(16) , \V28(16) , \V144(14) , \V28(17) , \V56(17) ,
    \V156(0) , \V28(19) , \V56(19) , \V156(1) , \V56(20) , \V28(20) ,
    \V156(2) , \V28(21) , \V56(21) , \V156(4) , \V28(23) , \V56(23) ,
    \V156(5) , \V56(24) , \V28(24) , \V156(6) , \V28(25) , \V56(25) ,
    \V156(8) , \V28(27) , \V56(27) , \V156(9) , \V120(0) , \V88(0) ,
    \V156(10) , \V88(1) , \V120(1) , \V156(12) , \V88(3) , \V120(3) ,
    \V156(13) , \V120(4) , \V88(4) , \V156(14) , \V88(5) , \V120(5) ,
    \V168(0) , \V88(7) , \V120(7) , \V168(1) , \V120(8) , \V88(8) ,
    \V168(2) , \V88(9) , \V120(9) , \V168(4) , \V88(11) , \V120(11) ,
    \V168(5) , \V120(12) , \V88(12) , \V168(6) , \V88(13) , \V120(13) ,
    \V168(8) , \V88(15) , \V120(15) , \V168(9) , \V120(16) , \V88(16) ,
    \V168(10) , \V88(17) , \V120(17) , \V168(12) , \V88(19) , \V120(19) ,
    \V168(13) , \V120(20) , \V88(20) , \V168(14) , \V88(21) , \V120(21) ,
    \V180(0) , \V88(23) , \V120(23) , \V180(1) , \V120(24) , \V88(24) ,
    \V180(2) , \V88(25) , \V120(25) , \V180(4) , \V88(27) , \V120(27) ,
    \V180(5) , \V120(28) , \V88(28) , \V180(6) , \V88(29) , \V120(29) ,
    \V180(8) , \V88(31) , \V120(31) , \V180(9) , \V132(0) , \V126(0) ,
    \V180(10) , \V126(1) , \V132(1) , \V180(12) , \V126(3) , \V132(3) ,
    \V180(13) , \V132(4) , \V126(4) , \V180(14) , \V126(5) , \V132(5) ,
    \V183(0) , \V183(1) , \V183(2) , \V186(0) , \V186(1) , \V186(2) ,
    \V189(0) , \V189(1) , \V189(2) , \V192(0) , \V192(1) , \V192(2) ;
  output \V194(0) , \V194(1) , \V198(0) , \V198(1) , \V198(2) , \V198(3) ;
  wire new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_;
  assign \V194(0)  = \V56(0)  & \V28(0) ;
  assign \V194(1)  = \V56(1)  & \V28(1) ;
  assign new_n201_ = \V144(12)  & \V144(14) ;
  assign new_n202_ = \V28(17)  & new_n201_;
  assign new_n203_ = \V56(17)  & new_n202_;
  assign new_n204_ = \V144(13)  & new_n203_;
  assign new_n205_ = \V144(12)  & \V28(15) ;
  assign new_n206_ = \V56(15)  & new_n205_;
  assign new_n207_ = \V56(14)  & \V28(14) ;
  assign new_n208_ = \V144(13)  & \V56(16) ;
  assign new_n209_ = \V28(16)  & new_n208_;
  assign new_n210_ = \V144(12)  & new_n209_;
  assign new_n211_ = ~new_n207_ & ~new_n210_;
  assign new_n212_ = ~new_n204_ & ~new_n206_;
  assign new_n213_ = new_n211_ & new_n212_;
  assign new_n214_ = \V183(0)  & \V183(2) ;
  assign new_n215_ = ~new_n213_ & new_n214_;
  assign new_n216_ = \V183(1)  & new_n215_;
  assign new_n217_ = \V144(4)  & \V144(6) ;
  assign new_n218_ = \V28(9)  & new_n217_;
  assign new_n219_ = \V56(9)  & new_n218_;
  assign new_n220_ = \V144(5)  & new_n219_;
  assign new_n221_ = \V144(4)  & \V28(7) ;
  assign new_n222_ = \V56(7)  & new_n221_;
  assign new_n223_ = \V56(6)  & \V28(6) ;
  assign new_n224_ = \V144(5)  & \V56(8) ;
  assign new_n225_ = \V28(8)  & new_n224_;
  assign new_n226_ = \V144(4)  & new_n225_;
  assign new_n227_ = ~new_n223_ & ~new_n226_;
  assign new_n228_ = ~new_n220_ & ~new_n222_;
  assign new_n229_ = new_n227_ & new_n228_;
  assign new_n230_ = \V183(0)  & ~new_n229_;
  assign new_n231_ = \V144(1)  & \V56(4) ;
  assign new_n232_ = \V28(4)  & new_n231_;
  assign new_n233_ = \V144(0)  & new_n232_;
  assign new_n234_ = \V56(2)  & \V28(2) ;
  assign new_n235_ = \V144(0)  & \V28(3) ;
  assign new_n236_ = \V56(3)  & new_n235_;
  assign new_n237_ = \V144(0)  & \V144(2) ;
  assign new_n238_ = \V28(5)  & new_n237_;
  assign new_n239_ = \V56(5)  & new_n238_;
  assign new_n240_ = \V144(1)  & new_n239_;
  assign new_n241_ = \V144(8)  & \V144(10) ;
  assign new_n242_ = \V28(13)  & new_n241_;
  assign new_n243_ = \V56(13)  & new_n242_;
  assign new_n244_ = \V144(9)  & new_n243_;
  assign new_n245_ = \V144(8)  & \V28(11) ;
  assign new_n246_ = \V56(11)  & new_n245_;
  assign new_n247_ = \V56(10)  & \V28(10) ;
  assign new_n248_ = \V144(9)  & \V56(12) ;
  assign new_n249_ = \V28(12)  & new_n248_;
  assign new_n250_ = \V144(8)  & new_n249_;
  assign new_n251_ = ~new_n247_ & ~new_n250_;
  assign new_n252_ = ~new_n244_ & ~new_n246_;
  assign new_n253_ = new_n251_ & new_n252_;
  assign new_n254_ = \V183(1)  & ~new_n253_;
  assign new_n255_ = \V183(0)  & new_n254_;
  assign new_n256_ = ~new_n233_ & ~new_n234_;
  assign new_n257_ = ~new_n216_ & ~new_n230_;
  assign new_n258_ = new_n256_ & new_n257_;
  assign new_n259_ = ~new_n236_ & ~new_n240_;
  assign new_n260_ = ~new_n255_ & new_n259_;
  assign \V198(0)  = ~new_n258_ | ~new_n260_;
  assign new_n262_ = \V156(12)  & \V156(14) ;
  assign new_n263_ = \V88(5)  & new_n262_;
  assign new_n264_ = \V120(5)  & new_n263_;
  assign new_n265_ = \V156(13)  & new_n264_;
  assign new_n266_ = \V156(12)  & \V88(3) ;
  assign new_n267_ = \V120(3)  & new_n266_;
  assign new_n268_ = \V120(2)  & \V88(2) ;
  assign new_n269_ = \V156(13)  & \V120(4) ;
  assign new_n270_ = \V88(4)  & new_n269_;
  assign new_n271_ = \V156(12)  & new_n270_;
  assign new_n272_ = ~new_n268_ & ~new_n271_;
  assign new_n273_ = ~new_n265_ & ~new_n267_;
  assign new_n274_ = new_n272_ & new_n273_;
  assign new_n275_ = \V186(0)  & \V186(2) ;
  assign new_n276_ = ~new_n274_ & new_n275_;
  assign new_n277_ = \V186(1)  & new_n276_;
  assign new_n278_ = \V156(4)  & \V156(6) ;
  assign new_n279_ = \V28(25)  & new_n278_;
  assign new_n280_ = \V56(25)  & new_n279_;
  assign new_n281_ = \V156(5)  & new_n280_;
  assign new_n282_ = \V156(4)  & \V28(23) ;
  assign new_n283_ = \V56(23)  & new_n282_;
  assign new_n284_ = \V56(22)  & \V28(22) ;
  assign new_n285_ = \V156(5)  & \V56(24) ;
  assign new_n286_ = \V28(24)  & new_n285_;
  assign new_n287_ = \V156(4)  & new_n286_;
  assign new_n288_ = ~new_n284_ & ~new_n287_;
  assign new_n289_ = ~new_n281_ & ~new_n283_;
  assign new_n290_ = new_n288_ & new_n289_;
  assign new_n291_ = \V186(0)  & ~new_n290_;
  assign new_n292_ = \V156(1)  & \V56(20) ;
  assign new_n293_ = \V28(20)  & new_n292_;
  assign new_n294_ = \V156(0)  & new_n293_;
  assign new_n295_ = \V56(18)  & \V28(18) ;
  assign new_n296_ = \V156(0)  & \V28(19) ;
  assign new_n297_ = \V56(19)  & new_n296_;
  assign new_n298_ = \V156(0)  & \V156(2) ;
  assign new_n299_ = \V28(21)  & new_n298_;
  assign new_n300_ = \V56(21)  & new_n299_;
  assign new_n301_ = \V156(1)  & new_n300_;
  assign new_n302_ = \V156(8)  & \V156(10) ;
  assign new_n303_ = \V88(1)  & new_n302_;
  assign new_n304_ = \V120(1)  & new_n303_;
  assign new_n305_ = \V156(9)  & new_n304_;
  assign new_n306_ = \V156(8)  & \V28(27) ;
  assign new_n307_ = \V56(27)  & new_n306_;
  assign new_n308_ = \V56(26)  & \V28(26) ;
  assign new_n309_ = \V156(9)  & \V120(0) ;
  assign new_n310_ = \V88(0)  & new_n309_;
  assign new_n311_ = \V156(8)  & new_n310_;
  assign new_n312_ = ~new_n308_ & ~new_n311_;
  assign new_n313_ = ~new_n305_ & ~new_n307_;
  assign new_n314_ = new_n312_ & new_n313_;
  assign new_n315_ = \V186(1)  & ~new_n314_;
  assign new_n316_ = \V186(0)  & new_n315_;
  assign new_n317_ = ~new_n294_ & ~new_n295_;
  assign new_n318_ = ~new_n277_ & ~new_n291_;
  assign new_n319_ = new_n317_ & new_n318_;
  assign new_n320_ = ~new_n297_ & ~new_n301_;
  assign new_n321_ = ~new_n316_ & new_n320_;
  assign \V198(1)  = ~new_n319_ | ~new_n321_;
  assign new_n323_ = \V168(12)  & \V168(14) ;
  assign new_n324_ = \V88(21)  & new_n323_;
  assign new_n325_ = \V120(21)  & new_n324_;
  assign new_n326_ = \V168(13)  & new_n325_;
  assign new_n327_ = \V168(12)  & \V88(19) ;
  assign new_n328_ = \V120(19)  & new_n327_;
  assign new_n329_ = \V120(18)  & \V88(18) ;
  assign new_n330_ = \V168(13)  & \V120(20) ;
  assign new_n331_ = \V88(20)  & new_n330_;
  assign new_n332_ = \V168(12)  & new_n331_;
  assign new_n333_ = ~new_n329_ & ~new_n332_;
  assign new_n334_ = ~new_n326_ & ~new_n328_;
  assign new_n335_ = new_n333_ & new_n334_;
  assign new_n336_ = \V189(0)  & \V189(2) ;
  assign new_n337_ = ~new_n335_ & new_n336_;
  assign new_n338_ = \V189(1)  & new_n337_;
  assign new_n339_ = \V168(4)  & \V168(6) ;
  assign new_n340_ = \V88(13)  & new_n339_;
  assign new_n341_ = \V120(13)  & new_n340_;
  assign new_n342_ = \V168(5)  & new_n341_;
  assign new_n343_ = \V168(4)  & \V88(11) ;
  assign new_n344_ = \V120(11)  & new_n343_;
  assign new_n345_ = \V120(10)  & \V88(10) ;
  assign new_n346_ = \V168(5)  & \V120(12) ;
  assign new_n347_ = \V88(12)  & new_n346_;
  assign new_n348_ = \V168(4)  & new_n347_;
  assign new_n349_ = ~new_n345_ & ~new_n348_;
  assign new_n350_ = ~new_n342_ & ~new_n344_;
  assign new_n351_ = new_n349_ & new_n350_;
  assign new_n352_ = \V189(0)  & ~new_n351_;
  assign new_n353_ = \V168(1)  & \V120(8) ;
  assign new_n354_ = \V88(8)  & new_n353_;
  assign new_n355_ = \V168(0)  & new_n354_;
  assign new_n356_ = \V120(6)  & \V88(6) ;
  assign new_n357_ = \V168(0)  & \V88(7) ;
  assign new_n358_ = \V120(7)  & new_n357_;
  assign new_n359_ = \V168(0)  & \V168(2) ;
  assign new_n360_ = \V88(9)  & new_n359_;
  assign new_n361_ = \V120(9)  & new_n360_;
  assign new_n362_ = \V168(1)  & new_n361_;
  assign new_n363_ = \V168(8)  & \V168(10) ;
  assign new_n364_ = \V88(17)  & new_n363_;
  assign new_n365_ = \V120(17)  & new_n364_;
  assign new_n366_ = \V168(9)  & new_n365_;
  assign new_n367_ = \V168(8)  & \V88(15) ;
  assign new_n368_ = \V120(15)  & new_n367_;
  assign new_n369_ = \V120(14)  & \V88(14) ;
  assign new_n370_ = \V168(9)  & \V120(16) ;
  assign new_n371_ = \V88(16)  & new_n370_;
  assign new_n372_ = \V168(8)  & new_n371_;
  assign new_n373_ = ~new_n369_ & ~new_n372_;
  assign new_n374_ = ~new_n366_ & ~new_n368_;
  assign new_n375_ = new_n373_ & new_n374_;
  assign new_n376_ = \V189(1)  & ~new_n375_;
  assign new_n377_ = \V189(0)  & new_n376_;
  assign new_n378_ = ~new_n355_ & ~new_n356_;
  assign new_n379_ = ~new_n338_ & ~new_n352_;
  assign new_n380_ = new_n378_ & new_n379_;
  assign new_n381_ = ~new_n358_ & ~new_n362_;
  assign new_n382_ = ~new_n377_ & new_n381_;
  assign \V198(2)  = ~new_n380_ | ~new_n382_;
  assign new_n384_ = \V180(12)  & \V180(14) ;
  assign new_n385_ = \V126(5)  & new_n384_;
  assign new_n386_ = \V132(5)  & new_n385_;
  assign new_n387_ = \V180(13)  & new_n386_;
  assign new_n388_ = \V180(12)  & \V126(3) ;
  assign new_n389_ = \V132(3)  & new_n388_;
  assign new_n390_ = \V132(2)  & \V126(2) ;
  assign new_n391_ = \V180(13)  & \V132(4) ;
  assign new_n392_ = \V126(4)  & new_n391_;
  assign new_n393_ = \V180(12)  & new_n392_;
  assign new_n394_ = ~new_n390_ & ~new_n393_;
  assign new_n395_ = ~new_n387_ & ~new_n389_;
  assign new_n396_ = new_n394_ & new_n395_;
  assign new_n397_ = \V192(0)  & \V192(2) ;
  assign new_n398_ = ~new_n396_ & new_n397_;
  assign new_n399_ = \V192(1)  & new_n398_;
  assign new_n400_ = \V180(4)  & \V180(6) ;
  assign new_n401_ = \V88(29)  & new_n400_;
  assign new_n402_ = \V120(29)  & new_n401_;
  assign new_n403_ = \V180(5)  & new_n402_;
  assign new_n404_ = \V180(4)  & \V88(27) ;
  assign new_n405_ = \V120(27)  & new_n404_;
  assign new_n406_ = \V120(26)  & \V88(26) ;
  assign new_n407_ = \V180(5)  & \V120(28) ;
  assign new_n408_ = \V88(28)  & new_n407_;
  assign new_n409_ = \V180(4)  & new_n408_;
  assign new_n410_ = ~new_n406_ & ~new_n409_;
  assign new_n411_ = ~new_n403_ & ~new_n405_;
  assign new_n412_ = new_n410_ & new_n411_;
  assign new_n413_ = \V192(0)  & ~new_n412_;
  assign new_n414_ = \V180(1)  & \V120(24) ;
  assign new_n415_ = \V88(24)  & new_n414_;
  assign new_n416_ = \V180(0)  & new_n415_;
  assign new_n417_ = \V120(22)  & \V88(22) ;
  assign new_n418_ = \V180(0)  & \V88(23) ;
  assign new_n419_ = \V120(23)  & new_n418_;
  assign new_n420_ = \V180(0)  & \V180(2) ;
  assign new_n421_ = \V88(25)  & new_n420_;
  assign new_n422_ = \V120(25)  & new_n421_;
  assign new_n423_ = \V180(1)  & new_n422_;
  assign new_n424_ = \V180(8)  & \V180(10) ;
  assign new_n425_ = \V126(1)  & new_n424_;
  assign new_n426_ = \V132(1)  & new_n425_;
  assign new_n427_ = \V180(9)  & new_n426_;
  assign new_n428_ = \V180(8)  & \V88(31) ;
  assign new_n429_ = \V120(31)  & new_n428_;
  assign new_n430_ = \V120(30)  & \V88(30) ;
  assign new_n431_ = \V180(9)  & \V132(0) ;
  assign new_n432_ = \V126(0)  & new_n431_;
  assign new_n433_ = \V180(8)  & new_n432_;
  assign new_n434_ = ~new_n430_ & ~new_n433_;
  assign new_n435_ = ~new_n427_ & ~new_n429_;
  assign new_n436_ = new_n434_ & new_n435_;
  assign new_n437_ = \V192(1)  & ~new_n436_;
  assign new_n438_ = \V192(0)  & new_n437_;
  assign new_n439_ = ~new_n416_ & ~new_n417_;
  assign new_n440_ = ~new_n399_ & ~new_n413_;
  assign new_n441_ = new_n439_ & new_n440_;
  assign new_n442_ = ~new_n419_ & ~new_n423_;
  assign new_n443_ = ~new_n438_ & new_n442_;
  assign \V198(3)  = ~new_n441_ | ~new_n443_;
endmodule


