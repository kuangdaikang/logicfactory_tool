// Benchmark "top" written by ABC on Fri Feb 25 15:09:03 2022

module dec ( 
    \count[0] , \count[1] , \count[2] , \count[3] , \count[4] , \count[5] ,
    \count[6] , \count[7] ,
    \selectp1[0] , \selectp1[1] , \selectp1[2] , \selectp1[3] ,
    \selectp1[4] , \selectp1[5] , \selectp1[6] , \selectp1[7] ,
    \selectp1[8] , \selectp1[9] , \selectp1[10] , \selectp1[11] ,
    \selectp1[12] , \selectp1[13] , \selectp1[14] , \selectp1[15] ,
    \selectp1[16] , \selectp1[17] , \selectp1[18] , \selectp1[19] ,
    \selectp1[20] , \selectp1[21] , \selectp1[22] , \selectp1[23] ,
    \selectp1[24] , \selectp1[25] , \selectp1[26] , \selectp1[27] ,
    \selectp1[28] , \selectp1[29] , \selectp1[30] , \selectp1[31] ,
    \selectp1[32] , \selectp1[33] , \selectp1[34] , \selectp1[35] ,
    \selectp1[36] , \selectp1[37] , \selectp1[38] , \selectp1[39] ,
    \selectp1[40] , \selectp1[41] , \selectp1[42] , \selectp1[43] ,
    \selectp1[44] , \selectp1[45] , \selectp1[46] , \selectp1[47] ,
    \selectp1[48] , \selectp1[49] , \selectp1[50] , \selectp1[51] ,
    \selectp1[52] , \selectp1[53] , \selectp1[54] , \selectp1[55] ,
    \selectp1[56] , \selectp1[57] , \selectp1[58] , \selectp1[59] ,
    \selectp1[60] , \selectp1[61] , \selectp1[62] , \selectp1[63] ,
    \selectp1[64] , \selectp1[65] , \selectp1[66] , \selectp1[67] ,
    \selectp1[68] , \selectp1[69] , \selectp1[70] , \selectp1[71] ,
    \selectp1[72] , \selectp1[73] , \selectp1[74] , \selectp1[75] ,
    \selectp1[76] , \selectp1[77] , \selectp1[78] , \selectp1[79] ,
    \selectp1[80] , \selectp1[81] , \selectp1[82] , \selectp1[83] ,
    \selectp1[84] , \selectp1[85] , \selectp1[86] , \selectp1[87] ,
    \selectp1[88] , \selectp1[89] , \selectp1[90] , \selectp1[91] ,
    \selectp1[92] , \selectp1[93] , \selectp1[94] , \selectp1[95] ,
    \selectp1[96] , \selectp1[97] , \selectp1[98] , \selectp1[99] ,
    \selectp1[100] , \selectp1[101] , \selectp1[102] , \selectp1[103] ,
    \selectp1[104] , \selectp1[105] , \selectp1[106] , \selectp1[107] ,
    \selectp1[108] , \selectp1[109] , \selectp1[110] , \selectp1[111] ,
    \selectp1[112] , \selectp1[113] , \selectp1[114] , \selectp1[115] ,
    \selectp1[116] , \selectp1[117] , \selectp1[118] , \selectp1[119] ,
    \selectp1[120] , \selectp1[121] , \selectp1[122] , \selectp1[123] ,
    \selectp1[124] , \selectp1[125] , \selectp1[126] , \selectp1[127] ,
    \selectp2[0] , \selectp2[1] , \selectp2[2] , \selectp2[3] ,
    \selectp2[4] , \selectp2[5] , \selectp2[6] , \selectp2[7] ,
    \selectp2[8] , \selectp2[9] , \selectp2[10] , \selectp2[11] ,
    \selectp2[12] , \selectp2[13] , \selectp2[14] , \selectp2[15] ,
    \selectp2[16] , \selectp2[17] , \selectp2[18] , \selectp2[19] ,
    \selectp2[20] , \selectp2[21] , \selectp2[22] , \selectp2[23] ,
    \selectp2[24] , \selectp2[25] , \selectp2[26] , \selectp2[27] ,
    \selectp2[28] , \selectp2[29] , \selectp2[30] , \selectp2[31] ,
    \selectp2[32] , \selectp2[33] , \selectp2[34] , \selectp2[35] ,
    \selectp2[36] , \selectp2[37] , \selectp2[38] , \selectp2[39] ,
    \selectp2[40] , \selectp2[41] , \selectp2[42] , \selectp2[43] ,
    \selectp2[44] , \selectp2[45] , \selectp2[46] , \selectp2[47] ,
    \selectp2[48] , \selectp2[49] , \selectp2[50] , \selectp2[51] ,
    \selectp2[52] , \selectp2[53] , \selectp2[54] , \selectp2[55] ,
    \selectp2[56] , \selectp2[57] , \selectp2[58] , \selectp2[59] ,
    \selectp2[60] , \selectp2[61] , \selectp2[62] , \selectp2[63] ,
    \selectp2[64] , \selectp2[65] , \selectp2[66] , \selectp2[67] ,
    \selectp2[68] , \selectp2[69] , \selectp2[70] , \selectp2[71] ,
    \selectp2[72] , \selectp2[73] , \selectp2[74] , \selectp2[75] ,
    \selectp2[76] , \selectp2[77] , \selectp2[78] , \selectp2[79] ,
    \selectp2[80] , \selectp2[81] , \selectp2[82] , \selectp2[83] ,
    \selectp2[84] , \selectp2[85] , \selectp2[86] , \selectp2[87] ,
    \selectp2[88] , \selectp2[89] , \selectp2[90] , \selectp2[91] ,
    \selectp2[92] , \selectp2[93] , \selectp2[94] , \selectp2[95] ,
    \selectp2[96] , \selectp2[97] , \selectp2[98] , \selectp2[99] ,
    \selectp2[100] , \selectp2[101] , \selectp2[102] , \selectp2[103] ,
    \selectp2[104] , \selectp2[105] , \selectp2[106] , \selectp2[107] ,
    \selectp2[108] , \selectp2[109] , \selectp2[110] , \selectp2[111] ,
    \selectp2[112] , \selectp2[113] , \selectp2[114] , \selectp2[115] ,
    \selectp2[116] , \selectp2[117] , \selectp2[118] , \selectp2[119] ,
    \selectp2[120] , \selectp2[121] , \selectp2[122] , \selectp2[123] ,
    \selectp2[124] , \selectp2[125] , \selectp2[126] , \selectp2[127]   );
  input  \count[0] , \count[1] , \count[2] , \count[3] , \count[4] ,
    \count[5] , \count[6] , \count[7] ;
  output \selectp1[0] , \selectp1[1] , \selectp1[2] , \selectp1[3] ,
    \selectp1[4] , \selectp1[5] , \selectp1[6] , \selectp1[7] ,
    \selectp1[8] , \selectp1[9] , \selectp1[10] , \selectp1[11] ,
    \selectp1[12] , \selectp1[13] , \selectp1[14] , \selectp1[15] ,
    \selectp1[16] , \selectp1[17] , \selectp1[18] , \selectp1[19] ,
    \selectp1[20] , \selectp1[21] , \selectp1[22] , \selectp1[23] ,
    \selectp1[24] , \selectp1[25] , \selectp1[26] , \selectp1[27] ,
    \selectp1[28] , \selectp1[29] , \selectp1[30] , \selectp1[31] ,
    \selectp1[32] , \selectp1[33] , \selectp1[34] , \selectp1[35] ,
    \selectp1[36] , \selectp1[37] , \selectp1[38] , \selectp1[39] ,
    \selectp1[40] , \selectp1[41] , \selectp1[42] , \selectp1[43] ,
    \selectp1[44] , \selectp1[45] , \selectp1[46] , \selectp1[47] ,
    \selectp1[48] , \selectp1[49] , \selectp1[50] , \selectp1[51] ,
    \selectp1[52] , \selectp1[53] , \selectp1[54] , \selectp1[55] ,
    \selectp1[56] , \selectp1[57] , \selectp1[58] , \selectp1[59] ,
    \selectp1[60] , \selectp1[61] , \selectp1[62] , \selectp1[63] ,
    \selectp1[64] , \selectp1[65] , \selectp1[66] , \selectp1[67] ,
    \selectp1[68] , \selectp1[69] , \selectp1[70] , \selectp1[71] ,
    \selectp1[72] , \selectp1[73] , \selectp1[74] , \selectp1[75] ,
    \selectp1[76] , \selectp1[77] , \selectp1[78] , \selectp1[79] ,
    \selectp1[80] , \selectp1[81] , \selectp1[82] , \selectp1[83] ,
    \selectp1[84] , \selectp1[85] , \selectp1[86] , \selectp1[87] ,
    \selectp1[88] , \selectp1[89] , \selectp1[90] , \selectp1[91] ,
    \selectp1[92] , \selectp1[93] , \selectp1[94] , \selectp1[95] ,
    \selectp1[96] , \selectp1[97] , \selectp1[98] , \selectp1[99] ,
    \selectp1[100] , \selectp1[101] , \selectp1[102] , \selectp1[103] ,
    \selectp1[104] , \selectp1[105] , \selectp1[106] , \selectp1[107] ,
    \selectp1[108] , \selectp1[109] , \selectp1[110] , \selectp1[111] ,
    \selectp1[112] , \selectp1[113] , \selectp1[114] , \selectp1[115] ,
    \selectp1[116] , \selectp1[117] , \selectp1[118] , \selectp1[119] ,
    \selectp1[120] , \selectp1[121] , \selectp1[122] , \selectp1[123] ,
    \selectp1[124] , \selectp1[125] , \selectp1[126] , \selectp1[127] ,
    \selectp2[0] , \selectp2[1] , \selectp2[2] , \selectp2[3] ,
    \selectp2[4] , \selectp2[5] , \selectp2[6] , \selectp2[7] ,
    \selectp2[8] , \selectp2[9] , \selectp2[10] , \selectp2[11] ,
    \selectp2[12] , \selectp2[13] , \selectp2[14] , \selectp2[15] ,
    \selectp2[16] , \selectp2[17] , \selectp2[18] , \selectp2[19] ,
    \selectp2[20] , \selectp2[21] , \selectp2[22] , \selectp2[23] ,
    \selectp2[24] , \selectp2[25] , \selectp2[26] , \selectp2[27] ,
    \selectp2[28] , \selectp2[29] , \selectp2[30] , \selectp2[31] ,
    \selectp2[32] , \selectp2[33] , \selectp2[34] , \selectp2[35] ,
    \selectp2[36] , \selectp2[37] , \selectp2[38] , \selectp2[39] ,
    \selectp2[40] , \selectp2[41] , \selectp2[42] , \selectp2[43] ,
    \selectp2[44] , \selectp2[45] , \selectp2[46] , \selectp2[47] ,
    \selectp2[48] , \selectp2[49] , \selectp2[50] , \selectp2[51] ,
    \selectp2[52] , \selectp2[53] , \selectp2[54] , \selectp2[55] ,
    \selectp2[56] , \selectp2[57] , \selectp2[58] , \selectp2[59] ,
    \selectp2[60] , \selectp2[61] , \selectp2[62] , \selectp2[63] ,
    \selectp2[64] , \selectp2[65] , \selectp2[66] , \selectp2[67] ,
    \selectp2[68] , \selectp2[69] , \selectp2[70] , \selectp2[71] ,
    \selectp2[72] , \selectp2[73] , \selectp2[74] , \selectp2[75] ,
    \selectp2[76] , \selectp2[77] , \selectp2[78] , \selectp2[79] ,
    \selectp2[80] , \selectp2[81] , \selectp2[82] , \selectp2[83] ,
    \selectp2[84] , \selectp2[85] , \selectp2[86] , \selectp2[87] ,
    \selectp2[88] , \selectp2[89] , \selectp2[90] , \selectp2[91] ,
    \selectp2[92] , \selectp2[93] , \selectp2[94] , \selectp2[95] ,
    \selectp2[96] , \selectp2[97] , \selectp2[98] , \selectp2[99] ,
    \selectp2[100] , \selectp2[101] , \selectp2[102] , \selectp2[103] ,
    \selectp2[104] , \selectp2[105] , \selectp2[106] , \selectp2[107] ,
    \selectp2[108] , \selectp2[109] , \selectp2[110] , \selectp2[111] ,
    \selectp2[112] , \selectp2[113] , \selectp2[114] , \selectp2[115] ,
    \selectp2[116] , \selectp2[117] , \selectp2[118] , \selectp2[119] ,
    \selectp2[120] , \selectp2[121] , \selectp2[122] , \selectp2[123] ,
    \selectp2[124] , \selectp2[125] , \selectp2[126] , \selectp2[127] ;
  wire new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n272_, new_n273_, new_n275_, new_n276_, new_n278_, new_n280_,
    new_n281_, new_n283_, new_n284_, new_n286_, new_n288_, new_n290_,
    new_n291_, new_n293_, new_n295_, new_n296_, new_n298_, new_n300_,
    new_n302_, new_n304_, new_n306_, new_n308_, new_n309_, new_n326_,
    new_n327_, new_n344_, new_n345_, new_n362_, new_n363_, new_n380_,
    new_n397_, new_n414_, new_n431_, new_n432_, new_n449_, new_n466_,
    new_n483_, new_n500_, new_n501_, new_n518_, new_n535_, new_n552_;
  assign new_n265_ = ~\count[4]  & ~\count[5] ;
  assign new_n266_ = ~\count[6]  & \count[7] ;
  assign new_n267_ = new_n265_ & new_n266_;
  assign new_n268_ = ~\count[0]  & ~\count[2] ;
  assign new_n269_ = ~\count[1]  & ~\count[3] ;
  assign new_n270_ = new_n268_ & new_n269_;
  assign \selectp1[0]  = new_n267_ & new_n270_;
  assign new_n272_ = \count[0]  & ~\count[2] ;
  assign new_n273_ = new_n269_ & new_n272_;
  assign \selectp1[1]  = new_n267_ & new_n273_;
  assign new_n275_ = \count[1]  & ~\count[3] ;
  assign new_n276_ = new_n268_ & new_n275_;
  assign \selectp1[2]  = new_n267_ & new_n276_;
  assign new_n278_ = new_n272_ & new_n275_;
  assign \selectp1[3]  = new_n267_ & new_n278_;
  assign new_n280_ = ~\count[0]  & \count[2] ;
  assign new_n281_ = new_n269_ & new_n280_;
  assign \selectp1[4]  = new_n267_ & new_n281_;
  assign new_n283_ = \count[0]  & \count[2] ;
  assign new_n284_ = new_n269_ & new_n283_;
  assign \selectp1[5]  = new_n267_ & new_n284_;
  assign new_n286_ = new_n275_ & new_n280_;
  assign \selectp1[6]  = new_n267_ & new_n286_;
  assign new_n288_ = new_n275_ & new_n283_;
  assign \selectp1[7]  = new_n267_ & new_n288_;
  assign new_n290_ = ~\count[1]  & \count[3] ;
  assign new_n291_ = new_n268_ & new_n290_;
  assign \selectp1[8]  = new_n267_ & new_n291_;
  assign new_n293_ = new_n272_ & new_n290_;
  assign \selectp1[9]  = new_n267_ & new_n293_;
  assign new_n295_ = \count[1]  & \count[3] ;
  assign new_n296_ = new_n268_ & new_n295_;
  assign \selectp1[10]  = new_n267_ & new_n296_;
  assign new_n298_ = new_n272_ & new_n295_;
  assign \selectp1[11]  = new_n267_ & new_n298_;
  assign new_n300_ = new_n280_ & new_n290_;
  assign \selectp1[12]  = new_n267_ & new_n300_;
  assign new_n302_ = new_n283_ & new_n290_;
  assign \selectp1[13]  = new_n267_ & new_n302_;
  assign new_n304_ = new_n280_ & new_n295_;
  assign \selectp1[14]  = new_n267_ & new_n304_;
  assign new_n306_ = new_n283_ & new_n295_;
  assign \selectp1[15]  = new_n267_ & new_n306_;
  assign new_n308_ = \count[4]  & ~\count[5] ;
  assign new_n309_ = new_n266_ & new_n308_;
  assign \selectp1[16]  = new_n270_ & new_n309_;
  assign \selectp1[17]  = new_n273_ & new_n309_;
  assign \selectp1[18]  = new_n276_ & new_n309_;
  assign \selectp1[19]  = new_n278_ & new_n309_;
  assign \selectp1[20]  = new_n281_ & new_n309_;
  assign \selectp1[21]  = new_n284_ & new_n309_;
  assign \selectp1[22]  = new_n286_ & new_n309_;
  assign \selectp1[23]  = new_n288_ & new_n309_;
  assign \selectp1[24]  = new_n291_ & new_n309_;
  assign \selectp1[25]  = new_n293_ & new_n309_;
  assign \selectp1[26]  = new_n296_ & new_n309_;
  assign \selectp1[27]  = new_n298_ & new_n309_;
  assign \selectp1[28]  = new_n300_ & new_n309_;
  assign \selectp1[29]  = new_n302_ & new_n309_;
  assign \selectp1[30]  = new_n304_ & new_n309_;
  assign \selectp1[31]  = new_n306_ & new_n309_;
  assign new_n326_ = ~\count[4]  & \count[5] ;
  assign new_n327_ = new_n266_ & new_n326_;
  assign \selectp1[32]  = new_n270_ & new_n327_;
  assign \selectp1[33]  = new_n273_ & new_n327_;
  assign \selectp1[34]  = new_n276_ & new_n327_;
  assign \selectp1[35]  = new_n278_ & new_n327_;
  assign \selectp1[36]  = new_n281_ & new_n327_;
  assign \selectp1[37]  = new_n284_ & new_n327_;
  assign \selectp1[38]  = new_n286_ & new_n327_;
  assign \selectp1[39]  = new_n288_ & new_n327_;
  assign \selectp1[40]  = new_n291_ & new_n327_;
  assign \selectp1[41]  = new_n293_ & new_n327_;
  assign \selectp1[42]  = new_n296_ & new_n327_;
  assign \selectp1[43]  = new_n298_ & new_n327_;
  assign \selectp1[44]  = new_n300_ & new_n327_;
  assign \selectp1[45]  = new_n302_ & new_n327_;
  assign \selectp1[46]  = new_n304_ & new_n327_;
  assign \selectp1[47]  = new_n306_ & new_n327_;
  assign new_n344_ = \count[4]  & \count[5] ;
  assign new_n345_ = new_n266_ & new_n344_;
  assign \selectp1[48]  = new_n270_ & new_n345_;
  assign \selectp1[49]  = new_n273_ & new_n345_;
  assign \selectp1[50]  = new_n276_ & new_n345_;
  assign \selectp1[51]  = new_n278_ & new_n345_;
  assign \selectp1[52]  = new_n281_ & new_n345_;
  assign \selectp1[53]  = new_n284_ & new_n345_;
  assign \selectp1[54]  = new_n286_ & new_n345_;
  assign \selectp1[55]  = new_n288_ & new_n345_;
  assign \selectp1[56]  = new_n291_ & new_n345_;
  assign \selectp1[57]  = new_n293_ & new_n345_;
  assign \selectp1[58]  = new_n296_ & new_n345_;
  assign \selectp1[59]  = new_n298_ & new_n345_;
  assign \selectp1[60]  = new_n300_ & new_n345_;
  assign \selectp1[61]  = new_n302_ & new_n345_;
  assign \selectp1[62]  = new_n304_ & new_n345_;
  assign \selectp1[63]  = new_n306_ & new_n345_;
  assign new_n362_ = \count[6]  & \count[7] ;
  assign new_n363_ = new_n265_ & new_n362_;
  assign \selectp1[64]  = new_n270_ & new_n363_;
  assign \selectp1[65]  = new_n273_ & new_n363_;
  assign \selectp1[66]  = new_n276_ & new_n363_;
  assign \selectp1[67]  = new_n278_ & new_n363_;
  assign \selectp1[68]  = new_n281_ & new_n363_;
  assign \selectp1[69]  = new_n284_ & new_n363_;
  assign \selectp1[70]  = new_n286_ & new_n363_;
  assign \selectp1[71]  = new_n288_ & new_n363_;
  assign \selectp1[72]  = new_n291_ & new_n363_;
  assign \selectp1[73]  = new_n293_ & new_n363_;
  assign \selectp1[74]  = new_n296_ & new_n363_;
  assign \selectp1[75]  = new_n298_ & new_n363_;
  assign \selectp1[76]  = new_n300_ & new_n363_;
  assign \selectp1[77]  = new_n302_ & new_n363_;
  assign \selectp1[78]  = new_n304_ & new_n363_;
  assign \selectp1[79]  = new_n306_ & new_n363_;
  assign new_n380_ = new_n308_ & new_n362_;
  assign \selectp1[80]  = new_n270_ & new_n380_;
  assign \selectp1[81]  = new_n273_ & new_n380_;
  assign \selectp1[82]  = new_n276_ & new_n380_;
  assign \selectp1[83]  = new_n278_ & new_n380_;
  assign \selectp1[84]  = new_n281_ & new_n380_;
  assign \selectp1[85]  = new_n284_ & new_n380_;
  assign \selectp1[86]  = new_n286_ & new_n380_;
  assign \selectp1[87]  = new_n288_ & new_n380_;
  assign \selectp1[88]  = new_n291_ & new_n380_;
  assign \selectp1[89]  = new_n293_ & new_n380_;
  assign \selectp1[90]  = new_n296_ & new_n380_;
  assign \selectp1[91]  = new_n298_ & new_n380_;
  assign \selectp1[92]  = new_n300_ & new_n380_;
  assign \selectp1[93]  = new_n302_ & new_n380_;
  assign \selectp1[94]  = new_n304_ & new_n380_;
  assign \selectp1[95]  = new_n306_ & new_n380_;
  assign new_n397_ = new_n326_ & new_n362_;
  assign \selectp1[96]  = new_n270_ & new_n397_;
  assign \selectp1[97]  = new_n273_ & new_n397_;
  assign \selectp1[98]  = new_n276_ & new_n397_;
  assign \selectp1[99]  = new_n278_ & new_n397_;
  assign \selectp1[100]  = new_n281_ & new_n397_;
  assign \selectp1[101]  = new_n284_ & new_n397_;
  assign \selectp1[102]  = new_n286_ & new_n397_;
  assign \selectp1[103]  = new_n288_ & new_n397_;
  assign \selectp1[104]  = new_n291_ & new_n397_;
  assign \selectp1[105]  = new_n293_ & new_n397_;
  assign \selectp1[106]  = new_n296_ & new_n397_;
  assign \selectp1[107]  = new_n298_ & new_n397_;
  assign \selectp1[108]  = new_n300_ & new_n397_;
  assign \selectp1[109]  = new_n302_ & new_n397_;
  assign \selectp1[110]  = new_n304_ & new_n397_;
  assign \selectp1[111]  = new_n306_ & new_n397_;
  assign new_n414_ = new_n344_ & new_n362_;
  assign \selectp1[112]  = new_n270_ & new_n414_;
  assign \selectp1[113]  = new_n273_ & new_n414_;
  assign \selectp1[114]  = new_n276_ & new_n414_;
  assign \selectp1[115]  = new_n278_ & new_n414_;
  assign \selectp1[116]  = new_n281_ & new_n414_;
  assign \selectp1[117]  = new_n284_ & new_n414_;
  assign \selectp1[118]  = new_n286_ & new_n414_;
  assign \selectp1[119]  = new_n288_ & new_n414_;
  assign \selectp1[120]  = new_n291_ & new_n414_;
  assign \selectp1[121]  = new_n293_ & new_n414_;
  assign \selectp1[122]  = new_n296_ & new_n414_;
  assign \selectp1[123]  = new_n298_ & new_n414_;
  assign \selectp1[124]  = new_n300_ & new_n414_;
  assign \selectp1[125]  = new_n302_ & new_n414_;
  assign \selectp1[126]  = new_n304_ & new_n414_;
  assign \selectp1[127]  = new_n306_ & new_n414_;
  assign new_n431_ = ~\count[6]  & ~\count[7] ;
  assign new_n432_ = new_n265_ & new_n431_;
  assign \selectp2[0]  = new_n270_ & new_n432_;
  assign \selectp2[1]  = new_n273_ & new_n432_;
  assign \selectp2[2]  = new_n276_ & new_n432_;
  assign \selectp2[3]  = new_n278_ & new_n432_;
  assign \selectp2[4]  = new_n281_ & new_n432_;
  assign \selectp2[5]  = new_n284_ & new_n432_;
  assign \selectp2[6]  = new_n286_ & new_n432_;
  assign \selectp2[7]  = new_n288_ & new_n432_;
  assign \selectp2[8]  = new_n291_ & new_n432_;
  assign \selectp2[9]  = new_n293_ & new_n432_;
  assign \selectp2[10]  = new_n296_ & new_n432_;
  assign \selectp2[11]  = new_n298_ & new_n432_;
  assign \selectp2[12]  = new_n300_ & new_n432_;
  assign \selectp2[13]  = new_n302_ & new_n432_;
  assign \selectp2[14]  = new_n304_ & new_n432_;
  assign \selectp2[15]  = new_n306_ & new_n432_;
  assign new_n449_ = new_n308_ & new_n431_;
  assign \selectp2[16]  = new_n270_ & new_n449_;
  assign \selectp2[17]  = new_n273_ & new_n449_;
  assign \selectp2[18]  = new_n276_ & new_n449_;
  assign \selectp2[19]  = new_n278_ & new_n449_;
  assign \selectp2[20]  = new_n281_ & new_n449_;
  assign \selectp2[21]  = new_n284_ & new_n449_;
  assign \selectp2[22]  = new_n286_ & new_n449_;
  assign \selectp2[23]  = new_n288_ & new_n449_;
  assign \selectp2[24]  = new_n291_ & new_n449_;
  assign \selectp2[25]  = new_n293_ & new_n449_;
  assign \selectp2[26]  = new_n296_ & new_n449_;
  assign \selectp2[27]  = new_n298_ & new_n449_;
  assign \selectp2[28]  = new_n300_ & new_n449_;
  assign \selectp2[29]  = new_n302_ & new_n449_;
  assign \selectp2[30]  = new_n304_ & new_n449_;
  assign \selectp2[31]  = new_n306_ & new_n449_;
  assign new_n466_ = new_n326_ & new_n431_;
  assign \selectp2[32]  = new_n270_ & new_n466_;
  assign \selectp2[33]  = new_n273_ & new_n466_;
  assign \selectp2[34]  = new_n276_ & new_n466_;
  assign \selectp2[35]  = new_n278_ & new_n466_;
  assign \selectp2[36]  = new_n281_ & new_n466_;
  assign \selectp2[37]  = new_n284_ & new_n466_;
  assign \selectp2[38]  = new_n286_ & new_n466_;
  assign \selectp2[39]  = new_n288_ & new_n466_;
  assign \selectp2[40]  = new_n291_ & new_n466_;
  assign \selectp2[41]  = new_n293_ & new_n466_;
  assign \selectp2[42]  = new_n296_ & new_n466_;
  assign \selectp2[43]  = new_n298_ & new_n466_;
  assign \selectp2[44]  = new_n300_ & new_n466_;
  assign \selectp2[45]  = new_n302_ & new_n466_;
  assign \selectp2[46]  = new_n304_ & new_n466_;
  assign \selectp2[47]  = new_n306_ & new_n466_;
  assign new_n483_ = new_n344_ & new_n431_;
  assign \selectp2[48]  = new_n270_ & new_n483_;
  assign \selectp2[49]  = new_n273_ & new_n483_;
  assign \selectp2[50]  = new_n276_ & new_n483_;
  assign \selectp2[51]  = new_n278_ & new_n483_;
  assign \selectp2[52]  = new_n281_ & new_n483_;
  assign \selectp2[53]  = new_n284_ & new_n483_;
  assign \selectp2[54]  = new_n286_ & new_n483_;
  assign \selectp2[55]  = new_n288_ & new_n483_;
  assign \selectp2[56]  = new_n291_ & new_n483_;
  assign \selectp2[57]  = new_n293_ & new_n483_;
  assign \selectp2[58]  = new_n296_ & new_n483_;
  assign \selectp2[59]  = new_n298_ & new_n483_;
  assign \selectp2[60]  = new_n300_ & new_n483_;
  assign \selectp2[61]  = new_n302_ & new_n483_;
  assign \selectp2[62]  = new_n304_ & new_n483_;
  assign \selectp2[63]  = new_n306_ & new_n483_;
  assign new_n500_ = \count[6]  & ~\count[7] ;
  assign new_n501_ = new_n265_ & new_n500_;
  assign \selectp2[64]  = new_n270_ & new_n501_;
  assign \selectp2[65]  = new_n273_ & new_n501_;
  assign \selectp2[66]  = new_n276_ & new_n501_;
  assign \selectp2[67]  = new_n278_ & new_n501_;
  assign \selectp2[68]  = new_n281_ & new_n501_;
  assign \selectp2[69]  = new_n284_ & new_n501_;
  assign \selectp2[70]  = new_n286_ & new_n501_;
  assign \selectp2[71]  = new_n288_ & new_n501_;
  assign \selectp2[72]  = new_n291_ & new_n501_;
  assign \selectp2[73]  = new_n293_ & new_n501_;
  assign \selectp2[74]  = new_n296_ & new_n501_;
  assign \selectp2[75]  = new_n298_ & new_n501_;
  assign \selectp2[76]  = new_n300_ & new_n501_;
  assign \selectp2[77]  = new_n302_ & new_n501_;
  assign \selectp2[78]  = new_n304_ & new_n501_;
  assign \selectp2[79]  = new_n306_ & new_n501_;
  assign new_n518_ = new_n308_ & new_n500_;
  assign \selectp2[80]  = new_n270_ & new_n518_;
  assign \selectp2[81]  = new_n273_ & new_n518_;
  assign \selectp2[82]  = new_n276_ & new_n518_;
  assign \selectp2[83]  = new_n278_ & new_n518_;
  assign \selectp2[84]  = new_n281_ & new_n518_;
  assign \selectp2[85]  = new_n284_ & new_n518_;
  assign \selectp2[86]  = new_n286_ & new_n518_;
  assign \selectp2[87]  = new_n288_ & new_n518_;
  assign \selectp2[88]  = new_n291_ & new_n518_;
  assign \selectp2[89]  = new_n293_ & new_n518_;
  assign \selectp2[90]  = new_n296_ & new_n518_;
  assign \selectp2[91]  = new_n298_ & new_n518_;
  assign \selectp2[92]  = new_n300_ & new_n518_;
  assign \selectp2[93]  = new_n302_ & new_n518_;
  assign \selectp2[94]  = new_n304_ & new_n518_;
  assign \selectp2[95]  = new_n306_ & new_n518_;
  assign new_n535_ = new_n326_ & new_n500_;
  assign \selectp2[96]  = new_n270_ & new_n535_;
  assign \selectp2[97]  = new_n273_ & new_n535_;
  assign \selectp2[98]  = new_n276_ & new_n535_;
  assign \selectp2[99]  = new_n278_ & new_n535_;
  assign \selectp2[100]  = new_n281_ & new_n535_;
  assign \selectp2[101]  = new_n284_ & new_n535_;
  assign \selectp2[102]  = new_n286_ & new_n535_;
  assign \selectp2[103]  = new_n288_ & new_n535_;
  assign \selectp2[104]  = new_n291_ & new_n535_;
  assign \selectp2[105]  = new_n293_ & new_n535_;
  assign \selectp2[106]  = new_n296_ & new_n535_;
  assign \selectp2[107]  = new_n298_ & new_n535_;
  assign \selectp2[108]  = new_n300_ & new_n535_;
  assign \selectp2[109]  = new_n302_ & new_n535_;
  assign \selectp2[110]  = new_n304_ & new_n535_;
  assign \selectp2[111]  = new_n306_ & new_n535_;
  assign new_n552_ = new_n344_ & new_n500_;
  assign \selectp2[112]  = new_n270_ & new_n552_;
  assign \selectp2[113]  = new_n273_ & new_n552_;
  assign \selectp2[114]  = new_n276_ & new_n552_;
  assign \selectp2[115]  = new_n278_ & new_n552_;
  assign \selectp2[116]  = new_n281_ & new_n552_;
  assign \selectp2[117]  = new_n284_ & new_n552_;
  assign \selectp2[118]  = new_n286_ & new_n552_;
  assign \selectp2[119]  = new_n288_ & new_n552_;
  assign \selectp2[120]  = new_n291_ & new_n552_;
  assign \selectp2[121]  = new_n293_ & new_n552_;
  assign \selectp2[122]  = new_n296_ & new_n552_;
  assign \selectp2[123]  = new_n298_ & new_n552_;
  assign \selectp2[124]  = new_n300_ & new_n552_;
  assign \selectp2[125]  = new_n302_ & new_n552_;
  assign \selectp2[126]  = new_n304_ & new_n552_;
  assign \selectp2[127]  = new_n306_ & new_n552_;
endmodule


