// Benchmark "top" written by ABC on Fri Sep 15 19:21:44 2023

module top ( 
    n_1, n_2, n_3, n_4,
    n_5  );
  input  n_1, n_2, n_3, n_4;
  output n_5;
  assign n_5 = n_1 & n_4;
endmodule


