// Benchmark "i9" written by ABC on Fri Feb 25 15:13:06 2022

module i9 ( 
    \V9(3) , \V9(1) , \V9(2) , \V9(10) , \V9(0) , \V9(5) , \V9(6) ,
    \V9(7) , \V9(8) , \V56(31) , \V56(30) , \V56(29) , \V56(28) ,
    \V56(27) , \V56(26) , \V56(25) , \V56(24) , \V56(23) , \V56(22) ,
    \V56(21) , \V56(20) , \V56(19) , \V56(18) , \V56(17) , \V56(16) ,
    \V56(15) , \V56(14) , \V56(13) , \V56(12) , \V56(11) , \V56(10) ,
    \V56(9) , \V56(8) , \V56(7) , \V56(6) , \V56(5) , \V56(4) , \V56(3) ,
    \V56(2) , \V56(1) , \V56(0) , \V88(11) , \V88(10) , \V88(9) , \V88(8) ,
    \V88(7) , \V88(6) , \V88(5) , \V88(4) , \V88(3) , \V88(2) , \V88(1) ,
    \V24(14) , \V24(13) , \V24(12) , \V24(11) , \V24(10) , \V24(9) ,
    \V24(8) , \V24(7) , \V24(6) , \V24(5) , \V24(4) , \V24(3) , \V24(2) ,
    \V24(1) , \V24(0) , \V88(31) , \V88(30) , \V88(29) , \V88(28) ,
    \V88(27) , \V88(26) , \V88(25) , \V88(24) , \V88(23) , \V88(22) ,
    \V88(21) , \V88(20) , \V88(19) , \V88(18) , \V88(17) , \V88(16) ,
    \V88(15) , \V88(14) , \V88(13) , \V88(12) , \V88(0) ,
    \V119(30) , \V119(29) , \V119(28) , \V119(27) , \V119(26) , \V119(25) ,
    \V119(24) , \V119(23) , \V119(22) , \V119(21) , \V119(20) , \V119(19) ,
    \V119(18) , \V119(17) , \V119(16) , \V119(15) , \V119(14) , \V119(13) ,
    \V119(12) , \V119(11) , \V119(10) , \V119(9) , \V119(8) , \V119(7) ,
    \V119(6) , \V119(5) , \V119(4) , \V119(3) , \V119(2) , \V119(1) ,
    \V119(0) , \V151(15) , \V151(14) , \V151(13) , \V151(12) , \V151(11) ,
    \V151(10) , \V151(9) , \V151(8) , \V151(7) , \V151(6) , \V151(5) ,
    \V151(4) , \V151(3) , \V151(2) , \V151(1) , \V151(0) , \V151(31) ,
    \V151(30) , \V151(29) , \V151(28) , \V151(27) , \V151(26) , \V151(25) ,
    \V151(24) , \V151(23) , \V151(22) , \V151(21) , \V151(20) , \V151(19) ,
    \V151(18) , \V151(17) , \V151(16)   );
  input  \V9(3) , \V9(1) , \V9(2) , \V9(10) , \V9(0) , \V9(5) , \V9(6) ,
    \V9(7) , \V9(8) , \V56(31) , \V56(30) , \V56(29) , \V56(28) ,
    \V56(27) , \V56(26) , \V56(25) , \V56(24) , \V56(23) , \V56(22) ,
    \V56(21) , \V56(20) , \V56(19) , \V56(18) , \V56(17) , \V56(16) ,
    \V56(15) , \V56(14) , \V56(13) , \V56(12) , \V56(11) , \V56(10) ,
    \V56(9) , \V56(8) , \V56(7) , \V56(6) , \V56(5) , \V56(4) , \V56(3) ,
    \V56(2) , \V56(1) , \V56(0) , \V88(11) , \V88(10) , \V88(9) , \V88(8) ,
    \V88(7) , \V88(6) , \V88(5) , \V88(4) , \V88(3) , \V88(2) , \V88(1) ,
    \V24(14) , \V24(13) , \V24(12) , \V24(11) , \V24(10) , \V24(9) ,
    \V24(8) , \V24(7) , \V24(6) , \V24(5) , \V24(4) , \V24(3) , \V24(2) ,
    \V24(1) , \V24(0) , \V88(31) , \V88(30) , \V88(29) , \V88(28) ,
    \V88(27) , \V88(26) , \V88(25) , \V88(24) , \V88(23) , \V88(22) ,
    \V88(21) , \V88(20) , \V88(19) , \V88(18) , \V88(17) , \V88(16) ,
    \V88(15) , \V88(14) , \V88(13) , \V88(12) , \V88(0) ;
  output \V119(30) , \V119(29) , \V119(28) , \V119(27) , \V119(26) ,
    \V119(25) , \V119(24) , \V119(23) , \V119(22) , \V119(21) , \V119(20) ,
    \V119(19) , \V119(18) , \V119(17) , \V119(16) , \V119(15) , \V119(14) ,
    \V119(13) , \V119(12) , \V119(11) , \V119(10) , \V119(9) , \V119(8) ,
    \V119(7) , \V119(6) , \V119(5) , \V119(4) , \V119(3) , \V119(2) ,
    \V119(1) , \V119(0) , \V151(15) , \V151(14) , \V151(13) , \V151(12) ,
    \V151(11) , \V151(10) , \V151(9) , \V151(8) , \V151(7) , \V151(6) ,
    \V151(5) , \V151(4) , \V151(3) , \V151(2) , \V151(1) , \V151(0) ,
    \V151(31) , \V151(30) , \V151(29) , \V151(28) , \V151(27) , \V151(26) ,
    \V151(25) , \V151(24) , \V151(23) , \V151(22) , \V151(21) , \V151(20) ,
    \V151(19) , \V151(18) , \V151(17) , \V151(16) ;
  wire new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_;
  assign new_n152_ = ~\V9(1)  & \V9(10) ;
  assign new_n153_ = ~\V9(2)  & new_n152_;
  assign new_n154_ = ~\V9(1)  & \V9(7) ;
  assign new_n155_ = ~\V9(2)  & new_n154_;
  assign new_n156_ = ~\V9(2)  & ~\V9(6) ;
  assign new_n157_ = ~\V9(1)  & new_n156_;
  assign new_n158_ = ~\V9(5)  & new_n157_;
  assign new_n159_ = \V9(2)  & \V9(10) ;
  assign new_n160_ = \V9(1)  & \V9(10) ;
  assign new_n161_ = \V9(3)  & \V9(1) ;
  assign new_n162_ = \V9(2)  & new_n161_;
  assign new_n163_ = ~\V9(10)  & ~\V9(0) ;
  assign new_n164_ = \V9(7)  & new_n163_;
  assign new_n165_ = ~\V9(5)  & new_n163_;
  assign new_n166_ = ~\V9(10)  & ~\V9(5) ;
  assign new_n167_ = \V9(1)  & new_n166_;
  assign new_n168_ = ~\V9(2)  & new_n167_;
  assign new_n169_ = ~\V9(6)  & new_n168_;
  assign new_n170_ = \V9(1)  & ~\V9(10) ;
  assign new_n171_ = \V9(8)  & new_n170_;
  assign new_n172_ = \V9(2)  & ~\V9(10) ;
  assign new_n173_ = \V9(1)  & new_n172_;
  assign new_n174_ = ~\V9(3)  & new_n173_;
  assign new_n175_ = ~\V9(1)  & new_n166_;
  assign new_n176_ = \V9(0)  & new_n175_;
  assign new_n177_ = \V9(2)  & new_n176_;
  assign new_n178_ = ~\V9(6)  & new_n177_;
  assign new_n179_ = ~\V9(1)  & new_n172_;
  assign new_n180_ = \V9(8)  & new_n179_;
  assign new_n181_ = ~new_n174_ & ~new_n178_;
  assign new_n182_ = ~new_n180_ & new_n181_;
  assign new_n183_ = ~new_n165_ & ~new_n169_;
  assign new_n184_ = ~new_n171_ & new_n183_;
  assign new_n185_ = new_n182_ & new_n184_;
  assign new_n186_ = ~new_n160_ & ~new_n162_;
  assign new_n187_ = ~new_n164_ & new_n186_;
  assign new_n188_ = ~new_n158_ & ~new_n159_;
  assign new_n189_ = ~new_n153_ & ~new_n155_;
  assign new_n190_ = new_n188_ & new_n189_;
  assign new_n191_ = new_n187_ & new_n190_;
  assign new_n192_ = new_n185_ & new_n191_;
  assign new_n193_ = ~new_n155_ & ~new_n158_;
  assign new_n194_ = ~new_n153_ & new_n193_;
  assign new_n195_ = ~new_n164_ & ~new_n171_;
  assign new_n196_ = new_n183_ & new_n195_;
  assign new_n197_ = new_n194_ & new_n196_;
  assign new_n198_ = ~new_n178_ & ~new_n180_;
  assign new_n199_ = ~new_n174_ & new_n198_;
  assign new_n200_ = new_n194_ & new_n199_;
  assign new_n201_ = \V56(31)  & new_n197_;
  assign new_n202_ = new_n200_ & new_n201_;
  assign new_n203_ = ~new_n192_ & new_n202_;
  assign new_n204_ = ~new_n192_ & new_n200_;
  assign new_n205_ = ~new_n197_ & new_n204_;
  assign new_n206_ = \V56(23)  & new_n205_;
  assign new_n207_ = \V56(20)  & new_n197_;
  assign new_n208_ = ~new_n200_ & new_n207_;
  assign new_n209_ = ~new_n192_ & new_n208_;
  assign new_n210_ = \V56(16)  & ~new_n197_;
  assign new_n211_ = ~new_n200_ & new_n210_;
  assign new_n212_ = ~new_n192_ & new_n211_;
  assign new_n213_ = ~new_n209_ & ~new_n212_;
  assign new_n214_ = ~new_n192_ & ~new_n203_;
  assign new_n215_ = ~new_n206_ & new_n214_;
  assign \V119(30)  = ~new_n213_ | ~new_n215_;
  assign new_n217_ = \V56(30)  & new_n197_;
  assign new_n218_ = new_n200_ & new_n217_;
  assign new_n219_ = ~new_n192_ & new_n218_;
  assign new_n220_ = \V56(22)  & new_n205_;
  assign new_n221_ = \V56(19)  & new_n197_;
  assign new_n222_ = ~new_n200_ & new_n221_;
  assign new_n223_ = ~new_n192_ & new_n222_;
  assign new_n224_ = \V56(15)  & ~new_n197_;
  assign new_n225_ = ~new_n200_ & new_n224_;
  assign new_n226_ = ~new_n192_ & new_n225_;
  assign new_n227_ = ~new_n223_ & ~new_n226_;
  assign new_n228_ = ~new_n192_ & ~new_n219_;
  assign new_n229_ = ~new_n220_ & new_n228_;
  assign \V119(29)  = ~new_n227_ | ~new_n229_;
  assign new_n231_ = \V56(29)  & new_n197_;
  assign new_n232_ = new_n200_ & new_n231_;
  assign new_n233_ = ~new_n192_ & new_n232_;
  assign new_n234_ = \V56(21)  & new_n205_;
  assign new_n235_ = \V56(18)  & new_n197_;
  assign new_n236_ = ~new_n200_ & new_n235_;
  assign new_n237_ = ~new_n192_ & new_n236_;
  assign new_n238_ = \V56(14)  & ~new_n197_;
  assign new_n239_ = ~new_n200_ & new_n238_;
  assign new_n240_ = ~new_n192_ & new_n239_;
  assign new_n241_ = ~new_n237_ & ~new_n240_;
  assign new_n242_ = ~new_n192_ & ~new_n233_;
  assign new_n243_ = ~new_n234_ & new_n242_;
  assign \V119(28)  = ~new_n241_ | ~new_n243_;
  assign new_n245_ = \V56(28)  & new_n197_;
  assign new_n246_ = new_n200_ & new_n245_;
  assign new_n247_ = ~new_n192_ & new_n246_;
  assign new_n248_ = \V56(20)  & new_n205_;
  assign new_n249_ = \V56(17)  & new_n197_;
  assign new_n250_ = ~new_n200_ & new_n249_;
  assign new_n251_ = ~new_n192_ & new_n250_;
  assign new_n252_ = \V56(13)  & ~new_n197_;
  assign new_n253_ = ~new_n200_ & new_n252_;
  assign new_n254_ = ~new_n192_ & new_n253_;
  assign new_n255_ = ~new_n251_ & ~new_n254_;
  assign new_n256_ = ~new_n192_ & ~new_n247_;
  assign new_n257_ = ~new_n248_ & new_n256_;
  assign \V119(27)  = ~new_n255_ | ~new_n257_;
  assign new_n259_ = \V56(27)  & new_n197_;
  assign new_n260_ = new_n200_ & new_n259_;
  assign new_n261_ = ~new_n192_ & new_n260_;
  assign new_n262_ = \V56(19)  & new_n205_;
  assign new_n263_ = \V56(16)  & new_n197_;
  assign new_n264_ = ~new_n200_ & new_n263_;
  assign new_n265_ = ~new_n192_ & new_n264_;
  assign new_n266_ = \V56(12)  & ~new_n197_;
  assign new_n267_ = ~new_n200_ & new_n266_;
  assign new_n268_ = ~new_n192_ & new_n267_;
  assign new_n269_ = ~new_n265_ & ~new_n268_;
  assign new_n270_ = ~new_n192_ & ~new_n261_;
  assign new_n271_ = ~new_n262_ & new_n270_;
  assign \V119(26)  = ~new_n269_ | ~new_n271_;
  assign new_n273_ = \V56(26)  & new_n197_;
  assign new_n274_ = new_n200_ & new_n273_;
  assign new_n275_ = ~new_n192_ & new_n274_;
  assign new_n276_ = \V56(18)  & new_n205_;
  assign new_n277_ = \V56(15)  & new_n197_;
  assign new_n278_ = ~new_n200_ & new_n277_;
  assign new_n279_ = ~new_n192_ & new_n278_;
  assign new_n280_ = \V56(11)  & ~new_n197_;
  assign new_n281_ = ~new_n200_ & new_n280_;
  assign new_n282_ = ~new_n192_ & new_n281_;
  assign new_n283_ = ~new_n279_ & ~new_n282_;
  assign new_n284_ = ~new_n192_ & ~new_n275_;
  assign new_n285_ = ~new_n276_ & new_n284_;
  assign \V119(25)  = ~new_n283_ | ~new_n285_;
  assign new_n287_ = \V56(25)  & new_n197_;
  assign new_n288_ = new_n200_ & new_n287_;
  assign new_n289_ = ~new_n192_ & new_n288_;
  assign new_n290_ = \V56(17)  & new_n205_;
  assign new_n291_ = \V56(14)  & new_n197_;
  assign new_n292_ = ~new_n200_ & new_n291_;
  assign new_n293_ = ~new_n192_ & new_n292_;
  assign new_n294_ = \V56(10)  & ~new_n197_;
  assign new_n295_ = ~new_n200_ & new_n294_;
  assign new_n296_ = ~new_n192_ & new_n295_;
  assign new_n297_ = ~new_n293_ & ~new_n296_;
  assign new_n298_ = ~new_n192_ & ~new_n289_;
  assign new_n299_ = ~new_n290_ & new_n298_;
  assign \V119(24)  = ~new_n297_ | ~new_n299_;
  assign new_n301_ = \V56(24)  & new_n197_;
  assign new_n302_ = new_n200_ & new_n301_;
  assign new_n303_ = ~new_n192_ & new_n302_;
  assign new_n304_ = \V56(16)  & new_n205_;
  assign new_n305_ = \V56(13)  & new_n197_;
  assign new_n306_ = ~new_n200_ & new_n305_;
  assign new_n307_ = ~new_n192_ & new_n306_;
  assign new_n308_ = \V56(9)  & ~new_n197_;
  assign new_n309_ = ~new_n200_ & new_n308_;
  assign new_n310_ = ~new_n192_ & new_n309_;
  assign new_n311_ = ~new_n307_ & ~new_n310_;
  assign new_n312_ = ~new_n192_ & ~new_n303_;
  assign new_n313_ = ~new_n304_ & new_n312_;
  assign \V119(23)  = ~new_n311_ | ~new_n313_;
  assign new_n315_ = \V56(23)  & new_n197_;
  assign new_n316_ = new_n200_ & new_n315_;
  assign new_n317_ = ~new_n192_ & new_n316_;
  assign new_n318_ = \V56(15)  & new_n205_;
  assign new_n319_ = \V56(12)  & new_n197_;
  assign new_n320_ = ~new_n200_ & new_n319_;
  assign new_n321_ = ~new_n192_ & new_n320_;
  assign new_n322_ = \V56(8)  & ~new_n197_;
  assign new_n323_ = ~new_n200_ & new_n322_;
  assign new_n324_ = ~new_n192_ & new_n323_;
  assign new_n325_ = ~new_n321_ & ~new_n324_;
  assign new_n326_ = ~new_n192_ & ~new_n317_;
  assign new_n327_ = ~new_n318_ & new_n326_;
  assign \V119(22)  = ~new_n325_ | ~new_n327_;
  assign new_n329_ = \V56(22)  & new_n197_;
  assign new_n330_ = new_n200_ & new_n329_;
  assign new_n331_ = ~new_n192_ & new_n330_;
  assign new_n332_ = \V56(14)  & new_n205_;
  assign new_n333_ = \V56(11)  & new_n197_;
  assign new_n334_ = ~new_n200_ & new_n333_;
  assign new_n335_ = ~new_n192_ & new_n334_;
  assign new_n336_ = \V56(7)  & ~new_n197_;
  assign new_n337_ = ~new_n200_ & new_n336_;
  assign new_n338_ = ~new_n192_ & new_n337_;
  assign new_n339_ = ~new_n335_ & ~new_n338_;
  assign new_n340_ = ~new_n192_ & ~new_n331_;
  assign new_n341_ = ~new_n332_ & new_n340_;
  assign \V119(21)  = ~new_n339_ | ~new_n341_;
  assign new_n343_ = \V56(21)  & new_n197_;
  assign new_n344_ = new_n200_ & new_n343_;
  assign new_n345_ = ~new_n192_ & new_n344_;
  assign new_n346_ = \V56(13)  & new_n205_;
  assign new_n347_ = \V56(10)  & new_n197_;
  assign new_n348_ = ~new_n200_ & new_n347_;
  assign new_n349_ = ~new_n192_ & new_n348_;
  assign new_n350_ = \V56(6)  & ~new_n197_;
  assign new_n351_ = ~new_n200_ & new_n350_;
  assign new_n352_ = ~new_n192_ & new_n351_;
  assign new_n353_ = ~new_n349_ & ~new_n352_;
  assign new_n354_ = ~new_n192_ & ~new_n345_;
  assign new_n355_ = ~new_n346_ & new_n354_;
  assign \V119(20)  = ~new_n353_ | ~new_n355_;
  assign new_n357_ = new_n200_ & new_n207_;
  assign new_n358_ = ~new_n192_ & new_n357_;
  assign new_n359_ = \V56(12)  & new_n205_;
  assign new_n360_ = \V56(9)  & new_n197_;
  assign new_n361_ = ~new_n200_ & new_n360_;
  assign new_n362_ = ~new_n192_ & new_n361_;
  assign new_n363_ = \V56(5)  & ~new_n197_;
  assign new_n364_ = ~new_n200_ & new_n363_;
  assign new_n365_ = ~new_n192_ & new_n364_;
  assign new_n366_ = ~new_n362_ & ~new_n365_;
  assign new_n367_ = ~new_n192_ & ~new_n358_;
  assign new_n368_ = ~new_n359_ & new_n367_;
  assign \V119(19)  = ~new_n366_ | ~new_n368_;
  assign new_n370_ = new_n200_ & new_n221_;
  assign new_n371_ = ~new_n192_ & new_n370_;
  assign new_n372_ = \V56(11)  & new_n205_;
  assign new_n373_ = \V56(8)  & new_n197_;
  assign new_n374_ = ~new_n200_ & new_n373_;
  assign new_n375_ = ~new_n192_ & new_n374_;
  assign new_n376_ = \V56(4)  & ~new_n197_;
  assign new_n377_ = ~new_n200_ & new_n376_;
  assign new_n378_ = ~new_n192_ & new_n377_;
  assign new_n379_ = ~new_n375_ & ~new_n378_;
  assign new_n380_ = ~new_n192_ & ~new_n371_;
  assign new_n381_ = ~new_n372_ & new_n380_;
  assign \V119(18)  = ~new_n379_ | ~new_n381_;
  assign new_n383_ = new_n200_ & new_n235_;
  assign new_n384_ = ~new_n192_ & new_n383_;
  assign new_n385_ = \V56(10)  & new_n205_;
  assign new_n386_ = \V56(7)  & new_n197_;
  assign new_n387_ = ~new_n200_ & new_n386_;
  assign new_n388_ = ~new_n192_ & new_n387_;
  assign new_n389_ = \V56(3)  & ~new_n197_;
  assign new_n390_ = ~new_n200_ & new_n389_;
  assign new_n391_ = ~new_n192_ & new_n390_;
  assign new_n392_ = ~new_n388_ & ~new_n391_;
  assign new_n393_ = ~new_n192_ & ~new_n384_;
  assign new_n394_ = ~new_n385_ & new_n393_;
  assign \V119(17)  = ~new_n392_ | ~new_n394_;
  assign new_n396_ = new_n200_ & new_n249_;
  assign new_n397_ = ~new_n192_ & new_n396_;
  assign new_n398_ = \V56(9)  & new_n205_;
  assign new_n399_ = \V56(6)  & new_n197_;
  assign new_n400_ = ~new_n200_ & new_n399_;
  assign new_n401_ = ~new_n192_ & new_n400_;
  assign new_n402_ = \V56(2)  & ~new_n197_;
  assign new_n403_ = ~new_n200_ & new_n402_;
  assign new_n404_ = ~new_n192_ & new_n403_;
  assign new_n405_ = ~new_n401_ & ~new_n404_;
  assign new_n406_ = ~new_n192_ & ~new_n397_;
  assign new_n407_ = ~new_n398_ & new_n406_;
  assign \V119(16)  = ~new_n405_ | ~new_n407_;
  assign new_n409_ = new_n200_ & new_n263_;
  assign new_n410_ = ~new_n192_ & new_n409_;
  assign new_n411_ = \V56(8)  & new_n205_;
  assign new_n412_ = \V56(5)  & new_n197_;
  assign new_n413_ = ~new_n200_ & new_n412_;
  assign new_n414_ = ~new_n192_ & new_n413_;
  assign new_n415_ = \V56(1)  & ~new_n197_;
  assign new_n416_ = ~new_n200_ & new_n415_;
  assign new_n417_ = ~new_n192_ & new_n416_;
  assign new_n418_ = ~new_n414_ & ~new_n417_;
  assign new_n419_ = ~new_n192_ & ~new_n410_;
  assign new_n420_ = ~new_n411_ & new_n419_;
  assign \V119(15)  = ~new_n418_ | ~new_n420_;
  assign new_n422_ = new_n200_ & new_n277_;
  assign new_n423_ = ~new_n192_ & new_n422_;
  assign new_n424_ = \V56(7)  & new_n205_;
  assign new_n425_ = \V56(4)  & new_n197_;
  assign new_n426_ = ~new_n200_ & new_n425_;
  assign new_n427_ = ~new_n192_ & new_n426_;
  assign new_n428_ = \V24(14)  & ~new_n197_;
  assign new_n429_ = ~new_n200_ & new_n428_;
  assign new_n430_ = ~new_n192_ & new_n429_;
  assign new_n431_ = ~new_n427_ & ~new_n430_;
  assign new_n432_ = ~new_n192_ & ~new_n423_;
  assign new_n433_ = ~new_n424_ & new_n432_;
  assign \V119(14)  = ~new_n431_ | ~new_n433_;
  assign new_n435_ = new_n200_ & new_n291_;
  assign new_n436_ = ~new_n192_ & new_n435_;
  assign new_n437_ = \V56(6)  & new_n205_;
  assign new_n438_ = \V56(3)  & new_n197_;
  assign new_n439_ = ~new_n200_ & new_n438_;
  assign new_n440_ = ~new_n192_ & new_n439_;
  assign new_n441_ = \V24(13)  & ~new_n197_;
  assign new_n442_ = ~new_n200_ & new_n441_;
  assign new_n443_ = ~new_n192_ & new_n442_;
  assign new_n444_ = ~new_n440_ & ~new_n443_;
  assign new_n445_ = ~new_n192_ & ~new_n436_;
  assign new_n446_ = ~new_n437_ & new_n445_;
  assign \V119(13)  = ~new_n444_ | ~new_n446_;
  assign new_n448_ = new_n200_ & new_n305_;
  assign new_n449_ = ~new_n192_ & new_n448_;
  assign new_n450_ = \V56(5)  & new_n205_;
  assign new_n451_ = \V56(2)  & new_n197_;
  assign new_n452_ = ~new_n200_ & new_n451_;
  assign new_n453_ = ~new_n192_ & new_n452_;
  assign new_n454_ = \V24(12)  & ~new_n197_;
  assign new_n455_ = ~new_n200_ & new_n454_;
  assign new_n456_ = ~new_n192_ & new_n455_;
  assign new_n457_ = ~new_n453_ & ~new_n456_;
  assign new_n458_ = ~new_n192_ & ~new_n449_;
  assign new_n459_ = ~new_n450_ & new_n458_;
  assign \V119(12)  = ~new_n457_ | ~new_n459_;
  assign new_n461_ = new_n200_ & new_n319_;
  assign new_n462_ = ~new_n192_ & new_n461_;
  assign new_n463_ = \V56(4)  & new_n205_;
  assign new_n464_ = \V56(1)  & new_n197_;
  assign new_n465_ = ~new_n200_ & new_n464_;
  assign new_n466_ = ~new_n192_ & new_n465_;
  assign new_n467_ = \V24(11)  & ~new_n197_;
  assign new_n468_ = ~new_n200_ & new_n467_;
  assign new_n469_ = ~new_n192_ & new_n468_;
  assign new_n470_ = ~new_n466_ & ~new_n469_;
  assign new_n471_ = ~new_n192_ & ~new_n462_;
  assign new_n472_ = ~new_n463_ & new_n471_;
  assign \V119(11)  = ~new_n470_ | ~new_n472_;
  assign new_n474_ = new_n200_ & new_n333_;
  assign new_n475_ = ~new_n192_ & new_n474_;
  assign new_n476_ = \V56(3)  & new_n205_;
  assign new_n477_ = \V88(11)  & new_n197_;
  assign new_n478_ = ~new_n200_ & new_n477_;
  assign new_n479_ = ~new_n192_ & new_n478_;
  assign new_n480_ = \V24(10)  & ~new_n197_;
  assign new_n481_ = ~new_n200_ & new_n480_;
  assign new_n482_ = ~new_n192_ & new_n481_;
  assign new_n483_ = ~new_n479_ & ~new_n482_;
  assign new_n484_ = ~new_n192_ & ~new_n475_;
  assign new_n485_ = ~new_n476_ & new_n484_;
  assign \V119(10)  = ~new_n483_ | ~new_n485_;
  assign new_n487_ = new_n200_ & new_n347_;
  assign new_n488_ = ~new_n192_ & new_n487_;
  assign new_n489_ = \V56(2)  & new_n205_;
  assign new_n490_ = \V88(10)  & new_n197_;
  assign new_n491_ = ~new_n200_ & new_n490_;
  assign new_n492_ = ~new_n192_ & new_n491_;
  assign new_n493_ = \V24(9)  & ~new_n197_;
  assign new_n494_ = ~new_n200_ & new_n493_;
  assign new_n495_ = ~new_n192_ & new_n494_;
  assign new_n496_ = ~new_n492_ & ~new_n495_;
  assign new_n497_ = ~new_n192_ & ~new_n488_;
  assign new_n498_ = ~new_n489_ & new_n497_;
  assign \V119(9)  = ~new_n496_ | ~new_n498_;
  assign new_n500_ = new_n200_ & new_n360_;
  assign new_n501_ = ~new_n192_ & new_n500_;
  assign new_n502_ = \V56(1)  & new_n205_;
  assign new_n503_ = \V88(9)  & new_n197_;
  assign new_n504_ = ~new_n200_ & new_n503_;
  assign new_n505_ = ~new_n192_ & new_n504_;
  assign new_n506_ = \V24(8)  & ~new_n197_;
  assign new_n507_ = ~new_n200_ & new_n506_;
  assign new_n508_ = ~new_n192_ & new_n507_;
  assign new_n509_ = ~new_n505_ & ~new_n508_;
  assign new_n510_ = ~new_n192_ & ~new_n501_;
  assign new_n511_ = ~new_n502_ & new_n510_;
  assign \V119(8)  = ~new_n509_ | ~new_n511_;
  assign new_n513_ = new_n200_ & new_n373_;
  assign new_n514_ = ~new_n192_ & new_n513_;
  assign new_n515_ = \V56(0)  & new_n205_;
  assign new_n516_ = \V88(8)  & new_n197_;
  assign new_n517_ = ~new_n200_ & new_n516_;
  assign new_n518_ = ~new_n192_ & new_n517_;
  assign new_n519_ = \V24(7)  & ~new_n197_;
  assign new_n520_ = ~new_n200_ & new_n519_;
  assign new_n521_ = ~new_n192_ & new_n520_;
  assign new_n522_ = ~new_n518_ & ~new_n521_;
  assign new_n523_ = ~new_n192_ & ~new_n514_;
  assign new_n524_ = ~new_n515_ & new_n523_;
  assign \V119(7)  = ~new_n522_ | ~new_n524_;
  assign new_n526_ = new_n200_ & new_n386_;
  assign new_n527_ = ~new_n192_ & new_n526_;
  assign new_n528_ = \V88(7)  & new_n197_;
  assign new_n529_ = ~new_n200_ & new_n528_;
  assign new_n530_ = ~new_n192_ & new_n529_;
  assign new_n531_ = \V24(6)  & ~new_n197_;
  assign new_n532_ = ~new_n200_ & new_n531_;
  assign new_n533_ = ~new_n192_ & new_n532_;
  assign new_n534_ = ~new_n530_ & ~new_n533_;
  assign new_n535_ = ~new_n192_ & ~new_n527_;
  assign new_n536_ = ~new_n205_ & new_n535_;
  assign \V119(6)  = ~new_n534_ | ~new_n536_;
  assign new_n538_ = new_n200_ & new_n399_;
  assign new_n539_ = ~new_n192_ & new_n538_;
  assign new_n540_ = \V88(6)  & new_n197_;
  assign new_n541_ = ~new_n200_ & new_n540_;
  assign new_n542_ = ~new_n192_ & new_n541_;
  assign new_n543_ = \V24(5)  & ~new_n197_;
  assign new_n544_ = ~new_n200_ & new_n543_;
  assign new_n545_ = ~new_n192_ & new_n544_;
  assign new_n546_ = ~new_n542_ & ~new_n545_;
  assign new_n547_ = ~new_n192_ & ~new_n539_;
  assign new_n548_ = ~new_n205_ & new_n547_;
  assign \V119(5)  = ~new_n546_ | ~new_n548_;
  assign new_n550_ = new_n200_ & new_n412_;
  assign new_n551_ = ~new_n192_ & new_n550_;
  assign new_n552_ = \V88(5)  & new_n197_;
  assign new_n553_ = ~new_n200_ & new_n552_;
  assign new_n554_ = ~new_n192_ & new_n553_;
  assign new_n555_ = \V24(4)  & ~new_n197_;
  assign new_n556_ = ~new_n200_ & new_n555_;
  assign new_n557_ = ~new_n192_ & new_n556_;
  assign new_n558_ = ~new_n554_ & ~new_n557_;
  assign new_n559_ = ~new_n192_ & ~new_n551_;
  assign new_n560_ = ~new_n205_ & new_n559_;
  assign \V119(4)  = ~new_n558_ | ~new_n560_;
  assign new_n562_ = new_n200_ & new_n425_;
  assign new_n563_ = ~new_n192_ & new_n562_;
  assign new_n564_ = \V88(4)  & new_n197_;
  assign new_n565_ = ~new_n200_ & new_n564_;
  assign new_n566_ = ~new_n192_ & new_n565_;
  assign new_n567_ = \V24(3)  & ~new_n197_;
  assign new_n568_ = ~new_n200_ & new_n567_;
  assign new_n569_ = ~new_n192_ & new_n568_;
  assign new_n570_ = ~new_n566_ & ~new_n569_;
  assign new_n571_ = ~new_n192_ & ~new_n563_;
  assign new_n572_ = ~new_n205_ & new_n571_;
  assign \V119(3)  = ~new_n570_ | ~new_n572_;
  assign new_n574_ = new_n200_ & new_n438_;
  assign new_n575_ = ~new_n192_ & new_n574_;
  assign new_n576_ = \V88(3)  & new_n197_;
  assign new_n577_ = ~new_n200_ & new_n576_;
  assign new_n578_ = ~new_n192_ & new_n577_;
  assign new_n579_ = \V24(2)  & ~new_n197_;
  assign new_n580_ = ~new_n200_ & new_n579_;
  assign new_n581_ = ~new_n192_ & new_n580_;
  assign new_n582_ = ~new_n578_ & ~new_n581_;
  assign new_n583_ = ~new_n192_ & ~new_n575_;
  assign new_n584_ = ~new_n205_ & new_n583_;
  assign \V119(2)  = ~new_n582_ | ~new_n584_;
  assign new_n586_ = new_n200_ & new_n451_;
  assign new_n587_ = ~new_n192_ & new_n586_;
  assign new_n588_ = \V88(2)  & new_n197_;
  assign new_n589_ = ~new_n200_ & new_n588_;
  assign new_n590_ = ~new_n192_ & new_n589_;
  assign new_n591_ = \V24(1)  & ~new_n197_;
  assign new_n592_ = ~new_n200_ & new_n591_;
  assign new_n593_ = ~new_n192_ & new_n592_;
  assign new_n594_ = ~new_n590_ & ~new_n593_;
  assign new_n595_ = ~new_n192_ & ~new_n587_;
  assign new_n596_ = ~new_n205_ & new_n595_;
  assign \V119(1)  = ~new_n594_ | ~new_n596_;
  assign new_n598_ = new_n200_ & new_n464_;
  assign new_n599_ = ~new_n192_ & new_n598_;
  assign new_n600_ = \V88(1)  & new_n197_;
  assign new_n601_ = ~new_n200_ & new_n600_;
  assign new_n602_ = ~new_n192_ & new_n601_;
  assign new_n603_ = \V24(0)  & ~new_n197_;
  assign new_n604_ = ~new_n200_ & new_n603_;
  assign new_n605_ = ~new_n192_ & new_n604_;
  assign new_n606_ = ~new_n602_ & ~new_n605_;
  assign new_n607_ = ~new_n192_ & ~new_n599_;
  assign new_n608_ = ~new_n205_ & new_n607_;
  assign \V119(0)  = ~new_n606_ | ~new_n608_;
  assign new_n610_ = new_n192_ & new_n200_;
  assign new_n611_ = new_n197_ & new_n610_;
  assign new_n612_ = ~new_n197_ & new_n610_;
  assign new_n613_ = new_n192_ & ~new_n200_;
  assign new_n614_ = new_n197_ & new_n613_;
  assign new_n615_ = ~new_n197_ & new_n613_;
  assign new_n616_ = \V88(15)  & new_n197_;
  assign new_n617_ = new_n200_ & new_n616_;
  assign new_n618_ = ~new_n192_ & new_n617_;
  assign new_n619_ = \V88(7)  & ~new_n197_;
  assign new_n620_ = new_n200_ & new_n619_;
  assign new_n621_ = ~new_n192_ & new_n620_;
  assign new_n622_ = \V88(0)  & ~new_n197_;
  assign new_n623_ = ~new_n200_ & new_n622_;
  assign new_n624_ = ~new_n192_ & new_n623_;
  assign new_n625_ = ~new_n614_ & ~new_n615_;
  assign new_n626_ = ~new_n611_ & ~new_n612_;
  assign new_n627_ = new_n625_ & new_n626_;
  assign new_n628_ = ~new_n618_ & ~new_n621_;
  assign new_n629_ = ~new_n566_ & ~new_n624_;
  assign new_n630_ = new_n628_ & new_n629_;
  assign \V151(15)  = ~new_n627_ | ~new_n630_;
  assign new_n632_ = \V88(14)  & new_n197_;
  assign new_n633_ = new_n200_ & new_n632_;
  assign new_n634_ = ~new_n192_ & new_n633_;
  assign new_n635_ = \V88(6)  & ~new_n197_;
  assign new_n636_ = new_n200_ & new_n635_;
  assign new_n637_ = ~new_n192_ & new_n636_;
  assign new_n638_ = \V56(31)  & ~new_n197_;
  assign new_n639_ = ~new_n200_ & new_n638_;
  assign new_n640_ = ~new_n192_ & new_n639_;
  assign new_n641_ = ~new_n634_ & ~new_n637_;
  assign new_n642_ = ~new_n578_ & ~new_n640_;
  assign new_n643_ = new_n641_ & new_n642_;
  assign \V151(14)  = ~new_n627_ | ~new_n643_;
  assign new_n645_ = \V88(13)  & new_n197_;
  assign new_n646_ = new_n200_ & new_n645_;
  assign new_n647_ = ~new_n192_ & new_n646_;
  assign new_n648_ = \V88(5)  & ~new_n197_;
  assign new_n649_ = new_n200_ & new_n648_;
  assign new_n650_ = ~new_n192_ & new_n649_;
  assign new_n651_ = \V56(30)  & ~new_n197_;
  assign new_n652_ = ~new_n200_ & new_n651_;
  assign new_n653_ = ~new_n192_ & new_n652_;
  assign new_n654_ = ~new_n647_ & ~new_n650_;
  assign new_n655_ = ~new_n590_ & ~new_n653_;
  assign new_n656_ = new_n654_ & new_n655_;
  assign \V151(13)  = ~new_n627_ | ~new_n656_;
  assign new_n658_ = \V88(12)  & new_n197_;
  assign new_n659_ = new_n200_ & new_n658_;
  assign new_n660_ = ~new_n192_ & new_n659_;
  assign new_n661_ = \V88(4)  & ~new_n197_;
  assign new_n662_ = new_n200_ & new_n661_;
  assign new_n663_ = ~new_n192_ & new_n662_;
  assign new_n664_ = \V56(29)  & ~new_n197_;
  assign new_n665_ = ~new_n200_ & new_n664_;
  assign new_n666_ = ~new_n192_ & new_n665_;
  assign new_n667_ = ~new_n660_ & ~new_n663_;
  assign new_n668_ = ~new_n602_ & ~new_n666_;
  assign new_n669_ = new_n667_ & new_n668_;
  assign \V151(12)  = ~new_n627_ | ~new_n669_;
  assign new_n671_ = new_n200_ & new_n477_;
  assign new_n672_ = ~new_n192_ & new_n671_;
  assign new_n673_ = \V88(3)  & ~new_n197_;
  assign new_n674_ = new_n200_ & new_n673_;
  assign new_n675_ = ~new_n192_ & new_n674_;
  assign new_n676_ = \V88(0)  & new_n197_;
  assign new_n677_ = ~new_n200_ & new_n676_;
  assign new_n678_ = ~new_n192_ & new_n677_;
  assign new_n679_ = \V56(28)  & ~new_n197_;
  assign new_n680_ = ~new_n200_ & new_n679_;
  assign new_n681_ = ~new_n192_ & new_n680_;
  assign new_n682_ = ~new_n672_ & ~new_n675_;
  assign new_n683_ = ~new_n678_ & ~new_n681_;
  assign new_n684_ = new_n682_ & new_n683_;
  assign \V151(11)  = ~new_n627_ | ~new_n684_;
  assign new_n686_ = new_n200_ & new_n490_;
  assign new_n687_ = ~new_n192_ & new_n686_;
  assign new_n688_ = \V88(2)  & ~new_n197_;
  assign new_n689_ = new_n200_ & new_n688_;
  assign new_n690_ = ~new_n192_ & new_n689_;
  assign new_n691_ = ~new_n200_ & new_n201_;
  assign new_n692_ = ~new_n192_ & new_n691_;
  assign new_n693_ = \V56(27)  & ~new_n197_;
  assign new_n694_ = ~new_n200_ & new_n693_;
  assign new_n695_ = ~new_n192_ & new_n694_;
  assign new_n696_ = ~new_n687_ & ~new_n690_;
  assign new_n697_ = ~new_n692_ & ~new_n695_;
  assign new_n698_ = new_n696_ & new_n697_;
  assign \V151(10)  = ~new_n627_ | ~new_n698_;
  assign new_n700_ = new_n200_ & new_n503_;
  assign new_n701_ = ~new_n192_ & new_n700_;
  assign new_n702_ = \V88(1)  & ~new_n197_;
  assign new_n703_ = new_n200_ & new_n702_;
  assign new_n704_ = ~new_n192_ & new_n703_;
  assign new_n705_ = ~new_n200_ & new_n217_;
  assign new_n706_ = ~new_n192_ & new_n705_;
  assign new_n707_ = \V56(26)  & ~new_n197_;
  assign new_n708_ = ~new_n200_ & new_n707_;
  assign new_n709_ = ~new_n192_ & new_n708_;
  assign new_n710_ = ~new_n701_ & ~new_n704_;
  assign new_n711_ = ~new_n706_ & ~new_n709_;
  assign new_n712_ = new_n710_ & new_n711_;
  assign \V151(9)  = ~new_n627_ | ~new_n712_;
  assign new_n714_ = new_n200_ & new_n516_;
  assign new_n715_ = ~new_n192_ & new_n714_;
  assign new_n716_ = new_n200_ & new_n622_;
  assign new_n717_ = ~new_n192_ & new_n716_;
  assign new_n718_ = ~new_n200_ & new_n231_;
  assign new_n719_ = ~new_n192_ & new_n718_;
  assign new_n720_ = \V56(25)  & ~new_n197_;
  assign new_n721_ = ~new_n200_ & new_n720_;
  assign new_n722_ = ~new_n192_ & new_n721_;
  assign new_n723_ = ~new_n715_ & ~new_n717_;
  assign new_n724_ = ~new_n719_ & ~new_n722_;
  assign new_n725_ = new_n723_ & new_n724_;
  assign \V151(8)  = ~new_n627_ | ~new_n725_;
  assign new_n727_ = new_n200_ & new_n528_;
  assign new_n728_ = ~new_n192_ & new_n727_;
  assign new_n729_ = new_n200_ & new_n638_;
  assign new_n730_ = ~new_n192_ & new_n729_;
  assign new_n731_ = ~new_n200_ & new_n245_;
  assign new_n732_ = ~new_n192_ & new_n731_;
  assign new_n733_ = \V56(24)  & ~new_n197_;
  assign new_n734_ = ~new_n200_ & new_n733_;
  assign new_n735_ = ~new_n192_ & new_n734_;
  assign new_n736_ = ~new_n728_ & ~new_n730_;
  assign new_n737_ = ~new_n732_ & ~new_n735_;
  assign new_n738_ = new_n736_ & new_n737_;
  assign \V151(7)  = ~new_n627_ | ~new_n738_;
  assign new_n740_ = new_n200_ & new_n540_;
  assign new_n741_ = ~new_n192_ & new_n740_;
  assign new_n742_ = new_n200_ & new_n651_;
  assign new_n743_ = ~new_n192_ & new_n742_;
  assign new_n744_ = ~new_n200_ & new_n259_;
  assign new_n745_ = ~new_n192_ & new_n744_;
  assign new_n746_ = \V56(23)  & ~new_n197_;
  assign new_n747_ = ~new_n200_ & new_n746_;
  assign new_n748_ = ~new_n192_ & new_n747_;
  assign new_n749_ = ~new_n741_ & ~new_n743_;
  assign new_n750_ = ~new_n745_ & ~new_n748_;
  assign new_n751_ = new_n749_ & new_n750_;
  assign \V151(6)  = ~new_n627_ | ~new_n751_;
  assign new_n753_ = new_n200_ & new_n552_;
  assign new_n754_ = ~new_n192_ & new_n753_;
  assign new_n755_ = new_n200_ & new_n664_;
  assign new_n756_ = ~new_n192_ & new_n755_;
  assign new_n757_ = ~new_n200_ & new_n273_;
  assign new_n758_ = ~new_n192_ & new_n757_;
  assign new_n759_ = \V56(22)  & ~new_n197_;
  assign new_n760_ = ~new_n200_ & new_n759_;
  assign new_n761_ = ~new_n192_ & new_n760_;
  assign new_n762_ = ~new_n754_ & ~new_n756_;
  assign new_n763_ = ~new_n758_ & ~new_n761_;
  assign new_n764_ = new_n762_ & new_n763_;
  assign \V151(5)  = ~new_n627_ | ~new_n764_;
  assign new_n766_ = new_n200_ & new_n564_;
  assign new_n767_ = ~new_n192_ & new_n766_;
  assign new_n768_ = new_n200_ & new_n679_;
  assign new_n769_ = ~new_n192_ & new_n768_;
  assign new_n770_ = ~new_n200_ & new_n287_;
  assign new_n771_ = ~new_n192_ & new_n770_;
  assign new_n772_ = \V56(21)  & ~new_n197_;
  assign new_n773_ = ~new_n200_ & new_n772_;
  assign new_n774_ = ~new_n192_ & new_n773_;
  assign new_n775_ = ~new_n767_ & ~new_n769_;
  assign new_n776_ = ~new_n771_ & ~new_n774_;
  assign new_n777_ = new_n775_ & new_n776_;
  assign \V151(4)  = ~new_n627_ | ~new_n777_;
  assign new_n779_ = new_n200_ & new_n576_;
  assign new_n780_ = ~new_n192_ & new_n779_;
  assign new_n781_ = new_n200_ & new_n693_;
  assign new_n782_ = ~new_n192_ & new_n781_;
  assign new_n783_ = ~new_n200_ & new_n301_;
  assign new_n784_ = ~new_n192_ & new_n783_;
  assign new_n785_ = \V56(20)  & ~new_n197_;
  assign new_n786_ = ~new_n200_ & new_n785_;
  assign new_n787_ = ~new_n192_ & new_n786_;
  assign new_n788_ = ~new_n780_ & ~new_n782_;
  assign new_n789_ = ~new_n784_ & ~new_n787_;
  assign new_n790_ = new_n788_ & new_n789_;
  assign \V151(3)  = ~new_n627_ | ~new_n790_;
  assign new_n792_ = new_n200_ & new_n588_;
  assign new_n793_ = ~new_n192_ & new_n792_;
  assign new_n794_ = new_n200_ & new_n707_;
  assign new_n795_ = ~new_n192_ & new_n794_;
  assign new_n796_ = ~new_n200_ & new_n315_;
  assign new_n797_ = ~new_n192_ & new_n796_;
  assign new_n798_ = \V56(19)  & ~new_n197_;
  assign new_n799_ = ~new_n200_ & new_n798_;
  assign new_n800_ = ~new_n192_ & new_n799_;
  assign new_n801_ = ~new_n793_ & ~new_n795_;
  assign new_n802_ = ~new_n797_ & ~new_n800_;
  assign new_n803_ = new_n801_ & new_n802_;
  assign \V151(2)  = ~new_n627_ | ~new_n803_;
  assign new_n805_ = new_n200_ & new_n600_;
  assign new_n806_ = ~new_n192_ & new_n805_;
  assign new_n807_ = new_n200_ & new_n720_;
  assign new_n808_ = ~new_n192_ & new_n807_;
  assign new_n809_ = ~new_n200_ & new_n329_;
  assign new_n810_ = ~new_n192_ & new_n809_;
  assign new_n811_ = \V56(18)  & ~new_n197_;
  assign new_n812_ = ~new_n200_ & new_n811_;
  assign new_n813_ = ~new_n192_ & new_n812_;
  assign new_n814_ = ~new_n806_ & ~new_n808_;
  assign new_n815_ = ~new_n810_ & ~new_n813_;
  assign new_n816_ = new_n814_ & new_n815_;
  assign \V151(1)  = ~new_n627_ | ~new_n816_;
  assign new_n818_ = new_n200_ & new_n676_;
  assign new_n819_ = ~new_n192_ & new_n818_;
  assign new_n820_ = new_n200_ & new_n733_;
  assign new_n821_ = ~new_n192_ & new_n820_;
  assign new_n822_ = ~new_n200_ & new_n343_;
  assign new_n823_ = ~new_n192_ & new_n822_;
  assign new_n824_ = \V56(17)  & ~new_n197_;
  assign new_n825_ = ~new_n200_ & new_n824_;
  assign new_n826_ = ~new_n192_ & new_n825_;
  assign new_n827_ = ~new_n819_ & ~new_n821_;
  assign new_n828_ = ~new_n823_ & ~new_n826_;
  assign new_n829_ = new_n827_ & new_n828_;
  assign \V151(0)  = ~new_n627_ | ~new_n829_;
  assign new_n831_ = \V88(31)  & new_n197_;
  assign new_n832_ = new_n200_ & new_n831_;
  assign new_n833_ = ~new_n192_ & new_n832_;
  assign new_n834_ = \V88(23)  & ~new_n197_;
  assign new_n835_ = new_n200_ & new_n834_;
  assign new_n836_ = ~new_n192_ & new_n835_;
  assign new_n837_ = \V88(20)  & new_n197_;
  assign new_n838_ = ~new_n200_ & new_n837_;
  assign new_n839_ = ~new_n192_ & new_n838_;
  assign new_n840_ = \V88(16)  & ~new_n197_;
  assign new_n841_ = ~new_n200_ & new_n840_;
  assign new_n842_ = ~new_n192_ & new_n841_;
  assign new_n843_ = ~new_n833_ & ~new_n836_;
  assign new_n844_ = ~new_n839_ & ~new_n842_;
  assign new_n845_ = new_n843_ & new_n844_;
  assign \V151(31)  = ~new_n627_ | ~new_n845_;
  assign new_n847_ = \V88(30)  & new_n197_;
  assign new_n848_ = new_n200_ & new_n847_;
  assign new_n849_ = ~new_n192_ & new_n848_;
  assign new_n850_ = \V88(22)  & ~new_n197_;
  assign new_n851_ = new_n200_ & new_n850_;
  assign new_n852_ = ~new_n192_ & new_n851_;
  assign new_n853_ = \V88(19)  & new_n197_;
  assign new_n854_ = ~new_n200_ & new_n853_;
  assign new_n855_ = ~new_n192_ & new_n854_;
  assign new_n856_ = \V88(15)  & ~new_n197_;
  assign new_n857_ = ~new_n200_ & new_n856_;
  assign new_n858_ = ~new_n192_ & new_n857_;
  assign new_n859_ = ~new_n849_ & ~new_n852_;
  assign new_n860_ = ~new_n855_ & ~new_n858_;
  assign new_n861_ = new_n859_ & new_n860_;
  assign \V151(30)  = ~new_n627_ | ~new_n861_;
  assign new_n863_ = \V88(29)  & new_n197_;
  assign new_n864_ = new_n200_ & new_n863_;
  assign new_n865_ = ~new_n192_ & new_n864_;
  assign new_n866_ = \V88(21)  & ~new_n197_;
  assign new_n867_ = new_n200_ & new_n866_;
  assign new_n868_ = ~new_n192_ & new_n867_;
  assign new_n869_ = \V88(18)  & new_n197_;
  assign new_n870_ = ~new_n200_ & new_n869_;
  assign new_n871_ = ~new_n192_ & new_n870_;
  assign new_n872_ = \V88(14)  & ~new_n197_;
  assign new_n873_ = ~new_n200_ & new_n872_;
  assign new_n874_ = ~new_n192_ & new_n873_;
  assign new_n875_ = ~new_n865_ & ~new_n868_;
  assign new_n876_ = ~new_n871_ & ~new_n874_;
  assign new_n877_ = new_n875_ & new_n876_;
  assign \V151(29)  = ~new_n627_ | ~new_n877_;
  assign new_n879_ = \V88(28)  & new_n197_;
  assign new_n880_ = new_n200_ & new_n879_;
  assign new_n881_ = ~new_n192_ & new_n880_;
  assign new_n882_ = \V88(20)  & ~new_n197_;
  assign new_n883_ = new_n200_ & new_n882_;
  assign new_n884_ = ~new_n192_ & new_n883_;
  assign new_n885_ = \V88(17)  & new_n197_;
  assign new_n886_ = ~new_n200_ & new_n885_;
  assign new_n887_ = ~new_n192_ & new_n886_;
  assign new_n888_ = \V88(13)  & ~new_n197_;
  assign new_n889_ = ~new_n200_ & new_n888_;
  assign new_n890_ = ~new_n192_ & new_n889_;
  assign new_n891_ = ~new_n881_ & ~new_n884_;
  assign new_n892_ = ~new_n887_ & ~new_n890_;
  assign new_n893_ = new_n891_ & new_n892_;
  assign \V151(28)  = ~new_n627_ | ~new_n893_;
  assign new_n895_ = \V88(27)  & new_n197_;
  assign new_n896_ = new_n200_ & new_n895_;
  assign new_n897_ = ~new_n192_ & new_n896_;
  assign new_n898_ = \V88(19)  & ~new_n197_;
  assign new_n899_ = new_n200_ & new_n898_;
  assign new_n900_ = ~new_n192_ & new_n899_;
  assign new_n901_ = \V88(16)  & new_n197_;
  assign new_n902_ = ~new_n200_ & new_n901_;
  assign new_n903_ = ~new_n192_ & new_n902_;
  assign new_n904_ = \V88(12)  & ~new_n197_;
  assign new_n905_ = ~new_n200_ & new_n904_;
  assign new_n906_ = ~new_n192_ & new_n905_;
  assign new_n907_ = ~new_n897_ & ~new_n900_;
  assign new_n908_ = ~new_n903_ & ~new_n906_;
  assign new_n909_ = new_n907_ & new_n908_;
  assign \V151(27)  = ~new_n627_ | ~new_n909_;
  assign new_n911_ = \V88(26)  & new_n197_;
  assign new_n912_ = new_n200_ & new_n911_;
  assign new_n913_ = ~new_n192_ & new_n912_;
  assign new_n914_ = \V88(18)  & ~new_n197_;
  assign new_n915_ = new_n200_ & new_n914_;
  assign new_n916_ = ~new_n192_ & new_n915_;
  assign new_n917_ = ~new_n200_ & new_n616_;
  assign new_n918_ = ~new_n192_ & new_n917_;
  assign new_n919_ = \V88(11)  & ~new_n197_;
  assign new_n920_ = ~new_n200_ & new_n919_;
  assign new_n921_ = ~new_n192_ & new_n920_;
  assign new_n922_ = ~new_n913_ & ~new_n916_;
  assign new_n923_ = ~new_n918_ & ~new_n921_;
  assign new_n924_ = new_n922_ & new_n923_;
  assign \V151(26)  = ~new_n627_ | ~new_n924_;
  assign new_n926_ = \V88(25)  & new_n197_;
  assign new_n927_ = new_n200_ & new_n926_;
  assign new_n928_ = ~new_n192_ & new_n927_;
  assign new_n929_ = \V88(17)  & ~new_n197_;
  assign new_n930_ = new_n200_ & new_n929_;
  assign new_n931_ = ~new_n192_ & new_n930_;
  assign new_n932_ = ~new_n200_ & new_n632_;
  assign new_n933_ = ~new_n192_ & new_n932_;
  assign new_n934_ = \V88(10)  & ~new_n197_;
  assign new_n935_ = ~new_n200_ & new_n934_;
  assign new_n936_ = ~new_n192_ & new_n935_;
  assign new_n937_ = ~new_n928_ & ~new_n931_;
  assign new_n938_ = ~new_n933_ & ~new_n936_;
  assign new_n939_ = new_n937_ & new_n938_;
  assign \V151(25)  = ~new_n627_ | ~new_n939_;
  assign new_n941_ = \V88(24)  & new_n197_;
  assign new_n942_ = new_n200_ & new_n941_;
  assign new_n943_ = ~new_n192_ & new_n942_;
  assign new_n944_ = new_n200_ & new_n840_;
  assign new_n945_ = ~new_n192_ & new_n944_;
  assign new_n946_ = ~new_n200_ & new_n645_;
  assign new_n947_ = ~new_n192_ & new_n946_;
  assign new_n948_ = \V88(9)  & ~new_n197_;
  assign new_n949_ = ~new_n200_ & new_n948_;
  assign new_n950_ = ~new_n192_ & new_n949_;
  assign new_n951_ = ~new_n943_ & ~new_n945_;
  assign new_n952_ = ~new_n947_ & ~new_n950_;
  assign new_n953_ = new_n951_ & new_n952_;
  assign \V151(24)  = ~new_n627_ | ~new_n953_;
  assign new_n955_ = \V88(23)  & new_n197_;
  assign new_n956_ = new_n200_ & new_n955_;
  assign new_n957_ = ~new_n192_ & new_n956_;
  assign new_n958_ = new_n200_ & new_n856_;
  assign new_n959_ = ~new_n192_ & new_n958_;
  assign new_n960_ = ~new_n200_ & new_n658_;
  assign new_n961_ = ~new_n192_ & new_n960_;
  assign new_n962_ = \V88(8)  & ~new_n197_;
  assign new_n963_ = ~new_n200_ & new_n962_;
  assign new_n964_ = ~new_n192_ & new_n963_;
  assign new_n965_ = ~new_n957_ & ~new_n959_;
  assign new_n966_ = ~new_n961_ & ~new_n964_;
  assign new_n967_ = new_n965_ & new_n966_;
  assign \V151(23)  = ~new_n627_ | ~new_n967_;
  assign new_n969_ = \V88(22)  & new_n197_;
  assign new_n970_ = new_n200_ & new_n969_;
  assign new_n971_ = ~new_n192_ & new_n970_;
  assign new_n972_ = new_n200_ & new_n872_;
  assign new_n973_ = ~new_n192_ & new_n972_;
  assign new_n974_ = ~new_n200_ & new_n619_;
  assign new_n975_ = ~new_n192_ & new_n974_;
  assign new_n976_ = ~new_n971_ & ~new_n973_;
  assign new_n977_ = ~new_n479_ & ~new_n975_;
  assign new_n978_ = new_n976_ & new_n977_;
  assign \V151(22)  = ~new_n627_ | ~new_n978_;
  assign new_n980_ = \V88(21)  & new_n197_;
  assign new_n981_ = new_n200_ & new_n980_;
  assign new_n982_ = ~new_n192_ & new_n981_;
  assign new_n983_ = new_n200_ & new_n888_;
  assign new_n984_ = ~new_n192_ & new_n983_;
  assign new_n985_ = ~new_n200_ & new_n635_;
  assign new_n986_ = ~new_n192_ & new_n985_;
  assign new_n987_ = ~new_n982_ & ~new_n984_;
  assign new_n988_ = ~new_n492_ & ~new_n986_;
  assign new_n989_ = new_n987_ & new_n988_;
  assign \V151(21)  = ~new_n627_ | ~new_n989_;
  assign new_n991_ = new_n200_ & new_n837_;
  assign new_n992_ = ~new_n192_ & new_n991_;
  assign new_n993_ = new_n200_ & new_n904_;
  assign new_n994_ = ~new_n192_ & new_n993_;
  assign new_n995_ = ~new_n200_ & new_n648_;
  assign new_n996_ = ~new_n192_ & new_n995_;
  assign new_n997_ = ~new_n992_ & ~new_n994_;
  assign new_n998_ = ~new_n505_ & ~new_n996_;
  assign new_n999_ = new_n997_ & new_n998_;
  assign \V151(20)  = ~new_n627_ | ~new_n999_;
  assign new_n1001_ = new_n200_ & new_n853_;
  assign new_n1002_ = ~new_n192_ & new_n1001_;
  assign new_n1003_ = new_n200_ & new_n919_;
  assign new_n1004_ = ~new_n192_ & new_n1003_;
  assign new_n1005_ = ~new_n200_ & new_n661_;
  assign new_n1006_ = ~new_n192_ & new_n1005_;
  assign new_n1007_ = ~new_n1002_ & ~new_n1004_;
  assign new_n1008_ = ~new_n518_ & ~new_n1006_;
  assign new_n1009_ = new_n1007_ & new_n1008_;
  assign \V151(19)  = ~new_n627_ | ~new_n1009_;
  assign new_n1011_ = new_n200_ & new_n869_;
  assign new_n1012_ = ~new_n192_ & new_n1011_;
  assign new_n1013_ = new_n200_ & new_n934_;
  assign new_n1014_ = ~new_n192_ & new_n1013_;
  assign new_n1015_ = ~new_n200_ & new_n673_;
  assign new_n1016_ = ~new_n192_ & new_n1015_;
  assign new_n1017_ = ~new_n1012_ & ~new_n1014_;
  assign new_n1018_ = ~new_n530_ & ~new_n1016_;
  assign new_n1019_ = new_n1017_ & new_n1018_;
  assign \V151(18)  = ~new_n627_ | ~new_n1019_;
  assign new_n1021_ = new_n200_ & new_n885_;
  assign new_n1022_ = ~new_n192_ & new_n1021_;
  assign new_n1023_ = new_n200_ & new_n948_;
  assign new_n1024_ = ~new_n192_ & new_n1023_;
  assign new_n1025_ = ~new_n200_ & new_n688_;
  assign new_n1026_ = ~new_n192_ & new_n1025_;
  assign new_n1027_ = ~new_n1022_ & ~new_n1024_;
  assign new_n1028_ = ~new_n542_ & ~new_n1026_;
  assign new_n1029_ = new_n1027_ & new_n1028_;
  assign \V151(17)  = ~new_n627_ | ~new_n1029_;
  assign new_n1031_ = new_n200_ & new_n901_;
  assign new_n1032_ = ~new_n192_ & new_n1031_;
  assign new_n1033_ = new_n200_ & new_n962_;
  assign new_n1034_ = ~new_n192_ & new_n1033_;
  assign new_n1035_ = ~new_n200_ & new_n702_;
  assign new_n1036_ = ~new_n192_ & new_n1035_;
  assign new_n1037_ = ~new_n1032_ & ~new_n1034_;
  assign new_n1038_ = ~new_n554_ & ~new_n1036_;
  assign new_n1039_ = new_n1037_ & new_n1038_;
  assign \V151(16)  = ~new_n627_ | ~new_n1039_;
endmodule


