// Benchmark "square" written by ABC on Thu Sep 14 23:16:29 2023

module square ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ;
  output \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127] ;
  wire new_n194_, new_n196_, new_n197_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n527_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n599_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1764_, new_n1765_,
    new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_,
    new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_,
    new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1948_,
    new_n1949_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_,
    new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_,
    new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_,
    new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_,
    new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_,
    new_n2582_, new_n2583_, new_n2584_, new_n2586_, new_n2587_, new_n2588_,
    new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_,
    new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_,
    new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_,
    new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_,
    new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_,
    new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_,
    new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_,
    new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_,
    new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_,
    new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_,
    new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_,
    new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_,
    new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_,
    new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_,
    new_n2679_, new_n2680_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_,
    new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_,
    new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_,
    new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_,
    new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3020_, new_n3021_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_,
    new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_,
    new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_,
    new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_,
    new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_,
    new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_,
    new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_,
    new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_,
    new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_,
    new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_,
    new_n3173_, new_n3174_, new_n3175_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3382_,
    new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_,
    new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_,
    new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_,
    new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_,
    new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_,
    new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_,
    new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_,
    new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_,
    new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_,
    new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_,
    new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_,
    new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_,
    new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_,
    new_n3461_, new_n3462_, new_n3463_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_,
    new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_,
    new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_,
    new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_,
    new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_,
    new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_,
    new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_,
    new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_,
    new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_,
    new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_,
    new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_,
    new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_,
    new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_,
    new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_,
    new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_,
    new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_,
    new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_,
    new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3728_, new_n3729_,
    new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_,
    new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_,
    new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_,
    new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_,
    new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_,
    new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_,
    new_n3767_, new_n3768_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_,
    new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_,
    new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_,
    new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_,
    new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_,
    new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_,
    new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_,
    new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_,
    new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_,
    new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_,
    new_n3943_, new_n3944_, new_n3945_, new_n3947_, new_n3948_, new_n3949_,
    new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_,
    new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_,
    new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_,
    new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_,
    new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_,
    new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_,
    new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_,
    new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_,
    new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_,
    new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_,
    new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_,
    new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_,
    new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_,
    new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_,
    new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_,
    new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_,
    new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_,
    new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_,
    new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_,
    new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_,
    new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_,
    new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_,
    new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_,
    new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_,
    new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_,
    new_n4112_, new_n4113_, new_n4115_, new_n4116_, new_n4117_, new_n4118_,
    new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_,
    new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_,
    new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_,
    new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_,
    new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_,
    new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_,
    new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_,
    new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_,
    new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_,
    new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_,
    new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_,
    new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_,
    new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_,
    new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_,
    new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_,
    new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_,
    new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_,
    new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_,
    new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_,
    new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_,
    new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_,
    new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_,
    new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_,
    new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_,
    new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_,
    new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_,
    new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_,
    new_n4683_, new_n4684_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_,
    new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_,
    new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_,
    new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_,
    new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_,
    new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_,
    new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_,
    new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_,
    new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_,
    new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_,
    new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_,
    new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_,
    new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_,
    new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_,
    new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_,
    new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_,
    new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4857_, new_n4858_,
    new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_,
    new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_,
    new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_,
    new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_,
    new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_,
    new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_,
    new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_,
    new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_,
    new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_,
    new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_,
    new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_,
    new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_,
    new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_,
    new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_,
    new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_,
    new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_,
    new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_,
    new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_,
    new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_,
    new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_,
    new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_,
    new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_,
    new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_,
    new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_,
    new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_,
    new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5229_, new_n5230_, new_n5231_, new_n5232_,
    new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_,
    new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_,
    new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_,
    new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_,
    new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_,
    new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_,
    new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_,
    new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_,
    new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_,
    new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_,
    new_n5293_, new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_,
    new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_,
    new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_,
    new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_,
    new_n5320_, new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_,
    new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_,
    new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_,
    new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_,
    new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_,
    new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_,
    new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_,
    new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_,
    new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_,
    new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_,
    new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_,
    new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_,
    new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_,
    new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_,
    new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_,
    new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_,
    new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_,
    new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_,
    new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_,
    new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_,
    new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_,
    new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_,
    new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_,
    new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_,
    new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_,
    new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_,
    new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_,
    new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_,
    new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_,
    new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_,
    new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_,
    new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_,
    new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_,
    new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_,
    new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_,
    new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_,
    new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_,
    new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_,
    new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_,
    new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_,
    new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_,
    new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_,
    new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_,
    new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_,
    new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_,
    new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_,
    new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_,
    new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_,
    new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_,
    new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_,
    new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_,
    new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_,
    new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_,
    new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_,
    new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_,
    new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_,
    new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_,
    new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_,
    new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_,
    new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_,
    new_n5785_, new_n5786_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_,
    new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_,
    new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5833_, new_n5834_,
    new_n5835_, new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_,
    new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_,
    new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_,
    new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_,
    new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_,
    new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_,
    new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_,
    new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_,
    new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_,
    new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_,
    new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_,
    new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_,
    new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_,
    new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_,
    new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_,
    new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_,
    new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_,
    new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_, new_n5943_,
    new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_, new_n5949_,
    new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5955_,
    new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5961_,
    new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_, new_n5967_,
    new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_, new_n5973_,
    new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_,
    new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_,
    new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_,
    new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_,
    new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_,
    new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_,
    new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_,
    new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_,
    new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_,
    new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_,
    new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_,
    new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_,
    new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_,
    new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_,
    new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_,
    new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_,
    new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_,
    new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_,
    new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_,
    new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_,
    new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_,
    new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_,
    new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_,
    new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_,
    new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_,
    new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_,
    new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_,
    new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_,
    new_n6244_, new_n6245_, new_n6247_, new_n6248_, new_n6249_, new_n6250_,
    new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_,
    new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_,
    new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_,
    new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_,
    new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_,
    new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_,
    new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_,
    new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_,
    new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_,
    new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_,
    new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_,
    new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_,
    new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_,
    new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_,
    new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_,
    new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_,
    new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_,
    new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_,
    new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_,
    new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_,
    new_n6407_, new_n6411_, new_n6412_, new_n6413_, new_n6419_, new_n6420_,
    new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_,
    new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_,
    new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_,
    new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_,
    new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_,
    new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_,
    new_n6457_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_,
    new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_,
    new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_,
    new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_,
    new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_,
    new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_,
    new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_,
    new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_,
    new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6674_, new_n6675_,
    new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_,
    new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6690_,
    new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_,
    new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_,
    new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_,
    new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_,
    new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_,
    new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_,
    new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_,
    new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_,
    new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_,
    new_n6745_, new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_,
    new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_, new_n6759_,
    new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_, new_n6765_,
    new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_, new_n6771_,
    new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_, new_n6777_,
    new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_, new_n6783_,
    new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_,
    new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_, new_n6795_,
    new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n6801_,
    new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_, new_n6807_,
    new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_,
    new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_, new_n6819_,
    new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_, new_n6825_,
    new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_, new_n6831_,
    new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_, new_n6837_,
    new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_, new_n6843_,
    new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6849_,
    new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_, new_n6855_,
    new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_, new_n6861_,
    new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_, new_n6867_,
    new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_, new_n6873_,
    new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_, new_n6879_,
    new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_, new_n6885_,
    new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_, new_n6891_,
    new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_, new_n6897_,
    new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_, new_n6903_,
    new_n6904_, new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_,
    new_n6911_, new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_,
    new_n6917_, new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_,
    new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_,
    new_n6929_, new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_,
    new_n6935_, new_n6936_, new_n6937_, new_n6938_, new_n6939_, new_n6940_,
    new_n6941_, new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_,
    new_n6947_, new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_,
    new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_,
    new_n6959_, new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_,
    new_n6965_, new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_,
    new_n6971_, new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_,
    new_n6977_, new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_,
    new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_,
    new_n6989_, new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_,
    new_n6995_, new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_,
    new_n7001_, new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_,
    new_n7007_, new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_,
    new_n7013_, new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_,
    new_n7019_, new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_,
    new_n7025_, new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_,
    new_n7031_, new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_,
    new_n7037_, new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_,
    new_n7043_, new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_,
    new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_,
    new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_,
    new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_,
    new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_,
    new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_,
    new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_,
    new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_,
    new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_,
    new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_,
    new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_,
    new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_,
    new_n7115_, new_n7116_, new_n7117_, new_n7119_, new_n7120_, new_n7121_,
    new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_,
    new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_,
    new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_,
    new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_,
    new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_,
    new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_,
    new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_,
    new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_,
    new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_,
    new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_,
    new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_,
    new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_,
    new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_,
    new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_,
    new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_,
    new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_,
    new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_,
    new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_,
    new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_,
    new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_,
    new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_,
    new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_,
    new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_,
    new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_,
    new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_,
    new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_,
    new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_,
    new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_,
    new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_,
    new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_,
    new_n7350_, new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_,
    new_n7356_, new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_,
    new_n7362_, new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_,
    new_n7368_, new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_,
    new_n7374_, new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_,
    new_n7380_, new_n7381_, new_n7382_, new_n7384_, new_n7385_, new_n7386_,
    new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_,
    new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_,
    new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_,
    new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_,
    new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_,
    new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_,
    new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_,
    new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_,
    new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_,
    new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_,
    new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_,
    new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_,
    new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_,
    new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_,
    new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_,
    new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_,
    new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_,
    new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_,
    new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_,
    new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_,
    new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_,
    new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_,
    new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_,
    new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_,
    new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_,
    new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_,
    new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7646_,
    new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_,
    new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_,
    new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_,
    new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_,
    new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_,
    new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_,
    new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_,
    new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_,
    new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_,
    new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_,
    new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_,
    new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_,
    new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_,
    new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_,
    new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_,
    new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_,
    new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_,
    new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_,
    new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_,
    new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_,
    new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_,
    new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_,
    new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_,
    new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_,
    new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_,
    new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_,
    new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_,
    new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_,
    new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_,
    new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_,
    new_n7881_, new_n7882_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_,
    new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_,
    new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_,
    new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_,
    new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_,
    new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_,
    new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_,
    new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_,
    new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_,
    new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_,
    new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_,
    new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_,
    new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_,
    new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_,
    new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_,
    new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_,
    new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_,
    new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_,
    new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_,
    new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8031_, new_n8032_,
    new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_,
    new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_,
    new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_,
    new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_,
    new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_,
    new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_,
    new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_,
    new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_,
    new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_,
    new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_,
    new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_,
    new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_,
    new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_,
    new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_,
    new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8177_, new_n8178_,
    new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_,
    new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_,
    new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_,
    new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_,
    new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_,
    new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_,
    new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_,
    new_n8221_, new_n8222_, new_n8226_, new_n8227_, new_n8228_, new_n8229_,
    new_n8230_, new_n8231_, new_n8233_, new_n8234_, new_n8235_, new_n8236_,
    new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_,
    new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_,
    new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_,
    new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_,
    new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_,
    new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_,
    new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_,
    new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_,
    new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_,
    new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_,
    new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_,
    new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_,
    new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_,
    new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_,
    new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_,
    new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_,
    new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_,
    new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_,
    new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_,
    new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_,
    new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_,
    new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_,
    new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8452_, new_n8453_, new_n8454_, new_n8455_, new_n8456_,
    new_n8457_, new_n8458_, new_n8459_, new_n8460_, new_n8461_, new_n8462_,
    new_n8463_, new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_,
    new_n8469_, new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_,
    new_n8475_, new_n8476_, new_n8477_, new_n8478_, new_n8479_, new_n8480_,
    new_n8481_, new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_,
    new_n8487_, new_n8488_, new_n8489_, new_n8490_, new_n8491_, new_n8492_,
    new_n8493_, new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8498_,
    new_n8499_, new_n8500_, new_n8501_, new_n8502_, new_n8503_, new_n8504_,
    new_n8505_, new_n8506_, new_n8507_, new_n8508_, new_n8509_, new_n8510_,
    new_n8511_, new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_,
    new_n8517_, new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_,
    new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_,
    new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_,
    new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_,
    new_n8541_, new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_,
    new_n8547_, new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_,
    new_n8553_, new_n8554_, new_n8555_, new_n8556_, new_n8557_, new_n8558_,
    new_n8559_, new_n8560_, new_n8561_, new_n8562_, new_n8563_, new_n8564_,
    new_n8565_, new_n8566_, new_n8570_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_,
    new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_,
    new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_,
    new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_,
    new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_,
    new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_,
    new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_,
    new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_,
    new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_,
    new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_,
    new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_,
    new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_,
    new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_,
    new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_,
    new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8665_,
    new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_,
    new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_,
    new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_,
    new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_,
    new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_,
    new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_, new_n8701_,
    new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_,
    new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_,
    new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_,
    new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8725_, new_n8726_,
    new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_, new_n8732_,
    new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_, new_n8738_,
    new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_, new_n8744_,
    new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8751_,
    new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_,
    new_n8758_, new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_,
    new_n8764_, new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_,
    new_n8770_, new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_,
    new_n8776_, new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_,
    new_n8782_, new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_,
    new_n8788_, new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_,
    new_n8794_, new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_,
    new_n8800_, new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_,
    new_n8806_, new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_,
    new_n8812_, new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_,
    new_n8818_, new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_,
    new_n8824_, new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_,
    new_n8830_, new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_,
    new_n8836_, new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_,
    new_n8842_, new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_,
    new_n8848_, new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_,
    new_n8854_, new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_,
    new_n8860_, new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_,
    new_n8866_, new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_,
    new_n8872_, new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8877_,
    new_n8878_, new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_,
    new_n8884_, new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_,
    new_n8890_, new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_,
    new_n8896_, new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_,
    new_n8902_, new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_,
    new_n8908_, new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_,
    new_n8914_, new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_,
    new_n8920_, new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_,
    new_n8926_, new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_,
    new_n8932_, new_n8933_, new_n8934_, new_n8935_, new_n8939_, new_n8940_,
    new_n8941_, new_n8942_, new_n8946_, new_n8947_, new_n8948_, new_n8949_,
    new_n8950_, new_n8951_, new_n8952_, new_n8953_, new_n8954_, new_n8955_,
    new_n8956_, new_n8957_, new_n8958_, new_n8959_, new_n8960_, new_n8961_,
    new_n8962_, new_n8963_, new_n8964_, new_n8965_, new_n8966_, new_n8967_,
    new_n8968_, new_n8969_, new_n8970_, new_n8971_, new_n8972_, new_n8973_,
    new_n8974_, new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_,
    new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_,
    new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_,
    new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_,
    new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_,
    new_n9004_, new_n9005_, new_n9006_, new_n9007_, new_n9008_, new_n9009_,
    new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_,
    new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_,
    new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_,
    new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_,
    new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_, new_n9039_,
    new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_, new_n9045_,
    new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_, new_n9051_,
    new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_,
    new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_, new_n9063_,
    new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_, new_n9069_,
    new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_, new_n9075_,
    new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_,
    new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_,
    new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_,
    new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_,
    new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9105_,
    new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_, new_n9111_,
    new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_,
    new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_, new_n9123_,
    new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_, new_n9129_,
    new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_, new_n9135_,
    new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_,
    new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_,
    new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_,
    new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_,
    new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_,
    new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_,
    new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_,
    new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_,
    new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_,
    new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_,
    new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9208_,
    new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_,
    new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_, new_n9220_,
    new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_,
    new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_, new_n9232_,
    new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_, new_n9238_,
    new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_, new_n9244_,
    new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_, new_n9250_,
    new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_,
    new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_,
    new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_,
    new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_,
    new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_,
    new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_,
    new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_,
    new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_,
    new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_,
    new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_,
    new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_,
    new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_,
    new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_,
    new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_,
    new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_,
    new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_,
    new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_,
    new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_,
    new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_,
    new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_,
    new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_,
    new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_,
    new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_,
    new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_,
    new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_,
    new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_,
    new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_,
    new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_,
    new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_,
    new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_,
    new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_,
    new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_,
    new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_,
    new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_,
    new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_,
    new_n9461_, new_n9462_, new_n9464_, new_n9465_, new_n9466_, new_n9467_,
    new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_,
    new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_,
    new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_,
    new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_,
    new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_,
    new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_,
    new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_,
    new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_,
    new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_,
    new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_,
    new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_,
    new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_,
    new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_,
    new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_,
    new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_,
    new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_,
    new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_,
    new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_,
    new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_,
    new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_,
    new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_,
    new_n9732_, new_n9733_, new_n9734_, new_n9736_, new_n9737_, new_n9738_,
    new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_,
    new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_,
    new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_,
    new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_,
    new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_,
    new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_,
    new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_,
    new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_,
    new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_,
    new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_,
    new_n9799_, new_n9800_, new_n9805_, new_n9806_, new_n9807_, new_n9808_,
    new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_,
    new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_,
    new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_,
    new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_,
    new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_,
    new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_,
    new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_,
    new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_,
    new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_,
    new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_,
    new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_,
    new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_,
    new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_,
    new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_,
    new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_,
    new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_,
    new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_,
    new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_,
    new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_,
    new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_,
    new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_,
    new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_,
    new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_,
    new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_,
    new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_,
    new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_,
    new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_,
    new_n9971_, new_n9972_, new_n9973_, new_n9975_, new_n9976_, new_n9977_,
    new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10464_, new_n10465_, new_n10466_,
    new_n10467_, new_n10468_, new_n10469_, new_n10470_, new_n10471_,
    new_n10472_, new_n10473_, new_n10474_, new_n10475_, new_n10476_,
    new_n10477_, new_n10478_, new_n10479_, new_n10480_, new_n10481_,
    new_n10482_, new_n10483_, new_n10484_, new_n10485_, new_n10486_,
    new_n10487_, new_n10488_, new_n10489_, new_n10490_, new_n10491_,
    new_n10492_, new_n10493_, new_n10494_, new_n10495_, new_n10496_,
    new_n10497_, new_n10498_, new_n10499_, new_n10500_, new_n10501_,
    new_n10502_, new_n10503_, new_n10504_, new_n10505_, new_n10506_,
    new_n10507_, new_n10508_, new_n10509_, new_n10510_, new_n10511_,
    new_n10512_, new_n10513_, new_n10514_, new_n10515_, new_n10516_,
    new_n10517_, new_n10518_, new_n10519_, new_n10520_, new_n10521_,
    new_n10522_, new_n10523_, new_n10524_, new_n10525_, new_n10526_,
    new_n10527_, new_n10528_, new_n10529_, new_n10530_, new_n10531_,
    new_n10532_, new_n10533_, new_n10534_, new_n10535_, new_n10536_,
    new_n10537_, new_n10538_, new_n10539_, new_n10540_, new_n10541_,
    new_n10542_, new_n10543_, new_n10544_, new_n10545_, new_n10546_,
    new_n10547_, new_n10548_, new_n10549_, new_n10550_, new_n10551_,
    new_n10552_, new_n10553_, new_n10554_, new_n10555_, new_n10556_,
    new_n10557_, new_n10558_, new_n10559_, new_n10560_, new_n10561_,
    new_n10562_, new_n10563_, new_n10564_, new_n10565_, new_n10566_,
    new_n10567_, new_n10568_, new_n10569_, new_n10570_, new_n10571_,
    new_n10572_, new_n10573_, new_n10574_, new_n10575_, new_n10576_,
    new_n10577_, new_n10578_, new_n10579_, new_n10580_, new_n10581_,
    new_n10582_, new_n10583_, new_n10584_, new_n10585_, new_n10586_,
    new_n10587_, new_n10588_, new_n10589_, new_n10590_, new_n10591_,
    new_n10592_, new_n10593_, new_n10594_, new_n10595_, new_n10596_,
    new_n10597_, new_n10598_, new_n10599_, new_n10600_, new_n10601_,
    new_n10602_, new_n10603_, new_n10604_, new_n10605_, new_n10606_,
    new_n10607_, new_n10608_, new_n10609_, new_n10610_, new_n10611_,
    new_n10612_, new_n10613_, new_n10614_, new_n10615_, new_n10616_,
    new_n10617_, new_n10618_, new_n10619_, new_n10620_, new_n10621_,
    new_n10622_, new_n10623_, new_n10624_, new_n10625_, new_n10626_,
    new_n10627_, new_n10628_, new_n10629_, new_n10630_, new_n10631_,
    new_n10632_, new_n10633_, new_n10634_, new_n10635_, new_n10636_,
    new_n10637_, new_n10638_, new_n10639_, new_n10640_, new_n10641_,
    new_n10642_, new_n10643_, new_n10644_, new_n10645_, new_n10646_,
    new_n10647_, new_n10648_, new_n10649_, new_n10650_, new_n10651_,
    new_n10652_, new_n10653_, new_n10654_, new_n10655_, new_n10656_,
    new_n10657_, new_n10658_, new_n10659_, new_n10660_, new_n10661_,
    new_n10662_, new_n10663_, new_n10664_, new_n10665_, new_n10666_,
    new_n10667_, new_n10668_, new_n10669_, new_n10670_, new_n10671_,
    new_n10672_, new_n10673_, new_n10674_, new_n10675_, new_n10676_,
    new_n10677_, new_n10678_, new_n10679_, new_n10680_, new_n10681_,
    new_n10682_, new_n10683_, new_n10684_, new_n10685_, new_n10686_,
    new_n10687_, new_n10688_, new_n10689_, new_n10690_, new_n10691_,
    new_n10692_, new_n10693_, new_n10694_, new_n10695_, new_n10696_,
    new_n10697_, new_n10698_, new_n10699_, new_n10700_, new_n10701_,
    new_n10702_, new_n10704_, new_n10705_, new_n10706_, new_n10707_,
    new_n10708_, new_n10709_, new_n10710_, new_n10711_, new_n10712_,
    new_n10713_, new_n10714_, new_n10715_, new_n10716_, new_n10717_,
    new_n10718_, new_n10719_, new_n10720_, new_n10721_, new_n10722_,
    new_n10723_, new_n10724_, new_n10725_, new_n10726_, new_n10727_,
    new_n10728_, new_n10729_, new_n10730_, new_n10731_, new_n10732_,
    new_n10733_, new_n10734_, new_n10735_, new_n10736_, new_n10737_,
    new_n10738_, new_n10739_, new_n10740_, new_n10741_, new_n10742_,
    new_n10743_, new_n10744_, new_n10745_, new_n10746_, new_n10747_,
    new_n10748_, new_n10749_, new_n10750_, new_n10751_, new_n10752_,
    new_n10753_, new_n10754_, new_n10755_, new_n10756_, new_n10757_,
    new_n10758_, new_n10759_, new_n10760_, new_n10761_, new_n10762_,
    new_n10763_, new_n10764_, new_n10765_, new_n10766_, new_n10767_,
    new_n10768_, new_n10769_, new_n10770_, new_n10771_, new_n10772_,
    new_n10773_, new_n10774_, new_n10775_, new_n10776_, new_n10777_,
    new_n10778_, new_n10779_, new_n10780_, new_n10781_, new_n10782_,
    new_n10783_, new_n10784_, new_n10785_, new_n10786_, new_n10787_,
    new_n10788_, new_n10789_, new_n10790_, new_n10791_, new_n10792_,
    new_n10793_, new_n10794_, new_n10795_, new_n10796_, new_n10797_,
    new_n10798_, new_n10799_, new_n10800_, new_n10801_, new_n10802_,
    new_n10803_, new_n10804_, new_n10805_, new_n10806_, new_n10807_,
    new_n10808_, new_n10809_, new_n10810_, new_n10811_, new_n10812_,
    new_n10813_, new_n10814_, new_n10815_, new_n10816_, new_n10817_,
    new_n10818_, new_n10819_, new_n10820_, new_n10821_, new_n10822_,
    new_n10823_, new_n10824_, new_n10825_, new_n10826_, new_n10827_,
    new_n10828_, new_n10829_, new_n10830_, new_n10831_, new_n10832_,
    new_n10833_, new_n10834_, new_n10835_, new_n10836_, new_n10837_,
    new_n10838_, new_n10839_, new_n10840_, new_n10841_, new_n10842_,
    new_n10843_, new_n10844_, new_n10845_, new_n10846_, new_n10847_,
    new_n10848_, new_n10849_, new_n10850_, new_n10851_, new_n10852_,
    new_n10853_, new_n10854_, new_n10855_, new_n10856_, new_n10857_,
    new_n10858_, new_n10859_, new_n10860_, new_n10861_, new_n10862_,
    new_n10863_, new_n10864_, new_n10865_, new_n10866_, new_n10867_,
    new_n10868_, new_n10869_, new_n10870_, new_n10871_, new_n10872_,
    new_n10873_, new_n10874_, new_n10875_, new_n10876_, new_n10877_,
    new_n10878_, new_n10879_, new_n10880_, new_n10881_, new_n10882_,
    new_n10883_, new_n10884_, new_n10885_, new_n10886_, new_n10887_,
    new_n10888_, new_n10889_, new_n10890_, new_n10891_, new_n10892_,
    new_n10893_, new_n10894_, new_n10895_, new_n10896_, new_n10897_,
    new_n10898_, new_n10899_, new_n10900_, new_n10901_, new_n10902_,
    new_n10903_, new_n10904_, new_n10905_, new_n10906_, new_n10907_,
    new_n10908_, new_n10909_, new_n10910_, new_n10911_, new_n10912_,
    new_n10913_, new_n10914_, new_n10915_, new_n10916_, new_n10917_,
    new_n10918_, new_n10919_, new_n10920_, new_n10921_, new_n10922_,
    new_n10923_, new_n10924_, new_n10925_, new_n10926_, new_n10927_,
    new_n10928_, new_n10929_, new_n10930_, new_n10931_, new_n10932_,
    new_n10933_, new_n10934_, new_n10935_, new_n10936_, new_n10937_,
    new_n10938_, new_n10939_, new_n10941_, new_n10942_, new_n10943_,
    new_n10944_, new_n10945_, new_n10946_, new_n10947_, new_n10948_,
    new_n10949_, new_n10950_, new_n10951_, new_n10952_, new_n10953_,
    new_n10954_, new_n10955_, new_n10956_, new_n10957_, new_n10958_,
    new_n10959_, new_n10960_, new_n10961_, new_n10962_, new_n10963_,
    new_n10964_, new_n10965_, new_n10966_, new_n10967_, new_n10968_,
    new_n10969_, new_n10970_, new_n10971_, new_n10972_, new_n10973_,
    new_n10974_, new_n10975_, new_n10976_, new_n10977_, new_n10978_,
    new_n10979_, new_n10980_, new_n10981_, new_n10982_, new_n10983_,
    new_n10984_, new_n10985_, new_n10986_, new_n10987_, new_n10988_,
    new_n10989_, new_n10990_, new_n10991_, new_n10992_, new_n10993_,
    new_n10994_, new_n10995_, new_n10996_, new_n10997_, new_n10998_,
    new_n10999_, new_n11000_, new_n11001_, new_n11002_, new_n11003_,
    new_n11004_, new_n11005_, new_n11006_, new_n11007_, new_n11008_,
    new_n11009_, new_n11010_, new_n11011_, new_n11012_, new_n11013_,
    new_n11014_, new_n11015_, new_n11016_, new_n11017_, new_n11018_,
    new_n11019_, new_n11020_, new_n11021_, new_n11022_, new_n11023_,
    new_n11024_, new_n11025_, new_n11026_, new_n11027_, new_n11028_,
    new_n11029_, new_n11030_, new_n11031_, new_n11032_, new_n11033_,
    new_n11034_, new_n11035_, new_n11036_, new_n11037_, new_n11038_,
    new_n11039_, new_n11040_, new_n11041_, new_n11042_, new_n11043_,
    new_n11044_, new_n11045_, new_n11046_, new_n11047_, new_n11048_,
    new_n11049_, new_n11050_, new_n11051_, new_n11052_, new_n11053_,
    new_n11054_, new_n11055_, new_n11056_, new_n11057_, new_n11058_,
    new_n11059_, new_n11060_, new_n11061_, new_n11062_, new_n11063_,
    new_n11064_, new_n11065_, new_n11066_, new_n11067_, new_n11068_,
    new_n11069_, new_n11070_, new_n11071_, new_n11072_, new_n11073_,
    new_n11074_, new_n11075_, new_n11076_, new_n11077_, new_n11078_,
    new_n11079_, new_n11080_, new_n11081_, new_n11082_, new_n11083_,
    new_n11084_, new_n11085_, new_n11086_, new_n11087_, new_n11088_,
    new_n11089_, new_n11090_, new_n11091_, new_n11092_, new_n11093_,
    new_n11094_, new_n11095_, new_n11096_, new_n11097_, new_n11098_,
    new_n11099_, new_n11100_, new_n11101_, new_n11102_, new_n11103_,
    new_n11104_, new_n11105_, new_n11106_, new_n11107_, new_n11108_,
    new_n11109_, new_n11110_, new_n11111_, new_n11112_, new_n11113_,
    new_n11114_, new_n11115_, new_n11116_, new_n11117_, new_n11118_,
    new_n11119_, new_n11120_, new_n11121_, new_n11122_, new_n11123_,
    new_n11124_, new_n11125_, new_n11126_, new_n11127_, new_n11128_,
    new_n11129_, new_n11130_, new_n11131_, new_n11132_, new_n11133_,
    new_n11134_, new_n11135_, new_n11136_, new_n11137_, new_n11138_,
    new_n11139_, new_n11140_, new_n11141_, new_n11142_, new_n11143_,
    new_n11144_, new_n11145_, new_n11146_, new_n11147_, new_n11148_,
    new_n11149_, new_n11150_, new_n11151_, new_n11152_, new_n11154_,
    new_n11155_, new_n11156_, new_n11157_, new_n11158_, new_n11159_,
    new_n11160_, new_n11161_, new_n11162_, new_n11163_, new_n11164_,
    new_n11165_, new_n11166_, new_n11167_, new_n11168_, new_n11169_,
    new_n11170_, new_n11171_, new_n11172_, new_n11173_, new_n11174_,
    new_n11175_, new_n11176_, new_n11177_, new_n11178_, new_n11179_,
    new_n11180_, new_n11181_, new_n11182_, new_n11183_, new_n11184_,
    new_n11185_, new_n11186_, new_n11187_, new_n11188_, new_n11189_,
    new_n11190_, new_n11191_, new_n11192_, new_n11193_, new_n11194_,
    new_n11195_, new_n11196_, new_n11197_, new_n11198_, new_n11199_,
    new_n11200_, new_n11201_, new_n11202_, new_n11203_, new_n11204_,
    new_n11205_, new_n11206_, new_n11207_, new_n11208_, new_n11209_,
    new_n11210_, new_n11211_, new_n11212_, new_n11213_, new_n11214_,
    new_n11215_, new_n11216_, new_n11217_, new_n11218_, new_n11219_,
    new_n11220_, new_n11221_, new_n11222_, new_n11223_, new_n11224_,
    new_n11225_, new_n11226_, new_n11227_, new_n11228_, new_n11229_,
    new_n11230_, new_n11231_, new_n11232_, new_n11233_, new_n11234_,
    new_n11235_, new_n11236_, new_n11237_, new_n11238_, new_n11239_,
    new_n11240_, new_n11241_, new_n11242_, new_n11243_, new_n11244_,
    new_n11245_, new_n11246_, new_n11247_, new_n11248_, new_n11249_,
    new_n11250_, new_n11251_, new_n11252_, new_n11253_, new_n11254_,
    new_n11255_, new_n11256_, new_n11257_, new_n11258_, new_n11259_,
    new_n11260_, new_n11261_, new_n11262_, new_n11263_, new_n11264_,
    new_n11265_, new_n11266_, new_n11267_, new_n11268_, new_n11269_,
    new_n11270_, new_n11271_, new_n11272_, new_n11273_, new_n11274_,
    new_n11275_, new_n11276_, new_n11277_, new_n11278_, new_n11279_,
    new_n11280_, new_n11281_, new_n11282_, new_n11283_, new_n11284_,
    new_n11285_, new_n11286_, new_n11287_, new_n11288_, new_n11289_,
    new_n11290_, new_n11291_, new_n11292_, new_n11293_, new_n11294_,
    new_n11295_, new_n11296_, new_n11297_, new_n11298_, new_n11299_,
    new_n11300_, new_n11301_, new_n11302_, new_n11303_, new_n11304_,
    new_n11305_, new_n11306_, new_n11307_, new_n11308_, new_n11309_,
    new_n11310_, new_n11311_, new_n11312_, new_n11313_, new_n11314_,
    new_n11315_, new_n11316_, new_n11317_, new_n11318_, new_n11319_,
    new_n11320_, new_n11321_, new_n11322_, new_n11323_, new_n11324_,
    new_n11325_, new_n11326_, new_n11327_, new_n11328_, new_n11329_,
    new_n11330_, new_n11331_, new_n11332_, new_n11333_, new_n11334_,
    new_n11335_, new_n11336_, new_n11337_, new_n11338_, new_n11339_,
    new_n11340_, new_n11341_, new_n11342_, new_n11343_, new_n11344_,
    new_n11345_, new_n11346_, new_n11347_, new_n11348_, new_n11349_,
    new_n11350_, new_n11351_, new_n11352_, new_n11353_, new_n11354_,
    new_n11355_, new_n11356_, new_n11357_, new_n11358_, new_n11359_,
    new_n11360_, new_n11361_, new_n11362_, new_n11363_, new_n11364_,
    new_n11365_, new_n11366_, new_n11367_, new_n11368_, new_n11369_,
    new_n11370_, new_n11371_, new_n11372_, new_n11374_, new_n11375_,
    new_n11376_, new_n11377_, new_n11378_, new_n11379_, new_n11380_,
    new_n11381_, new_n11382_, new_n11383_, new_n11384_, new_n11385_,
    new_n11386_, new_n11387_, new_n11388_, new_n11389_, new_n11390_,
    new_n11391_, new_n11392_, new_n11393_, new_n11394_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11421_, new_n11422_, new_n11423_, new_n11424_, new_n11425_,
    new_n11426_, new_n11427_, new_n11428_, new_n11429_, new_n11430_,
    new_n11431_, new_n11432_, new_n11433_, new_n11434_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11447_, new_n11448_, new_n11449_, new_n11450_,
    new_n11451_, new_n11452_, new_n11453_, new_n11454_, new_n11455_,
    new_n11456_, new_n11457_, new_n11458_, new_n11459_, new_n11460_,
    new_n11461_, new_n11462_, new_n11463_, new_n11464_, new_n11465_,
    new_n11466_, new_n11467_, new_n11468_, new_n11469_, new_n11470_,
    new_n11471_, new_n11472_, new_n11473_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11491_, new_n11492_, new_n11493_, new_n11494_, new_n11495_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11579_, new_n11580_, new_n11581_,
    new_n11582_, new_n11583_, new_n11584_, new_n11585_, new_n11586_,
    new_n11587_, new_n11588_, new_n11589_, new_n11590_, new_n11591_,
    new_n11592_, new_n11593_, new_n11594_, new_n11595_, new_n11596_,
    new_n11597_, new_n11598_, new_n11599_, new_n11600_, new_n11601_,
    new_n11602_, new_n11603_, new_n11604_, new_n11605_, new_n11606_,
    new_n11607_, new_n11608_, new_n11609_, new_n11610_, new_n11611_,
    new_n11612_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11667_, new_n11668_, new_n11669_, new_n11670_, new_n11671_,
    new_n11672_, new_n11673_, new_n11674_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11728_, new_n11729_, new_n11730_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11740_, new_n11741_,
    new_n11742_, new_n11743_, new_n11744_, new_n11745_, new_n11746_,
    new_n11747_, new_n11748_, new_n11749_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11762_, new_n11763_, new_n11764_, new_n11765_, new_n11766_,
    new_n11767_, new_n11768_, new_n11769_, new_n11770_, new_n11771_,
    new_n11772_, new_n11773_, new_n11774_, new_n11775_, new_n11776_,
    new_n11777_, new_n11778_, new_n11779_, new_n11780_, new_n11781_,
    new_n11782_, new_n11783_, new_n11784_, new_n11785_, new_n11786_,
    new_n11787_, new_n11788_, new_n11789_, new_n11791_, new_n11792_,
    new_n11793_, new_n11794_, new_n11795_, new_n11796_, new_n11797_,
    new_n11798_, new_n11799_, new_n11800_, new_n11801_, new_n11802_,
    new_n11803_, new_n11804_, new_n11805_, new_n11806_, new_n11807_,
    new_n11808_, new_n11809_, new_n11810_, new_n11811_, new_n11812_,
    new_n11813_, new_n11814_, new_n11815_, new_n11816_, new_n11817_,
    new_n11818_, new_n11819_, new_n11820_, new_n11821_, new_n11822_,
    new_n11823_, new_n11824_, new_n11825_, new_n11826_, new_n11827_,
    new_n11828_, new_n11829_, new_n11830_, new_n11831_, new_n11832_,
    new_n11833_, new_n11834_, new_n11835_, new_n11836_, new_n11837_,
    new_n11838_, new_n11839_, new_n11840_, new_n11841_, new_n11842_,
    new_n11843_, new_n11844_, new_n11845_, new_n11846_, new_n11847_,
    new_n11848_, new_n11849_, new_n11850_, new_n11851_, new_n11852_,
    new_n11853_, new_n11854_, new_n11855_, new_n11856_, new_n11857_,
    new_n11858_, new_n11859_, new_n11860_, new_n11861_, new_n11862_,
    new_n11863_, new_n11864_, new_n11865_, new_n11866_, new_n11867_,
    new_n11868_, new_n11869_, new_n11870_, new_n11871_, new_n11872_,
    new_n11873_, new_n11874_, new_n11875_, new_n11876_, new_n11877_,
    new_n11878_, new_n11879_, new_n11880_, new_n11881_, new_n11882_,
    new_n11883_, new_n11884_, new_n11885_, new_n11886_, new_n11887_,
    new_n11888_, new_n11889_, new_n11890_, new_n11891_, new_n11892_,
    new_n11893_, new_n11894_, new_n11895_, new_n11896_, new_n11897_,
    new_n11898_, new_n11899_, new_n11900_, new_n11901_, new_n11902_,
    new_n11903_, new_n11904_, new_n11905_, new_n11906_, new_n11907_,
    new_n11908_, new_n11909_, new_n11910_, new_n11911_, new_n11912_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11918_, new_n11919_, new_n11920_, new_n11921_, new_n11922_,
    new_n11923_, new_n11924_, new_n11925_, new_n11926_, new_n11927_,
    new_n11928_, new_n11929_, new_n11930_, new_n11931_, new_n11932_,
    new_n11933_, new_n11934_, new_n11935_, new_n11936_, new_n11937_,
    new_n11938_, new_n11939_, new_n11940_, new_n11941_, new_n11942_,
    new_n11943_, new_n11944_, new_n11945_, new_n11946_, new_n11947_,
    new_n11948_, new_n11949_, new_n11950_, new_n11951_, new_n11952_,
    new_n11953_, new_n11954_, new_n11955_, new_n11956_, new_n11957_,
    new_n11959_, new_n11960_, new_n11961_, new_n11962_, new_n11963_,
    new_n11964_, new_n11965_, new_n11966_, new_n11967_, new_n11968_,
    new_n11969_, new_n11970_, new_n11971_, new_n11972_, new_n11973_,
    new_n11974_, new_n11975_, new_n11976_, new_n11977_, new_n11978_,
    new_n11979_, new_n11980_, new_n11981_, new_n11982_, new_n11983_,
    new_n11984_, new_n11985_, new_n11986_, new_n11987_, new_n11988_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11996_, new_n11997_, new_n11998_,
    new_n11999_, new_n12000_, new_n12001_, new_n12002_, new_n12003_,
    new_n12004_, new_n12005_, new_n12006_, new_n12008_, new_n12009_,
    new_n12010_, new_n12011_, new_n12012_, new_n12013_, new_n12014_,
    new_n12015_, new_n12016_, new_n12017_, new_n12018_, new_n12019_,
    new_n12020_, new_n12021_, new_n12022_, new_n12023_, new_n12024_,
    new_n12025_, new_n12026_, new_n12027_, new_n12028_, new_n12029_,
    new_n12030_, new_n12031_, new_n12032_, new_n12033_, new_n12034_,
    new_n12035_, new_n12036_, new_n12037_, new_n12038_, new_n12039_,
    new_n12040_, new_n12041_, new_n12042_, new_n12043_, new_n12044_,
    new_n12045_, new_n12046_, new_n12047_, new_n12048_, new_n12049_,
    new_n12050_, new_n12051_, new_n12052_, new_n12053_, new_n12054_,
    new_n12055_, new_n12056_, new_n12057_, new_n12058_, new_n12059_,
    new_n12060_, new_n12061_, new_n12062_, new_n12063_, new_n12064_,
    new_n12065_, new_n12066_, new_n12067_, new_n12068_, new_n12069_,
    new_n12070_, new_n12071_, new_n12072_, new_n12073_, new_n12074_,
    new_n12075_, new_n12076_, new_n12077_, new_n12078_, new_n12079_,
    new_n12080_, new_n12081_, new_n12082_, new_n12083_, new_n12084_,
    new_n12085_, new_n12086_, new_n12087_, new_n12088_, new_n12089_,
    new_n12090_, new_n12091_, new_n12092_, new_n12093_, new_n12094_,
    new_n12095_, new_n12096_, new_n12097_, new_n12098_, new_n12099_,
    new_n12100_, new_n12101_, new_n12102_, new_n12103_, new_n12104_,
    new_n12105_, new_n12106_, new_n12107_, new_n12108_, new_n12109_,
    new_n12110_, new_n12111_, new_n12112_, new_n12113_, new_n12114_,
    new_n12115_, new_n12116_, new_n12117_, new_n12118_, new_n12119_,
    new_n12120_, new_n12121_, new_n12122_, new_n12123_, new_n12124_,
    new_n12125_, new_n12126_, new_n12127_, new_n12128_, new_n12129_,
    new_n12130_, new_n12131_, new_n12132_, new_n12133_, new_n12134_,
    new_n12135_, new_n12136_, new_n12137_, new_n12138_, new_n12139_,
    new_n12140_, new_n12141_, new_n12142_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12156_, new_n12157_, new_n12158_, new_n12159_,
    new_n12160_, new_n12161_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12171_, new_n12172_, new_n12173_, new_n12174_,
    new_n12175_, new_n12176_, new_n12177_, new_n12178_, new_n12179_,
    new_n12180_, new_n12181_, new_n12182_, new_n12183_, new_n12184_,
    new_n12185_, new_n12186_, new_n12187_, new_n12188_, new_n12189_,
    new_n12190_, new_n12191_, new_n12192_, new_n12193_, new_n12194_,
    new_n12195_, new_n12196_, new_n12197_, new_n12198_, new_n12199_,
    new_n12200_, new_n12201_, new_n12202_, new_n12203_, new_n12204_,
    new_n12205_, new_n12206_, new_n12207_, new_n12208_, new_n12210_,
    new_n12211_, new_n12212_, new_n12213_, new_n12214_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12243_, new_n12244_, new_n12245_,
    new_n12246_, new_n12247_, new_n12248_, new_n12249_, new_n12250_,
    new_n12251_, new_n12252_, new_n12253_, new_n12254_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12307_, new_n12308_, new_n12309_, new_n12310_,
    new_n12311_, new_n12312_, new_n12313_, new_n12314_, new_n12315_,
    new_n12316_, new_n12317_, new_n12318_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12323_, new_n12324_, new_n12325_,
    new_n12326_, new_n12327_, new_n12328_, new_n12329_, new_n12330_,
    new_n12331_, new_n12332_, new_n12333_, new_n12337_, new_n12338_,
    new_n12339_, new_n12340_, new_n12341_, new_n12342_, new_n12343_,
    new_n12344_, new_n12345_, new_n12346_, new_n12347_, new_n12348_,
    new_n12349_, new_n12350_, new_n12351_, new_n12352_, new_n12353_,
    new_n12354_, new_n12355_, new_n12356_, new_n12357_, new_n12358_,
    new_n12359_, new_n12360_, new_n12361_, new_n12362_, new_n12363_,
    new_n12364_, new_n12365_, new_n12366_, new_n12367_, new_n12368_,
    new_n12369_, new_n12370_, new_n12371_, new_n12372_, new_n12373_,
    new_n12374_, new_n12375_, new_n12376_, new_n12377_, new_n12378_,
    new_n12379_, new_n12380_, new_n12381_, new_n12382_, new_n12383_,
    new_n12384_, new_n12385_, new_n12386_, new_n12387_, new_n12388_,
    new_n12389_, new_n12390_, new_n12391_, new_n12392_, new_n12393_,
    new_n12394_, new_n12395_, new_n12396_, new_n12397_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12438_, new_n12439_,
    new_n12440_, new_n12441_, new_n12442_, new_n12443_, new_n12444_,
    new_n12445_, new_n12446_, new_n12447_, new_n12448_, new_n12449_,
    new_n12450_, new_n12451_, new_n12452_, new_n12453_, new_n12454_,
    new_n12455_, new_n12456_, new_n12457_, new_n12458_, new_n12459_,
    new_n12460_, new_n12461_, new_n12462_, new_n12463_, new_n12464_,
    new_n12465_, new_n12466_, new_n12467_, new_n12468_, new_n12469_,
    new_n12470_, new_n12471_, new_n12472_, new_n12473_, new_n12474_,
    new_n12475_, new_n12476_, new_n12477_, new_n12478_, new_n12479_,
    new_n12480_, new_n12481_, new_n12482_, new_n12483_, new_n12484_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12491_, new_n12492_, new_n12493_, new_n12494_,
    new_n12495_, new_n12496_, new_n12497_, new_n12498_, new_n12499_,
    new_n12500_, new_n12501_, new_n12502_, new_n12503_, new_n12504_,
    new_n12505_, new_n12506_, new_n12507_, new_n12508_, new_n12509_,
    new_n12510_, new_n12511_, new_n12512_, new_n12513_, new_n12514_,
    new_n12515_, new_n12516_, new_n12517_, new_n12518_, new_n12519_,
    new_n12520_, new_n12521_, new_n12522_, new_n12523_, new_n12524_,
    new_n12525_, new_n12526_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12532_, new_n12533_, new_n12534_,
    new_n12535_, new_n12536_, new_n12537_, new_n12538_, new_n12539_,
    new_n12540_, new_n12541_, new_n12542_, new_n12543_, new_n12544_,
    new_n12545_, new_n12546_, new_n12547_, new_n12548_, new_n12549_,
    new_n12550_, new_n12551_, new_n12552_, new_n12553_, new_n12554_,
    new_n12555_, new_n12556_, new_n12557_, new_n12558_, new_n12559_,
    new_n12560_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12604_, new_n12605_, new_n12606_,
    new_n12607_, new_n12608_, new_n12609_, new_n12610_, new_n12611_,
    new_n12612_, new_n12613_, new_n12614_, new_n12615_, new_n12616_,
    new_n12617_, new_n12618_, new_n12619_, new_n12620_, new_n12621_,
    new_n12622_, new_n12623_, new_n12624_, new_n12625_, new_n12626_,
    new_n12627_, new_n12628_, new_n12629_, new_n12630_, new_n12631_,
    new_n12632_, new_n12633_, new_n12634_, new_n12635_, new_n12636_,
    new_n12637_, new_n12638_, new_n12639_, new_n12640_, new_n12641_,
    new_n12642_, new_n12643_, new_n12644_, new_n12645_, new_n12646_,
    new_n12647_, new_n12648_, new_n12649_, new_n12650_, new_n12651_,
    new_n12652_, new_n12653_, new_n12654_, new_n12655_, new_n12656_,
    new_n12657_, new_n12658_, new_n12659_, new_n12660_, new_n12661_,
    new_n12662_, new_n12663_, new_n12664_, new_n12665_, new_n12666_,
    new_n12667_, new_n12668_, new_n12669_, new_n12670_, new_n12671_,
    new_n12672_, new_n12673_, new_n12674_, new_n12675_, new_n12676_,
    new_n12677_, new_n12678_, new_n12679_, new_n12680_, new_n12681_,
    new_n12682_, new_n12683_, new_n12684_, new_n12685_, new_n12686_,
    new_n12687_, new_n12688_, new_n12689_, new_n12690_, new_n12691_,
    new_n12692_, new_n12693_, new_n12694_, new_n12695_, new_n12696_,
    new_n12697_, new_n12698_, new_n12699_, new_n12700_, new_n12701_,
    new_n12702_, new_n12703_, new_n12704_, new_n12705_, new_n12706_,
    new_n12707_, new_n12708_, new_n12709_, new_n12710_, new_n12711_,
    new_n12712_, new_n12713_, new_n12714_, new_n12715_, new_n12716_,
    new_n12717_, new_n12718_, new_n12719_, new_n12720_, new_n12721_,
    new_n12722_, new_n12723_, new_n12724_, new_n12725_, new_n12726_,
    new_n12727_, new_n12728_, new_n12729_, new_n12730_, new_n12731_,
    new_n12732_, new_n12733_, new_n12734_, new_n12735_, new_n12736_,
    new_n12737_, new_n12738_, new_n12739_, new_n12740_, new_n12741_,
    new_n12742_, new_n12743_, new_n12744_, new_n12745_, new_n12746_,
    new_n12747_, new_n12748_, new_n12749_, new_n12750_, new_n12751_,
    new_n12752_, new_n12753_, new_n12754_, new_n12755_, new_n12756_,
    new_n12757_, new_n12758_, new_n12759_, new_n12760_, new_n12761_,
    new_n12762_, new_n12763_, new_n12764_, new_n12765_, new_n12766_,
    new_n12767_, new_n12768_, new_n12769_, new_n12770_, new_n12771_,
    new_n12772_, new_n12773_, new_n12774_, new_n12775_, new_n12776_,
    new_n12777_, new_n12778_, new_n12779_, new_n12780_, new_n12781_,
    new_n12782_, new_n12783_, new_n12784_, new_n12785_, new_n12787_,
    new_n12788_, new_n12789_, new_n12790_, new_n12792_, new_n12793_,
    new_n12794_, new_n12795_, new_n12796_, new_n12797_, new_n12798_,
    new_n12799_, new_n12800_, new_n12801_, new_n12802_, new_n12803_,
    new_n12804_, new_n12805_, new_n12806_, new_n12807_, new_n12808_,
    new_n12809_, new_n12810_, new_n12811_, new_n12812_, new_n12813_,
    new_n12814_, new_n12815_, new_n12816_, new_n12817_, new_n12818_,
    new_n12819_, new_n12820_, new_n12821_, new_n12822_, new_n12823_,
    new_n12824_, new_n12825_, new_n12826_, new_n12827_, new_n12828_,
    new_n12829_, new_n12830_, new_n12831_, new_n12832_, new_n12833_,
    new_n12834_, new_n12835_, new_n12836_, new_n12837_, new_n12838_,
    new_n12839_, new_n12840_, new_n12841_, new_n12842_, new_n12843_,
    new_n12844_, new_n12845_, new_n12846_, new_n12847_, new_n12848_,
    new_n12849_, new_n12850_, new_n12851_, new_n12852_, new_n12853_,
    new_n12854_, new_n12855_, new_n12856_, new_n12857_, new_n12858_,
    new_n12859_, new_n12860_, new_n12861_, new_n12862_, new_n12863_,
    new_n12864_, new_n12865_, new_n12866_, new_n12867_, new_n12868_,
    new_n12869_, new_n12870_, new_n12871_, new_n12872_, new_n12873_,
    new_n12874_, new_n12875_, new_n12876_, new_n12877_, new_n12878_,
    new_n12879_, new_n12880_, new_n12881_, new_n12882_, new_n12883_,
    new_n12884_, new_n12885_, new_n12886_, new_n12887_, new_n12888_,
    new_n12889_, new_n12890_, new_n12891_, new_n12892_, new_n12893_,
    new_n12894_, new_n12895_, new_n12896_, new_n12897_, new_n12898_,
    new_n12899_, new_n12900_, new_n12901_, new_n12902_, new_n12903_,
    new_n12904_, new_n12905_, new_n12906_, new_n12907_, new_n12908_,
    new_n12909_, new_n12910_, new_n12911_, new_n12912_, new_n12913_,
    new_n12914_, new_n12915_, new_n12916_, new_n12917_, new_n12918_,
    new_n12919_, new_n12920_, new_n12921_, new_n12922_, new_n12923_,
    new_n12924_, new_n12925_, new_n12926_, new_n12927_, new_n12928_,
    new_n12929_, new_n12930_, new_n12931_, new_n12932_, new_n12933_,
    new_n12934_, new_n12935_, new_n12936_, new_n12937_, new_n12938_,
    new_n12939_, new_n12940_, new_n12941_, new_n12942_, new_n12943_,
    new_n12944_, new_n12945_, new_n12946_, new_n12947_, new_n12948_,
    new_n12949_, new_n12950_, new_n12951_, new_n12952_, new_n12953_,
    new_n12954_, new_n12955_, new_n12956_, new_n12957_, new_n12958_,
    new_n12959_, new_n12960_, new_n12961_, new_n12962_, new_n12964_,
    new_n12965_, new_n12969_, new_n12970_, new_n12971_, new_n12972_,
    new_n12973_, new_n12974_, new_n12975_, new_n12976_, new_n12977_,
    new_n12978_, new_n12979_, new_n12980_, new_n12981_, new_n12982_,
    new_n12983_, new_n12984_, new_n12985_, new_n12986_, new_n12987_,
    new_n12988_, new_n12989_, new_n12990_, new_n12991_, new_n12992_,
    new_n12993_, new_n12994_, new_n12995_, new_n12996_, new_n12997_,
    new_n12998_, new_n12999_, new_n13000_, new_n13001_, new_n13002_,
    new_n13003_, new_n13004_, new_n13005_, new_n13006_, new_n13007_,
    new_n13008_, new_n13009_, new_n13010_, new_n13011_, new_n13012_,
    new_n13013_, new_n13014_, new_n13015_, new_n13016_, new_n13017_,
    new_n13018_, new_n13019_, new_n13020_, new_n13021_, new_n13022_,
    new_n13023_, new_n13024_, new_n13025_, new_n13026_, new_n13027_,
    new_n13028_, new_n13029_, new_n13030_, new_n13031_, new_n13032_,
    new_n13033_, new_n13034_, new_n13035_, new_n13036_, new_n13037_,
    new_n13038_, new_n13039_, new_n13040_, new_n13041_, new_n13042_,
    new_n13043_, new_n13044_, new_n13045_, new_n13046_, new_n13047_,
    new_n13048_, new_n13049_, new_n13050_, new_n13051_, new_n13052_,
    new_n13053_, new_n13054_, new_n13055_, new_n13056_, new_n13057_,
    new_n13058_, new_n13059_, new_n13060_, new_n13061_, new_n13062_,
    new_n13063_, new_n13064_, new_n13065_, new_n13066_, new_n13067_,
    new_n13068_, new_n13069_, new_n13070_, new_n13071_, new_n13072_,
    new_n13073_, new_n13074_, new_n13075_, new_n13076_, new_n13077_,
    new_n13078_, new_n13079_, new_n13080_, new_n13081_, new_n13082_,
    new_n13083_, new_n13084_, new_n13085_, new_n13086_, new_n13087_,
    new_n13088_, new_n13089_, new_n13090_, new_n13091_, new_n13092_,
    new_n13093_, new_n13094_, new_n13095_, new_n13096_, new_n13097_,
    new_n13098_, new_n13099_, new_n13100_, new_n13101_, new_n13102_,
    new_n13103_, new_n13104_, new_n13105_, new_n13106_, new_n13107_,
    new_n13108_, new_n13109_, new_n13110_, new_n13111_, new_n13112_,
    new_n13113_, new_n13114_, new_n13115_, new_n13116_, new_n13117_,
    new_n13118_, new_n13119_, new_n13120_, new_n13121_, new_n13122_,
    new_n13123_, new_n13124_, new_n13125_, new_n13126_, new_n13127_,
    new_n13128_, new_n13129_, new_n13130_, new_n13131_, new_n13132_,
    new_n13133_, new_n13134_, new_n13135_, new_n13136_, new_n13137_,
    new_n13138_, new_n13139_, new_n13140_, new_n13141_, new_n13142_,
    new_n13143_, new_n13145_, new_n13146_, new_n13147_, new_n13148_,
    new_n13149_, new_n13150_, new_n13151_, new_n13152_, new_n13153_,
    new_n13154_, new_n13155_, new_n13156_, new_n13157_, new_n13158_,
    new_n13159_, new_n13160_, new_n13161_, new_n13162_, new_n13163_,
    new_n13164_, new_n13165_, new_n13166_, new_n13167_, new_n13168_,
    new_n13169_, new_n13170_, new_n13171_, new_n13172_, new_n13173_,
    new_n13174_, new_n13175_, new_n13176_, new_n13177_, new_n13178_,
    new_n13179_, new_n13180_, new_n13181_, new_n13182_, new_n13183_,
    new_n13184_, new_n13185_, new_n13186_, new_n13187_, new_n13188_,
    new_n13189_, new_n13190_, new_n13191_, new_n13192_, new_n13193_,
    new_n13194_, new_n13195_, new_n13196_, new_n13197_, new_n13198_,
    new_n13199_, new_n13200_, new_n13201_, new_n13202_, new_n13203_,
    new_n13204_, new_n13205_, new_n13206_, new_n13207_, new_n13208_,
    new_n13209_, new_n13210_, new_n13211_, new_n13212_, new_n13213_,
    new_n13214_, new_n13215_, new_n13216_, new_n13217_, new_n13218_,
    new_n13219_, new_n13220_, new_n13221_, new_n13222_, new_n13223_,
    new_n13224_, new_n13225_, new_n13226_, new_n13227_, new_n13228_,
    new_n13229_, new_n13230_, new_n13231_, new_n13232_, new_n13233_,
    new_n13234_, new_n13235_, new_n13236_, new_n13237_, new_n13238_,
    new_n13239_, new_n13240_, new_n13241_, new_n13242_, new_n13243_,
    new_n13244_, new_n13245_, new_n13246_, new_n13247_, new_n13248_,
    new_n13249_, new_n13250_, new_n13251_, new_n13252_, new_n13253_,
    new_n13254_, new_n13255_, new_n13256_, new_n13257_, new_n13258_,
    new_n13259_, new_n13260_, new_n13261_, new_n13262_, new_n13263_,
    new_n13264_, new_n13265_, new_n13266_, new_n13267_, new_n13268_,
    new_n13269_, new_n13270_, new_n13271_, new_n13272_, new_n13273_,
    new_n13274_, new_n13275_, new_n13276_, new_n13277_, new_n13278_,
    new_n13279_, new_n13280_, new_n13281_, new_n13282_, new_n13283_,
    new_n13284_, new_n13285_, new_n13286_, new_n13287_, new_n13288_,
    new_n13289_, new_n13290_, new_n13291_, new_n13292_, new_n13293_,
    new_n13294_, new_n13295_, new_n13296_, new_n13297_, new_n13298_,
    new_n13299_, new_n13300_, new_n13301_, new_n13302_, new_n13303_,
    new_n13304_, new_n13305_, new_n13306_, new_n13307_, new_n13308_,
    new_n13309_, new_n13310_, new_n13311_, new_n13312_, new_n13313_,
    new_n13314_, new_n13315_, new_n13316_, new_n13317_, new_n13318_,
    new_n13319_, new_n13321_, new_n13322_, new_n13323_, new_n13324_,
    new_n13325_, new_n13326_, new_n13327_, new_n13328_, new_n13329_,
    new_n13330_, new_n13331_, new_n13332_, new_n13333_, new_n13334_,
    new_n13335_, new_n13336_, new_n13337_, new_n13338_, new_n13339_,
    new_n13340_, new_n13341_, new_n13342_, new_n13343_, new_n13344_,
    new_n13345_, new_n13346_, new_n13347_, new_n13348_, new_n13349_,
    new_n13350_, new_n13351_, new_n13352_, new_n13353_, new_n13354_,
    new_n13355_, new_n13356_, new_n13357_, new_n13358_, new_n13359_,
    new_n13360_, new_n13361_, new_n13362_, new_n13363_, new_n13364_,
    new_n13365_, new_n13366_, new_n13367_, new_n13368_, new_n13369_,
    new_n13370_, new_n13371_, new_n13372_, new_n13373_, new_n13374_,
    new_n13375_, new_n13376_, new_n13377_, new_n13378_, new_n13379_,
    new_n13380_, new_n13381_, new_n13382_, new_n13383_, new_n13384_,
    new_n13385_, new_n13386_, new_n13387_, new_n13388_, new_n13389_,
    new_n13390_, new_n13391_, new_n13392_, new_n13393_, new_n13394_,
    new_n13395_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13489_, new_n13490_, new_n13491_,
    new_n13492_, new_n13493_, new_n13494_, new_n13495_, new_n13496_,
    new_n13497_, new_n13498_, new_n13499_, new_n13500_, new_n13501_,
    new_n13502_, new_n13503_, new_n13504_, new_n13505_, new_n13506_,
    new_n13507_, new_n13508_, new_n13509_, new_n13510_, new_n13511_,
    new_n13512_, new_n13513_, new_n13514_, new_n13515_, new_n13516_,
    new_n13517_, new_n13518_, new_n13519_, new_n13520_, new_n13521_,
    new_n13522_, new_n13523_, new_n13524_, new_n13525_, new_n13526_,
    new_n13527_, new_n13528_, new_n13529_, new_n13530_, new_n13531_,
    new_n13532_, new_n13533_, new_n13534_, new_n13535_, new_n13536_,
    new_n13537_, new_n13538_, new_n13539_, new_n13540_, new_n13541_,
    new_n13542_, new_n13543_, new_n13544_, new_n13545_, new_n13546_,
    new_n13547_, new_n13548_, new_n13549_, new_n13550_, new_n13551_,
    new_n13552_, new_n13553_, new_n13554_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13639_, new_n13640_, new_n13641_,
    new_n13642_, new_n13643_, new_n13644_, new_n13645_, new_n13646_,
    new_n13647_, new_n13648_, new_n13649_, new_n13650_, new_n13651_,
    new_n13652_, new_n13653_, new_n13654_, new_n13655_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13666_, new_n13667_,
    new_n13668_, new_n13669_, new_n13670_, new_n13671_, new_n13672_,
    new_n13673_, new_n13674_, new_n13675_, new_n13676_, new_n13677_,
    new_n13678_, new_n13679_, new_n13680_, new_n13681_, new_n13682_,
    new_n13683_, new_n13684_, new_n13685_, new_n13686_, new_n13687_,
    new_n13688_, new_n13689_, new_n13690_, new_n13691_, new_n13692_,
    new_n13693_, new_n13694_, new_n13695_, new_n13696_, new_n13697_,
    new_n13698_, new_n13699_, new_n13700_, new_n13701_, new_n13702_,
    new_n13703_, new_n13704_, new_n13705_, new_n13706_, new_n13707_,
    new_n13708_, new_n13709_, new_n13710_, new_n13711_, new_n13712_,
    new_n13713_, new_n13714_, new_n13715_, new_n13716_, new_n13717_,
    new_n13718_, new_n13719_, new_n13720_, new_n13721_, new_n13722_,
    new_n13723_, new_n13724_, new_n13725_, new_n13726_, new_n13727_,
    new_n13728_, new_n13729_, new_n13730_, new_n13731_, new_n13732_,
    new_n13733_, new_n13734_, new_n13735_, new_n13736_, new_n13737_,
    new_n13738_, new_n13739_, new_n13740_, new_n13741_, new_n13742_,
    new_n13743_, new_n13744_, new_n13745_, new_n13746_, new_n13747_,
    new_n13748_, new_n13749_, new_n13750_, new_n13751_, new_n13752_,
    new_n13753_, new_n13754_, new_n13755_, new_n13756_, new_n13757_,
    new_n13758_, new_n13759_, new_n13760_, new_n13761_, new_n13762_,
    new_n13763_, new_n13764_, new_n13765_, new_n13766_, new_n13767_,
    new_n13768_, new_n13769_, new_n13770_, new_n13771_, new_n13772_,
    new_n13773_, new_n13774_, new_n13775_, new_n13776_, new_n13777_,
    new_n13778_, new_n13779_, new_n13780_, new_n13781_, new_n13782_,
    new_n13783_, new_n13784_, new_n13785_, new_n13786_, new_n13787_,
    new_n13788_, new_n13789_, new_n13790_, new_n13791_, new_n13792_,
    new_n13793_, new_n13794_, new_n13795_, new_n13796_, new_n13797_,
    new_n13798_, new_n13799_, new_n13800_, new_n13801_, new_n13802_,
    new_n13803_, new_n13804_, new_n13805_, new_n13806_, new_n13807_,
    new_n13808_, new_n13809_, new_n13810_, new_n13811_, new_n13812_,
    new_n13813_, new_n13814_, new_n13815_, new_n13816_, new_n13817_,
    new_n13818_, new_n13819_, new_n13820_, new_n13821_, new_n13822_,
    new_n13824_, new_n13825_, new_n13826_, new_n13828_, new_n13829_,
    new_n13830_, new_n13831_, new_n13832_, new_n13833_, new_n13834_,
    new_n13835_, new_n13836_, new_n13837_, new_n13838_, new_n13839_,
    new_n13840_, new_n13841_, new_n13842_, new_n13843_, new_n13844_,
    new_n13845_, new_n13846_, new_n13847_, new_n13848_, new_n13849_,
    new_n13850_, new_n13851_, new_n13852_, new_n13853_, new_n13854_,
    new_n13855_, new_n13856_, new_n13857_, new_n13858_, new_n13859_,
    new_n13860_, new_n13861_, new_n13862_, new_n13863_, new_n13864_,
    new_n13865_, new_n13866_, new_n13867_, new_n13868_, new_n13869_,
    new_n13870_, new_n13871_, new_n13872_, new_n13873_, new_n13874_,
    new_n13875_, new_n13876_, new_n13877_, new_n13878_, new_n13879_,
    new_n13880_, new_n13881_, new_n13882_, new_n13883_, new_n13884_,
    new_n13885_, new_n13886_, new_n13887_, new_n13888_, new_n13889_,
    new_n13890_, new_n13891_, new_n13892_, new_n13893_, new_n13894_,
    new_n13895_, new_n13896_, new_n13897_, new_n13898_, new_n13899_,
    new_n13900_, new_n13901_, new_n13902_, new_n13903_, new_n13904_,
    new_n13905_, new_n13906_, new_n13907_, new_n13908_, new_n13909_,
    new_n13910_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13917_, new_n13918_, new_n13919_, new_n13920_,
    new_n13921_, new_n13922_, new_n13923_, new_n13924_, new_n13925_,
    new_n13926_, new_n13927_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13933_, new_n13934_, new_n13935_,
    new_n13936_, new_n13937_, new_n13938_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13944_, new_n13945_,
    new_n13946_, new_n13947_, new_n13948_, new_n13949_, new_n13950_,
    new_n13951_, new_n13952_, new_n13953_, new_n13954_, new_n13955_,
    new_n13956_, new_n13957_, new_n13958_, new_n13959_, new_n13960_,
    new_n13961_, new_n13962_, new_n13963_, new_n13964_, new_n13965_,
    new_n13966_, new_n13967_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14013_, new_n14014_, new_n14015_,
    new_n14016_, new_n14017_, new_n14018_, new_n14019_, new_n14020_,
    new_n14021_, new_n14022_, new_n14023_, new_n14024_, new_n14025_,
    new_n14026_, new_n14027_, new_n14028_, new_n14029_, new_n14030_,
    new_n14031_, new_n14032_, new_n14033_, new_n14034_, new_n14035_,
    new_n14036_, new_n14037_, new_n14038_, new_n14039_, new_n14040_,
    new_n14041_, new_n14042_, new_n14043_, new_n14044_, new_n14045_,
    new_n14046_, new_n14047_, new_n14048_, new_n14049_, new_n14050_,
    new_n14051_, new_n14052_, new_n14053_, new_n14054_, new_n14055_,
    new_n14056_, new_n14057_, new_n14058_, new_n14059_, new_n14060_,
    new_n14061_, new_n14062_, new_n14063_, new_n14064_, new_n14065_,
    new_n14066_, new_n14067_, new_n14068_, new_n14069_, new_n14070_,
    new_n14071_, new_n14072_, new_n14073_, new_n14074_, new_n14075_,
    new_n14076_, new_n14077_, new_n14078_, new_n14079_, new_n14080_,
    new_n14081_, new_n14082_, new_n14086_, new_n14087_, new_n14088_,
    new_n14089_, new_n14090_, new_n14091_, new_n14092_, new_n14093_,
    new_n14094_, new_n14095_, new_n14096_, new_n14097_, new_n14098_,
    new_n14099_, new_n14100_, new_n14101_, new_n14102_, new_n14103_,
    new_n14104_, new_n14105_, new_n14106_, new_n14107_, new_n14108_,
    new_n14109_, new_n14110_, new_n14111_, new_n14112_, new_n14113_,
    new_n14114_, new_n14115_, new_n14116_, new_n14117_, new_n14118_,
    new_n14119_, new_n14120_, new_n14121_, new_n14122_, new_n14123_,
    new_n14124_, new_n14125_, new_n14127_, new_n14128_, new_n14129_,
    new_n14130_, new_n14131_, new_n14132_, new_n14133_, new_n14134_,
    new_n14135_, new_n14136_, new_n14137_, new_n14138_, new_n14139_,
    new_n14140_, new_n14141_, new_n14142_, new_n14143_, new_n14144_,
    new_n14145_, new_n14146_, new_n14147_, new_n14148_, new_n14149_,
    new_n14150_, new_n14151_, new_n14152_, new_n14153_, new_n14154_,
    new_n14155_, new_n14156_, new_n14157_, new_n14158_, new_n14159_,
    new_n14160_, new_n14161_, new_n14162_, new_n14163_, new_n14164_,
    new_n14165_, new_n14166_, new_n14167_, new_n14168_, new_n14169_,
    new_n14170_, new_n14171_, new_n14172_, new_n14173_, new_n14174_,
    new_n14175_, new_n14176_, new_n14177_, new_n14178_, new_n14179_,
    new_n14180_, new_n14181_, new_n14182_, new_n14183_, new_n14184_,
    new_n14185_, new_n14186_, new_n14187_, new_n14188_, new_n14189_,
    new_n14190_, new_n14191_, new_n14192_, new_n14193_, new_n14194_,
    new_n14195_, new_n14196_, new_n14197_, new_n14198_, new_n14199_,
    new_n14200_, new_n14201_, new_n14202_, new_n14203_, new_n14204_,
    new_n14205_, new_n14206_, new_n14207_, new_n14208_, new_n14209_,
    new_n14210_, new_n14211_, new_n14212_, new_n14213_, new_n14214_,
    new_n14215_, new_n14216_, new_n14217_, new_n14218_, new_n14219_,
    new_n14220_, new_n14221_, new_n14222_, new_n14223_, new_n14224_,
    new_n14225_, new_n14226_, new_n14227_, new_n14228_, new_n14229_,
    new_n14230_, new_n14231_, new_n14232_, new_n14233_, new_n14234_,
    new_n14235_, new_n14236_, new_n14237_, new_n14238_, new_n14239_,
    new_n14240_, new_n14241_, new_n14242_, new_n14243_, new_n14244_,
    new_n14245_, new_n14246_, new_n14247_, new_n14248_, new_n14249_,
    new_n14250_, new_n14251_, new_n14252_, new_n14253_, new_n14254_,
    new_n14255_, new_n14256_, new_n14257_, new_n14258_, new_n14259_,
    new_n14260_, new_n14261_, new_n14262_, new_n14263_, new_n14264_,
    new_n14265_, new_n14266_, new_n14267_, new_n14268_, new_n14269_,
    new_n14270_, new_n14271_, new_n14272_, new_n14273_, new_n14274_,
    new_n14276_, new_n14277_, new_n14278_, new_n14279_, new_n14280_,
    new_n14281_, new_n14282_, new_n14283_, new_n14284_, new_n14285_,
    new_n14286_, new_n14287_, new_n14288_, new_n14289_, new_n14290_,
    new_n14291_, new_n14292_, new_n14293_, new_n14294_, new_n14295_,
    new_n14296_, new_n14297_, new_n14298_, new_n14299_, new_n14300_,
    new_n14301_, new_n14302_, new_n14303_, new_n14304_, new_n14305_,
    new_n14306_, new_n14307_, new_n14308_, new_n14309_, new_n14310_,
    new_n14311_, new_n14312_, new_n14313_, new_n14314_, new_n14315_,
    new_n14316_, new_n14317_, new_n14318_, new_n14319_, new_n14320_,
    new_n14321_, new_n14322_, new_n14323_, new_n14324_, new_n14325_,
    new_n14326_, new_n14327_, new_n14328_, new_n14329_, new_n14330_,
    new_n14331_, new_n14332_, new_n14333_, new_n14334_, new_n14335_,
    new_n14336_, new_n14337_, new_n14338_, new_n14339_, new_n14340_,
    new_n14341_, new_n14342_, new_n14343_, new_n14344_, new_n14345_,
    new_n14346_, new_n14347_, new_n14348_, new_n14349_, new_n14350_,
    new_n14351_, new_n14352_, new_n14353_, new_n14354_, new_n14355_,
    new_n14356_, new_n14357_, new_n14358_, new_n14359_, new_n14360_,
    new_n14361_, new_n14362_, new_n14363_, new_n14364_, new_n14365_,
    new_n14366_, new_n14367_, new_n14368_, new_n14369_, new_n14370_,
    new_n14371_, new_n14372_, new_n14373_, new_n14374_, new_n14375_,
    new_n14376_, new_n14377_, new_n14378_, new_n14379_, new_n14380_,
    new_n14381_, new_n14382_, new_n14383_, new_n14384_, new_n14385_,
    new_n14386_, new_n14387_, new_n14388_, new_n14389_, new_n14390_,
    new_n14391_, new_n14392_, new_n14393_, new_n14394_, new_n14395_,
    new_n14396_, new_n14397_, new_n14398_, new_n14399_, new_n14400_,
    new_n14401_, new_n14402_, new_n14403_, new_n14404_, new_n14405_,
    new_n14406_, new_n14407_, new_n14408_, new_n14409_, new_n14410_,
    new_n14411_, new_n14412_, new_n14413_, new_n14414_, new_n14415_,
    new_n14417_, new_n14418_, new_n14419_, new_n14420_, new_n14421_,
    new_n14422_, new_n14423_, new_n14424_, new_n14425_, new_n14426_,
    new_n14427_, new_n14428_, new_n14429_, new_n14430_, new_n14431_,
    new_n14432_, new_n14433_, new_n14434_, new_n14435_, new_n14436_,
    new_n14437_, new_n14438_, new_n14439_, new_n14440_, new_n14441_,
    new_n14442_, new_n14443_, new_n14444_, new_n14445_, new_n14446_,
    new_n14447_, new_n14448_, new_n14449_, new_n14450_, new_n14451_,
    new_n14452_, new_n14453_, new_n14454_, new_n14455_, new_n14456_,
    new_n14457_, new_n14458_, new_n14459_, new_n14460_, new_n14461_,
    new_n14462_, new_n14463_, new_n14464_, new_n14465_, new_n14466_,
    new_n14467_, new_n14468_, new_n14469_, new_n14470_, new_n14471_,
    new_n14472_, new_n14473_, new_n14474_, new_n14475_, new_n14476_,
    new_n14477_, new_n14478_, new_n14479_, new_n14480_, new_n14481_,
    new_n14482_, new_n14483_, new_n14484_, new_n14485_, new_n14486_,
    new_n14487_, new_n14488_, new_n14489_, new_n14490_, new_n14491_,
    new_n14492_, new_n14493_, new_n14494_, new_n14495_, new_n14496_,
    new_n14497_, new_n14498_, new_n14499_, new_n14500_, new_n14501_,
    new_n14502_, new_n14503_, new_n14504_, new_n14505_, new_n14506_,
    new_n14507_, new_n14508_, new_n14509_, new_n14510_, new_n14511_,
    new_n14512_, new_n14513_, new_n14514_, new_n14515_, new_n14516_,
    new_n14517_, new_n14518_, new_n14519_, new_n14520_, new_n14521_,
    new_n14522_, new_n14523_, new_n14524_, new_n14525_, new_n14526_,
    new_n14527_, new_n14528_, new_n14529_, new_n14530_, new_n14531_,
    new_n14532_, new_n14533_, new_n14534_, new_n14535_, new_n14536_,
    new_n14537_, new_n14538_, new_n14539_, new_n14540_, new_n14541_,
    new_n14542_, new_n14543_, new_n14544_, new_n14545_, new_n14546_,
    new_n14547_, new_n14548_, new_n14549_, new_n14550_, new_n14551_,
    new_n14552_, new_n14553_, new_n14554_, new_n14555_, new_n14556_,
    new_n14557_, new_n14558_, new_n14559_, new_n14560_, new_n14561_,
    new_n14562_, new_n14563_, new_n14564_, new_n14565_, new_n14566_,
    new_n14567_, new_n14568_, new_n14569_, new_n14570_, new_n14571_,
    new_n14572_, new_n14573_, new_n14574_, new_n14575_, new_n14576_,
    new_n14577_, new_n14578_, new_n14579_, new_n14580_, new_n14582_,
    new_n14583_, new_n14584_, new_n14585_, new_n14586_, new_n14587_,
    new_n14588_, new_n14589_, new_n14590_, new_n14591_, new_n14592_,
    new_n14593_, new_n14594_, new_n14595_, new_n14596_, new_n14597_,
    new_n14598_, new_n14599_, new_n14600_, new_n14601_, new_n14602_,
    new_n14603_, new_n14604_, new_n14605_, new_n14606_, new_n14607_,
    new_n14608_, new_n14609_, new_n14610_, new_n14611_, new_n14612_,
    new_n14613_, new_n14614_, new_n14615_, new_n14616_, new_n14617_,
    new_n14618_, new_n14619_, new_n14620_, new_n14621_, new_n14622_,
    new_n14623_, new_n14624_, new_n14625_, new_n14626_, new_n14627_,
    new_n14628_, new_n14629_, new_n14630_, new_n14631_, new_n14632_,
    new_n14633_, new_n14634_, new_n14635_, new_n14636_, new_n14637_,
    new_n14638_, new_n14639_, new_n14640_, new_n14641_, new_n14642_,
    new_n14643_, new_n14644_, new_n14645_, new_n14646_, new_n14647_,
    new_n14648_, new_n14649_, new_n14650_, new_n14651_, new_n14652_,
    new_n14653_, new_n14654_, new_n14655_, new_n14656_, new_n14657_,
    new_n14658_, new_n14659_, new_n14660_, new_n14661_, new_n14662_,
    new_n14663_, new_n14664_, new_n14665_, new_n14666_, new_n14667_,
    new_n14668_, new_n14669_, new_n14670_, new_n14671_, new_n14672_,
    new_n14673_, new_n14674_, new_n14675_, new_n14676_, new_n14677_,
    new_n14678_, new_n14679_, new_n14680_, new_n14681_, new_n14682_,
    new_n14683_, new_n14684_, new_n14685_, new_n14686_, new_n14687_,
    new_n14688_, new_n14689_, new_n14690_, new_n14691_, new_n14692_,
    new_n14693_, new_n14694_, new_n14695_, new_n14696_, new_n14697_,
    new_n14698_, new_n14699_, new_n14700_, new_n14701_, new_n14702_,
    new_n14703_, new_n14704_, new_n14705_, new_n14706_, new_n14707_,
    new_n14708_, new_n14709_, new_n14710_, new_n14711_, new_n14713_,
    new_n14714_, new_n14716_, new_n14717_, new_n14718_, new_n14719_,
    new_n14720_, new_n14721_, new_n14722_, new_n14723_, new_n14724_,
    new_n14725_, new_n14726_, new_n14727_, new_n14728_, new_n14730_,
    new_n14731_, new_n14732_, new_n14733_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14739_, new_n14740_,
    new_n14741_, new_n14742_, new_n14743_, new_n14744_, new_n14745_,
    new_n14746_, new_n14747_, new_n14748_, new_n14749_, new_n14750_,
    new_n14751_, new_n14752_, new_n14753_, new_n14754_, new_n14755_,
    new_n14756_, new_n14757_, new_n14758_, new_n14759_, new_n14760_,
    new_n14761_, new_n14762_, new_n14763_, new_n14764_, new_n14765_,
    new_n14766_, new_n14767_, new_n14768_, new_n14769_, new_n14770_,
    new_n14771_, new_n14772_, new_n14773_, new_n14774_, new_n14775_,
    new_n14776_, new_n14777_, new_n14778_, new_n14779_, new_n14780_,
    new_n14781_, new_n14782_, new_n14783_, new_n14784_, new_n14785_,
    new_n14786_, new_n14787_, new_n14788_, new_n14789_, new_n14790_,
    new_n14791_, new_n14792_, new_n14793_, new_n14794_, new_n14795_,
    new_n14796_, new_n14797_, new_n14798_, new_n14799_, new_n14800_,
    new_n14801_, new_n14802_, new_n14803_, new_n14804_, new_n14805_,
    new_n14806_, new_n14807_, new_n14808_, new_n14809_, new_n14810_,
    new_n14811_, new_n14812_, new_n14813_, new_n14814_, new_n14815_,
    new_n14816_, new_n14817_, new_n14818_, new_n14819_, new_n14820_,
    new_n14821_, new_n14822_, new_n14823_, new_n14824_, new_n14825_,
    new_n14826_, new_n14827_, new_n14828_, new_n14829_, new_n14830_,
    new_n14831_, new_n14832_, new_n14833_, new_n14834_, new_n14835_,
    new_n14836_, new_n14837_, new_n14838_, new_n14839_, new_n14840_,
    new_n14841_, new_n14842_, new_n14843_, new_n14844_, new_n14845_,
    new_n14846_, new_n14847_, new_n14848_, new_n14849_, new_n14850_,
    new_n14851_, new_n14852_, new_n14853_, new_n14854_, new_n14855_,
    new_n14856_, new_n14857_, new_n14858_, new_n14859_, new_n14860_,
    new_n14861_, new_n14862_, new_n14863_, new_n14864_, new_n14865_,
    new_n14866_, new_n14867_, new_n14868_, new_n14869_, new_n14870_,
    new_n14871_, new_n14872_, new_n14873_, new_n14874_, new_n14875_,
    new_n14876_, new_n14877_, new_n14878_, new_n14879_, new_n14880_,
    new_n14881_, new_n14882_, new_n14883_, new_n14884_, new_n14885_,
    new_n14886_, new_n14887_, new_n14888_, new_n14889_, new_n14890_,
    new_n14891_, new_n14892_, new_n14893_, new_n14894_, new_n14895_,
    new_n14896_, new_n14897_, new_n14898_, new_n14899_, new_n14900_,
    new_n14901_, new_n14902_, new_n14903_, new_n14904_, new_n14905_,
    new_n14906_, new_n14907_, new_n14908_, new_n14909_, new_n14910_,
    new_n14911_, new_n14912_, new_n14913_, new_n14914_, new_n14915_,
    new_n14916_, new_n14917_, new_n14918_, new_n14919_, new_n14920_,
    new_n14921_, new_n14922_, new_n14923_, new_n14924_, new_n14925_,
    new_n14926_, new_n14927_, new_n14928_, new_n14929_, new_n14930_,
    new_n14931_, new_n14932_, new_n14933_, new_n14934_, new_n14935_,
    new_n14936_, new_n14937_, new_n14938_, new_n14939_, new_n14940_,
    new_n14941_, new_n14942_, new_n14943_, new_n14944_, new_n14945_,
    new_n14946_, new_n14947_, new_n14948_, new_n14949_, new_n14950_,
    new_n14951_, new_n14952_, new_n14953_, new_n14954_, new_n14955_,
    new_n14956_, new_n14957_, new_n14958_, new_n14959_, new_n14960_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14981_, new_n14983_, new_n14984_, new_n14985_, new_n14986_,
    new_n14987_, new_n14988_, new_n14989_, new_n14990_, new_n14991_,
    new_n14992_, new_n14993_, new_n14994_, new_n14995_, new_n14996_,
    new_n14997_, new_n14998_, new_n14999_, new_n15000_, new_n15001_,
    new_n15002_, new_n15003_, new_n15004_, new_n15005_, new_n15006_,
    new_n15007_, new_n15008_, new_n15009_, new_n15010_, new_n15011_,
    new_n15012_, new_n15013_, new_n15014_, new_n15015_, new_n15016_,
    new_n15017_, new_n15018_, new_n15019_, new_n15020_, new_n15021_,
    new_n15022_, new_n15023_, new_n15024_, new_n15025_, new_n15026_,
    new_n15027_, new_n15028_, new_n15029_, new_n15030_, new_n15031_,
    new_n15032_, new_n15033_, new_n15034_, new_n15035_, new_n15036_,
    new_n15037_, new_n15038_, new_n15039_, new_n15040_, new_n15041_,
    new_n15042_, new_n15043_, new_n15044_, new_n15045_, new_n15046_,
    new_n15047_, new_n15048_, new_n15049_, new_n15050_, new_n15051_,
    new_n15052_, new_n15053_, new_n15054_, new_n15055_, new_n15056_,
    new_n15057_, new_n15058_, new_n15059_, new_n15060_, new_n15061_,
    new_n15062_, new_n15063_, new_n15064_, new_n15065_, new_n15066_,
    new_n15067_, new_n15068_, new_n15069_, new_n15070_, new_n15071_,
    new_n15072_, new_n15073_, new_n15074_, new_n15075_, new_n15076_,
    new_n15077_, new_n15078_, new_n15079_, new_n15080_, new_n15081_,
    new_n15082_, new_n15083_, new_n15084_, new_n15085_, new_n15086_,
    new_n15087_, new_n15088_, new_n15089_, new_n15090_, new_n15091_,
    new_n15092_, new_n15093_, new_n15094_, new_n15095_, new_n15096_,
    new_n15097_, new_n15098_, new_n15099_, new_n15100_, new_n15101_,
    new_n15102_, new_n15103_, new_n15104_, new_n15105_, new_n15106_,
    new_n15108_, new_n15109_, new_n15110_, new_n15111_, new_n15112_,
    new_n15113_, new_n15114_, new_n15115_, new_n15116_, new_n15117_,
    new_n15118_, new_n15119_, new_n15120_, new_n15121_, new_n15122_,
    new_n15123_, new_n15124_, new_n15125_, new_n15126_, new_n15127_,
    new_n15128_, new_n15129_, new_n15130_, new_n15131_, new_n15132_,
    new_n15133_, new_n15134_, new_n15135_, new_n15136_, new_n15137_,
    new_n15138_, new_n15139_, new_n15140_, new_n15141_, new_n15142_,
    new_n15143_, new_n15144_, new_n15145_, new_n15146_, new_n15147_,
    new_n15148_, new_n15149_, new_n15150_, new_n15152_, new_n15153_,
    new_n15154_, new_n15155_, new_n15156_, new_n15157_, new_n15158_,
    new_n15159_, new_n15160_, new_n15161_, new_n15162_, new_n15163_,
    new_n15164_, new_n15165_, new_n15166_, new_n15167_, new_n15168_,
    new_n15169_, new_n15170_, new_n15171_, new_n15172_, new_n15173_,
    new_n15174_, new_n15175_, new_n15176_, new_n15177_, new_n15178_,
    new_n15179_, new_n15180_, new_n15181_, new_n15182_, new_n15183_,
    new_n15184_, new_n15185_, new_n15186_, new_n15187_, new_n15188_,
    new_n15189_, new_n15190_, new_n15191_, new_n15192_, new_n15193_,
    new_n15194_, new_n15195_, new_n15196_, new_n15197_, new_n15198_,
    new_n15199_, new_n15200_, new_n15201_, new_n15202_, new_n15203_,
    new_n15204_, new_n15205_, new_n15206_, new_n15207_, new_n15208_,
    new_n15209_, new_n15210_, new_n15211_, new_n15212_, new_n15213_,
    new_n15214_, new_n15215_, new_n15216_, new_n15217_, new_n15218_,
    new_n15219_, new_n15220_, new_n15221_, new_n15222_, new_n15223_,
    new_n15224_, new_n15225_, new_n15226_, new_n15227_, new_n15228_,
    new_n15229_, new_n15230_, new_n15231_, new_n15233_, new_n15234_,
    new_n15235_, new_n15236_, new_n15237_, new_n15238_, new_n15239_,
    new_n15240_, new_n15241_, new_n15242_, new_n15243_, new_n15244_,
    new_n15245_, new_n15246_, new_n15247_, new_n15248_, new_n15249_,
    new_n15250_, new_n15251_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15267_, new_n15268_, new_n15269_,
    new_n15270_, new_n15271_, new_n15272_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15300_, new_n15301_, new_n15302_, new_n15303_, new_n15304_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15335_, new_n15336_, new_n15337_, new_n15338_, new_n15339_,
    new_n15340_, new_n15341_, new_n15342_, new_n15343_, new_n15344_,
    new_n15345_, new_n15346_, new_n15347_, new_n15348_, new_n15349_,
    new_n15350_, new_n15351_, new_n15352_, new_n15353_, new_n15354_,
    new_n15355_, new_n15356_, new_n15357_, new_n15358_, new_n15359_,
    new_n15360_, new_n15361_, new_n15362_, new_n15363_, new_n15364_,
    new_n15365_, new_n15366_, new_n15367_, new_n15368_, new_n15370_,
    new_n15371_, new_n15372_, new_n15373_, new_n15374_, new_n15375_,
    new_n15376_, new_n15377_, new_n15378_, new_n15379_, new_n15380_,
    new_n15381_, new_n15382_, new_n15383_, new_n15384_, new_n15385_,
    new_n15386_, new_n15387_, new_n15388_, new_n15389_, new_n15390_,
    new_n15391_, new_n15392_, new_n15393_, new_n15394_, new_n15395_,
    new_n15396_, new_n15397_, new_n15398_, new_n15399_, new_n15400_,
    new_n15401_, new_n15402_, new_n15403_, new_n15404_, new_n15405_,
    new_n15406_, new_n15407_, new_n15408_, new_n15409_, new_n15410_,
    new_n15411_, new_n15412_, new_n15413_, new_n15414_, new_n15415_,
    new_n15416_, new_n15417_, new_n15418_, new_n15419_, new_n15420_,
    new_n15421_, new_n15422_, new_n15423_, new_n15424_, new_n15425_,
    new_n15426_, new_n15427_, new_n15428_, new_n15429_, new_n15430_,
    new_n15431_, new_n15432_, new_n15433_, new_n15434_, new_n15435_,
    new_n15436_, new_n15437_, new_n15439_, new_n15440_, new_n15441_,
    new_n15442_, new_n15443_, new_n15444_, new_n15445_, new_n15446_,
    new_n15447_, new_n15448_, new_n15449_, new_n15450_, new_n15451_,
    new_n15452_, new_n15453_, new_n15454_, new_n15455_, new_n15456_,
    new_n15457_, new_n15458_, new_n15459_, new_n15460_, new_n15461_,
    new_n15462_, new_n15463_, new_n15464_, new_n15465_, new_n15466_,
    new_n15467_, new_n15468_, new_n15469_, new_n15471_, new_n15472_,
    new_n15473_, new_n15474_, new_n15475_, new_n15476_, new_n15477_,
    new_n15478_, new_n15479_, new_n15480_, new_n15481_, new_n15482_,
    new_n15483_, new_n15484_, new_n15485_, new_n15486_, new_n15487_,
    new_n15488_, new_n15489_, new_n15490_, new_n15491_, new_n15492_,
    new_n15493_, new_n15494_, new_n15495_, new_n15496_, new_n15497_,
    new_n15498_, new_n15499_, new_n15500_, new_n15501_, new_n15502_,
    new_n15503_, new_n15504_, new_n15505_, new_n15506_, new_n15507_,
    new_n15508_, new_n15509_, new_n15510_, new_n15511_, new_n15512_,
    new_n15513_, new_n15514_, new_n15515_, new_n15516_, new_n15517_,
    new_n15518_, new_n15519_, new_n15520_, new_n15521_, new_n15522_,
    new_n15523_, new_n15524_, new_n15525_, new_n15526_, new_n15527_,
    new_n15528_, new_n15529_, new_n15530_, new_n15531_, new_n15532_,
    new_n15533_, new_n15534_, new_n15535_, new_n15536_, new_n15537_,
    new_n15538_, new_n15539_, new_n15540_, new_n15541_, new_n15542_,
    new_n15543_, new_n15544_, new_n15545_, new_n15546_, new_n15547_,
    new_n15548_, new_n15549_, new_n15550_, new_n15551_, new_n15552_,
    new_n15553_, new_n15554_, new_n15555_, new_n15556_, new_n15557_,
    new_n15558_, new_n15559_, new_n15560_, new_n15561_, new_n15562_,
    new_n15563_, new_n15564_, new_n15565_, new_n15566_, new_n15567_,
    new_n15568_, new_n15569_, new_n15570_, new_n15571_, new_n15572_,
    new_n15573_, new_n15574_, new_n15575_, new_n15576_, new_n15577_,
    new_n15578_, new_n15579_, new_n15580_, new_n15581_, new_n15582_,
    new_n15583_, new_n15584_, new_n15585_, new_n15586_, new_n15587_,
    new_n15588_, new_n15589_, new_n15591_, new_n15592_, new_n15593_,
    new_n15594_, new_n15595_, new_n15596_, new_n15597_, new_n15598_,
    new_n15599_, new_n15600_, new_n15601_, new_n15602_, new_n15603_,
    new_n15604_, new_n15605_, new_n15606_, new_n15607_, new_n15608_,
    new_n15609_, new_n15610_, new_n15611_, new_n15612_, new_n15613_,
    new_n15614_, new_n15615_, new_n15616_, new_n15617_, new_n15618_,
    new_n15619_, new_n15620_, new_n15621_, new_n15622_, new_n15623_,
    new_n15624_, new_n15625_, new_n15626_, new_n15627_, new_n15628_,
    new_n15629_, new_n15630_, new_n15631_, new_n15632_, new_n15633_,
    new_n15634_, new_n15635_, new_n15636_, new_n15637_, new_n15638_,
    new_n15639_, new_n15640_, new_n15641_, new_n15642_, new_n15643_,
    new_n15644_, new_n15645_, new_n15646_, new_n15647_, new_n15648_,
    new_n15649_, new_n15650_, new_n15651_, new_n15652_, new_n15653_,
    new_n15654_, new_n15655_, new_n15656_, new_n15657_, new_n15658_,
    new_n15659_, new_n15660_, new_n15661_, new_n15662_, new_n15663_,
    new_n15664_, new_n15665_, new_n15666_, new_n15667_, new_n15668_,
    new_n15669_, new_n15670_, new_n15671_, new_n15672_, new_n15673_,
    new_n15674_, new_n15675_, new_n15676_, new_n15677_, new_n15678_,
    new_n15679_, new_n15680_, new_n15681_, new_n15682_, new_n15683_,
    new_n15684_, new_n15685_, new_n15686_, new_n15687_, new_n15688_,
    new_n15689_, new_n15690_, new_n15691_, new_n15692_, new_n15693_,
    new_n15694_, new_n15695_, new_n15696_, new_n15697_, new_n15698_,
    new_n15699_, new_n15700_, new_n15701_, new_n15702_, new_n15703_,
    new_n15704_, new_n15705_, new_n15706_, new_n15707_, new_n15708_,
    new_n15710_, new_n15711_, new_n15712_, new_n15713_, new_n15714_,
    new_n15715_, new_n15716_, new_n15717_, new_n15718_, new_n15719_,
    new_n15720_, new_n15721_, new_n15722_, new_n15723_, new_n15724_,
    new_n15725_, new_n15726_, new_n15727_, new_n15728_, new_n15729_,
    new_n15730_, new_n15731_, new_n15732_, new_n15733_, new_n15734_,
    new_n15735_, new_n15736_, new_n15737_, new_n15738_, new_n15739_,
    new_n15740_, new_n15741_, new_n15742_, new_n15743_, new_n15744_,
    new_n15745_, new_n15746_, new_n15747_, new_n15748_, new_n15749_,
    new_n15750_, new_n15751_, new_n15752_, new_n15753_, new_n15754_,
    new_n15755_, new_n15756_, new_n15757_, new_n15758_, new_n15759_,
    new_n15760_, new_n15761_, new_n15762_, new_n15763_, new_n15764_,
    new_n15765_, new_n15766_, new_n15767_, new_n15768_, new_n15769_,
    new_n15770_, new_n15771_, new_n15772_, new_n15773_, new_n15774_,
    new_n15775_, new_n15776_, new_n15777_, new_n15778_, new_n15779_,
    new_n15780_, new_n15781_, new_n15782_, new_n15783_, new_n15784_,
    new_n15785_, new_n15786_, new_n15787_, new_n15788_, new_n15789_,
    new_n15790_, new_n15791_, new_n15792_, new_n15793_, new_n15794_,
    new_n15795_, new_n15796_, new_n15797_, new_n15798_, new_n15799_,
    new_n15800_, new_n15801_, new_n15802_, new_n15803_, new_n15804_,
    new_n15805_, new_n15806_, new_n15807_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15840_,
    new_n15841_, new_n15842_, new_n15843_, new_n15844_, new_n15845_,
    new_n15846_, new_n15847_, new_n15848_, new_n15849_, new_n15850_,
    new_n15851_, new_n15852_, new_n15853_, new_n15857_, new_n15859_,
    new_n15863_, new_n15864_, new_n15865_, new_n15866_, new_n15867_,
    new_n15868_, new_n15869_, new_n15870_, new_n15871_, new_n15872_,
    new_n15873_, new_n15874_, new_n15875_, new_n15876_, new_n15877_,
    new_n15878_, new_n15879_, new_n15880_, new_n15881_, new_n15882_,
    new_n15883_, new_n15884_, new_n15885_, new_n15886_, new_n15887_,
    new_n15888_, new_n15889_, new_n15890_, new_n15891_, new_n15892_,
    new_n15893_, new_n15894_, new_n15895_, new_n15896_, new_n15897_,
    new_n15898_, new_n15899_, new_n15900_, new_n15901_, new_n15902_,
    new_n15903_, new_n15904_, new_n15905_, new_n15906_, new_n15907_,
    new_n15908_, new_n15909_, new_n15911_, new_n15912_, new_n15913_,
    new_n15914_, new_n15915_, new_n15916_, new_n15917_, new_n15918_,
    new_n15919_, new_n15920_, new_n15921_, new_n15922_, new_n15923_,
    new_n15924_, new_n15925_, new_n15926_, new_n15927_, new_n15928_,
    new_n15929_, new_n15930_, new_n15931_, new_n15932_, new_n15933_,
    new_n15934_, new_n15935_, new_n15936_, new_n15937_, new_n15938_,
    new_n15939_, new_n15940_, new_n15941_, new_n15942_, new_n15943_,
    new_n15944_, new_n15945_, new_n15946_, new_n15947_, new_n15948_,
    new_n15949_, new_n15950_, new_n15951_, new_n15952_, new_n15953_,
    new_n15954_, new_n15955_, new_n15956_, new_n15957_, new_n15958_,
    new_n15959_, new_n15960_, new_n15961_, new_n15962_, new_n15963_,
    new_n15964_, new_n15965_, new_n15966_, new_n15967_, new_n15968_,
    new_n15969_, new_n15970_, new_n15971_, new_n15972_, new_n15973_,
    new_n15974_, new_n15975_, new_n15976_, new_n15977_, new_n15978_,
    new_n15979_, new_n15980_, new_n15981_, new_n15982_, new_n15986_,
    new_n15987_, new_n15988_, new_n15989_, new_n15990_, new_n15991_,
    new_n15992_, new_n15993_, new_n15994_, new_n15995_, new_n15996_,
    new_n15997_, new_n15998_, new_n15999_, new_n16000_, new_n16001_,
    new_n16002_, new_n16003_, new_n16004_, new_n16005_, new_n16006_,
    new_n16007_, new_n16008_, new_n16009_, new_n16010_, new_n16012_,
    new_n16013_, new_n16014_, new_n16015_, new_n16016_, new_n16017_,
    new_n16018_, new_n16019_, new_n16020_, new_n16021_, new_n16022_,
    new_n16023_, new_n16024_, new_n16025_, new_n16026_, new_n16027_,
    new_n16028_, new_n16029_, new_n16030_, new_n16031_, new_n16032_,
    new_n16033_, new_n16034_, new_n16035_, new_n16036_, new_n16037_,
    new_n16038_, new_n16039_, new_n16040_, new_n16041_, new_n16042_,
    new_n16043_, new_n16044_, new_n16045_, new_n16046_, new_n16047_,
    new_n16048_, new_n16049_, new_n16050_, new_n16051_, new_n16052_,
    new_n16053_, new_n16054_, new_n16055_, new_n16056_, new_n16057_,
    new_n16058_, new_n16059_, new_n16060_, new_n16061_, new_n16062_,
    new_n16063_, new_n16064_, new_n16065_, new_n16066_, new_n16067_,
    new_n16068_, new_n16069_, new_n16070_, new_n16071_, new_n16072_,
    new_n16073_, new_n16074_, new_n16075_, new_n16076_, new_n16077_,
    new_n16078_, new_n16079_, new_n16080_, new_n16081_, new_n16082_,
    new_n16083_, new_n16084_, new_n16085_, new_n16086_, new_n16087_,
    new_n16088_, new_n16089_, new_n16090_, new_n16091_, new_n16092_,
    new_n16093_, new_n16094_, new_n16095_, new_n16096_, new_n16097_,
    new_n16098_, new_n16099_, new_n16101_, new_n16102_, new_n16103_,
    new_n16104_, new_n16105_, new_n16106_, new_n16107_, new_n16108_,
    new_n16109_, new_n16110_, new_n16111_, new_n16112_, new_n16113_,
    new_n16114_, new_n16115_, new_n16116_, new_n16117_, new_n16118_,
    new_n16119_, new_n16120_, new_n16121_, new_n16122_, new_n16123_,
    new_n16124_, new_n16125_, new_n16126_, new_n16127_, new_n16128_,
    new_n16129_, new_n16130_, new_n16131_, new_n16132_, new_n16133_,
    new_n16134_, new_n16135_, new_n16136_, new_n16137_, new_n16138_,
    new_n16139_, new_n16140_, new_n16141_, new_n16142_, new_n16143_,
    new_n16144_, new_n16145_, new_n16146_, new_n16147_, new_n16148_,
    new_n16149_, new_n16150_, new_n16151_, new_n16152_, new_n16153_,
    new_n16154_, new_n16155_, new_n16156_, new_n16157_, new_n16158_,
    new_n16159_, new_n16160_, new_n16161_, new_n16162_, new_n16163_,
    new_n16164_, new_n16165_, new_n16166_, new_n16167_, new_n16168_,
    new_n16169_, new_n16170_, new_n16171_, new_n16172_, new_n16173_,
    new_n16174_, new_n16175_, new_n16177_, new_n16178_, new_n16179_,
    new_n16180_, new_n16181_, new_n16182_, new_n16183_, new_n16184_,
    new_n16185_, new_n16186_, new_n16187_, new_n16188_, new_n16189_,
    new_n16190_, new_n16191_, new_n16192_, new_n16193_, new_n16194_,
    new_n16195_, new_n16196_, new_n16197_, new_n16198_, new_n16199_,
    new_n16200_, new_n16201_, new_n16202_, new_n16203_, new_n16204_,
    new_n16205_, new_n16206_, new_n16207_, new_n16208_, new_n16209_,
    new_n16210_, new_n16211_, new_n16212_, new_n16213_, new_n16214_,
    new_n16215_, new_n16216_, new_n16217_, new_n16218_, new_n16219_,
    new_n16220_, new_n16221_, new_n16222_, new_n16223_, new_n16224_,
    new_n16225_, new_n16226_, new_n16227_, new_n16228_, new_n16229_,
    new_n16230_, new_n16231_, new_n16232_, new_n16233_, new_n16234_,
    new_n16235_, new_n16236_, new_n16237_, new_n16238_, new_n16239_,
    new_n16240_, new_n16241_, new_n16242_, new_n16243_, new_n16244_,
    new_n16245_, new_n16246_, new_n16247_, new_n16248_, new_n16249_,
    new_n16250_, new_n16251_, new_n16252_, new_n16253_, new_n16254_,
    new_n16255_, new_n16256_, new_n16257_, new_n16258_, new_n16259_,
    new_n16260_, new_n16261_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16269_, new_n16270_,
    new_n16271_, new_n16272_, new_n16273_, new_n16274_, new_n16275_,
    new_n16276_, new_n16277_, new_n16278_, new_n16279_, new_n16280_,
    new_n16281_, new_n16282_, new_n16283_, new_n16284_, new_n16285_,
    new_n16286_, new_n16287_, new_n16288_, new_n16289_, new_n16290_,
    new_n16291_, new_n16292_, new_n16293_, new_n16294_, new_n16295_,
    new_n16296_, new_n16297_, new_n16298_, new_n16299_, new_n16300_,
    new_n16301_, new_n16302_, new_n16303_, new_n16304_, new_n16305_,
    new_n16306_, new_n16307_, new_n16308_, new_n16309_, new_n16310_,
    new_n16311_, new_n16312_, new_n16313_, new_n16314_, new_n16315_,
    new_n16316_, new_n16317_, new_n16318_, new_n16319_, new_n16320_,
    new_n16321_, new_n16322_, new_n16323_, new_n16324_, new_n16325_,
    new_n16326_, new_n16327_, new_n16328_, new_n16329_, new_n16330_,
    new_n16331_, new_n16332_, new_n16333_, new_n16334_, new_n16335_,
    new_n16336_, new_n16337_, new_n16338_, new_n16339_, new_n16340_,
    new_n16341_, new_n16342_, new_n16343_, new_n16344_, new_n16345_,
    new_n16346_, new_n16347_, new_n16348_, new_n16350_, new_n16351_,
    new_n16352_, new_n16353_, new_n16354_, new_n16355_, new_n16356_,
    new_n16357_, new_n16358_, new_n16359_, new_n16360_, new_n16361_,
    new_n16362_, new_n16363_, new_n16364_, new_n16365_, new_n16366_,
    new_n16367_, new_n16368_, new_n16369_, new_n16370_, new_n16371_,
    new_n16372_, new_n16373_, new_n16374_, new_n16375_, new_n16376_,
    new_n16377_, new_n16378_, new_n16379_, new_n16380_, new_n16381_,
    new_n16382_, new_n16383_, new_n16384_, new_n16385_, new_n16386_,
    new_n16387_, new_n16388_, new_n16389_, new_n16390_, new_n16391_,
    new_n16392_, new_n16393_, new_n16394_, new_n16395_, new_n16396_,
    new_n16397_, new_n16398_, new_n16399_, new_n16400_, new_n16401_,
    new_n16402_, new_n16403_, new_n16404_, new_n16405_, new_n16406_,
    new_n16407_, new_n16408_, new_n16409_, new_n16410_, new_n16411_,
    new_n16412_, new_n16413_, new_n16414_, new_n16415_, new_n16416_,
    new_n16417_, new_n16418_, new_n16419_, new_n16420_, new_n16421_,
    new_n16422_, new_n16423_, new_n16424_, new_n16425_, new_n16427_,
    new_n16428_, new_n16429_, new_n16430_, new_n16431_, new_n16432_,
    new_n16433_, new_n16434_, new_n16435_, new_n16436_, new_n16437_,
    new_n16438_, new_n16439_, new_n16440_, new_n16441_, new_n16442_,
    new_n16443_, new_n16444_, new_n16445_, new_n16446_, new_n16447_,
    new_n16448_, new_n16449_, new_n16450_, new_n16451_, new_n16452_,
    new_n16453_, new_n16454_, new_n16455_, new_n16456_, new_n16457_,
    new_n16458_, new_n16459_, new_n16460_, new_n16461_, new_n16462_,
    new_n16463_, new_n16464_, new_n16465_, new_n16466_, new_n16467_,
    new_n16468_, new_n16469_, new_n16470_, new_n16471_, new_n16472_,
    new_n16473_, new_n16474_, new_n16475_, new_n16476_, new_n16477_,
    new_n16478_, new_n16479_, new_n16480_, new_n16481_, new_n16482_,
    new_n16483_, new_n16484_, new_n16485_, new_n16486_, new_n16487_,
    new_n16488_, new_n16489_, new_n16490_, new_n16491_, new_n16492_,
    new_n16493_, new_n16494_, new_n16495_, new_n16496_, new_n16497_,
    new_n16498_, new_n16499_, new_n16500_, new_n16501_, new_n16502_,
    new_n16504_, new_n16505_, new_n16506_, new_n16507_, new_n16508_,
    new_n16509_, new_n16510_, new_n16511_, new_n16512_, new_n16513_,
    new_n16514_, new_n16515_, new_n16516_, new_n16517_, new_n16518_,
    new_n16519_, new_n16520_, new_n16521_, new_n16522_, new_n16523_,
    new_n16524_, new_n16525_, new_n16526_, new_n16527_, new_n16528_,
    new_n16529_, new_n16530_, new_n16531_, new_n16532_, new_n16533_,
    new_n16534_, new_n16535_, new_n16536_, new_n16537_, new_n16538_,
    new_n16539_, new_n16540_, new_n16541_, new_n16542_, new_n16543_,
    new_n16544_, new_n16545_, new_n16546_, new_n16547_, new_n16548_,
    new_n16549_, new_n16550_, new_n16551_, new_n16552_, new_n16553_,
    new_n16554_, new_n16555_, new_n16556_, new_n16558_, new_n16559_,
    new_n16560_, new_n16562_, new_n16563_, new_n16564_, new_n16565_,
    new_n16566_, new_n16567_, new_n16568_, new_n16569_, new_n16570_,
    new_n16571_, new_n16572_, new_n16573_, new_n16574_, new_n16575_,
    new_n16576_, new_n16577_, new_n16578_, new_n16579_, new_n16580_,
    new_n16581_, new_n16582_, new_n16583_, new_n16584_, new_n16585_,
    new_n16586_, new_n16587_, new_n16588_, new_n16589_, new_n16590_,
    new_n16591_, new_n16592_, new_n16593_, new_n16594_, new_n16595_,
    new_n16596_, new_n16597_, new_n16598_, new_n16599_, new_n16600_,
    new_n16601_, new_n16602_, new_n16603_, new_n16604_, new_n16605_,
    new_n16606_, new_n16607_, new_n16608_, new_n16609_, new_n16610_,
    new_n16611_, new_n16612_, new_n16613_, new_n16614_, new_n16615_,
    new_n16616_, new_n16617_, new_n16618_, new_n16619_, new_n16620_,
    new_n16621_, new_n16622_, new_n16623_, new_n16624_, new_n16625_,
    new_n16626_, new_n16627_, new_n16628_, new_n16629_, new_n16630_,
    new_n16631_, new_n16632_, new_n16633_, new_n16634_, new_n16635_,
    new_n16636_, new_n16637_, new_n16638_, new_n16639_, new_n16640_,
    new_n16641_, new_n16642_, new_n16643_, new_n16644_, new_n16645_,
    new_n16646_, new_n16647_, new_n16648_, new_n16649_, new_n16650_,
    new_n16651_, new_n16652_, new_n16653_, new_n16654_, new_n16655_,
    new_n16656_, new_n16657_, new_n16658_, new_n16659_, new_n16660_,
    new_n16661_, new_n16662_, new_n16664_, new_n16665_, new_n16666_,
    new_n16667_, new_n16668_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16722_, new_n16723_, new_n16724_, new_n16725_, new_n16726_,
    new_n16727_, new_n16728_, new_n16730_, new_n16731_, new_n16732_,
    new_n16733_, new_n16734_, new_n16735_, new_n16736_, new_n16737_,
    new_n16738_, new_n16739_, new_n16740_, new_n16741_, new_n16742_,
    new_n16743_, new_n16744_, new_n16745_, new_n16746_, new_n16747_,
    new_n16748_, new_n16749_, new_n16750_, new_n16751_, new_n16752_,
    new_n16753_, new_n16754_, new_n16755_, new_n16756_, new_n16757_,
    new_n16758_, new_n16759_, new_n16760_, new_n16761_, new_n16762_,
    new_n16763_, new_n16764_, new_n16765_, new_n16766_, new_n16767_,
    new_n16768_, new_n16769_, new_n16770_, new_n16771_, new_n16772_,
    new_n16773_, new_n16774_, new_n16775_, new_n16776_, new_n16777_,
    new_n16778_, new_n16779_, new_n16780_, new_n16782_, new_n16783_,
    new_n16784_, new_n16785_, new_n16786_, new_n16787_, new_n16788_,
    new_n16789_, new_n16790_, new_n16791_, new_n16792_, new_n16793_,
    new_n16794_, new_n16795_, new_n16796_, new_n16797_, new_n16798_,
    new_n16799_, new_n16800_, new_n16801_, new_n16802_, new_n16803_,
    new_n16804_, new_n16805_, new_n16806_, new_n16807_, new_n16808_,
    new_n16809_, new_n16810_, new_n16811_, new_n16812_, new_n16813_,
    new_n16814_, new_n16815_, new_n16816_, new_n16817_, new_n16818_,
    new_n16819_, new_n16820_, new_n16821_, new_n16822_, new_n16823_,
    new_n16824_, new_n16825_, new_n16826_, new_n16827_, new_n16828_,
    new_n16829_, new_n16830_, new_n16831_, new_n16832_, new_n16833_,
    new_n16834_, new_n16835_, new_n16836_, new_n16838_, new_n16839_,
    new_n16840_, new_n16841_, new_n16842_, new_n16843_, new_n16844_,
    new_n16845_, new_n16846_, new_n16847_, new_n16848_, new_n16849_,
    new_n16850_, new_n16851_, new_n16852_, new_n16853_, new_n16854_,
    new_n16855_, new_n16856_, new_n16857_, new_n16858_, new_n16859_,
    new_n16860_, new_n16861_, new_n16862_, new_n16863_, new_n16864_,
    new_n16865_, new_n16866_, new_n16867_, new_n16868_, new_n16869_,
    new_n16870_, new_n16871_, new_n16872_, new_n16873_, new_n16874_,
    new_n16876_, new_n16877_, new_n16878_, new_n16879_, new_n16880_,
    new_n16881_, new_n16883_, new_n16884_, new_n16885_, new_n16886_,
    new_n16887_, new_n16888_, new_n16889_, new_n16890_, new_n16891_,
    new_n16892_, new_n16893_, new_n16894_, new_n16895_, new_n16896_,
    new_n16897_, new_n16898_, new_n16899_, new_n16900_, new_n16901_,
    new_n16902_, new_n16903_, new_n16904_, new_n16905_, new_n16906_,
    new_n16907_, new_n16908_, new_n16909_, new_n16910_, new_n16911_,
    new_n16912_, new_n16913_, new_n16914_, new_n16915_, new_n16916_,
    new_n16917_, new_n16918_, new_n16919_, new_n16920_, new_n16921_,
    new_n16922_, new_n16923_, new_n16924_, new_n16925_, new_n16926_,
    new_n16927_, new_n16928_, new_n16929_, new_n16930_, new_n16931_,
    new_n16932_, new_n16934_, new_n16935_, new_n16936_, new_n16937_,
    new_n16938_, new_n16939_, new_n16940_, new_n16941_, new_n16942_,
    new_n16943_, new_n16944_, new_n16945_, new_n16946_, new_n16947_,
    new_n16948_, new_n16949_, new_n16950_, new_n16951_, new_n16952_,
    new_n16953_, new_n16954_, new_n16955_, new_n16956_, new_n16957_,
    new_n16958_, new_n16959_, new_n16960_, new_n16961_, new_n16962_,
    new_n16963_, new_n16964_, new_n16965_, new_n16967_, new_n16968_,
    new_n16969_, new_n16970_, new_n16971_, new_n16972_, new_n16973_,
    new_n16974_, new_n16975_, new_n16976_, new_n16977_, new_n16978_,
    new_n16979_, new_n16980_, new_n16981_, new_n16982_, new_n16983_,
    new_n16984_, new_n16985_, new_n16986_, new_n16987_, new_n16988_,
    new_n16989_, new_n16990_, new_n16991_, new_n16992_, new_n16993_,
    new_n16994_, new_n16995_, new_n16997_, new_n16998_, new_n16999_,
    new_n17000_, new_n17001_, new_n17002_, new_n17003_, new_n17004_,
    new_n17005_, new_n17006_, new_n17007_, new_n17008_, new_n17009_,
    new_n17010_, new_n17011_, new_n17012_, new_n17013_, new_n17014_,
    new_n17015_, new_n17016_, new_n17017_, new_n17018_, new_n17019_,
    new_n17020_, new_n17021_, new_n17022_, new_n17023_, new_n17025_,
    new_n17026_, new_n17027_, new_n17028_, new_n17029_, new_n17030_,
    new_n17031_, new_n17032_, new_n17033_, new_n17034_, new_n17035_,
    new_n17036_, new_n17037_, new_n17038_, new_n17040_, new_n17041_,
    new_n17042_, new_n17043_, new_n17044_, new_n17045_, new_n17046_,
    new_n17047_, new_n17048_, new_n17049_, new_n17050_, new_n17051_,
    new_n17052_, new_n17053_, new_n17054_, new_n17056_, new_n17057_,
    new_n17058_, new_n17059_, new_n17060_, new_n17061_, new_n17062_,
    new_n17063_, new_n17064_, new_n17065_, new_n17066_, new_n17067_,
    new_n17068_, new_n17069_, new_n17071_, new_n17072_, new_n17073_,
    new_n17074_, new_n17075_, new_n17076_, new_n17077_, new_n17078_,
    new_n17079_, new_n17080_, new_n17082_, new_n17083_, new_n17084_,
    new_n17085_, new_n17086_, new_n17087_, new_n17088_, new_n17089_,
    new_n17090_, new_n17092_;
  INV_X1     g00000(.I(\a[1] ), .ZN(new_n194_));
  NOR2_X1    g00001(.A1(new_n194_), .A2(\a[0] ), .ZN(\asquared[2] ));
  NAND2_X1   g00002(.A1(\a[0] ), .A2(\a[1] ), .ZN(new_n196_));
  NAND2_X1   g00003(.A1(\a[0] ), .A2(\a[2] ), .ZN(new_n197_));
  XOR2_X1    g00004(.A1(new_n196_), .A2(new_n197_), .Z(\asquared[3] ));
  INV_X1     g00005(.I(\a[0] ), .ZN(new_n199_));
  INV_X1     g00006(.I(\a[3] ), .ZN(new_n200_));
  INV_X1     g00007(.I(\a[2] ), .ZN(new_n201_));
  NOR2_X1    g00008(.A1(new_n194_), .A2(new_n201_), .ZN(new_n202_));
  NAND2_X1   g00009(.A1(new_n202_), .A2(new_n200_), .ZN(new_n203_));
  OAI21_X1   g00010(.A1(new_n194_), .A2(new_n201_), .B(\a[3] ), .ZN(new_n204_));
  AOI22_X1   g00011(.A1(new_n203_), .A2(new_n204_), .B1(new_n199_), .B2(new_n194_), .ZN(\asquared[4] ));
  NAND2_X1   g00012(.A1(\a[1] ), .A2(\a[4] ), .ZN(new_n206_));
  INV_X1     g00013(.I(new_n206_), .ZN(new_n207_));
  NOR4_X1    g00014(.A1(new_n207_), .A2(new_n199_), .A3(new_n201_), .A4(new_n200_), .ZN(new_n208_));
  XOR2_X1    g00015(.A1(new_n208_), .A2(new_n194_), .Z(new_n209_));
  XOR2_X1    g00016(.A1(new_n209_), .A2(new_n201_), .Z(\asquared[5] ));
  NAND2_X1   g00017(.A1(\a[4] ), .A2(\a[5] ), .ZN(new_n211_));
  NAND2_X1   g00018(.A1(\a[3] ), .A2(\a[4] ), .ZN(new_n212_));
  MUX2_X1    g00019(.I0(new_n212_), .I1(new_n196_), .S(new_n211_), .Z(new_n213_));
  NAND2_X1   g00020(.A1(\a[0] ), .A2(\a[3] ), .ZN(new_n214_));
  NAND2_X1   g00021(.A1(new_n207_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1     g00022(.I(new_n214_), .ZN(new_n216_));
  NAND2_X1   g00023(.A1(new_n216_), .A2(new_n206_), .ZN(new_n217_));
  INV_X1     g00024(.I(new_n197_), .ZN(new_n218_));
  NAND2_X1   g00025(.A1(new_n218_), .A2(\a[3] ), .ZN(new_n219_));
  NAND3_X1   g00026(.A1(new_n215_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  AOI21_X1   g00027(.A1(new_n220_), .A2(new_n202_), .B(new_n208_), .ZN(new_n221_));
  NOR2_X1    g00028(.A1(new_n221_), .A2(new_n213_), .ZN(new_n222_));
  XOR2_X1    g00029(.A1(new_n222_), .A2(new_n201_), .Z(new_n223_));
  XOR2_X1    g00030(.A1(new_n223_), .A2(new_n200_), .Z(\asquared[6] ));
  NAND2_X1   g00031(.A1(\a[2] ), .A2(\a[3] ), .ZN(new_n225_));
  AOI21_X1   g00032(.A1(new_n221_), .A2(new_n213_), .B(new_n225_), .ZN(new_n226_));
  NOR2_X1    g00033(.A1(new_n226_), .A2(new_n222_), .ZN(new_n227_));
  INV_X1     g00034(.I(new_n196_), .ZN(new_n228_));
  INV_X1     g00035(.I(new_n211_), .ZN(new_n229_));
  OAI21_X1   g00036(.A1(new_n196_), .A2(new_n211_), .B(new_n212_), .ZN(new_n230_));
  OAI21_X1   g00037(.A1(new_n228_), .A2(new_n229_), .B(new_n230_), .ZN(new_n231_));
  INV_X1     g00038(.I(new_n225_), .ZN(new_n232_));
  NAND2_X1   g00039(.A1(\a[2] ), .A2(\a[5] ), .ZN(new_n233_));
  XOR2_X1    g00040(.A1(new_n206_), .A2(new_n233_), .Z(new_n234_));
  NAND3_X1   g00041(.A1(new_n234_), .A2(new_n199_), .A3(new_n232_), .ZN(new_n235_));
  NOR2_X1    g00042(.A1(new_n207_), .A2(new_n233_), .ZN(new_n236_));
  INV_X1     g00043(.I(new_n233_), .ZN(new_n237_));
  NOR2_X1    g00044(.A1(new_n237_), .A2(new_n206_), .ZN(new_n238_));
  OAI21_X1   g00045(.A1(new_n236_), .A2(new_n238_), .B(new_n232_), .ZN(new_n239_));
  NAND2_X1   g00046(.A1(new_n239_), .A2(\a[0] ), .ZN(new_n240_));
  AOI21_X1   g00047(.A1(new_n240_), .A2(new_n235_), .B(\a[6] ), .ZN(new_n241_));
  INV_X1     g00048(.I(\a[6] ), .ZN(new_n242_));
  NOR2_X1    g00049(.A1(new_n239_), .A2(\a[0] ), .ZN(new_n243_));
  AOI21_X1   g00050(.A1(new_n234_), .A2(new_n232_), .B(new_n199_), .ZN(new_n244_));
  NOR3_X1    g00051(.A1(new_n243_), .A2(new_n244_), .A3(new_n242_), .ZN(new_n245_));
  NOR2_X1    g00052(.A1(new_n245_), .A2(new_n241_), .ZN(new_n246_));
  XOR2_X1    g00053(.A1(new_n246_), .A2(new_n231_), .Z(new_n247_));
  OAI21_X1   g00054(.A1(new_n245_), .A2(new_n241_), .B(new_n231_), .ZN(new_n248_));
  INV_X1     g00055(.I(new_n231_), .ZN(new_n249_));
  NAND2_X1   g00056(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1   g00057(.A1(new_n250_), .A2(new_n248_), .ZN(new_n251_));
  NAND2_X1   g00058(.A1(new_n251_), .A2(new_n227_), .ZN(new_n252_));
  OAI21_X1   g00059(.A1(new_n227_), .A2(new_n247_), .B(new_n252_), .ZN(\asquared[7] ));
  NOR2_X1    g00060(.A1(new_n246_), .A2(new_n249_), .ZN(new_n254_));
  OAI21_X1   g00061(.A1(new_n227_), .A2(new_n254_), .B(new_n250_), .ZN(new_n255_));
  NAND2_X1   g00062(.A1(new_n211_), .A2(new_n225_), .ZN(new_n256_));
  NAND2_X1   g00063(.A1(\a[0] ), .A2(\a[4] ), .ZN(new_n257_));
  NAND2_X1   g00064(.A1(\a[3] ), .A2(\a[7] ), .ZN(new_n258_));
  NOR2_X1    g00065(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1   g00066(.A1(\a[2] ), .A2(\a[4] ), .ZN(new_n260_));
  NAND2_X1   g00067(.A1(\a[3] ), .A2(\a[5] ), .ZN(new_n261_));
  NOR2_X1    g00068(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1   g00069(.A1(\a[0] ), .A2(\a[5] ), .ZN(new_n263_));
  NAND2_X1   g00070(.A1(\a[2] ), .A2(\a[7] ), .ZN(new_n264_));
  NOR2_X1    g00071(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND4_X1   g00072(.A1(new_n259_), .A2(new_n262_), .A3(new_n265_), .A4(new_n256_), .ZN(new_n266_));
  INV_X1     g00073(.I(new_n212_), .ZN(new_n267_));
  INV_X1     g00074(.I(\a[7] ), .ZN(new_n268_));
  NOR4_X1    g00075(.A1(new_n260_), .A2(new_n261_), .A3(new_n199_), .A4(new_n268_), .ZN(new_n269_));
  OAI21_X1   g00076(.A1(new_n269_), .A2(new_n265_), .B(new_n267_), .ZN(new_n270_));
  NAND2_X1   g00077(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1     g00078(.I(new_n271_), .ZN(new_n272_));
  INV_X1     g00079(.I(new_n239_), .ZN(new_n273_));
  NOR2_X1    g00080(.A1(new_n236_), .A2(new_n238_), .ZN(new_n274_));
  NOR2_X1    g00081(.A1(new_n199_), .A2(new_n242_), .ZN(new_n275_));
  INV_X1     g00082(.I(new_n275_), .ZN(new_n276_));
  AOI21_X1   g00083(.A1(new_n274_), .A2(new_n225_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1   g00084(.A1(\a[1] ), .A2(\a[6] ), .ZN(new_n278_));
  NOR2_X1    g00085(.A1(new_n206_), .A2(new_n233_), .ZN(new_n279_));
  INV_X1     g00086(.I(new_n279_), .ZN(new_n280_));
  OAI21_X1   g00087(.A1(new_n233_), .A2(new_n194_), .B(\a[4] ), .ZN(new_n281_));
  INV_X1     g00088(.I(\a[4] ), .ZN(new_n282_));
  NOR2_X1    g00089(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  AOI22_X1   g00090(.A1(new_n280_), .A2(new_n283_), .B1(new_n278_), .B2(new_n281_), .ZN(new_n284_));
  NOR3_X1    g00091(.A1(new_n277_), .A2(new_n273_), .A3(new_n284_), .ZN(new_n285_));
  OAI21_X1   g00092(.A1(new_n234_), .A2(new_n232_), .B(new_n275_), .ZN(new_n286_));
  NAND2_X1   g00093(.A1(new_n281_), .A2(new_n278_), .ZN(new_n287_));
  INV_X1     g00094(.I(new_n283_), .ZN(new_n288_));
  OAI21_X1   g00095(.A1(new_n279_), .A2(new_n288_), .B(new_n287_), .ZN(new_n289_));
  AOI21_X1   g00096(.A1(new_n286_), .A2(new_n239_), .B(new_n289_), .ZN(new_n290_));
  NOR2_X1    g00097(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1    g00098(.A1(new_n291_), .A2(new_n272_), .Z(new_n292_));
  NAND2_X1   g00099(.A1(new_n255_), .A2(new_n292_), .ZN(new_n293_));
  XOR2_X1    g00100(.A1(new_n291_), .A2(new_n272_), .Z(new_n294_));
  OAI21_X1   g00101(.A1(new_n255_), .A2(new_n294_), .B(new_n293_), .ZN(\asquared[8] ));
  NOR2_X1    g00102(.A1(new_n266_), .A2(new_n270_), .ZN(new_n296_));
  OAI21_X1   g00103(.A1(new_n285_), .A2(new_n290_), .B(new_n296_), .ZN(new_n297_));
  OAI21_X1   g00104(.A1(new_n297_), .A2(new_n246_), .B(new_n231_), .ZN(new_n298_));
  AOI21_X1   g00105(.A1(new_n246_), .A2(new_n297_), .B(new_n227_), .ZN(new_n299_));
  NAND2_X1   g00106(.A1(new_n299_), .A2(new_n298_), .ZN(new_n300_));
  OAI21_X1   g00107(.A1(new_n285_), .A2(new_n290_), .B(new_n271_), .ZN(new_n301_));
  INV_X1     g00108(.I(new_n301_), .ZN(new_n302_));
  NOR3_X1    g00109(.A1(new_n259_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n303_));
  NAND3_X1   g00110(.A1(new_n197_), .A2(\a[6] ), .A3(\a[8] ), .ZN(new_n304_));
  NAND2_X1   g00111(.A1(\a[6] ), .A2(\a[8] ), .ZN(new_n305_));
  NAND2_X1   g00112(.A1(new_n218_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1   g00113(.A1(\a[1] ), .A2(\a[7] ), .ZN(new_n307_));
  INV_X1     g00114(.I(new_n307_), .ZN(new_n308_));
  NAND3_X1   g00115(.A1(new_n306_), .A2(new_n304_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1   g00116(.A1(new_n306_), .A2(new_n304_), .B(new_n308_), .ZN(new_n310_));
  INV_X1     g00117(.I(new_n310_), .ZN(new_n311_));
  AOI21_X1   g00118(.A1(new_n311_), .A2(new_n309_), .B(new_n303_), .ZN(new_n312_));
  INV_X1     g00119(.I(new_n303_), .ZN(new_n313_));
  INV_X1     g00120(.I(new_n309_), .ZN(new_n314_));
  NOR3_X1    g00121(.A1(new_n314_), .A2(new_n313_), .A3(new_n310_), .ZN(new_n315_));
  OAI21_X1   g00122(.A1(new_n312_), .A2(new_n315_), .B(new_n261_), .ZN(new_n316_));
  INV_X1     g00123(.I(new_n261_), .ZN(new_n317_));
  OAI21_X1   g00124(.A1(new_n314_), .A2(new_n310_), .B(new_n313_), .ZN(new_n318_));
  NAND3_X1   g00125(.A1(new_n311_), .A2(new_n303_), .A3(new_n309_), .ZN(new_n319_));
  NAND3_X1   g00126(.A1(new_n318_), .A2(new_n319_), .A3(new_n317_), .ZN(new_n320_));
  NAND2_X1   g00127(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1     g00128(.I(new_n278_), .ZN(new_n322_));
  OAI22_X1   g00129(.A1(new_n277_), .A2(new_n273_), .B1(new_n322_), .B2(new_n280_), .ZN(new_n323_));
  NOR2_X1    g00130(.A1(new_n322_), .A2(\a[4] ), .ZN(new_n324_));
  OAI21_X1   g00131(.A1(new_n283_), .A2(new_n324_), .B(new_n280_), .ZN(new_n325_));
  NAND2_X1   g00132(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1   g00133(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  XOR2_X1    g00134(.A1(new_n327_), .A2(new_n302_), .Z(new_n328_));
  XOR2_X1    g00135(.A1(new_n328_), .A2(new_n300_), .Z(\asquared[9] ));
  NAND2_X1   g00136(.A1(new_n321_), .A2(new_n302_), .ZN(new_n330_));
  NAND3_X1   g00137(.A1(new_n301_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n331_));
  NAND4_X1   g00138(.A1(new_n299_), .A2(new_n298_), .A3(new_n331_), .A4(new_n326_), .ZN(new_n332_));
  NAND2_X1   g00139(.A1(new_n332_), .A2(new_n330_), .ZN(new_n333_));
  INV_X1     g00140(.I(new_n333_), .ZN(new_n334_));
  NAND2_X1   g00141(.A1(new_n306_), .A2(new_n304_), .ZN(new_n335_));
  INV_X1     g00142(.I(new_n335_), .ZN(new_n336_));
  NOR2_X1    g00143(.A1(new_n336_), .A2(new_n313_), .ZN(new_n337_));
  NAND2_X1   g00144(.A1(new_n336_), .A2(new_n313_), .ZN(new_n338_));
  XOR2_X1    g00145(.A1(new_n261_), .A2(new_n307_), .Z(new_n339_));
  AOI21_X1   g00146(.A1(new_n338_), .A2(new_n339_), .B(new_n337_), .ZN(new_n340_));
  NAND2_X1   g00147(.A1(\a[6] ), .A2(\a[8] ), .ZN(new_n341_));
  INV_X1     g00148(.I(new_n341_), .ZN(new_n342_));
  AOI21_X1   g00149(.A1(new_n283_), .A2(new_n218_), .B(new_n342_), .ZN(new_n343_));
  INV_X1     g00150(.I(new_n264_), .ZN(new_n344_));
  NAND4_X1   g00151(.A1(\a[2] ), .A2(\a[4] ), .A3(\a[5] ), .A4(\a[7] ), .ZN(new_n345_));
  NAND4_X1   g00152(.A1(\a[2] ), .A2(\a[3] ), .A3(\a[6] ), .A4(\a[7] ), .ZN(new_n346_));
  NAND2_X1   g00153(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1     g00154(.I(new_n347_), .ZN(new_n348_));
  NAND4_X1   g00155(.A1(\a[3] ), .A2(\a[4] ), .A3(\a[5] ), .A4(\a[6] ), .ZN(new_n349_));
  AOI21_X1   g00156(.A1(\a[3] ), .A2(\a[6] ), .B(new_n229_), .ZN(new_n350_));
  NOR4_X1    g00157(.A1(new_n348_), .A2(new_n350_), .A3(new_n344_), .A4(new_n349_), .ZN(new_n351_));
  NAND4_X1   g00158(.A1(\a[1] ), .A2(\a[3] ), .A3(\a[5] ), .A4(\a[7] ), .ZN(new_n352_));
  INV_X1     g00159(.I(\a[5] ), .ZN(new_n353_));
  NAND2_X1   g00160(.A1(\a[1] ), .A2(\a[8] ), .ZN(new_n354_));
  NAND2_X1   g00161(.A1(new_n354_), .A2(new_n353_), .ZN(new_n355_));
  NAND3_X1   g00162(.A1(\a[1] ), .A2(\a[5] ), .A3(\a[8] ), .ZN(new_n356_));
  AOI21_X1   g00163(.A1(new_n355_), .A2(new_n356_), .B(new_n352_), .ZN(new_n357_));
  NAND2_X1   g00164(.A1(new_n357_), .A2(new_n199_), .ZN(new_n358_));
  INV_X1     g00165(.I(\a[8] ), .ZN(new_n359_));
  NOR2_X1    g00166(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  AOI22_X1   g00167(.A1(new_n360_), .A2(\a[1] ), .B1(new_n353_), .B2(new_n354_), .ZN(new_n361_));
  OAI21_X1   g00168(.A1(new_n361_), .A2(new_n352_), .B(\a[0] ), .ZN(new_n362_));
  AOI21_X1   g00169(.A1(new_n362_), .A2(new_n358_), .B(\a[9] ), .ZN(new_n363_));
  INV_X1     g00170(.I(\a[9] ), .ZN(new_n364_));
  NOR3_X1    g00171(.A1(new_n361_), .A2(\a[0] ), .A3(new_n352_), .ZN(new_n365_));
  NOR2_X1    g00172(.A1(new_n357_), .A2(new_n199_), .ZN(new_n366_));
  NOR3_X1    g00173(.A1(new_n365_), .A2(new_n366_), .A3(new_n364_), .ZN(new_n367_));
  OAI21_X1   g00174(.A1(new_n367_), .A2(new_n363_), .B(new_n351_), .ZN(new_n368_));
  NOR3_X1    g00175(.A1(new_n350_), .A2(new_n344_), .A3(new_n349_), .ZN(new_n369_));
  NAND2_X1   g00176(.A1(new_n369_), .A2(new_n347_), .ZN(new_n370_));
  OAI21_X1   g00177(.A1(new_n365_), .A2(new_n366_), .B(new_n364_), .ZN(new_n371_));
  NAND3_X1   g00178(.A1(new_n362_), .A2(new_n358_), .A3(\a[9] ), .ZN(new_n372_));
  NAND3_X1   g00179(.A1(new_n371_), .A2(new_n372_), .A3(new_n370_), .ZN(new_n373_));
  AOI21_X1   g00180(.A1(new_n368_), .A2(new_n373_), .B(new_n343_), .ZN(new_n374_));
  INV_X1     g00181(.I(new_n343_), .ZN(new_n375_));
  OAI21_X1   g00182(.A1(new_n367_), .A2(new_n363_), .B(new_n370_), .ZN(new_n376_));
  NAND3_X1   g00183(.A1(new_n371_), .A2(new_n372_), .A3(new_n351_), .ZN(new_n377_));
  AOI21_X1   g00184(.A1(new_n376_), .A2(new_n377_), .B(new_n375_), .ZN(new_n378_));
  NOR2_X1    g00185(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  XOR2_X1    g00186(.A1(new_n379_), .A2(new_n340_), .Z(new_n380_));
  INV_X1     g00187(.I(new_n340_), .ZN(new_n381_));
  NOR2_X1    g00188(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1     g00189(.I(new_n382_), .ZN(new_n383_));
  NAND2_X1   g00190(.A1(new_n379_), .A2(new_n381_), .ZN(new_n384_));
  NAND2_X1   g00191(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1   g00192(.A1(new_n385_), .A2(new_n334_), .ZN(new_n386_));
  OAI21_X1   g00193(.A1(new_n334_), .A2(new_n380_), .B(new_n386_), .ZN(\asquared[10] ));
  OAI21_X1   g00194(.A1(new_n334_), .A2(new_n382_), .B(new_n384_), .ZN(new_n388_));
  AOI21_X1   g00195(.A1(new_n371_), .A2(new_n372_), .B(new_n351_), .ZN(new_n389_));
  OAI21_X1   g00196(.A1(new_n343_), .A2(new_n389_), .B(new_n377_), .ZN(new_n390_));
  NAND2_X1   g00197(.A1(\a[8] ), .A2(\a[10] ), .ZN(new_n391_));
  NAND2_X1   g00198(.A1(\a[7] ), .A2(\a[8] ), .ZN(new_n392_));
  OAI22_X1   g00199(.A1(new_n197_), .A2(new_n392_), .B1(new_n225_), .B2(new_n391_), .ZN(new_n393_));
  INV_X1     g00200(.I(new_n393_), .ZN(new_n394_));
  NAND2_X1   g00201(.A1(\a[0] ), .A2(\a[10] ), .ZN(new_n395_));
  XNOR2_X1   g00202(.A1(new_n258_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1   g00203(.A1(new_n395_), .A2(\a[3] ), .A3(\a[7] ), .ZN(new_n397_));
  NOR2_X1    g00204(.A1(new_n201_), .A2(new_n359_), .ZN(new_n398_));
  INV_X1     g00205(.I(new_n398_), .ZN(new_n399_));
  AOI22_X1   g00206(.A1(new_n396_), .A2(new_n399_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n400_));
  INV_X1     g00207(.I(new_n400_), .ZN(new_n401_));
  NAND3_X1   g00208(.A1(new_n355_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n402_));
  NOR2_X1    g00209(.A1(new_n199_), .A2(new_n364_), .ZN(new_n403_));
  AOI21_X1   g00210(.A1(new_n402_), .A2(new_n403_), .B(new_n357_), .ZN(new_n404_));
  INV_X1     g00211(.I(new_n404_), .ZN(new_n405_));
  AOI21_X1   g00212(.A1(new_n345_), .A2(new_n349_), .B(new_n346_), .ZN(new_n406_));
  INV_X1     g00213(.I(new_n406_), .ZN(new_n407_));
  NOR2_X1    g00214(.A1(new_n354_), .A2(new_n353_), .ZN(new_n408_));
  INV_X1     g00215(.I(new_n408_), .ZN(new_n409_));
  NAND3_X1   g00216(.A1(new_n278_), .A2(\a[4] ), .A3(\a[9] ), .ZN(new_n410_));
  INV_X1     g00217(.I(new_n410_), .ZN(new_n411_));
  AOI21_X1   g00218(.A1(\a[4] ), .A2(\a[9] ), .B(new_n278_), .ZN(new_n412_));
  OAI21_X1   g00219(.A1(new_n411_), .A2(new_n412_), .B(new_n409_), .ZN(new_n413_));
  NAND2_X1   g00220(.A1(\a[4] ), .A2(\a[9] ), .ZN(new_n414_));
  NAND2_X1   g00221(.A1(new_n322_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1   g00222(.A1(new_n415_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n416_));
  AOI21_X1   g00223(.A1(new_n413_), .A2(new_n416_), .B(new_n407_), .ZN(new_n417_));
  OAI21_X1   g00224(.A1(new_n411_), .A2(new_n412_), .B(new_n408_), .ZN(new_n418_));
  NAND3_X1   g00225(.A1(new_n409_), .A2(new_n415_), .A3(new_n410_), .ZN(new_n419_));
  AOI21_X1   g00226(.A1(new_n418_), .A2(new_n419_), .B(new_n406_), .ZN(new_n420_));
  OAI21_X1   g00227(.A1(new_n417_), .A2(new_n420_), .B(new_n405_), .ZN(new_n421_));
  AOI21_X1   g00228(.A1(new_n415_), .A2(new_n410_), .B(new_n408_), .ZN(new_n422_));
  INV_X1     g00229(.I(new_n416_), .ZN(new_n423_));
  OAI21_X1   g00230(.A1(new_n423_), .A2(new_n422_), .B(new_n406_), .ZN(new_n424_));
  AOI21_X1   g00231(.A1(new_n415_), .A2(new_n410_), .B(new_n409_), .ZN(new_n425_));
  NOR3_X1    g00232(.A1(new_n411_), .A2(new_n408_), .A3(new_n412_), .ZN(new_n426_));
  OAI21_X1   g00233(.A1(new_n425_), .A2(new_n426_), .B(new_n407_), .ZN(new_n427_));
  NAND3_X1   g00234(.A1(new_n424_), .A2(new_n427_), .A3(new_n404_), .ZN(new_n428_));
  AOI21_X1   g00235(.A1(new_n428_), .A2(new_n421_), .B(new_n401_), .ZN(new_n429_));
  OAI21_X1   g00236(.A1(new_n417_), .A2(new_n420_), .B(new_n404_), .ZN(new_n430_));
  NAND3_X1   g00237(.A1(new_n424_), .A2(new_n427_), .A3(new_n405_), .ZN(new_n431_));
  AOI21_X1   g00238(.A1(new_n431_), .A2(new_n430_), .B(new_n400_), .ZN(new_n432_));
  NOR2_X1    g00239(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  XOR2_X1    g00240(.A1(new_n433_), .A2(new_n390_), .Z(new_n434_));
  NAND2_X1   g00241(.A1(new_n388_), .A2(new_n434_), .ZN(new_n435_));
  NOR3_X1    g00242(.A1(new_n367_), .A2(new_n363_), .A3(new_n370_), .ZN(new_n436_));
  AOI21_X1   g00243(.A1(new_n375_), .A2(new_n376_), .B(new_n436_), .ZN(new_n437_));
  OAI21_X1   g00244(.A1(new_n429_), .A2(new_n432_), .B(new_n437_), .ZN(new_n438_));
  AOI21_X1   g00245(.A1(new_n424_), .A2(new_n427_), .B(new_n404_), .ZN(new_n439_));
  NOR3_X1    g00246(.A1(new_n417_), .A2(new_n420_), .A3(new_n405_), .ZN(new_n440_));
  OAI21_X1   g00247(.A1(new_n439_), .A2(new_n440_), .B(new_n400_), .ZN(new_n441_));
  AOI21_X1   g00248(.A1(new_n424_), .A2(new_n427_), .B(new_n405_), .ZN(new_n442_));
  NOR3_X1    g00249(.A1(new_n417_), .A2(new_n420_), .A3(new_n404_), .ZN(new_n443_));
  OAI21_X1   g00250(.A1(new_n442_), .A2(new_n443_), .B(new_n401_), .ZN(new_n444_));
  NAND3_X1   g00251(.A1(new_n390_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  AND2_X2    g00252(.A1(new_n438_), .A2(new_n445_), .Z(new_n446_));
  OAI21_X1   g00253(.A1(new_n388_), .A2(new_n446_), .B(new_n435_), .ZN(\asquared[11] ));
  NAND2_X1   g00254(.A1(new_n445_), .A2(new_n379_), .ZN(new_n448_));
  OAI21_X1   g00255(.A1(new_n445_), .A2(new_n379_), .B(new_n340_), .ZN(new_n449_));
  NAND3_X1   g00256(.A1(new_n333_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  NOR2_X1    g00257(.A1(new_n258_), .A2(new_n395_), .ZN(new_n451_));
  NOR2_X1    g00258(.A1(new_n394_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1   g00259(.A1(\a[8] ), .A2(\a[9] ), .ZN(new_n453_));
  INV_X1     g00260(.I(new_n453_), .ZN(new_n454_));
  NAND4_X1   g00261(.A1(\a[1] ), .A2(\a[4] ), .A3(\a[6] ), .A4(\a[9] ), .ZN(new_n455_));
  NAND2_X1   g00262(.A1(new_n454_), .A2(new_n225_), .ZN(new_n457_));
  NAND2_X1   g00263(.A1(\a[8] ), .A2(\a[9] ), .ZN(new_n458_));
  NAND2_X1   g00264(.A1(new_n232_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1   g00265(.A1(\a[1] ), .A2(\a[10] ), .B(\a[6] ), .ZN(new_n460_));
  INV_X1     g00266(.I(\a[10] ), .ZN(new_n461_));
  NOR2_X1    g00267(.A1(new_n242_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1   g00268(.A1(new_n462_), .A2(\a[1] ), .B(new_n460_), .ZN(new_n463_));
  AOI21_X1   g00269(.A1(new_n457_), .A2(new_n459_), .B(new_n463_), .ZN(new_n464_));
  NOR2_X1    g00270(.A1(new_n232_), .A2(new_n458_), .ZN(new_n465_));
  NOR2_X1    g00271(.A1(new_n454_), .A2(new_n225_), .ZN(new_n466_));
  NOR2_X1    g00272(.A1(new_n194_), .A2(new_n461_), .ZN(new_n467_));
  NAND3_X1   g00273(.A1(\a[1] ), .A2(\a[6] ), .A3(\a[10] ), .ZN(new_n468_));
  OAI21_X1   g00274(.A1(new_n467_), .A2(\a[6] ), .B(new_n468_), .ZN(new_n469_));
  NOR3_X1    g00275(.A1(new_n469_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n470_));
  OAI21_X1   g00276(.A1(new_n464_), .A2(new_n470_), .B(new_n452_), .ZN(new_n471_));
  OAI21_X1   g00277(.A1(new_n258_), .A2(new_n395_), .B(new_n393_), .ZN(new_n472_));
  NOR3_X1    g00278(.A1(new_n463_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n473_));
  AOI21_X1   g00279(.A1(new_n457_), .A2(new_n459_), .B(new_n469_), .ZN(new_n474_));
  OAI21_X1   g00280(.A1(new_n474_), .A2(new_n473_), .B(new_n472_), .ZN(new_n475_));
  OAI21_X1   g00281(.A1(new_n425_), .A2(new_n407_), .B(new_n419_), .ZN(new_n476_));
  INV_X1     g00282(.I(new_n476_), .ZN(new_n477_));
  NAND2_X1   g00283(.A1(\a[6] ), .A2(\a[7] ), .ZN(new_n478_));
  INV_X1     g00284(.I(new_n478_), .ZN(new_n479_));
  NAND2_X1   g00285(.A1(\a[4] ), .A2(\a[7] ), .ZN(new_n480_));
  NAND2_X1   g00286(.A1(\a[5] ), .A2(\a[6] ), .ZN(new_n481_));
  NAND2_X1   g00287(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1   g00288(.A1(\a[0] ), .A2(\a[11] ), .ZN(new_n483_));
  NAND2_X1   g00289(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1   g00290(.A1(new_n484_), .A2(new_n211_), .A3(new_n479_), .ZN(new_n485_));
  NAND2_X1   g00291(.A1(new_n484_), .A2(new_n479_), .ZN(new_n486_));
  NAND2_X1   g00292(.A1(new_n486_), .A2(new_n229_), .ZN(new_n487_));
  NAND2_X1   g00293(.A1(new_n487_), .A2(new_n485_), .ZN(new_n488_));
  NAND2_X1   g00294(.A1(new_n477_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1   g00295(.A1(new_n476_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n490_));
  AOI22_X1   g00296(.A1(new_n489_), .A2(new_n490_), .B1(new_n471_), .B2(new_n475_), .ZN(new_n491_));
  NAND2_X1   g00297(.A1(new_n471_), .A2(new_n475_), .ZN(new_n492_));
  NAND2_X1   g00298(.A1(new_n488_), .A2(new_n476_), .ZN(new_n493_));
  NAND3_X1   g00299(.A1(new_n477_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n494_));
  AOI21_X1   g00300(.A1(new_n494_), .A2(new_n493_), .B(new_n492_), .ZN(new_n495_));
  NOR2_X1    g00301(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1   g00302(.A1(new_n400_), .A2(new_n430_), .B(new_n443_), .ZN(new_n497_));
  NOR2_X1    g00303(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XOR2_X1    g00304(.A1(new_n450_), .A2(new_n498_), .Z(new_n499_));
  XOR2_X1    g00305(.A1(new_n499_), .A2(new_n438_), .Z(\asquared[12] ));
  OR2_X2     g00306(.A1(new_n438_), .A2(new_n496_), .Z(new_n501_));
  AOI21_X1   g00307(.A1(new_n438_), .A2(new_n496_), .B(new_n497_), .ZN(new_n502_));
  NAND4_X1   g00308(.A1(new_n333_), .A2(new_n502_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n503_));
  NAND2_X1   g00309(.A1(new_n503_), .A2(new_n501_), .ZN(new_n504_));
  NAND2_X1   g00310(.A1(new_n494_), .A2(new_n492_), .ZN(new_n505_));
  AND2_X2    g00311(.A1(new_n505_), .A2(new_n493_), .Z(new_n506_));
  INV_X1     g00312(.I(new_n506_), .ZN(new_n507_));
  NOR2_X1    g00313(.A1(new_n278_), .A2(new_n461_), .ZN(new_n508_));
  NAND2_X1   g00314(.A1(\a[5] ), .A2(\a[11] ), .ZN(new_n509_));
  AOI21_X1   g00315(.A1(\a[1] ), .A2(\a[7] ), .B(new_n509_), .ZN(new_n510_));
  AOI21_X1   g00316(.A1(\a[5] ), .A2(\a[11] ), .B(new_n307_), .ZN(new_n511_));
  OAI21_X1   g00317(.A1(new_n510_), .A2(new_n511_), .B(new_n508_), .ZN(new_n512_));
  NOR2_X1    g00318(.A1(new_n512_), .A2(\a[4] ), .ZN(new_n513_));
  NAND3_X1   g00319(.A1(new_n307_), .A2(\a[5] ), .A3(\a[11] ), .ZN(new_n514_));
  NAND3_X1   g00320(.A1(new_n509_), .A2(\a[1] ), .A3(\a[7] ), .ZN(new_n515_));
  NAND2_X1   g00321(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1   g00322(.A1(new_n516_), .A2(new_n508_), .B(new_n282_), .ZN(new_n517_));
  OAI21_X1   g00323(.A1(new_n513_), .A2(new_n517_), .B(new_n359_), .ZN(new_n518_));
  NAND3_X1   g00324(.A1(new_n516_), .A2(new_n282_), .A3(new_n508_), .ZN(new_n519_));
  NAND2_X1   g00325(.A1(new_n512_), .A2(\a[4] ), .ZN(new_n520_));
  NAND3_X1   g00326(.A1(new_n520_), .A2(new_n519_), .A3(\a[8] ), .ZN(new_n521_));
  NAND2_X1   g00327(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1   g00328(.A1(\a[10] ), .A2(\a[12] ), .ZN(new_n523_));
  NOR2_X1    g00329(.A1(new_n200_), .A2(new_n364_), .ZN(new_n524_));
  NAND2_X1   g00330(.A1(\a[9] ), .A2(\a[10] ), .ZN(new_n525_));
  NAND2_X1   g00331(.A1(\a[0] ), .A2(\a[12] ), .ZN(new_n527_));
  NOR2_X1    g00332(.A1(new_n197_), .A2(new_n523_), .ZN(new_n531_));
  INV_X1     g00333(.I(new_n531_), .ZN(new_n532_));
  OAI21_X1   g00334(.A1(new_n455_), .A2(new_n453_), .B(new_n225_), .ZN(new_n533_));
  NAND3_X1   g00335(.A1(new_n479_), .A2(\a[0] ), .A3(\a[11] ), .ZN(new_n534_));
  NAND3_X1   g00336(.A1(new_n229_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n535_));
  AOI21_X1   g00337(.A1(new_n534_), .A2(new_n535_), .B(new_n533_), .ZN(new_n536_));
  NAND3_X1   g00338(.A1(new_n534_), .A2(new_n535_), .A3(new_n533_), .ZN(new_n537_));
  INV_X1     g00339(.I(new_n537_), .ZN(new_n538_));
  NOR2_X1    g00340(.A1(new_n538_), .A2(new_n536_), .ZN(new_n539_));
  OAI21_X1   g00341(.A1(new_n465_), .A2(new_n466_), .B(new_n469_), .ZN(new_n540_));
  OAI21_X1   g00342(.A1(new_n472_), .A2(new_n470_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1   g00343(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1     g00344(.I(new_n542_), .ZN(new_n543_));
  NOR2_X1    g00345(.A1(new_n539_), .A2(new_n541_), .ZN(new_n544_));
  OAI21_X1   g00346(.A1(new_n543_), .A2(new_n544_), .B(new_n532_), .ZN(new_n545_));
  INV_X1     g00347(.I(new_n544_), .ZN(new_n546_));
  NAND3_X1   g00348(.A1(new_n546_), .A2(new_n531_), .A3(new_n542_), .ZN(new_n547_));
  AOI21_X1   g00349(.A1(new_n545_), .A2(new_n547_), .B(new_n522_), .ZN(new_n548_));
  AND3_X2    g00350(.A1(new_n545_), .A2(new_n547_), .A3(new_n522_), .Z(new_n549_));
  NOR2_X1    g00351(.A1(new_n549_), .A2(new_n548_), .ZN(new_n550_));
  XOR2_X1    g00352(.A1(new_n550_), .A2(new_n507_), .Z(new_n551_));
  OAI21_X1   g00353(.A1(new_n549_), .A2(new_n548_), .B(new_n506_), .ZN(new_n552_));
  NAND2_X1   g00354(.A1(new_n550_), .A2(new_n507_), .ZN(new_n553_));
  NAND2_X1   g00355(.A1(new_n553_), .A2(new_n552_), .ZN(new_n554_));
  MUX2_X1    g00356(.I0(new_n554_), .I1(new_n551_), .S(new_n504_), .Z(\asquared[13] ));
  NAND2_X1   g00357(.A1(new_n504_), .A2(new_n552_), .ZN(new_n556_));
  NAND2_X1   g00358(.A1(new_n556_), .A2(new_n553_), .ZN(new_n557_));
  NAND2_X1   g00359(.A1(new_n534_), .A2(new_n535_), .ZN(new_n558_));
  NOR2_X1    g00360(.A1(new_n558_), .A2(new_n533_), .ZN(new_n559_));
  INV_X1     g00361(.I(new_n559_), .ZN(new_n560_));
  INV_X1     g00362(.I(new_n536_), .ZN(new_n561_));
  AOI21_X1   g00363(.A1(new_n561_), .A2(new_n537_), .B(new_n531_), .ZN(new_n562_));
  OAI22_X1   g00364(.A1(new_n197_), .A2(new_n523_), .B1(new_n225_), .B2(new_n525_), .ZN(new_n563_));
  NAND2_X1   g00365(.A1(\a[1] ), .A2(\a[12] ), .ZN(new_n564_));
  INV_X1     g00366(.I(new_n564_), .ZN(new_n565_));
  INV_X1     g00367(.I(\a[12] ), .ZN(new_n566_));
  NAND3_X1   g00368(.A1(new_n509_), .A2(\a[7] ), .A3(new_n566_), .ZN(new_n567_));
  NOR2_X1    g00369(.A1(new_n567_), .A2(new_n565_), .ZN(new_n568_));
  NOR2_X1    g00370(.A1(new_n268_), .A2(\a[12] ), .ZN(new_n569_));
  AOI21_X1   g00371(.A1(new_n569_), .A2(new_n509_), .B(new_n564_), .ZN(new_n570_));
  NOR2_X1    g00372(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1    g00373(.A1(new_n571_), .A2(new_n563_), .Z(new_n572_));
  NAND3_X1   g00374(.A1(new_n463_), .A2(new_n459_), .A3(new_n457_), .ZN(new_n573_));
  AOI21_X1   g00375(.A1(new_n452_), .A2(new_n573_), .B(new_n464_), .ZN(new_n574_));
  AOI21_X1   g00376(.A1(new_n518_), .A2(new_n521_), .B(new_n574_), .ZN(new_n575_));
  NAND3_X1   g00377(.A1(new_n518_), .A2(new_n521_), .A3(new_n574_), .ZN(new_n576_));
  OAI21_X1   g00378(.A1(new_n538_), .A2(new_n536_), .B(new_n532_), .ZN(new_n577_));
  NAND3_X1   g00379(.A1(new_n561_), .A2(new_n531_), .A3(new_n537_), .ZN(new_n578_));
  NAND2_X1   g00380(.A1(new_n578_), .A2(new_n577_), .ZN(new_n579_));
  AOI21_X1   g00381(.A1(new_n576_), .A2(new_n579_), .B(new_n575_), .ZN(new_n580_));
  NOR3_X1    g00382(.A1(new_n580_), .A2(new_n562_), .A3(new_n572_), .ZN(new_n581_));
  INV_X1     g00383(.I(new_n572_), .ZN(new_n582_));
  AOI21_X1   g00384(.A1(new_n520_), .A2(new_n519_), .B(\a[8] ), .ZN(new_n583_));
  NOR3_X1    g00385(.A1(new_n513_), .A2(new_n359_), .A3(new_n517_), .ZN(new_n584_));
  OAI21_X1   g00386(.A1(new_n584_), .A2(new_n583_), .B(new_n541_), .ZN(new_n585_));
  NOR3_X1    g00387(.A1(new_n583_), .A2(new_n584_), .A3(new_n541_), .ZN(new_n586_));
  NOR3_X1    g00388(.A1(new_n538_), .A2(new_n532_), .A3(new_n536_), .ZN(new_n587_));
  NOR2_X1    g00389(.A1(new_n562_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1   g00390(.A1(new_n586_), .A2(new_n588_), .B(new_n585_), .ZN(new_n589_));
  AOI21_X1   g00391(.A1(new_n589_), .A2(new_n582_), .B(new_n577_), .ZN(new_n590_));
  OAI21_X1   g00392(.A1(new_n581_), .A2(new_n590_), .B(new_n560_), .ZN(new_n591_));
  NAND3_X1   g00393(.A1(new_n589_), .A2(new_n577_), .A3(new_n582_), .ZN(new_n592_));
  OAI21_X1   g00394(.A1(new_n580_), .A2(new_n572_), .B(new_n562_), .ZN(new_n593_));
  NAND3_X1   g00395(.A1(new_n593_), .A2(new_n592_), .A3(new_n559_), .ZN(new_n594_));
  AND2_X2    g00396(.A1(new_n591_), .A2(new_n594_), .Z(new_n595_));
  NAND2_X1   g00397(.A1(\a[9] ), .A2(\a[13] ), .ZN(new_n596_));
  INV_X1     g00398(.I(new_n525_), .ZN(new_n597_));
  INV_X1     g00399(.I(\a[13] ), .ZN(new_n599_));
  NOR2_X1    g00400(.A1(new_n257_), .A2(new_n596_), .ZN(new_n603_));
  INV_X1     g00401(.I(new_n512_), .ZN(new_n604_));
  NOR2_X1    g00402(.A1(new_n516_), .A2(new_n508_), .ZN(new_n605_));
  NOR3_X1    g00403(.A1(new_n605_), .A2(new_n282_), .A3(new_n359_), .ZN(new_n606_));
  NOR2_X1    g00404(.A1(new_n606_), .A2(new_n604_), .ZN(new_n607_));
  INV_X1     g00405(.I(new_n481_), .ZN(new_n608_));
  AND2_X2    g00406(.A1(\a[7] ), .A2(\a[8] ), .Z(new_n609_));
  NAND2_X1   g00407(.A1(\a[2] ), .A2(\a[11] ), .ZN(new_n610_));
  OAI21_X1   g00408(.A1(new_n360_), .A2(new_n479_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1   g00409(.A1(new_n611_), .A2(new_n609_), .ZN(new_n612_));
  XOR2_X1    g00410(.A1(new_n612_), .A2(new_n608_), .Z(new_n613_));
  XOR2_X1    g00411(.A1(new_n613_), .A2(new_n607_), .Z(new_n614_));
  OR2_X2     g00412(.A1(new_n613_), .A2(new_n607_), .Z(new_n615_));
  NAND2_X1   g00413(.A1(new_n613_), .A2(new_n607_), .ZN(new_n616_));
  AOI21_X1   g00414(.A1(new_n615_), .A2(new_n616_), .B(new_n603_), .ZN(new_n617_));
  AOI21_X1   g00415(.A1(new_n614_), .A2(new_n603_), .B(new_n617_), .ZN(new_n618_));
  XOR2_X1    g00416(.A1(new_n595_), .A2(new_n618_), .Z(new_n619_));
  NAND2_X1   g00417(.A1(new_n557_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1   g00418(.A1(new_n591_), .A2(new_n594_), .B(new_n618_), .ZN(new_n621_));
  NAND3_X1   g00419(.A1(new_n591_), .A2(new_n594_), .A3(new_n618_), .ZN(new_n622_));
  INV_X1     g00420(.I(new_n622_), .ZN(new_n623_));
  NOR2_X1    g00421(.A1(new_n623_), .A2(new_n621_), .ZN(new_n624_));
  OAI21_X1   g00422(.A1(new_n557_), .A2(new_n624_), .B(new_n620_), .ZN(\asquared[14] ));
  OAI21_X1   g00423(.A1(new_n622_), .A2(new_n550_), .B(new_n506_), .ZN(new_n626_));
  NAND2_X1   g00424(.A1(new_n622_), .A2(new_n550_), .ZN(new_n627_));
  NAND4_X1   g00425(.A1(new_n626_), .A2(new_n504_), .A3(new_n627_), .A4(new_n621_), .ZN(new_n628_));
  INV_X1     g00426(.I(new_n628_), .ZN(\asquared[15] ));
  OAI22_X1   g00427(.A1(new_n212_), .A2(new_n525_), .B1(new_n257_), .B2(new_n596_), .ZN(new_n630_));
  NAND4_X1   g00428(.A1(new_n268_), .A2(new_n359_), .A3(\a[5] ), .A4(\a[6] ), .ZN(new_n631_));
  OAI21_X1   g00429(.A1(new_n392_), .A2(new_n610_), .B(new_n631_), .ZN(new_n632_));
  NAND2_X1   g00430(.A1(\a[1] ), .A2(\a[13] ), .ZN(new_n633_));
  XNOR2_X1   g00431(.A1(new_n341_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1    g00432(.A1(new_n634_), .A2(new_n632_), .ZN(new_n635_));
  NOR2_X1    g00433(.A1(new_n392_), .A2(new_n610_), .ZN(new_n636_));
  INV_X1     g00434(.I(new_n631_), .ZN(new_n637_));
  NOR2_X1    g00435(.A1(new_n637_), .A2(new_n636_), .ZN(new_n638_));
  XOR2_X1    g00436(.A1(new_n341_), .A2(new_n633_), .Z(new_n639_));
  NOR2_X1    g00437(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1    g00438(.A1(new_n640_), .A2(new_n635_), .ZN(new_n641_));
  NOR2_X1    g00439(.A1(new_n641_), .A2(new_n630_), .ZN(new_n642_));
  XOR2_X1    g00440(.A1(new_n634_), .A2(new_n632_), .Z(new_n643_));
  AOI21_X1   g00441(.A1(new_n630_), .A2(new_n643_), .B(new_n642_), .ZN(new_n644_));
  NOR2_X1    g00442(.A1(new_n613_), .A2(new_n607_), .ZN(new_n645_));
  AOI21_X1   g00443(.A1(new_n603_), .A2(new_n616_), .B(new_n645_), .ZN(new_n646_));
  NOR2_X1    g00444(.A1(new_n646_), .A2(new_n644_), .ZN(new_n647_));
  NAND3_X1   g00445(.A1(new_n308_), .A2(\a[5] ), .A3(\a[11] ), .ZN(new_n648_));
  OAI22_X1   g00446(.A1(new_n571_), .A2(new_n566_), .B1(new_n563_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1     g00447(.I(\a[14] ), .ZN(new_n650_));
  NAND2_X1   g00448(.A1(\a[11] ), .A2(\a[12] ), .ZN(new_n651_));
  NOR2_X1    g00449(.A1(new_n225_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1   g00450(.A1(\a[12] ), .A2(\a[14] ), .ZN(new_n653_));
  INV_X1     g00451(.I(new_n653_), .ZN(new_n654_));
  NAND2_X1   g00452(.A1(\a[3] ), .A2(\a[14] ), .ZN(new_n655_));
  NAND4_X1   g00453(.A1(\a[2] ), .A2(\a[3] ), .A3(\a[11] ), .A4(\a[12] ), .ZN(new_n659_));
  NOR2_X1    g00454(.A1(new_n307_), .A2(new_n566_), .ZN(new_n660_));
  NAND2_X1   g00455(.A1(new_n597_), .A2(new_n211_), .ZN(new_n661_));
  NAND2_X1   g00456(.A1(new_n229_), .A2(new_n525_), .ZN(new_n662_));
  NAND2_X1   g00457(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  XOR2_X1    g00458(.A1(new_n663_), .A2(new_n659_), .Z(new_n664_));
  INV_X1     g00459(.I(new_n664_), .ZN(new_n665_));
  AOI21_X1   g00460(.A1(new_n661_), .A2(new_n662_), .B(new_n659_), .ZN(new_n666_));
  INV_X1     g00461(.I(new_n666_), .ZN(new_n667_));
  NAND3_X1   g00462(.A1(new_n661_), .A2(new_n662_), .A3(new_n659_), .ZN(new_n668_));
  AOI21_X1   g00463(.A1(new_n667_), .A2(new_n668_), .B(new_n649_), .ZN(new_n669_));
  AOI21_X1   g00464(.A1(new_n649_), .A2(new_n665_), .B(new_n669_), .ZN(new_n670_));
  NAND2_X1   g00465(.A1(new_n646_), .A2(new_n644_), .ZN(new_n671_));
  AOI21_X1   g00466(.A1(new_n670_), .A2(new_n671_), .B(new_n647_), .ZN(new_n672_));
  AOI21_X1   g00467(.A1(new_n638_), .A2(new_n639_), .B(new_n630_), .ZN(new_n673_));
  NOR2_X1    g00468(.A1(new_n673_), .A2(new_n640_), .ZN(new_n674_));
  INV_X1     g00469(.I(\a[11] ), .ZN(new_n675_));
  NAND4_X1   g00470(.A1(\a[1] ), .A2(\a[6] ), .A3(\a[8] ), .A4(\a[13] ), .ZN(new_n676_));
  AND3_X2    g00471(.A1(\a[1] ), .A2(\a[8] ), .A3(\a[14] ), .Z(new_n677_));
  AOI21_X1   g00472(.A1(\a[1] ), .A2(\a[14] ), .B(\a[8] ), .ZN(new_n678_));
  NOR2_X1    g00473(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NOR3_X1    g00474(.A1(new_n679_), .A2(\a[4] ), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1   g00475(.A1(\a[1] ), .A2(\a[14] ), .ZN(new_n681_));
  NOR4_X1    g00476(.A1(new_n633_), .A2(new_n681_), .A3(new_n242_), .A4(new_n359_), .ZN(new_n682_));
  NOR2_X1    g00477(.A1(new_n682_), .A2(new_n282_), .ZN(new_n683_));
  OAI21_X1   g00478(.A1(new_n680_), .A2(new_n683_), .B(new_n675_), .ZN(new_n684_));
  NAND2_X1   g00479(.A1(new_n682_), .A2(new_n282_), .ZN(new_n685_));
  OAI21_X1   g00480(.A1(new_n679_), .A2(new_n676_), .B(\a[4] ), .ZN(new_n686_));
  NAND3_X1   g00481(.A1(new_n686_), .A2(\a[11] ), .A3(new_n685_), .ZN(new_n687_));
  NAND2_X1   g00482(.A1(\a[6] ), .A2(\a[9] ), .ZN(new_n688_));
  NOR3_X1    g00483(.A1(new_n392_), .A2(new_n688_), .A3(\a[2] ), .ZN(new_n689_));
  AND2_X2    g00484(.A1(\a[6] ), .A2(\a[9] ), .Z(new_n690_));
  AOI21_X1   g00485(.A1(new_n609_), .A2(new_n690_), .B(new_n201_), .ZN(new_n691_));
  OAI21_X1   g00486(.A1(new_n691_), .A2(new_n689_), .B(new_n599_), .ZN(new_n692_));
  NAND3_X1   g00487(.A1(new_n609_), .A2(new_n690_), .A3(new_n201_), .ZN(new_n693_));
  OAI21_X1   g00488(.A1(new_n392_), .A2(new_n688_), .B(\a[2] ), .ZN(new_n694_));
  NAND3_X1   g00489(.A1(new_n693_), .A2(\a[13] ), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1   g00490(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1   g00491(.A1(new_n684_), .A2(new_n696_), .A3(new_n687_), .ZN(new_n697_));
  AOI21_X1   g00492(.A1(new_n686_), .A2(new_n685_), .B(\a[11] ), .ZN(new_n698_));
  NOR3_X1    g00493(.A1(new_n680_), .A2(new_n675_), .A3(new_n683_), .ZN(new_n699_));
  AOI21_X1   g00494(.A1(new_n693_), .A2(new_n694_), .B(\a[13] ), .ZN(new_n700_));
  NOR3_X1    g00495(.A1(new_n691_), .A2(new_n599_), .A3(new_n689_), .ZN(new_n701_));
  NOR2_X1    g00496(.A1(new_n701_), .A2(new_n700_), .ZN(new_n702_));
  OAI21_X1   g00497(.A1(new_n698_), .A2(new_n699_), .B(new_n702_), .ZN(new_n703_));
  AOI21_X1   g00498(.A1(new_n703_), .A2(new_n697_), .B(new_n674_), .ZN(new_n704_));
  NAND2_X1   g00499(.A1(new_n634_), .A2(new_n632_), .ZN(new_n705_));
  OAI21_X1   g00500(.A1(new_n630_), .A2(new_n635_), .B(new_n705_), .ZN(new_n706_));
  OAI21_X1   g00501(.A1(new_n698_), .A2(new_n699_), .B(new_n696_), .ZN(new_n707_));
  NAND3_X1   g00502(.A1(new_n684_), .A2(new_n702_), .A3(new_n687_), .ZN(new_n708_));
  AOI21_X1   g00503(.A1(new_n707_), .A2(new_n708_), .B(new_n706_), .ZN(new_n709_));
  NOR2_X1    g00504(.A1(new_n704_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1     g00505(.I(new_n710_), .ZN(new_n711_));
  NAND3_X1   g00506(.A1(new_n569_), .A2(new_n509_), .A3(new_n564_), .ZN(new_n712_));
  NAND2_X1   g00507(.A1(new_n567_), .A2(new_n565_), .ZN(new_n713_));
  AOI21_X1   g00508(.A1(new_n713_), .A2(new_n712_), .B(new_n566_), .ZN(new_n714_));
  NOR2_X1    g00509(.A1(new_n648_), .A2(new_n563_), .ZN(new_n715_));
  OAI21_X1   g00510(.A1(new_n714_), .A2(new_n715_), .B(new_n668_), .ZN(new_n716_));
  NAND2_X1   g00511(.A1(new_n716_), .A2(new_n667_), .ZN(new_n717_));
  AOI21_X1   g00512(.A1(new_n218_), .A2(new_n654_), .B(new_n652_), .ZN(new_n718_));
  NAND3_X1   g00513(.A1(\a[10] ), .A2(\a[12] ), .A3(\a[15] ), .ZN(new_n719_));
  NAND2_X1   g00514(.A1(new_n719_), .A2(new_n214_), .ZN(new_n720_));
  NOR2_X1    g00515(.A1(\a[5] ), .A2(\a[10] ), .ZN(new_n721_));
  NAND4_X1   g00516(.A1(\a[0] ), .A2(\a[3] ), .A3(\a[12] ), .A4(\a[15] ), .ZN(new_n722_));
  NOR2_X1    g00517(.A1(new_n722_), .A2(new_n721_), .ZN(new_n723_));
  NAND2_X1   g00518(.A1(new_n723_), .A2(new_n720_), .ZN(new_n724_));
  NAND3_X1   g00519(.A1(new_n719_), .A2(new_n214_), .A3(\a[5] ), .ZN(new_n725_));
  AOI22_X1   g00520(.A1(\a[0] ), .A2(\a[3] ), .B1(\a[12] ), .B2(\a[15] ), .ZN(new_n726_));
  NAND3_X1   g00521(.A1(new_n725_), .A2(new_n722_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1   g00522(.A1(new_n727_), .A2(new_n724_), .ZN(new_n728_));
  AOI21_X1   g00523(.A1(new_n660_), .A2(new_n597_), .B(new_n229_), .ZN(new_n729_));
  NOR2_X1    g00524(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1     g00525(.I(new_n729_), .ZN(new_n731_));
  AOI21_X1   g00526(.A1(new_n724_), .A2(new_n727_), .B(new_n731_), .ZN(new_n732_));
  OAI21_X1   g00527(.A1(new_n730_), .A2(new_n732_), .B(new_n718_), .ZN(new_n733_));
  INV_X1     g00528(.I(new_n718_), .ZN(new_n734_));
  AOI21_X1   g00529(.A1(new_n727_), .A2(new_n724_), .B(new_n729_), .ZN(new_n735_));
  NAND3_X1   g00530(.A1(new_n727_), .A2(new_n724_), .A3(new_n729_), .ZN(new_n736_));
  INV_X1     g00531(.I(new_n736_), .ZN(new_n737_));
  OAI21_X1   g00532(.A1(new_n737_), .A2(new_n735_), .B(new_n734_), .ZN(new_n738_));
  AOI21_X1   g00533(.A1(new_n733_), .A2(new_n738_), .B(new_n717_), .ZN(new_n739_));
  AOI21_X1   g00534(.A1(new_n649_), .A2(new_n668_), .B(new_n666_), .ZN(new_n740_));
  NAND3_X1   g00535(.A1(new_n731_), .A2(new_n727_), .A3(new_n724_), .ZN(new_n741_));
  NAND2_X1   g00536(.A1(new_n728_), .A2(new_n729_), .ZN(new_n742_));
  AOI21_X1   g00537(.A1(new_n742_), .A2(new_n741_), .B(new_n734_), .ZN(new_n743_));
  INV_X1     g00538(.I(new_n720_), .ZN(new_n744_));
  NOR3_X1    g00539(.A1(new_n744_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n745_));
  INV_X1     g00540(.I(new_n727_), .ZN(new_n746_));
  OAI21_X1   g00541(.A1(new_n746_), .A2(new_n745_), .B(new_n731_), .ZN(new_n747_));
  AOI21_X1   g00542(.A1(new_n747_), .A2(new_n736_), .B(new_n718_), .ZN(new_n748_));
  NOR3_X1    g00543(.A1(new_n743_), .A2(new_n748_), .A3(new_n740_), .ZN(new_n749_));
  OAI22_X1   g00544(.A1(new_n739_), .A2(new_n749_), .B1(new_n704_), .B2(new_n709_), .ZN(new_n750_));
  AOI21_X1   g00545(.A1(new_n733_), .A2(new_n738_), .B(new_n740_), .ZN(new_n751_));
  NOR3_X1    g00546(.A1(new_n743_), .A2(new_n748_), .A3(new_n717_), .ZN(new_n752_));
  NOR2_X1    g00547(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1   g00548(.A1(new_n711_), .A2(new_n753_), .B(new_n750_), .ZN(new_n754_));
  XOR2_X1    g00549(.A1(new_n672_), .A2(new_n754_), .Z(new_n755_));
  INV_X1     g00550(.I(new_n672_), .ZN(new_n756_));
  NAND2_X1   g00551(.A1(new_n756_), .A2(new_n754_), .ZN(new_n757_));
  INV_X1     g00552(.I(new_n754_), .ZN(new_n758_));
  NAND2_X1   g00553(.A1(new_n758_), .A2(new_n672_), .ZN(new_n759_));
  NAND2_X1   g00554(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1   g00555(.A1(new_n628_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1   g00556(.A1(new_n628_), .A2(new_n755_), .B(new_n761_), .ZN(\asquared[16] ));
  NAND2_X1   g00557(.A1(\asquared[15] ), .A2(new_n759_), .ZN(new_n763_));
  NAND2_X1   g00558(.A1(new_n763_), .A2(new_n757_), .ZN(new_n764_));
  INV_X1     g00559(.I(new_n751_), .ZN(new_n765_));
  OAI21_X1   g00560(.A1(new_n711_), .A2(new_n752_), .B(new_n765_), .ZN(new_n766_));
  INV_X1     g00561(.I(new_n681_), .ZN(new_n767_));
  NOR2_X1    g00562(.A1(new_n392_), .A2(new_n688_), .ZN(new_n768_));
  NAND2_X1   g00563(.A1(\a[2] ), .A2(\a[13] ), .ZN(new_n769_));
  AOI21_X1   g00564(.A1(new_n392_), .A2(new_n688_), .B(new_n769_), .ZN(new_n770_));
  NOR2_X1    g00565(.A1(new_n770_), .A2(new_n768_), .ZN(new_n771_));
  NAND2_X1   g00566(.A1(\a[7] ), .A2(\a[9] ), .ZN(new_n772_));
  NAND2_X1   g00567(.A1(\a[1] ), .A2(\a[15] ), .ZN(new_n773_));
  XNOR2_X1   g00568(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NOR3_X1    g00569(.A1(new_n774_), .A2(new_n767_), .A3(new_n771_), .ZN(new_n775_));
  INV_X1     g00570(.I(new_n775_), .ZN(new_n776_));
  OAI21_X1   g00571(.A1(new_n774_), .A2(new_n771_), .B(new_n767_), .ZN(new_n777_));
  AOI21_X1   g00572(.A1(new_n776_), .A2(new_n777_), .B(\a[8] ), .ZN(new_n778_));
  INV_X1     g00573(.I(new_n777_), .ZN(new_n779_));
  NOR3_X1    g00574(.A1(new_n779_), .A2(new_n359_), .A3(new_n775_), .ZN(new_n780_));
  NOR2_X1    g00575(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1   g00576(.A1(new_n728_), .A2(new_n729_), .B(new_n734_), .ZN(new_n782_));
  NAND3_X1   g00577(.A1(\a[12] ), .A2(\a[13] ), .A3(\a[14] ), .ZN(new_n783_));
  NAND3_X1   g00578(.A1(\a[2] ), .A2(\a[3] ), .A3(\a[4] ), .ZN(new_n784_));
  NAND2_X1   g00579(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1   g00580(.A1(\a[13] ), .A2(\a[14] ), .ZN(new_n786_));
  INV_X1     g00581(.I(new_n786_), .ZN(new_n787_));
  NAND2_X1   g00582(.A1(\a[4] ), .A2(\a[12] ), .ZN(new_n788_));
  NOR4_X1    g00583(.A1(new_n785_), .A2(new_n232_), .A3(new_n787_), .A4(new_n788_), .ZN(new_n789_));
  OAI21_X1   g00584(.A1(new_n782_), .A2(new_n730_), .B(new_n789_), .ZN(new_n790_));
  NAND2_X1   g00585(.A1(new_n742_), .A2(new_n718_), .ZN(new_n791_));
  INV_X1     g00586(.I(new_n789_), .ZN(new_n792_));
  NAND3_X1   g00587(.A1(new_n791_), .A2(new_n741_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1   g00588(.A1(new_n793_), .A2(new_n790_), .ZN(new_n794_));
  NAND2_X1   g00589(.A1(new_n708_), .A2(new_n706_), .ZN(new_n795_));
  NAND2_X1   g00590(.A1(\a[10] ), .A2(\a[11] ), .ZN(new_n796_));
  INV_X1     g00591(.I(new_n796_), .ZN(new_n797_));
  NAND2_X1   g00592(.A1(\a[6] ), .A2(\a[16] ), .ZN(new_n798_));
  NOR2_X1    g00593(.A1(new_n395_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1     g00594(.I(\a[16] ), .ZN(new_n800_));
  NAND4_X1   g00595(.A1(\a[0] ), .A2(\a[6] ), .A3(\a[10] ), .A4(\a[16] ), .ZN(new_n805_));
  INV_X1     g00596(.I(new_n805_), .ZN(new_n806_));
  NAND2_X1   g00597(.A1(new_n725_), .A2(new_n722_), .ZN(new_n807_));
  NAND3_X1   g00598(.A1(\a[1] ), .A2(\a[8] ), .A3(\a[14] ), .ZN(new_n808_));
  NAND2_X1   g00599(.A1(new_n681_), .A2(new_n359_), .ZN(new_n809_));
  NAND3_X1   g00600(.A1(new_n809_), .A2(new_n676_), .A3(new_n808_), .ZN(new_n810_));
  NAND2_X1   g00601(.A1(\a[4] ), .A2(\a[11] ), .ZN(new_n811_));
  INV_X1     g00602(.I(new_n811_), .ZN(new_n812_));
  AOI21_X1   g00603(.A1(new_n810_), .A2(new_n812_), .B(new_n682_), .ZN(new_n813_));
  NOR2_X1    g00604(.A1(new_n813_), .A2(new_n807_), .ZN(new_n814_));
  INV_X1     g00605(.I(new_n807_), .ZN(new_n815_));
  AOI21_X1   g00606(.A1(new_n679_), .A2(new_n676_), .B(new_n811_), .ZN(new_n816_));
  NOR3_X1    g00607(.A1(new_n815_), .A2(new_n816_), .A3(new_n682_), .ZN(new_n817_));
  OAI21_X1   g00608(.A1(new_n817_), .A2(new_n814_), .B(new_n806_), .ZN(new_n818_));
  NOR3_X1    g00609(.A1(new_n816_), .A2(new_n682_), .A3(new_n807_), .ZN(new_n819_));
  NOR2_X1    g00610(.A1(new_n813_), .A2(new_n815_), .ZN(new_n820_));
  OAI21_X1   g00611(.A1(new_n820_), .A2(new_n819_), .B(new_n805_), .ZN(new_n821_));
  NAND2_X1   g00612(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1   g00613(.A1(new_n822_), .A2(new_n795_), .A3(new_n707_), .ZN(new_n823_));
  NOR3_X1    g00614(.A1(new_n699_), .A2(new_n696_), .A3(new_n698_), .ZN(new_n824_));
  OAI21_X1   g00615(.A1(new_n674_), .A2(new_n824_), .B(new_n707_), .ZN(new_n825_));
  OAI21_X1   g00616(.A1(new_n682_), .A2(new_n816_), .B(new_n815_), .ZN(new_n826_));
  NAND2_X1   g00617(.A1(new_n813_), .A2(new_n807_), .ZN(new_n827_));
  AOI21_X1   g00618(.A1(new_n826_), .A2(new_n827_), .B(new_n805_), .ZN(new_n828_));
  NAND2_X1   g00619(.A1(new_n813_), .A2(new_n815_), .ZN(new_n829_));
  OAI21_X1   g00620(.A1(new_n816_), .A2(new_n682_), .B(new_n807_), .ZN(new_n830_));
  AOI21_X1   g00621(.A1(new_n829_), .A2(new_n830_), .B(new_n806_), .ZN(new_n831_));
  NOR2_X1    g00622(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1   g00623(.A1(new_n825_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1   g00624(.A1(new_n833_), .A2(new_n823_), .B(new_n794_), .ZN(new_n834_));
  INV_X1     g00625(.I(new_n790_), .ZN(new_n835_));
  NOR3_X1    g00626(.A1(new_n782_), .A2(new_n730_), .A3(new_n789_), .ZN(new_n836_));
  NOR2_X1    g00627(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1     g00628(.I(new_n707_), .ZN(new_n838_));
  NOR2_X1    g00629(.A1(new_n824_), .A2(new_n674_), .ZN(new_n839_));
  NOR3_X1    g00630(.A1(new_n832_), .A2(new_n839_), .A3(new_n838_), .ZN(new_n840_));
  AOI21_X1   g00631(.A1(new_n707_), .A2(new_n795_), .B(new_n822_), .ZN(new_n841_));
  NOR3_X1    g00632(.A1(new_n841_), .A2(new_n840_), .A3(new_n837_), .ZN(new_n842_));
  OAI21_X1   g00633(.A1(new_n842_), .A2(new_n834_), .B(new_n781_), .ZN(new_n843_));
  INV_X1     g00634(.I(new_n781_), .ZN(new_n844_));
  OAI21_X1   g00635(.A1(new_n841_), .A2(new_n840_), .B(new_n837_), .ZN(new_n845_));
  NAND3_X1   g00636(.A1(new_n833_), .A2(new_n823_), .A3(new_n794_), .ZN(new_n846_));
  NAND3_X1   g00637(.A1(new_n845_), .A2(new_n846_), .A3(new_n844_), .ZN(new_n847_));
  AND2_X2    g00638(.A1(new_n843_), .A2(new_n847_), .Z(new_n848_));
  XOR2_X1    g00639(.A1(new_n848_), .A2(new_n766_), .Z(new_n849_));
  NAND2_X1   g00640(.A1(new_n764_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1   g00641(.A1(new_n843_), .A2(new_n847_), .B(new_n766_), .ZN(new_n851_));
  NAND3_X1   g00642(.A1(new_n843_), .A2(new_n847_), .A3(new_n766_), .ZN(new_n852_));
  INV_X1     g00643(.I(new_n852_), .ZN(new_n853_));
  NOR2_X1    g00644(.A1(new_n853_), .A2(new_n851_), .ZN(new_n854_));
  OAI21_X1   g00645(.A1(new_n764_), .A2(new_n854_), .B(new_n850_), .ZN(\asquared[17] ));
  NAND2_X1   g00646(.A1(new_n852_), .A2(new_n758_), .ZN(new_n856_));
  NAND4_X1   g00647(.A1(new_n843_), .A2(new_n847_), .A3(new_n754_), .A4(new_n766_), .ZN(new_n857_));
  NAND2_X1   g00648(.A1(new_n857_), .A2(new_n672_), .ZN(new_n858_));
  NAND2_X1   g00649(.A1(new_n858_), .A2(new_n856_), .ZN(new_n859_));
  NOR2_X1    g00650(.A1(new_n628_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1     g00651(.I(new_n825_), .ZN(new_n861_));
  NOR2_X1    g00652(.A1(new_n861_), .A2(new_n832_), .ZN(new_n862_));
  NAND2_X1   g00653(.A1(new_n861_), .A2(new_n832_), .ZN(new_n863_));
  NAND2_X1   g00654(.A1(new_n844_), .A2(new_n837_), .ZN(new_n864_));
  NAND2_X1   g00655(.A1(new_n794_), .A2(new_n781_), .ZN(new_n865_));
  NAND2_X1   g00656(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1   g00657(.A1(new_n866_), .A2(new_n863_), .B(new_n862_), .ZN(new_n867_));
  NAND2_X1   g00658(.A1(\a[11] ), .A2(\a[15] ), .ZN(new_n868_));
  NOR2_X1    g00659(.A1(new_n868_), .A2(new_n282_), .ZN(new_n869_));
  NAND2_X1   g00660(.A1(\a[11] ), .A2(\a[13] ), .ZN(new_n870_));
  OAI21_X1   g00661(.A1(new_n870_), .A2(new_n201_), .B(new_n242_), .ZN(new_n871_));
  NOR2_X1    g00662(.A1(new_n871_), .A2(new_n869_), .ZN(new_n872_));
  NAND2_X1   g00663(.A1(\a[13] ), .A2(\a[15] ), .ZN(new_n873_));
  NOR3_X1    g00664(.A1(new_n872_), .A2(new_n260_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1     g00665(.I(\a[15] ), .ZN(new_n875_));
  NOR3_X1    g00666(.A1(new_n260_), .A2(new_n599_), .A3(new_n875_), .ZN(new_n877_));
  INV_X1     g00667(.I(new_n877_), .ZN(new_n878_));
  NAND2_X1   g00668(.A1(\a[6] ), .A2(\a[11] ), .ZN(new_n879_));
  INV_X1     g00669(.I(new_n879_), .ZN(new_n880_));
  NAND2_X1   g00670(.A1(new_n260_), .A2(new_n873_), .ZN(new_n881_));
  AOI22_X1   g00671(.A1(new_n874_), .A2(new_n878_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1     g00672(.I(new_n882_), .ZN(new_n883_));
  NOR2_X1    g00673(.A1(new_n772_), .A2(new_n773_), .ZN(new_n884_));
  INV_X1     g00674(.I(\a[17] ), .ZN(new_n885_));
  NOR2_X1    g00675(.A1(new_n199_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1   g00676(.A1(new_n884_), .A2(new_n353_), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1   g00677(.A1(new_n884_), .A2(new_n886_), .ZN(new_n888_));
  NAND2_X1   g00678(.A1(new_n888_), .A2(\a[5] ), .ZN(new_n889_));
  AOI21_X1   g00679(.A1(new_n889_), .A2(new_n887_), .B(\a[12] ), .ZN(new_n890_));
  NAND3_X1   g00680(.A1(new_n889_), .A2(\a[12] ), .A3(new_n887_), .ZN(new_n891_));
  INV_X1     g00681(.I(new_n891_), .ZN(new_n892_));
  OAI21_X1   g00682(.A1(new_n268_), .A2(new_n461_), .B(new_n453_), .ZN(new_n893_));
  AOI21_X1   g00683(.A1(new_n893_), .A2(new_n655_), .B(new_n525_), .ZN(new_n894_));
  NAND2_X1   g00684(.A1(new_n894_), .A2(new_n392_), .ZN(new_n895_));
  INV_X1     g00685(.I(new_n895_), .ZN(new_n896_));
  NOR2_X1    g00686(.A1(new_n894_), .A2(new_n392_), .ZN(new_n897_));
  OAI22_X1   g00687(.A1(new_n892_), .A2(new_n890_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1     g00688(.I(new_n898_), .ZN(new_n899_));
  INV_X1     g00689(.I(new_n897_), .ZN(new_n900_));
  NAND2_X1   g00690(.A1(new_n900_), .A2(new_n895_), .ZN(new_n901_));
  NOR3_X1    g00691(.A1(new_n901_), .A2(new_n892_), .A3(new_n890_), .ZN(new_n902_));
  OAI21_X1   g00692(.A1(new_n899_), .A2(new_n902_), .B(new_n883_), .ZN(new_n903_));
  NOR2_X1    g00693(.A1(new_n892_), .A2(new_n890_), .ZN(new_n904_));
  XOR2_X1    g00694(.A1(new_n904_), .A2(new_n901_), .Z(new_n905_));
  OAI21_X1   g00695(.A1(new_n905_), .A2(new_n883_), .B(new_n903_), .ZN(new_n906_));
  NOR2_X1    g00696(.A1(new_n782_), .A2(new_n730_), .ZN(new_n907_));
  INV_X1     g00697(.I(new_n907_), .ZN(new_n908_));
  OAI21_X1   g00698(.A1(new_n779_), .A2(new_n775_), .B(new_n359_), .ZN(new_n909_));
  NAND3_X1   g00699(.A1(new_n776_), .A2(\a[8] ), .A3(new_n777_), .ZN(new_n910_));
  AOI21_X1   g00700(.A1(new_n909_), .A2(new_n910_), .B(new_n792_), .ZN(new_n911_));
  NAND3_X1   g00701(.A1(new_n909_), .A2(new_n910_), .A3(new_n792_), .ZN(new_n912_));
  AOI21_X1   g00702(.A1(new_n908_), .A2(new_n912_), .B(new_n911_), .ZN(new_n913_));
  AOI21_X1   g00703(.A1(new_n806_), .A2(new_n827_), .B(new_n814_), .ZN(new_n914_));
  INV_X1     g00704(.I(new_n914_), .ZN(new_n915_));
  AOI21_X1   g00705(.A1(new_n608_), .A2(new_n797_), .B(new_n799_), .ZN(new_n916_));
  AOI22_X1   g00706(.A1(new_n232_), .A2(new_n787_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n917_));
  NAND2_X1   g00707(.A1(\a[1] ), .A2(\a[16] ), .ZN(new_n918_));
  XOR2_X1    g00708(.A1(new_n918_), .A2(\a[9] ), .Z(new_n919_));
  NOR2_X1    g00709(.A1(new_n919_), .A2(new_n917_), .ZN(new_n920_));
  NAND2_X1   g00710(.A1(new_n919_), .A2(new_n917_), .ZN(new_n921_));
  INV_X1     g00711(.I(new_n921_), .ZN(new_n922_));
  OAI21_X1   g00712(.A1(new_n922_), .A2(new_n920_), .B(new_n916_), .ZN(new_n923_));
  INV_X1     g00713(.I(new_n916_), .ZN(new_n924_));
  INV_X1     g00714(.I(new_n917_), .ZN(new_n925_));
  NOR2_X1    g00715(.A1(new_n925_), .A2(new_n919_), .ZN(new_n926_));
  XOR2_X1    g00716(.A1(new_n918_), .A2(new_n364_), .Z(new_n927_));
  NOR2_X1    g00717(.A1(new_n927_), .A2(new_n917_), .ZN(new_n928_));
  OAI21_X1   g00718(.A1(new_n926_), .A2(new_n928_), .B(new_n924_), .ZN(new_n929_));
  NOR2_X1    g00719(.A1(new_n774_), .A2(new_n771_), .ZN(new_n930_));
  AOI21_X1   g00720(.A1(new_n774_), .A2(new_n771_), .B(new_n808_), .ZN(new_n931_));
  NOR2_X1    g00721(.A1(new_n931_), .A2(new_n930_), .ZN(new_n932_));
  INV_X1     g00722(.I(new_n932_), .ZN(new_n933_));
  NAND3_X1   g00723(.A1(new_n933_), .A2(new_n923_), .A3(new_n929_), .ZN(new_n934_));
  INV_X1     g00724(.I(new_n934_), .ZN(new_n935_));
  AOI21_X1   g00725(.A1(new_n923_), .A2(new_n929_), .B(new_n933_), .ZN(new_n936_));
  OAI21_X1   g00726(.A1(new_n935_), .A2(new_n936_), .B(new_n915_), .ZN(new_n937_));
  AOI21_X1   g00727(.A1(new_n923_), .A2(new_n929_), .B(new_n932_), .ZN(new_n938_));
  NAND3_X1   g00728(.A1(new_n923_), .A2(new_n929_), .A3(new_n932_), .ZN(new_n939_));
  INV_X1     g00729(.I(new_n939_), .ZN(new_n940_));
  OAI21_X1   g00730(.A1(new_n940_), .A2(new_n938_), .B(new_n914_), .ZN(new_n941_));
  AOI21_X1   g00731(.A1(new_n937_), .A2(new_n941_), .B(new_n913_), .ZN(new_n942_));
  OAI21_X1   g00732(.A1(new_n778_), .A2(new_n780_), .B(new_n789_), .ZN(new_n943_));
  NOR3_X1    g00733(.A1(new_n778_), .A2(new_n780_), .A3(new_n789_), .ZN(new_n944_));
  OAI21_X1   g00734(.A1(new_n907_), .A2(new_n944_), .B(new_n943_), .ZN(new_n945_));
  NAND2_X1   g00735(.A1(new_n923_), .A2(new_n929_), .ZN(new_n946_));
  NAND2_X1   g00736(.A1(new_n946_), .A2(new_n932_), .ZN(new_n947_));
  AOI21_X1   g00737(.A1(new_n947_), .A2(new_n934_), .B(new_n914_), .ZN(new_n948_));
  INV_X1     g00738(.I(new_n938_), .ZN(new_n949_));
  AOI21_X1   g00739(.A1(new_n949_), .A2(new_n939_), .B(new_n915_), .ZN(new_n950_));
  NOR3_X1    g00740(.A1(new_n945_), .A2(new_n950_), .A3(new_n948_), .ZN(new_n951_));
  OAI21_X1   g00741(.A1(new_n942_), .A2(new_n951_), .B(new_n906_), .ZN(new_n952_));
  INV_X1     g00742(.I(new_n902_), .ZN(new_n953_));
  AOI21_X1   g00743(.A1(new_n953_), .A2(new_n898_), .B(new_n882_), .ZN(new_n954_));
  NOR2_X1    g00744(.A1(new_n896_), .A2(new_n897_), .ZN(new_n955_));
  XOR2_X1    g00745(.A1(new_n904_), .A2(new_n955_), .Z(new_n956_));
  AOI21_X1   g00746(.A1(new_n956_), .A2(new_n882_), .B(new_n954_), .ZN(new_n957_));
  AOI21_X1   g00747(.A1(new_n937_), .A2(new_n941_), .B(new_n945_), .ZN(new_n958_));
  NOR3_X1    g00748(.A1(new_n913_), .A2(new_n950_), .A3(new_n948_), .ZN(new_n959_));
  OAI21_X1   g00749(.A1(new_n958_), .A2(new_n959_), .B(new_n957_), .ZN(new_n960_));
  AOI21_X1   g00750(.A1(new_n960_), .A2(new_n952_), .B(new_n867_), .ZN(new_n961_));
  XOR2_X1    g00751(.A1(new_n860_), .A2(new_n961_), .Z(new_n962_));
  XOR2_X1    g00752(.A1(new_n962_), .A2(new_n851_), .Z(\asquared[18] ));
  NAND3_X1   g00753(.A1(new_n960_), .A2(new_n952_), .A3(new_n867_), .ZN(new_n964_));
  NAND2_X1   g00754(.A1(new_n964_), .A2(new_n851_), .ZN(new_n965_));
  NOR3_X1    g00755(.A1(new_n628_), .A2(new_n859_), .A3(new_n965_), .ZN(new_n966_));
  NOR2_X1    g00756(.A1(new_n966_), .A2(new_n961_), .ZN(new_n967_));
  INV_X1     g00757(.I(new_n890_), .ZN(new_n968_));
  NAND2_X1   g00758(.A1(new_n968_), .A2(new_n891_), .ZN(new_n969_));
  OAI21_X1   g00759(.A1(new_n969_), .A2(new_n901_), .B(new_n883_), .ZN(new_n970_));
  NAND2_X1   g00760(.A1(\a[5] ), .A2(\a[12] ), .ZN(new_n971_));
  INV_X1     g00761(.I(new_n971_), .ZN(new_n972_));
  OAI21_X1   g00762(.A1(new_n884_), .A2(new_n886_), .B(new_n972_), .ZN(new_n973_));
  NAND2_X1   g00763(.A1(new_n973_), .A2(new_n888_), .ZN(new_n974_));
  INV_X1     g00764(.I(new_n974_), .ZN(new_n975_));
  OAI22_X1   g00765(.A1(new_n893_), .A2(new_n392_), .B1(new_n525_), .B2(new_n655_), .ZN(new_n976_));
  NAND2_X1   g00766(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  INV_X1     g00767(.I(new_n976_), .ZN(new_n978_));
  NAND2_X1   g00768(.A1(new_n978_), .A2(new_n974_), .ZN(new_n979_));
  AOI21_X1   g00769(.A1(new_n977_), .A2(new_n979_), .B(new_n877_), .ZN(new_n980_));
  NAND2_X1   g00770(.A1(new_n974_), .A2(new_n976_), .ZN(new_n981_));
  NOR2_X1    g00771(.A1(new_n974_), .A2(new_n976_), .ZN(new_n982_));
  INV_X1     g00772(.I(new_n982_), .ZN(new_n983_));
  AOI21_X1   g00773(.A1(new_n983_), .A2(new_n981_), .B(new_n878_), .ZN(new_n984_));
  OAI21_X1   g00774(.A1(new_n924_), .A2(new_n920_), .B(new_n921_), .ZN(new_n985_));
  OAI21_X1   g00775(.A1(new_n984_), .A2(new_n980_), .B(new_n985_), .ZN(new_n986_));
  NOR2_X1    g00776(.A1(new_n978_), .A2(new_n974_), .ZN(new_n987_));
  NOR2_X1    g00777(.A1(new_n975_), .A2(new_n976_), .ZN(new_n988_));
  OAI21_X1   g00778(.A1(new_n988_), .A2(new_n987_), .B(new_n878_), .ZN(new_n989_));
  INV_X1     g00779(.I(new_n981_), .ZN(new_n990_));
  OAI21_X1   g00780(.A1(new_n990_), .A2(new_n982_), .B(new_n877_), .ZN(new_n991_));
  INV_X1     g00781(.I(new_n985_), .ZN(new_n992_));
  NAND3_X1   g00782(.A1(new_n989_), .A2(new_n991_), .A3(new_n992_), .ZN(new_n993_));
  AOI22_X1   g00783(.A1(new_n986_), .A2(new_n993_), .B1(new_n898_), .B2(new_n970_), .ZN(new_n994_));
  OAI21_X1   g00784(.A1(new_n902_), .A2(new_n882_), .B(new_n898_), .ZN(new_n995_));
  NAND3_X1   g00785(.A1(new_n989_), .A2(new_n991_), .A3(new_n985_), .ZN(new_n996_));
  OAI21_X1   g00786(.A1(new_n984_), .A2(new_n980_), .B(new_n992_), .ZN(new_n997_));
  AOI21_X1   g00787(.A1(new_n996_), .A2(new_n997_), .B(new_n995_), .ZN(new_n998_));
  NOR2_X1    g00788(.A1(new_n998_), .A2(new_n994_), .ZN(new_n999_));
  NAND2_X1   g00789(.A1(\a[5] ), .A2(\a[7] ), .ZN(new_n1000_));
  INV_X1     g00790(.I(new_n870_), .ZN(new_n1001_));
  NAND2_X1   g00791(.A1(\a[13] ), .A2(\a[18] ), .ZN(new_n1002_));
  NOR2_X1    g00792(.A1(new_n263_), .A2(new_n1002_), .ZN(new_n1003_));
  NAND2_X1   g00793(.A1(\a[7] ), .A2(\a[18] ), .ZN(new_n1004_));
  NOR2_X1    g00794(.A1(new_n483_), .A2(new_n1004_), .ZN(new_n1005_));
  AOI21_X1   g00795(.A1(new_n1003_), .A2(new_n1005_), .B(new_n1001_), .ZN(new_n1006_));
  NOR2_X1    g00796(.A1(new_n1006_), .A2(new_n1000_), .ZN(new_n1007_));
  INV_X1     g00797(.I(new_n1007_), .ZN(new_n1008_));
  NOR2_X1    g00798(.A1(new_n268_), .A2(new_n675_), .ZN(new_n1009_));
  NOR2_X1    g00799(.A1(new_n1007_), .A2(new_n1003_), .ZN(new_n1010_));
  INV_X1     g00800(.I(new_n263_), .ZN(new_n1011_));
  INV_X1     g00801(.I(new_n1002_), .ZN(new_n1012_));
  NOR2_X1    g00802(.A1(new_n1011_), .A2(new_n1012_), .ZN(new_n1013_));
  AOI22_X1   g00803(.A1(new_n1010_), .A2(new_n1013_), .B1(new_n1008_), .B2(new_n1009_), .ZN(new_n1014_));
  INV_X1     g00804(.I(new_n1014_), .ZN(new_n1015_));
  INV_X1     g00805(.I(new_n784_), .ZN(new_n1016_));
  NAND2_X1   g00806(.A1(\a[14] ), .A2(\a[16] ), .ZN(new_n1017_));
  NAND2_X1   g00807(.A1(\a[14] ), .A2(\a[15] ), .ZN(new_n1018_));
  NOR2_X1    g00808(.A1(new_n1017_), .A2(new_n1018_), .ZN(new_n1019_));
  NOR2_X1    g00809(.A1(new_n1019_), .A2(new_n1016_), .ZN(new_n1020_));
  NAND2_X1   g00810(.A1(\a[15] ), .A2(\a[16] ), .ZN(new_n1021_));
  NOR2_X1    g00811(.A1(new_n225_), .A2(new_n1021_), .ZN(new_n1022_));
  NOR2_X1    g00812(.A1(new_n282_), .A2(new_n650_), .ZN(new_n1023_));
  INV_X1     g00813(.I(new_n1023_), .ZN(new_n1024_));
  NOR2_X1    g00814(.A1(new_n201_), .A2(new_n800_), .ZN(new_n1025_));
  AOI21_X1   g00815(.A1(\a[3] ), .A2(\a[15] ), .B(new_n1025_), .ZN(new_n1026_));
  NOR3_X1    g00816(.A1(new_n1026_), .A2(new_n1022_), .A3(new_n1024_), .ZN(new_n1027_));
  AND2_X2    g00817(.A1(new_n1027_), .A2(new_n1020_), .Z(new_n1028_));
  NOR2_X1    g00818(.A1(new_n364_), .A2(new_n800_), .ZN(new_n1029_));
  NAND2_X1   g00819(.A1(new_n1029_), .A2(\a[1] ), .ZN(new_n1030_));
  OAI21_X1   g00820(.A1(new_n194_), .A2(new_n885_), .B(new_n391_), .ZN(new_n1031_));
  INV_X1     g00821(.I(new_n1031_), .ZN(new_n1032_));
  NOR3_X1    g00822(.A1(new_n391_), .A2(new_n194_), .A3(new_n885_), .ZN(new_n1033_));
  NOR2_X1    g00823(.A1(new_n1032_), .A2(new_n1033_), .ZN(new_n1034_));
  NOR2_X1    g00824(.A1(new_n1034_), .A2(new_n1030_), .ZN(new_n1035_));
  NAND2_X1   g00825(.A1(new_n1035_), .A2(new_n242_), .ZN(new_n1036_));
  INV_X1     g00826(.I(new_n1030_), .ZN(new_n1037_));
  INV_X1     g00827(.I(new_n1033_), .ZN(new_n1038_));
  NAND2_X1   g00828(.A1(new_n1038_), .A2(new_n1031_), .ZN(new_n1039_));
  NAND2_X1   g00829(.A1(new_n1039_), .A2(new_n1037_), .ZN(new_n1040_));
  NAND2_X1   g00830(.A1(new_n1040_), .A2(\a[6] ), .ZN(new_n1041_));
  AOI21_X1   g00831(.A1(new_n1036_), .A2(new_n1041_), .B(\a[12] ), .ZN(new_n1042_));
  NOR2_X1    g00832(.A1(new_n1040_), .A2(\a[6] ), .ZN(new_n1043_));
  NOR2_X1    g00833(.A1(new_n1035_), .A2(new_n242_), .ZN(new_n1044_));
  NOR3_X1    g00834(.A1(new_n1044_), .A2(new_n566_), .A3(new_n1043_), .ZN(new_n1045_));
  OAI21_X1   g00835(.A1(new_n1045_), .A2(new_n1042_), .B(new_n1028_), .ZN(new_n1046_));
  INV_X1     g00836(.I(new_n1028_), .ZN(new_n1047_));
  OAI21_X1   g00837(.A1(new_n1044_), .A2(new_n1043_), .B(new_n566_), .ZN(new_n1048_));
  NAND3_X1   g00838(.A1(new_n1036_), .A2(\a[12] ), .A3(new_n1041_), .ZN(new_n1049_));
  NAND3_X1   g00839(.A1(new_n1048_), .A2(new_n1049_), .A3(new_n1047_), .ZN(new_n1050_));
  AOI21_X1   g00840(.A1(new_n1046_), .A2(new_n1050_), .B(new_n1015_), .ZN(new_n1051_));
  OAI21_X1   g00841(.A1(new_n1045_), .A2(new_n1042_), .B(new_n1047_), .ZN(new_n1052_));
  NAND3_X1   g00842(.A1(new_n1048_), .A2(new_n1049_), .A3(new_n1028_), .ZN(new_n1053_));
  AOI21_X1   g00843(.A1(new_n1052_), .A2(new_n1053_), .B(new_n1014_), .ZN(new_n1054_));
  AOI21_X1   g00844(.A1(new_n915_), .A2(new_n939_), .B(new_n938_), .ZN(new_n1055_));
  INV_X1     g00845(.I(new_n1055_), .ZN(new_n1056_));
  OAI21_X1   g00846(.A1(new_n1051_), .A2(new_n1054_), .B(new_n1056_), .ZN(new_n1057_));
  AOI21_X1   g00847(.A1(new_n1048_), .A2(new_n1049_), .B(new_n1047_), .ZN(new_n1058_));
  NOR3_X1    g00848(.A1(new_n1045_), .A2(new_n1042_), .A3(new_n1028_), .ZN(new_n1059_));
  OAI21_X1   g00849(.A1(new_n1059_), .A2(new_n1058_), .B(new_n1014_), .ZN(new_n1060_));
  AOI21_X1   g00850(.A1(new_n1048_), .A2(new_n1049_), .B(new_n1028_), .ZN(new_n1061_));
  NOR3_X1    g00851(.A1(new_n1045_), .A2(new_n1042_), .A3(new_n1047_), .ZN(new_n1062_));
  OAI21_X1   g00852(.A1(new_n1062_), .A2(new_n1061_), .B(new_n1015_), .ZN(new_n1063_));
  NAND3_X1   g00853(.A1(new_n1060_), .A2(new_n1063_), .A3(new_n1055_), .ZN(new_n1064_));
  AOI21_X1   g00854(.A1(new_n1057_), .A2(new_n1064_), .B(new_n999_), .ZN(new_n1065_));
  NAND2_X1   g00855(.A1(new_n986_), .A2(new_n993_), .ZN(new_n1066_));
  NAND2_X1   g00856(.A1(new_n1066_), .A2(new_n995_), .ZN(new_n1067_));
  AOI21_X1   g00857(.A1(new_n904_), .A2(new_n955_), .B(new_n882_), .ZN(new_n1068_));
  NOR2_X1    g00858(.A1(new_n899_), .A2(new_n1068_), .ZN(new_n1069_));
  NOR3_X1    g00859(.A1(new_n984_), .A2(new_n980_), .A3(new_n992_), .ZN(new_n1070_));
  AOI21_X1   g00860(.A1(new_n989_), .A2(new_n991_), .B(new_n985_), .ZN(new_n1071_));
  OAI21_X1   g00861(.A1(new_n1070_), .A2(new_n1071_), .B(new_n1069_), .ZN(new_n1072_));
  NAND2_X1   g00862(.A1(new_n1072_), .A2(new_n1067_), .ZN(new_n1073_));
  NOR3_X1    g00863(.A1(new_n1051_), .A2(new_n1054_), .A3(new_n1055_), .ZN(new_n1074_));
  INV_X1     g00864(.I(new_n1074_), .ZN(new_n1075_));
  OAI21_X1   g00865(.A1(new_n1051_), .A2(new_n1054_), .B(new_n1055_), .ZN(new_n1076_));
  AOI21_X1   g00866(.A1(new_n1075_), .A2(new_n1076_), .B(new_n1073_), .ZN(new_n1077_));
  NOR2_X1    g00867(.A1(new_n1077_), .A2(new_n1065_), .ZN(new_n1078_));
  NOR2_X1    g00868(.A1(new_n958_), .A2(new_n957_), .ZN(new_n1079_));
  NOR2_X1    g00869(.A1(new_n1079_), .A2(new_n959_), .ZN(new_n1080_));
  XOR2_X1    g00870(.A1(new_n1078_), .A2(new_n1080_), .Z(new_n1081_));
  INV_X1     g00871(.I(new_n1057_), .ZN(new_n1082_));
  NOR3_X1    g00872(.A1(new_n1051_), .A2(new_n1054_), .A3(new_n1056_), .ZN(new_n1083_));
  OAI21_X1   g00873(.A1(new_n1082_), .A2(new_n1083_), .B(new_n1073_), .ZN(new_n1084_));
  AOI21_X1   g00874(.A1(new_n1060_), .A2(new_n1063_), .B(new_n1056_), .ZN(new_n1085_));
  OAI21_X1   g00875(.A1(new_n1074_), .A2(new_n1085_), .B(new_n999_), .ZN(new_n1086_));
  NAND3_X1   g00876(.A1(new_n945_), .A2(new_n937_), .A3(new_n941_), .ZN(new_n1087_));
  OAI21_X1   g00877(.A1(new_n957_), .A2(new_n958_), .B(new_n1087_), .ZN(new_n1088_));
  NAND3_X1   g00878(.A1(new_n1084_), .A2(new_n1088_), .A3(new_n1086_), .ZN(new_n1089_));
  OAI21_X1   g00879(.A1(new_n1077_), .A2(new_n1065_), .B(new_n1080_), .ZN(new_n1090_));
  NAND2_X1   g00880(.A1(new_n1090_), .A2(new_n1089_), .ZN(new_n1091_));
  NAND2_X1   g00881(.A1(new_n967_), .A2(new_n1091_), .ZN(new_n1092_));
  OAI21_X1   g00882(.A1(new_n967_), .A2(new_n1081_), .B(new_n1092_), .ZN(\asquared[19] ));
  NAND2_X1   g00883(.A1(new_n967_), .A2(new_n1089_), .ZN(new_n1094_));
  NAND2_X1   g00884(.A1(new_n1094_), .A2(new_n1090_), .ZN(new_n1095_));
  AOI21_X1   g00885(.A1(new_n1014_), .A2(new_n1050_), .B(new_n1058_), .ZN(new_n1096_));
  INV_X1     g00886(.I(new_n1010_), .ZN(new_n1097_));
  NOR2_X1    g00887(.A1(new_n1039_), .A2(new_n1037_), .ZN(new_n1098_));
  NAND2_X1   g00888(.A1(\a[6] ), .A2(\a[12] ), .ZN(new_n1099_));
  OAI21_X1   g00889(.A1(new_n1098_), .A2(new_n1099_), .B(new_n1040_), .ZN(new_n1100_));
  NAND2_X1   g00890(.A1(\a[8] ), .A2(\a[11] ), .ZN(new_n1101_));
  NOR2_X1    g00891(.A1(new_n525_), .A2(new_n1101_), .ZN(new_n1102_));
  NAND2_X1   g00892(.A1(new_n1102_), .A2(new_n200_), .ZN(new_n1103_));
  OAI21_X1   g00893(.A1(new_n525_), .A2(new_n1101_), .B(\a[3] ), .ZN(new_n1104_));
  AOI21_X1   g00894(.A1(new_n1103_), .A2(new_n1104_), .B(\a[16] ), .ZN(new_n1105_));
  AND3_X2    g00895(.A1(new_n1103_), .A2(\a[16] ), .A3(new_n1104_), .Z(new_n1106_));
  NOR2_X1    g00896(.A1(new_n1106_), .A2(new_n1105_), .ZN(new_n1107_));
  INV_X1     g00897(.I(new_n1107_), .ZN(new_n1108_));
  NAND2_X1   g00898(.A1(new_n1108_), .A2(new_n1100_), .ZN(new_n1109_));
  AOI21_X1   g00899(.A1(new_n1034_), .A2(new_n1030_), .B(new_n1099_), .ZN(new_n1110_));
  NOR2_X1    g00900(.A1(new_n1110_), .A2(new_n1035_), .ZN(new_n1111_));
  NAND2_X1   g00901(.A1(new_n1111_), .A2(new_n1107_), .ZN(new_n1112_));
  AOI21_X1   g00902(.A1(new_n1109_), .A2(new_n1112_), .B(new_n1097_), .ZN(new_n1113_));
  NOR2_X1    g00903(.A1(new_n1100_), .A2(new_n1107_), .ZN(new_n1114_));
  INV_X1     g00904(.I(new_n1114_), .ZN(new_n1115_));
  NAND2_X1   g00905(.A1(new_n1100_), .A2(new_n1107_), .ZN(new_n1116_));
  AOI21_X1   g00906(.A1(new_n1115_), .A2(new_n1116_), .B(new_n1010_), .ZN(new_n1117_));
  OAI22_X1   g00907(.A1(new_n1019_), .A2(new_n1016_), .B1(new_n225_), .B2(new_n1021_), .ZN(new_n1118_));
  NAND2_X1   g00908(.A1(\a[1] ), .A2(\a[18] ), .ZN(new_n1119_));
  NOR3_X1    g00909(.A1(new_n1118_), .A2(new_n1033_), .A3(new_n1119_), .ZN(new_n1120_));
  INV_X1     g00910(.I(new_n1120_), .ZN(new_n1121_));
  OAI21_X1   g00911(.A1(new_n1118_), .A2(new_n1119_), .B(new_n1033_), .ZN(new_n1122_));
  AOI21_X1   g00912(.A1(new_n1121_), .A2(new_n1122_), .B(\a[10] ), .ZN(new_n1123_));
  INV_X1     g00913(.I(new_n1122_), .ZN(new_n1124_));
  NOR3_X1    g00914(.A1(new_n1124_), .A2(new_n461_), .A3(new_n1120_), .ZN(new_n1125_));
  NOR2_X1    g00915(.A1(new_n1123_), .A2(new_n1125_), .ZN(new_n1126_));
  INV_X1     g00916(.I(new_n1126_), .ZN(new_n1127_));
  OAI21_X1   g00917(.A1(new_n1117_), .A2(new_n1113_), .B(new_n1127_), .ZN(new_n1128_));
  NOR2_X1    g00918(.A1(new_n1111_), .A2(new_n1107_), .ZN(new_n1129_));
  NOR2_X1    g00919(.A1(new_n1108_), .A2(new_n1100_), .ZN(new_n1130_));
  OAI21_X1   g00920(.A1(new_n1130_), .A2(new_n1129_), .B(new_n1010_), .ZN(new_n1131_));
  INV_X1     g00921(.I(new_n1116_), .ZN(new_n1132_));
  OAI21_X1   g00922(.A1(new_n1132_), .A2(new_n1114_), .B(new_n1097_), .ZN(new_n1133_));
  NAND3_X1   g00923(.A1(new_n1133_), .A2(new_n1131_), .A3(new_n1126_), .ZN(new_n1134_));
  AOI21_X1   g00924(.A1(new_n1128_), .A2(new_n1134_), .B(new_n1096_), .ZN(new_n1135_));
  OAI21_X1   g00925(.A1(new_n1015_), .A2(new_n1059_), .B(new_n1046_), .ZN(new_n1136_));
  NAND3_X1   g00926(.A1(new_n1133_), .A2(new_n1131_), .A3(new_n1127_), .ZN(new_n1137_));
  OAI21_X1   g00927(.A1(new_n1117_), .A2(new_n1113_), .B(new_n1126_), .ZN(new_n1138_));
  AOI21_X1   g00928(.A1(new_n1138_), .A2(new_n1137_), .B(new_n1136_), .ZN(new_n1139_));
  OAI21_X1   g00929(.A1(new_n1069_), .A2(new_n1071_), .B(new_n996_), .ZN(new_n1140_));
  NAND2_X1   g00930(.A1(\a[15] ), .A2(\a[17] ), .ZN(new_n1141_));
  NOR2_X1    g00931(.A1(new_n197_), .A2(new_n257_), .ZN(new_n1142_));
  INV_X1     g00932(.I(new_n1141_), .ZN(new_n1143_));
  NOR3_X1    g00933(.A1(new_n1142_), .A2(\a[19] ), .A3(new_n1143_), .ZN(new_n1144_));
  OR3_X2     g00934(.A1(new_n1144_), .A2(new_n260_), .A3(new_n1141_), .Z(new_n1145_));
  NAND3_X1   g00935(.A1(new_n1145_), .A2(\a[0] ), .A3(\a[19] ), .ZN(new_n1146_));
  NAND2_X1   g00936(.A1(new_n260_), .A2(new_n1141_), .ZN(new_n1147_));
  NAND2_X1   g00937(.A1(new_n1146_), .A2(new_n1147_), .ZN(new_n1148_));
  NOR2_X1    g00938(.A1(new_n982_), .A2(new_n877_), .ZN(new_n1149_));
  NAND2_X1   g00939(.A1(\a[12] ), .A2(\a[13] ), .ZN(new_n1150_));
  INV_X1     g00940(.I(new_n1000_), .ZN(new_n1151_));
  AOI22_X1   g00941(.A1(new_n608_), .A2(new_n654_), .B1(new_n787_), .B2(new_n1151_), .ZN(new_n1152_));
  NOR2_X1    g00942(.A1(new_n353_), .A2(new_n650_), .ZN(new_n1153_));
  NAND4_X1   g00943(.A1(new_n1152_), .A2(new_n478_), .A3(new_n1150_), .A4(new_n1153_), .ZN(new_n1154_));
  NOR3_X1    g00944(.A1(new_n1149_), .A2(new_n990_), .A3(new_n1154_), .ZN(new_n1155_));
  INV_X1     g00945(.I(new_n1155_), .ZN(new_n1156_));
  OAI21_X1   g00946(.A1(new_n1149_), .A2(new_n990_), .B(new_n1154_), .ZN(new_n1157_));
  AOI21_X1   g00947(.A1(new_n1156_), .A2(new_n1157_), .B(new_n1148_), .ZN(new_n1158_));
  INV_X1     g00948(.I(new_n1148_), .ZN(new_n1159_));
  INV_X1     g00949(.I(new_n1154_), .ZN(new_n1160_));
  OAI21_X1   g00950(.A1(new_n1149_), .A2(new_n990_), .B(new_n1160_), .ZN(new_n1161_));
  NOR3_X1    g00951(.A1(new_n1149_), .A2(new_n990_), .A3(new_n1160_), .ZN(new_n1162_));
  INV_X1     g00952(.I(new_n1162_), .ZN(new_n1163_));
  AOI21_X1   g00953(.A1(new_n1163_), .A2(new_n1161_), .B(new_n1159_), .ZN(new_n1164_));
  NOR2_X1    g00954(.A1(new_n1164_), .A2(new_n1158_), .ZN(new_n1165_));
  NOR2_X1    g00955(.A1(new_n1165_), .A2(new_n1140_), .ZN(new_n1166_));
  AOI21_X1   g00956(.A1(new_n995_), .A2(new_n997_), .B(new_n1070_), .ZN(new_n1167_));
  NOR3_X1    g00957(.A1(new_n1167_), .A2(new_n1158_), .A3(new_n1164_), .ZN(new_n1168_));
  OAI22_X1   g00958(.A1(new_n1135_), .A2(new_n1139_), .B1(new_n1166_), .B2(new_n1168_), .ZN(new_n1169_));
  AOI21_X1   g00959(.A1(new_n1133_), .A2(new_n1131_), .B(new_n1126_), .ZN(new_n1170_));
  NOR3_X1    g00960(.A1(new_n1117_), .A2(new_n1113_), .A3(new_n1127_), .ZN(new_n1171_));
  OAI21_X1   g00961(.A1(new_n1171_), .A2(new_n1170_), .B(new_n1136_), .ZN(new_n1172_));
  NOR3_X1    g00962(.A1(new_n1117_), .A2(new_n1113_), .A3(new_n1126_), .ZN(new_n1173_));
  AOI21_X1   g00963(.A1(new_n1133_), .A2(new_n1131_), .B(new_n1127_), .ZN(new_n1174_));
  OAI21_X1   g00964(.A1(new_n1173_), .A2(new_n1174_), .B(new_n1096_), .ZN(new_n1175_));
  AOI21_X1   g00965(.A1(new_n898_), .A2(new_n970_), .B(new_n1071_), .ZN(new_n1176_));
  OAI22_X1   g00966(.A1(new_n1176_), .A2(new_n1070_), .B1(new_n1158_), .B2(new_n1164_), .ZN(new_n1177_));
  INV_X1     g00967(.I(new_n1157_), .ZN(new_n1178_));
  OAI21_X1   g00968(.A1(new_n1178_), .A2(new_n1155_), .B(new_n1159_), .ZN(new_n1179_));
  INV_X1     g00969(.I(new_n1161_), .ZN(new_n1180_));
  OAI21_X1   g00970(.A1(new_n1180_), .A2(new_n1162_), .B(new_n1148_), .ZN(new_n1181_));
  NAND3_X1   g00971(.A1(new_n1167_), .A2(new_n1179_), .A3(new_n1181_), .ZN(new_n1182_));
  NAND2_X1   g00972(.A1(new_n1177_), .A2(new_n1182_), .ZN(new_n1183_));
  NAND3_X1   g00973(.A1(new_n1183_), .A2(new_n1172_), .A3(new_n1175_), .ZN(new_n1184_));
  NAND2_X1   g00974(.A1(new_n1184_), .A2(new_n1169_), .ZN(new_n1185_));
  OAI21_X1   g00975(.A1(new_n1073_), .A2(new_n1083_), .B(new_n1057_), .ZN(new_n1186_));
  XNOR2_X1   g00976(.A1(new_n1185_), .A2(new_n1186_), .ZN(new_n1187_));
  NAND3_X1   g00977(.A1(new_n1184_), .A2(new_n1169_), .A3(new_n1186_), .ZN(new_n1188_));
  AOI21_X1   g00978(.A1(new_n1184_), .A2(new_n1169_), .B(new_n1186_), .ZN(new_n1189_));
  INV_X1     g00979(.I(new_n1189_), .ZN(new_n1190_));
  NAND2_X1   g00980(.A1(new_n1190_), .A2(new_n1188_), .ZN(new_n1191_));
  MUX2_X1    g00981(.I0(new_n1187_), .I1(new_n1191_), .S(new_n1095_), .Z(\asquared[20] ));
  OAI21_X1   g00982(.A1(new_n1188_), .A2(new_n1090_), .B(new_n1089_), .ZN(new_n1193_));
  OAI21_X1   g00983(.A1(new_n966_), .A2(new_n961_), .B(new_n1193_), .ZN(new_n1194_));
  NOR4_X1    g00984(.A1(new_n971_), .A2(new_n359_), .A3(new_n650_), .A4(new_n875_), .ZN(new_n1195_));
  NOR3_X1    g00985(.A1(new_n341_), .A2(new_n481_), .A3(new_n653_), .ZN(new_n1196_));
  NOR2_X1    g00986(.A1(new_n1196_), .A2(new_n1195_), .ZN(new_n1197_));
  NOR2_X1    g00987(.A1(new_n242_), .A2(new_n650_), .ZN(new_n1198_));
  INV_X1     g00988(.I(new_n1198_), .ZN(new_n1199_));
  OAI21_X1   g00989(.A1(new_n481_), .A2(new_n1018_), .B(new_n1197_), .ZN(new_n1200_));
  OAI21_X1   g00990(.A1(new_n1200_), .A2(new_n1199_), .B(new_n875_), .ZN(new_n1201_));
  NAND2_X1   g00991(.A1(new_n1201_), .A2(\a[5] ), .ZN(new_n1202_));
  NOR2_X1    g00992(.A1(\a[8] ), .A2(\a[12] ), .ZN(new_n1203_));
  AOI21_X1   g00993(.A1(new_n1202_), .A2(new_n1203_), .B(new_n1197_), .ZN(new_n1204_));
  INV_X1     g00994(.I(new_n1152_), .ZN(new_n1205_));
  OAI21_X1   g00995(.A1(new_n478_), .A2(new_n1150_), .B(new_n1205_), .ZN(new_n1206_));
  NOR2_X1    g00996(.A1(new_n1119_), .A2(new_n461_), .ZN(new_n1207_));
  INV_X1     g00997(.I(new_n1207_), .ZN(new_n1208_));
  NAND2_X1   g00998(.A1(\a[7] ), .A2(\a[13] ), .ZN(new_n1209_));
  NOR2_X1    g00999(.A1(new_n1208_), .A2(new_n1209_), .ZN(new_n1210_));
  NAND2_X1   g01000(.A1(new_n1210_), .A2(new_n199_), .ZN(new_n1211_));
  NAND3_X1   g01001(.A1(new_n1207_), .A2(\a[7] ), .A3(\a[13] ), .ZN(new_n1212_));
  NAND2_X1   g01002(.A1(new_n1212_), .A2(\a[0] ), .ZN(new_n1213_));
  AOI21_X1   g01003(.A1(new_n1211_), .A2(new_n1213_), .B(\a[20] ), .ZN(new_n1214_));
  INV_X1     g01004(.I(\a[20] ), .ZN(new_n1215_));
  NOR2_X1    g01005(.A1(new_n1212_), .A2(\a[0] ), .ZN(new_n1216_));
  INV_X1     g01006(.I(new_n1213_), .ZN(new_n1217_));
  NOR3_X1    g01007(.A1(new_n1217_), .A2(new_n1215_), .A3(new_n1216_), .ZN(new_n1218_));
  OAI21_X1   g01008(.A1(new_n1218_), .A2(new_n1214_), .B(new_n1206_), .ZN(new_n1219_));
  INV_X1     g01009(.I(new_n1150_), .ZN(new_n1220_));
  AOI21_X1   g01010(.A1(new_n479_), .A2(new_n1220_), .B(new_n1152_), .ZN(new_n1221_));
  OAI21_X1   g01011(.A1(new_n1217_), .A2(new_n1216_), .B(new_n1215_), .ZN(new_n1222_));
  NAND3_X1   g01012(.A1(new_n1211_), .A2(\a[20] ), .A3(new_n1213_), .ZN(new_n1223_));
  NAND3_X1   g01013(.A1(new_n1222_), .A2(new_n1223_), .A3(new_n1221_), .ZN(new_n1224_));
  NAND2_X1   g01014(.A1(new_n1219_), .A2(new_n1224_), .ZN(new_n1225_));
  AOI21_X1   g01015(.A1(new_n1222_), .A2(new_n1223_), .B(new_n1206_), .ZN(new_n1226_));
  NOR3_X1    g01016(.A1(new_n1218_), .A2(new_n1214_), .A3(new_n1221_), .ZN(new_n1227_));
  NOR2_X1    g01017(.A1(new_n1227_), .A2(new_n1226_), .ZN(new_n1228_));
  NOR2_X1    g01018(.A1(new_n1228_), .A2(new_n1204_), .ZN(new_n1229_));
  AOI21_X1   g01019(.A1(new_n1204_), .A2(new_n1225_), .B(new_n1229_), .ZN(new_n1230_));
  NOR2_X1    g01020(.A1(new_n1162_), .A2(new_n1148_), .ZN(new_n1231_));
  NOR2_X1    g01021(.A1(new_n1231_), .A2(new_n1180_), .ZN(new_n1232_));
  NOR2_X1    g01022(.A1(new_n260_), .A2(new_n1141_), .ZN(new_n1233_));
  NAND2_X1   g01023(.A1(\a[3] ), .A2(\a[16] ), .ZN(new_n1234_));
  AOI21_X1   g01024(.A1(new_n525_), .A2(new_n1101_), .B(new_n1234_), .ZN(new_n1235_));
  NAND2_X1   g01025(.A1(\a[9] ), .A2(\a[11] ), .ZN(new_n1236_));
  NAND2_X1   g01026(.A1(\a[1] ), .A2(\a[19] ), .ZN(new_n1237_));
  XNOR2_X1   g01027(.A1(new_n1236_), .A2(new_n1237_), .ZN(new_n1238_));
  NOR3_X1    g01028(.A1(new_n1238_), .A2(new_n1102_), .A3(new_n1235_), .ZN(new_n1239_));
  NOR2_X1    g01029(.A1(new_n1235_), .A2(new_n1102_), .ZN(new_n1240_));
  INV_X1     g01030(.I(new_n1238_), .ZN(new_n1241_));
  NOR2_X1    g01031(.A1(new_n1241_), .A2(new_n1240_), .ZN(new_n1242_));
  NOR2_X1    g01032(.A1(new_n1242_), .A2(new_n1239_), .ZN(new_n1243_));
  XNOR2_X1   g01033(.A1(new_n1238_), .A2(new_n1240_), .ZN(new_n1244_));
  NAND2_X1   g01034(.A1(new_n1244_), .A2(new_n1233_), .ZN(new_n1245_));
  OAI21_X1   g01035(.A1(new_n1233_), .A2(new_n1243_), .B(new_n1245_), .ZN(new_n1246_));
  NAND2_X1   g01036(.A1(new_n1232_), .A2(new_n1246_), .ZN(new_n1247_));
  INV_X1     g01037(.I(new_n1246_), .ZN(new_n1248_));
  OAI21_X1   g01038(.A1(new_n1231_), .A2(new_n1180_), .B(new_n1248_), .ZN(new_n1249_));
  AOI21_X1   g01039(.A1(new_n1247_), .A2(new_n1249_), .B(new_n1230_), .ZN(new_n1250_));
  NAND2_X1   g01040(.A1(new_n1225_), .A2(new_n1204_), .ZN(new_n1251_));
  OAI21_X1   g01041(.A1(new_n1204_), .A2(new_n1228_), .B(new_n1251_), .ZN(new_n1252_));
  OAI21_X1   g01042(.A1(new_n1180_), .A2(new_n1231_), .B(new_n1246_), .ZN(new_n1253_));
  NOR3_X1    g01043(.A1(new_n1246_), .A2(new_n1231_), .A3(new_n1180_), .ZN(new_n1254_));
  INV_X1     g01044(.I(new_n1254_), .ZN(new_n1255_));
  AOI21_X1   g01045(.A1(new_n1253_), .A2(new_n1255_), .B(new_n1252_), .ZN(new_n1256_));
  NOR2_X1    g01046(.A1(new_n1250_), .A2(new_n1256_), .ZN(new_n1257_));
  INV_X1     g01047(.I(new_n1257_), .ZN(new_n1258_));
  AOI21_X1   g01048(.A1(new_n1136_), .A2(new_n1137_), .B(new_n1174_), .ZN(new_n1259_));
  OAI21_X1   g01049(.A1(new_n1097_), .A2(new_n1130_), .B(new_n1109_), .ZN(new_n1260_));
  INV_X1     g01050(.I(new_n1118_), .ZN(new_n1261_));
  INV_X1     g01051(.I(new_n1119_), .ZN(new_n1262_));
  OAI21_X1   g01052(.A1(new_n1038_), .A2(new_n1262_), .B(new_n1261_), .ZN(new_n1263_));
  NOR2_X1    g01053(.A1(new_n1262_), .A2(\a[10] ), .ZN(new_n1264_));
  OAI21_X1   g01054(.A1(new_n1207_), .A2(new_n1264_), .B(new_n1038_), .ZN(new_n1265_));
  NAND2_X1   g01055(.A1(new_n1263_), .A2(new_n1265_), .ZN(new_n1266_));
  NAND2_X1   g01056(.A1(\a[16] ), .A2(\a[18] ), .ZN(new_n1267_));
  NAND2_X1   g01057(.A1(\a[17] ), .A2(\a[18] ), .ZN(new_n1268_));
  NOR2_X1    g01058(.A1(new_n1267_), .A2(new_n1268_), .ZN(new_n1269_));
  INV_X1     g01059(.I(new_n1269_), .ZN(new_n1270_));
  NOR2_X1    g01060(.A1(new_n225_), .A2(new_n260_), .ZN(new_n1271_));
  INV_X1     g01061(.I(new_n1271_), .ZN(new_n1272_));
  NAND2_X1   g01062(.A1(new_n1270_), .A2(new_n1272_), .ZN(new_n1273_));
  NAND2_X1   g01063(.A1(\a[16] ), .A2(\a[17] ), .ZN(new_n1274_));
  INV_X1     g01064(.I(new_n1274_), .ZN(new_n1275_));
  INV_X1     g01065(.I(\a[18] ), .ZN(new_n1276_));
  NOR2_X1    g01066(.A1(new_n201_), .A2(new_n1276_), .ZN(new_n1277_));
  INV_X1     g01067(.I(new_n1277_), .ZN(new_n1278_));
  NOR4_X1    g01068(.A1(new_n1273_), .A2(new_n267_), .A3(new_n1275_), .A4(new_n1278_), .ZN(new_n1279_));
  XOR2_X1    g01069(.A1(new_n1266_), .A2(new_n1279_), .Z(new_n1280_));
  NAND2_X1   g01070(.A1(new_n1266_), .A2(new_n1279_), .ZN(new_n1281_));
  INV_X1     g01071(.I(new_n1281_), .ZN(new_n1282_));
  NOR2_X1    g01072(.A1(new_n1266_), .A2(new_n1279_), .ZN(new_n1283_));
  NOR2_X1    g01073(.A1(new_n1282_), .A2(new_n1283_), .ZN(new_n1284_));
  NOR2_X1    g01074(.A1(new_n1284_), .A2(new_n1260_), .ZN(new_n1285_));
  AOI21_X1   g01075(.A1(new_n1260_), .A2(new_n1280_), .B(new_n1285_), .ZN(new_n1286_));
  NOR2_X1    g01076(.A1(new_n1286_), .A2(new_n1259_), .ZN(new_n1287_));
  OAI21_X1   g01077(.A1(new_n1096_), .A2(new_n1173_), .B(new_n1138_), .ZN(new_n1288_));
  NAND2_X1   g01078(.A1(new_n1280_), .A2(new_n1260_), .ZN(new_n1289_));
  OAI21_X1   g01079(.A1(new_n1260_), .A2(new_n1284_), .B(new_n1289_), .ZN(new_n1290_));
  NOR2_X1    g01080(.A1(new_n1288_), .A2(new_n1290_), .ZN(new_n1291_));
  OAI22_X1   g01081(.A1(new_n1287_), .A2(new_n1291_), .B1(new_n1250_), .B2(new_n1256_), .ZN(new_n1292_));
  NOR2_X1    g01082(.A1(new_n1286_), .A2(new_n1288_), .ZN(new_n1293_));
  NOR2_X1    g01083(.A1(new_n1259_), .A2(new_n1290_), .ZN(new_n1294_));
  NOR2_X1    g01084(.A1(new_n1293_), .A2(new_n1294_), .ZN(new_n1295_));
  OAI21_X1   g01085(.A1(new_n1258_), .A2(new_n1295_), .B(new_n1292_), .ZN(new_n1296_));
  NAND2_X1   g01086(.A1(new_n1172_), .A2(new_n1175_), .ZN(new_n1297_));
  INV_X1     g01087(.I(new_n1168_), .ZN(new_n1298_));
  OAI21_X1   g01088(.A1(new_n1297_), .A2(new_n1166_), .B(new_n1298_), .ZN(new_n1299_));
  NAND2_X1   g01089(.A1(new_n1296_), .A2(new_n1299_), .ZN(new_n1300_));
  XOR2_X1    g01090(.A1(new_n1194_), .A2(new_n1300_), .Z(new_n1301_));
  XOR2_X1    g01091(.A1(new_n1301_), .A2(new_n1189_), .Z(\asquared[21] ));
  NAND2_X1   g01092(.A1(new_n1296_), .A2(new_n1189_), .ZN(new_n1303_));
  OAI21_X1   g01093(.A1(new_n1296_), .A2(new_n1189_), .B(new_n1299_), .ZN(new_n1304_));
  OAI21_X1   g01094(.A1(new_n1194_), .A2(new_n1304_), .B(new_n1303_), .ZN(new_n1305_));
  INV_X1     g01095(.I(new_n1294_), .ZN(new_n1306_));
  OAI21_X1   g01096(.A1(new_n1258_), .A2(new_n1293_), .B(new_n1306_), .ZN(new_n1307_));
  INV_X1     g01097(.I(new_n1224_), .ZN(new_n1308_));
  AOI21_X1   g01098(.A1(new_n1204_), .A2(new_n1219_), .B(new_n1308_), .ZN(new_n1309_));
  NOR2_X1    g01099(.A1(new_n1239_), .A2(new_n1233_), .ZN(new_n1310_));
  NOR2_X1    g01100(.A1(new_n1310_), .A2(new_n1242_), .ZN(new_n1311_));
  INV_X1     g01101(.I(new_n1311_), .ZN(new_n1312_));
  INV_X1     g01102(.I(\a[21] ), .ZN(new_n1313_));
  NOR2_X1    g01103(.A1(new_n1236_), .A2(new_n1237_), .ZN(new_n1314_));
  NOR2_X1    g01104(.A1(new_n194_), .A2(new_n1215_), .ZN(new_n1315_));
  NAND2_X1   g01105(.A1(\a[11] ), .A2(\a[20] ), .ZN(new_n1316_));
  OAI22_X1   g01106(.A1(new_n1315_), .A2(\a[11] ), .B1(new_n194_), .B2(new_n1316_), .ZN(new_n1317_));
  NAND2_X1   g01107(.A1(new_n1317_), .A2(new_n1314_), .ZN(new_n1318_));
  XOR2_X1    g01108(.A1(new_n1318_), .A2(new_n199_), .Z(new_n1319_));
  NAND2_X1   g01109(.A1(new_n1319_), .A2(new_n1313_), .ZN(new_n1320_));
  XOR2_X1    g01110(.A1(new_n1318_), .A2(\a[0] ), .Z(new_n1321_));
  NAND2_X1   g01111(.A1(new_n1321_), .A2(\a[21] ), .ZN(new_n1322_));
  NAND2_X1   g01112(.A1(new_n1320_), .A2(new_n1322_), .ZN(new_n1323_));
  NAND2_X1   g01113(.A1(new_n1323_), .A2(new_n1312_), .ZN(new_n1324_));
  NOR2_X1    g01114(.A1(new_n1321_), .A2(\a[21] ), .ZN(new_n1325_));
  NOR2_X1    g01115(.A1(new_n1319_), .A2(new_n1313_), .ZN(new_n1326_));
  NOR2_X1    g01116(.A1(new_n1325_), .A2(new_n1326_), .ZN(new_n1327_));
  NAND2_X1   g01117(.A1(new_n1327_), .A2(new_n1311_), .ZN(new_n1328_));
  AOI21_X1   g01118(.A1(new_n1328_), .A2(new_n1324_), .B(new_n1309_), .ZN(new_n1329_));
  NAND2_X1   g01119(.A1(new_n1204_), .A2(new_n1219_), .ZN(new_n1330_));
  NAND2_X1   g01120(.A1(new_n1330_), .A2(new_n1224_), .ZN(new_n1331_));
  NAND2_X1   g01121(.A1(new_n1323_), .A2(new_n1311_), .ZN(new_n1332_));
  NAND2_X1   g01122(.A1(new_n1327_), .A2(new_n1312_), .ZN(new_n1333_));
  AOI21_X1   g01123(.A1(new_n1332_), .A2(new_n1333_), .B(new_n1331_), .ZN(new_n1334_));
  OAI21_X1   g01124(.A1(new_n1230_), .A2(new_n1254_), .B(new_n1253_), .ZN(new_n1335_));
  AOI21_X1   g01125(.A1(new_n1010_), .A2(new_n1112_), .B(new_n1129_), .ZN(new_n1336_));
  OAI21_X1   g01126(.A1(new_n1336_), .A2(new_n1283_), .B(new_n1281_), .ZN(new_n1337_));
  NOR3_X1    g01127(.A1(new_n201_), .A2(new_n800_), .A3(new_n1276_), .ZN(new_n1338_));
  INV_X1     g01128(.I(\a[19] ), .ZN(new_n1339_));
  NOR2_X1    g01129(.A1(new_n200_), .A2(new_n1339_), .ZN(new_n1340_));
  NOR3_X1    g01130(.A1(new_n1338_), .A2(\a[5] ), .A3(new_n1340_), .ZN(new_n1341_));
  NAND2_X1   g01131(.A1(\a[18] ), .A2(\a[19] ), .ZN(new_n1342_));
  OR3_X2     g01132(.A1(new_n1341_), .A2(new_n225_), .A3(new_n1342_), .Z(new_n1343_));
  NOR2_X1    g01133(.A1(new_n353_), .A2(new_n800_), .ZN(new_n1344_));
  OAI21_X1   g01134(.A1(new_n1276_), .A2(new_n1339_), .B(new_n225_), .ZN(new_n1345_));
  INV_X1     g01135(.I(new_n1345_), .ZN(new_n1346_));
  AOI21_X1   g01136(.A1(new_n1343_), .A2(new_n1344_), .B(new_n1346_), .ZN(new_n1347_));
  INV_X1     g01137(.I(new_n1347_), .ZN(new_n1348_));
  OAI22_X1   g01138(.A1(new_n341_), .A2(new_n1018_), .B1(new_n478_), .B2(new_n873_), .ZN(new_n1349_));
  NAND2_X1   g01139(.A1(\a[6] ), .A2(\a[15] ), .ZN(new_n1350_));
  NOR4_X1    g01140(.A1(new_n1349_), .A2(new_n609_), .A3(new_n787_), .A4(new_n1350_), .ZN(new_n1351_));
  INV_X1     g01141(.I(new_n1351_), .ZN(new_n1352_));
  OAI21_X1   g01142(.A1(new_n364_), .A2(new_n566_), .B(new_n796_), .ZN(new_n1353_));
  NAND2_X1   g01143(.A1(\a[4] ), .A2(\a[17] ), .ZN(new_n1354_));
  AOI21_X1   g01144(.A1(new_n1353_), .A2(new_n1354_), .B(new_n651_), .ZN(new_n1355_));
  NAND2_X1   g01145(.A1(new_n1355_), .A2(new_n525_), .ZN(new_n1356_));
  OR2_X2     g01146(.A1(new_n1355_), .A2(new_n525_), .Z(new_n1357_));
  AOI21_X1   g01147(.A1(new_n1357_), .A2(new_n1356_), .B(new_n1352_), .ZN(new_n1358_));
  INV_X1     g01148(.I(new_n1358_), .ZN(new_n1359_));
  NAND3_X1   g01149(.A1(new_n1357_), .A2(new_n1352_), .A3(new_n1356_), .ZN(new_n1360_));
  AOI21_X1   g01150(.A1(new_n1359_), .A2(new_n1360_), .B(new_n1348_), .ZN(new_n1361_));
  AOI21_X1   g01151(.A1(new_n1357_), .A2(new_n1356_), .B(new_n1351_), .ZN(new_n1362_));
  INV_X1     g01152(.I(new_n1362_), .ZN(new_n1363_));
  NAND3_X1   g01153(.A1(new_n1357_), .A2(new_n1351_), .A3(new_n1356_), .ZN(new_n1364_));
  AOI21_X1   g01154(.A1(new_n1363_), .A2(new_n1364_), .B(new_n1347_), .ZN(new_n1365_));
  INV_X1     g01155(.I(new_n1200_), .ZN(new_n1366_));
  AOI22_X1   g01156(.A1(new_n1270_), .A2(new_n1272_), .B1(new_n267_), .B2(new_n1275_), .ZN(new_n1367_));
  NAND2_X1   g01157(.A1(\a[0] ), .A2(\a[20] ), .ZN(new_n1368_));
  AOI21_X1   g01158(.A1(new_n1208_), .A2(new_n1209_), .B(new_n1368_), .ZN(new_n1369_));
  NOR2_X1    g01159(.A1(new_n1369_), .A2(new_n1210_), .ZN(new_n1370_));
  NOR2_X1    g01160(.A1(new_n1370_), .A2(new_n1367_), .ZN(new_n1371_));
  NAND2_X1   g01161(.A1(new_n1370_), .A2(new_n1367_), .ZN(new_n1372_));
  INV_X1     g01162(.I(new_n1372_), .ZN(new_n1373_));
  OAI21_X1   g01163(.A1(new_n1373_), .A2(new_n1371_), .B(new_n1366_), .ZN(new_n1374_));
  INV_X1     g01164(.I(new_n1367_), .ZN(new_n1375_));
  NOR2_X1    g01165(.A1(new_n1375_), .A2(new_n1370_), .ZN(new_n1376_));
  OR2_X2     g01166(.A1(new_n1369_), .A2(new_n1210_), .Z(new_n1377_));
  NOR2_X1    g01167(.A1(new_n1377_), .A2(new_n1367_), .ZN(new_n1378_));
  OAI21_X1   g01168(.A1(new_n1378_), .A2(new_n1376_), .B(new_n1200_), .ZN(new_n1379_));
  NAND2_X1   g01169(.A1(new_n1374_), .A2(new_n1379_), .ZN(new_n1380_));
  OAI21_X1   g01170(.A1(new_n1361_), .A2(new_n1365_), .B(new_n1380_), .ZN(new_n1381_));
  INV_X1     g01171(.I(new_n1360_), .ZN(new_n1382_));
  OAI21_X1   g01172(.A1(new_n1382_), .A2(new_n1358_), .B(new_n1347_), .ZN(new_n1383_));
  INV_X1     g01173(.I(new_n1364_), .ZN(new_n1384_));
  OAI21_X1   g01174(.A1(new_n1384_), .A2(new_n1362_), .B(new_n1348_), .ZN(new_n1385_));
  INV_X1     g01175(.I(new_n1371_), .ZN(new_n1386_));
  AOI21_X1   g01176(.A1(new_n1386_), .A2(new_n1372_), .B(new_n1200_), .ZN(new_n1387_));
  NAND2_X1   g01177(.A1(new_n1377_), .A2(new_n1367_), .ZN(new_n1388_));
  NAND2_X1   g01178(.A1(new_n1375_), .A2(new_n1370_), .ZN(new_n1389_));
  AOI21_X1   g01179(.A1(new_n1388_), .A2(new_n1389_), .B(new_n1366_), .ZN(new_n1390_));
  NOR2_X1    g01180(.A1(new_n1387_), .A2(new_n1390_), .ZN(new_n1391_));
  NAND3_X1   g01181(.A1(new_n1391_), .A2(new_n1383_), .A3(new_n1385_), .ZN(new_n1392_));
  NAND2_X1   g01182(.A1(new_n1381_), .A2(new_n1392_), .ZN(new_n1393_));
  NAND2_X1   g01183(.A1(new_n1393_), .A2(new_n1337_), .ZN(new_n1394_));
  INV_X1     g01184(.I(new_n1283_), .ZN(new_n1395_));
  AOI21_X1   g01185(.A1(new_n1260_), .A2(new_n1395_), .B(new_n1282_), .ZN(new_n1396_));
  NOR3_X1    g01186(.A1(new_n1391_), .A2(new_n1361_), .A3(new_n1365_), .ZN(new_n1397_));
  AOI21_X1   g01187(.A1(new_n1383_), .A2(new_n1385_), .B(new_n1380_), .ZN(new_n1398_));
  OAI21_X1   g01188(.A1(new_n1398_), .A2(new_n1397_), .B(new_n1396_), .ZN(new_n1399_));
  AOI21_X1   g01189(.A1(new_n1394_), .A2(new_n1399_), .B(new_n1335_), .ZN(new_n1400_));
  NOR2_X1    g01190(.A1(new_n1248_), .A2(new_n1232_), .ZN(new_n1401_));
  AOI21_X1   g01191(.A1(new_n1252_), .A2(new_n1255_), .B(new_n1401_), .ZN(new_n1402_));
  AOI21_X1   g01192(.A1(new_n1381_), .A2(new_n1392_), .B(new_n1396_), .ZN(new_n1403_));
  NAND3_X1   g01193(.A1(new_n1380_), .A2(new_n1383_), .A3(new_n1385_), .ZN(new_n1404_));
  OAI21_X1   g01194(.A1(new_n1361_), .A2(new_n1365_), .B(new_n1391_), .ZN(new_n1405_));
  AOI21_X1   g01195(.A1(new_n1405_), .A2(new_n1404_), .B(new_n1337_), .ZN(new_n1406_));
  NOR3_X1    g01196(.A1(new_n1402_), .A2(new_n1403_), .A3(new_n1406_), .ZN(new_n1407_));
  OAI22_X1   g01197(.A1(new_n1400_), .A2(new_n1407_), .B1(new_n1329_), .B2(new_n1334_), .ZN(new_n1408_));
  NOR2_X1    g01198(.A1(new_n1334_), .A2(new_n1329_), .ZN(new_n1409_));
  AOI21_X1   g01199(.A1(new_n1394_), .A2(new_n1399_), .B(new_n1402_), .ZN(new_n1410_));
  NOR3_X1    g01200(.A1(new_n1335_), .A2(new_n1403_), .A3(new_n1406_), .ZN(new_n1411_));
  OAI21_X1   g01201(.A1(new_n1410_), .A2(new_n1411_), .B(new_n1409_), .ZN(new_n1412_));
  NAND2_X1   g01202(.A1(new_n1408_), .A2(new_n1412_), .ZN(new_n1413_));
  XNOR2_X1   g01203(.A1(new_n1413_), .A2(new_n1307_), .ZN(new_n1414_));
  INV_X1     g01204(.I(new_n1307_), .ZN(new_n1415_));
  NAND2_X1   g01205(.A1(new_n1415_), .A2(new_n1413_), .ZN(new_n1416_));
  NAND3_X1   g01206(.A1(new_n1307_), .A2(new_n1408_), .A3(new_n1412_), .ZN(new_n1417_));
  NAND2_X1   g01207(.A1(new_n1416_), .A2(new_n1417_), .ZN(new_n1418_));
  MUX2_X1    g01208(.I0(new_n1418_), .I1(new_n1414_), .S(new_n1305_), .Z(\asquared[22] ));
  NAND2_X1   g01209(.A1(new_n1305_), .A2(new_n1416_), .ZN(new_n1420_));
  NAND2_X1   g01210(.A1(new_n1420_), .A2(new_n1417_), .ZN(new_n1421_));
  OAI21_X1   g01211(.A1(new_n1403_), .A2(new_n1406_), .B(new_n1402_), .ZN(new_n1422_));
  AOI21_X1   g01212(.A1(new_n1422_), .A2(new_n1409_), .B(new_n1407_), .ZN(new_n1423_));
  NOR2_X1    g01213(.A1(new_n1327_), .A2(new_n1312_), .ZN(new_n1424_));
  OAI21_X1   g01214(.A1(new_n1309_), .A2(new_n1424_), .B(new_n1333_), .ZN(new_n1425_));
  NAND3_X1   g01215(.A1(new_n232_), .A2(\a[18] ), .A3(\a[19] ), .ZN(new_n1426_));
  INV_X1     g01216(.I(new_n1426_), .ZN(new_n1427_));
  OAI21_X1   g01217(.A1(new_n392_), .A2(new_n786_), .B(new_n1349_), .ZN(new_n1428_));
  NOR2_X1    g01218(.A1(new_n199_), .A2(new_n1313_), .ZN(new_n1429_));
  OAI21_X1   g01219(.A1(new_n1317_), .A2(new_n1314_), .B(new_n1429_), .ZN(new_n1430_));
  NAND2_X1   g01220(.A1(new_n1430_), .A2(new_n1318_), .ZN(new_n1431_));
  XOR2_X1    g01221(.A1(new_n1431_), .A2(new_n1428_), .Z(new_n1432_));
  NOR2_X1    g01222(.A1(new_n1432_), .A2(new_n1427_), .ZN(new_n1433_));
  INV_X1     g01223(.I(new_n1428_), .ZN(new_n1434_));
  NAND2_X1   g01224(.A1(new_n1431_), .A2(new_n1434_), .ZN(new_n1435_));
  INV_X1     g01225(.I(new_n1435_), .ZN(new_n1436_));
  NOR2_X1    g01226(.A1(new_n1431_), .A2(new_n1434_), .ZN(new_n1437_));
  OAI21_X1   g01227(.A1(new_n1436_), .A2(new_n1437_), .B(new_n1427_), .ZN(new_n1438_));
  INV_X1     g01228(.I(new_n1438_), .ZN(new_n1439_));
  NOR2_X1    g01229(.A1(new_n1439_), .A2(new_n1433_), .ZN(new_n1440_));
  INV_X1     g01230(.I(new_n1268_), .ZN(new_n1441_));
  NOR2_X1    g01231(.A1(new_n211_), .A2(new_n1268_), .ZN(new_n1445_));
  INV_X1     g01232(.I(new_n1445_), .ZN(new_n1446_));
  INV_X1     g01233(.I(new_n1018_), .ZN(new_n1447_));
  NAND2_X1   g01234(.A1(new_n1447_), .A2(new_n609_), .ZN(new_n1448_));
  NAND2_X1   g01235(.A1(\a[0] ), .A2(\a[22] ), .ZN(new_n1449_));
  XNOR2_X1   g01236(.A1(new_n1448_), .A2(new_n1449_), .ZN(new_n1450_));
  INV_X1     g01237(.I(new_n1450_), .ZN(new_n1451_));
  NOR2_X1    g01238(.A1(new_n596_), .A2(new_n798_), .ZN(new_n1452_));
  XOR2_X1    g01239(.A1(new_n1452_), .A2(\a[2] ), .Z(new_n1453_));
  NAND2_X1   g01240(.A1(new_n1453_), .A2(new_n1215_), .ZN(new_n1454_));
  XOR2_X1    g01241(.A1(new_n1452_), .A2(new_n201_), .Z(new_n1455_));
  NAND2_X1   g01242(.A1(new_n1455_), .A2(\a[20] ), .ZN(new_n1456_));
  NAND2_X1   g01243(.A1(new_n1454_), .A2(new_n1456_), .ZN(new_n1457_));
  NAND2_X1   g01244(.A1(new_n1457_), .A2(new_n1451_), .ZN(new_n1458_));
  NAND3_X1   g01245(.A1(new_n1454_), .A2(new_n1456_), .A3(new_n1450_), .ZN(new_n1459_));
  AOI21_X1   g01246(.A1(new_n1458_), .A2(new_n1459_), .B(new_n1446_), .ZN(new_n1460_));
  NAND2_X1   g01247(.A1(new_n1457_), .A2(new_n1450_), .ZN(new_n1461_));
  NAND3_X1   g01248(.A1(new_n1451_), .A2(new_n1454_), .A3(new_n1456_), .ZN(new_n1462_));
  AOI21_X1   g01249(.A1(new_n1461_), .A2(new_n1462_), .B(new_n1445_), .ZN(new_n1463_));
  NOR2_X1    g01250(.A1(new_n1460_), .A2(new_n1463_), .ZN(new_n1464_));
  NOR2_X1    g01251(.A1(new_n1464_), .A2(new_n1440_), .ZN(new_n1465_));
  OAI21_X1   g01252(.A1(new_n1427_), .A2(new_n1432_), .B(new_n1438_), .ZN(new_n1466_));
  NOR3_X1    g01253(.A1(new_n1466_), .A2(new_n1460_), .A3(new_n1463_), .ZN(new_n1467_));
  OAI21_X1   g01254(.A1(new_n1465_), .A2(new_n1467_), .B(new_n1425_), .ZN(new_n1468_));
  NOR2_X1    g01255(.A1(new_n1323_), .A2(new_n1311_), .ZN(new_n1469_));
  AOI21_X1   g01256(.A1(new_n1331_), .A2(new_n1332_), .B(new_n1469_), .ZN(new_n1470_));
  NOR2_X1    g01257(.A1(new_n1464_), .A2(new_n1466_), .ZN(new_n1471_));
  NOR3_X1    g01258(.A1(new_n1440_), .A2(new_n1460_), .A3(new_n1463_), .ZN(new_n1472_));
  OAI21_X1   g01259(.A1(new_n1471_), .A2(new_n1472_), .B(new_n1470_), .ZN(new_n1473_));
  AOI21_X1   g01260(.A1(new_n1337_), .A2(new_n1404_), .B(new_n1398_), .ZN(new_n1474_));
  AOI21_X1   g01261(.A1(new_n1347_), .A2(new_n1360_), .B(new_n1358_), .ZN(new_n1475_));
  INV_X1     g01262(.I(new_n1475_), .ZN(new_n1476_));
  AOI21_X1   g01263(.A1(new_n1366_), .A2(new_n1389_), .B(new_n1376_), .ZN(new_n1477_));
  NAND2_X1   g01264(.A1(\a[1] ), .A2(\a[21] ), .ZN(new_n1478_));
  INV_X1     g01265(.I(new_n523_), .ZN(new_n1479_));
  NOR2_X1    g01266(.A1(new_n651_), .A2(new_n1354_), .ZN(new_n1480_));
  NOR4_X1    g01267(.A1(new_n364_), .A2(new_n461_), .A3(\a[11] ), .A4(\a[12] ), .ZN(new_n1481_));
  NOR2_X1    g01268(.A1(new_n1480_), .A2(new_n1481_), .ZN(new_n1482_));
  NAND2_X1   g01269(.A1(new_n1315_), .A2(\a[11] ), .ZN(new_n1483_));
  XNOR2_X1   g01270(.A1(new_n1482_), .A2(new_n1483_), .ZN(new_n1484_));
  NOR2_X1    g01271(.A1(new_n1484_), .A2(new_n1479_), .ZN(new_n1485_));
  XOR2_X1    g01272(.A1(new_n1482_), .A2(new_n1483_), .Z(new_n1486_));
  NOR2_X1    g01273(.A1(new_n1486_), .A2(new_n523_), .ZN(new_n1487_));
  OAI21_X1   g01274(.A1(new_n1485_), .A2(new_n1487_), .B(new_n1478_), .ZN(new_n1488_));
  INV_X1     g01275(.I(new_n1478_), .ZN(new_n1489_));
  NAND2_X1   g01276(.A1(new_n1486_), .A2(new_n523_), .ZN(new_n1490_));
  NAND2_X1   g01277(.A1(new_n1484_), .A2(new_n1479_), .ZN(new_n1491_));
  NAND3_X1   g01278(.A1(new_n1491_), .A2(new_n1490_), .A3(new_n1489_), .ZN(new_n1492_));
  AOI21_X1   g01279(.A1(new_n1488_), .A2(new_n1492_), .B(new_n1477_), .ZN(new_n1493_));
  OAI21_X1   g01280(.A1(new_n1200_), .A2(new_n1378_), .B(new_n1388_), .ZN(new_n1494_));
  AOI21_X1   g01281(.A1(new_n1491_), .A2(new_n1490_), .B(new_n1489_), .ZN(new_n1495_));
  NOR3_X1    g01282(.A1(new_n1485_), .A2(new_n1487_), .A3(new_n1478_), .ZN(new_n1496_));
  NOR3_X1    g01283(.A1(new_n1495_), .A2(new_n1496_), .A3(new_n1494_), .ZN(new_n1497_));
  OAI21_X1   g01284(.A1(new_n1497_), .A2(new_n1493_), .B(new_n1476_), .ZN(new_n1498_));
  AOI21_X1   g01285(.A1(new_n1488_), .A2(new_n1492_), .B(new_n1494_), .ZN(new_n1499_));
  NOR3_X1    g01286(.A1(new_n1496_), .A2(new_n1495_), .A3(new_n1477_), .ZN(new_n1500_));
  OAI21_X1   g01287(.A1(new_n1499_), .A2(new_n1500_), .B(new_n1475_), .ZN(new_n1501_));
  NAND2_X1   g01288(.A1(new_n1501_), .A2(new_n1498_), .ZN(new_n1502_));
  NAND2_X1   g01289(.A1(new_n1502_), .A2(new_n1474_), .ZN(new_n1503_));
  OAI21_X1   g01290(.A1(new_n1396_), .A2(new_n1397_), .B(new_n1405_), .ZN(new_n1504_));
  NAND3_X1   g01291(.A1(new_n1504_), .A2(new_n1498_), .A3(new_n1501_), .ZN(new_n1505_));
  AOI22_X1   g01292(.A1(new_n1503_), .A2(new_n1505_), .B1(new_n1473_), .B2(new_n1468_), .ZN(new_n1506_));
  NAND2_X1   g01293(.A1(new_n1473_), .A2(new_n1468_), .ZN(new_n1507_));
  NAND2_X1   g01294(.A1(new_n1404_), .A2(new_n1337_), .ZN(new_n1508_));
  AOI22_X1   g01295(.A1(new_n1508_), .A2(new_n1405_), .B1(new_n1501_), .B2(new_n1498_), .ZN(new_n1509_));
  NOR2_X1    g01296(.A1(new_n1502_), .A2(new_n1504_), .ZN(new_n1510_));
  NOR2_X1    g01297(.A1(new_n1510_), .A2(new_n1509_), .ZN(new_n1511_));
  NOR2_X1    g01298(.A1(new_n1511_), .A2(new_n1507_), .ZN(new_n1512_));
  OAI21_X1   g01299(.A1(new_n1512_), .A2(new_n1506_), .B(new_n1423_), .ZN(new_n1513_));
  INV_X1     g01300(.I(new_n1513_), .ZN(new_n1514_));
  NOR3_X1    g01301(.A1(new_n1512_), .A2(new_n1423_), .A3(new_n1506_), .ZN(new_n1515_));
  NOR2_X1    g01302(.A1(new_n1514_), .A2(new_n1515_), .ZN(new_n1516_));
  XNOR2_X1   g01303(.A1(new_n1421_), .A2(new_n1516_), .ZN(\asquared[23] ));
  NOR2_X1    g01304(.A1(new_n1515_), .A2(new_n1413_), .ZN(new_n1518_));
  AOI21_X1   g01305(.A1(new_n1515_), .A2(new_n1413_), .B(new_n1307_), .ZN(new_n1519_));
  NOR2_X1    g01306(.A1(new_n1519_), .A2(new_n1518_), .ZN(new_n1520_));
  NAND2_X1   g01307(.A1(new_n1305_), .A2(new_n1520_), .ZN(new_n1521_));
  INV_X1     g01308(.I(new_n1507_), .ZN(new_n1522_));
  INV_X1     g01309(.I(new_n1505_), .ZN(new_n1523_));
  AOI21_X1   g01310(.A1(new_n1522_), .A2(new_n1503_), .B(new_n1523_), .ZN(new_n1524_));
  NAND2_X1   g01311(.A1(new_n1464_), .A2(new_n1466_), .ZN(new_n1525_));
  AOI21_X1   g01312(.A1(new_n1425_), .A2(new_n1525_), .B(new_n1471_), .ZN(new_n1526_));
  INV_X1     g01313(.I(new_n1500_), .ZN(new_n1527_));
  OAI21_X1   g01314(.A1(new_n1496_), .A2(new_n1495_), .B(new_n1477_), .ZN(new_n1528_));
  NAND2_X1   g01315(.A1(new_n1528_), .A2(new_n1476_), .ZN(new_n1529_));
  NAND2_X1   g01316(.A1(new_n1529_), .A2(new_n1527_), .ZN(new_n1530_));
  NOR2_X1    g01317(.A1(new_n353_), .A2(new_n1276_), .ZN(new_n1531_));
  INV_X1     g01318(.I(new_n1531_), .ZN(new_n1532_));
  NAND2_X1   g01319(.A1(\a[3] ), .A2(\a[6] ), .ZN(new_n1533_));
  NAND2_X1   g01320(.A1(\a[17] ), .A2(\a[20] ), .ZN(new_n1534_));
  OAI22_X1   g01321(.A1(new_n1533_), .A2(new_n1534_), .B1(new_n481_), .B2(new_n1268_), .ZN(new_n1535_));
  NAND2_X1   g01322(.A1(\a[18] ), .A2(\a[20] ), .ZN(new_n1536_));
  NOR2_X1    g01323(.A1(new_n261_), .A2(new_n1536_), .ZN(new_n1537_));
  NOR2_X1    g01324(.A1(new_n1535_), .A2(new_n1537_), .ZN(new_n1538_));
  INV_X1     g01325(.I(new_n1538_), .ZN(new_n1539_));
  OAI21_X1   g01326(.A1(new_n1539_), .A2(new_n1532_), .B(new_n1215_), .ZN(new_n1540_));
  NAND2_X1   g01327(.A1(new_n1540_), .A2(\a[3] ), .ZN(new_n1541_));
  NOR2_X1    g01328(.A1(\a[6] ), .A2(\a[17] ), .ZN(new_n1542_));
  INV_X1     g01329(.I(new_n1537_), .ZN(new_n1543_));
  NAND2_X1   g01330(.A1(new_n1543_), .A2(new_n1535_), .ZN(new_n1544_));
  AOI21_X1   g01331(.A1(new_n1541_), .A2(new_n1542_), .B(new_n1544_), .ZN(new_n1545_));
  INV_X1     g01332(.I(new_n1545_), .ZN(new_n1546_));
  NOR2_X1    g01333(.A1(new_n1482_), .A2(new_n1483_), .ZN(new_n1547_));
  XNOR2_X1   g01334(.A1(new_n523_), .A2(new_n1478_), .ZN(new_n1548_));
  AOI21_X1   g01335(.A1(new_n1482_), .A2(new_n1483_), .B(new_n1548_), .ZN(new_n1549_));
  NOR2_X1    g01336(.A1(new_n1549_), .A2(new_n1547_), .ZN(new_n1550_));
  OAI21_X1   g01337(.A1(new_n461_), .A2(new_n599_), .B(new_n651_), .ZN(new_n1551_));
  INV_X1     g01338(.I(new_n1551_), .ZN(new_n1552_));
  NAND3_X1   g01339(.A1(new_n1552_), .A2(new_n1220_), .A3(new_n797_), .ZN(new_n1553_));
  NAND2_X1   g01340(.A1(\a[4] ), .A2(\a[19] ), .ZN(new_n1554_));
  XOR2_X1    g01341(.A1(new_n1553_), .A2(new_n1554_), .Z(new_n1555_));
  XOR2_X1    g01342(.A1(new_n1555_), .A2(new_n1550_), .Z(new_n1556_));
  NOR2_X1    g01343(.A1(new_n1556_), .A2(new_n1546_), .ZN(new_n1557_));
  XNOR2_X1   g01344(.A1(new_n1553_), .A2(new_n1554_), .ZN(new_n1558_));
  NOR2_X1    g01345(.A1(new_n1558_), .A2(new_n1550_), .ZN(new_n1559_));
  INV_X1     g01346(.I(new_n1559_), .ZN(new_n1560_));
  NAND2_X1   g01347(.A1(new_n1558_), .A2(new_n1550_), .ZN(new_n1561_));
  AOI21_X1   g01348(.A1(new_n1560_), .A2(new_n1561_), .B(new_n1545_), .ZN(new_n1562_));
  NOR2_X1    g01349(.A1(\a[0] ), .A2(\a[22] ), .ZN(new_n1563_));
  OAI21_X1   g01350(.A1(new_n392_), .A2(new_n1018_), .B(new_n1563_), .ZN(new_n1564_));
  OAI21_X1   g01351(.A1(new_n609_), .A2(new_n1447_), .B(new_n1564_), .ZN(new_n1565_));
  NAND2_X1   g01352(.A1(\a[21] ), .A2(\a[23] ), .ZN(new_n1566_));
  XNOR2_X1   g01353(.A1(new_n197_), .A2(new_n1566_), .ZN(new_n1567_));
  OAI22_X1   g01354(.A1(new_n392_), .A2(new_n1017_), .B1(new_n772_), .B2(new_n1021_), .ZN(new_n1568_));
  NAND4_X1   g01355(.A1(new_n453_), .A2(new_n1018_), .A3(\a[7] ), .A4(\a[16] ), .ZN(new_n1569_));
  NOR2_X1    g01356(.A1(new_n1568_), .A2(new_n1569_), .ZN(new_n1570_));
  XOR2_X1    g01357(.A1(new_n1570_), .A2(new_n1567_), .Z(new_n1571_));
  NOR2_X1    g01358(.A1(new_n1571_), .A2(new_n1565_), .ZN(new_n1572_));
  INV_X1     g01359(.I(new_n1567_), .ZN(new_n1573_));
  NAND2_X1   g01360(.A1(new_n1573_), .A2(new_n1570_), .ZN(new_n1574_));
  NOR2_X1    g01361(.A1(new_n1573_), .A2(new_n1570_), .ZN(new_n1575_));
  INV_X1     g01362(.I(new_n1575_), .ZN(new_n1576_));
  NAND2_X1   g01363(.A1(new_n1576_), .A2(new_n1574_), .ZN(new_n1577_));
  AOI21_X1   g01364(.A1(new_n1565_), .A2(new_n1577_), .B(new_n1572_), .ZN(new_n1578_));
  NOR3_X1    g01365(.A1(new_n1557_), .A2(new_n1562_), .A3(new_n1578_), .ZN(new_n1579_));
  OAI21_X1   g01366(.A1(new_n1557_), .A2(new_n1562_), .B(new_n1578_), .ZN(new_n1580_));
  INV_X1     g01367(.I(new_n1580_), .ZN(new_n1581_));
  OAI21_X1   g01368(.A1(new_n1581_), .A2(new_n1579_), .B(new_n1530_), .ZN(new_n1582_));
  AOI21_X1   g01369(.A1(new_n1476_), .A2(new_n1528_), .B(new_n1500_), .ZN(new_n1583_));
  XOR2_X1    g01370(.A1(new_n1558_), .A2(new_n1550_), .Z(new_n1584_));
  NAND2_X1   g01371(.A1(new_n1584_), .A2(new_n1545_), .ZN(new_n1585_));
  INV_X1     g01372(.I(new_n1561_), .ZN(new_n1586_));
  OAI21_X1   g01373(.A1(new_n1586_), .A2(new_n1559_), .B(new_n1546_), .ZN(new_n1587_));
  AOI21_X1   g01374(.A1(new_n1585_), .A2(new_n1587_), .B(new_n1578_), .ZN(new_n1588_));
  INV_X1     g01375(.I(new_n1578_), .ZN(new_n1589_));
  NOR3_X1    g01376(.A1(new_n1557_), .A2(new_n1562_), .A3(new_n1589_), .ZN(new_n1590_));
  OAI21_X1   g01377(.A1(new_n1588_), .A2(new_n1590_), .B(new_n1583_), .ZN(new_n1591_));
  OAI21_X1   g01378(.A1(new_n1427_), .A2(new_n1437_), .B(new_n1435_), .ZN(new_n1592_));
  NAND2_X1   g01379(.A1(new_n1459_), .A2(new_n1445_), .ZN(new_n1593_));
  NAND2_X1   g01380(.A1(new_n1593_), .A2(new_n1458_), .ZN(new_n1594_));
  INV_X1     g01381(.I(new_n1594_), .ZN(new_n1595_));
  AOI22_X1   g01382(.A1(\a[6] ), .A2(\a[16] ), .B1(\a[9] ), .B2(\a[13] ), .ZN(new_n1596_));
  NAND2_X1   g01383(.A1(\a[2] ), .A2(\a[20] ), .ZN(new_n1597_));
  NOR2_X1    g01384(.A1(new_n1596_), .A2(new_n1597_), .ZN(new_n1598_));
  NOR2_X1    g01385(.A1(new_n1598_), .A2(new_n1452_), .ZN(new_n1599_));
  OAI22_X1   g01386(.A1(new_n211_), .A2(new_n1268_), .B1(new_n212_), .B2(new_n1342_), .ZN(new_n1600_));
  NAND2_X1   g01387(.A1(\a[1] ), .A2(\a[22] ), .ZN(new_n1601_));
  XOR2_X1    g01388(.A1(new_n1600_), .A2(new_n1601_), .Z(new_n1602_));
  XOR2_X1    g01389(.A1(new_n1602_), .A2(new_n1599_), .Z(new_n1603_));
  XOR2_X1    g01390(.A1(new_n1603_), .A2(\a[12] ), .Z(new_n1604_));
  NOR2_X1    g01391(.A1(new_n1604_), .A2(new_n1595_), .ZN(new_n1605_));
  XNOR2_X1   g01392(.A1(new_n1602_), .A2(new_n1599_), .ZN(new_n1606_));
  NAND2_X1   g01393(.A1(new_n1606_), .A2(new_n566_), .ZN(new_n1607_));
  NAND2_X1   g01394(.A1(new_n1603_), .A2(\a[12] ), .ZN(new_n1608_));
  NAND2_X1   g01395(.A1(new_n1607_), .A2(new_n1608_), .ZN(new_n1609_));
  NOR2_X1    g01396(.A1(new_n1609_), .A2(new_n1594_), .ZN(new_n1610_));
  OAI21_X1   g01397(.A1(new_n1605_), .A2(new_n1610_), .B(new_n1592_), .ZN(new_n1611_));
  INV_X1     g01398(.I(new_n1592_), .ZN(new_n1612_));
  NOR2_X1    g01399(.A1(new_n1604_), .A2(new_n1594_), .ZN(new_n1613_));
  NAND3_X1   g01400(.A1(new_n1594_), .A2(new_n1607_), .A3(new_n1608_), .ZN(new_n1614_));
  INV_X1     g01401(.I(new_n1614_), .ZN(new_n1615_));
  OAI21_X1   g01402(.A1(new_n1613_), .A2(new_n1615_), .B(new_n1612_), .ZN(new_n1616_));
  NAND2_X1   g01403(.A1(new_n1611_), .A2(new_n1616_), .ZN(new_n1617_));
  NAND3_X1   g01404(.A1(new_n1617_), .A2(new_n1582_), .A3(new_n1591_), .ZN(new_n1618_));
  NAND3_X1   g01405(.A1(new_n1585_), .A2(new_n1587_), .A3(new_n1589_), .ZN(new_n1619_));
  AOI21_X1   g01406(.A1(new_n1619_), .A2(new_n1580_), .B(new_n1583_), .ZN(new_n1620_));
  OAI21_X1   g01407(.A1(new_n1557_), .A2(new_n1562_), .B(new_n1589_), .ZN(new_n1621_));
  NAND3_X1   g01408(.A1(new_n1585_), .A2(new_n1587_), .A3(new_n1578_), .ZN(new_n1622_));
  AOI21_X1   g01409(.A1(new_n1622_), .A2(new_n1621_), .B(new_n1530_), .ZN(new_n1623_));
  NAND2_X1   g01410(.A1(new_n1609_), .A2(new_n1594_), .ZN(new_n1624_));
  NAND2_X1   g01411(.A1(new_n1604_), .A2(new_n1595_), .ZN(new_n1625_));
  AOI21_X1   g01412(.A1(new_n1625_), .A2(new_n1624_), .B(new_n1612_), .ZN(new_n1626_));
  NAND2_X1   g01413(.A1(new_n1609_), .A2(new_n1595_), .ZN(new_n1627_));
  AOI21_X1   g01414(.A1(new_n1627_), .A2(new_n1614_), .B(new_n1592_), .ZN(new_n1628_));
  NOR2_X1    g01415(.A1(new_n1626_), .A2(new_n1628_), .ZN(new_n1629_));
  OAI21_X1   g01416(.A1(new_n1620_), .A2(new_n1623_), .B(new_n1629_), .ZN(new_n1630_));
  AOI21_X1   g01417(.A1(new_n1630_), .A2(new_n1618_), .B(new_n1526_), .ZN(new_n1631_));
  INV_X1     g01418(.I(new_n1526_), .ZN(new_n1632_));
  OAI22_X1   g01419(.A1(new_n1623_), .A2(new_n1620_), .B1(new_n1626_), .B2(new_n1628_), .ZN(new_n1633_));
  NAND3_X1   g01420(.A1(new_n1582_), .A2(new_n1629_), .A3(new_n1591_), .ZN(new_n1634_));
  AOI21_X1   g01421(.A1(new_n1634_), .A2(new_n1633_), .B(new_n1632_), .ZN(new_n1635_));
  NOR2_X1    g01422(.A1(new_n1631_), .A2(new_n1635_), .ZN(new_n1636_));
  OR2_X2     g01423(.A1(new_n1636_), .A2(new_n1524_), .Z(new_n1637_));
  XOR2_X1    g01424(.A1(new_n1521_), .A2(new_n1637_), .Z(new_n1638_));
  XOR2_X1    g01425(.A1(new_n1638_), .A2(new_n1514_), .Z(\asquared[24] ));
  AOI21_X1   g01426(.A1(new_n1636_), .A2(new_n1524_), .B(new_n1513_), .ZN(new_n1640_));
  NAND3_X1   g01427(.A1(new_n1305_), .A2(new_n1520_), .A3(new_n1640_), .ZN(new_n1641_));
  NAND2_X1   g01428(.A1(new_n1641_), .A2(new_n1637_), .ZN(new_n1642_));
  NAND2_X1   g01429(.A1(new_n1633_), .A2(new_n1632_), .ZN(new_n1643_));
  NAND2_X1   g01430(.A1(new_n1643_), .A2(new_n1634_), .ZN(new_n1644_));
  AOI21_X1   g01431(.A1(new_n1530_), .A2(new_n1621_), .B(new_n1590_), .ZN(new_n1645_));
  INV_X1     g01432(.I(new_n1645_), .ZN(new_n1646_));
  AOI21_X1   g01433(.A1(new_n1545_), .A2(new_n1561_), .B(new_n1559_), .ZN(new_n1647_));
  INV_X1     g01434(.I(new_n1647_), .ZN(new_n1648_));
  NAND2_X1   g01435(.A1(new_n1220_), .A2(new_n797_), .ZN(new_n1649_));
  NOR2_X1    g01436(.A1(\a[4] ), .A2(\a[19] ), .ZN(new_n1650_));
  AOI21_X1   g01437(.A1(new_n1649_), .A2(new_n1650_), .B(new_n1551_), .ZN(new_n1651_));
  OAI21_X1   g01438(.A1(new_n453_), .A2(new_n1018_), .B(new_n1568_), .ZN(new_n1652_));
  XOR2_X1    g01439(.A1(new_n1652_), .A2(new_n1651_), .Z(new_n1653_));
  NOR2_X1    g01440(.A1(new_n1653_), .A2(new_n1539_), .ZN(new_n1654_));
  INV_X1     g01441(.I(new_n1651_), .ZN(new_n1655_));
  NOR2_X1    g01442(.A1(new_n1655_), .A2(new_n1652_), .ZN(new_n1656_));
  INV_X1     g01443(.I(new_n1656_), .ZN(new_n1657_));
  NAND2_X1   g01444(.A1(new_n1655_), .A2(new_n1652_), .ZN(new_n1658_));
  AOI21_X1   g01445(.A1(new_n1657_), .A2(new_n1658_), .B(new_n1538_), .ZN(new_n1659_));
  NOR2_X1    g01446(.A1(new_n1659_), .A2(new_n1654_), .ZN(new_n1660_));
  OAI21_X1   g01447(.A1(new_n1565_), .A2(new_n1575_), .B(new_n1574_), .ZN(new_n1661_));
  XOR2_X1    g01448(.A1(new_n1660_), .A2(new_n1661_), .Z(new_n1662_));
  NAND2_X1   g01449(.A1(new_n1662_), .A2(new_n1648_), .ZN(new_n1663_));
  NAND2_X1   g01450(.A1(new_n1660_), .A2(new_n1661_), .ZN(new_n1664_));
  NOR2_X1    g01451(.A1(new_n1660_), .A2(new_n1661_), .ZN(new_n1665_));
  INV_X1     g01452(.I(new_n1665_), .ZN(new_n1666_));
  AOI21_X1   g01453(.A1(new_n1666_), .A2(new_n1664_), .B(new_n1648_), .ZN(new_n1667_));
  INV_X1     g01454(.I(new_n1667_), .ZN(new_n1668_));
  NAND2_X1   g01455(.A1(new_n1668_), .A2(new_n1663_), .ZN(new_n1669_));
  NOR2_X1    g01456(.A1(new_n1599_), .A2(new_n1600_), .ZN(new_n1670_));
  XOR2_X1    g01457(.A1(new_n1601_), .A2(\a[12] ), .Z(new_n1671_));
  AOI21_X1   g01458(.A1(new_n1599_), .A2(new_n1600_), .B(new_n1671_), .ZN(new_n1672_));
  NOR2_X1    g01459(.A1(new_n1672_), .A2(new_n1670_), .ZN(new_n1673_));
  INV_X1     g01460(.I(\a[22] ), .ZN(new_n1674_));
  NOR2_X1    g01461(.A1(new_n1276_), .A2(new_n1674_), .ZN(new_n1675_));
  INV_X1     g01462(.I(new_n1675_), .ZN(new_n1676_));
  NOR3_X1    g01463(.A1(new_n1676_), .A2(new_n201_), .A3(new_n242_), .ZN(new_n1681_));
  INV_X1     g01464(.I(new_n1681_), .ZN(new_n1682_));
  NOR2_X1    g01465(.A1(new_n1601_), .A2(new_n566_), .ZN(new_n1683_));
  NAND2_X1   g01466(.A1(\a[1] ), .A2(\a[23] ), .ZN(new_n1684_));
  INV_X1     g01467(.I(new_n1684_), .ZN(new_n1685_));
  NOR2_X1    g01468(.A1(new_n1001_), .A2(new_n1685_), .ZN(new_n1686_));
  NOR2_X1    g01469(.A1(new_n870_), .A2(new_n1684_), .ZN(new_n1687_));
  OAI21_X1   g01470(.A1(new_n1686_), .A2(new_n1687_), .B(new_n1683_), .ZN(new_n1688_));
  XOR2_X1    g01471(.A1(new_n1688_), .A2(\a[0] ), .Z(new_n1689_));
  NOR2_X1    g01472(.A1(new_n1689_), .A2(\a[24] ), .ZN(new_n1690_));
  INV_X1     g01473(.I(\a[24] ), .ZN(new_n1691_));
  XOR2_X1    g01474(.A1(new_n1688_), .A2(new_n199_), .Z(new_n1692_));
  NOR2_X1    g01475(.A1(new_n1692_), .A2(new_n1691_), .ZN(new_n1693_));
  OAI21_X1   g01476(.A1(new_n1690_), .A2(new_n1693_), .B(new_n1682_), .ZN(new_n1694_));
  NAND2_X1   g01477(.A1(new_n1692_), .A2(new_n1691_), .ZN(new_n1695_));
  NAND2_X1   g01478(.A1(new_n1689_), .A2(\a[24] ), .ZN(new_n1696_));
  NAND3_X1   g01479(.A1(new_n1695_), .A2(new_n1696_), .A3(new_n1681_), .ZN(new_n1697_));
  AOI21_X1   g01480(.A1(new_n1694_), .A2(new_n1697_), .B(new_n1673_), .ZN(new_n1698_));
  INV_X1     g01481(.I(new_n1673_), .ZN(new_n1699_));
  OAI21_X1   g01482(.A1(new_n1690_), .A2(new_n1693_), .B(new_n1681_), .ZN(new_n1700_));
  NAND3_X1   g01483(.A1(new_n1695_), .A2(new_n1696_), .A3(new_n1682_), .ZN(new_n1701_));
  AOI21_X1   g01484(.A1(new_n1700_), .A2(new_n1701_), .B(new_n1699_), .ZN(new_n1702_));
  NOR2_X1    g01485(.A1(new_n1698_), .A2(new_n1702_), .ZN(new_n1703_));
  INV_X1     g01486(.I(new_n1703_), .ZN(new_n1704_));
  AOI21_X1   g01487(.A1(new_n1609_), .A2(new_n1595_), .B(new_n1612_), .ZN(new_n1705_));
  NAND2_X1   g01488(.A1(\a[21] ), .A2(\a[23] ), .ZN(new_n1706_));
  INV_X1     g01489(.I(new_n1706_), .ZN(new_n1707_));
  NOR2_X1    g01490(.A1(new_n523_), .A2(new_n1478_), .ZN(new_n1708_));
  AOI21_X1   g01491(.A1(new_n1708_), .A2(new_n218_), .B(new_n1707_), .ZN(new_n1709_));
  NAND2_X1   g01492(.A1(\a[19] ), .A2(\a[21] ), .ZN(new_n1710_));
  NAND2_X1   g01493(.A1(\a[20] ), .A2(\a[21] ), .ZN(new_n1711_));
  NOR2_X1    g01494(.A1(new_n1710_), .A2(new_n1711_), .ZN(new_n1712_));
  NOR2_X1    g01495(.A1(new_n212_), .A2(new_n261_), .ZN(new_n1713_));
  NOR2_X1    g01496(.A1(new_n1712_), .A2(new_n1713_), .ZN(new_n1714_));
  NAND2_X1   g01497(.A1(\a[19] ), .A2(\a[20] ), .ZN(new_n1715_));
  NOR2_X1    g01498(.A1(new_n200_), .A2(new_n1313_), .ZN(new_n1716_));
  NAND4_X1   g01499(.A1(new_n1714_), .A2(new_n211_), .A3(new_n1715_), .A4(new_n1716_), .ZN(new_n1717_));
  INV_X1     g01500(.I(new_n1017_), .ZN(new_n1718_));
  INV_X1     g01501(.I(new_n1021_), .ZN(new_n1719_));
  NOR2_X1    g01502(.A1(new_n391_), .A2(new_n453_), .ZN(new_n1720_));
  AOI21_X1   g01503(.A1(new_n1718_), .A2(new_n1719_), .B(new_n1720_), .ZN(new_n1721_));
  NOR2_X1    g01504(.A1(new_n359_), .A2(new_n800_), .ZN(new_n1722_));
  NAND4_X1   g01505(.A1(new_n1721_), .A2(new_n525_), .A3(new_n1018_), .A4(new_n1722_), .ZN(new_n1723_));
  XNOR2_X1   g01506(.A1(new_n1723_), .A2(new_n1717_), .ZN(new_n1724_));
  NOR2_X1    g01507(.A1(new_n1724_), .A2(new_n1709_), .ZN(new_n1725_));
  INV_X1     g01508(.I(new_n1709_), .ZN(new_n1726_));
  OR2_X2     g01509(.A1(new_n1723_), .A2(new_n1717_), .Z(new_n1727_));
  NAND2_X1   g01510(.A1(new_n1723_), .A2(new_n1717_), .ZN(new_n1728_));
  AOI21_X1   g01511(.A1(new_n1727_), .A2(new_n1728_), .B(new_n1726_), .ZN(new_n1729_));
  NOR2_X1    g01512(.A1(new_n1725_), .A2(new_n1729_), .ZN(new_n1730_));
  NOR3_X1    g01513(.A1(new_n1705_), .A2(new_n1615_), .A3(new_n1730_), .ZN(new_n1731_));
  OAI21_X1   g01514(.A1(new_n1604_), .A2(new_n1594_), .B(new_n1592_), .ZN(new_n1732_));
  INV_X1     g01515(.I(new_n1730_), .ZN(new_n1733_));
  AOI21_X1   g01516(.A1(new_n1732_), .A2(new_n1614_), .B(new_n1733_), .ZN(new_n1734_));
  OAI21_X1   g01517(.A1(new_n1734_), .A2(new_n1731_), .B(new_n1704_), .ZN(new_n1735_));
  AOI21_X1   g01518(.A1(new_n1732_), .A2(new_n1614_), .B(new_n1730_), .ZN(new_n1736_));
  NOR3_X1    g01519(.A1(new_n1705_), .A2(new_n1615_), .A3(new_n1733_), .ZN(new_n1737_));
  OAI21_X1   g01520(.A1(new_n1736_), .A2(new_n1737_), .B(new_n1703_), .ZN(new_n1738_));
  AOI21_X1   g01521(.A1(new_n1735_), .A2(new_n1738_), .B(new_n1669_), .ZN(new_n1739_));
  AOI21_X1   g01522(.A1(new_n1662_), .A2(new_n1648_), .B(new_n1667_), .ZN(new_n1740_));
  NAND3_X1   g01523(.A1(new_n1732_), .A2(new_n1614_), .A3(new_n1733_), .ZN(new_n1741_));
  OAI21_X1   g01524(.A1(new_n1705_), .A2(new_n1615_), .B(new_n1730_), .ZN(new_n1742_));
  AOI21_X1   g01525(.A1(new_n1741_), .A2(new_n1742_), .B(new_n1703_), .ZN(new_n1743_));
  OAI21_X1   g01526(.A1(new_n1705_), .A2(new_n1615_), .B(new_n1733_), .ZN(new_n1744_));
  NAND3_X1   g01527(.A1(new_n1732_), .A2(new_n1614_), .A3(new_n1730_), .ZN(new_n1745_));
  AOI21_X1   g01528(.A1(new_n1745_), .A2(new_n1744_), .B(new_n1704_), .ZN(new_n1746_));
  NOR3_X1    g01529(.A1(new_n1743_), .A2(new_n1746_), .A3(new_n1740_), .ZN(new_n1747_));
  OAI21_X1   g01530(.A1(new_n1739_), .A2(new_n1747_), .B(new_n1646_), .ZN(new_n1748_));
  AOI21_X1   g01531(.A1(new_n1735_), .A2(new_n1738_), .B(new_n1740_), .ZN(new_n1749_));
  NOR3_X1    g01532(.A1(new_n1743_), .A2(new_n1746_), .A3(new_n1669_), .ZN(new_n1750_));
  OAI21_X1   g01533(.A1(new_n1749_), .A2(new_n1750_), .B(new_n1645_), .ZN(new_n1751_));
  AOI21_X1   g01534(.A1(new_n1751_), .A2(new_n1748_), .B(new_n1644_), .ZN(new_n1752_));
  NOR3_X1    g01535(.A1(new_n1617_), .A2(new_n1620_), .A3(new_n1623_), .ZN(new_n1753_));
  AOI21_X1   g01536(.A1(new_n1632_), .A2(new_n1633_), .B(new_n1753_), .ZN(new_n1754_));
  OAI21_X1   g01537(.A1(new_n1743_), .A2(new_n1746_), .B(new_n1740_), .ZN(new_n1755_));
  NAND3_X1   g01538(.A1(new_n1735_), .A2(new_n1738_), .A3(new_n1669_), .ZN(new_n1756_));
  AOI21_X1   g01539(.A1(new_n1756_), .A2(new_n1755_), .B(new_n1645_), .ZN(new_n1757_));
  OAI21_X1   g01540(.A1(new_n1743_), .A2(new_n1746_), .B(new_n1669_), .ZN(new_n1758_));
  NAND3_X1   g01541(.A1(new_n1735_), .A2(new_n1738_), .A3(new_n1740_), .ZN(new_n1759_));
  AOI21_X1   g01542(.A1(new_n1758_), .A2(new_n1759_), .B(new_n1646_), .ZN(new_n1760_));
  NOR3_X1    g01543(.A1(new_n1757_), .A2(new_n1760_), .A3(new_n1754_), .ZN(new_n1761_));
  NOR2_X1    g01544(.A1(new_n1752_), .A2(new_n1761_), .ZN(new_n1762_));
  XNOR2_X1   g01545(.A1(new_n1642_), .A2(new_n1762_), .ZN(\asquared[25] ));
  INV_X1     g01546(.I(new_n1752_), .ZN(new_n1764_));
  OAI21_X1   g01547(.A1(new_n1642_), .A2(new_n1761_), .B(new_n1764_), .ZN(new_n1765_));
  AOI21_X1   g01548(.A1(new_n1646_), .A2(new_n1758_), .B(new_n1750_), .ZN(new_n1766_));
  OAI21_X1   g01549(.A1(new_n1647_), .A2(new_n1665_), .B(new_n1664_), .ZN(new_n1767_));
  INV_X1     g01550(.I(new_n1767_), .ZN(new_n1768_));
  INV_X1     g01551(.I(new_n1710_), .ZN(new_n1769_));
  NAND2_X1   g01552(.A1(\a[4] ), .A2(\a[22] ), .ZN(new_n1770_));
  NAND2_X1   g01553(.A1(new_n1770_), .A2(new_n242_), .ZN(new_n1771_));
  AOI21_X1   g01554(.A1(new_n1340_), .A2(new_n1769_), .B(new_n1771_), .ZN(new_n1772_));
  NAND2_X1   g01555(.A1(\a[21] ), .A2(\a[22] ), .ZN(new_n1773_));
  OR3_X2     g01556(.A1(new_n1772_), .A2(new_n212_), .A3(new_n1773_), .Z(new_n1774_));
  NOR2_X1    g01557(.A1(new_n242_), .A2(new_n1339_), .ZN(new_n1775_));
  AOI21_X1   g01558(.A1(\a[21] ), .A2(\a[22] ), .B(new_n267_), .ZN(new_n1776_));
  AOI21_X1   g01559(.A1(new_n1774_), .A2(new_n1775_), .B(new_n1776_), .ZN(new_n1777_));
  INV_X1     g01560(.I(new_n772_), .ZN(new_n1778_));
  NAND2_X1   g01561(.A1(new_n1778_), .A2(new_n609_), .ZN(new_n1779_));
  NAND2_X1   g01562(.A1(new_n1270_), .A2(new_n1779_), .ZN(new_n1780_));
  NOR2_X1    g01563(.A1(new_n453_), .A2(new_n1274_), .ZN(new_n1781_));
  AOI21_X1   g01564(.A1(\a[8] ), .A2(\a[17] ), .B(new_n1029_), .ZN(new_n1782_));
  OR3_X2     g01565(.A1(new_n1782_), .A2(new_n1004_), .A3(new_n1781_), .Z(new_n1783_));
  NOR2_X1    g01566(.A1(new_n1783_), .A2(new_n1780_), .ZN(new_n1784_));
  NAND2_X1   g01567(.A1(\a[10] ), .A2(\a[15] ), .ZN(new_n1785_));
  INV_X1     g01568(.I(new_n1785_), .ZN(new_n1786_));
  NAND2_X1   g01569(.A1(\a[23] ), .A2(\a[25] ), .ZN(new_n1787_));
  XNOR2_X1   g01570(.A1(new_n197_), .A2(new_n1787_), .ZN(new_n1788_));
  INV_X1     g01571(.I(new_n1788_), .ZN(new_n1789_));
  NAND2_X1   g01572(.A1(new_n1784_), .A2(new_n1789_), .ZN(new_n1790_));
  INV_X1     g01573(.I(new_n1790_), .ZN(new_n1791_));
  NOR2_X1    g01574(.A1(new_n1784_), .A2(new_n1789_), .ZN(new_n1792_));
  OAI21_X1   g01575(.A1(new_n1791_), .A2(new_n1792_), .B(new_n1777_), .ZN(new_n1793_));
  INV_X1     g01576(.I(new_n1777_), .ZN(new_n1794_));
  XOR2_X1    g01577(.A1(new_n1784_), .A2(new_n1789_), .Z(new_n1795_));
  NAND2_X1   g01578(.A1(new_n1795_), .A2(new_n1794_), .ZN(new_n1796_));
  NAND2_X1   g01579(.A1(new_n1796_), .A2(new_n1793_), .ZN(new_n1797_));
  INV_X1     g01580(.I(new_n1715_), .ZN(new_n1798_));
  AOI21_X1   g01581(.A1(new_n229_), .A2(new_n1798_), .B(new_n1714_), .ZN(new_n1799_));
  INV_X1     g01582(.I(new_n1687_), .ZN(new_n1800_));
  NAND2_X1   g01583(.A1(\a[1] ), .A2(\a[24] ), .ZN(new_n1801_));
  XOR2_X1    g01584(.A1(new_n1801_), .A2(\a[13] ), .Z(new_n1802_));
  XOR2_X1    g01585(.A1(new_n1802_), .A2(new_n1800_), .Z(new_n1803_));
  NAND2_X1   g01586(.A1(new_n1803_), .A2(new_n1799_), .ZN(new_n1804_));
  INV_X1     g01587(.I(new_n1799_), .ZN(new_n1805_));
  NOR2_X1    g01588(.A1(new_n1802_), .A2(new_n1800_), .ZN(new_n1806_));
  NAND2_X1   g01589(.A1(new_n1802_), .A2(new_n1800_), .ZN(new_n1807_));
  INV_X1     g01590(.I(new_n1807_), .ZN(new_n1808_));
  OAI21_X1   g01591(.A1(new_n1806_), .A2(new_n1808_), .B(new_n1805_), .ZN(new_n1809_));
  AOI21_X1   g01592(.A1(new_n1655_), .A2(new_n1652_), .B(new_n1539_), .ZN(new_n1810_));
  NOR2_X1    g01593(.A1(new_n1810_), .A2(new_n1656_), .ZN(new_n1811_));
  NAND2_X1   g01594(.A1(\a[11] ), .A2(\a[14] ), .ZN(new_n1812_));
  NOR2_X1    g01595(.A1(new_n1150_), .A2(new_n1812_), .ZN(new_n1813_));
  XOR2_X1    g01596(.A1(new_n1813_), .A2(new_n353_), .Z(new_n1814_));
  XOR2_X1    g01597(.A1(new_n1814_), .A2(\a[20] ), .Z(new_n1815_));
  INV_X1     g01598(.I(new_n1815_), .ZN(new_n1816_));
  NAND2_X1   g01599(.A1(new_n1816_), .A2(new_n1811_), .ZN(new_n1817_));
  INV_X1     g01600(.I(new_n1811_), .ZN(new_n1818_));
  NAND2_X1   g01601(.A1(new_n1818_), .A2(new_n1815_), .ZN(new_n1819_));
  AOI22_X1   g01602(.A1(new_n1817_), .A2(new_n1819_), .B1(new_n1804_), .B2(new_n1809_), .ZN(new_n1820_));
  NAND2_X1   g01603(.A1(new_n1809_), .A2(new_n1804_), .ZN(new_n1821_));
  NOR2_X1    g01604(.A1(new_n1815_), .A2(new_n1811_), .ZN(new_n1822_));
  INV_X1     g01605(.I(new_n1822_), .ZN(new_n1823_));
  NAND2_X1   g01606(.A1(new_n1815_), .A2(new_n1811_), .ZN(new_n1824_));
  AOI21_X1   g01607(.A1(new_n1823_), .A2(new_n1824_), .B(new_n1821_), .ZN(new_n1825_));
  OAI21_X1   g01608(.A1(new_n1820_), .A2(new_n1825_), .B(new_n1797_), .ZN(new_n1826_));
  INV_X1     g01609(.I(new_n1792_), .ZN(new_n1827_));
  AOI21_X1   g01610(.A1(new_n1827_), .A2(new_n1790_), .B(new_n1794_), .ZN(new_n1828_));
  AOI21_X1   g01611(.A1(new_n1795_), .A2(new_n1794_), .B(new_n1828_), .ZN(new_n1829_));
  NOR2_X1    g01612(.A1(new_n1820_), .A2(new_n1825_), .ZN(new_n1830_));
  NAND2_X1   g01613(.A1(new_n1830_), .A2(new_n1829_), .ZN(new_n1831_));
  AOI21_X1   g01614(.A1(new_n1831_), .A2(new_n1826_), .B(new_n1768_), .ZN(new_n1832_));
  NOR2_X1    g01615(.A1(new_n1830_), .A2(new_n1797_), .ZN(new_n1833_));
  NOR3_X1    g01616(.A1(new_n1829_), .A2(new_n1820_), .A3(new_n1825_), .ZN(new_n1834_));
  OAI21_X1   g01617(.A1(new_n1833_), .A2(new_n1834_), .B(new_n1768_), .ZN(new_n1835_));
  INV_X1     g01618(.I(new_n1835_), .ZN(new_n1836_));
  NOR2_X1    g01619(.A1(new_n1836_), .A2(new_n1832_), .ZN(new_n1837_));
  NAND2_X1   g01620(.A1(new_n1701_), .A2(new_n1699_), .ZN(new_n1838_));
  NAND2_X1   g01621(.A1(new_n1838_), .A2(new_n1700_), .ZN(new_n1839_));
  NAND3_X1   g01622(.A1(new_n1675_), .A2(\a[2] ), .A3(\a[6] ), .ZN(new_n1840_));
  OAI21_X1   g01623(.A1(new_n478_), .A2(new_n1268_), .B(new_n1840_), .ZN(new_n1841_));
  INV_X1     g01624(.I(new_n1841_), .ZN(new_n1842_));
  AOI21_X1   g01625(.A1(new_n597_), .A2(new_n1447_), .B(new_n1721_), .ZN(new_n1843_));
  NOR3_X1    g01626(.A1(new_n1686_), .A2(new_n1683_), .A3(new_n1687_), .ZN(new_n1844_));
  NAND2_X1   g01627(.A1(\a[0] ), .A2(\a[24] ), .ZN(new_n1845_));
  OAI21_X1   g01628(.A1(new_n1844_), .A2(new_n1845_), .B(new_n1688_), .ZN(new_n1846_));
  INV_X1     g01629(.I(new_n1846_), .ZN(new_n1847_));
  NOR2_X1    g01630(.A1(new_n1847_), .A2(new_n1843_), .ZN(new_n1848_));
  INV_X1     g01631(.I(new_n1843_), .ZN(new_n1849_));
  NOR2_X1    g01632(.A1(new_n1849_), .A2(new_n1846_), .ZN(new_n1850_));
  OAI21_X1   g01633(.A1(new_n1848_), .A2(new_n1850_), .B(new_n1842_), .ZN(new_n1851_));
  INV_X1     g01634(.I(new_n1851_), .ZN(new_n1852_));
  NAND2_X1   g01635(.A1(new_n1846_), .A2(new_n1843_), .ZN(new_n1853_));
  NOR2_X1    g01636(.A1(new_n1846_), .A2(new_n1843_), .ZN(new_n1854_));
  INV_X1     g01637(.I(new_n1854_), .ZN(new_n1855_));
  AOI21_X1   g01638(.A1(new_n1855_), .A2(new_n1853_), .B(new_n1842_), .ZN(new_n1856_));
  NOR2_X1    g01639(.A1(new_n1852_), .A2(new_n1856_), .ZN(new_n1857_));
  NAND2_X1   g01640(.A1(new_n1728_), .A2(new_n1726_), .ZN(new_n1858_));
  NAND2_X1   g01641(.A1(new_n1858_), .A2(new_n1727_), .ZN(new_n1859_));
  INV_X1     g01642(.I(new_n1859_), .ZN(new_n1860_));
  NOR2_X1    g01643(.A1(new_n1857_), .A2(new_n1860_), .ZN(new_n1861_));
  INV_X1     g01644(.I(new_n1856_), .ZN(new_n1862_));
  NAND2_X1   g01645(.A1(new_n1862_), .A2(new_n1851_), .ZN(new_n1863_));
  NOR2_X1    g01646(.A1(new_n1863_), .A2(new_n1859_), .ZN(new_n1864_));
  OAI21_X1   g01647(.A1(new_n1861_), .A2(new_n1864_), .B(new_n1839_), .ZN(new_n1865_));
  INV_X1     g01648(.I(new_n1700_), .ZN(new_n1866_));
  AOI21_X1   g01649(.A1(new_n1699_), .A2(new_n1701_), .B(new_n1866_), .ZN(new_n1867_));
  NAND2_X1   g01650(.A1(new_n1857_), .A2(new_n1859_), .ZN(new_n1868_));
  INV_X1     g01651(.I(new_n1868_), .ZN(new_n1869_));
  NOR2_X1    g01652(.A1(new_n1857_), .A2(new_n1859_), .ZN(new_n1870_));
  OAI21_X1   g01653(.A1(new_n1869_), .A2(new_n1870_), .B(new_n1867_), .ZN(new_n1871_));
  NAND2_X1   g01654(.A1(new_n1871_), .A2(new_n1865_), .ZN(new_n1872_));
  OAI21_X1   g01655(.A1(new_n1704_), .A2(new_n1731_), .B(new_n1742_), .ZN(new_n1873_));
  NAND2_X1   g01656(.A1(new_n1872_), .A2(new_n1873_), .ZN(new_n1874_));
  NAND2_X1   g01657(.A1(new_n1863_), .A2(new_n1859_), .ZN(new_n1875_));
  NAND2_X1   g01658(.A1(new_n1857_), .A2(new_n1860_), .ZN(new_n1876_));
  AOI21_X1   g01659(.A1(new_n1875_), .A2(new_n1876_), .B(new_n1867_), .ZN(new_n1877_));
  NAND2_X1   g01660(.A1(new_n1863_), .A2(new_n1860_), .ZN(new_n1878_));
  AOI21_X1   g01661(.A1(new_n1868_), .A2(new_n1878_), .B(new_n1839_), .ZN(new_n1879_));
  NOR2_X1    g01662(.A1(new_n1877_), .A2(new_n1879_), .ZN(new_n1880_));
  INV_X1     g01663(.I(new_n1873_), .ZN(new_n1881_));
  NAND2_X1   g01664(.A1(new_n1881_), .A2(new_n1880_), .ZN(new_n1882_));
  AOI21_X1   g01665(.A1(new_n1882_), .A2(new_n1874_), .B(new_n1837_), .ZN(new_n1883_));
  INV_X1     g01666(.I(new_n1883_), .ZN(new_n1884_));
  NAND2_X1   g01667(.A1(new_n1880_), .A2(new_n1873_), .ZN(new_n1885_));
  NAND2_X1   g01668(.A1(new_n1881_), .A2(new_n1872_), .ZN(new_n1886_));
  NAND2_X1   g01669(.A1(new_n1886_), .A2(new_n1885_), .ZN(new_n1887_));
  NAND2_X1   g01670(.A1(new_n1887_), .A2(new_n1837_), .ZN(new_n1888_));
  NAND2_X1   g01671(.A1(new_n1884_), .A2(new_n1888_), .ZN(new_n1889_));
  XNOR2_X1   g01672(.A1(new_n1889_), .A2(new_n1766_), .ZN(new_n1890_));
  NAND2_X1   g01673(.A1(new_n1889_), .A2(new_n1766_), .ZN(new_n1891_));
  INV_X1     g01674(.I(new_n1832_), .ZN(new_n1892_));
  NAND2_X1   g01675(.A1(new_n1892_), .A2(new_n1835_), .ZN(new_n1893_));
  AOI21_X1   g01676(.A1(new_n1886_), .A2(new_n1885_), .B(new_n1893_), .ZN(new_n1894_));
  NOR3_X1    g01677(.A1(new_n1883_), .A2(new_n1894_), .A3(new_n1766_), .ZN(new_n1895_));
  INV_X1     g01678(.I(new_n1895_), .ZN(new_n1896_));
  NAND2_X1   g01679(.A1(new_n1891_), .A2(new_n1896_), .ZN(new_n1897_));
  NAND2_X1   g01680(.A1(new_n1765_), .A2(new_n1897_), .ZN(new_n1898_));
  OAI21_X1   g01681(.A1(new_n1765_), .A2(new_n1890_), .B(new_n1898_), .ZN(\asquared[26] ));
  AOI21_X1   g01682(.A1(new_n1895_), .A2(new_n1752_), .B(new_n1761_), .ZN(new_n1900_));
  AOI21_X1   g01683(.A1(new_n1641_), .A2(new_n1637_), .B(new_n1900_), .ZN(new_n1901_));
  INV_X1     g01684(.I(new_n1885_), .ZN(new_n1902_));
  AOI21_X1   g01685(.A1(new_n1893_), .A2(new_n1886_), .B(new_n1902_), .ZN(new_n1903_));
  AOI21_X1   g01686(.A1(new_n1839_), .A2(new_n1878_), .B(new_n1869_), .ZN(new_n1904_));
  INV_X1     g01687(.I(new_n1904_), .ZN(new_n1905_));
  OAI21_X1   g01688(.A1(new_n1841_), .A2(new_n1854_), .B(new_n1853_), .ZN(new_n1906_));
  INV_X1     g01689(.I(new_n1906_), .ZN(new_n1907_));
  OAI21_X1   g01690(.A1(new_n1805_), .A2(new_n1806_), .B(new_n1807_), .ZN(new_n1908_));
  INV_X1     g01691(.I(new_n1908_), .ZN(new_n1909_));
  AOI21_X1   g01692(.A1(new_n1270_), .A2(new_n1779_), .B(new_n1781_), .ZN(new_n1910_));
  INV_X1     g01693(.I(new_n1910_), .ZN(new_n1911_));
  NAND2_X1   g01694(.A1(\a[23] ), .A2(\a[25] ), .ZN(new_n1912_));
  INV_X1     g01695(.I(new_n1912_), .ZN(new_n1913_));
  AOI21_X1   g01696(.A1(new_n218_), .A2(new_n1786_), .B(new_n1913_), .ZN(new_n1914_));
  INV_X1     g01697(.I(new_n1914_), .ZN(new_n1915_));
  INV_X1     g01698(.I(\a[26] ), .ZN(new_n1916_));
  NOR2_X1    g01699(.A1(new_n633_), .A2(new_n1691_), .ZN(new_n1917_));
  NOR2_X1    g01700(.A1(new_n359_), .A2(new_n1276_), .ZN(new_n1918_));
  NAND2_X1   g01701(.A1(new_n1917_), .A2(new_n1918_), .ZN(new_n1919_));
  XOR2_X1    g01702(.A1(new_n1919_), .A2(new_n199_), .Z(new_n1920_));
  NAND2_X1   g01703(.A1(new_n1920_), .A2(new_n1916_), .ZN(new_n1921_));
  XOR2_X1    g01704(.A1(new_n1919_), .A2(\a[0] ), .Z(new_n1922_));
  NAND2_X1   g01705(.A1(new_n1922_), .A2(\a[26] ), .ZN(new_n1923_));
  NAND2_X1   g01706(.A1(new_n1921_), .A2(new_n1923_), .ZN(new_n1924_));
  NAND2_X1   g01707(.A1(new_n1924_), .A2(new_n1915_), .ZN(new_n1925_));
  NOR2_X1    g01708(.A1(new_n1922_), .A2(\a[26] ), .ZN(new_n1926_));
  NOR2_X1    g01709(.A1(new_n1920_), .A2(new_n1916_), .ZN(new_n1927_));
  NOR2_X1    g01710(.A1(new_n1926_), .A2(new_n1927_), .ZN(new_n1928_));
  NAND2_X1   g01711(.A1(new_n1928_), .A2(new_n1914_), .ZN(new_n1929_));
  AOI21_X1   g01712(.A1(new_n1929_), .A2(new_n1925_), .B(new_n1911_), .ZN(new_n1930_));
  NAND2_X1   g01713(.A1(new_n1924_), .A2(new_n1914_), .ZN(new_n1931_));
  NAND2_X1   g01714(.A1(new_n1928_), .A2(new_n1915_), .ZN(new_n1932_));
  AOI21_X1   g01715(.A1(new_n1932_), .A2(new_n1931_), .B(new_n1910_), .ZN(new_n1933_));
  OAI21_X1   g01716(.A1(new_n1933_), .A2(new_n1930_), .B(new_n1909_), .ZN(new_n1934_));
  NOR2_X1    g01717(.A1(new_n1928_), .A2(new_n1914_), .ZN(new_n1935_));
  NOR2_X1    g01718(.A1(new_n1924_), .A2(new_n1915_), .ZN(new_n1936_));
  OAI21_X1   g01719(.A1(new_n1935_), .A2(new_n1936_), .B(new_n1910_), .ZN(new_n1937_));
  NOR2_X1    g01720(.A1(new_n1928_), .A2(new_n1915_), .ZN(new_n1938_));
  NOR2_X1    g01721(.A1(new_n1924_), .A2(new_n1914_), .ZN(new_n1939_));
  OAI21_X1   g01722(.A1(new_n1938_), .A2(new_n1939_), .B(new_n1911_), .ZN(new_n1940_));
  NAND3_X1   g01723(.A1(new_n1937_), .A2(new_n1940_), .A3(new_n1908_), .ZN(new_n1941_));
  AOI21_X1   g01724(.A1(new_n1934_), .A2(new_n1941_), .B(new_n1907_), .ZN(new_n1942_));
  OAI21_X1   g01725(.A1(new_n1933_), .A2(new_n1930_), .B(new_n1908_), .ZN(new_n1943_));
  NAND3_X1   g01726(.A1(new_n1937_), .A2(new_n1940_), .A3(new_n1909_), .ZN(new_n1944_));
  AOI21_X1   g01727(.A1(new_n1943_), .A2(new_n1944_), .B(new_n1906_), .ZN(new_n1945_));
  NAND2_X1   g01728(.A1(\a[4] ), .A2(\a[6] ), .ZN(new_n1948_));
  NAND2_X1   g01729(.A1(\a[20] ), .A2(\a[22] ), .ZN(new_n1949_));
  NOR2_X1    g01730(.A1(new_n481_), .A2(new_n1711_), .ZN(new_n1953_));
  INV_X1     g01731(.I(new_n1953_), .ZN(new_n1954_));
  NAND2_X1   g01732(.A1(\a[19] ), .A2(\a[24] ), .ZN(new_n1955_));
  NAND2_X1   g01733(.A1(\a[23] ), .A2(\a[24] ), .ZN(new_n1956_));
  OAI22_X1   g01734(.A1(new_n225_), .A2(new_n264_), .B1(new_n1955_), .B2(new_n1956_), .ZN(new_n1957_));
  INV_X1     g01735(.I(new_n1957_), .ZN(new_n1958_));
  NAND2_X1   g01736(.A1(\a[3] ), .A2(\a[23] ), .ZN(new_n1959_));
  INV_X1     g01737(.I(new_n1959_), .ZN(new_n1960_));
  NAND2_X1   g01738(.A1(\a[7] ), .A2(\a[19] ), .ZN(new_n1961_));
  OAI21_X1   g01739(.A1(new_n1960_), .A2(new_n1961_), .B(new_n1958_), .ZN(new_n1962_));
  XNOR2_X1   g01740(.A1(new_n1959_), .A2(new_n1961_), .ZN(new_n1963_));
  OAI21_X1   g01741(.A1(new_n201_), .A2(new_n1691_), .B(new_n1963_), .ZN(new_n1964_));
  NAND2_X1   g01742(.A1(\a[9] ), .A2(\a[17] ), .ZN(new_n1965_));
  OAI22_X1   g01743(.A1(new_n525_), .A2(new_n1965_), .B1(new_n868_), .B2(new_n1274_), .ZN(new_n1966_));
  NOR2_X1    g01744(.A1(new_n796_), .A2(new_n1021_), .ZN(new_n1967_));
  INV_X1     g01745(.I(new_n868_), .ZN(new_n1968_));
  AOI21_X1   g01746(.A1(\a[10] ), .A2(\a[16] ), .B(new_n1968_), .ZN(new_n1969_));
  NOR4_X1    g01747(.A1(new_n1969_), .A2(new_n1965_), .A3(new_n1966_), .A4(new_n1967_), .ZN(new_n1970_));
  NAND3_X1   g01748(.A1(new_n1964_), .A2(new_n1962_), .A3(new_n1970_), .ZN(new_n1971_));
  NAND2_X1   g01749(.A1(new_n1964_), .A2(new_n1962_), .ZN(new_n1972_));
  INV_X1     g01750(.I(new_n1970_), .ZN(new_n1973_));
  NAND2_X1   g01751(.A1(new_n1972_), .A2(new_n1973_), .ZN(new_n1974_));
  AOI21_X1   g01752(.A1(new_n1974_), .A2(new_n1971_), .B(new_n1954_), .ZN(new_n1975_));
  XOR2_X1    g01753(.A1(new_n1972_), .A2(new_n1970_), .Z(new_n1976_));
  NOR2_X1    g01754(.A1(new_n1976_), .A2(new_n1953_), .ZN(new_n1977_));
  NOR2_X1    g01755(.A1(new_n1977_), .A2(new_n1975_), .ZN(new_n1978_));
  NOR3_X1    g01756(.A1(new_n1942_), .A2(new_n1945_), .A3(new_n1978_), .ZN(new_n1979_));
  INV_X1     g01757(.I(new_n1934_), .ZN(new_n1980_));
  NOR3_X1    g01758(.A1(new_n1933_), .A2(new_n1930_), .A3(new_n1909_), .ZN(new_n1981_));
  OAI21_X1   g01759(.A1(new_n1980_), .A2(new_n1981_), .B(new_n1906_), .ZN(new_n1982_));
  AOI21_X1   g01760(.A1(new_n1940_), .A2(new_n1937_), .B(new_n1909_), .ZN(new_n1983_));
  NOR3_X1    g01761(.A1(new_n1933_), .A2(new_n1930_), .A3(new_n1908_), .ZN(new_n1984_));
  OAI21_X1   g01762(.A1(new_n1983_), .A2(new_n1984_), .B(new_n1907_), .ZN(new_n1985_));
  INV_X1     g01763(.I(new_n1978_), .ZN(new_n1986_));
  AOI21_X1   g01764(.A1(new_n1982_), .A2(new_n1985_), .B(new_n1986_), .ZN(new_n1987_));
  OAI21_X1   g01765(.A1(new_n1987_), .A2(new_n1979_), .B(new_n1905_), .ZN(new_n1988_));
  AOI21_X1   g01766(.A1(new_n1982_), .A2(new_n1985_), .B(new_n1978_), .ZN(new_n1989_));
  NOR3_X1    g01767(.A1(new_n1942_), .A2(new_n1945_), .A3(new_n1986_), .ZN(new_n1990_));
  OAI21_X1   g01768(.A1(new_n1989_), .A2(new_n1990_), .B(new_n1904_), .ZN(new_n1991_));
  NAND2_X1   g01769(.A1(new_n1988_), .A2(new_n1991_), .ZN(new_n1992_));
  INV_X1     g01770(.I(new_n1826_), .ZN(new_n1993_));
  AOI21_X1   g01771(.A1(new_n1767_), .A2(new_n1831_), .B(new_n1993_), .ZN(new_n1994_));
  OAI21_X1   g01772(.A1(new_n1794_), .A2(new_n1792_), .B(new_n1790_), .ZN(new_n1995_));
  INV_X1     g01773(.I(new_n1824_), .ZN(new_n1996_));
  NOR2_X1    g01774(.A1(new_n1996_), .A2(new_n1821_), .ZN(new_n1997_));
  NOR2_X1    g01775(.A1(new_n1997_), .A2(new_n1822_), .ZN(new_n1998_));
  INV_X1     g01776(.I(\a[25] ), .ZN(new_n1999_));
  NOR2_X1    g01777(.A1(new_n194_), .A2(new_n1999_), .ZN(new_n2000_));
  NAND2_X1   g01778(.A1(\a[5] ), .A2(\a[20] ), .ZN(new_n2001_));
  AOI21_X1   g01779(.A1(new_n1150_), .A2(new_n1812_), .B(new_n2001_), .ZN(new_n2002_));
  NOR2_X1    g01780(.A1(new_n2002_), .A2(new_n1813_), .ZN(new_n2003_));
  NOR3_X1    g01781(.A1(new_n212_), .A2(new_n1313_), .A3(new_n1674_), .ZN(new_n2004_));
  XOR2_X1    g01782(.A1(new_n2004_), .A2(new_n653_), .Z(new_n2005_));
  XOR2_X1    g01783(.A1(new_n2005_), .A2(new_n2003_), .Z(new_n2006_));
  XOR2_X1    g01784(.A1(new_n2006_), .A2(new_n2000_), .Z(new_n2007_));
  NOR2_X1    g01785(.A1(new_n1998_), .A2(new_n2007_), .ZN(new_n2008_));
  OAI21_X1   g01786(.A1(new_n1821_), .A2(new_n1996_), .B(new_n1823_), .ZN(new_n2009_));
  INV_X1     g01787(.I(new_n2007_), .ZN(new_n2010_));
  NOR2_X1    g01788(.A1(new_n2009_), .A2(new_n2010_), .ZN(new_n2011_));
  OAI21_X1   g01789(.A1(new_n2008_), .A2(new_n2011_), .B(new_n1995_), .ZN(new_n2012_));
  INV_X1     g01790(.I(new_n1995_), .ZN(new_n2013_));
  NOR2_X1    g01791(.A1(new_n2009_), .A2(new_n2007_), .ZN(new_n2014_));
  NOR2_X1    g01792(.A1(new_n1998_), .A2(new_n2010_), .ZN(new_n2015_));
  OAI21_X1   g01793(.A1(new_n2015_), .A2(new_n2014_), .B(new_n2013_), .ZN(new_n2016_));
  NAND2_X1   g01794(.A1(new_n2012_), .A2(new_n2016_), .ZN(new_n2017_));
  NAND2_X1   g01795(.A1(new_n2017_), .A2(new_n1994_), .ZN(new_n2018_));
  INV_X1     g01796(.I(new_n2018_), .ZN(new_n2019_));
  NOR2_X1    g01797(.A1(new_n2017_), .A2(new_n1994_), .ZN(new_n2020_));
  NOR2_X1    g01798(.A1(new_n2019_), .A2(new_n2020_), .ZN(new_n2021_));
  XNOR2_X1   g01799(.A1(new_n2017_), .A2(new_n1994_), .ZN(new_n2022_));
  MUX2_X1    g01800(.I0(new_n2022_), .I1(new_n2021_), .S(new_n1992_), .Z(new_n2023_));
  NOR2_X1    g01801(.A1(new_n2023_), .A2(new_n1903_), .ZN(new_n2024_));
  XNOR2_X1   g01802(.A1(new_n1901_), .A2(new_n2024_), .ZN(new_n2025_));
  XOR2_X1    g01803(.A1(new_n2025_), .A2(new_n1891_), .Z(\asquared[27] ));
  NOR2_X1    g01804(.A1(new_n1891_), .A2(new_n1903_), .ZN(new_n2027_));
  AOI21_X1   g01805(.A1(new_n1891_), .A2(new_n1903_), .B(new_n2023_), .ZN(new_n2028_));
  AOI21_X1   g01806(.A1(new_n1901_), .A2(new_n2028_), .B(new_n2027_), .ZN(new_n2029_));
  AOI21_X1   g01807(.A1(new_n1992_), .A2(new_n2018_), .B(new_n2020_), .ZN(new_n2030_));
  OAI21_X1   g01808(.A1(new_n1942_), .A2(new_n1945_), .B(new_n1978_), .ZN(new_n2031_));
  AOI21_X1   g01809(.A1(new_n1905_), .A2(new_n2031_), .B(new_n1979_), .ZN(new_n2032_));
  NOR2_X1    g01810(.A1(new_n2014_), .A2(new_n2013_), .ZN(new_n2033_));
  NOR2_X1    g01811(.A1(new_n2033_), .A2(new_n2015_), .ZN(new_n2034_));
  NOR2_X1    g01812(.A1(new_n2003_), .A2(new_n2004_), .ZN(new_n2035_));
  NAND2_X1   g01813(.A1(new_n2003_), .A2(new_n2004_), .ZN(new_n2036_));
  XOR2_X1    g01814(.A1(new_n2000_), .A2(new_n653_), .Z(new_n2037_));
  INV_X1     g01815(.I(new_n2037_), .ZN(new_n2038_));
  AOI21_X1   g01816(.A1(new_n2038_), .A2(new_n2036_), .B(new_n2035_), .ZN(new_n2039_));
  NAND2_X1   g01817(.A1(new_n1974_), .A2(new_n1953_), .ZN(new_n2040_));
  NAND2_X1   g01818(.A1(new_n2040_), .A2(new_n1971_), .ZN(new_n2041_));
  INV_X1     g01819(.I(new_n2041_), .ZN(new_n2042_));
  OAI21_X1   g01820(.A1(new_n1911_), .A2(new_n1936_), .B(new_n1925_), .ZN(new_n2043_));
  NAND2_X1   g01821(.A1(new_n2043_), .A2(new_n2042_), .ZN(new_n2044_));
  AOI21_X1   g01822(.A1(new_n1928_), .A2(new_n1914_), .B(new_n1911_), .ZN(new_n2045_));
  NOR2_X1    g01823(.A1(new_n2045_), .A2(new_n1935_), .ZN(new_n2046_));
  NAND2_X1   g01824(.A1(new_n2046_), .A2(new_n2041_), .ZN(new_n2047_));
  AOI21_X1   g01825(.A1(new_n2044_), .A2(new_n2047_), .B(new_n2039_), .ZN(new_n2048_));
  INV_X1     g01826(.I(new_n2039_), .ZN(new_n2049_));
  NAND2_X1   g01827(.A1(new_n2043_), .A2(new_n2041_), .ZN(new_n2050_));
  NOR3_X1    g01828(.A1(new_n2041_), .A2(new_n2045_), .A3(new_n1935_), .ZN(new_n2051_));
  INV_X1     g01829(.I(new_n2051_), .ZN(new_n2052_));
  AOI21_X1   g01830(.A1(new_n2052_), .A2(new_n2050_), .B(new_n2049_), .ZN(new_n2053_));
  NAND2_X1   g01831(.A1(\a[7] ), .A2(\a[25] ), .ZN(new_n2054_));
  XNOR2_X1   g01832(.A1(new_n1597_), .A2(new_n2054_), .ZN(new_n2055_));
  INV_X1     g01833(.I(new_n2055_), .ZN(new_n2056_));
  NOR2_X1    g01834(.A1(new_n199_), .A2(new_n1916_), .ZN(new_n2057_));
  OAI21_X1   g01835(.A1(new_n1917_), .A2(new_n1918_), .B(new_n2057_), .ZN(new_n2058_));
  NAND2_X1   g01836(.A1(new_n2058_), .A2(new_n1919_), .ZN(new_n2059_));
  NOR2_X1    g01837(.A1(new_n359_), .A2(new_n1339_), .ZN(new_n2060_));
  NOR2_X1    g01838(.A1(new_n525_), .A2(new_n1268_), .ZN(new_n2061_));
  NOR2_X1    g01839(.A1(new_n461_), .A2(new_n885_), .ZN(new_n2062_));
  NOR2_X1    g01840(.A1(new_n525_), .A2(new_n1268_), .ZN(new_n2065_));
  NAND2_X1   g01841(.A1(\a[11] ), .A2(\a[16] ), .ZN(new_n2066_));
  XOR2_X1    g01842(.A1(new_n2065_), .A2(new_n2066_), .Z(new_n2067_));
  XOR2_X1    g01843(.A1(new_n2067_), .A2(new_n2059_), .Z(new_n2068_));
  XOR2_X1    g01844(.A1(new_n2068_), .A2(new_n2056_), .Z(new_n2069_));
  INV_X1     g01845(.I(new_n2069_), .ZN(new_n2070_));
  OAI21_X1   g01846(.A1(new_n2053_), .A2(new_n2048_), .B(new_n2070_), .ZN(new_n2071_));
  NOR2_X1    g01847(.A1(new_n2046_), .A2(new_n2041_), .ZN(new_n2072_));
  NOR2_X1    g01848(.A1(new_n2043_), .A2(new_n2042_), .ZN(new_n2073_));
  OAI21_X1   g01849(.A1(new_n2073_), .A2(new_n2072_), .B(new_n2049_), .ZN(new_n2074_));
  NOR2_X1    g01850(.A1(new_n2042_), .A2(new_n2046_), .ZN(new_n2075_));
  OAI21_X1   g01851(.A1(new_n2075_), .A2(new_n2051_), .B(new_n2039_), .ZN(new_n2076_));
  NAND3_X1   g01852(.A1(new_n2074_), .A2(new_n2076_), .A3(new_n2069_), .ZN(new_n2077_));
  AOI21_X1   g01853(.A1(new_n2071_), .A2(new_n2077_), .B(new_n2034_), .ZN(new_n2078_));
  NAND2_X1   g01854(.A1(new_n2009_), .A2(new_n2007_), .ZN(new_n2079_));
  OAI21_X1   g01855(.A1(new_n2013_), .A2(new_n2014_), .B(new_n2079_), .ZN(new_n2080_));
  NAND3_X1   g01856(.A1(new_n2074_), .A2(new_n2076_), .A3(new_n2070_), .ZN(new_n2081_));
  OAI21_X1   g01857(.A1(new_n2053_), .A2(new_n2048_), .B(new_n2069_), .ZN(new_n2082_));
  AOI21_X1   g01858(.A1(new_n2082_), .A2(new_n2081_), .B(new_n2080_), .ZN(new_n2083_));
  NOR2_X1    g01859(.A1(new_n2078_), .A2(new_n2083_), .ZN(new_n2084_));
  OAI21_X1   g01860(.A1(new_n1907_), .A2(new_n1984_), .B(new_n1943_), .ZN(new_n2085_));
  NOR4_X1    g01861(.A1(new_n200_), .A2(new_n242_), .A3(new_n1313_), .A4(new_n1691_), .ZN(new_n2086_));
  NAND4_X1   g01862(.A1(new_n2086_), .A2(\a[4] ), .A3(\a[6] ), .A4(new_n1707_), .ZN(new_n2087_));
  AOI21_X1   g01863(.A1(new_n2087_), .A2(new_n212_), .B(new_n1956_), .ZN(new_n2088_));
  NAND2_X1   g01864(.A1(\a[3] ), .A2(\a[24] ), .ZN(new_n2089_));
  OAI22_X1   g01865(.A1(new_n212_), .A2(new_n1956_), .B1(new_n1948_), .B2(new_n1706_), .ZN(new_n2090_));
  NAND2_X1   g01866(.A1(new_n1948_), .A2(new_n1706_), .ZN(new_n2091_));
  OAI22_X1   g01867(.A1(new_n2088_), .A2(new_n2089_), .B1(new_n2090_), .B2(new_n2091_), .ZN(new_n2092_));
  INV_X1     g01868(.I(new_n2092_), .ZN(new_n2093_));
  AOI21_X1   g01869(.A1(\a[12] ), .A2(\a[15] ), .B(new_n787_), .ZN(new_n2094_));
  NAND3_X1   g01870(.A1(new_n2094_), .A2(new_n1220_), .A3(new_n1447_), .ZN(new_n2095_));
  NOR2_X1    g01871(.A1(new_n353_), .A2(new_n1674_), .ZN(new_n2096_));
  XOR2_X1    g01872(.A1(new_n2095_), .A2(new_n2096_), .Z(new_n2097_));
  INV_X1     g01873(.I(\a[27] ), .ZN(new_n2098_));
  NAND2_X1   g01874(.A1(new_n2000_), .A2(new_n654_), .ZN(new_n2099_));
  AOI21_X1   g01875(.A1(\a[1] ), .A2(\a[26] ), .B(\a[14] ), .ZN(new_n2100_));
  NOR2_X1    g01876(.A1(new_n681_), .A2(new_n1916_), .ZN(new_n2101_));
  NOR2_X1    g01877(.A1(new_n2101_), .A2(new_n2100_), .ZN(new_n2102_));
  NOR2_X1    g01878(.A1(new_n2102_), .A2(new_n2099_), .ZN(new_n2103_));
  XOR2_X1    g01879(.A1(new_n2103_), .A2(new_n199_), .Z(new_n2104_));
  XOR2_X1    g01880(.A1(new_n2104_), .A2(new_n2098_), .Z(new_n2105_));
  NAND2_X1   g01881(.A1(new_n2105_), .A2(new_n2097_), .ZN(new_n2106_));
  INV_X1     g01882(.I(new_n2106_), .ZN(new_n2107_));
  NOR2_X1    g01883(.A1(new_n2105_), .A2(new_n2097_), .ZN(new_n2108_));
  OAI21_X1   g01884(.A1(new_n2107_), .A2(new_n2108_), .B(new_n2093_), .ZN(new_n2109_));
  INV_X1     g01885(.I(new_n2097_), .ZN(new_n2110_));
  NAND2_X1   g01886(.A1(new_n2105_), .A2(new_n2110_), .ZN(new_n2111_));
  INV_X1     g01887(.I(new_n2111_), .ZN(new_n2112_));
  NOR2_X1    g01888(.A1(new_n2105_), .A2(new_n2110_), .ZN(new_n2113_));
  OAI21_X1   g01889(.A1(new_n2112_), .A2(new_n2113_), .B(new_n2092_), .ZN(new_n2114_));
  OAI22_X1   g01890(.A1(new_n211_), .A2(new_n1773_), .B1(new_n481_), .B2(new_n1711_), .ZN(new_n2115_));
  OAI21_X1   g01891(.A1(new_n1959_), .A2(new_n1961_), .B(new_n1957_), .ZN(new_n2116_));
  OAI21_X1   g01892(.A1(new_n796_), .A2(new_n1021_), .B(new_n1966_), .ZN(new_n2117_));
  XNOR2_X1   g01893(.A1(new_n2116_), .A2(new_n2117_), .ZN(new_n2118_));
  NOR2_X1    g01894(.A1(new_n2118_), .A2(new_n2115_), .ZN(new_n2119_));
  INV_X1     g01895(.I(new_n2115_), .ZN(new_n2120_));
  NOR2_X1    g01896(.A1(new_n2116_), .A2(new_n2117_), .ZN(new_n2121_));
  INV_X1     g01897(.I(new_n2121_), .ZN(new_n2122_));
  NAND2_X1   g01898(.A1(new_n2116_), .A2(new_n2117_), .ZN(new_n2123_));
  AOI21_X1   g01899(.A1(new_n2122_), .A2(new_n2123_), .B(new_n2120_), .ZN(new_n2124_));
  NOR2_X1    g01900(.A1(new_n2119_), .A2(new_n2124_), .ZN(new_n2125_));
  AOI21_X1   g01901(.A1(new_n2109_), .A2(new_n2114_), .B(new_n2125_), .ZN(new_n2126_));
  INV_X1     g01902(.I(new_n2108_), .ZN(new_n2127_));
  AOI21_X1   g01903(.A1(new_n2127_), .A2(new_n2106_), .B(new_n2092_), .ZN(new_n2128_));
  OR2_X2     g01904(.A1(new_n2105_), .A2(new_n2110_), .Z(new_n2129_));
  AOI21_X1   g01905(.A1(new_n2129_), .A2(new_n2111_), .B(new_n2093_), .ZN(new_n2130_));
  INV_X1     g01906(.I(new_n2125_), .ZN(new_n2131_));
  NOR3_X1    g01907(.A1(new_n2128_), .A2(new_n2130_), .A3(new_n2131_), .ZN(new_n2132_));
  OAI21_X1   g01908(.A1(new_n2126_), .A2(new_n2132_), .B(new_n2085_), .ZN(new_n2133_));
  AOI21_X1   g01909(.A1(new_n1906_), .A2(new_n1944_), .B(new_n1983_), .ZN(new_n2134_));
  NOR3_X1    g01910(.A1(new_n2128_), .A2(new_n2130_), .A3(new_n2125_), .ZN(new_n2135_));
  AOI21_X1   g01911(.A1(new_n2109_), .A2(new_n2114_), .B(new_n2131_), .ZN(new_n2136_));
  OAI21_X1   g01912(.A1(new_n2136_), .A2(new_n2135_), .B(new_n2134_), .ZN(new_n2137_));
  NAND2_X1   g01913(.A1(new_n2137_), .A2(new_n2133_), .ZN(new_n2138_));
  NAND2_X1   g01914(.A1(new_n2084_), .A2(new_n2138_), .ZN(new_n2139_));
  AOI21_X1   g01915(.A1(new_n2074_), .A2(new_n2076_), .B(new_n2069_), .ZN(new_n2140_));
  NOR3_X1    g01916(.A1(new_n2053_), .A2(new_n2048_), .A3(new_n2070_), .ZN(new_n2141_));
  OAI21_X1   g01917(.A1(new_n2141_), .A2(new_n2140_), .B(new_n2080_), .ZN(new_n2142_));
  NOR3_X1    g01918(.A1(new_n2053_), .A2(new_n2048_), .A3(new_n2069_), .ZN(new_n2143_));
  AOI21_X1   g01919(.A1(new_n2074_), .A2(new_n2076_), .B(new_n2070_), .ZN(new_n2144_));
  OAI21_X1   g01920(.A1(new_n2143_), .A2(new_n2144_), .B(new_n2034_), .ZN(new_n2145_));
  NAND2_X1   g01921(.A1(new_n2145_), .A2(new_n2142_), .ZN(new_n2146_));
  OAI21_X1   g01922(.A1(new_n2128_), .A2(new_n2130_), .B(new_n2131_), .ZN(new_n2147_));
  NAND3_X1   g01923(.A1(new_n2109_), .A2(new_n2114_), .A3(new_n2125_), .ZN(new_n2148_));
  AOI21_X1   g01924(.A1(new_n2147_), .A2(new_n2148_), .B(new_n2134_), .ZN(new_n2149_));
  NAND3_X1   g01925(.A1(new_n2109_), .A2(new_n2114_), .A3(new_n2131_), .ZN(new_n2150_));
  OAI21_X1   g01926(.A1(new_n2128_), .A2(new_n2130_), .B(new_n2125_), .ZN(new_n2151_));
  AOI21_X1   g01927(.A1(new_n2151_), .A2(new_n2150_), .B(new_n2085_), .ZN(new_n2152_));
  NOR2_X1    g01928(.A1(new_n2149_), .A2(new_n2152_), .ZN(new_n2153_));
  NAND2_X1   g01929(.A1(new_n2146_), .A2(new_n2153_), .ZN(new_n2154_));
  AOI21_X1   g01930(.A1(new_n2139_), .A2(new_n2154_), .B(new_n2032_), .ZN(new_n2155_));
  NAND3_X1   g01931(.A1(new_n1982_), .A2(new_n1985_), .A3(new_n1986_), .ZN(new_n2156_));
  OAI21_X1   g01932(.A1(new_n1904_), .A2(new_n1987_), .B(new_n2156_), .ZN(new_n2157_));
  NAND2_X1   g01933(.A1(new_n2146_), .A2(new_n2138_), .ZN(new_n2158_));
  NAND2_X1   g01934(.A1(new_n2084_), .A2(new_n2153_), .ZN(new_n2159_));
  AOI21_X1   g01935(.A1(new_n2158_), .A2(new_n2159_), .B(new_n2157_), .ZN(new_n2160_));
  NOR2_X1    g01936(.A1(new_n2155_), .A2(new_n2160_), .ZN(new_n2161_));
  XOR2_X1    g01937(.A1(new_n2161_), .A2(new_n2030_), .Z(new_n2162_));
  OAI21_X1   g01938(.A1(new_n2155_), .A2(new_n2160_), .B(new_n2030_), .ZN(new_n2163_));
  INV_X1     g01939(.I(new_n2030_), .ZN(new_n2164_));
  NAND2_X1   g01940(.A1(new_n2161_), .A2(new_n2164_), .ZN(new_n2165_));
  NAND2_X1   g01941(.A1(new_n2165_), .A2(new_n2163_), .ZN(new_n2166_));
  NAND2_X1   g01942(.A1(new_n2029_), .A2(new_n2166_), .ZN(new_n2167_));
  OAI21_X1   g01943(.A1(new_n2029_), .A2(new_n2162_), .B(new_n2167_), .ZN(\asquared[28] ));
  NOR2_X1    g01944(.A1(new_n2161_), .A2(new_n2164_), .ZN(new_n2169_));
  OAI21_X1   g01945(.A1(new_n2029_), .A2(new_n2169_), .B(new_n2165_), .ZN(new_n2170_));
  NOR2_X1    g01946(.A1(new_n2146_), .A2(new_n2138_), .ZN(new_n2171_));
  AOI21_X1   g01947(.A1(new_n2146_), .A2(new_n2138_), .B(new_n2032_), .ZN(new_n2172_));
  OAI21_X1   g01948(.A1(new_n2034_), .A2(new_n2144_), .B(new_n2081_), .ZN(new_n2173_));
  OAI21_X1   g01949(.A1(new_n2043_), .A2(new_n2041_), .B(new_n2049_), .ZN(new_n2174_));
  NAND2_X1   g01950(.A1(new_n2174_), .A2(new_n2050_), .ZN(new_n2175_));
  NAND2_X1   g01951(.A1(\a[16] ), .A2(\a[28] ), .ZN(new_n2176_));
  INV_X1     g01952(.I(new_n2176_), .ZN(new_n2177_));
  INV_X1     g01953(.I(\a[28] ), .ZN(new_n2178_));
  NOR2_X1    g01954(.A1(new_n675_), .A2(new_n2178_), .ZN(new_n2179_));
  INV_X1     g01955(.I(new_n2179_), .ZN(new_n2180_));
  NOR3_X1    g01956(.A1(new_n2180_), .A2(new_n199_), .A3(new_n885_), .ZN(new_n2181_));
  NAND4_X1   g01957(.A1(new_n2181_), .A2(\a[0] ), .A3(\a[12] ), .A4(new_n2177_), .ZN(new_n2182_));
  AOI21_X1   g01958(.A1(new_n2182_), .A2(new_n1274_), .B(new_n651_), .ZN(new_n2183_));
  NAND2_X1   g01959(.A1(\a[11] ), .A2(\a[17] ), .ZN(new_n2184_));
  OAI22_X1   g01960(.A1(new_n527_), .A2(new_n2176_), .B1(new_n651_), .B2(new_n1274_), .ZN(new_n2185_));
  NAND2_X1   g01961(.A1(new_n527_), .A2(new_n2176_), .ZN(new_n2186_));
  OAI22_X1   g01962(.A1(new_n2183_), .A2(new_n2184_), .B1(new_n2185_), .B2(new_n2186_), .ZN(new_n2187_));
  AOI21_X1   g01963(.A1(new_n2116_), .A2(new_n2117_), .B(new_n2115_), .ZN(new_n2188_));
  NOR2_X1    g01964(.A1(new_n2188_), .A2(new_n2121_), .ZN(new_n2189_));
  NAND2_X1   g01965(.A1(\a[2] ), .A2(\a[26] ), .ZN(new_n2190_));
  INV_X1     g01966(.I(new_n2190_), .ZN(new_n2191_));
  XNOR2_X1   g01967(.A1(new_n525_), .A2(new_n1342_), .ZN(new_n2192_));
  INV_X1     g01968(.I(new_n2192_), .ZN(new_n2193_));
  NAND2_X1   g01969(.A1(new_n2189_), .A2(new_n2193_), .ZN(new_n2194_));
  INV_X1     g01970(.I(new_n2189_), .ZN(new_n2195_));
  NAND2_X1   g01971(.A1(new_n2195_), .A2(new_n2192_), .ZN(new_n2196_));
  AOI21_X1   g01972(.A1(new_n2196_), .A2(new_n2194_), .B(new_n2187_), .ZN(new_n2197_));
  INV_X1     g01973(.I(new_n2197_), .ZN(new_n2198_));
  NOR2_X1    g01974(.A1(new_n2189_), .A2(new_n2192_), .ZN(new_n2199_));
  NAND2_X1   g01975(.A1(new_n2189_), .A2(new_n2192_), .ZN(new_n2200_));
  INV_X1     g01976(.I(new_n2200_), .ZN(new_n2201_));
  OAI21_X1   g01977(.A1(new_n2201_), .A2(new_n2199_), .B(new_n2187_), .ZN(new_n2202_));
  NAND2_X1   g01978(.A1(new_n2198_), .A2(new_n2202_), .ZN(new_n2203_));
  INV_X1     g01979(.I(new_n2061_), .ZN(new_n2204_));
  OAI21_X1   g01980(.A1(new_n453_), .A2(new_n1342_), .B(new_n2204_), .ZN(new_n2205_));
  INV_X1     g01981(.I(new_n2090_), .ZN(new_n2206_));
  NAND3_X1   g01982(.A1(new_n344_), .A2(\a[20] ), .A3(\a[25] ), .ZN(new_n2207_));
  OAI21_X1   g01983(.A1(new_n2055_), .A2(new_n2066_), .B(new_n2207_), .ZN(new_n2208_));
  XOR2_X1    g01984(.A1(new_n2208_), .A2(new_n2206_), .Z(new_n2209_));
  NOR2_X1    g01985(.A1(new_n2209_), .A2(new_n2205_), .ZN(new_n2210_));
  INV_X1     g01986(.I(new_n2205_), .ZN(new_n2211_));
  OR2_X2     g01987(.A1(new_n2208_), .A2(new_n2090_), .Z(new_n2212_));
  NAND2_X1   g01988(.A1(new_n2208_), .A2(new_n2090_), .ZN(new_n2213_));
  AOI21_X1   g01989(.A1(new_n2212_), .A2(new_n2213_), .B(new_n2211_), .ZN(new_n2214_));
  NOR2_X1    g01990(.A1(new_n2210_), .A2(new_n2214_), .ZN(new_n2215_));
  NOR2_X1    g01991(.A1(new_n2203_), .A2(new_n2215_), .ZN(new_n2216_));
  INV_X1     g01992(.I(new_n2202_), .ZN(new_n2217_));
  NOR2_X1    g01993(.A1(new_n2217_), .A2(new_n2197_), .ZN(new_n2218_));
  INV_X1     g01994(.I(new_n2215_), .ZN(new_n2219_));
  NOR2_X1    g01995(.A1(new_n2218_), .A2(new_n2219_), .ZN(new_n2220_));
  OAI21_X1   g01996(.A1(new_n2220_), .A2(new_n2216_), .B(new_n2175_), .ZN(new_n2221_));
  AOI21_X1   g01997(.A1(new_n2049_), .A2(new_n2052_), .B(new_n2075_), .ZN(new_n2222_));
  NOR2_X1    g01998(.A1(new_n2218_), .A2(new_n2215_), .ZN(new_n2223_));
  NOR2_X1    g01999(.A1(new_n2203_), .A2(new_n2219_), .ZN(new_n2224_));
  OAI21_X1   g02000(.A1(new_n2223_), .A2(new_n2224_), .B(new_n2222_), .ZN(new_n2225_));
  NAND2_X1   g02001(.A1(new_n2225_), .A2(new_n2221_), .ZN(new_n2226_));
  NAND2_X1   g02002(.A1(new_n2173_), .A2(new_n2226_), .ZN(new_n2227_));
  NAND2_X1   g02003(.A1(new_n2082_), .A2(new_n2080_), .ZN(new_n2228_));
  NAND2_X1   g02004(.A1(new_n2218_), .A2(new_n2219_), .ZN(new_n2229_));
  NAND2_X1   g02005(.A1(new_n2203_), .A2(new_n2215_), .ZN(new_n2230_));
  AOI21_X1   g02006(.A1(new_n2229_), .A2(new_n2230_), .B(new_n2222_), .ZN(new_n2231_));
  NAND2_X1   g02007(.A1(new_n2203_), .A2(new_n2219_), .ZN(new_n2232_));
  NAND2_X1   g02008(.A1(new_n2218_), .A2(new_n2215_), .ZN(new_n2233_));
  AOI21_X1   g02009(.A1(new_n2233_), .A2(new_n2232_), .B(new_n2175_), .ZN(new_n2234_));
  NOR2_X1    g02010(.A1(new_n2231_), .A2(new_n2234_), .ZN(new_n2235_));
  NAND3_X1   g02011(.A1(new_n2235_), .A2(new_n2228_), .A3(new_n2081_), .ZN(new_n2236_));
  NAND2_X1   g02012(.A1(new_n2236_), .A2(new_n2227_), .ZN(new_n2237_));
  OAI21_X1   g02013(.A1(new_n2172_), .A2(new_n2171_), .B(new_n2237_), .ZN(new_n2238_));
  OAI21_X1   g02014(.A1(new_n2084_), .A2(new_n2153_), .B(new_n2157_), .ZN(new_n2239_));
  NAND3_X1   g02015(.A1(new_n2226_), .A2(new_n2228_), .A3(new_n2081_), .ZN(new_n2240_));
  NAND2_X1   g02016(.A1(new_n2235_), .A2(new_n2173_), .ZN(new_n2241_));
  NAND2_X1   g02017(.A1(new_n2241_), .A2(new_n2240_), .ZN(new_n2242_));
  NAND3_X1   g02018(.A1(new_n2239_), .A2(new_n2242_), .A3(new_n2159_), .ZN(new_n2243_));
  AND2_X2    g02019(.A1(new_n2238_), .A2(new_n2243_), .Z(new_n2244_));
  AOI21_X1   g02020(.A1(new_n2085_), .A2(new_n2150_), .B(new_n2136_), .ZN(new_n2245_));
  AOI21_X1   g02021(.A1(new_n2093_), .A2(new_n2106_), .B(new_n2108_), .ZN(new_n2246_));
  INV_X1     g02022(.I(new_n2246_), .ZN(new_n2247_));
  INV_X1     g02023(.I(new_n2059_), .ZN(new_n2248_));
  INV_X1     g02024(.I(new_n2065_), .ZN(new_n2249_));
  NOR2_X1    g02025(.A1(new_n2248_), .A2(new_n2249_), .ZN(new_n2250_));
  NOR2_X1    g02026(.A1(new_n2059_), .A2(new_n2065_), .ZN(new_n2251_));
  INV_X1     g02027(.I(new_n2066_), .ZN(new_n2252_));
  XOR2_X1    g02028(.A1(new_n2055_), .A2(new_n2252_), .Z(new_n2253_));
  NOR2_X1    g02029(.A1(new_n2253_), .A2(new_n2251_), .ZN(new_n2254_));
  NOR2_X1    g02030(.A1(new_n2254_), .A2(new_n2250_), .ZN(new_n2255_));
  NAND2_X1   g02031(.A1(\a[1] ), .A2(\a[27] ), .ZN(new_n2256_));
  INV_X1     g02032(.I(new_n2256_), .ZN(new_n2257_));
  INV_X1     g02033(.I(new_n2101_), .ZN(new_n2258_));
  NOR2_X1    g02034(.A1(\a[5] ), .A2(\a[22] ), .ZN(new_n2259_));
  OAI21_X1   g02035(.A1(new_n1150_), .A2(new_n1018_), .B(new_n2259_), .ZN(new_n2260_));
  NAND2_X1   g02036(.A1(new_n2094_), .A2(new_n2260_), .ZN(new_n2261_));
  XOR2_X1    g02037(.A1(new_n2261_), .A2(new_n873_), .Z(new_n2262_));
  XOR2_X1    g02038(.A1(new_n2262_), .A2(new_n2258_), .Z(new_n2263_));
  NOR2_X1    g02039(.A1(new_n2263_), .A2(new_n2257_), .ZN(new_n2264_));
  XOR2_X1    g02040(.A1(new_n2262_), .A2(new_n2101_), .Z(new_n2265_));
  NOR2_X1    g02041(.A1(new_n2265_), .A2(new_n2256_), .ZN(new_n2266_));
  NOR2_X1    g02042(.A1(new_n2264_), .A2(new_n2266_), .ZN(new_n2267_));
  NOR2_X1    g02043(.A1(new_n2267_), .A2(new_n2255_), .ZN(new_n2268_));
  NAND2_X1   g02044(.A1(new_n2267_), .A2(new_n2255_), .ZN(new_n2269_));
  INV_X1     g02045(.I(new_n2269_), .ZN(new_n2270_));
  OAI21_X1   g02046(.A1(new_n2270_), .A2(new_n2268_), .B(new_n2247_), .ZN(new_n2271_));
  OAI21_X1   g02047(.A1(new_n2264_), .A2(new_n2266_), .B(new_n2255_), .ZN(new_n2272_));
  INV_X1     g02048(.I(new_n2272_), .ZN(new_n2273_));
  NOR3_X1    g02049(.A1(new_n2264_), .A2(new_n2266_), .A3(new_n2255_), .ZN(new_n2274_));
  OAI21_X1   g02050(.A1(new_n2273_), .A2(new_n2274_), .B(new_n2246_), .ZN(new_n2275_));
  NAND2_X1   g02051(.A1(\a[24] ), .A2(\a[25] ), .ZN(new_n2276_));
  INV_X1     g02052(.I(new_n2276_), .ZN(new_n2277_));
  NAND2_X1   g02053(.A1(new_n267_), .A2(new_n2277_), .ZN(new_n2278_));
  NAND2_X1   g02054(.A1(\a[8] ), .A2(\a[20] ), .ZN(new_n2279_));
  XNOR2_X1   g02055(.A1(new_n2278_), .A2(new_n2279_), .ZN(new_n2280_));
  NAND2_X1   g02056(.A1(\a[0] ), .A2(\a[27] ), .ZN(new_n2281_));
  AOI21_X1   g02057(.A1(new_n2102_), .A2(new_n2099_), .B(new_n2281_), .ZN(new_n2282_));
  NOR2_X1    g02058(.A1(new_n2282_), .A2(new_n2103_), .ZN(new_n2283_));
  OAI22_X1   g02059(.A1(new_n478_), .A2(new_n1706_), .B1(new_n1000_), .B2(new_n1773_), .ZN(new_n2284_));
  NAND2_X1   g02060(.A1(\a[22] ), .A2(\a[23] ), .ZN(new_n2285_));
  INV_X1     g02061(.I(new_n2285_), .ZN(new_n2286_));
  NOR2_X1    g02062(.A1(new_n268_), .A2(new_n1313_), .ZN(new_n2287_));
  INV_X1     g02063(.I(new_n2287_), .ZN(new_n2288_));
  NOR4_X1    g02064(.A1(new_n2284_), .A2(new_n2288_), .A3(new_n608_), .A4(new_n2286_), .ZN(new_n2289_));
  XOR2_X1    g02065(.A1(new_n2283_), .A2(new_n2289_), .Z(new_n2290_));
  NOR2_X1    g02066(.A1(new_n2290_), .A2(new_n2280_), .ZN(new_n2291_));
  INV_X1     g02067(.I(new_n2280_), .ZN(new_n2292_));
  INV_X1     g02068(.I(new_n2289_), .ZN(new_n2293_));
  NOR2_X1    g02069(.A1(new_n2283_), .A2(new_n2293_), .ZN(new_n2294_));
  INV_X1     g02070(.I(new_n2294_), .ZN(new_n2295_));
  NAND2_X1   g02071(.A1(new_n2283_), .A2(new_n2293_), .ZN(new_n2296_));
  AOI21_X1   g02072(.A1(new_n2295_), .A2(new_n2296_), .B(new_n2292_), .ZN(new_n2297_));
  NOR2_X1    g02073(.A1(new_n2291_), .A2(new_n2297_), .ZN(new_n2298_));
  INV_X1     g02074(.I(new_n2298_), .ZN(new_n2299_));
  NAND3_X1   g02075(.A1(new_n2271_), .A2(new_n2275_), .A3(new_n2299_), .ZN(new_n2300_));
  INV_X1     g02076(.I(new_n2268_), .ZN(new_n2301_));
  AOI21_X1   g02077(.A1(new_n2301_), .A2(new_n2269_), .B(new_n2246_), .ZN(new_n2302_));
  INV_X1     g02078(.I(new_n2275_), .ZN(new_n2303_));
  OAI21_X1   g02079(.A1(new_n2302_), .A2(new_n2303_), .B(new_n2298_), .ZN(new_n2304_));
  AOI21_X1   g02080(.A1(new_n2304_), .A2(new_n2300_), .B(new_n2245_), .ZN(new_n2305_));
  INV_X1     g02081(.I(new_n2245_), .ZN(new_n2306_));
  OAI21_X1   g02082(.A1(new_n2302_), .A2(new_n2303_), .B(new_n2299_), .ZN(new_n2307_));
  NAND3_X1   g02083(.A1(new_n2271_), .A2(new_n2275_), .A3(new_n2298_), .ZN(new_n2308_));
  AOI21_X1   g02084(.A1(new_n2307_), .A2(new_n2308_), .B(new_n2306_), .ZN(new_n2309_));
  NOR2_X1    g02085(.A1(new_n2309_), .A2(new_n2305_), .ZN(new_n2310_));
  XOR2_X1    g02086(.A1(new_n2244_), .A2(new_n2310_), .Z(new_n2311_));
  NAND2_X1   g02087(.A1(new_n2170_), .A2(new_n2311_), .ZN(new_n2312_));
  AOI21_X1   g02088(.A1(new_n2238_), .A2(new_n2243_), .B(new_n2310_), .ZN(new_n2313_));
  NAND3_X1   g02089(.A1(new_n2238_), .A2(new_n2243_), .A3(new_n2310_), .ZN(new_n2314_));
  INV_X1     g02090(.I(new_n2314_), .ZN(new_n2315_));
  NOR2_X1    g02091(.A1(new_n2315_), .A2(new_n2313_), .ZN(new_n2316_));
  OAI21_X1   g02092(.A1(new_n2170_), .A2(new_n2316_), .B(new_n2312_), .ZN(\asquared[29] ));
  NAND2_X1   g02093(.A1(new_n2314_), .A2(new_n2161_), .ZN(new_n2318_));
  OAI21_X1   g02094(.A1(new_n2314_), .A2(new_n2161_), .B(new_n2030_), .ZN(new_n2319_));
  NAND2_X1   g02095(.A1(new_n2319_), .A2(new_n2318_), .ZN(new_n2320_));
  NOR2_X1    g02096(.A1(new_n2029_), .A2(new_n2320_), .ZN(new_n2321_));
  OAI21_X1   g02097(.A1(new_n2172_), .A2(new_n2171_), .B(new_n2240_), .ZN(new_n2322_));
  AND2_X2    g02098(.A1(new_n2322_), .A2(new_n2241_), .Z(new_n2323_));
  AOI21_X1   g02099(.A1(new_n2175_), .A2(new_n2232_), .B(new_n2224_), .ZN(new_n2324_));
  INV_X1     g02100(.I(new_n2199_), .ZN(new_n2325_));
  OAI21_X1   g02101(.A1(new_n2187_), .A2(new_n2201_), .B(new_n2325_), .ZN(new_n2326_));
  INV_X1     g02102(.I(new_n2326_), .ZN(new_n2327_));
  INV_X1     g02103(.I(new_n873_), .ZN(new_n2328_));
  NAND2_X1   g02104(.A1(\a[27] ), .A2(\a[29] ), .ZN(new_n2329_));
  XOR2_X1    g02105(.A1(new_n197_), .A2(new_n2329_), .Z(new_n2330_));
  INV_X1     g02106(.I(new_n1342_), .ZN(new_n2331_));
  AOI21_X1   g02107(.A1(new_n597_), .A2(new_n2191_), .B(new_n2331_), .ZN(new_n2332_));
  INV_X1     g02108(.I(new_n2332_), .ZN(new_n2333_));
  NAND2_X1   g02109(.A1(new_n2333_), .A2(new_n2330_), .ZN(new_n2334_));
  NOR2_X1    g02110(.A1(new_n2333_), .A2(new_n2330_), .ZN(new_n2335_));
  INV_X1     g02111(.I(new_n2335_), .ZN(new_n2336_));
  AOI21_X1   g02112(.A1(new_n2336_), .A2(new_n2334_), .B(new_n2185_), .ZN(new_n2337_));
  INV_X1     g02113(.I(new_n2185_), .ZN(new_n2338_));
  XOR2_X1    g02114(.A1(new_n2330_), .A2(new_n2332_), .Z(new_n2339_));
  NOR2_X1    g02115(.A1(new_n2339_), .A2(new_n2338_), .ZN(new_n2340_));
  NOR2_X1    g02116(.A1(new_n2340_), .A2(new_n2337_), .ZN(new_n2341_));
  AOI21_X1   g02117(.A1(new_n2283_), .A2(new_n2293_), .B(new_n2280_), .ZN(new_n2342_));
  NOR2_X1    g02118(.A1(new_n2342_), .A2(new_n2294_), .ZN(new_n2343_));
  XNOR2_X1   g02119(.A1(new_n2341_), .A2(new_n2343_), .ZN(new_n2344_));
  NOR2_X1    g02120(.A1(new_n2344_), .A2(new_n2327_), .ZN(new_n2345_));
  OAI22_X1   g02121(.A1(new_n2337_), .A2(new_n2340_), .B1(new_n2342_), .B2(new_n2294_), .ZN(new_n2346_));
  NAND2_X1   g02122(.A1(new_n2341_), .A2(new_n2343_), .ZN(new_n2347_));
  AOI21_X1   g02123(.A1(new_n2346_), .A2(new_n2347_), .B(new_n2326_), .ZN(new_n2348_));
  NOR2_X1    g02124(.A1(new_n2345_), .A2(new_n2348_), .ZN(new_n2349_));
  INV_X1     g02125(.I(new_n2274_), .ZN(new_n2350_));
  OAI21_X1   g02126(.A1(new_n2246_), .A2(new_n2273_), .B(new_n2350_), .ZN(new_n2351_));
  NAND2_X1   g02127(.A1(new_n2351_), .A2(new_n2349_), .ZN(new_n2352_));
  INV_X1     g02128(.I(new_n2349_), .ZN(new_n2353_));
  AOI21_X1   g02129(.A1(new_n2247_), .A2(new_n2272_), .B(new_n2274_), .ZN(new_n2354_));
  NAND2_X1   g02130(.A1(new_n2353_), .A2(new_n2354_), .ZN(new_n2355_));
  AOI21_X1   g02131(.A1(new_n2352_), .A2(new_n2355_), .B(new_n2324_), .ZN(new_n2356_));
  INV_X1     g02132(.I(new_n2356_), .ZN(new_n2357_));
  XNOR2_X1   g02133(.A1(new_n2354_), .A2(new_n2349_), .ZN(new_n2358_));
  NAND2_X1   g02134(.A1(new_n2358_), .A2(new_n2324_), .ZN(new_n2359_));
  NAND2_X1   g02135(.A1(new_n2359_), .A2(new_n2357_), .ZN(new_n2360_));
  NAND2_X1   g02136(.A1(new_n2307_), .A2(new_n2306_), .ZN(new_n2361_));
  NAND2_X1   g02137(.A1(new_n2213_), .A2(new_n2211_), .ZN(new_n2362_));
  NOR2_X1    g02138(.A1(new_n2261_), .A2(new_n2258_), .ZN(new_n2363_));
  NAND2_X1   g02139(.A1(new_n2257_), .A2(new_n873_), .ZN(new_n2364_));
  NAND2_X1   g02140(.A1(new_n2328_), .A2(new_n2256_), .ZN(new_n2365_));
  AOI22_X1   g02141(.A1(new_n2261_), .A2(new_n2258_), .B1(new_n2364_), .B2(new_n2365_), .ZN(new_n2366_));
  NOR2_X1    g02142(.A1(new_n2366_), .A2(new_n2363_), .ZN(new_n2367_));
  INV_X1     g02143(.I(\a[23] ), .ZN(new_n2368_));
  NOR3_X1    g02144(.A1(new_n1018_), .A2(new_n599_), .A3(new_n800_), .ZN(new_n2369_));
  XOR2_X1    g02145(.A1(new_n2369_), .A2(new_n242_), .Z(new_n2370_));
  XOR2_X1    g02146(.A1(new_n2370_), .A2(new_n2368_), .Z(new_n2371_));
  NAND2_X1   g02147(.A1(new_n2371_), .A2(new_n2367_), .ZN(new_n2372_));
  INV_X1     g02148(.I(new_n2367_), .ZN(new_n2373_));
  INV_X1     g02149(.I(new_n2371_), .ZN(new_n2374_));
  NAND2_X1   g02150(.A1(new_n2374_), .A2(new_n2373_), .ZN(new_n2375_));
  AOI22_X1   g02151(.A1(new_n2375_), .A2(new_n2372_), .B1(new_n2212_), .B2(new_n2362_), .ZN(new_n2376_));
  NAND2_X1   g02152(.A1(new_n2362_), .A2(new_n2212_), .ZN(new_n2377_));
  NAND2_X1   g02153(.A1(new_n2373_), .A2(new_n2371_), .ZN(new_n2378_));
  NAND2_X1   g02154(.A1(new_n2374_), .A2(new_n2367_), .ZN(new_n2379_));
  AOI21_X1   g02155(.A1(new_n2379_), .A2(new_n2378_), .B(new_n2377_), .ZN(new_n2380_));
  NOR2_X1    g02156(.A1(new_n2376_), .A2(new_n2380_), .ZN(new_n2381_));
  INV_X1     g02157(.I(new_n2381_), .ZN(new_n2382_));
  NOR2_X1    g02158(.A1(new_n1674_), .A2(new_n1691_), .ZN(new_n2383_));
  INV_X1     g02159(.I(new_n2383_), .ZN(new_n2384_));
  NOR2_X1    g02160(.A1(new_n282_), .A2(new_n1999_), .ZN(new_n2385_));
  NOR2_X1    g02161(.A1(new_n2384_), .A2(new_n1000_), .ZN(new_n2386_));
  NAND4_X1   g02162(.A1(new_n2386_), .A2(\a[7] ), .A3(new_n2385_), .A4(\a[22] ), .ZN(new_n2387_));
  AOI21_X1   g02163(.A1(new_n2387_), .A2(new_n2276_), .B(new_n211_), .ZN(new_n2388_));
  NOR2_X1    g02164(.A1(new_n2384_), .A2(new_n1000_), .ZN(new_n2389_));
  INV_X1     g02165(.I(new_n2389_), .ZN(new_n2390_));
  NOR2_X1    g02166(.A1(new_n1536_), .A2(new_n1715_), .ZN(new_n2391_));
  INV_X1     g02167(.I(new_n2391_), .ZN(new_n2392_));
  NOR2_X1    g02168(.A1(new_n525_), .A2(new_n1236_), .ZN(new_n2393_));
  INV_X1     g02169(.I(new_n2393_), .ZN(new_n2394_));
  NAND2_X1   g02170(.A1(new_n2392_), .A2(new_n2394_), .ZN(new_n2395_));
  NAND4_X1   g02171(.A1(new_n796_), .A2(new_n1342_), .A3(\a[9] ), .A4(\a[20] ), .ZN(new_n2396_));
  NOR2_X1    g02172(.A1(new_n2395_), .A2(new_n2396_), .ZN(new_n2397_));
  INV_X1     g02173(.I(new_n2397_), .ZN(new_n2398_));
  NAND2_X1   g02174(.A1(\a[3] ), .A2(\a[8] ), .ZN(new_n2399_));
  OAI21_X1   g02175(.A1(new_n1313_), .A2(new_n1916_), .B(new_n2399_), .ZN(new_n2400_));
  NOR4_X1    g02176(.A1(new_n200_), .A2(new_n359_), .A3(new_n1313_), .A4(new_n1916_), .ZN(new_n2401_));
  NAND2_X1   g02177(.A1(new_n2400_), .A2(new_n2401_), .ZN(new_n2402_));
  NAND2_X1   g02178(.A1(\a[12] ), .A2(\a[17] ), .ZN(new_n2403_));
  XNOR2_X1   g02179(.A1(new_n2402_), .A2(new_n2403_), .ZN(new_n2404_));
  NOR2_X1    g02180(.A1(new_n2404_), .A2(new_n2398_), .ZN(new_n2405_));
  INV_X1     g02181(.I(new_n2405_), .ZN(new_n2406_));
  NAND2_X1   g02182(.A1(new_n2404_), .A2(new_n2398_), .ZN(new_n2407_));
  AOI21_X1   g02183(.A1(new_n2406_), .A2(new_n2407_), .B(new_n2390_), .ZN(new_n2408_));
  XOR2_X1    g02184(.A1(new_n2404_), .A2(new_n2397_), .Z(new_n2409_));
  NOR2_X1    g02185(.A1(new_n2409_), .A2(new_n2389_), .ZN(new_n2410_));
  NOR2_X1    g02186(.A1(new_n2410_), .A2(new_n2408_), .ZN(new_n2411_));
  NAND2_X1   g02187(.A1(new_n267_), .A2(new_n2277_), .ZN(new_n2412_));
  NOR2_X1    g02188(.A1(new_n267_), .A2(new_n2277_), .ZN(new_n2413_));
  NOR2_X1    g02189(.A1(\a[8] ), .A2(\a[20] ), .ZN(new_n2414_));
  AOI21_X1   g02190(.A1(new_n2412_), .A2(new_n2414_), .B(new_n2413_), .ZN(new_n2415_));
  INV_X1     g02191(.I(new_n2415_), .ZN(new_n2416_));
  OAI21_X1   g02192(.A1(new_n481_), .A2(new_n2285_), .B(new_n2284_), .ZN(new_n2417_));
  NAND2_X1   g02193(.A1(\a[1] ), .A2(\a[28] ), .ZN(new_n2418_));
  XOR2_X1    g02194(.A1(new_n2418_), .A2(new_n875_), .Z(new_n2419_));
  XNOR2_X1   g02195(.A1(new_n2417_), .A2(new_n2419_), .ZN(new_n2420_));
  NOR2_X1    g02196(.A1(new_n2420_), .A2(new_n2416_), .ZN(new_n2421_));
  NAND2_X1   g02197(.A1(new_n2417_), .A2(new_n2419_), .ZN(new_n2422_));
  NOR2_X1    g02198(.A1(new_n2417_), .A2(new_n2419_), .ZN(new_n2423_));
  INV_X1     g02199(.I(new_n2423_), .ZN(new_n2424_));
  AOI21_X1   g02200(.A1(new_n2424_), .A2(new_n2422_), .B(new_n2415_), .ZN(new_n2425_));
  NOR2_X1    g02201(.A1(new_n2421_), .A2(new_n2425_), .ZN(new_n2426_));
  INV_X1     g02202(.I(new_n2426_), .ZN(new_n2427_));
  NAND2_X1   g02203(.A1(new_n2411_), .A2(new_n2427_), .ZN(new_n2428_));
  OAI21_X1   g02204(.A1(new_n2410_), .A2(new_n2408_), .B(new_n2426_), .ZN(new_n2429_));
  NAND2_X1   g02205(.A1(new_n2428_), .A2(new_n2429_), .ZN(new_n2430_));
  XOR2_X1    g02206(.A1(new_n2411_), .A2(new_n2426_), .Z(new_n2431_));
  NOR2_X1    g02207(.A1(new_n2431_), .A2(new_n2382_), .ZN(new_n2432_));
  AOI21_X1   g02208(.A1(new_n2382_), .A2(new_n2430_), .B(new_n2432_), .ZN(new_n2433_));
  AOI21_X1   g02209(.A1(new_n2361_), .A2(new_n2308_), .B(new_n2433_), .ZN(new_n2434_));
  INV_X1     g02210(.I(new_n2308_), .ZN(new_n2435_));
  AOI21_X1   g02211(.A1(new_n2271_), .A2(new_n2275_), .B(new_n2298_), .ZN(new_n2436_));
  NOR2_X1    g02212(.A1(new_n2436_), .A2(new_n2245_), .ZN(new_n2437_));
  INV_X1     g02213(.I(new_n2433_), .ZN(new_n2438_));
  NOR3_X1    g02214(.A1(new_n2437_), .A2(new_n2438_), .A3(new_n2435_), .ZN(new_n2439_));
  OAI21_X1   g02215(.A1(new_n2439_), .A2(new_n2434_), .B(new_n2360_), .ZN(new_n2440_));
  AOI21_X1   g02216(.A1(new_n2358_), .A2(new_n2324_), .B(new_n2356_), .ZN(new_n2441_));
  NOR3_X1    g02217(.A1(new_n2437_), .A2(new_n2435_), .A3(new_n2433_), .ZN(new_n2442_));
  AOI21_X1   g02218(.A1(new_n2361_), .A2(new_n2308_), .B(new_n2438_), .ZN(new_n2443_));
  OAI21_X1   g02219(.A1(new_n2443_), .A2(new_n2442_), .B(new_n2441_), .ZN(new_n2444_));
  AND2_X2    g02220(.A1(new_n2440_), .A2(new_n2444_), .Z(new_n2445_));
  NOR2_X1    g02221(.A1(new_n2445_), .A2(new_n2323_), .ZN(new_n2446_));
  XOR2_X1    g02222(.A1(new_n2321_), .A2(new_n2446_), .Z(new_n2447_));
  XOR2_X1    g02223(.A1(new_n2447_), .A2(new_n2313_), .Z(\asquared[30] ));
  NAND4_X1   g02224(.A1(new_n2440_), .A2(new_n2444_), .A3(new_n2241_), .A4(new_n2322_), .ZN(new_n2449_));
  NAND2_X1   g02225(.A1(new_n2449_), .A2(new_n2313_), .ZN(new_n2450_));
  NOR3_X1    g02226(.A1(new_n2029_), .A2(new_n2320_), .A3(new_n2450_), .ZN(new_n2451_));
  NOR2_X1    g02227(.A1(new_n2451_), .A2(new_n2446_), .ZN(new_n2452_));
  NOR2_X1    g02228(.A1(new_n2442_), .A2(new_n2441_), .ZN(new_n2453_));
  OR2_X2     g02229(.A1(new_n2453_), .A2(new_n2443_), .Z(new_n2454_));
  NAND2_X1   g02230(.A1(new_n2428_), .A2(new_n2381_), .ZN(new_n2455_));
  NAND2_X1   g02231(.A1(new_n2455_), .A2(new_n2429_), .ZN(new_n2456_));
  INV_X1     g02232(.I(new_n2456_), .ZN(new_n2457_));
  OAI21_X1   g02233(.A1(new_n2185_), .A2(new_n2335_), .B(new_n2334_), .ZN(new_n2458_));
  INV_X1     g02234(.I(new_n2458_), .ZN(new_n2459_));
  AOI21_X1   g02235(.A1(new_n2415_), .A2(new_n2422_), .B(new_n2423_), .ZN(new_n2460_));
  INV_X1     g02236(.I(\a[30] ), .ZN(new_n2461_));
  NAND2_X1   g02237(.A1(\a[1] ), .A2(\a[29] ), .ZN(new_n2462_));
  NAND2_X1   g02238(.A1(new_n1017_), .A2(new_n2462_), .ZN(new_n2463_));
  NAND3_X1   g02239(.A1(new_n1718_), .A2(\a[1] ), .A3(\a[29] ), .ZN(new_n2464_));
  NAND2_X1   g02240(.A1(new_n2464_), .A2(new_n2463_), .ZN(new_n2465_));
  NOR2_X1    g02241(.A1(new_n773_), .A2(new_n2178_), .ZN(new_n2466_));
  NAND2_X1   g02242(.A1(new_n2465_), .A2(new_n2466_), .ZN(new_n2467_));
  XOR2_X1    g02243(.A1(new_n2467_), .A2(new_n199_), .Z(new_n2468_));
  NAND2_X1   g02244(.A1(new_n2468_), .A2(new_n2461_), .ZN(new_n2469_));
  XOR2_X1    g02245(.A1(new_n2467_), .A2(\a[0] ), .Z(new_n2470_));
  NAND2_X1   g02246(.A1(new_n2470_), .A2(\a[30] ), .ZN(new_n2471_));
  NAND2_X1   g02247(.A1(new_n2469_), .A2(new_n2471_), .ZN(new_n2472_));
  XOR2_X1    g02248(.A1(new_n2472_), .A2(new_n2460_), .Z(new_n2473_));
  NOR2_X1    g02249(.A1(new_n2470_), .A2(\a[30] ), .ZN(new_n2474_));
  NOR2_X1    g02250(.A1(new_n2468_), .A2(new_n2461_), .ZN(new_n2475_));
  NOR2_X1    g02251(.A1(new_n2474_), .A2(new_n2475_), .ZN(new_n2476_));
  NOR2_X1    g02252(.A1(new_n2476_), .A2(new_n2460_), .ZN(new_n2477_));
  INV_X1     g02253(.I(new_n2460_), .ZN(new_n2478_));
  NOR2_X1    g02254(.A1(new_n2472_), .A2(new_n2478_), .ZN(new_n2479_));
  OAI21_X1   g02255(.A1(new_n2477_), .A2(new_n2479_), .B(new_n2459_), .ZN(new_n2480_));
  OAI21_X1   g02256(.A1(new_n2473_), .A2(new_n2459_), .B(new_n2480_), .ZN(new_n2481_));
  INV_X1     g02257(.I(new_n2481_), .ZN(new_n2482_));
  NOR2_X1    g02258(.A1(new_n2388_), .A2(new_n2386_), .ZN(new_n2483_));
  AOI21_X1   g02259(.A1(\a[13] ), .A2(\a[16] ), .B(new_n1447_), .ZN(new_n2484_));
  NOR3_X1    g02260(.A1(new_n2484_), .A2(new_n242_), .A3(new_n2368_), .ZN(new_n2485_));
  NOR2_X1    g02261(.A1(new_n2485_), .A2(new_n2369_), .ZN(new_n2486_));
  NAND4_X1   g02262(.A1(\a[2] ), .A2(\a[9] ), .A3(\a[21] ), .A4(\a[28] ), .ZN(new_n2487_));
  XOR2_X1    g02263(.A1(new_n2487_), .A2(\a[13] ), .Z(new_n2488_));
  XOR2_X1    g02264(.A1(new_n2488_), .A2(\a[17] ), .Z(new_n2489_));
  NOR2_X1    g02265(.A1(new_n2489_), .A2(new_n2486_), .ZN(new_n2490_));
  XOR2_X1    g02266(.A1(new_n2488_), .A2(new_n885_), .Z(new_n2491_));
  NOR3_X1    g02267(.A1(new_n2491_), .A2(new_n2369_), .A3(new_n2485_), .ZN(new_n2492_));
  OAI21_X1   g02268(.A1(new_n2492_), .A2(new_n2490_), .B(new_n2483_), .ZN(new_n2493_));
  XOR2_X1    g02269(.A1(new_n2491_), .A2(new_n2486_), .Z(new_n2494_));
  OAI21_X1   g02270(.A1(new_n2494_), .A2(new_n2483_), .B(new_n2493_), .ZN(new_n2495_));
  INV_X1     g02271(.I(new_n2495_), .ZN(new_n2496_));
  AOI21_X1   g02272(.A1(new_n2404_), .A2(new_n2398_), .B(new_n2390_), .ZN(new_n2497_));
  NOR2_X1    g02273(.A1(new_n2497_), .A2(new_n2405_), .ZN(new_n2498_));
  INV_X1     g02274(.I(\a[29] ), .ZN(new_n2499_));
  NOR2_X1    g02275(.A1(new_n2098_), .A2(new_n2499_), .ZN(new_n2500_));
  NOR2_X1    g02276(.A1(new_n873_), .A2(new_n2256_), .ZN(new_n2501_));
  AOI21_X1   g02277(.A1(new_n2501_), .A2(new_n218_), .B(new_n2500_), .ZN(new_n2502_));
  INV_X1     g02278(.I(new_n2502_), .ZN(new_n2503_));
  OAI22_X1   g02279(.A1(new_n2391_), .A2(new_n2393_), .B1(new_n796_), .B2(new_n1342_), .ZN(new_n2504_));
  NAND2_X1   g02280(.A1(new_n566_), .A2(new_n885_), .ZN(new_n2505_));
  OAI21_X1   g02281(.A1(new_n2401_), .A2(new_n2505_), .B(new_n2400_), .ZN(new_n2506_));
  XOR2_X1    g02282(.A1(new_n2506_), .A2(new_n2504_), .Z(new_n2507_));
  NAND2_X1   g02283(.A1(new_n2507_), .A2(new_n2503_), .ZN(new_n2508_));
  NOR2_X1    g02284(.A1(new_n2506_), .A2(new_n2504_), .ZN(new_n2509_));
  AND2_X2    g02285(.A1(new_n2506_), .A2(new_n2504_), .Z(new_n2510_));
  OAI21_X1   g02286(.A1(new_n2510_), .A2(new_n2509_), .B(new_n2502_), .ZN(new_n2511_));
  NAND2_X1   g02287(.A1(new_n2508_), .A2(new_n2511_), .ZN(new_n2512_));
  XNOR2_X1   g02288(.A1(new_n2498_), .A2(new_n2512_), .ZN(new_n2513_));
  NOR2_X1    g02289(.A1(new_n2496_), .A2(new_n2513_), .ZN(new_n2514_));
  NAND2_X1   g02290(.A1(new_n2498_), .A2(new_n2512_), .ZN(new_n2515_));
  OR2_X2     g02291(.A1(new_n2498_), .A2(new_n2512_), .Z(new_n2516_));
  AOI21_X1   g02292(.A1(new_n2516_), .A2(new_n2515_), .B(new_n2495_), .ZN(new_n2517_));
  NOR2_X1    g02293(.A1(new_n2514_), .A2(new_n2517_), .ZN(new_n2518_));
  INV_X1     g02294(.I(new_n2518_), .ZN(new_n2519_));
  NAND2_X1   g02295(.A1(new_n2482_), .A2(new_n2519_), .ZN(new_n2520_));
  NAND2_X1   g02296(.A1(new_n2481_), .A2(new_n2518_), .ZN(new_n2521_));
  AOI21_X1   g02297(.A1(new_n2520_), .A2(new_n2521_), .B(new_n2457_), .ZN(new_n2522_));
  NAND2_X1   g02298(.A1(new_n2519_), .A2(new_n2481_), .ZN(new_n2523_));
  NAND2_X1   g02299(.A1(new_n2482_), .A2(new_n2518_), .ZN(new_n2524_));
  AOI21_X1   g02300(.A1(new_n2524_), .A2(new_n2523_), .B(new_n2456_), .ZN(new_n2525_));
  NOR2_X1    g02301(.A1(new_n2351_), .A2(new_n2349_), .ZN(new_n2526_));
  OAI21_X1   g02302(.A1(new_n2324_), .A2(new_n2526_), .B(new_n2352_), .ZN(new_n2527_));
  NAND2_X1   g02303(.A1(new_n2326_), .A2(new_n2347_), .ZN(new_n2528_));
  NAND2_X1   g02304(.A1(new_n2528_), .A2(new_n2346_), .ZN(new_n2529_));
  NAND2_X1   g02305(.A1(new_n2379_), .A2(new_n2377_), .ZN(new_n2530_));
  NAND2_X1   g02306(.A1(new_n2530_), .A2(new_n2378_), .ZN(new_n2531_));
  NAND2_X1   g02307(.A1(\a[22] ), .A2(\a[27] ), .ZN(new_n2532_));
  NOR2_X1    g02308(.A1(new_n1916_), .A2(new_n2098_), .ZN(new_n2533_));
  INV_X1     g02309(.I(new_n2533_), .ZN(new_n2534_));
  OAI22_X1   g02310(.A1(new_n2534_), .A2(new_n212_), .B1(new_n2399_), .B2(new_n2532_), .ZN(new_n2535_));
  INV_X1     g02311(.I(new_n2535_), .ZN(new_n2536_));
  NAND2_X1   g02312(.A1(\a[4] ), .A2(\a[26] ), .ZN(new_n2537_));
  NAND2_X1   g02313(.A1(\a[8] ), .A2(\a[22] ), .ZN(new_n2538_));
  XOR2_X1    g02314(.A1(new_n2537_), .A2(new_n2538_), .Z(new_n2539_));
  AOI21_X1   g02315(.A1(\a[4] ), .A2(\a[26] ), .B(new_n2538_), .ZN(new_n2540_));
  NOR2_X1    g02316(.A1(new_n200_), .A2(new_n2098_), .ZN(new_n2541_));
  OAI22_X1   g02317(.A1(new_n2536_), .A2(new_n2540_), .B1(new_n2539_), .B2(new_n2541_), .ZN(new_n2542_));
  INV_X1     g02318(.I(new_n1956_), .ZN(new_n2543_));
  OAI22_X1   g02319(.A1(new_n481_), .A2(new_n1912_), .B1(new_n1000_), .B2(new_n2276_), .ZN(new_n2544_));
  NAND2_X1   g02320(.A1(\a[5] ), .A2(\a[25] ), .ZN(new_n2545_));
  NOR4_X1    g02321(.A1(new_n2544_), .A2(new_n479_), .A3(new_n2543_), .A4(new_n2545_), .ZN(new_n2546_));
  OAI22_X1   g02322(.A1(new_n523_), .A2(new_n1715_), .B1(new_n796_), .B2(new_n1536_), .ZN(new_n2547_));
  NOR2_X1    g02323(.A1(new_n461_), .A2(new_n1215_), .ZN(new_n2548_));
  NAND3_X1   g02324(.A1(new_n2548_), .A2(new_n651_), .A3(new_n1342_), .ZN(new_n2549_));
  NOR2_X1    g02325(.A1(new_n2549_), .A2(new_n2547_), .ZN(new_n2550_));
  NAND2_X1   g02326(.A1(new_n2546_), .A2(new_n2550_), .ZN(new_n2551_));
  NOR2_X1    g02327(.A1(new_n2546_), .A2(new_n2550_), .ZN(new_n2552_));
  INV_X1     g02328(.I(new_n2552_), .ZN(new_n2553_));
  AOI21_X1   g02329(.A1(new_n2553_), .A2(new_n2551_), .B(new_n2542_), .ZN(new_n2554_));
  XOR2_X1    g02330(.A1(new_n2546_), .A2(new_n2550_), .Z(new_n2555_));
  AND2_X2    g02331(.A1(new_n2555_), .A2(new_n2542_), .Z(new_n2556_));
  NOR2_X1    g02332(.A1(new_n2556_), .A2(new_n2554_), .ZN(new_n2557_));
  INV_X1     g02333(.I(new_n2557_), .ZN(new_n2558_));
  XOR2_X1    g02334(.A1(new_n2531_), .A2(new_n2558_), .Z(new_n2559_));
  NAND2_X1   g02335(.A1(new_n2559_), .A2(new_n2529_), .ZN(new_n2560_));
  INV_X1     g02336(.I(new_n2529_), .ZN(new_n2561_));
  NAND2_X1   g02337(.A1(new_n2531_), .A2(new_n2558_), .ZN(new_n2562_));
  INV_X1     g02338(.I(new_n2562_), .ZN(new_n2563_));
  NOR2_X1    g02339(.A1(new_n2531_), .A2(new_n2558_), .ZN(new_n2564_));
  OAI21_X1   g02340(.A1(new_n2563_), .A2(new_n2564_), .B(new_n2561_), .ZN(new_n2565_));
  NAND2_X1   g02341(.A1(new_n2560_), .A2(new_n2565_), .ZN(new_n2566_));
  INV_X1     g02342(.I(new_n2566_), .ZN(new_n2567_));
  NOR2_X1    g02343(.A1(new_n2527_), .A2(new_n2567_), .ZN(new_n2568_));
  INV_X1     g02344(.I(new_n2352_), .ZN(new_n2569_));
  NOR2_X1    g02345(.A1(new_n2526_), .A2(new_n2324_), .ZN(new_n2570_));
  NOR2_X1    g02346(.A1(new_n2570_), .A2(new_n2569_), .ZN(new_n2571_));
  NOR2_X1    g02347(.A1(new_n2571_), .A2(new_n2566_), .ZN(new_n2572_));
  OAI22_X1   g02348(.A1(new_n2572_), .A2(new_n2568_), .B1(new_n2522_), .B2(new_n2525_), .ZN(new_n2573_));
  NOR2_X1    g02349(.A1(new_n2522_), .A2(new_n2525_), .ZN(new_n2574_));
  NOR2_X1    g02350(.A1(new_n2571_), .A2(new_n2567_), .ZN(new_n2575_));
  NOR2_X1    g02351(.A1(new_n2527_), .A2(new_n2566_), .ZN(new_n2576_));
  OAI21_X1   g02352(.A1(new_n2575_), .A2(new_n2576_), .B(new_n2574_), .ZN(new_n2577_));
  NAND2_X1   g02353(.A1(new_n2573_), .A2(new_n2577_), .ZN(new_n2578_));
  XOR2_X1    g02354(.A1(new_n2454_), .A2(new_n2578_), .Z(new_n2579_));
  INV_X1     g02355(.I(new_n2454_), .ZN(new_n2580_));
  NAND2_X1   g02356(.A1(new_n2580_), .A2(new_n2578_), .ZN(new_n2581_));
  NAND3_X1   g02357(.A1(new_n2454_), .A2(new_n2573_), .A3(new_n2577_), .ZN(new_n2582_));
  NAND2_X1   g02358(.A1(new_n2581_), .A2(new_n2582_), .ZN(new_n2583_));
  NAND2_X1   g02359(.A1(new_n2452_), .A2(new_n2583_), .ZN(new_n2584_));
  OAI21_X1   g02360(.A1(new_n2452_), .A2(new_n2579_), .B(new_n2584_), .ZN(\asquared[31] ));
  OAI21_X1   g02361(.A1(new_n2451_), .A2(new_n2446_), .B(new_n2581_), .ZN(new_n2586_));
  NAND2_X1   g02362(.A1(new_n2586_), .A2(new_n2582_), .ZN(new_n2587_));
  OAI21_X1   g02363(.A1(new_n2561_), .A2(new_n2564_), .B(new_n2562_), .ZN(new_n2588_));
  NAND2_X1   g02364(.A1(new_n2476_), .A2(new_n2460_), .ZN(new_n2589_));
  AOI21_X1   g02365(.A1(new_n2458_), .A2(new_n2589_), .B(new_n2477_), .ZN(new_n2590_));
  NOR2_X1    g02366(.A1(new_n2537_), .A2(new_n2538_), .ZN(new_n2591_));
  NOR2_X1    g02367(.A1(new_n2535_), .A2(new_n2591_), .ZN(new_n2592_));
  INV_X1     g02368(.I(new_n2592_), .ZN(new_n2593_));
  OAI21_X1   g02369(.A1(new_n651_), .A2(new_n1342_), .B(new_n2547_), .ZN(new_n2594_));
  OAI22_X1   g02370(.A1(new_n201_), .A2(new_n2178_), .B1(new_n364_), .B2(new_n1313_), .ZN(new_n2595_));
  NAND3_X1   g02371(.A1(new_n2595_), .A2(\a[13] ), .A3(\a[17] ), .ZN(new_n2596_));
  NAND2_X1   g02372(.A1(new_n2596_), .A2(new_n2487_), .ZN(new_n2597_));
  XOR2_X1    g02373(.A1(new_n2597_), .A2(new_n2594_), .Z(new_n2598_));
  OR2_X2     g02374(.A1(new_n2598_), .A2(new_n2593_), .Z(new_n2599_));
  INV_X1     g02375(.I(new_n2597_), .ZN(new_n2600_));
  NOR2_X1    g02376(.A1(new_n2600_), .A2(new_n2594_), .ZN(new_n2601_));
  AND2_X2    g02377(.A1(new_n2600_), .A2(new_n2594_), .Z(new_n2602_));
  OAI21_X1   g02378(.A1(new_n2602_), .A2(new_n2601_), .B(new_n2593_), .ZN(new_n2603_));
  NAND2_X1   g02379(.A1(new_n2599_), .A2(new_n2603_), .ZN(new_n2604_));
  OAI21_X1   g02380(.A1(new_n2542_), .A2(new_n2552_), .B(new_n2551_), .ZN(new_n2605_));
  XOR2_X1    g02381(.A1(new_n2604_), .A2(new_n2605_), .Z(new_n2606_));
  NOR2_X1    g02382(.A1(new_n2606_), .A2(new_n2590_), .ZN(new_n2607_));
  NAND2_X1   g02383(.A1(new_n2472_), .A2(new_n2478_), .ZN(new_n2608_));
  OAI21_X1   g02384(.A1(new_n2459_), .A2(new_n2479_), .B(new_n2608_), .ZN(new_n2609_));
  NAND3_X1   g02385(.A1(new_n2599_), .A2(new_n2603_), .A3(new_n2605_), .ZN(new_n2610_));
  INV_X1     g02386(.I(new_n2605_), .ZN(new_n2611_));
  NAND2_X1   g02387(.A1(new_n2604_), .A2(new_n2611_), .ZN(new_n2612_));
  AOI21_X1   g02388(.A1(new_n2610_), .A2(new_n2612_), .B(new_n2609_), .ZN(new_n2613_));
  NOR2_X1    g02389(.A1(new_n2613_), .A2(new_n2607_), .ZN(new_n2614_));
  INV_X1     g02390(.I(new_n2614_), .ZN(new_n2615_));
  INV_X1     g02391(.I(new_n2483_), .ZN(new_n2616_));
  INV_X1     g02392(.I(new_n2490_), .ZN(new_n2617_));
  OAI21_X1   g02393(.A1(new_n2616_), .A2(new_n2492_), .B(new_n2617_), .ZN(new_n2618_));
  INV_X1     g02394(.I(new_n2618_), .ZN(new_n2619_));
  NOR2_X1    g02395(.A1(new_n2510_), .A2(new_n2502_), .ZN(new_n2620_));
  NOR2_X1    g02396(.A1(new_n2620_), .A2(new_n2509_), .ZN(new_n2621_));
  INV_X1     g02397(.I(new_n2621_), .ZN(new_n2622_));
  NAND2_X1   g02398(.A1(new_n479_), .A2(new_n2543_), .ZN(new_n2623_));
  NAND2_X1   g02399(.A1(new_n2623_), .A2(new_n2544_), .ZN(new_n2624_));
  NAND2_X1   g02400(.A1(\a[1] ), .A2(\a[30] ), .ZN(new_n2625_));
  INV_X1     g02401(.I(new_n2625_), .ZN(new_n2626_));
  XOR2_X1    g02402(.A1(new_n2624_), .A2(new_n2626_), .Z(new_n2627_));
  XOR2_X1    g02403(.A1(new_n2627_), .A2(new_n2464_), .Z(new_n2628_));
  NAND2_X1   g02404(.A1(new_n2628_), .A2(new_n800_), .ZN(new_n2629_));
  XNOR2_X1   g02405(.A1(new_n2627_), .A2(new_n2464_), .ZN(new_n2630_));
  NAND2_X1   g02406(.A1(new_n2630_), .A2(\a[16] ), .ZN(new_n2631_));
  NAND2_X1   g02407(.A1(new_n2631_), .A2(new_n2629_), .ZN(new_n2632_));
  NAND2_X1   g02408(.A1(new_n2632_), .A2(new_n2622_), .ZN(new_n2633_));
  XOR2_X1    g02409(.A1(new_n2628_), .A2(new_n800_), .Z(new_n2634_));
  NAND2_X1   g02410(.A1(new_n2634_), .A2(new_n2621_), .ZN(new_n2635_));
  AOI21_X1   g02411(.A1(new_n2635_), .A2(new_n2633_), .B(new_n2619_), .ZN(new_n2636_));
  NAND2_X1   g02412(.A1(new_n2632_), .A2(new_n2621_), .ZN(new_n2637_));
  NAND2_X1   g02413(.A1(new_n2634_), .A2(new_n2622_), .ZN(new_n2638_));
  AOI21_X1   g02414(.A1(new_n2638_), .A2(new_n2637_), .B(new_n2618_), .ZN(new_n2639_));
  NOR2_X1    g02415(.A1(new_n2636_), .A2(new_n2639_), .ZN(new_n2640_));
  NOR2_X1    g02416(.A1(new_n2615_), .A2(new_n2640_), .ZN(new_n2641_));
  OR2_X2     g02417(.A1(new_n2636_), .A2(new_n2639_), .Z(new_n2642_));
  NOR2_X1    g02418(.A1(new_n2642_), .A2(new_n2614_), .ZN(new_n2643_));
  OAI21_X1   g02419(.A1(new_n2643_), .A2(new_n2641_), .B(new_n2588_), .ZN(new_n2644_));
  INV_X1     g02420(.I(new_n2588_), .ZN(new_n2645_));
  NOR2_X1    g02421(.A1(new_n2640_), .A2(new_n2614_), .ZN(new_n2646_));
  NOR2_X1    g02422(.A1(new_n2642_), .A2(new_n2615_), .ZN(new_n2647_));
  OAI21_X1   g02423(.A1(new_n2647_), .A2(new_n2646_), .B(new_n2645_), .ZN(new_n2648_));
  NAND2_X1   g02424(.A1(new_n2523_), .A2(new_n2456_), .ZN(new_n2649_));
  NAND2_X1   g02425(.A1(new_n2495_), .A2(new_n2515_), .ZN(new_n2650_));
  NAND2_X1   g02426(.A1(new_n2650_), .A2(new_n2516_), .ZN(new_n2651_));
  INV_X1     g02427(.I(new_n2651_), .ZN(new_n2652_));
  NAND2_X1   g02428(.A1(\a[22] ), .A2(\a[31] ), .ZN(new_n2653_));
  INV_X1     g02429(.I(new_n2653_), .ZN(new_n2654_));
  INV_X1     g02430(.I(\a[31] ), .ZN(new_n2655_));
  NOR4_X1    g02431(.A1(new_n199_), .A2(new_n461_), .A3(new_n1313_), .A4(new_n2655_), .ZN(new_n2656_));
  NAND3_X1   g02432(.A1(new_n2656_), .A2(new_n403_), .A3(new_n2654_), .ZN(new_n2657_));
  AOI21_X1   g02433(.A1(new_n2657_), .A2(new_n1773_), .B(new_n525_), .ZN(new_n2658_));
  NOR3_X1    g02434(.A1(new_n2658_), .A2(new_n461_), .A3(new_n1313_), .ZN(new_n2659_));
  INV_X1     g02435(.I(new_n403_), .ZN(new_n2660_));
  OAI22_X1   g02436(.A1(new_n2660_), .A2(new_n2653_), .B1(new_n525_), .B2(new_n1773_), .ZN(new_n2661_));
  NOR3_X1    g02437(.A1(new_n2661_), .A2(new_n403_), .A3(new_n2654_), .ZN(new_n2662_));
  NOR2_X1    g02438(.A1(new_n2659_), .A2(new_n2662_), .ZN(new_n2663_));
  INV_X1     g02439(.I(new_n2663_), .ZN(new_n2664_));
  NOR2_X1    g02440(.A1(new_n199_), .A2(new_n2461_), .ZN(new_n2665_));
  OAI21_X1   g02441(.A1(new_n2465_), .A2(new_n2466_), .B(new_n2665_), .ZN(new_n2666_));
  NAND2_X1   g02442(.A1(new_n2666_), .A2(new_n2467_), .ZN(new_n2667_));
  NOR2_X1    g02443(.A1(new_n651_), .A2(new_n870_), .ZN(new_n2668_));
  INV_X1     g02444(.I(new_n2668_), .ZN(new_n2669_));
  NAND2_X1   g02445(.A1(new_n2392_), .A2(new_n2669_), .ZN(new_n2670_));
  NOR4_X1    g02446(.A1(new_n2670_), .A2(new_n1220_), .A3(new_n1316_), .A4(new_n2331_), .ZN(new_n2671_));
  XNOR2_X1   g02447(.A1(new_n2667_), .A2(new_n2671_), .ZN(new_n2672_));
  INV_X1     g02448(.I(new_n2667_), .ZN(new_n2673_));
  INV_X1     g02449(.I(new_n2671_), .ZN(new_n2674_));
  NOR2_X1    g02450(.A1(new_n2673_), .A2(new_n2674_), .ZN(new_n2675_));
  NOR2_X1    g02451(.A1(new_n2667_), .A2(new_n2671_), .ZN(new_n2676_));
  OAI21_X1   g02452(.A1(new_n2675_), .A2(new_n2676_), .B(new_n2664_), .ZN(new_n2677_));
  OAI21_X1   g02453(.A1(new_n2664_), .A2(new_n2672_), .B(new_n2677_), .ZN(new_n2678_));
  NAND2_X1   g02454(.A1(\a[24] ), .A2(\a[26] ), .ZN(new_n2679_));
  NAND2_X1   g02455(.A1(\a[23] ), .A2(\a[24] ), .ZN(new_n2680_));
  NOR2_X1    g02456(.A1(new_n1000_), .A2(new_n2679_), .ZN(new_n2682_));
  INV_X1     g02457(.I(new_n2682_), .ZN(new_n2683_));
  NAND2_X1   g02458(.A1(\a[14] ), .A2(\a[17] ), .ZN(new_n2684_));
  NAND4_X1   g02459(.A1(new_n1447_), .A2(new_n1275_), .A3(new_n1021_), .A4(new_n2684_), .ZN(new_n2685_));
  AND3_X2    g02460(.A1(new_n2685_), .A2(\a[6] ), .A3(\a[25] ), .Z(new_n2686_));
  AOI21_X1   g02461(.A1(\a[6] ), .A2(\a[25] ), .B(new_n2685_), .ZN(new_n2687_));
  NOR2_X1    g02462(.A1(new_n2686_), .A2(new_n2687_), .ZN(new_n2688_));
  NAND2_X1   g02463(.A1(\a[28] ), .A2(\a[29] ), .ZN(new_n2689_));
  INV_X1     g02464(.I(new_n2689_), .ZN(new_n2690_));
  AOI21_X1   g02465(.A1(new_n2500_), .A2(new_n2690_), .B(new_n1271_), .ZN(new_n2691_));
  NAND2_X1   g02466(.A1(\a[27] ), .A2(\a[28] ), .ZN(new_n2692_));
  NAND4_X1   g02467(.A1(new_n212_), .A2(new_n2692_), .A3(\a[2] ), .A4(\a[29] ), .ZN(new_n2693_));
  INV_X1     g02468(.I(new_n2693_), .ZN(new_n2694_));
  AND2_X2    g02469(.A1(new_n2691_), .A2(new_n2694_), .Z(new_n2695_));
  INV_X1     g02470(.I(new_n2695_), .ZN(new_n2696_));
  NOR2_X1    g02471(.A1(new_n2696_), .A2(new_n2688_), .ZN(new_n2697_));
  INV_X1     g02472(.I(new_n2697_), .ZN(new_n2698_));
  NAND2_X1   g02473(.A1(new_n2696_), .A2(new_n2688_), .ZN(new_n2699_));
  AOI21_X1   g02474(.A1(new_n2698_), .A2(new_n2699_), .B(new_n2683_), .ZN(new_n2700_));
  XOR2_X1    g02475(.A1(new_n2688_), .A2(new_n2695_), .Z(new_n2701_));
  NOR2_X1    g02476(.A1(new_n2701_), .A2(new_n2682_), .ZN(new_n2702_));
  NOR2_X1    g02477(.A1(new_n2702_), .A2(new_n2700_), .ZN(new_n2703_));
  XNOR2_X1   g02478(.A1(new_n2678_), .A2(new_n2703_), .ZN(new_n2704_));
  NOR2_X1    g02479(.A1(new_n2704_), .A2(new_n2652_), .ZN(new_n2705_));
  NOR2_X1    g02480(.A1(new_n2678_), .A2(new_n2703_), .ZN(new_n2706_));
  INV_X1     g02481(.I(new_n2706_), .ZN(new_n2707_));
  NAND2_X1   g02482(.A1(new_n2678_), .A2(new_n2703_), .ZN(new_n2708_));
  AOI21_X1   g02483(.A1(new_n2707_), .A2(new_n2708_), .B(new_n2651_), .ZN(new_n2709_));
  NOR2_X1    g02484(.A1(new_n2705_), .A2(new_n2709_), .ZN(new_n2710_));
  INV_X1     g02485(.I(new_n2710_), .ZN(new_n2711_));
  NAND3_X1   g02486(.A1(new_n2711_), .A2(new_n2649_), .A3(new_n2524_), .ZN(new_n2712_));
  INV_X1     g02487(.I(new_n2524_), .ZN(new_n2713_));
  AOI21_X1   g02488(.A1(new_n2481_), .A2(new_n2519_), .B(new_n2457_), .ZN(new_n2714_));
  OAI21_X1   g02489(.A1(new_n2714_), .A2(new_n2713_), .B(new_n2710_), .ZN(new_n2715_));
  AOI22_X1   g02490(.A1(new_n2644_), .A2(new_n2648_), .B1(new_n2715_), .B2(new_n2712_), .ZN(new_n2716_));
  NAND2_X1   g02491(.A1(new_n2644_), .A2(new_n2648_), .ZN(new_n2717_));
  AOI21_X1   g02492(.A1(new_n2649_), .A2(new_n2524_), .B(new_n2710_), .ZN(new_n2718_));
  NOR3_X1    g02493(.A1(new_n2711_), .A2(new_n2714_), .A3(new_n2713_), .ZN(new_n2719_));
  NOR2_X1    g02494(.A1(new_n2719_), .A2(new_n2718_), .ZN(new_n2720_));
  NOR2_X1    g02495(.A1(new_n2717_), .A2(new_n2720_), .ZN(new_n2721_));
  NOR2_X1    g02496(.A1(new_n2721_), .A2(new_n2716_), .ZN(new_n2722_));
  INV_X1     g02497(.I(new_n2568_), .ZN(new_n2723_));
  AOI21_X1   g02498(.A1(new_n2723_), .A2(new_n2574_), .B(new_n2572_), .ZN(new_n2724_));
  INV_X1     g02499(.I(new_n2724_), .ZN(new_n2725_));
  XOR2_X1    g02500(.A1(new_n2722_), .A2(new_n2725_), .Z(new_n2726_));
  NAND2_X1   g02501(.A1(new_n2587_), .A2(new_n2726_), .ZN(new_n2727_));
  NOR3_X1    g02502(.A1(new_n2721_), .A2(new_n2716_), .A3(new_n2724_), .ZN(new_n2728_));
  NOR2_X1    g02503(.A1(new_n2722_), .A2(new_n2725_), .ZN(new_n2729_));
  NOR2_X1    g02504(.A1(new_n2729_), .A2(new_n2728_), .ZN(new_n2730_));
  OAI21_X1   g02505(.A1(new_n2587_), .A2(new_n2730_), .B(new_n2727_), .ZN(\asquared[32] ));
  NOR2_X1    g02506(.A1(new_n2728_), .A2(new_n2578_), .ZN(new_n2732_));
  AOI21_X1   g02507(.A1(new_n2728_), .A2(new_n2578_), .B(new_n2454_), .ZN(new_n2733_));
  NOR2_X1    g02508(.A1(new_n2733_), .A2(new_n2732_), .ZN(new_n2734_));
  OAI21_X1   g02509(.A1(new_n2451_), .A2(new_n2446_), .B(new_n2734_), .ZN(new_n2735_));
  INV_X1     g02510(.I(new_n2717_), .ZN(new_n2736_));
  INV_X1     g02511(.I(new_n2715_), .ZN(new_n2737_));
  AOI21_X1   g02512(.A1(new_n2736_), .A2(new_n2712_), .B(new_n2737_), .ZN(new_n2738_));
  INV_X1     g02513(.I(new_n2738_), .ZN(new_n2739_));
  INV_X1     g02514(.I(new_n2647_), .ZN(new_n2740_));
  OAI21_X1   g02515(.A1(new_n2640_), .A2(new_n2614_), .B(new_n2588_), .ZN(new_n2741_));
  NAND2_X1   g02516(.A1(new_n2740_), .A2(new_n2741_), .ZN(new_n2742_));
  NAND2_X1   g02517(.A1(new_n2609_), .A2(new_n2612_), .ZN(new_n2743_));
  NAND2_X1   g02518(.A1(new_n2743_), .A2(new_n2610_), .ZN(new_n2744_));
  NOR2_X1    g02519(.A1(new_n2624_), .A2(new_n2464_), .ZN(new_n2745_));
  XOR2_X1    g02520(.A1(new_n2625_), .A2(\a[16] ), .Z(new_n2746_));
  AOI21_X1   g02521(.A1(new_n2624_), .A2(new_n2464_), .B(new_n2746_), .ZN(new_n2747_));
  NOR2_X1    g02522(.A1(new_n2747_), .A2(new_n2745_), .ZN(new_n2748_));
  NOR2_X1    g02523(.A1(new_n2276_), .A2(new_n2679_), .ZN(new_n2749_));
  NOR2_X1    g02524(.A1(new_n341_), .A2(new_n392_), .ZN(new_n2750_));
  NOR2_X1    g02525(.A1(new_n2749_), .A2(new_n2750_), .ZN(new_n2751_));
  NOR2_X1    g02526(.A1(new_n1999_), .A2(new_n1916_), .ZN(new_n2752_));
  INV_X1     g02527(.I(new_n2752_), .ZN(new_n2753_));
  NAND4_X1   g02528(.A1(new_n2753_), .A2(\a[8] ), .A3(\a[24] ), .A4(new_n478_), .ZN(new_n2754_));
  INV_X1     g02529(.I(new_n2754_), .ZN(new_n2755_));
  NAND2_X1   g02530(.A1(new_n2755_), .A2(new_n2751_), .ZN(new_n2756_));
  NOR2_X1    g02531(.A1(new_n364_), .A2(new_n2368_), .ZN(new_n2757_));
  XNOR2_X1   g02532(.A1(new_n211_), .A2(new_n2692_), .ZN(new_n2758_));
  INV_X1     g02533(.I(new_n2758_), .ZN(new_n2759_));
  XOR2_X1    g02534(.A1(new_n2756_), .A2(new_n2759_), .Z(new_n2760_));
  NOR2_X1    g02535(.A1(new_n2756_), .A2(new_n2758_), .ZN(new_n2761_));
  AOI21_X1   g02536(.A1(new_n2755_), .A2(new_n2751_), .B(new_n2759_), .ZN(new_n2762_));
  OAI21_X1   g02537(.A1(new_n2761_), .A2(new_n2762_), .B(new_n2748_), .ZN(new_n2763_));
  OAI21_X1   g02538(.A1(new_n2760_), .A2(new_n2748_), .B(new_n2763_), .ZN(new_n2764_));
  INV_X1     g02539(.I(\a[32] ), .ZN(new_n2765_));
  NOR2_X1    g02540(.A1(new_n2461_), .A2(new_n2765_), .ZN(new_n2766_));
  NOR2_X1    g02541(.A1(new_n2625_), .A2(new_n800_), .ZN(new_n2767_));
  XOR2_X1    g02542(.A1(new_n2766_), .A2(new_n197_), .Z(new_n2768_));
  INV_X1     g02543(.I(new_n1712_), .ZN(new_n2769_));
  NAND2_X1   g02544(.A1(new_n2769_), .A2(new_n2669_), .ZN(new_n2770_));
  NOR2_X1    g02545(.A1(new_n675_), .A2(new_n1313_), .ZN(new_n2771_));
  INV_X1     g02546(.I(new_n2771_), .ZN(new_n2772_));
  NOR4_X1    g02547(.A1(new_n2770_), .A2(new_n1220_), .A3(new_n1798_), .A4(new_n2772_), .ZN(new_n2773_));
  INV_X1     g02548(.I(new_n2773_), .ZN(new_n2774_));
  NAND4_X1   g02549(.A1(\a[3] ), .A2(\a[10] ), .A3(\a[22] ), .A4(\a[29] ), .ZN(new_n2775_));
  XOR2_X1    g02550(.A1(new_n2775_), .A2(\a[14] ), .Z(new_n2776_));
  XOR2_X1    g02551(.A1(new_n2776_), .A2(\a[18] ), .Z(new_n2777_));
  NOR2_X1    g02552(.A1(new_n2777_), .A2(new_n2774_), .ZN(new_n2778_));
  INV_X1     g02553(.I(new_n2778_), .ZN(new_n2779_));
  NAND2_X1   g02554(.A1(new_n2777_), .A2(new_n2774_), .ZN(new_n2780_));
  AOI21_X1   g02555(.A1(new_n2779_), .A2(new_n2780_), .B(new_n2768_), .ZN(new_n2781_));
  XOR2_X1    g02556(.A1(new_n2777_), .A2(new_n2773_), .Z(new_n2782_));
  INV_X1     g02557(.I(new_n2782_), .ZN(new_n2783_));
  AOI21_X1   g02558(.A1(new_n2783_), .A2(new_n2768_), .B(new_n2781_), .ZN(new_n2784_));
  XNOR2_X1   g02559(.A1(new_n2784_), .A2(new_n2764_), .ZN(new_n2785_));
  INV_X1     g02560(.I(new_n2785_), .ZN(new_n2786_));
  NOR2_X1    g02561(.A1(new_n2784_), .A2(new_n2764_), .ZN(new_n2787_));
  NAND2_X1   g02562(.A1(new_n2784_), .A2(new_n2764_), .ZN(new_n2788_));
  INV_X1     g02563(.I(new_n2788_), .ZN(new_n2789_));
  NOR2_X1    g02564(.A1(new_n2789_), .A2(new_n2787_), .ZN(new_n2790_));
  NOR2_X1    g02565(.A1(new_n2744_), .A2(new_n2790_), .ZN(new_n2791_));
  AOI21_X1   g02566(.A1(new_n2744_), .A2(new_n2786_), .B(new_n2791_), .ZN(new_n2792_));
  INV_X1     g02567(.I(new_n2792_), .ZN(new_n2793_));
  NOR2_X1    g02568(.A1(new_n2632_), .A2(new_n2621_), .ZN(new_n2794_));
  AOI21_X1   g02569(.A1(new_n2632_), .A2(new_n2621_), .B(new_n2619_), .ZN(new_n2795_));
  NOR2_X1    g02570(.A1(new_n2795_), .A2(new_n2794_), .ZN(new_n2796_));
  INV_X1     g02571(.I(new_n2692_), .ZN(new_n2797_));
  AOI21_X1   g02572(.A1(new_n267_), .A2(new_n2797_), .B(new_n2691_), .ZN(new_n2798_));
  AOI22_X1   g02573(.A1(new_n2392_), .A2(new_n2669_), .B1(new_n1220_), .B2(new_n2331_), .ZN(new_n2799_));
  XOR2_X1    g02574(.A1(new_n2798_), .A2(new_n2799_), .Z(new_n2800_));
  INV_X1     g02575(.I(new_n2800_), .ZN(new_n2801_));
  NAND2_X1   g02576(.A1(new_n2798_), .A2(new_n2799_), .ZN(new_n2802_));
  INV_X1     g02577(.I(new_n2802_), .ZN(new_n2803_));
  NOR2_X1    g02578(.A1(new_n2798_), .A2(new_n2799_), .ZN(new_n2804_));
  OAI21_X1   g02579(.A1(new_n2803_), .A2(new_n2804_), .B(new_n2661_), .ZN(new_n2805_));
  OAI21_X1   g02580(.A1(new_n2801_), .A2(new_n2661_), .B(new_n2805_), .ZN(new_n2806_));
  OAI22_X1   g02581(.A1(new_n392_), .A2(new_n2680_), .B1(new_n1000_), .B2(new_n2679_), .ZN(new_n2807_));
  INV_X1     g02582(.I(new_n2807_), .ZN(new_n2808_));
  NAND2_X1   g02583(.A1(new_n1447_), .A2(new_n1275_), .ZN(new_n2809_));
  NAND2_X1   g02584(.A1(new_n1021_), .A2(new_n2684_), .ZN(new_n2810_));
  NOR2_X1    g02585(.A1(\a[6] ), .A2(\a[25] ), .ZN(new_n2811_));
  AOI21_X1   g02586(.A1(new_n2809_), .A2(new_n2811_), .B(new_n2810_), .ZN(new_n2812_));
  NOR2_X1    g02587(.A1(new_n194_), .A2(new_n2655_), .ZN(new_n2813_));
  XOR2_X1    g02588(.A1(new_n2813_), .A2(new_n1141_), .Z(new_n2814_));
  XOR2_X1    g02589(.A1(new_n2814_), .A2(new_n2812_), .Z(new_n2815_));
  NOR2_X1    g02590(.A1(new_n2814_), .A2(new_n2812_), .ZN(new_n2816_));
  INV_X1     g02591(.I(new_n2816_), .ZN(new_n2817_));
  NAND2_X1   g02592(.A1(new_n2814_), .A2(new_n2812_), .ZN(new_n2818_));
  AOI21_X1   g02593(.A1(new_n2817_), .A2(new_n2818_), .B(new_n2808_), .ZN(new_n2819_));
  AOI21_X1   g02594(.A1(new_n2808_), .A2(new_n2815_), .B(new_n2819_), .ZN(new_n2820_));
  XOR2_X1    g02595(.A1(new_n2806_), .A2(new_n2820_), .Z(new_n2821_));
  NOR2_X1    g02596(.A1(new_n2796_), .A2(new_n2821_), .ZN(new_n2822_));
  INV_X1     g02597(.I(new_n2820_), .ZN(new_n2823_));
  NAND2_X1   g02598(.A1(new_n2806_), .A2(new_n2823_), .ZN(new_n2824_));
  NOR2_X1    g02599(.A1(new_n2806_), .A2(new_n2823_), .ZN(new_n2825_));
  INV_X1     g02600(.I(new_n2825_), .ZN(new_n2826_));
  NAND2_X1   g02601(.A1(new_n2826_), .A2(new_n2824_), .ZN(new_n2827_));
  AOI21_X1   g02602(.A1(new_n2796_), .A2(new_n2827_), .B(new_n2822_), .ZN(new_n2828_));
  INV_X1     g02603(.I(new_n2676_), .ZN(new_n2829_));
  AOI21_X1   g02604(.A1(new_n2663_), .A2(new_n2829_), .B(new_n2675_), .ZN(new_n2830_));
  INV_X1     g02605(.I(new_n2830_), .ZN(new_n2831_));
  AOI21_X1   g02606(.A1(new_n2696_), .A2(new_n2688_), .B(new_n2683_), .ZN(new_n2832_));
  NOR2_X1    g02607(.A1(new_n2832_), .A2(new_n2697_), .ZN(new_n2833_));
  NOR2_X1    g02608(.A1(new_n2602_), .A2(new_n2593_), .ZN(new_n2834_));
  NOR2_X1    g02609(.A1(new_n2834_), .A2(new_n2601_), .ZN(new_n2835_));
  XOR2_X1    g02610(.A1(new_n2835_), .A2(new_n2833_), .Z(new_n2836_));
  NAND2_X1   g02611(.A1(new_n2836_), .A2(new_n2831_), .ZN(new_n2837_));
  NOR2_X1    g02612(.A1(new_n2835_), .A2(new_n2833_), .ZN(new_n2838_));
  NOR4_X1    g02613(.A1(new_n2834_), .A2(new_n2601_), .A3(new_n2697_), .A4(new_n2832_), .ZN(new_n2839_));
  OAI21_X1   g02614(.A1(new_n2838_), .A2(new_n2839_), .B(new_n2830_), .ZN(new_n2840_));
  NAND2_X1   g02615(.A1(new_n2837_), .A2(new_n2840_), .ZN(new_n2841_));
  AOI21_X1   g02616(.A1(new_n2651_), .A2(new_n2708_), .B(new_n2706_), .ZN(new_n2842_));
  OR2_X2     g02617(.A1(new_n2842_), .A2(new_n2841_), .Z(new_n2843_));
  NAND2_X1   g02618(.A1(new_n2842_), .A2(new_n2841_), .ZN(new_n2844_));
  AOI21_X1   g02619(.A1(new_n2843_), .A2(new_n2844_), .B(new_n2828_), .ZN(new_n2845_));
  INV_X1     g02620(.I(new_n2828_), .ZN(new_n2846_));
  XNOR2_X1   g02621(.A1(new_n2842_), .A2(new_n2841_), .ZN(new_n2847_));
  NOR2_X1    g02622(.A1(new_n2846_), .A2(new_n2847_), .ZN(new_n2848_));
  NOR2_X1    g02623(.A1(new_n2848_), .A2(new_n2845_), .ZN(new_n2849_));
  NOR2_X1    g02624(.A1(new_n2849_), .A2(new_n2793_), .ZN(new_n2850_));
  INV_X1     g02625(.I(new_n2849_), .ZN(new_n2851_));
  NOR2_X1    g02626(.A1(new_n2851_), .A2(new_n2792_), .ZN(new_n2852_));
  OAI21_X1   g02627(.A1(new_n2852_), .A2(new_n2850_), .B(new_n2742_), .ZN(new_n2853_));
  INV_X1     g02628(.I(new_n2853_), .ZN(new_n2854_));
  INV_X1     g02629(.I(new_n2742_), .ZN(new_n2855_));
  NOR2_X1    g02630(.A1(new_n2849_), .A2(new_n2792_), .ZN(new_n2856_));
  NOR2_X1    g02631(.A1(new_n2851_), .A2(new_n2793_), .ZN(new_n2857_));
  OAI21_X1   g02632(.A1(new_n2857_), .A2(new_n2856_), .B(new_n2855_), .ZN(new_n2858_));
  INV_X1     g02633(.I(new_n2858_), .ZN(new_n2859_));
  OAI21_X1   g02634(.A1(new_n2854_), .A2(new_n2859_), .B(new_n2739_), .ZN(new_n2860_));
  XOR2_X1    g02635(.A1(new_n2735_), .A2(new_n2860_), .Z(new_n2861_));
  XOR2_X1    g02636(.A1(new_n2861_), .A2(new_n2729_), .Z(\asquared[33] ));
  NAND3_X1   g02637(.A1(new_n2853_), .A2(new_n2858_), .A3(new_n2738_), .ZN(new_n2863_));
  NAND2_X1   g02638(.A1(new_n2863_), .A2(new_n2729_), .ZN(new_n2864_));
  OAI21_X1   g02639(.A1(new_n2735_), .A2(new_n2864_), .B(new_n2860_), .ZN(new_n2865_));
  AOI21_X1   g02640(.A1(new_n2744_), .A2(new_n2788_), .B(new_n2787_), .ZN(new_n2866_));
  INV_X1     g02641(.I(new_n2866_), .ZN(new_n2867_));
  INV_X1     g02642(.I(\a[33] ), .ZN(new_n2868_));
  NOR2_X1    g02643(.A1(new_n2655_), .A2(new_n2868_), .ZN(new_n2869_));
  INV_X1     g02644(.I(new_n2869_), .ZN(new_n2870_));
  NAND2_X1   g02645(.A1(\a[22] ), .A2(\a[33] ), .ZN(new_n2871_));
  NOR2_X1    g02646(.A1(new_n483_), .A2(new_n2871_), .ZN(new_n2872_));
  NOR2_X1    g02647(.A1(new_n610_), .A2(new_n2653_), .ZN(new_n2873_));
  NAND2_X1   g02648(.A1(new_n2872_), .A2(new_n2873_), .ZN(new_n2874_));
  AOI21_X1   g02649(.A1(new_n2874_), .A2(new_n2870_), .B(new_n197_), .ZN(new_n2875_));
  NOR3_X1    g02650(.A1(new_n2875_), .A2(new_n201_), .A3(new_n2655_), .ZN(new_n2876_));
  OAI22_X1   g02651(.A1(new_n2870_), .A2(new_n197_), .B1(new_n483_), .B2(new_n2871_), .ZN(new_n2877_));
  INV_X1     g02652(.I(new_n2877_), .ZN(new_n2878_));
  AND3_X2    g02653(.A1(new_n2878_), .A2(new_n483_), .A3(new_n2871_), .Z(new_n2879_));
  NOR2_X1    g02654(.A1(new_n2879_), .A2(new_n2876_), .ZN(new_n2880_));
  OAI22_X1   g02655(.A1(new_n2753_), .A2(new_n478_), .B1(new_n2749_), .B2(new_n2750_), .ZN(new_n2881_));
  AOI21_X1   g02656(.A1(new_n229_), .A2(new_n2757_), .B(new_n2797_), .ZN(new_n2882_));
  NOR2_X1    g02657(.A1(new_n2881_), .A2(new_n2882_), .ZN(new_n2883_));
  INV_X1     g02658(.I(new_n2883_), .ZN(new_n2884_));
  NAND2_X1   g02659(.A1(new_n2881_), .A2(new_n2882_), .ZN(new_n2885_));
  NAND2_X1   g02660(.A1(new_n2884_), .A2(new_n2885_), .ZN(new_n2886_));
  XNOR2_X1   g02661(.A1(new_n2881_), .A2(new_n2882_), .ZN(new_n2887_));
  NOR2_X1    g02662(.A1(new_n2880_), .A2(new_n2887_), .ZN(new_n2888_));
  AOI21_X1   g02663(.A1(new_n2880_), .A2(new_n2886_), .B(new_n2888_), .ZN(new_n2889_));
  NOR2_X1    g02664(.A1(new_n1999_), .A2(new_n2098_), .ZN(new_n2890_));
  INV_X1     g02665(.I(new_n2890_), .ZN(new_n2891_));
  NOR2_X1    g02666(.A1(new_n353_), .A2(new_n2178_), .ZN(new_n2892_));
  NOR2_X1    g02667(.A1(new_n2891_), .A2(new_n341_), .ZN(new_n2896_));
  INV_X1     g02668(.I(new_n2896_), .ZN(new_n2897_));
  NOR2_X1    g02669(.A1(new_n2499_), .A2(new_n2461_), .ZN(new_n2898_));
  NOR2_X1    g02670(.A1(new_n1691_), .A2(new_n2461_), .ZN(new_n2899_));
  AOI22_X1   g02671(.A1(new_n524_), .A2(new_n2898_), .B1(new_n2899_), .B2(new_n267_), .ZN(new_n2900_));
  NAND2_X1   g02672(.A1(\a[4] ), .A2(\a[29] ), .ZN(new_n2901_));
  INV_X1     g02673(.I(new_n2901_), .ZN(new_n2902_));
  NAND2_X1   g02674(.A1(\a[9] ), .A2(\a[24] ), .ZN(new_n2903_));
  OAI21_X1   g02675(.A1(new_n2902_), .A2(new_n2903_), .B(new_n2900_), .ZN(new_n2904_));
  XNOR2_X1   g02676(.A1(new_n2901_), .A2(new_n2903_), .ZN(new_n2905_));
  NAND2_X1   g02677(.A1(\a[3] ), .A2(\a[30] ), .ZN(new_n2906_));
  NAND2_X1   g02678(.A1(new_n2905_), .A2(new_n2906_), .ZN(new_n2907_));
  NOR2_X1    g02679(.A1(new_n1021_), .A2(new_n1268_), .ZN(new_n2908_));
  AOI21_X1   g02680(.A1(\a[15] ), .A2(\a[18] ), .B(new_n1275_), .ZN(new_n2909_));
  NAND2_X1   g02681(.A1(new_n2909_), .A2(new_n2908_), .ZN(new_n2910_));
  NAND2_X1   g02682(.A1(\a[7] ), .A2(\a[26] ), .ZN(new_n2911_));
  XOR2_X1    g02683(.A1(new_n2910_), .A2(new_n2911_), .Z(new_n2912_));
  NAND3_X1   g02684(.A1(new_n2912_), .A2(new_n2904_), .A3(new_n2907_), .ZN(new_n2913_));
  NAND2_X1   g02685(.A1(new_n2904_), .A2(new_n2907_), .ZN(new_n2914_));
  INV_X1     g02686(.I(new_n2912_), .ZN(new_n2915_));
  NAND2_X1   g02687(.A1(new_n2915_), .A2(new_n2914_), .ZN(new_n2916_));
  AOI21_X1   g02688(.A1(new_n2916_), .A2(new_n2913_), .B(new_n2897_), .ZN(new_n2917_));
  XOR2_X1    g02689(.A1(new_n2912_), .A2(new_n2914_), .Z(new_n2918_));
  NOR2_X1    g02690(.A1(new_n2918_), .A2(new_n2896_), .ZN(new_n2919_));
  NOR2_X1    g02691(.A1(new_n2919_), .A2(new_n2917_), .ZN(new_n2920_));
  AOI21_X1   g02692(.A1(new_n2767_), .A2(new_n218_), .B(new_n2766_), .ZN(new_n2921_));
  OAI21_X1   g02693(.A1(new_n1150_), .A2(new_n1715_), .B(new_n2770_), .ZN(new_n2922_));
  INV_X1     g02694(.I(new_n2775_), .ZN(new_n2923_));
  AOI22_X1   g02695(.A1(\a[3] ), .A2(\a[29] ), .B1(\a[10] ), .B2(\a[22] ), .ZN(new_n2924_));
  NOR3_X1    g02696(.A1(new_n2924_), .A2(new_n650_), .A3(new_n1276_), .ZN(new_n2925_));
  NOR2_X1    g02697(.A1(new_n2925_), .A2(new_n2923_), .ZN(new_n2926_));
  INV_X1     g02698(.I(new_n2926_), .ZN(new_n2927_));
  XOR2_X1    g02699(.A1(new_n2922_), .A2(new_n2927_), .Z(new_n2928_));
  NOR2_X1    g02700(.A1(new_n2928_), .A2(new_n2921_), .ZN(new_n2929_));
  INV_X1     g02701(.I(new_n2921_), .ZN(new_n2930_));
  NOR2_X1    g02702(.A1(new_n2922_), .A2(new_n2926_), .ZN(new_n2931_));
  INV_X1     g02703(.I(new_n2931_), .ZN(new_n2932_));
  NAND2_X1   g02704(.A1(new_n2922_), .A2(new_n2926_), .ZN(new_n2933_));
  AOI21_X1   g02705(.A1(new_n2932_), .A2(new_n2933_), .B(new_n2930_), .ZN(new_n2934_));
  NOR2_X1    g02706(.A1(new_n2929_), .A2(new_n2934_), .ZN(new_n2935_));
  INV_X1     g02707(.I(new_n2935_), .ZN(new_n2936_));
  NAND2_X1   g02708(.A1(new_n2920_), .A2(new_n2936_), .ZN(new_n2937_));
  NOR2_X1    g02709(.A1(new_n2920_), .A2(new_n2936_), .ZN(new_n2938_));
  INV_X1     g02710(.I(new_n2938_), .ZN(new_n2939_));
  AOI21_X1   g02711(.A1(new_n2939_), .A2(new_n2937_), .B(new_n2889_), .ZN(new_n2940_));
  INV_X1     g02712(.I(new_n2889_), .ZN(new_n2941_));
  XOR2_X1    g02713(.A1(new_n2920_), .A2(new_n2935_), .Z(new_n2942_));
  NOR2_X1    g02714(.A1(new_n2942_), .A2(new_n2941_), .ZN(new_n2943_));
  NOR2_X1    g02715(.A1(new_n2943_), .A2(new_n2940_), .ZN(new_n2944_));
  OAI21_X1   g02716(.A1(new_n2661_), .A2(new_n2804_), .B(new_n2802_), .ZN(new_n2945_));
  NOR2_X1    g02717(.A1(new_n2748_), .A2(new_n2762_), .ZN(new_n2946_));
  NOR2_X1    g02718(.A1(new_n2946_), .A2(new_n2761_), .ZN(new_n2947_));
  AOI21_X1   g02719(.A1(new_n2777_), .A2(new_n2774_), .B(new_n2768_), .ZN(new_n2948_));
  NOR2_X1    g02720(.A1(new_n2948_), .A2(new_n2778_), .ZN(new_n2949_));
  XOR2_X1    g02721(.A1(new_n2949_), .A2(new_n2947_), .Z(new_n2950_));
  NAND2_X1   g02722(.A1(new_n2950_), .A2(new_n2945_), .ZN(new_n2951_));
  INV_X1     g02723(.I(new_n2945_), .ZN(new_n2952_));
  NOR2_X1    g02724(.A1(new_n2949_), .A2(new_n2947_), .ZN(new_n2953_));
  NOR4_X1    g02725(.A1(new_n2948_), .A2(new_n2778_), .A3(new_n2761_), .A4(new_n2946_), .ZN(new_n2954_));
  OAI21_X1   g02726(.A1(new_n2953_), .A2(new_n2954_), .B(new_n2952_), .ZN(new_n2955_));
  NAND2_X1   g02727(.A1(new_n2951_), .A2(new_n2955_), .ZN(new_n2956_));
  XOR2_X1    g02728(.A1(new_n2944_), .A2(new_n2956_), .Z(new_n2957_));
  AND2_X2    g02729(.A1(new_n2957_), .A2(new_n2867_), .Z(new_n2958_));
  NAND2_X1   g02730(.A1(new_n2944_), .A2(new_n2956_), .ZN(new_n2959_));
  NOR2_X1    g02731(.A1(new_n2944_), .A2(new_n2956_), .ZN(new_n2960_));
  INV_X1     g02732(.I(new_n2960_), .ZN(new_n2961_));
  AOI21_X1   g02733(.A1(new_n2961_), .A2(new_n2959_), .B(new_n2867_), .ZN(new_n2962_));
  NOR2_X1    g02734(.A1(new_n2839_), .A2(new_n2830_), .ZN(new_n2963_));
  NOR2_X1    g02735(.A1(new_n2963_), .A2(new_n2838_), .ZN(new_n2964_));
  OR2_X2     g02736(.A1(new_n2795_), .A2(new_n2794_), .Z(new_n2965_));
  AOI21_X1   g02737(.A1(new_n2965_), .A2(new_n2824_), .B(new_n2825_), .ZN(new_n2966_));
  INV_X1     g02738(.I(new_n2966_), .ZN(new_n2967_));
  OAI21_X1   g02739(.A1(new_n2807_), .A2(new_n2816_), .B(new_n2818_), .ZN(new_n2968_));
  NAND2_X1   g02740(.A1(new_n2813_), .A2(new_n1143_), .ZN(new_n2969_));
  NAND2_X1   g02741(.A1(\a[1] ), .A2(\a[32] ), .ZN(new_n2970_));
  NOR2_X1    g02742(.A1(new_n2970_), .A2(new_n885_), .ZN(new_n2971_));
  INV_X1     g02743(.I(new_n2970_), .ZN(new_n2972_));
  NOR2_X1    g02744(.A1(new_n2972_), .A2(\a[17] ), .ZN(new_n2973_));
  NOR2_X1    g02745(.A1(new_n2973_), .A2(new_n2971_), .ZN(new_n2974_));
  NOR2_X1    g02746(.A1(new_n2974_), .A2(new_n2969_), .ZN(new_n2975_));
  XOR2_X1    g02747(.A1(new_n2975_), .A2(new_n461_), .Z(new_n2976_));
  XOR2_X1    g02748(.A1(new_n2976_), .A2(new_n2368_), .Z(new_n2977_));
  INV_X1     g02749(.I(new_n1711_), .ZN(new_n2978_));
  AOI22_X1   g02750(.A1(new_n654_), .A2(new_n2978_), .B1(new_n1220_), .B2(new_n1769_), .ZN(new_n2979_));
  NOR2_X1    g02751(.A1(new_n566_), .A2(new_n1313_), .ZN(new_n2980_));
  NAND4_X1   g02752(.A1(new_n2979_), .A2(new_n786_), .A3(new_n1715_), .A4(new_n2980_), .ZN(new_n2981_));
  INV_X1     g02753(.I(new_n2981_), .ZN(new_n2982_));
  XOR2_X1    g02754(.A1(new_n2977_), .A2(new_n2982_), .Z(new_n2983_));
  NAND2_X1   g02755(.A1(new_n2983_), .A2(new_n2968_), .ZN(new_n2984_));
  INV_X1     g02756(.I(new_n2977_), .ZN(new_n2985_));
  NOR2_X1    g02757(.A1(new_n2985_), .A2(new_n2981_), .ZN(new_n2986_));
  NOR2_X1    g02758(.A1(new_n2977_), .A2(new_n2982_), .ZN(new_n2987_));
  NOR2_X1    g02759(.A1(new_n2986_), .A2(new_n2987_), .ZN(new_n2988_));
  OAI21_X1   g02760(.A1(new_n2968_), .A2(new_n2988_), .B(new_n2984_), .ZN(new_n2989_));
  NAND2_X1   g02761(.A1(new_n2967_), .A2(new_n2989_), .ZN(new_n2990_));
  INV_X1     g02762(.I(new_n2989_), .ZN(new_n2991_));
  NAND2_X1   g02763(.A1(new_n2991_), .A2(new_n2966_), .ZN(new_n2992_));
  AOI21_X1   g02764(.A1(new_n2990_), .A2(new_n2992_), .B(new_n2964_), .ZN(new_n2993_));
  INV_X1     g02765(.I(new_n2964_), .ZN(new_n2994_));
  NAND2_X1   g02766(.A1(new_n2966_), .A2(new_n2989_), .ZN(new_n2995_));
  NOR2_X1    g02767(.A1(new_n2966_), .A2(new_n2989_), .ZN(new_n2996_));
  INV_X1     g02768(.I(new_n2996_), .ZN(new_n2997_));
  AOI21_X1   g02769(.A1(new_n2997_), .A2(new_n2995_), .B(new_n2994_), .ZN(new_n2998_));
  NAND2_X1   g02770(.A1(new_n2828_), .A2(new_n2844_), .ZN(new_n2999_));
  NAND2_X1   g02771(.A1(new_n2999_), .A2(new_n2843_), .ZN(new_n3000_));
  INV_X1     g02772(.I(new_n3000_), .ZN(new_n3001_));
  NOR3_X1    g02773(.A1(new_n3001_), .A2(new_n2993_), .A3(new_n2998_), .ZN(new_n3002_));
  OAI21_X1   g02774(.A1(new_n2993_), .A2(new_n2998_), .B(new_n3001_), .ZN(new_n3003_));
  INV_X1     g02775(.I(new_n3003_), .ZN(new_n3004_));
  OAI22_X1   g02776(.A1(new_n3004_), .A2(new_n3002_), .B1(new_n2958_), .B2(new_n2962_), .ZN(new_n3005_));
  AOI21_X1   g02777(.A1(new_n2957_), .A2(new_n2867_), .B(new_n2962_), .ZN(new_n3006_));
  NOR2_X1    g02778(.A1(new_n2998_), .A2(new_n2993_), .ZN(new_n3007_));
  NOR2_X1    g02779(.A1(new_n3007_), .A2(new_n3001_), .ZN(new_n3008_));
  NOR3_X1    g02780(.A1(new_n2998_), .A2(new_n2993_), .A3(new_n3000_), .ZN(new_n3009_));
  OAI21_X1   g02781(.A1(new_n3008_), .A2(new_n3009_), .B(new_n3006_), .ZN(new_n3010_));
  NAND2_X1   g02782(.A1(new_n3005_), .A2(new_n3010_), .ZN(new_n3011_));
  INV_X1     g02783(.I(new_n2857_), .ZN(new_n3012_));
  OAI21_X1   g02784(.A1(new_n2855_), .A2(new_n2856_), .B(new_n3012_), .ZN(new_n3013_));
  XNOR2_X1   g02785(.A1(new_n3011_), .A2(new_n3013_), .ZN(new_n3014_));
  NAND3_X1   g02786(.A1(new_n3005_), .A2(new_n3010_), .A3(new_n3013_), .ZN(new_n3015_));
  INV_X1     g02787(.I(new_n3013_), .ZN(new_n3016_));
  NAND2_X1   g02788(.A1(new_n3016_), .A2(new_n3011_), .ZN(new_n3017_));
  NAND2_X1   g02789(.A1(new_n3017_), .A2(new_n3015_), .ZN(new_n3018_));
  MUX2_X1    g02790(.I0(new_n3018_), .I1(new_n3014_), .S(new_n2865_), .Z(\asquared[34] ));
  NAND2_X1   g02791(.A1(new_n2865_), .A2(new_n3017_), .ZN(new_n3020_));
  NAND2_X1   g02792(.A1(new_n3020_), .A2(new_n3015_), .ZN(new_n3021_));
  AOI21_X1   g02793(.A1(new_n3006_), .A2(new_n3003_), .B(new_n3002_), .ZN(new_n3022_));
  NAND2_X1   g02794(.A1(\a[9] ), .A2(\a[29] ), .ZN(new_n3023_));
  NOR2_X1    g02795(.A1(new_n2545_), .A2(new_n3023_), .ZN(new_n3024_));
  NAND2_X1   g02796(.A1(\a[5] ), .A2(\a[10] ), .ZN(new_n3025_));
  NOR3_X1    g02797(.A1(new_n3025_), .A2(new_n1691_), .A3(new_n2499_), .ZN(new_n3026_));
  NAND2_X1   g02798(.A1(new_n3026_), .A2(new_n3024_), .ZN(new_n3027_));
  AOI21_X1   g02799(.A1(new_n3027_), .A2(new_n525_), .B(new_n2276_), .ZN(new_n3028_));
  NOR3_X1    g02800(.A1(new_n3028_), .A2(new_n461_), .A3(new_n1691_), .ZN(new_n3029_));
  OAI22_X1   g02801(.A1(new_n525_), .A2(new_n2276_), .B1(new_n2545_), .B2(new_n3023_), .ZN(new_n3030_));
  OAI22_X1   g02802(.A1(new_n353_), .A2(new_n364_), .B1(new_n1999_), .B2(new_n2499_), .ZN(new_n3031_));
  NOR2_X1    g02803(.A1(new_n3030_), .A2(new_n3031_), .ZN(new_n3032_));
  NOR2_X1    g02804(.A1(new_n3029_), .A2(new_n3032_), .ZN(new_n3033_));
  OAI21_X1   g02805(.A1(new_n786_), .A2(new_n873_), .B(new_n2769_), .ZN(new_n3034_));
  NAND4_X1   g02806(.A1(new_n1018_), .A2(new_n1715_), .A3(\a[13] ), .A4(\a[21] ), .ZN(new_n3035_));
  NAND2_X1   g02807(.A1(\a[26] ), .A2(\a[28] ), .ZN(new_n3036_));
  INV_X1     g02808(.I(new_n3036_), .ZN(new_n3037_));
  NAND2_X1   g02809(.A1(new_n2797_), .A2(new_n3037_), .ZN(new_n3038_));
  NOR2_X1    g02810(.A1(new_n341_), .A2(new_n478_), .ZN(new_n3039_));
  INV_X1     g02811(.I(new_n3039_), .ZN(new_n3040_));
  NAND2_X1   g02812(.A1(new_n3040_), .A2(new_n3038_), .ZN(new_n3041_));
  NAND4_X1   g02813(.A1(new_n2534_), .A2(\a[6] ), .A3(\a[28] ), .A4(new_n392_), .ZN(new_n3042_));
  NOR4_X1    g02814(.A1(new_n3041_), .A2(new_n3034_), .A3(new_n3035_), .A4(new_n3042_), .ZN(new_n3043_));
  NOR2_X1    g02815(.A1(new_n3034_), .A2(new_n3035_), .ZN(new_n3044_));
  NOR2_X1    g02816(.A1(new_n3041_), .A2(new_n3042_), .ZN(new_n3045_));
  NOR2_X1    g02817(.A1(new_n3044_), .A2(new_n3045_), .ZN(new_n3046_));
  OAI21_X1   g02818(.A1(new_n3043_), .A2(new_n3046_), .B(new_n3033_), .ZN(new_n3047_));
  INV_X1     g02819(.I(new_n3033_), .ZN(new_n3048_));
  XOR2_X1    g02820(.A1(new_n3044_), .A2(new_n3045_), .Z(new_n3049_));
  NAND2_X1   g02821(.A1(new_n3049_), .A2(new_n3048_), .ZN(new_n3050_));
  NAND2_X1   g02822(.A1(new_n3050_), .A2(new_n3047_), .ZN(new_n3051_));
  INV_X1     g02823(.I(new_n3051_), .ZN(new_n3052_));
  INV_X1     g02824(.I(new_n2987_), .ZN(new_n3053_));
  AOI21_X1   g02825(.A1(new_n2968_), .A2(new_n3053_), .B(new_n2986_), .ZN(new_n3054_));
  NAND2_X1   g02826(.A1(\a[10] ), .A2(\a[23] ), .ZN(new_n3055_));
  AOI21_X1   g02827(.A1(new_n2974_), .A2(new_n2969_), .B(new_n3055_), .ZN(new_n3056_));
  NOR2_X1    g02828(.A1(new_n3056_), .A2(new_n2975_), .ZN(new_n3057_));
  NOR2_X1    g02829(.A1(new_n786_), .A2(new_n1715_), .ZN(new_n3058_));
  NOR2_X1    g02830(.A1(new_n2979_), .A2(new_n3058_), .ZN(new_n3059_));
  INV_X1     g02831(.I(new_n3059_), .ZN(new_n3060_));
  INV_X1     g02832(.I(new_n651_), .ZN(new_n3061_));
  NAND2_X1   g02833(.A1(new_n3061_), .A2(new_n2286_), .ZN(new_n3062_));
  NAND2_X1   g02834(.A1(\a[2] ), .A2(\a[32] ), .ZN(new_n3063_));
  XNOR2_X1   g02835(.A1(new_n3062_), .A2(new_n3063_), .ZN(new_n3064_));
  NOR2_X1    g02836(.A1(new_n3064_), .A2(new_n3060_), .ZN(new_n3065_));
  INV_X1     g02837(.I(new_n3065_), .ZN(new_n3066_));
  NAND2_X1   g02838(.A1(new_n3064_), .A2(new_n3060_), .ZN(new_n3067_));
  AOI21_X1   g02839(.A1(new_n3066_), .A2(new_n3067_), .B(new_n3057_), .ZN(new_n3068_));
  XOR2_X1    g02840(.A1(new_n3064_), .A2(new_n3060_), .Z(new_n3069_));
  AOI21_X1   g02841(.A1(new_n3069_), .A2(new_n3057_), .B(new_n3068_), .ZN(new_n3070_));
  XOR2_X1    g02842(.A1(new_n3054_), .A2(new_n3070_), .Z(new_n3071_));
  NAND2_X1   g02843(.A1(new_n2995_), .A2(new_n2994_), .ZN(new_n3072_));
  OAI22_X1   g02844(.A1(new_n2891_), .A2(new_n341_), .B1(new_n481_), .B2(new_n2692_), .ZN(new_n3073_));
  NOR2_X1    g02845(.A1(new_n2901_), .A2(new_n2903_), .ZN(new_n3074_));
  OR2_X2     g02846(.A1(new_n2900_), .A2(new_n3074_), .Z(new_n3075_));
  XNOR2_X1   g02847(.A1(new_n3075_), .A2(new_n3073_), .ZN(new_n3076_));
  NOR2_X1    g02848(.A1(new_n3075_), .A2(new_n3073_), .ZN(new_n3077_));
  NAND2_X1   g02849(.A1(new_n3075_), .A2(new_n3073_), .ZN(new_n3078_));
  INV_X1     g02850(.I(new_n3078_), .ZN(new_n3079_));
  OAI21_X1   g02851(.A1(new_n3079_), .A2(new_n3077_), .B(new_n2877_), .ZN(new_n3080_));
  OAI21_X1   g02852(.A1(new_n2877_), .A2(new_n3076_), .B(new_n3080_), .ZN(new_n3081_));
  INV_X1     g02853(.I(new_n2913_), .ZN(new_n3082_));
  AOI21_X1   g02854(.A1(new_n2915_), .A2(new_n2914_), .B(new_n2897_), .ZN(new_n3083_));
  NOR2_X1    g02855(.A1(new_n3083_), .A2(new_n3082_), .ZN(new_n3084_));
  INV_X1     g02856(.I(new_n3084_), .ZN(new_n3085_));
  NAND2_X1   g02857(.A1(new_n268_), .A2(new_n1916_), .ZN(new_n3086_));
  OAI21_X1   g02858(.A1(new_n2908_), .A2(new_n3086_), .B(new_n2909_), .ZN(new_n3087_));
  NAND2_X1   g02859(.A1(\a[1] ), .A2(\a[33] ), .ZN(new_n3088_));
  XNOR2_X1   g02860(.A1(new_n1267_), .A2(new_n3088_), .ZN(new_n3089_));
  NOR2_X1    g02861(.A1(new_n3087_), .A2(new_n3089_), .ZN(new_n3090_));
  XOR2_X1    g02862(.A1(new_n3090_), .A2(new_n2970_), .Z(new_n3091_));
  XOR2_X1    g02863(.A1(new_n3091_), .A2(\a[17] ), .Z(new_n3092_));
  NOR2_X1    g02864(.A1(new_n3092_), .A2(new_n3085_), .ZN(new_n3093_));
  INV_X1     g02865(.I(new_n3092_), .ZN(new_n3094_));
  NOR2_X1    g02866(.A1(new_n3094_), .A2(new_n3084_), .ZN(new_n3095_));
  OR2_X2     g02867(.A1(new_n3095_), .A2(new_n3093_), .Z(new_n3096_));
  XOR2_X1    g02868(.A1(new_n3092_), .A2(new_n3084_), .Z(new_n3097_));
  NOR2_X1    g02869(.A1(new_n3097_), .A2(new_n3081_), .ZN(new_n3098_));
  AOI21_X1   g02870(.A1(new_n3081_), .A2(new_n3096_), .B(new_n3098_), .ZN(new_n3099_));
  INV_X1     g02871(.I(new_n3099_), .ZN(new_n3100_));
  NAND3_X1   g02872(.A1(new_n3072_), .A2(new_n2997_), .A3(new_n3100_), .ZN(new_n3101_));
  AOI21_X1   g02873(.A1(new_n2966_), .A2(new_n2989_), .B(new_n2964_), .ZN(new_n3102_));
  OAI21_X1   g02874(.A1(new_n3102_), .A2(new_n2996_), .B(new_n3099_), .ZN(new_n3103_));
  AOI21_X1   g02875(.A1(new_n3101_), .A2(new_n3103_), .B(new_n3071_), .ZN(new_n3104_));
  INV_X1     g02876(.I(new_n3071_), .ZN(new_n3105_));
  NOR3_X1    g02877(.A1(new_n3102_), .A2(new_n2996_), .A3(new_n3099_), .ZN(new_n3106_));
  INV_X1     g02878(.I(new_n3103_), .ZN(new_n3107_));
  NOR3_X1    g02879(.A1(new_n3107_), .A2(new_n3105_), .A3(new_n3106_), .ZN(new_n3108_));
  OAI21_X1   g02880(.A1(new_n3108_), .A2(new_n3104_), .B(new_n3052_), .ZN(new_n3109_));
  OAI21_X1   g02881(.A1(new_n3107_), .A2(new_n3106_), .B(new_n3105_), .ZN(new_n3110_));
  NAND3_X1   g02882(.A1(new_n3101_), .A2(new_n3071_), .A3(new_n3103_), .ZN(new_n3111_));
  NAND3_X1   g02883(.A1(new_n3110_), .A2(new_n3111_), .A3(new_n3051_), .ZN(new_n3112_));
  AOI21_X1   g02884(.A1(new_n2944_), .A2(new_n2956_), .B(new_n2866_), .ZN(new_n3113_));
  NOR2_X1    g02885(.A1(new_n3113_), .A2(new_n2960_), .ZN(new_n3114_));
  AOI21_X1   g02886(.A1(new_n2941_), .A2(new_n2937_), .B(new_n2938_), .ZN(new_n3115_));
  AOI21_X1   g02887(.A1(new_n2880_), .A2(new_n2885_), .B(new_n2883_), .ZN(new_n3116_));
  AOI21_X1   g02888(.A1(new_n2922_), .A2(new_n2926_), .B(new_n2921_), .ZN(new_n3117_));
  NOR2_X1    g02889(.A1(new_n3117_), .A2(new_n2931_), .ZN(new_n3118_));
  NAND2_X1   g02890(.A1(\a[4] ), .A2(\a[31] ), .ZN(new_n3119_));
  XNOR2_X1   g02891(.A1(new_n2906_), .A2(new_n3119_), .ZN(new_n3120_));
  INV_X1     g02892(.I(new_n3120_), .ZN(new_n3121_));
  NAND2_X1   g02893(.A1(new_n216_), .A2(\a[31] ), .ZN(new_n3122_));
  INV_X1     g02894(.I(new_n257_), .ZN(new_n3123_));
  NAND2_X1   g02895(.A1(new_n3123_), .A2(\a[30] ), .ZN(new_n3124_));
  AOI21_X1   g02896(.A1(new_n3122_), .A2(new_n3124_), .B(\a[34] ), .ZN(new_n3125_));
  NOR2_X1    g02897(.A1(new_n2461_), .A2(new_n2655_), .ZN(new_n3126_));
  INV_X1     g02898(.I(new_n3126_), .ZN(new_n3127_));
  NOR3_X1    g02899(.A1(new_n3125_), .A2(new_n212_), .A3(new_n3127_), .ZN(new_n3128_));
  AOI21_X1   g02900(.A1(new_n3128_), .A2(new_n3121_), .B(\a[34] ), .ZN(new_n3129_));
  NOR2_X1    g02901(.A1(new_n3129_), .A2(new_n199_), .ZN(new_n3130_));
  XNOR2_X1   g02902(.A1(new_n3118_), .A2(new_n3130_), .ZN(new_n3131_));
  NOR4_X1    g02903(.A1(new_n3117_), .A2(new_n2931_), .A3(new_n199_), .A4(new_n3129_), .ZN(new_n3132_));
  NOR2_X1    g02904(.A1(new_n3118_), .A2(new_n3130_), .ZN(new_n3133_));
  OAI21_X1   g02905(.A1(new_n3132_), .A2(new_n3133_), .B(new_n3116_), .ZN(new_n3134_));
  OAI21_X1   g02906(.A1(new_n3116_), .A2(new_n3131_), .B(new_n3134_), .ZN(new_n3135_));
  NOR2_X1    g02907(.A1(new_n2954_), .A2(new_n2952_), .ZN(new_n3136_));
  NOR2_X1    g02908(.A1(new_n3136_), .A2(new_n2953_), .ZN(new_n3137_));
  XOR2_X1    g02909(.A1(new_n3135_), .A2(new_n3137_), .Z(new_n3138_));
  INV_X1     g02910(.I(new_n3138_), .ZN(new_n3139_));
  NOR2_X1    g02911(.A1(new_n3135_), .A2(new_n3137_), .ZN(new_n3140_));
  AND2_X2    g02912(.A1(new_n3135_), .A2(new_n3137_), .Z(new_n3141_));
  OAI21_X1   g02913(.A1(new_n3141_), .A2(new_n3140_), .B(new_n3115_), .ZN(new_n3142_));
  OAI21_X1   g02914(.A1(new_n3139_), .A2(new_n3115_), .B(new_n3142_), .ZN(new_n3143_));
  XOR2_X1    g02915(.A1(new_n3114_), .A2(new_n3143_), .Z(new_n3144_));
  AOI21_X1   g02916(.A1(new_n3109_), .A2(new_n3112_), .B(new_n3144_), .ZN(new_n3145_));
  AOI21_X1   g02917(.A1(new_n3110_), .A2(new_n3111_), .B(new_n3051_), .ZN(new_n3146_));
  NOR3_X1    g02918(.A1(new_n3108_), .A2(new_n3104_), .A3(new_n3052_), .ZN(new_n3147_));
  XNOR2_X1   g02919(.A1(new_n3114_), .A2(new_n3143_), .ZN(new_n3148_));
  NOR3_X1    g02920(.A1(new_n3147_), .A2(new_n3146_), .A3(new_n3148_), .ZN(new_n3149_));
  OAI21_X1   g02921(.A1(new_n3149_), .A2(new_n3145_), .B(new_n3022_), .ZN(new_n3150_));
  INV_X1     g02922(.I(new_n3150_), .ZN(new_n3151_));
  NOR3_X1    g02923(.A1(new_n3149_), .A2(new_n3145_), .A3(new_n3022_), .ZN(new_n3152_));
  NOR2_X1    g02924(.A1(new_n3151_), .A2(new_n3152_), .ZN(new_n3153_));
  XNOR2_X1   g02925(.A1(new_n3021_), .A2(new_n3153_), .ZN(\asquared[35] ));
  NOR2_X1    g02926(.A1(new_n3152_), .A2(new_n3011_), .ZN(new_n3155_));
  AOI21_X1   g02927(.A1(new_n3152_), .A2(new_n3011_), .B(new_n3013_), .ZN(new_n3156_));
  NOR2_X1    g02928(.A1(new_n3156_), .A2(new_n3155_), .ZN(new_n3157_));
  NAND2_X1   g02929(.A1(new_n2865_), .A2(new_n3157_), .ZN(new_n3158_));
  NOR2_X1    g02930(.A1(new_n3114_), .A2(new_n3143_), .ZN(new_n3159_));
  NAND2_X1   g02931(.A1(new_n3114_), .A2(new_n3143_), .ZN(new_n3160_));
  AND3_X2    g02932(.A1(new_n3109_), .A2(new_n3112_), .A3(new_n3160_), .Z(new_n3161_));
  NOR2_X1    g02933(.A1(new_n3102_), .A2(new_n2996_), .ZN(new_n3162_));
  NOR2_X1    g02934(.A1(new_n3162_), .A2(new_n3099_), .ZN(new_n3163_));
  NAND2_X1   g02935(.A1(new_n3162_), .A2(new_n3099_), .ZN(new_n3164_));
  XOR2_X1    g02936(.A1(new_n3071_), .A2(new_n3051_), .Z(new_n3165_));
  AOI21_X1   g02937(.A1(new_n3164_), .A2(new_n3165_), .B(new_n3163_), .ZN(new_n3166_));
  INV_X1     g02938(.I(new_n3166_), .ZN(new_n3167_));
  NOR2_X1    g02939(.A1(new_n3115_), .A2(new_n3141_), .ZN(new_n3168_));
  NOR2_X1    g02940(.A1(new_n3168_), .A2(new_n3140_), .ZN(new_n3169_));
  INV_X1     g02941(.I(new_n3169_), .ZN(new_n3170_));
  INV_X1     g02942(.I(new_n3133_), .ZN(new_n3171_));
  OAI21_X1   g02943(.A1(new_n3116_), .A2(new_n3132_), .B(new_n3171_), .ZN(new_n3172_));
  INV_X1     g02944(.I(new_n3172_), .ZN(new_n3173_));
  INV_X1     g02945(.I(new_n2500_), .ZN(new_n3174_));
  INV_X1     g02946(.I(new_n2898_), .ZN(new_n3175_));
  NOR2_X1    g02947(.A1(new_n3174_), .A2(new_n341_), .ZN(new_n3180_));
  INV_X1     g02948(.I(new_n3180_), .ZN(new_n3181_));
  NAND2_X1   g02949(.A1(new_n2752_), .A2(new_n597_), .ZN(new_n3182_));
  XOR2_X1    g02950(.A1(new_n3182_), .A2(new_n3119_), .Z(new_n3183_));
  NOR2_X1    g02951(.A1(new_n800_), .A2(new_n1339_), .ZN(new_n3184_));
  NAND2_X1   g02952(.A1(new_n3184_), .A2(new_n1441_), .ZN(new_n3185_));
  XOR2_X1    g02953(.A1(new_n3185_), .A2(new_n268_), .Z(new_n3186_));
  NAND2_X1   g02954(.A1(new_n3186_), .A2(new_n2178_), .ZN(new_n3187_));
  XOR2_X1    g02955(.A1(new_n3185_), .A2(\a[7] ), .Z(new_n3188_));
  NAND2_X1   g02956(.A1(new_n3188_), .A2(\a[28] ), .ZN(new_n3189_));
  NAND2_X1   g02957(.A1(new_n3187_), .A2(new_n3189_), .ZN(new_n3190_));
  NAND2_X1   g02958(.A1(new_n3190_), .A2(new_n3183_), .ZN(new_n3191_));
  INV_X1     g02959(.I(new_n3183_), .ZN(new_n3192_));
  INV_X1     g02960(.I(new_n3190_), .ZN(new_n3193_));
  NAND2_X1   g02961(.A1(new_n3193_), .A2(new_n3192_), .ZN(new_n3194_));
  AOI21_X1   g02962(.A1(new_n3194_), .A2(new_n3191_), .B(new_n3181_), .ZN(new_n3195_));
  XOR2_X1    g02963(.A1(new_n3190_), .A2(new_n3192_), .Z(new_n3196_));
  NOR2_X1    g02964(.A1(new_n3196_), .A2(new_n3180_), .ZN(new_n3197_));
  NOR2_X1    g02965(.A1(new_n3197_), .A2(new_n3195_), .ZN(new_n3198_));
  NOR2_X1    g02966(.A1(new_n1267_), .A2(new_n3088_), .ZN(new_n3199_));
  NAND2_X1   g02967(.A1(\a[33] ), .A2(\a[35] ), .ZN(new_n3200_));
  XNOR2_X1   g02968(.A1(new_n197_), .A2(new_n3200_), .ZN(new_n3201_));
  INV_X1     g02969(.I(new_n3201_), .ZN(new_n3202_));
  OAI22_X1   g02970(.A1(new_n786_), .A2(new_n1949_), .B1(new_n873_), .B2(new_n1773_), .ZN(new_n3203_));
  NAND4_X1   g02971(.A1(new_n1018_), .A2(new_n1711_), .A3(\a[13] ), .A4(\a[22] ), .ZN(new_n3204_));
  NOR2_X1    g02972(.A1(new_n3203_), .A2(new_n3204_), .ZN(new_n3205_));
  INV_X1     g02973(.I(new_n3205_), .ZN(new_n3206_));
  NAND2_X1   g02974(.A1(\a[3] ), .A2(\a[32] ), .ZN(new_n3207_));
  INV_X1     g02975(.I(new_n3207_), .ZN(new_n3208_));
  XNOR2_X1   g02976(.A1(new_n651_), .A2(new_n1956_), .ZN(new_n3209_));
  NOR2_X1    g02977(.A1(new_n3206_), .A2(new_n3209_), .ZN(new_n3210_));
  INV_X1     g02978(.I(new_n3209_), .ZN(new_n3211_));
  NOR2_X1    g02979(.A1(new_n3211_), .A2(new_n3205_), .ZN(new_n3212_));
  OAI21_X1   g02980(.A1(new_n3210_), .A2(new_n3212_), .B(new_n3202_), .ZN(new_n3213_));
  XNOR2_X1   g02981(.A1(new_n3205_), .A2(new_n3209_), .ZN(new_n3214_));
  NAND2_X1   g02982(.A1(new_n3214_), .A2(new_n3201_), .ZN(new_n3215_));
  NAND2_X1   g02983(.A1(new_n3215_), .A2(new_n3213_), .ZN(new_n3216_));
  XOR2_X1    g02984(.A1(new_n3198_), .A2(new_n3216_), .Z(new_n3217_));
  NOR2_X1    g02985(.A1(new_n3217_), .A2(new_n3173_), .ZN(new_n3218_));
  OAI21_X1   g02986(.A1(new_n3197_), .A2(new_n3195_), .B(new_n3216_), .ZN(new_n3219_));
  INV_X1     g02987(.I(new_n3216_), .ZN(new_n3220_));
  NAND2_X1   g02988(.A1(new_n3198_), .A2(new_n3220_), .ZN(new_n3221_));
  AOI21_X1   g02989(.A1(new_n3221_), .A2(new_n3219_), .B(new_n3172_), .ZN(new_n3222_));
  NOR2_X1    g02990(.A1(new_n3218_), .A2(new_n3222_), .ZN(new_n3223_));
  NOR2_X1    g02991(.A1(new_n3127_), .A2(new_n212_), .ZN(new_n3224_));
  NOR2_X1    g02992(.A1(new_n3061_), .A2(new_n2286_), .ZN(new_n3225_));
  NAND2_X1   g02993(.A1(new_n201_), .A2(new_n2765_), .ZN(new_n3226_));
  AOI21_X1   g02994(.A1(new_n3061_), .A2(new_n2286_), .B(new_n3226_), .ZN(new_n3227_));
  NOR2_X1    g02995(.A1(new_n3227_), .A2(new_n3225_), .ZN(new_n3228_));
  OAI21_X1   g02996(.A1(new_n1018_), .A2(new_n1715_), .B(new_n3034_), .ZN(new_n3229_));
  XOR2_X1    g02997(.A1(new_n3229_), .A2(new_n3228_), .Z(new_n3230_));
  NOR3_X1    g02998(.A1(new_n3230_), .A2(new_n3224_), .A3(new_n3128_), .ZN(new_n3231_));
  NOR2_X1    g02999(.A1(new_n3128_), .A2(new_n3224_), .ZN(new_n3232_));
  INV_X1     g03000(.I(new_n3228_), .ZN(new_n3233_));
  NOR2_X1    g03001(.A1(new_n3229_), .A2(new_n3233_), .ZN(new_n3234_));
  INV_X1     g03002(.I(new_n3234_), .ZN(new_n3235_));
  NAND2_X1   g03003(.A1(new_n3229_), .A2(new_n3233_), .ZN(new_n3236_));
  AOI21_X1   g03004(.A1(new_n3235_), .A2(new_n3236_), .B(new_n3232_), .ZN(new_n3237_));
  NOR2_X1    g03005(.A1(new_n3231_), .A2(new_n3237_), .ZN(new_n3238_));
  NOR2_X1    g03006(.A1(new_n3048_), .A2(new_n3046_), .ZN(new_n3239_));
  NOR2_X1    g03007(.A1(new_n3239_), .A2(new_n3043_), .ZN(new_n3240_));
  AOI22_X1   g03008(.A1(new_n3040_), .A2(new_n3038_), .B1(new_n609_), .B2(new_n2533_), .ZN(new_n3241_));
  NAND2_X1   g03009(.A1(\a[1] ), .A2(\a[34] ), .ZN(new_n3242_));
  XOR2_X1    g03010(.A1(new_n3242_), .A2(\a[18] ), .Z(new_n3243_));
  INV_X1     g03011(.I(new_n3243_), .ZN(new_n3244_));
  XOR2_X1    g03012(.A1(new_n3241_), .A2(new_n3244_), .Z(new_n3245_));
  NOR2_X1    g03013(.A1(new_n3245_), .A2(new_n3030_), .ZN(new_n3246_));
  INV_X1     g03014(.I(new_n3030_), .ZN(new_n3247_));
  OR2_X2     g03015(.A1(new_n3241_), .A2(new_n3243_), .Z(new_n3248_));
  NAND2_X1   g03016(.A1(new_n3241_), .A2(new_n3243_), .ZN(new_n3249_));
  AOI21_X1   g03017(.A1(new_n3248_), .A2(new_n3249_), .B(new_n3247_), .ZN(new_n3250_));
  NOR2_X1    g03018(.A1(new_n3246_), .A2(new_n3250_), .ZN(new_n3251_));
  INV_X1     g03019(.I(new_n3251_), .ZN(new_n3252_));
  NAND2_X1   g03020(.A1(new_n3252_), .A2(new_n3240_), .ZN(new_n3253_));
  NOR2_X1    g03021(.A1(new_n3252_), .A2(new_n3240_), .ZN(new_n3254_));
  INV_X1     g03022(.I(new_n3254_), .ZN(new_n3255_));
  AOI21_X1   g03023(.A1(new_n3255_), .A2(new_n3253_), .B(new_n3238_), .ZN(new_n3256_));
  INV_X1     g03024(.I(new_n3238_), .ZN(new_n3257_));
  XOR2_X1    g03025(.A1(new_n3240_), .A2(new_n3251_), .Z(new_n3258_));
  NOR2_X1    g03026(.A1(new_n3258_), .A2(new_n3257_), .ZN(new_n3259_));
  NOR2_X1    g03027(.A1(new_n3259_), .A2(new_n3256_), .ZN(new_n3260_));
  NOR2_X1    g03028(.A1(new_n3223_), .A2(new_n3260_), .ZN(new_n3261_));
  INV_X1     g03029(.I(new_n3222_), .ZN(new_n3262_));
  OAI21_X1   g03030(.A1(new_n3173_), .A2(new_n3217_), .B(new_n3262_), .ZN(new_n3263_));
  INV_X1     g03031(.I(new_n3260_), .ZN(new_n3264_));
  NOR2_X1    g03032(.A1(new_n3263_), .A2(new_n3264_), .ZN(new_n3265_));
  OAI21_X1   g03033(.A1(new_n3261_), .A2(new_n3265_), .B(new_n3170_), .ZN(new_n3266_));
  NOR2_X1    g03034(.A1(new_n3263_), .A2(new_n3260_), .ZN(new_n3267_));
  NOR2_X1    g03035(.A1(new_n3223_), .A2(new_n3264_), .ZN(new_n3268_));
  OAI21_X1   g03036(.A1(new_n3268_), .A2(new_n3267_), .B(new_n3169_), .ZN(new_n3269_));
  NOR2_X1    g03037(.A1(new_n3052_), .A2(new_n3070_), .ZN(new_n3270_));
  AOI21_X1   g03038(.A1(new_n3052_), .A2(new_n3070_), .B(new_n3054_), .ZN(new_n3271_));
  NOR2_X1    g03039(.A1(new_n3271_), .A2(new_n3270_), .ZN(new_n3272_));
  AOI21_X1   g03040(.A1(new_n2878_), .A2(new_n3078_), .B(new_n3077_), .ZN(new_n3273_));
  INV_X1     g03041(.I(new_n3273_), .ZN(new_n3274_));
  INV_X1     g03042(.I(new_n2971_), .ZN(new_n3275_));
  AOI21_X1   g03043(.A1(new_n3087_), .A2(new_n3089_), .B(new_n3275_), .ZN(new_n3276_));
  NOR2_X1    g03044(.A1(new_n3276_), .A2(new_n3090_), .ZN(new_n3277_));
  AOI21_X1   g03045(.A1(new_n3060_), .A2(new_n3064_), .B(new_n3057_), .ZN(new_n3278_));
  NOR2_X1    g03046(.A1(new_n3278_), .A2(new_n3065_), .ZN(new_n3279_));
  XOR2_X1    g03047(.A1(new_n3279_), .A2(new_n3277_), .Z(new_n3280_));
  NAND2_X1   g03048(.A1(new_n3280_), .A2(new_n3274_), .ZN(new_n3281_));
  NOR2_X1    g03049(.A1(new_n3279_), .A2(new_n3277_), .ZN(new_n3282_));
  NOR4_X1    g03050(.A1(new_n3278_), .A2(new_n3065_), .A3(new_n3090_), .A4(new_n3276_), .ZN(new_n3283_));
  OAI21_X1   g03051(.A1(new_n3282_), .A2(new_n3283_), .B(new_n3273_), .ZN(new_n3284_));
  NAND2_X1   g03052(.A1(new_n3281_), .A2(new_n3284_), .ZN(new_n3285_));
  INV_X1     g03053(.I(new_n3285_), .ZN(new_n3286_));
  NOR2_X1    g03054(.A1(new_n3093_), .A2(new_n3081_), .ZN(new_n3287_));
  NOR2_X1    g03055(.A1(new_n3287_), .A2(new_n3095_), .ZN(new_n3288_));
  XOR2_X1    g03056(.A1(new_n3288_), .A2(new_n3286_), .Z(new_n3289_));
  NOR2_X1    g03057(.A1(new_n3289_), .A2(new_n3272_), .ZN(new_n3290_));
  NOR2_X1    g03058(.A1(new_n3288_), .A2(new_n3285_), .ZN(new_n3291_));
  NOR3_X1    g03059(.A1(new_n3286_), .A2(new_n3095_), .A3(new_n3287_), .ZN(new_n3292_));
  OR2_X2     g03060(.A1(new_n3292_), .A2(new_n3291_), .Z(new_n3293_));
  AOI21_X1   g03061(.A1(new_n3272_), .A2(new_n3293_), .B(new_n3290_), .ZN(new_n3294_));
  AOI21_X1   g03062(.A1(new_n3269_), .A2(new_n3266_), .B(new_n3294_), .ZN(new_n3295_));
  AND3_X2    g03063(.A1(new_n3266_), .A2(new_n3269_), .A3(new_n3294_), .Z(new_n3296_));
  OAI21_X1   g03064(.A1(new_n3296_), .A2(new_n3295_), .B(new_n3167_), .ZN(new_n3297_));
  NAND2_X1   g03065(.A1(new_n3269_), .A2(new_n3266_), .ZN(new_n3298_));
  NOR2_X1    g03066(.A1(new_n3298_), .A2(new_n3294_), .ZN(new_n3299_));
  NAND2_X1   g03067(.A1(new_n3293_), .A2(new_n3272_), .ZN(new_n3300_));
  OAI21_X1   g03068(.A1(new_n3272_), .A2(new_n3289_), .B(new_n3300_), .ZN(new_n3301_));
  AOI21_X1   g03069(.A1(new_n3269_), .A2(new_n3266_), .B(new_n3301_), .ZN(new_n3302_));
  OAI21_X1   g03070(.A1(new_n3299_), .A2(new_n3302_), .B(new_n3166_), .ZN(new_n3303_));
  NAND2_X1   g03071(.A1(new_n3303_), .A2(new_n3297_), .ZN(new_n3304_));
  OAI21_X1   g03072(.A1(new_n3159_), .A2(new_n3161_), .B(new_n3304_), .ZN(new_n3305_));
  XOR2_X1    g03073(.A1(new_n3158_), .A2(new_n3305_), .Z(new_n3306_));
  XOR2_X1    g03074(.A1(new_n3306_), .A2(new_n3151_), .Z(\asquared[36] ));
  NOR3_X1    g03075(.A1(new_n3304_), .A2(new_n3159_), .A3(new_n3161_), .ZN(new_n3308_));
  NOR2_X1    g03076(.A1(new_n3308_), .A2(new_n3150_), .ZN(new_n3309_));
  NAND3_X1   g03077(.A1(new_n2865_), .A2(new_n3157_), .A3(new_n3309_), .ZN(new_n3310_));
  NAND2_X1   g03078(.A1(new_n3310_), .A2(new_n3305_), .ZN(new_n3311_));
  INV_X1     g03079(.I(new_n3302_), .ZN(new_n3312_));
  OAI21_X1   g03080(.A1(new_n3298_), .A2(new_n3294_), .B(new_n3167_), .ZN(new_n3313_));
  AND2_X2    g03081(.A1(new_n3313_), .A2(new_n3312_), .Z(new_n3314_));
  NOR2_X1    g03082(.A1(new_n3261_), .A2(new_n3169_), .ZN(new_n3315_));
  NOR2_X1    g03083(.A1(new_n3315_), .A2(new_n3265_), .ZN(new_n3316_));
  NAND2_X1   g03084(.A1(new_n3221_), .A2(new_n3172_), .ZN(new_n3317_));
  AOI21_X1   g03085(.A1(new_n3232_), .A2(new_n3236_), .B(new_n3234_), .ZN(new_n3318_));
  NAND2_X1   g03086(.A1(new_n3248_), .A2(new_n3247_), .ZN(new_n3319_));
  NAND2_X1   g03087(.A1(new_n3319_), .A2(new_n3249_), .ZN(new_n3320_));
  INV_X1     g03088(.I(new_n3210_), .ZN(new_n3321_));
  OAI21_X1   g03089(.A1(new_n3205_), .A2(new_n3211_), .B(new_n3202_), .ZN(new_n3322_));
  NAND2_X1   g03090(.A1(new_n3321_), .A2(new_n3322_), .ZN(new_n3323_));
  XNOR2_X1   g03091(.A1(new_n3320_), .A2(new_n3323_), .ZN(new_n3324_));
  NOR2_X1    g03092(.A1(new_n3324_), .A2(new_n3318_), .ZN(new_n3325_));
  INV_X1     g03093(.I(new_n3318_), .ZN(new_n3326_));
  NAND2_X1   g03094(.A1(new_n3320_), .A2(new_n3323_), .ZN(new_n3327_));
  NOR2_X1    g03095(.A1(new_n3320_), .A2(new_n3323_), .ZN(new_n3328_));
  INV_X1     g03096(.I(new_n3328_), .ZN(new_n3329_));
  AOI21_X1   g03097(.A1(new_n3329_), .A2(new_n3327_), .B(new_n3326_), .ZN(new_n3330_));
  NOR2_X1    g03098(.A1(new_n3325_), .A2(new_n3330_), .ZN(new_n3331_));
  AOI21_X1   g03099(.A1(new_n3240_), .A2(new_n3252_), .B(new_n3257_), .ZN(new_n3332_));
  NOR2_X1    g03100(.A1(new_n3332_), .A2(new_n3254_), .ZN(new_n3333_));
  XOR2_X1    g03101(.A1(new_n3333_), .A2(new_n3331_), .Z(new_n3334_));
  AOI21_X1   g03102(.A1(new_n3219_), .A2(new_n3317_), .B(new_n3334_), .ZN(new_n3335_));
  NAND2_X1   g03103(.A1(new_n3317_), .A2(new_n3219_), .ZN(new_n3336_));
  OAI21_X1   g03104(.A1(new_n3254_), .A2(new_n3332_), .B(new_n3331_), .ZN(new_n3337_));
  OAI21_X1   g03105(.A1(new_n3325_), .A2(new_n3330_), .B(new_n3333_), .ZN(new_n3338_));
  AOI21_X1   g03106(.A1(new_n3338_), .A2(new_n3337_), .B(new_n3336_), .ZN(new_n3339_));
  NOR2_X1    g03107(.A1(new_n3335_), .A2(new_n3339_), .ZN(new_n3340_));
  NOR2_X1    g03108(.A1(new_n3272_), .A2(new_n3292_), .ZN(new_n3341_));
  NOR2_X1    g03109(.A1(new_n3341_), .A2(new_n3291_), .ZN(new_n3342_));
  NOR2_X1    g03110(.A1(new_n461_), .A2(new_n2655_), .ZN(new_n3343_));
  NOR4_X1    g03111(.A1(new_n353_), .A2(new_n364_), .A3(new_n2098_), .A4(new_n2655_), .ZN(new_n3344_));
  NAND4_X1   g03112(.A1(new_n3344_), .A2(\a[5] ), .A3(\a[26] ), .A4(new_n3343_), .ZN(new_n3345_));
  AOI21_X1   g03113(.A1(new_n3345_), .A2(new_n2534_), .B(new_n525_), .ZN(new_n3346_));
  NOR3_X1    g03114(.A1(new_n3346_), .A2(new_n461_), .A3(new_n1916_), .ZN(new_n3347_));
  NOR2_X1    g03115(.A1(new_n3346_), .A2(new_n3344_), .ZN(new_n3348_));
  AOI22_X1   g03116(.A1(\a[5] ), .A2(\a[9] ), .B1(\a[27] ), .B2(\a[31] ), .ZN(new_n3349_));
  AOI21_X1   g03117(.A1(new_n3348_), .A2(new_n3349_), .B(new_n3347_), .ZN(new_n3350_));
  NOR2_X1    g03118(.A1(new_n1150_), .A2(new_n1956_), .ZN(new_n3351_));
  NAND2_X1   g03119(.A1(\a[2] ), .A2(\a[34] ), .ZN(new_n3352_));
  XOR2_X1    g03120(.A1(new_n3351_), .A2(new_n3352_), .Z(new_n3353_));
  NOR2_X1    g03121(.A1(new_n2178_), .A2(new_n2461_), .ZN(new_n3354_));
  INV_X1     g03122(.I(new_n3354_), .ZN(new_n3355_));
  NOR2_X1    g03123(.A1(new_n3175_), .A2(new_n3355_), .ZN(new_n3356_));
  NOR2_X1    g03124(.A1(new_n3356_), .A2(new_n3039_), .ZN(new_n3357_));
  NOR2_X1    g03125(.A1(new_n242_), .A2(new_n2461_), .ZN(new_n3358_));
  NAND4_X1   g03126(.A1(new_n3357_), .A2(new_n392_), .A3(new_n2689_), .A4(new_n3358_), .ZN(new_n3359_));
  NOR2_X1    g03127(.A1(new_n3359_), .A2(new_n3353_), .ZN(new_n3360_));
  NAND2_X1   g03128(.A1(new_n3359_), .A2(new_n3353_), .ZN(new_n3361_));
  INV_X1     g03129(.I(new_n3361_), .ZN(new_n3362_));
  NOR2_X1    g03130(.A1(new_n3362_), .A2(new_n3360_), .ZN(new_n3363_));
  INV_X1     g03131(.I(new_n3363_), .ZN(new_n3364_));
  XNOR2_X1   g03132(.A1(new_n3359_), .A2(new_n3353_), .ZN(new_n3365_));
  NOR2_X1    g03133(.A1(new_n3365_), .A2(new_n3350_), .ZN(new_n3366_));
  AOI21_X1   g03134(.A1(new_n3350_), .A2(new_n3364_), .B(new_n3366_), .ZN(new_n3367_));
  INV_X1     g03135(.I(new_n3367_), .ZN(new_n3368_));
  NOR2_X1    g03136(.A1(new_n3283_), .A2(new_n3273_), .ZN(new_n3369_));
  NOR2_X1    g03137(.A1(new_n3369_), .A2(new_n3282_), .ZN(new_n3370_));
  INV_X1     g03138(.I(\a[34] ), .ZN(new_n3371_));
  NOR2_X1    g03139(.A1(new_n1119_), .A2(new_n3371_), .ZN(new_n3372_));
  NAND2_X1   g03140(.A1(\a[17] ), .A2(\a[19] ), .ZN(new_n3373_));
  NAND2_X1   g03141(.A1(\a[1] ), .A2(\a[35] ), .ZN(new_n3374_));
  NAND2_X1   g03142(.A1(new_n3373_), .A2(new_n3374_), .ZN(new_n3375_));
  INV_X1     g03143(.I(new_n3375_), .ZN(new_n3376_));
  NOR2_X1    g03144(.A1(new_n3373_), .A2(new_n3374_), .ZN(new_n3377_));
  OAI21_X1   g03145(.A1(new_n3376_), .A2(new_n3377_), .B(new_n3372_), .ZN(new_n3378_));
  XOR2_X1    g03146(.A1(new_n3378_), .A2(\a[0] ), .Z(new_n3379_));
  XOR2_X1    g03147(.A1(new_n3379_), .A2(\a[36] ), .Z(new_n3380_));
  NAND4_X1   g03148(.A1(\a[3] ), .A2(\a[4] ), .A3(\a[32] ), .A4(\a[33] ), .ZN(new_n3382_));
  INV_X1     g03149(.I(new_n1019_), .ZN(new_n3383_));
  OAI21_X1   g03150(.A1(new_n1773_), .A2(new_n1949_), .B(new_n3383_), .ZN(new_n3384_));
  NAND4_X1   g03151(.A1(new_n1021_), .A2(new_n1711_), .A3(\a[14] ), .A4(\a[22] ), .ZN(new_n3385_));
  NOR2_X1    g03152(.A1(new_n3384_), .A2(new_n3385_), .ZN(new_n3386_));
  INV_X1     g03153(.I(new_n3386_), .ZN(new_n3387_));
  NOR2_X1    g03154(.A1(new_n3387_), .A2(new_n3382_), .ZN(new_n3388_));
  INV_X1     g03155(.I(new_n3382_), .ZN(new_n3389_));
  NOR2_X1    g03156(.A1(new_n3386_), .A2(new_n3389_), .ZN(new_n3390_));
  NOR2_X1    g03157(.A1(new_n3388_), .A2(new_n3390_), .ZN(new_n3391_));
  NOR2_X1    g03158(.A1(new_n3380_), .A2(new_n3391_), .ZN(new_n3392_));
  INV_X1     g03159(.I(\a[36] ), .ZN(new_n3393_));
  XOR2_X1    g03160(.A1(new_n3379_), .A2(new_n3393_), .Z(new_n3394_));
  NAND2_X1   g03161(.A1(new_n3386_), .A2(new_n3382_), .ZN(new_n3395_));
  NAND2_X1   g03162(.A1(new_n3387_), .A2(new_n3389_), .ZN(new_n3396_));
  AOI21_X1   g03163(.A1(new_n3395_), .A2(new_n3396_), .B(new_n3394_), .ZN(new_n3397_));
  NOR2_X1    g03164(.A1(new_n3397_), .A2(new_n3392_), .ZN(new_n3398_));
  NOR2_X1    g03165(.A1(new_n3398_), .A2(new_n3370_), .ZN(new_n3399_));
  NOR4_X1    g03166(.A1(new_n3397_), .A2(new_n3282_), .A3(new_n3369_), .A4(new_n3392_), .ZN(new_n3400_));
  OAI21_X1   g03167(.A1(new_n3399_), .A2(new_n3400_), .B(new_n3368_), .ZN(new_n3401_));
  XNOR2_X1   g03168(.A1(new_n3398_), .A2(new_n3370_), .ZN(new_n3402_));
  OAI21_X1   g03169(.A1(new_n3402_), .A2(new_n3368_), .B(new_n3401_), .ZN(new_n3403_));
  OAI22_X1   g03170(.A1(new_n341_), .A2(new_n3174_), .B1(new_n3175_), .B2(new_n481_), .ZN(new_n3404_));
  NAND2_X1   g03171(.A1(new_n2752_), .A2(new_n597_), .ZN(new_n3405_));
  NOR2_X1    g03172(.A1(new_n2752_), .A2(new_n597_), .ZN(new_n3406_));
  NOR2_X1    g03173(.A1(\a[4] ), .A2(\a[31] ), .ZN(new_n3407_));
  AOI21_X1   g03174(.A1(new_n3405_), .A2(new_n3407_), .B(new_n3406_), .ZN(new_n3408_));
  NOR2_X1    g03175(.A1(new_n3184_), .A2(new_n1441_), .ZN(new_n3409_));
  NAND2_X1   g03176(.A1(\a[7] ), .A2(\a[28] ), .ZN(new_n3410_));
  OAI21_X1   g03177(.A1(new_n3409_), .A2(new_n3410_), .B(new_n3185_), .ZN(new_n3411_));
  XNOR2_X1   g03178(.A1(new_n3408_), .A2(new_n3411_), .ZN(new_n3412_));
  NOR2_X1    g03179(.A1(new_n3412_), .A2(new_n3404_), .ZN(new_n3413_));
  INV_X1     g03180(.I(new_n3404_), .ZN(new_n3414_));
  NAND2_X1   g03181(.A1(new_n3408_), .A2(new_n3411_), .ZN(new_n3415_));
  OR2_X2     g03182(.A1(new_n3408_), .A2(new_n3411_), .Z(new_n3416_));
  AOI21_X1   g03183(.A1(new_n3416_), .A2(new_n3415_), .B(new_n3414_), .ZN(new_n3417_));
  NOR2_X1    g03184(.A1(new_n3413_), .A2(new_n3417_), .ZN(new_n3418_));
  INV_X1     g03185(.I(new_n3418_), .ZN(new_n3419_));
  INV_X1     g03186(.I(new_n3191_), .ZN(new_n3420_));
  AOI21_X1   g03187(.A1(new_n3193_), .A2(new_n3192_), .B(new_n3181_), .ZN(new_n3421_));
  NOR2_X1    g03188(.A1(new_n3421_), .A2(new_n3420_), .ZN(new_n3422_));
  INV_X1     g03189(.I(\a[35] ), .ZN(new_n3423_));
  NOR2_X1    g03190(.A1(new_n2868_), .A2(new_n3423_), .ZN(new_n3424_));
  AOI21_X1   g03191(.A1(new_n3199_), .A2(new_n218_), .B(new_n3424_), .ZN(new_n3425_));
  OAI21_X1   g03192(.A1(new_n1018_), .A2(new_n1711_), .B(new_n3203_), .ZN(new_n3426_));
  OAI21_X1   g03193(.A1(new_n651_), .A2(new_n3207_), .B(new_n1956_), .ZN(new_n3427_));
  XOR2_X1    g03194(.A1(new_n3426_), .A2(new_n3427_), .Z(new_n3428_));
  INV_X1     g03195(.I(new_n3427_), .ZN(new_n3429_));
  NOR2_X1    g03196(.A1(new_n3426_), .A2(new_n3429_), .ZN(new_n3430_));
  AND2_X2    g03197(.A1(new_n3426_), .A2(new_n3429_), .Z(new_n3431_));
  OAI21_X1   g03198(.A1(new_n3431_), .A2(new_n3430_), .B(new_n3425_), .ZN(new_n3432_));
  OAI21_X1   g03199(.A1(new_n3425_), .A2(new_n3428_), .B(new_n3432_), .ZN(new_n3433_));
  NAND2_X1   g03200(.A1(new_n3422_), .A2(new_n3433_), .ZN(new_n3434_));
  INV_X1     g03201(.I(new_n3433_), .ZN(new_n3435_));
  OAI21_X1   g03202(.A1(new_n3421_), .A2(new_n3420_), .B(new_n3435_), .ZN(new_n3436_));
  NAND2_X1   g03203(.A1(new_n3434_), .A2(new_n3436_), .ZN(new_n3437_));
  XOR2_X1    g03204(.A1(new_n3422_), .A2(new_n3435_), .Z(new_n3438_));
  NOR2_X1    g03205(.A1(new_n3438_), .A2(new_n3419_), .ZN(new_n3439_));
  AOI21_X1   g03206(.A1(new_n3419_), .A2(new_n3437_), .B(new_n3439_), .ZN(new_n3440_));
  XNOR2_X1   g03207(.A1(new_n3440_), .A2(new_n3403_), .ZN(new_n3441_));
  NOR2_X1    g03208(.A1(new_n3441_), .A2(new_n3342_), .ZN(new_n3442_));
  OR2_X2     g03209(.A1(new_n3440_), .A2(new_n3403_), .Z(new_n3443_));
  NAND2_X1   g03210(.A1(new_n3440_), .A2(new_n3403_), .ZN(new_n3444_));
  NAND2_X1   g03211(.A1(new_n3443_), .A2(new_n3444_), .ZN(new_n3445_));
  NAND2_X1   g03212(.A1(new_n3445_), .A2(new_n3342_), .ZN(new_n3446_));
  INV_X1     g03213(.I(new_n3446_), .ZN(new_n3447_));
  OAI21_X1   g03214(.A1(new_n3447_), .A2(new_n3442_), .B(new_n3340_), .ZN(new_n3448_));
  INV_X1     g03215(.I(new_n3340_), .ZN(new_n3449_));
  INV_X1     g03216(.I(new_n3442_), .ZN(new_n3450_));
  NAND3_X1   g03217(.A1(new_n3450_), .A2(new_n3446_), .A3(new_n3449_), .ZN(new_n3451_));
  AOI21_X1   g03218(.A1(new_n3448_), .A2(new_n3451_), .B(new_n3316_), .ZN(new_n3452_));
  INV_X1     g03219(.I(new_n3316_), .ZN(new_n3453_));
  OAI21_X1   g03220(.A1(new_n3447_), .A2(new_n3442_), .B(new_n3449_), .ZN(new_n3454_));
  NAND3_X1   g03221(.A1(new_n3450_), .A2(new_n3446_), .A3(new_n3340_), .ZN(new_n3455_));
  AOI21_X1   g03222(.A1(new_n3454_), .A2(new_n3455_), .B(new_n3453_), .ZN(new_n3456_));
  NOR2_X1    g03223(.A1(new_n3452_), .A2(new_n3456_), .ZN(new_n3457_));
  XNOR2_X1   g03224(.A1(new_n3314_), .A2(new_n3457_), .ZN(new_n3458_));
  NAND2_X1   g03225(.A1(new_n3311_), .A2(new_n3458_), .ZN(new_n3459_));
  OAI21_X1   g03226(.A1(new_n3452_), .A2(new_n3456_), .B(new_n3314_), .ZN(new_n3460_));
  INV_X1     g03227(.I(new_n3314_), .ZN(new_n3461_));
  NAND2_X1   g03228(.A1(new_n3461_), .A2(new_n3457_), .ZN(new_n3462_));
  AND2_X2    g03229(.A1(new_n3462_), .A2(new_n3460_), .Z(new_n3463_));
  OAI21_X1   g03230(.A1(new_n3311_), .A2(new_n3463_), .B(new_n3459_), .ZN(\asquared[37] ));
  NAND2_X1   g03231(.A1(new_n3311_), .A2(new_n3460_), .ZN(new_n3465_));
  NAND2_X1   g03232(.A1(new_n3465_), .A2(new_n3462_), .ZN(new_n3466_));
  NAND2_X1   g03233(.A1(new_n3454_), .A2(new_n3453_), .ZN(new_n3467_));
  NAND2_X1   g03234(.A1(new_n3338_), .A2(new_n3336_), .ZN(new_n3468_));
  NAND2_X1   g03235(.A1(new_n3468_), .A2(new_n3337_), .ZN(new_n3469_));
  OAI21_X1   g03236(.A1(new_n3318_), .A2(new_n3328_), .B(new_n3327_), .ZN(new_n3470_));
  INV_X1     g03237(.I(new_n3470_), .ZN(new_n3471_));
  OAI22_X1   g03238(.A1(new_n1999_), .A2(new_n527_), .B1(new_n257_), .B2(new_n2868_), .ZN(new_n3472_));
  INV_X1     g03239(.I(new_n788_), .ZN(new_n3473_));
  NOR2_X1    g03240(.A1(new_n1999_), .A2(new_n2868_), .ZN(new_n3474_));
  NAND2_X1   g03241(.A1(new_n3474_), .A2(new_n3473_), .ZN(new_n3475_));
  NAND3_X1   g03242(.A1(new_n3475_), .A2(new_n3472_), .A3(\a[37] ), .ZN(new_n3476_));
  NAND3_X1   g03243(.A1(new_n3476_), .A2(\a[0] ), .A3(\a[37] ), .ZN(new_n3477_));
  AOI22_X1   g03244(.A1(new_n3472_), .A2(\a[37] ), .B1(new_n3473_), .B2(new_n3474_), .ZN(new_n3478_));
  NOR2_X1    g03245(.A1(new_n3474_), .A2(new_n3473_), .ZN(new_n3479_));
  NAND2_X1   g03246(.A1(new_n3478_), .A2(new_n3479_), .ZN(new_n3480_));
  NAND2_X1   g03247(.A1(new_n3477_), .A2(new_n3480_), .ZN(new_n3481_));
  NOR2_X1    g03248(.A1(new_n364_), .A2(new_n2178_), .ZN(new_n3482_));
  NOR2_X1    g03249(.A1(new_n3127_), .A2(new_n478_), .ZN(new_n3483_));
  NAND4_X1   g03250(.A1(new_n3483_), .A2(\a[6] ), .A3(new_n3482_), .A4(\a[31] ), .ZN(new_n3484_));
  AOI21_X1   g03251(.A1(new_n3484_), .A2(new_n3355_), .B(new_n772_), .ZN(new_n3485_));
  NOR2_X1    g03252(.A1(new_n3127_), .A2(new_n478_), .ZN(new_n3486_));
  NOR2_X1    g03253(.A1(new_n3371_), .A2(new_n3423_), .ZN(new_n3487_));
  NAND2_X1   g03254(.A1(new_n3487_), .A2(new_n232_), .ZN(new_n3488_));
  NAND2_X1   g03255(.A1(\a[16] ), .A2(\a[21] ), .ZN(new_n3489_));
  XOR2_X1    g03256(.A1(new_n3488_), .A2(new_n3489_), .Z(new_n3490_));
  NAND2_X1   g03257(.A1(new_n3490_), .A2(new_n3486_), .ZN(new_n3491_));
  NOR2_X1    g03258(.A1(new_n3490_), .A2(new_n3486_), .ZN(new_n3492_));
  INV_X1     g03259(.I(new_n3492_), .ZN(new_n3493_));
  AOI21_X1   g03260(.A1(new_n3493_), .A2(new_n3491_), .B(new_n3481_), .ZN(new_n3494_));
  XNOR2_X1   g03261(.A1(new_n3490_), .A2(new_n3486_), .ZN(new_n3495_));
  AOI21_X1   g03262(.A1(new_n3477_), .A2(new_n3480_), .B(new_n3495_), .ZN(new_n3496_));
  NOR2_X1    g03263(.A1(new_n3496_), .A2(new_n3494_), .ZN(new_n3497_));
  NOR2_X1    g03264(.A1(new_n3431_), .A2(new_n3425_), .ZN(new_n3498_));
  NOR2_X1    g03265(.A1(new_n3498_), .A2(new_n3430_), .ZN(new_n3499_));
  NAND2_X1   g03266(.A1(\a[26] ), .A2(\a[32] ), .ZN(new_n3500_));
  OAI22_X1   g03267(.A1(new_n2534_), .A2(new_n3500_), .B1(new_n509_), .B2(new_n796_), .ZN(new_n3501_));
  NAND4_X1   g03268(.A1(\a[5] ), .A2(\a[10] ), .A3(\a[27] ), .A4(\a[32] ), .ZN(new_n3502_));
  NOR2_X1    g03269(.A1(new_n675_), .A2(new_n1916_), .ZN(new_n3503_));
  NAND2_X1   g03270(.A1(\a[27] ), .A2(\a[32] ), .ZN(new_n3504_));
  NAND4_X1   g03271(.A1(new_n3503_), .A2(new_n3502_), .A3(new_n3025_), .A4(new_n3504_), .ZN(new_n3505_));
  NOR2_X1    g03272(.A1(new_n3501_), .A2(new_n3505_), .ZN(new_n3506_));
  INV_X1     g03273(.I(new_n3506_), .ZN(new_n3507_));
  AOI21_X1   g03274(.A1(\a[17] ), .A2(\a[20] ), .B(new_n2331_), .ZN(new_n3508_));
  NAND3_X1   g03275(.A1(new_n3508_), .A2(new_n1441_), .A3(new_n1798_), .ZN(new_n3509_));
  NAND2_X1   g03276(.A1(\a[8] ), .A2(\a[29] ), .ZN(new_n3510_));
  XOR2_X1    g03277(.A1(new_n3509_), .A2(new_n3510_), .Z(new_n3511_));
  XOR2_X1    g03278(.A1(new_n3511_), .A2(new_n3507_), .Z(new_n3512_));
  NOR2_X1    g03279(.A1(new_n3512_), .A2(new_n3499_), .ZN(new_n3513_));
  INV_X1     g03280(.I(new_n3499_), .ZN(new_n3514_));
  NAND2_X1   g03281(.A1(new_n3511_), .A2(new_n3506_), .ZN(new_n3515_));
  NOR2_X1    g03282(.A1(new_n3511_), .A2(new_n3506_), .ZN(new_n3516_));
  INV_X1     g03283(.I(new_n3516_), .ZN(new_n3517_));
  AOI21_X1   g03284(.A1(new_n3515_), .A2(new_n3517_), .B(new_n3514_), .ZN(new_n3518_));
  NOR2_X1    g03285(.A1(new_n3513_), .A2(new_n3518_), .ZN(new_n3519_));
  XOR2_X1    g03286(.A1(new_n3519_), .A2(new_n3497_), .Z(new_n3520_));
  NOR2_X1    g03287(.A1(new_n3520_), .A2(new_n3471_), .ZN(new_n3521_));
  OAI21_X1   g03288(.A1(new_n3513_), .A2(new_n3518_), .B(new_n3497_), .ZN(new_n3522_));
  OAI21_X1   g03289(.A1(new_n3494_), .A2(new_n3496_), .B(new_n3519_), .ZN(new_n3523_));
  AOI21_X1   g03290(.A1(new_n3523_), .A2(new_n3522_), .B(new_n3470_), .ZN(new_n3524_));
  NOR2_X1    g03291(.A1(new_n3521_), .A2(new_n3524_), .ZN(new_n3525_));
  INV_X1     g03292(.I(new_n3348_), .ZN(new_n3526_));
  INV_X1     g03293(.I(new_n3378_), .ZN(new_n3527_));
  NOR3_X1    g03294(.A1(new_n3376_), .A2(new_n3372_), .A3(new_n3377_), .ZN(new_n3528_));
  NOR3_X1    g03295(.A1(new_n3528_), .A2(new_n199_), .A3(new_n3393_), .ZN(new_n3529_));
  NOR2_X1    g03296(.A1(new_n3529_), .A2(new_n3527_), .ZN(new_n3530_));
  AOI22_X1   g03297(.A1(new_n787_), .A2(new_n2383_), .B1(new_n2328_), .B2(new_n2543_), .ZN(new_n3531_));
  NOR2_X1    g03298(.A1(new_n599_), .A2(new_n1691_), .ZN(new_n3532_));
  NAND4_X1   g03299(.A1(new_n3531_), .A2(new_n1018_), .A3(new_n2285_), .A4(new_n3532_), .ZN(new_n3533_));
  NOR2_X1    g03300(.A1(new_n3530_), .A2(new_n3533_), .ZN(new_n3534_));
  INV_X1     g03301(.I(new_n3534_), .ZN(new_n3535_));
  NAND2_X1   g03302(.A1(new_n3530_), .A2(new_n3533_), .ZN(new_n3536_));
  AOI21_X1   g03303(.A1(new_n3535_), .A2(new_n3536_), .B(new_n3526_), .ZN(new_n3537_));
  XNOR2_X1   g03304(.A1(new_n3530_), .A2(new_n3533_), .ZN(new_n3538_));
  NOR2_X1    g03305(.A1(new_n3538_), .A2(new_n3348_), .ZN(new_n3539_));
  NOR2_X1    g03306(.A1(new_n3539_), .A2(new_n3537_), .ZN(new_n3540_));
  NAND2_X1   g03307(.A1(new_n1220_), .A2(new_n2543_), .ZN(new_n3541_));
  NOR2_X1    g03308(.A1(new_n1220_), .A2(new_n2543_), .ZN(new_n3542_));
  NOR2_X1    g03309(.A1(\a[2] ), .A2(\a[34] ), .ZN(new_n3543_));
  AOI21_X1   g03310(.A1(new_n3541_), .A2(new_n3543_), .B(new_n3542_), .ZN(new_n3544_));
  INV_X1     g03311(.I(new_n3544_), .ZN(new_n3545_));
  NAND4_X1   g03312(.A1(\a[3] ), .A2(\a[4] ), .A3(\a[32] ), .A4(\a[33] ), .ZN(new_n3546_));
  INV_X1     g03313(.I(new_n3546_), .ZN(new_n3547_));
  NAND2_X1   g03314(.A1(new_n1719_), .A2(new_n2978_), .ZN(new_n3548_));
  NAND2_X1   g03315(.A1(new_n3384_), .A2(new_n3548_), .ZN(new_n3549_));
  XOR2_X1    g03316(.A1(new_n3549_), .A2(new_n3547_), .Z(new_n3550_));
  NOR2_X1    g03317(.A1(new_n3549_), .A2(new_n3546_), .ZN(new_n3551_));
  INV_X1     g03318(.I(new_n3549_), .ZN(new_n3552_));
  NOR2_X1    g03319(.A1(new_n3552_), .A2(new_n3547_), .ZN(new_n3553_));
  OAI21_X1   g03320(.A1(new_n3553_), .A2(new_n3551_), .B(new_n3545_), .ZN(new_n3554_));
  OAI21_X1   g03321(.A1(new_n3550_), .A2(new_n3545_), .B(new_n3554_), .ZN(new_n3555_));
  INV_X1     g03322(.I(new_n3390_), .ZN(new_n3556_));
  AOI21_X1   g03323(.A1(new_n3394_), .A2(new_n3556_), .B(new_n3388_), .ZN(new_n3557_));
  NOR2_X1    g03324(.A1(new_n3557_), .A2(new_n3555_), .ZN(new_n3558_));
  INV_X1     g03325(.I(new_n3558_), .ZN(new_n3559_));
  NAND2_X1   g03326(.A1(new_n3557_), .A2(new_n3555_), .ZN(new_n3560_));
  AOI21_X1   g03327(.A1(new_n3559_), .A2(new_n3560_), .B(new_n3540_), .ZN(new_n3561_));
  XNOR2_X1   g03328(.A1(new_n3557_), .A2(new_n3555_), .ZN(new_n3562_));
  NOR3_X1    g03329(.A1(new_n3562_), .A2(new_n3537_), .A3(new_n3539_), .ZN(new_n3563_));
  NOR2_X1    g03330(.A1(new_n3563_), .A2(new_n3561_), .ZN(new_n3564_));
  XNOR2_X1   g03331(.A1(new_n3525_), .A2(new_n3564_), .ZN(new_n3565_));
  NAND2_X1   g03332(.A1(new_n3565_), .A2(new_n3469_), .ZN(new_n3566_));
  INV_X1     g03333(.I(new_n3469_), .ZN(new_n3567_));
  NOR3_X1    g03334(.A1(new_n3564_), .A2(new_n3521_), .A3(new_n3524_), .ZN(new_n3568_));
  NOR3_X1    g03335(.A1(new_n3525_), .A2(new_n3561_), .A3(new_n3563_), .ZN(new_n3569_));
  OAI21_X1   g03336(.A1(new_n3569_), .A2(new_n3568_), .B(new_n3567_), .ZN(new_n3570_));
  NAND2_X1   g03337(.A1(new_n3566_), .A2(new_n3570_), .ZN(new_n3571_));
  OAI21_X1   g03338(.A1(new_n3291_), .A2(new_n3341_), .B(new_n3443_), .ZN(new_n3572_));
  NAND2_X1   g03339(.A1(new_n3572_), .A2(new_n3444_), .ZN(new_n3573_));
  NOR2_X1    g03340(.A1(new_n3400_), .A2(new_n3367_), .ZN(new_n3574_));
  NOR2_X1    g03341(.A1(new_n3574_), .A2(new_n3399_), .ZN(new_n3575_));
  AOI21_X1   g03342(.A1(new_n3350_), .A2(new_n3361_), .B(new_n3360_), .ZN(new_n3576_));
  NAND2_X1   g03343(.A1(new_n3416_), .A2(new_n3414_), .ZN(new_n3577_));
  NAND2_X1   g03344(.A1(new_n3577_), .A2(new_n3415_), .ZN(new_n3578_));
  OAI22_X1   g03345(.A1(new_n3356_), .A2(new_n3039_), .B1(new_n392_), .B2(new_n2689_), .ZN(new_n3579_));
  INV_X1     g03346(.I(new_n3579_), .ZN(new_n3580_));
  INV_X1     g03347(.I(new_n3377_), .ZN(new_n3581_));
  NAND2_X1   g03348(.A1(\a[1] ), .A2(\a[36] ), .ZN(new_n3582_));
  XOR2_X1    g03349(.A1(new_n3582_), .A2(\a[19] ), .Z(new_n3583_));
  XOR2_X1    g03350(.A1(new_n3583_), .A2(new_n3581_), .Z(new_n3584_));
  NAND2_X1   g03351(.A1(new_n3584_), .A2(new_n3580_), .ZN(new_n3585_));
  NOR2_X1    g03352(.A1(new_n3583_), .A2(new_n3581_), .ZN(new_n3586_));
  NAND2_X1   g03353(.A1(new_n3583_), .A2(new_n3581_), .ZN(new_n3587_));
  INV_X1     g03354(.I(new_n3587_), .ZN(new_n3588_));
  OAI21_X1   g03355(.A1(new_n3588_), .A2(new_n3586_), .B(new_n3579_), .ZN(new_n3589_));
  NAND2_X1   g03356(.A1(new_n3585_), .A2(new_n3589_), .ZN(new_n3590_));
  XOR2_X1    g03357(.A1(new_n3578_), .A2(new_n3590_), .Z(new_n3591_));
  AOI21_X1   g03358(.A1(new_n3585_), .A2(new_n3589_), .B(new_n3578_), .ZN(new_n3592_));
  AOI21_X1   g03359(.A1(new_n3415_), .A2(new_n3577_), .B(new_n3590_), .ZN(new_n3593_));
  OAI21_X1   g03360(.A1(new_n3592_), .A2(new_n3593_), .B(new_n3576_), .ZN(new_n3594_));
  OAI21_X1   g03361(.A1(new_n3576_), .A2(new_n3591_), .B(new_n3594_), .ZN(new_n3595_));
  NAND2_X1   g03362(.A1(new_n3434_), .A2(new_n3418_), .ZN(new_n3596_));
  NAND2_X1   g03363(.A1(new_n3596_), .A2(new_n3436_), .ZN(new_n3597_));
  XOR2_X1    g03364(.A1(new_n3597_), .A2(new_n3595_), .Z(new_n3598_));
  NOR2_X1    g03365(.A1(new_n3598_), .A2(new_n3575_), .ZN(new_n3599_));
  INV_X1     g03366(.I(new_n3595_), .ZN(new_n3600_));
  NAND2_X1   g03367(.A1(new_n3597_), .A2(new_n3600_), .ZN(new_n3601_));
  NAND3_X1   g03368(.A1(new_n3596_), .A2(new_n3595_), .A3(new_n3436_), .ZN(new_n3602_));
  NAND2_X1   g03369(.A1(new_n3601_), .A2(new_n3602_), .ZN(new_n3603_));
  AOI21_X1   g03370(.A1(new_n3575_), .A2(new_n3603_), .B(new_n3599_), .ZN(new_n3604_));
  NOR2_X1    g03371(.A1(new_n3573_), .A2(new_n3604_), .ZN(new_n3605_));
  NAND2_X1   g03372(.A1(new_n3573_), .A2(new_n3604_), .ZN(new_n3606_));
  INV_X1     g03373(.I(new_n3606_), .ZN(new_n3607_));
  OAI21_X1   g03374(.A1(new_n3607_), .A2(new_n3605_), .B(new_n3571_), .ZN(new_n3608_));
  INV_X1     g03375(.I(new_n3571_), .ZN(new_n3609_));
  AOI21_X1   g03376(.A1(new_n3572_), .A2(new_n3444_), .B(new_n3604_), .ZN(new_n3610_));
  INV_X1     g03377(.I(new_n3604_), .ZN(new_n3611_));
  NOR2_X1    g03378(.A1(new_n3573_), .A2(new_n3611_), .ZN(new_n3612_));
  OAI21_X1   g03379(.A1(new_n3612_), .A2(new_n3610_), .B(new_n3609_), .ZN(new_n3613_));
  NAND2_X1   g03380(.A1(new_n3613_), .A2(new_n3608_), .ZN(new_n3614_));
  NAND3_X1   g03381(.A1(new_n3614_), .A2(new_n3455_), .A3(new_n3467_), .ZN(new_n3615_));
  NAND2_X1   g03382(.A1(new_n3467_), .A2(new_n3455_), .ZN(new_n3616_));
  NAND3_X1   g03383(.A1(new_n3616_), .A2(new_n3613_), .A3(new_n3608_), .ZN(new_n3617_));
  NAND2_X1   g03384(.A1(new_n3615_), .A2(new_n3617_), .ZN(new_n3618_));
  XOR2_X1    g03385(.A1(new_n3466_), .A2(new_n3618_), .Z(\asquared[38] ));
  NAND2_X1   g03386(.A1(new_n3617_), .A2(new_n3457_), .ZN(new_n3620_));
  OAI21_X1   g03387(.A1(new_n3617_), .A2(new_n3457_), .B(new_n3314_), .ZN(new_n3621_));
  NAND2_X1   g03388(.A1(new_n3621_), .A2(new_n3620_), .ZN(new_n3622_));
  AOI21_X1   g03389(.A1(new_n3310_), .A2(new_n3305_), .B(new_n3622_), .ZN(new_n3623_));
  OAI21_X1   g03390(.A1(new_n3571_), .A2(new_n3605_), .B(new_n3606_), .ZN(new_n3624_));
  INV_X1     g03391(.I(new_n3624_), .ZN(new_n3625_));
  NOR2_X1    g03392(.A1(new_n3567_), .A2(new_n3569_), .ZN(new_n3626_));
  NOR2_X1    g03393(.A1(new_n3626_), .A2(new_n3568_), .ZN(new_n3627_));
  INV_X1     g03394(.I(new_n3602_), .ZN(new_n3628_));
  OAI21_X1   g03395(.A1(new_n3575_), .A2(new_n3628_), .B(new_n3601_), .ZN(new_n3629_));
  NOR2_X1    g03396(.A1(new_n3592_), .A2(new_n3576_), .ZN(new_n3630_));
  OAI21_X1   g03397(.A1(new_n3579_), .A2(new_n3586_), .B(new_n3587_), .ZN(new_n3631_));
  INV_X1     g03398(.I(new_n3631_), .ZN(new_n3632_));
  INV_X1     g03399(.I(new_n3551_), .ZN(new_n3633_));
  OAI21_X1   g03400(.A1(new_n3552_), .A2(new_n3547_), .B(new_n3544_), .ZN(new_n3634_));
  NAND2_X1   g03401(.A1(new_n3634_), .A2(new_n3633_), .ZN(new_n3635_));
  NAND2_X1   g03402(.A1(\a[12] ), .A2(\a[34] ), .ZN(new_n3636_));
  OAI22_X1   g03403(.A1(new_n2534_), .A2(new_n2537_), .B1(new_n651_), .B2(new_n3636_), .ZN(new_n3637_));
  NOR2_X1    g03404(.A1(new_n2098_), .A2(new_n3371_), .ZN(new_n3638_));
  NOR2_X1    g03405(.A1(new_n566_), .A2(new_n1916_), .ZN(new_n3639_));
  INV_X1     g03406(.I(new_n3639_), .ZN(new_n3640_));
  NOR4_X1    g03407(.A1(new_n3637_), .A2(new_n3640_), .A3(new_n812_), .A4(new_n3638_), .ZN(new_n3641_));
  INV_X1     g03408(.I(new_n3641_), .ZN(new_n3642_));
  XOR2_X1    g03409(.A1(new_n3635_), .A2(new_n3642_), .Z(new_n3643_));
  NOR2_X1    g03410(.A1(new_n3643_), .A2(new_n3632_), .ZN(new_n3644_));
  NAND2_X1   g03411(.A1(new_n3635_), .A2(new_n3641_), .ZN(new_n3645_));
  NAND3_X1   g03412(.A1(new_n3634_), .A2(new_n3633_), .A3(new_n3642_), .ZN(new_n3646_));
  AOI21_X1   g03413(.A1(new_n3645_), .A2(new_n3646_), .B(new_n3631_), .ZN(new_n3647_));
  NOR2_X1    g03414(.A1(new_n3644_), .A2(new_n3647_), .ZN(new_n3648_));
  NAND2_X1   g03415(.A1(new_n3501_), .A2(new_n3502_), .ZN(new_n3649_));
  NOR2_X1    g03416(.A1(new_n786_), .A2(new_n2276_), .ZN(new_n3650_));
  NAND2_X1   g03417(.A1(\a[3] ), .A2(\a[35] ), .ZN(new_n3651_));
  XOR2_X1    g03418(.A1(new_n3650_), .A2(new_n3651_), .Z(new_n3652_));
  NOR2_X1    g03419(.A1(new_n1237_), .A2(new_n3393_), .ZN(new_n3653_));
  NAND2_X1   g03420(.A1(\a[36] ), .A2(\a[38] ), .ZN(new_n3654_));
  XNOR2_X1   g03421(.A1(new_n197_), .A2(new_n3654_), .ZN(new_n3655_));
  XNOR2_X1   g03422(.A1(new_n3652_), .A2(new_n3655_), .ZN(new_n3656_));
  NOR2_X1    g03423(.A1(new_n3656_), .A2(new_n3649_), .ZN(new_n3657_));
  INV_X1     g03424(.I(new_n3649_), .ZN(new_n3658_));
  NOR2_X1    g03425(.A1(new_n3652_), .A2(new_n3655_), .ZN(new_n3659_));
  INV_X1     g03426(.I(new_n3659_), .ZN(new_n3660_));
  NAND2_X1   g03427(.A1(new_n3652_), .A2(new_n3655_), .ZN(new_n3661_));
  AOI21_X1   g03428(.A1(new_n3660_), .A2(new_n3661_), .B(new_n3658_), .ZN(new_n3662_));
  NOR2_X1    g03429(.A1(new_n3657_), .A2(new_n3662_), .ZN(new_n3663_));
  XOR2_X1    g03430(.A1(new_n3648_), .A2(new_n3663_), .Z(new_n3664_));
  OAI21_X1   g03431(.A1(new_n3593_), .A2(new_n3630_), .B(new_n3664_), .ZN(new_n3665_));
  NOR2_X1    g03432(.A1(new_n3630_), .A2(new_n3593_), .ZN(new_n3666_));
  NOR2_X1    g03433(.A1(new_n3648_), .A2(new_n3663_), .ZN(new_n3667_));
  NAND2_X1   g03434(.A1(new_n3648_), .A2(new_n3663_), .ZN(new_n3668_));
  INV_X1     g03435(.I(new_n3668_), .ZN(new_n3669_));
  OAI21_X1   g03436(.A1(new_n3669_), .A2(new_n3667_), .B(new_n3666_), .ZN(new_n3670_));
  NAND2_X1   g03437(.A1(new_n3665_), .A2(new_n3670_), .ZN(new_n3671_));
  OAI21_X1   g03438(.A1(new_n3481_), .A2(new_n3492_), .B(new_n3491_), .ZN(new_n3672_));
  AOI21_X1   g03439(.A1(new_n3530_), .A2(new_n3533_), .B(new_n3526_), .ZN(new_n3673_));
  NOR2_X1    g03440(.A1(new_n3673_), .A2(new_n3534_), .ZN(new_n3674_));
  NOR2_X1    g03441(.A1(\a[8] ), .A2(\a[29] ), .ZN(new_n3675_));
  OAI21_X1   g03442(.A1(new_n1268_), .A2(new_n1715_), .B(new_n3675_), .ZN(new_n3676_));
  NAND2_X1   g03443(.A1(new_n3508_), .A2(new_n3676_), .ZN(new_n3677_));
  NAND2_X1   g03444(.A1(\a[1] ), .A2(\a[37] ), .ZN(new_n3678_));
  XNOR2_X1   g03445(.A1(new_n1536_), .A2(new_n3678_), .ZN(new_n3679_));
  XOR2_X1    g03446(.A1(new_n3677_), .A2(new_n3679_), .Z(new_n3680_));
  NOR3_X1    g03447(.A1(new_n3680_), .A2(new_n3483_), .A3(new_n3485_), .ZN(new_n3681_));
  NOR2_X1    g03448(.A1(new_n3485_), .A2(new_n3483_), .ZN(new_n3682_));
  INV_X1     g03449(.I(new_n3679_), .ZN(new_n3683_));
  NAND2_X1   g03450(.A1(new_n3683_), .A2(new_n3677_), .ZN(new_n3684_));
  NOR2_X1    g03451(.A1(new_n3683_), .A2(new_n3677_), .ZN(new_n3685_));
  INV_X1     g03452(.I(new_n3685_), .ZN(new_n3686_));
  AOI21_X1   g03453(.A1(new_n3686_), .A2(new_n3684_), .B(new_n3682_), .ZN(new_n3687_));
  NOR2_X1    g03454(.A1(new_n3687_), .A2(new_n3681_), .ZN(new_n3688_));
  XNOR2_X1   g03455(.A1(new_n3688_), .A2(new_n3674_), .ZN(new_n3689_));
  NAND2_X1   g03456(.A1(new_n3689_), .A2(new_n3672_), .ZN(new_n3690_));
  INV_X1     g03457(.I(new_n3688_), .ZN(new_n3691_));
  NAND2_X1   g03458(.A1(new_n3691_), .A2(new_n3674_), .ZN(new_n3692_));
  NOR2_X1    g03459(.A1(new_n3691_), .A2(new_n3674_), .ZN(new_n3693_));
  INV_X1     g03460(.I(new_n3693_), .ZN(new_n3694_));
  AOI21_X1   g03461(.A1(new_n3694_), .A2(new_n3692_), .B(new_n3672_), .ZN(new_n3695_));
  INV_X1     g03462(.I(new_n3695_), .ZN(new_n3696_));
  NAND2_X1   g03463(.A1(new_n3696_), .A2(new_n3690_), .ZN(new_n3697_));
  XOR2_X1    g03464(.A1(new_n3671_), .A2(new_n3697_), .Z(new_n3698_));
  NAND2_X1   g03465(.A1(new_n3698_), .A2(new_n3629_), .ZN(new_n3699_));
  INV_X1     g03466(.I(new_n3629_), .ZN(new_n3700_));
  INV_X1     g03467(.I(new_n3671_), .ZN(new_n3701_));
  INV_X1     g03468(.I(new_n3697_), .ZN(new_n3702_));
  NOR2_X1    g03469(.A1(new_n3701_), .A2(new_n3702_), .ZN(new_n3703_));
  NOR2_X1    g03470(.A1(new_n3671_), .A2(new_n3697_), .ZN(new_n3704_));
  OAI21_X1   g03471(.A1(new_n3703_), .A2(new_n3704_), .B(new_n3700_), .ZN(new_n3705_));
  NAND2_X1   g03472(.A1(new_n3699_), .A2(new_n3705_), .ZN(new_n3706_));
  NAND2_X1   g03473(.A1(new_n3522_), .A2(new_n3470_), .ZN(new_n3707_));
  AOI21_X1   g03474(.A1(new_n3555_), .A2(new_n3557_), .B(new_n3540_), .ZN(new_n3708_));
  NOR2_X1    g03475(.A1(new_n3708_), .A2(new_n3558_), .ZN(new_n3709_));
  NOR2_X1    g03476(.A1(new_n1018_), .A2(new_n2285_), .ZN(new_n3710_));
  NOR2_X1    g03477(.A1(new_n3531_), .A2(new_n3710_), .ZN(new_n3711_));
  INV_X1     g03478(.I(new_n3487_), .ZN(new_n3712_));
  NAND2_X1   g03479(.A1(new_n3712_), .A2(new_n225_), .ZN(new_n3713_));
  NOR2_X1    g03480(.A1(\a[16] ), .A2(\a[21] ), .ZN(new_n3714_));
  OAI21_X1   g03481(.A1(new_n225_), .A2(new_n3712_), .B(new_n3714_), .ZN(new_n3715_));
  NAND2_X1   g03482(.A1(new_n3715_), .A2(new_n3713_), .ZN(new_n3716_));
  XNOR2_X1   g03483(.A1(new_n3716_), .A2(new_n3711_), .ZN(new_n3717_));
  NAND3_X1   g03484(.A1(new_n3711_), .A2(new_n3713_), .A3(new_n3715_), .ZN(new_n3718_));
  OAI21_X1   g03485(.A1(new_n3531_), .A2(new_n3710_), .B(new_n3716_), .ZN(new_n3719_));
  AOI21_X1   g03486(.A1(new_n3719_), .A2(new_n3718_), .B(new_n3478_), .ZN(new_n3720_));
  AOI21_X1   g03487(.A1(new_n3717_), .A2(new_n3478_), .B(new_n3720_), .ZN(new_n3721_));
  OAI21_X1   g03488(.A1(new_n3499_), .A2(new_n3516_), .B(new_n3515_), .ZN(new_n3722_));
  INV_X1     g03489(.I(new_n3722_), .ZN(new_n3723_));
  NOR2_X1    g03490(.A1(new_n1274_), .A2(new_n1773_), .ZN(new_n3724_));
  NOR2_X1    g03491(.A1(new_n1274_), .A2(new_n1773_), .ZN(new_n3728_));
  INV_X1     g03492(.I(new_n3728_), .ZN(new_n3729_));
  NAND4_X1   g03493(.A1(\a[5] ), .A2(\a[6] ), .A3(\a[32] ), .A4(\a[33] ), .ZN(new_n3731_));
  INV_X1     g03494(.I(new_n3731_), .ZN(new_n3732_));
  NOR2_X1    g03495(.A1(new_n2499_), .A2(new_n2655_), .ZN(new_n3733_));
  INV_X1     g03496(.I(new_n3733_), .ZN(new_n3734_));
  OAI22_X1   g03497(.A1(new_n453_), .A2(new_n3734_), .B1(new_n3175_), .B2(new_n772_), .ZN(new_n3735_));
  NAND4_X1   g03498(.A1(new_n3127_), .A2(\a[9] ), .A3(\a[29] ), .A4(new_n392_), .ZN(new_n3736_));
  NOR2_X1    g03499(.A1(new_n3735_), .A2(new_n3736_), .ZN(new_n3737_));
  NAND2_X1   g03500(.A1(new_n3737_), .A2(new_n3732_), .ZN(new_n3738_));
  OAI21_X1   g03501(.A1(new_n3735_), .A2(new_n3736_), .B(new_n3731_), .ZN(new_n3739_));
  AOI21_X1   g03502(.A1(new_n3738_), .A2(new_n3739_), .B(new_n3729_), .ZN(new_n3740_));
  XOR2_X1    g03503(.A1(new_n3737_), .A2(new_n3731_), .Z(new_n3741_));
  NOR2_X1    g03504(.A1(new_n3741_), .A2(new_n3728_), .ZN(new_n3742_));
  NOR2_X1    g03505(.A1(new_n3742_), .A2(new_n3740_), .ZN(new_n3743_));
  NOR2_X1    g03506(.A1(new_n3723_), .A2(new_n3743_), .ZN(new_n3744_));
  INV_X1     g03507(.I(new_n3744_), .ZN(new_n3745_));
  NAND2_X1   g03508(.A1(new_n3723_), .A2(new_n3743_), .ZN(new_n3746_));
  AOI21_X1   g03509(.A1(new_n3745_), .A2(new_n3746_), .B(new_n3721_), .ZN(new_n3747_));
  INV_X1     g03510(.I(new_n3721_), .ZN(new_n3748_));
  XOR2_X1    g03511(.A1(new_n3743_), .A2(new_n3722_), .Z(new_n3749_));
  NOR2_X1    g03512(.A1(new_n3749_), .A2(new_n3748_), .ZN(new_n3750_));
  OAI21_X1   g03513(.A1(new_n3747_), .A2(new_n3750_), .B(new_n3709_), .ZN(new_n3751_));
  NOR2_X1    g03514(.A1(new_n3750_), .A2(new_n3747_), .ZN(new_n3752_));
  OAI21_X1   g03515(.A1(new_n3558_), .A2(new_n3708_), .B(new_n3752_), .ZN(new_n3753_));
  AOI22_X1   g03516(.A1(new_n3753_), .A2(new_n3751_), .B1(new_n3523_), .B2(new_n3707_), .ZN(new_n3754_));
  NAND2_X1   g03517(.A1(new_n3707_), .A2(new_n3523_), .ZN(new_n3755_));
  XOR2_X1    g03518(.A1(new_n3752_), .A2(new_n3709_), .Z(new_n3756_));
  NOR2_X1    g03519(.A1(new_n3756_), .A2(new_n3755_), .ZN(new_n3757_));
  NOR2_X1    g03520(.A1(new_n3757_), .A2(new_n3754_), .ZN(new_n3758_));
  INV_X1     g03521(.I(new_n3758_), .ZN(new_n3759_));
  XOR2_X1    g03522(.A1(new_n3706_), .A2(new_n3759_), .Z(new_n3760_));
  NOR2_X1    g03523(.A1(new_n3760_), .A2(new_n3627_), .ZN(new_n3761_));
  INV_X1     g03524(.I(new_n3627_), .ZN(new_n3762_));
  NAND3_X1   g03525(.A1(new_n3699_), .A2(new_n3705_), .A3(new_n3759_), .ZN(new_n3763_));
  NAND2_X1   g03526(.A1(new_n3706_), .A2(new_n3758_), .ZN(new_n3764_));
  AOI21_X1   g03527(.A1(new_n3764_), .A2(new_n3763_), .B(new_n3762_), .ZN(new_n3765_));
  NOR2_X1    g03528(.A1(new_n3761_), .A2(new_n3765_), .ZN(new_n3766_));
  NOR2_X1    g03529(.A1(new_n3766_), .A2(new_n3625_), .ZN(new_n3767_));
  XNOR2_X1   g03530(.A1(new_n3623_), .A2(new_n3767_), .ZN(new_n3768_));
  XOR2_X1    g03531(.A1(new_n3768_), .A2(new_n3615_), .Z(\asquared[39] ));
  AOI21_X1   g03532(.A1(new_n3766_), .A2(new_n3625_), .B(new_n3615_), .ZN(new_n3770_));
  AOI21_X1   g03533(.A1(new_n3623_), .A2(new_n3770_), .B(new_n3767_), .ZN(new_n3771_));
  NAND2_X1   g03534(.A1(new_n3764_), .A2(new_n3762_), .ZN(new_n3772_));
  AND2_X2    g03535(.A1(new_n3772_), .A2(new_n3763_), .Z(new_n3773_));
  INV_X1     g03536(.I(new_n3704_), .ZN(new_n3774_));
  OAI21_X1   g03537(.A1(new_n3700_), .A2(new_n3703_), .B(new_n3774_), .ZN(new_n3775_));
  INV_X1     g03538(.I(new_n3775_), .ZN(new_n3776_));
  OAI21_X1   g03539(.A1(new_n3666_), .A2(new_n3667_), .B(new_n3668_), .ZN(new_n3777_));
  INV_X1     g03540(.I(new_n3777_), .ZN(new_n3778_));
  AOI21_X1   g03541(.A1(new_n3682_), .A2(new_n3684_), .B(new_n3685_), .ZN(new_n3779_));
  INV_X1     g03542(.I(new_n3779_), .ZN(new_n3780_));
  NAND2_X1   g03543(.A1(new_n3719_), .A2(new_n3478_), .ZN(new_n3781_));
  NAND2_X1   g03544(.A1(new_n3781_), .A2(new_n3718_), .ZN(new_n3782_));
  INV_X1     g03545(.I(\a[39] ), .ZN(new_n3783_));
  NOR2_X1    g03546(.A1(new_n1536_), .A2(new_n3678_), .ZN(new_n3784_));
  INV_X1     g03547(.I(new_n3784_), .ZN(new_n3785_));
  AOI21_X1   g03548(.A1(\a[1] ), .A2(\a[38] ), .B(\a[20] ), .ZN(new_n3786_));
  NAND2_X1   g03549(.A1(new_n1315_), .A2(\a[38] ), .ZN(new_n3787_));
  INV_X1     g03550(.I(new_n3787_), .ZN(new_n3788_));
  NOR2_X1    g03551(.A1(new_n3788_), .A2(new_n3786_), .ZN(new_n3789_));
  NOR2_X1    g03552(.A1(new_n3789_), .A2(new_n3785_), .ZN(new_n3790_));
  XOR2_X1    g03553(.A1(new_n3790_), .A2(new_n199_), .Z(new_n3791_));
  XOR2_X1    g03554(.A1(new_n3791_), .A2(new_n3783_), .Z(new_n3792_));
  XOR2_X1    g03555(.A1(new_n3792_), .A2(new_n3782_), .Z(new_n3793_));
  NAND2_X1   g03556(.A1(new_n3793_), .A2(new_n3780_), .ZN(new_n3794_));
  AND2_X2    g03557(.A1(new_n3792_), .A2(new_n3782_), .Z(new_n3795_));
  NOR2_X1    g03558(.A1(new_n3792_), .A2(new_n3782_), .ZN(new_n3796_));
  OAI21_X1   g03559(.A1(new_n3795_), .A2(new_n3796_), .B(new_n3779_), .ZN(new_n3797_));
  NAND2_X1   g03560(.A1(new_n3794_), .A2(new_n3797_), .ZN(new_n3798_));
  AOI21_X1   g03561(.A1(new_n1719_), .A2(new_n2286_), .B(new_n3724_), .ZN(new_n3799_));
  INV_X1     g03562(.I(new_n3799_), .ZN(new_n3800_));
  NOR2_X1    g03563(.A1(\a[3] ), .A2(\a[35] ), .ZN(new_n3801_));
  OAI21_X1   g03564(.A1(new_n786_), .A2(new_n2276_), .B(new_n3801_), .ZN(new_n3802_));
  OAI21_X1   g03565(.A1(new_n787_), .A2(new_n2277_), .B(new_n3802_), .ZN(new_n3803_));
  INV_X1     g03566(.I(\a[38] ), .ZN(new_n3804_));
  NOR2_X1    g03567(.A1(new_n3393_), .A2(new_n3804_), .ZN(new_n3805_));
  AOI21_X1   g03568(.A1(new_n3653_), .A2(new_n218_), .B(new_n3805_), .ZN(new_n3806_));
  XNOR2_X1   g03569(.A1(new_n3803_), .A2(new_n3806_), .ZN(new_n3807_));
  NOR2_X1    g03570(.A1(new_n3807_), .A2(new_n3800_), .ZN(new_n3808_));
  NOR2_X1    g03571(.A1(new_n3803_), .A2(new_n3806_), .ZN(new_n3809_));
  INV_X1     g03572(.I(new_n3809_), .ZN(new_n3810_));
  NAND2_X1   g03573(.A1(new_n3803_), .A2(new_n3806_), .ZN(new_n3811_));
  AOI21_X1   g03574(.A1(new_n3810_), .A2(new_n3811_), .B(new_n3799_), .ZN(new_n3812_));
  NOR2_X1    g03575(.A1(new_n3808_), .A2(new_n3812_), .ZN(new_n3813_));
  NAND2_X1   g03576(.A1(new_n3739_), .A2(new_n3728_), .ZN(new_n3814_));
  NAND2_X1   g03577(.A1(new_n3814_), .A2(new_n3738_), .ZN(new_n3815_));
  INV_X1     g03578(.I(new_n3815_), .ZN(new_n3816_));
  NAND2_X1   g03579(.A1(new_n3658_), .A2(new_n3661_), .ZN(new_n3817_));
  NAND2_X1   g03580(.A1(new_n3817_), .A2(new_n3660_), .ZN(new_n3818_));
  INV_X1     g03581(.I(new_n3818_), .ZN(new_n3819_));
  NOR2_X1    g03582(.A1(new_n3819_), .A2(new_n3816_), .ZN(new_n3820_));
  NOR2_X1    g03583(.A1(new_n3818_), .A2(new_n3815_), .ZN(new_n3821_));
  NOR2_X1    g03584(.A1(new_n3820_), .A2(new_n3821_), .ZN(new_n3822_));
  NOR2_X1    g03585(.A1(new_n3822_), .A2(new_n3813_), .ZN(new_n3823_));
  XNOR2_X1   g03586(.A1(new_n3818_), .A2(new_n3815_), .ZN(new_n3824_));
  INV_X1     g03587(.I(new_n3824_), .ZN(new_n3825_));
  AOI21_X1   g03588(.A1(new_n3813_), .A2(new_n3825_), .B(new_n3823_), .ZN(new_n3826_));
  XOR2_X1    g03589(.A1(new_n3798_), .A2(new_n3826_), .Z(new_n3827_));
  NOR2_X1    g03590(.A1(new_n3827_), .A2(new_n3778_), .ZN(new_n3828_));
  INV_X1     g03591(.I(new_n3798_), .ZN(new_n3829_));
  NOR2_X1    g03592(.A1(new_n3829_), .A2(new_n3826_), .ZN(new_n3830_));
  INV_X1     g03593(.I(new_n3830_), .ZN(new_n3831_));
  NAND2_X1   g03594(.A1(new_n3829_), .A2(new_n3826_), .ZN(new_n3832_));
  AOI21_X1   g03595(.A1(new_n3831_), .A2(new_n3832_), .B(new_n3777_), .ZN(new_n3833_));
  NOR2_X1    g03596(.A1(new_n3833_), .A2(new_n3828_), .ZN(new_n3834_));
  NAND2_X1   g03597(.A1(new_n3751_), .A2(new_n3755_), .ZN(new_n3835_));
  AOI21_X1   g03598(.A1(new_n3672_), .A2(new_n3692_), .B(new_n3693_), .ZN(new_n3836_));
  INV_X1     g03599(.I(\a[37] ), .ZN(new_n3837_));
  NOR2_X1    g03600(.A1(new_n3393_), .A2(new_n3837_), .ZN(new_n3838_));
  INV_X1     g03601(.I(new_n3838_), .ZN(new_n3839_));
  NAND2_X1   g03602(.A1(\a[13] ), .A2(\a[36] ), .ZN(new_n3840_));
  NOR3_X1    g03603(.A1(new_n3840_), .A2(new_n200_), .A3(new_n1916_), .ZN(new_n3841_));
  NAND4_X1   g03604(.A1(new_n3841_), .A2(\a[13] ), .A3(new_n2191_), .A4(\a[37] ), .ZN(new_n3842_));
  AOI21_X1   g03605(.A1(new_n3842_), .A2(new_n3839_), .B(new_n225_), .ZN(new_n3843_));
  NOR3_X1    g03606(.A1(new_n3843_), .A2(new_n201_), .A3(new_n3837_), .ZN(new_n3844_));
  OR2_X2     g03607(.A1(new_n3843_), .A2(new_n3841_), .Z(new_n3845_));
  INV_X1     g03608(.I(new_n3845_), .ZN(new_n3846_));
  AOI22_X1   g03609(.A1(\a[3] ), .A2(\a[13] ), .B1(\a[26] ), .B2(\a[36] ), .ZN(new_n3847_));
  AOI21_X1   g03610(.A1(new_n3846_), .A2(new_n3847_), .B(new_n3844_), .ZN(new_n3848_));
  INV_X1     g03611(.I(new_n2766_), .ZN(new_n3849_));
  NOR2_X1    g03612(.A1(new_n242_), .A2(new_n2868_), .ZN(new_n3850_));
  NOR2_X1    g03613(.A1(new_n2765_), .A2(new_n2868_), .ZN(new_n3851_));
  INV_X1     g03614(.I(new_n3851_), .ZN(new_n3852_));
  NOR2_X1    g03615(.A1(new_n3849_), .A2(new_n772_), .ZN(new_n3853_));
  NAND4_X1   g03616(.A1(new_n3853_), .A2(\a[9] ), .A3(new_n3850_), .A4(\a[30] ), .ZN(new_n3854_));
  AOI21_X1   g03617(.A1(new_n3854_), .A2(new_n3852_), .B(new_n478_), .ZN(new_n3855_));
  NOR2_X1    g03618(.A1(new_n3849_), .A2(new_n772_), .ZN(new_n3856_));
  INV_X1     g03619(.I(new_n3856_), .ZN(new_n3857_));
  AOI22_X1   g03620(.A1(new_n1718_), .A2(new_n2277_), .B1(new_n1447_), .B2(new_n1913_), .ZN(new_n3858_));
  NOR4_X1    g03621(.A1(new_n1719_), .A2(new_n2543_), .A3(new_n650_), .A4(new_n1999_), .ZN(new_n3859_));
  NAND2_X1   g03622(.A1(new_n3858_), .A2(new_n3859_), .ZN(new_n3860_));
  NOR2_X1    g03623(.A1(new_n3860_), .A2(new_n3857_), .ZN(new_n3861_));
  INV_X1     g03624(.I(new_n3861_), .ZN(new_n3862_));
  NAND2_X1   g03625(.A1(new_n3860_), .A2(new_n3857_), .ZN(new_n3863_));
  NAND2_X1   g03626(.A1(new_n3862_), .A2(new_n3863_), .ZN(new_n3864_));
  NAND2_X1   g03627(.A1(new_n3848_), .A2(new_n3864_), .ZN(new_n3865_));
  XOR2_X1    g03628(.A1(new_n3860_), .A2(new_n3856_), .Z(new_n3866_));
  OAI21_X1   g03629(.A1(new_n3848_), .A2(new_n3866_), .B(new_n3865_), .ZN(new_n3867_));
  AOI21_X1   g03630(.A1(new_n3723_), .A2(new_n3743_), .B(new_n3748_), .ZN(new_n3868_));
  NOR2_X1    g03631(.A1(new_n3868_), .A2(new_n3744_), .ZN(new_n3869_));
  XOR2_X1    g03632(.A1(new_n3869_), .A2(new_n3867_), .Z(new_n3870_));
  INV_X1     g03633(.I(new_n3869_), .ZN(new_n3871_));
  NAND2_X1   g03634(.A1(new_n3871_), .A2(new_n3867_), .ZN(new_n3872_));
  INV_X1     g03635(.I(new_n3872_), .ZN(new_n3873_));
  NOR2_X1    g03636(.A1(new_n3871_), .A2(new_n3867_), .ZN(new_n3874_));
  OAI21_X1   g03637(.A1(new_n3873_), .A2(new_n3874_), .B(new_n3836_), .ZN(new_n3875_));
  OAI21_X1   g03638(.A1(new_n3836_), .A2(new_n3870_), .B(new_n3875_), .ZN(new_n3876_));
  NAND2_X1   g03639(.A1(new_n3646_), .A2(new_n3631_), .ZN(new_n3877_));
  NAND2_X1   g03640(.A1(new_n3877_), .A2(new_n3645_), .ZN(new_n3878_));
  INV_X1     g03641(.I(new_n3878_), .ZN(new_n3879_));
  NAND2_X1   g03642(.A1(\a[10] ), .A2(\a[11] ), .ZN(new_n3881_));
  NOR2_X1    g03643(.A1(new_n2689_), .A2(new_n3881_), .ZN(new_n3882_));
  NOR4_X1    g03644(.A1(new_n353_), .A2(new_n461_), .A3(new_n2499_), .A4(new_n3371_), .ZN(new_n3883_));
  NOR2_X1    g03645(.A1(new_n3883_), .A2(new_n3882_), .ZN(new_n3884_));
  INV_X1     g03646(.I(new_n3884_), .ZN(new_n3885_));
  OAI21_X1   g03647(.A1(new_n2499_), .A2(new_n3371_), .B(new_n3025_), .ZN(new_n3886_));
  OAI22_X1   g03648(.A1(new_n3885_), .A2(new_n3886_), .B1(new_n2180_), .B2(new_n3882_), .ZN(new_n3887_));
  NAND2_X1   g03649(.A1(new_n2331_), .A2(new_n2978_), .ZN(new_n3888_));
  NAND2_X1   g03650(.A1(\a[18] ), .A2(\a[21] ), .ZN(new_n3889_));
  NAND2_X1   g03651(.A1(new_n1715_), .A2(new_n3889_), .ZN(new_n3890_));
  NOR2_X1    g03652(.A1(new_n3888_), .A2(new_n3890_), .ZN(new_n3891_));
  NOR2_X1    g03653(.A1(new_n359_), .A2(new_n2655_), .ZN(new_n3892_));
  XNOR2_X1   g03654(.A1(new_n3891_), .A2(new_n3892_), .ZN(new_n3893_));
  NOR2_X1    g03655(.A1(new_n566_), .A2(new_n2098_), .ZN(new_n3894_));
  NAND3_X1   g03656(.A1(new_n3894_), .A2(\a[17] ), .A3(\a[22] ), .ZN(new_n3895_));
  XOR2_X1    g03657(.A1(new_n3895_), .A2(\a[4] ), .Z(new_n3896_));
  NOR2_X1    g03658(.A1(new_n3896_), .A2(\a[35] ), .ZN(new_n3897_));
  AND2_X2    g03659(.A1(new_n3896_), .A2(\a[35] ), .Z(new_n3898_));
  NOR2_X1    g03660(.A1(new_n3898_), .A2(new_n3897_), .ZN(new_n3899_));
  NOR2_X1    g03661(.A1(new_n3899_), .A2(new_n3893_), .ZN(new_n3900_));
  INV_X1     g03662(.I(new_n3900_), .ZN(new_n3901_));
  NAND2_X1   g03663(.A1(new_n3899_), .A2(new_n3893_), .ZN(new_n3902_));
  AOI21_X1   g03664(.A1(new_n3901_), .A2(new_n3902_), .B(new_n3887_), .ZN(new_n3903_));
  INV_X1     g03665(.I(new_n3887_), .ZN(new_n3904_));
  XNOR2_X1   g03666(.A1(new_n3899_), .A2(new_n3893_), .ZN(new_n3905_));
  NOR2_X1    g03667(.A1(new_n3905_), .A2(new_n3904_), .ZN(new_n3906_));
  NOR2_X1    g03668(.A1(new_n3906_), .A2(new_n3903_), .ZN(new_n3907_));
  NOR4_X1    g03669(.A1(new_n353_), .A2(new_n242_), .A3(new_n2765_), .A4(new_n2868_), .ZN(new_n3908_));
  INV_X1     g03670(.I(new_n3908_), .ZN(new_n3909_));
  OAI21_X1   g03671(.A1(new_n392_), .A2(new_n3127_), .B(new_n3735_), .ZN(new_n3910_));
  NAND2_X1   g03672(.A1(new_n3638_), .A2(new_n812_), .ZN(new_n3911_));
  NAND2_X1   g03673(.A1(new_n3637_), .A2(new_n3911_), .ZN(new_n3912_));
  XNOR2_X1   g03674(.A1(new_n3910_), .A2(new_n3912_), .ZN(new_n3913_));
  NOR2_X1    g03675(.A1(new_n3913_), .A2(new_n3909_), .ZN(new_n3914_));
  NOR2_X1    g03676(.A1(new_n3910_), .A2(new_n3912_), .ZN(new_n3915_));
  INV_X1     g03677(.I(new_n3915_), .ZN(new_n3916_));
  NAND2_X1   g03678(.A1(new_n3910_), .A2(new_n3912_), .ZN(new_n3917_));
  AOI21_X1   g03679(.A1(new_n3916_), .A2(new_n3917_), .B(new_n3908_), .ZN(new_n3918_));
  NOR2_X1    g03680(.A1(new_n3914_), .A2(new_n3918_), .ZN(new_n3919_));
  XOR2_X1    g03681(.A1(new_n3907_), .A2(new_n3919_), .Z(new_n3920_));
  INV_X1     g03682(.I(new_n3907_), .ZN(new_n3921_));
  NOR2_X1    g03683(.A1(new_n3921_), .A2(new_n3919_), .ZN(new_n3922_));
  INV_X1     g03684(.I(new_n3919_), .ZN(new_n3923_));
  NOR2_X1    g03685(.A1(new_n3907_), .A2(new_n3923_), .ZN(new_n3924_));
  OAI21_X1   g03686(.A1(new_n3922_), .A2(new_n3924_), .B(new_n3879_), .ZN(new_n3925_));
  OAI21_X1   g03687(.A1(new_n3879_), .A2(new_n3920_), .B(new_n3925_), .ZN(new_n3926_));
  NAND2_X1   g03688(.A1(new_n3876_), .A2(new_n3926_), .ZN(new_n3927_));
  OR2_X2     g03689(.A1(new_n3876_), .A2(new_n3926_), .Z(new_n3928_));
  AOI22_X1   g03690(.A1(new_n3928_), .A2(new_n3927_), .B1(new_n3753_), .B2(new_n3835_), .ZN(new_n3929_));
  NAND2_X1   g03691(.A1(new_n3835_), .A2(new_n3753_), .ZN(new_n3930_));
  XNOR2_X1   g03692(.A1(new_n3876_), .A2(new_n3926_), .ZN(new_n3931_));
  NOR2_X1    g03693(.A1(new_n3931_), .A2(new_n3930_), .ZN(new_n3932_));
  NOR2_X1    g03694(.A1(new_n3932_), .A2(new_n3929_), .ZN(new_n3933_));
  XOR2_X1    g03695(.A1(new_n3933_), .A2(new_n3834_), .Z(new_n3934_));
  NOR2_X1    g03696(.A1(new_n3934_), .A2(new_n3776_), .ZN(new_n3935_));
  OAI21_X1   g03697(.A1(new_n3932_), .A2(new_n3929_), .B(new_n3834_), .ZN(new_n3936_));
  OAI21_X1   g03698(.A1(new_n3828_), .A2(new_n3833_), .B(new_n3933_), .ZN(new_n3937_));
  AOI21_X1   g03699(.A1(new_n3937_), .A2(new_n3936_), .B(new_n3775_), .ZN(new_n3938_));
  NOR2_X1    g03700(.A1(new_n3935_), .A2(new_n3938_), .ZN(new_n3939_));
  XOR2_X1    g03701(.A1(new_n3939_), .A2(new_n3773_), .Z(new_n3940_));
  OAI21_X1   g03702(.A1(new_n3935_), .A2(new_n3938_), .B(new_n3773_), .ZN(new_n3941_));
  INV_X1     g03703(.I(new_n3773_), .ZN(new_n3942_));
  NAND2_X1   g03704(.A1(new_n3942_), .A2(new_n3939_), .ZN(new_n3943_));
  NAND2_X1   g03705(.A1(new_n3943_), .A2(new_n3941_), .ZN(new_n3944_));
  NAND2_X1   g03706(.A1(new_n3771_), .A2(new_n3944_), .ZN(new_n3945_));
  OAI21_X1   g03707(.A1(new_n3771_), .A2(new_n3940_), .B(new_n3945_), .ZN(\asquared[40] ));
  NOR2_X1    g03708(.A1(new_n3942_), .A2(new_n3939_), .ZN(new_n3947_));
  OAI21_X1   g03709(.A1(new_n3771_), .A2(new_n3947_), .B(new_n3943_), .ZN(new_n3948_));
  NAND2_X1   g03710(.A1(new_n3937_), .A2(new_n3775_), .ZN(new_n3949_));
  NAND2_X1   g03711(.A1(new_n3949_), .A2(new_n3936_), .ZN(new_n3950_));
  OAI21_X1   g03712(.A1(new_n3778_), .A2(new_n3830_), .B(new_n3832_), .ZN(new_n3951_));
  NOR2_X1    g03713(.A1(new_n3796_), .A2(new_n3779_), .ZN(new_n3952_));
  AOI21_X1   g03714(.A1(new_n1719_), .A2(new_n2543_), .B(new_n3858_), .ZN(new_n3953_));
  NAND2_X1   g03715(.A1(\a[0] ), .A2(\a[39] ), .ZN(new_n3954_));
  AOI21_X1   g03716(.A1(new_n3789_), .A2(new_n3785_), .B(new_n3954_), .ZN(new_n3955_));
  NOR2_X1    g03717(.A1(new_n3955_), .A2(new_n3790_), .ZN(new_n3956_));
  XOR2_X1    g03718(.A1(new_n3956_), .A2(new_n3953_), .Z(new_n3957_));
  NOR3_X1    g03719(.A1(new_n3957_), .A2(new_n3853_), .A3(new_n3855_), .ZN(new_n3958_));
  NOR2_X1    g03720(.A1(new_n3855_), .A2(new_n3853_), .ZN(new_n3959_));
  INV_X1     g03721(.I(new_n3953_), .ZN(new_n3960_));
  NOR2_X1    g03722(.A1(new_n3956_), .A2(new_n3960_), .ZN(new_n3961_));
  INV_X1     g03723(.I(new_n3961_), .ZN(new_n3962_));
  NAND2_X1   g03724(.A1(new_n3956_), .A2(new_n3960_), .ZN(new_n3963_));
  AOI21_X1   g03725(.A1(new_n3962_), .A2(new_n3963_), .B(new_n3959_), .ZN(new_n3964_));
  NOR2_X1    g03726(.A1(new_n3958_), .A2(new_n3964_), .ZN(new_n3965_));
  NOR2_X1    g03727(.A1(new_n3423_), .A2(new_n3393_), .ZN(new_n3966_));
  INV_X1     g03728(.I(new_n3966_), .ZN(new_n3967_));
  NOR2_X1    g03729(.A1(new_n566_), .A2(new_n3423_), .ZN(new_n3968_));
  NOR2_X1    g03730(.A1(new_n566_), .A2(new_n3393_), .ZN(new_n3969_));
  NAND2_X1   g03731(.A1(\a[4] ), .A2(\a[5] ), .ZN(new_n3970_));
  NOR2_X1    g03732(.A1(new_n3967_), .A2(new_n3970_), .ZN(new_n3971_));
  INV_X1     g03733(.I(new_n3971_), .ZN(new_n3972_));
  NOR2_X1    g03734(.A1(new_n282_), .A2(new_n3393_), .ZN(new_n3973_));
  NAND2_X1   g03735(.A1(new_n2892_), .A2(new_n3968_), .ZN(new_n3974_));
  NAND2_X1   g03736(.A1(new_n3972_), .A2(new_n3974_), .ZN(new_n3975_));
  INV_X1     g03737(.I(new_n3975_), .ZN(new_n3976_));
  AOI21_X1   g03738(.A1(\a[28] ), .A2(\a[35] ), .B(new_n972_), .ZN(new_n3977_));
  AOI22_X1   g03739(.A1(new_n3976_), .A2(new_n3977_), .B1(new_n3972_), .B2(new_n3973_), .ZN(new_n3978_));
  NAND2_X1   g03740(.A1(new_n2869_), .A2(new_n3851_), .ZN(new_n3979_));
  NAND2_X1   g03741(.A1(new_n3979_), .A2(new_n1779_), .ZN(new_n3980_));
  NOR2_X1    g03742(.A1(new_n2655_), .A2(new_n2765_), .ZN(new_n3981_));
  NOR4_X1    g03743(.A1(new_n3981_), .A2(new_n454_), .A3(new_n268_), .A4(new_n2868_), .ZN(new_n3982_));
  INV_X1     g03744(.I(new_n3982_), .ZN(new_n3983_));
  NOR2_X1    g03745(.A1(new_n3983_), .A2(new_n3980_), .ZN(new_n3984_));
  INV_X1     g03746(.I(new_n3984_), .ZN(new_n3985_));
  NAND2_X1   g03747(.A1(\a[38] ), .A2(\a[40] ), .ZN(new_n3986_));
  XNOR2_X1   g03748(.A1(new_n197_), .A2(new_n3986_), .ZN(new_n3987_));
  NOR2_X1    g03749(.A1(new_n3985_), .A2(new_n3987_), .ZN(new_n3988_));
  INV_X1     g03750(.I(new_n3987_), .ZN(new_n3989_));
  NOR2_X1    g03751(.A1(new_n3984_), .A2(new_n3989_), .ZN(new_n3990_));
  NOR2_X1    g03752(.A1(new_n3988_), .A2(new_n3990_), .ZN(new_n3991_));
  XOR2_X1    g03753(.A1(new_n3984_), .A2(new_n3987_), .Z(new_n3992_));
  MUX2_X1    g03754(.I0(new_n3992_), .I1(new_n3991_), .S(new_n3978_), .Z(new_n3993_));
  XNOR2_X1   g03755(.A1(new_n3965_), .A2(new_n3993_), .ZN(new_n3994_));
  OAI21_X1   g03756(.A1(new_n3795_), .A2(new_n3952_), .B(new_n3994_), .ZN(new_n3995_));
  NOR2_X1    g03757(.A1(new_n3952_), .A2(new_n3795_), .ZN(new_n3996_));
  INV_X1     g03758(.I(new_n3965_), .ZN(new_n3997_));
  NOR2_X1    g03759(.A1(new_n3997_), .A2(new_n3993_), .ZN(new_n3998_));
  NAND2_X1   g03760(.A1(new_n3997_), .A2(new_n3993_), .ZN(new_n3999_));
  INV_X1     g03761(.I(new_n3999_), .ZN(new_n4000_));
  OAI21_X1   g03762(.A1(new_n4000_), .A2(new_n3998_), .B(new_n3996_), .ZN(new_n4001_));
  NAND2_X1   g03763(.A1(new_n3995_), .A2(new_n4001_), .ZN(new_n4002_));
  INV_X1     g03764(.I(new_n4002_), .ZN(new_n4003_));
  INV_X1     g03765(.I(new_n3821_), .ZN(new_n4004_));
  AOI21_X1   g03766(.A1(new_n3813_), .A2(new_n4004_), .B(new_n3820_), .ZN(new_n4005_));
  AOI21_X1   g03767(.A1(new_n3799_), .A2(new_n3811_), .B(new_n3809_), .ZN(new_n4006_));
  INV_X1     g03768(.I(new_n4006_), .ZN(new_n4007_));
  AOI21_X1   g03769(.A1(new_n3910_), .A2(new_n3912_), .B(new_n3909_), .ZN(new_n4008_));
  NOR2_X1    g03770(.A1(new_n4008_), .A2(new_n3915_), .ZN(new_n4009_));
  INV_X1     g03771(.I(new_n4009_), .ZN(new_n4010_));
  NOR2_X1    g03772(.A1(\a[8] ), .A2(\a[31] ), .ZN(new_n4011_));
  AOI21_X1   g03773(.A1(new_n3888_), .A2(new_n4011_), .B(new_n3890_), .ZN(new_n4012_));
  INV_X1     g03774(.I(new_n4012_), .ZN(new_n4013_));
  NAND2_X1   g03775(.A1(\a[1] ), .A2(\a[39] ), .ZN(new_n4014_));
  INV_X1     g03776(.I(new_n4014_), .ZN(new_n4015_));
  NOR2_X1    g03777(.A1(new_n4015_), .A2(new_n1710_), .ZN(new_n4016_));
  NOR2_X1    g03778(.A1(new_n1769_), .A2(new_n4014_), .ZN(new_n4017_));
  NOR2_X1    g03779(.A1(new_n4016_), .A2(new_n4017_), .ZN(new_n4018_));
  XOR2_X1    g03780(.A1(new_n4018_), .A2(new_n3788_), .Z(new_n4019_));
  NOR2_X1    g03781(.A1(new_n4019_), .A2(new_n4013_), .ZN(new_n4020_));
  INV_X1     g03782(.I(new_n4018_), .ZN(new_n4021_));
  NAND2_X1   g03783(.A1(new_n4021_), .A2(new_n3788_), .ZN(new_n4022_));
  NOR2_X1    g03784(.A1(new_n4021_), .A2(new_n3788_), .ZN(new_n4023_));
  INV_X1     g03785(.I(new_n4023_), .ZN(new_n4024_));
  AOI21_X1   g03786(.A1(new_n4024_), .A2(new_n4022_), .B(new_n4012_), .ZN(new_n4025_));
  NOR2_X1    g03787(.A1(new_n4025_), .A2(new_n4020_), .ZN(new_n4026_));
  XOR2_X1    g03788(.A1(new_n4026_), .A2(new_n4010_), .Z(new_n4027_));
  NAND2_X1   g03789(.A1(new_n4027_), .A2(new_n4007_), .ZN(new_n4028_));
  NOR2_X1    g03790(.A1(new_n4026_), .A2(new_n4010_), .ZN(new_n4029_));
  NOR3_X1    g03791(.A1(new_n4009_), .A2(new_n4025_), .A3(new_n4020_), .ZN(new_n4030_));
  OAI21_X1   g03792(.A1(new_n4029_), .A2(new_n4030_), .B(new_n4006_), .ZN(new_n4031_));
  NAND2_X1   g03793(.A1(new_n4028_), .A2(new_n4031_), .ZN(new_n4032_));
  NOR4_X1    g03794(.A1(new_n242_), .A2(new_n461_), .A3(new_n2461_), .A4(new_n3371_), .ZN(new_n4033_));
  NOR3_X1    g03795(.A1(new_n879_), .A2(new_n2499_), .A3(new_n3371_), .ZN(new_n4034_));
  NAND2_X1   g03796(.A1(new_n4033_), .A2(new_n4034_), .ZN(new_n4035_));
  AOI21_X1   g03797(.A1(new_n4035_), .A2(new_n796_), .B(new_n3175_), .ZN(new_n4036_));
  NAND2_X1   g03798(.A1(\a[11] ), .A2(\a[29] ), .ZN(new_n4037_));
  INV_X1     g03799(.I(new_n4033_), .ZN(new_n4038_));
  OAI21_X1   g03800(.A1(new_n796_), .A2(new_n3175_), .B(new_n4038_), .ZN(new_n4039_));
  NOR2_X1    g03801(.A1(new_n2461_), .A2(new_n3371_), .ZN(new_n4040_));
  INV_X1     g03802(.I(new_n4040_), .ZN(new_n4041_));
  OAI21_X1   g03803(.A1(new_n242_), .A2(new_n461_), .B(new_n4041_), .ZN(new_n4042_));
  OAI22_X1   g03804(.A1(new_n4036_), .A2(new_n4037_), .B1(new_n4039_), .B2(new_n4042_), .ZN(new_n4043_));
  NAND2_X1   g03805(.A1(new_n2533_), .A2(new_n787_), .ZN(new_n4044_));
  NAND2_X1   g03806(.A1(\a[3] ), .A2(\a[37] ), .ZN(new_n4045_));
  XNOR2_X1   g03807(.A1(new_n4044_), .A2(new_n4045_), .ZN(new_n4046_));
  INV_X1     g03808(.I(new_n4046_), .ZN(new_n4047_));
  NOR2_X1    g03809(.A1(new_n1912_), .A2(new_n2276_), .ZN(new_n4048_));
  NOR2_X1    g03810(.A1(new_n1021_), .A2(new_n1141_), .ZN(new_n4049_));
  NAND4_X1   g03811(.A1(new_n1274_), .A2(new_n1956_), .A3(\a[15] ), .A4(\a[25] ), .ZN(new_n4050_));
  NOR3_X1    g03812(.A1(new_n4050_), .A2(new_n4048_), .A3(new_n4049_), .ZN(new_n4051_));
  NAND2_X1   g03813(.A1(new_n4047_), .A2(new_n4051_), .ZN(new_n4052_));
  INV_X1     g03814(.I(new_n4052_), .ZN(new_n4053_));
  NOR2_X1    g03815(.A1(new_n4047_), .A2(new_n4051_), .ZN(new_n4054_));
  NOR2_X1    g03816(.A1(new_n4053_), .A2(new_n4054_), .ZN(new_n4055_));
  NOR2_X1    g03817(.A1(new_n4055_), .A2(new_n4043_), .ZN(new_n4056_));
  XOR2_X1    g03818(.A1(new_n4046_), .A2(new_n4051_), .Z(new_n4057_));
  INV_X1     g03819(.I(new_n4057_), .ZN(new_n4058_));
  AOI21_X1   g03820(.A1(new_n4043_), .A2(new_n4058_), .B(new_n4056_), .ZN(new_n4059_));
  INV_X1     g03821(.I(new_n4059_), .ZN(new_n4060_));
  XOR2_X1    g03822(.A1(new_n4032_), .A2(new_n4060_), .Z(new_n4061_));
  NOR2_X1    g03823(.A1(new_n4061_), .A2(new_n4005_), .ZN(new_n4062_));
  INV_X1     g03824(.I(new_n4005_), .ZN(new_n4063_));
  NAND3_X1   g03825(.A1(new_n4028_), .A2(new_n4031_), .A3(new_n4060_), .ZN(new_n4064_));
  NAND2_X1   g03826(.A1(new_n4032_), .A2(new_n4059_), .ZN(new_n4065_));
  AOI21_X1   g03827(.A1(new_n4065_), .A2(new_n4064_), .B(new_n4063_), .ZN(new_n4066_));
  NOR2_X1    g03828(.A1(new_n4062_), .A2(new_n4066_), .ZN(new_n4067_));
  XOR2_X1    g03829(.A1(new_n4067_), .A2(new_n4003_), .Z(new_n4068_));
  NOR2_X1    g03830(.A1(new_n4067_), .A2(new_n4003_), .ZN(new_n4069_));
  INV_X1     g03831(.I(new_n4069_), .ZN(new_n4070_));
  NAND2_X1   g03832(.A1(new_n4067_), .A2(new_n4003_), .ZN(new_n4071_));
  AOI21_X1   g03833(.A1(new_n4070_), .A2(new_n4071_), .B(new_n3951_), .ZN(new_n4072_));
  AOI21_X1   g03834(.A1(new_n4068_), .A2(new_n3951_), .B(new_n4072_), .ZN(new_n4073_));
  OAI21_X1   g03835(.A1(new_n3836_), .A2(new_n3874_), .B(new_n3872_), .ZN(new_n4074_));
  AOI21_X1   g03836(.A1(new_n3848_), .A2(new_n3863_), .B(new_n3861_), .ZN(new_n4075_));
  INV_X1     g03837(.I(new_n3895_), .ZN(new_n4076_));
  AOI21_X1   g03838(.A1(\a[17] ), .A2(\a[22] ), .B(new_n3894_), .ZN(new_n4077_));
  NOR3_X1    g03839(.A1(new_n4077_), .A2(new_n282_), .A3(new_n3423_), .ZN(new_n4078_));
  NOR2_X1    g03840(.A1(new_n4078_), .A2(new_n4076_), .ZN(new_n4079_));
  XOR2_X1    g03841(.A1(new_n4079_), .A2(new_n3885_), .Z(new_n4080_));
  NAND2_X1   g03842(.A1(new_n4080_), .A2(new_n3846_), .ZN(new_n4081_));
  NOR2_X1    g03843(.A1(new_n4079_), .A2(new_n3885_), .ZN(new_n4082_));
  NOR3_X1    g03844(.A1(new_n4078_), .A2(new_n4076_), .A3(new_n3884_), .ZN(new_n4083_));
  OAI21_X1   g03845(.A1(new_n4083_), .A2(new_n4082_), .B(new_n3845_), .ZN(new_n4084_));
  NAND2_X1   g03846(.A1(new_n4081_), .A2(new_n4084_), .ZN(new_n4085_));
  AOI21_X1   g03847(.A1(new_n3904_), .A2(new_n3902_), .B(new_n3900_), .ZN(new_n4086_));
  XNOR2_X1   g03848(.A1(new_n4086_), .A2(new_n4085_), .ZN(new_n4087_));
  NOR2_X1    g03849(.A1(new_n4087_), .A2(new_n4075_), .ZN(new_n4088_));
  INV_X1     g03850(.I(new_n4075_), .ZN(new_n4089_));
  NOR2_X1    g03851(.A1(new_n4086_), .A2(new_n4085_), .ZN(new_n4090_));
  INV_X1     g03852(.I(new_n4090_), .ZN(new_n4091_));
  NAND2_X1   g03853(.A1(new_n4086_), .A2(new_n4085_), .ZN(new_n4092_));
  AOI21_X1   g03854(.A1(new_n4091_), .A2(new_n4092_), .B(new_n4089_), .ZN(new_n4093_));
  NOR2_X1    g03855(.A1(new_n4088_), .A2(new_n4093_), .ZN(new_n4094_));
  INV_X1     g03856(.I(new_n3924_), .ZN(new_n4095_));
  OAI21_X1   g03857(.A1(new_n3879_), .A2(new_n3922_), .B(new_n4095_), .ZN(new_n4096_));
  XOR2_X1    g03858(.A1(new_n4096_), .A2(new_n4094_), .Z(new_n4097_));
  NAND2_X1   g03859(.A1(new_n4096_), .A2(new_n4094_), .ZN(new_n4098_));
  NOR2_X1    g03860(.A1(new_n3922_), .A2(new_n3879_), .ZN(new_n4099_));
  OR3_X2     g03861(.A1(new_n4099_), .A2(new_n3924_), .A3(new_n4094_), .Z(new_n4100_));
  AOI21_X1   g03862(.A1(new_n4100_), .A2(new_n4098_), .B(new_n4074_), .ZN(new_n4101_));
  AOI21_X1   g03863(.A1(new_n4074_), .A2(new_n4097_), .B(new_n4101_), .ZN(new_n4102_));
  NAND2_X1   g03864(.A1(new_n3927_), .A2(new_n3930_), .ZN(new_n4103_));
  NAND2_X1   g03865(.A1(new_n4103_), .A2(new_n3928_), .ZN(new_n4104_));
  NAND2_X1   g03866(.A1(new_n4104_), .A2(new_n4102_), .ZN(new_n4105_));
  OR2_X2     g03867(.A1(new_n4104_), .A2(new_n4102_), .Z(new_n4106_));
  AOI21_X1   g03868(.A1(new_n4106_), .A2(new_n4105_), .B(new_n4073_), .ZN(new_n4107_));
  XOR2_X1    g03869(.A1(new_n4104_), .A2(new_n4102_), .Z(new_n4108_));
  AOI21_X1   g03870(.A1(new_n4073_), .A2(new_n4108_), .B(new_n4107_), .ZN(new_n4109_));
  NOR2_X1    g03871(.A1(new_n3950_), .A2(new_n4109_), .ZN(new_n4110_));
  INV_X1     g03872(.I(new_n4110_), .ZN(new_n4111_));
  NAND2_X1   g03873(.A1(new_n3950_), .A2(new_n4109_), .ZN(new_n4112_));
  NAND2_X1   g03874(.A1(new_n4111_), .A2(new_n4112_), .ZN(new_n4113_));
  XOR2_X1    g03875(.A1(new_n3948_), .A2(new_n4113_), .Z(\asquared[41] ));
  NAND2_X1   g03876(.A1(new_n3939_), .A2(new_n4112_), .ZN(new_n4115_));
  OAI21_X1   g03877(.A1(new_n3939_), .A2(new_n4112_), .B(new_n3773_), .ZN(new_n4116_));
  NAND2_X1   g03878(.A1(new_n4116_), .A2(new_n4115_), .ZN(new_n4117_));
  NOR2_X1    g03879(.A1(new_n3771_), .A2(new_n4117_), .ZN(new_n4118_));
  INV_X1     g03880(.I(new_n4105_), .ZN(new_n4119_));
  AOI21_X1   g03881(.A1(new_n4073_), .A2(new_n4106_), .B(new_n4119_), .ZN(new_n4120_));
  INV_X1     g03882(.I(new_n4071_), .ZN(new_n4121_));
  AOI21_X1   g03883(.A1(new_n3951_), .A2(new_n4070_), .B(new_n4121_), .ZN(new_n4122_));
  NAND2_X1   g03884(.A1(new_n4100_), .A2(new_n4074_), .ZN(new_n4123_));
  NAND2_X1   g03885(.A1(new_n4123_), .A2(new_n4098_), .ZN(new_n4124_));
  INV_X1     g03886(.I(new_n4124_), .ZN(new_n4125_));
  AOI21_X1   g03887(.A1(new_n4089_), .A2(new_n4092_), .B(new_n4090_), .ZN(new_n4126_));
  AOI21_X1   g03888(.A1(new_n3959_), .A2(new_n3963_), .B(new_n3961_), .ZN(new_n4127_));
  INV_X1     g03889(.I(new_n4127_), .ZN(new_n4128_));
  INV_X1     g03890(.I(new_n4082_), .ZN(new_n4129_));
  OAI21_X1   g03891(.A1(new_n3845_), .A2(new_n4083_), .B(new_n4129_), .ZN(new_n4130_));
  OAI21_X1   g03892(.A1(new_n4043_), .A2(new_n4054_), .B(new_n4052_), .ZN(new_n4131_));
  XOR2_X1    g03893(.A1(new_n4131_), .A2(new_n4130_), .Z(new_n4132_));
  NAND2_X1   g03894(.A1(new_n4132_), .A2(new_n4128_), .ZN(new_n4133_));
  AND2_X2    g03895(.A1(new_n4131_), .A2(new_n4130_), .Z(new_n4134_));
  NOR2_X1    g03896(.A1(new_n4131_), .A2(new_n4130_), .ZN(new_n4135_));
  OAI21_X1   g03897(.A1(new_n4134_), .A2(new_n4135_), .B(new_n4127_), .ZN(new_n4136_));
  NAND2_X1   g03898(.A1(new_n4133_), .A2(new_n4136_), .ZN(new_n4137_));
  NOR2_X1    g03899(.A1(new_n873_), .A2(new_n3036_), .ZN(new_n4138_));
  NAND2_X1   g03900(.A1(\a[3] ), .A2(\a[38] ), .ZN(new_n4139_));
  XOR2_X1    g03901(.A1(new_n4138_), .A2(new_n4139_), .Z(new_n4140_));
  NAND2_X1   g03902(.A1(\a[2] ), .A2(\a[41] ), .ZN(new_n4141_));
  XOR2_X1    g03903(.A1(new_n3954_), .A2(new_n4141_), .Z(new_n4142_));
  NAND2_X1   g03904(.A1(new_n4142_), .A2(new_n4015_), .ZN(new_n4143_));
  XOR2_X1    g03905(.A1(new_n4143_), .A2(new_n1769_), .Z(new_n4144_));
  INV_X1     g03906(.I(new_n4144_), .ZN(new_n4145_));
  NAND2_X1   g03907(.A1(new_n4145_), .A2(new_n4140_), .ZN(new_n4146_));
  NOR2_X1    g03908(.A1(new_n4145_), .A2(new_n4140_), .ZN(new_n4147_));
  INV_X1     g03909(.I(new_n4147_), .ZN(new_n4148_));
  AOI21_X1   g03910(.A1(new_n4148_), .A2(new_n4146_), .B(new_n3975_), .ZN(new_n4149_));
  XOR2_X1    g03911(.A1(new_n4144_), .A2(new_n4140_), .Z(new_n4150_));
  NOR2_X1    g03912(.A1(new_n4150_), .A2(new_n3976_), .ZN(new_n4151_));
  NOR2_X1    g03913(.A1(new_n4149_), .A2(new_n4151_), .ZN(new_n4152_));
  INV_X1     g03914(.I(new_n4152_), .ZN(new_n4153_));
  XOR2_X1    g03915(.A1(new_n4137_), .A2(new_n4153_), .Z(new_n4154_));
  NOR2_X1    g03916(.A1(new_n4154_), .A2(new_n4126_), .ZN(new_n4155_));
  INV_X1     g03917(.I(new_n4126_), .ZN(new_n4156_));
  NAND3_X1   g03918(.A1(new_n4153_), .A2(new_n4133_), .A3(new_n4136_), .ZN(new_n4157_));
  NAND2_X1   g03919(.A1(new_n4137_), .A2(new_n4152_), .ZN(new_n4158_));
  AOI21_X1   g03920(.A1(new_n4158_), .A2(new_n4157_), .B(new_n4156_), .ZN(new_n4159_));
  NOR2_X1    g03921(.A1(new_n4155_), .A2(new_n4159_), .ZN(new_n4160_));
  NOR2_X1    g03922(.A1(new_n4029_), .A2(new_n4006_), .ZN(new_n4161_));
  NOR2_X1    g03923(.A1(new_n4161_), .A2(new_n4030_), .ZN(new_n4162_));
  NOR2_X1    g03924(.A1(new_n2461_), .A2(new_n3423_), .ZN(new_n4163_));
  INV_X1     g03925(.I(new_n4163_), .ZN(new_n4164_));
  NOR2_X1    g03926(.A1(new_n4164_), .A2(new_n879_), .ZN(new_n4169_));
  INV_X1     g03927(.I(new_n4169_), .ZN(new_n4170_));
  AOI21_X1   g03928(.A1(new_n3788_), .A2(new_n4021_), .B(new_n4013_), .ZN(new_n4171_));
  NOR2_X1    g03929(.A1(new_n4171_), .A2(new_n4023_), .ZN(new_n4172_));
  NOR2_X1    g03930(.A1(new_n1339_), .A2(new_n1674_), .ZN(new_n4173_));
  NAND2_X1   g03931(.A1(new_n4173_), .A2(new_n2978_), .ZN(new_n4174_));
  XOR2_X1    g03932(.A1(new_n4174_), .A2(\a[8] ), .Z(new_n4175_));
  XOR2_X1    g03933(.A1(new_n4175_), .A2(new_n2868_), .Z(new_n4176_));
  XOR2_X1    g03934(.A1(new_n4176_), .A2(new_n4172_), .Z(new_n4177_));
  INV_X1     g03935(.I(new_n4176_), .ZN(new_n4178_));
  NOR2_X1    g03936(.A1(new_n4178_), .A2(new_n4172_), .ZN(new_n4179_));
  INV_X1     g03937(.I(new_n4172_), .ZN(new_n4180_));
  NOR2_X1    g03938(.A1(new_n4180_), .A2(new_n4176_), .ZN(new_n4181_));
  OAI21_X1   g03939(.A1(new_n4179_), .A2(new_n4181_), .B(new_n4170_), .ZN(new_n4182_));
  OAI21_X1   g03940(.A1(new_n4170_), .A2(new_n4177_), .B(new_n4182_), .ZN(new_n4183_));
  INV_X1     g03941(.I(new_n3981_), .ZN(new_n4184_));
  NOR3_X1    g03942(.A1(new_n772_), .A2(new_n2765_), .A3(new_n3371_), .ZN(new_n4185_));
  NAND4_X1   g03943(.A1(new_n4185_), .A2(\a[7] ), .A3(new_n3343_), .A4(\a[34] ), .ZN(new_n4186_));
  AOI21_X1   g03944(.A1(new_n4186_), .A2(new_n4184_), .B(new_n525_), .ZN(new_n4187_));
  NOR3_X1    g03945(.A1(new_n772_), .A2(new_n2765_), .A3(new_n3371_), .ZN(new_n4188_));
  INV_X1     g03946(.I(new_n4188_), .ZN(new_n4189_));
  NOR2_X1    g03947(.A1(new_n2098_), .A2(new_n3837_), .ZN(new_n4190_));
  AOI22_X1   g03948(.A1(new_n1023_), .A2(new_n2500_), .B1(new_n4190_), .B2(new_n654_), .ZN(new_n4191_));
  NAND2_X1   g03949(.A1(\a[4] ), .A2(\a[37] ), .ZN(new_n4192_));
  INV_X1     g03950(.I(new_n4192_), .ZN(new_n4193_));
  NAND2_X1   g03951(.A1(\a[12] ), .A2(\a[29] ), .ZN(new_n4194_));
  OAI21_X1   g03952(.A1(new_n4193_), .A2(new_n4194_), .B(new_n4191_), .ZN(new_n4195_));
  XNOR2_X1   g03953(.A1(new_n4192_), .A2(new_n4194_), .ZN(new_n4196_));
  OAI21_X1   g03954(.A1(new_n650_), .A2(new_n2098_), .B(new_n4196_), .ZN(new_n4197_));
  NAND2_X1   g03955(.A1(new_n4197_), .A2(new_n4195_), .ZN(new_n4198_));
  INV_X1     g03956(.I(new_n4048_), .ZN(new_n4199_));
  INV_X1     g03957(.I(new_n1267_), .ZN(new_n4200_));
  NAND2_X1   g03958(.A1(new_n4200_), .A2(new_n1275_), .ZN(new_n4201_));
  NOR4_X1    g03959(.A1(new_n1441_), .A2(new_n2543_), .A3(new_n800_), .A4(new_n1999_), .ZN(new_n4202_));
  NAND3_X1   g03960(.A1(new_n4202_), .A2(new_n4199_), .A3(new_n4201_), .ZN(new_n4203_));
  NOR2_X1    g03961(.A1(new_n4198_), .A2(new_n4203_), .ZN(new_n4204_));
  INV_X1     g03962(.I(new_n4204_), .ZN(new_n4205_));
  NAND2_X1   g03963(.A1(new_n4198_), .A2(new_n4203_), .ZN(new_n4206_));
  AOI21_X1   g03964(.A1(new_n4205_), .A2(new_n4206_), .B(new_n4189_), .ZN(new_n4207_));
  XNOR2_X1   g03965(.A1(new_n4198_), .A2(new_n4203_), .ZN(new_n4208_));
  NOR2_X1    g03966(.A1(new_n4208_), .A2(new_n4188_), .ZN(new_n4209_));
  NOR2_X1    g03967(.A1(new_n4209_), .A2(new_n4207_), .ZN(new_n4210_));
  XNOR2_X1   g03968(.A1(new_n4183_), .A2(new_n4210_), .ZN(new_n4211_));
  NOR2_X1    g03969(.A1(new_n4211_), .A2(new_n4162_), .ZN(new_n4212_));
  INV_X1     g03970(.I(new_n4162_), .ZN(new_n4213_));
  NOR2_X1    g03971(.A1(new_n4183_), .A2(new_n4210_), .ZN(new_n4214_));
  INV_X1     g03972(.I(new_n4214_), .ZN(new_n4215_));
  NAND2_X1   g03973(.A1(new_n4183_), .A2(new_n4210_), .ZN(new_n4216_));
  AOI21_X1   g03974(.A1(new_n4215_), .A2(new_n4216_), .B(new_n4213_), .ZN(new_n4217_));
  NOR2_X1    g03975(.A1(new_n4212_), .A2(new_n4217_), .ZN(new_n4218_));
  INV_X1     g03976(.I(new_n4218_), .ZN(new_n4219_));
  XOR2_X1    g03977(.A1(new_n4160_), .A2(new_n4219_), .Z(new_n4220_));
  NOR2_X1    g03978(.A1(new_n4220_), .A2(new_n4125_), .ZN(new_n4221_));
  NOR2_X1    g03979(.A1(new_n4160_), .A2(new_n4218_), .ZN(new_n4222_));
  NOR3_X1    g03980(.A1(new_n4219_), .A2(new_n4155_), .A3(new_n4159_), .ZN(new_n4223_));
  NOR2_X1    g03981(.A1(new_n4223_), .A2(new_n4222_), .ZN(new_n4224_));
  NOR2_X1    g03982(.A1(new_n4224_), .A2(new_n4124_), .ZN(new_n4225_));
  NOR2_X1    g03983(.A1(new_n4221_), .A2(new_n4225_), .ZN(new_n4226_));
  NOR2_X1    g03984(.A1(new_n4032_), .A2(new_n4059_), .ZN(new_n4227_));
  AOI21_X1   g03985(.A1(new_n4063_), .A2(new_n4065_), .B(new_n4227_), .ZN(new_n4228_));
  NOR2_X1    g03986(.A1(new_n4000_), .A2(new_n3996_), .ZN(new_n4229_));
  NOR2_X1    g03987(.A1(new_n4229_), .A2(new_n3998_), .ZN(new_n4230_));
  INV_X1     g03988(.I(new_n3990_), .ZN(new_n4231_));
  AOI21_X1   g03989(.A1(new_n3978_), .A2(new_n4231_), .B(new_n3988_), .ZN(new_n4232_));
  INV_X1     g03990(.I(new_n4232_), .ZN(new_n4233_));
  NAND2_X1   g03991(.A1(new_n2533_), .A2(new_n787_), .ZN(new_n4234_));
  NOR2_X1    g03992(.A1(new_n2533_), .A2(new_n787_), .ZN(new_n4235_));
  NOR2_X1    g03993(.A1(\a[3] ), .A2(\a[37] ), .ZN(new_n4236_));
  AOI21_X1   g03994(.A1(new_n4234_), .A2(new_n4236_), .B(new_n4235_), .ZN(new_n4237_));
  NOR2_X1    g03995(.A1(new_n4048_), .A2(new_n4049_), .ZN(new_n4238_));
  AOI21_X1   g03996(.A1(new_n1275_), .A2(new_n2543_), .B(new_n4238_), .ZN(new_n4239_));
  INV_X1     g03997(.I(\a[40] ), .ZN(new_n4240_));
  NOR2_X1    g03998(.A1(new_n3804_), .A2(new_n4240_), .ZN(new_n4241_));
  AOI21_X1   g03999(.A1(new_n218_), .A2(new_n1675_), .B(new_n4241_), .ZN(new_n4242_));
  XOR2_X1    g04000(.A1(new_n4239_), .A2(new_n4242_), .Z(new_n4243_));
  INV_X1     g04001(.I(new_n4243_), .ZN(new_n4244_));
  INV_X1     g04002(.I(new_n4239_), .ZN(new_n4245_));
  NOR2_X1    g04003(.A1(new_n4245_), .A2(new_n4242_), .ZN(new_n4246_));
  INV_X1     g04004(.I(new_n4246_), .ZN(new_n4247_));
  NAND2_X1   g04005(.A1(new_n4245_), .A2(new_n4242_), .ZN(new_n4248_));
  AOI21_X1   g04006(.A1(new_n4247_), .A2(new_n4248_), .B(new_n4237_), .ZN(new_n4249_));
  AOI21_X1   g04007(.A1(new_n4237_), .A2(new_n4244_), .B(new_n4249_), .ZN(new_n4250_));
  OAI21_X1   g04008(.A1(new_n453_), .A2(new_n4184_), .B(new_n3980_), .ZN(new_n4251_));
  NAND2_X1   g04009(.A1(\a[1] ), .A2(\a[40] ), .ZN(new_n4252_));
  XOR2_X1    g04010(.A1(new_n4252_), .A2(\a[21] ), .Z(new_n4253_));
  XOR2_X1    g04011(.A1(new_n4039_), .A2(new_n4253_), .Z(new_n4254_));
  NOR2_X1    g04012(.A1(new_n4254_), .A2(new_n4251_), .ZN(new_n4255_));
  INV_X1     g04013(.I(new_n4039_), .ZN(new_n4256_));
  NOR2_X1    g04014(.A1(new_n4256_), .A2(new_n4253_), .ZN(new_n4257_));
  INV_X1     g04015(.I(new_n4257_), .ZN(new_n4258_));
  NAND2_X1   g04016(.A1(new_n4256_), .A2(new_n4253_), .ZN(new_n4259_));
  NAND2_X1   g04017(.A1(new_n4258_), .A2(new_n4259_), .ZN(new_n4260_));
  AOI21_X1   g04018(.A1(new_n4251_), .A2(new_n4260_), .B(new_n4255_), .ZN(new_n4261_));
  XOR2_X1    g04019(.A1(new_n4250_), .A2(new_n4261_), .Z(new_n4262_));
  NAND2_X1   g04020(.A1(new_n4262_), .A2(new_n4233_), .ZN(new_n4263_));
  NOR2_X1    g04021(.A1(new_n4250_), .A2(new_n4261_), .ZN(new_n4264_));
  NAND2_X1   g04022(.A1(new_n4250_), .A2(new_n4261_), .ZN(new_n4265_));
  INV_X1     g04023(.I(new_n4265_), .ZN(new_n4266_));
  OAI21_X1   g04024(.A1(new_n4266_), .A2(new_n4264_), .B(new_n4232_), .ZN(new_n4267_));
  NAND2_X1   g04025(.A1(new_n4263_), .A2(new_n4267_), .ZN(new_n4268_));
  INV_X1     g04026(.I(new_n4268_), .ZN(new_n4269_));
  XOR2_X1    g04027(.A1(new_n4230_), .A2(new_n4269_), .Z(new_n4270_));
  NOR3_X1    g04028(.A1(new_n4269_), .A2(new_n3998_), .A3(new_n4229_), .ZN(new_n4271_));
  NOR2_X1    g04029(.A1(new_n4230_), .A2(new_n4268_), .ZN(new_n4272_));
  OAI21_X1   g04030(.A1(new_n4272_), .A2(new_n4271_), .B(new_n4228_), .ZN(new_n4273_));
  OAI21_X1   g04031(.A1(new_n4270_), .A2(new_n4228_), .B(new_n4273_), .ZN(new_n4274_));
  XOR2_X1    g04032(.A1(new_n4226_), .A2(new_n4274_), .Z(new_n4275_));
  INV_X1     g04033(.I(new_n4274_), .ZN(new_n4276_));
  NOR2_X1    g04034(.A1(new_n4226_), .A2(new_n4276_), .ZN(new_n4277_));
  NOR3_X1    g04035(.A1(new_n4221_), .A2(new_n4225_), .A3(new_n4274_), .ZN(new_n4278_));
  OAI21_X1   g04036(.A1(new_n4277_), .A2(new_n4278_), .B(new_n4122_), .ZN(new_n4279_));
  OAI21_X1   g04037(.A1(new_n4275_), .A2(new_n4122_), .B(new_n4279_), .ZN(new_n4280_));
  INV_X1     g04038(.I(new_n4280_), .ZN(new_n4281_));
  NOR2_X1    g04039(.A1(new_n4281_), .A2(new_n4120_), .ZN(new_n4282_));
  XOR2_X1    g04040(.A1(new_n4118_), .A2(new_n4282_), .Z(new_n4283_));
  XOR2_X1    g04041(.A1(new_n4283_), .A2(new_n4110_), .Z(\asquared[42] ));
  NAND2_X1   g04042(.A1(new_n4281_), .A2(new_n4120_), .ZN(new_n4285_));
  NAND2_X1   g04043(.A1(new_n4285_), .A2(new_n4110_), .ZN(new_n4286_));
  NOR3_X1    g04044(.A1(new_n3771_), .A2(new_n4117_), .A3(new_n4286_), .ZN(new_n4287_));
  NOR2_X1    g04045(.A1(new_n4287_), .A2(new_n4282_), .ZN(new_n4288_));
  INV_X1     g04046(.I(new_n4278_), .ZN(new_n4289_));
  OAI21_X1   g04047(.A1(new_n4122_), .A2(new_n4277_), .B(new_n4289_), .ZN(new_n4290_));
  INV_X1     g04048(.I(new_n4290_), .ZN(new_n4291_));
  INV_X1     g04049(.I(new_n4222_), .ZN(new_n4292_));
  AOI21_X1   g04050(.A1(new_n4292_), .A2(new_n4124_), .B(new_n4223_), .ZN(new_n4293_));
  INV_X1     g04051(.I(new_n4293_), .ZN(new_n4294_));
  NOR2_X1    g04052(.A1(new_n4137_), .A2(new_n4152_), .ZN(new_n4295_));
  AOI21_X1   g04053(.A1(new_n4156_), .A2(new_n4158_), .B(new_n4295_), .ZN(new_n4296_));
  NAND2_X1   g04054(.A1(new_n4216_), .A2(new_n4213_), .ZN(new_n4297_));
  NAND2_X1   g04055(.A1(new_n4297_), .A2(new_n4215_), .ZN(new_n4298_));
  AOI21_X1   g04056(.A1(new_n4188_), .A2(new_n4206_), .B(new_n4204_), .ZN(new_n4299_));
  AOI21_X1   g04057(.A1(new_n4237_), .A2(new_n4248_), .B(new_n4246_), .ZN(new_n4300_));
  AOI21_X1   g04058(.A1(new_n3976_), .A2(new_n4146_), .B(new_n4147_), .ZN(new_n4301_));
  XNOR2_X1   g04059(.A1(new_n4301_), .A2(new_n4300_), .ZN(new_n4302_));
  NOR2_X1    g04060(.A1(new_n4302_), .A2(new_n4299_), .ZN(new_n4303_));
  INV_X1     g04061(.I(new_n4299_), .ZN(new_n4304_));
  NOR2_X1    g04062(.A1(new_n4301_), .A2(new_n4300_), .ZN(new_n4305_));
  INV_X1     g04063(.I(new_n4305_), .ZN(new_n4306_));
  NAND2_X1   g04064(.A1(new_n4301_), .A2(new_n4300_), .ZN(new_n4307_));
  AOI21_X1   g04065(.A1(new_n4306_), .A2(new_n4307_), .B(new_n4304_), .ZN(new_n4308_));
  NOR2_X1    g04066(.A1(new_n4303_), .A2(new_n4308_), .ZN(new_n4309_));
  XNOR2_X1   g04067(.A1(new_n4298_), .A2(new_n4309_), .ZN(new_n4310_));
  NOR2_X1    g04068(.A1(new_n4298_), .A2(new_n4309_), .ZN(new_n4311_));
  NAND2_X1   g04069(.A1(new_n4298_), .A2(new_n4309_), .ZN(new_n4312_));
  INV_X1     g04070(.I(new_n4312_), .ZN(new_n4313_));
  OAI21_X1   g04071(.A1(new_n4313_), .A2(new_n4311_), .B(new_n4296_), .ZN(new_n4314_));
  OAI21_X1   g04072(.A1(new_n4310_), .A2(new_n4296_), .B(new_n4314_), .ZN(new_n4315_));
  INV_X1     g04073(.I(new_n4272_), .ZN(new_n4316_));
  OAI21_X1   g04074(.A1(new_n4228_), .A2(new_n4271_), .B(new_n4316_), .ZN(new_n4317_));
  INV_X1     g04075(.I(new_n4317_), .ZN(new_n4318_));
  NOR2_X1    g04076(.A1(new_n4135_), .A2(new_n4127_), .ZN(new_n4319_));
  NOR2_X1    g04077(.A1(new_n4319_), .A2(new_n4134_), .ZN(new_n4320_));
  NAND2_X1   g04078(.A1(\a[39] ), .A2(\a[40] ), .ZN(new_n4321_));
  NAND2_X1   g04079(.A1(\a[16] ), .A2(\a[39] ), .ZN(new_n4322_));
  NOR3_X1    g04080(.A1(new_n4322_), .A2(new_n200_), .A3(new_n1916_), .ZN(new_n4323_));
  NAND4_X1   g04081(.A1(new_n4323_), .A2(\a[16] ), .A3(new_n2191_), .A4(\a[40] ), .ZN(new_n4324_));
  AOI21_X1   g04082(.A1(new_n4324_), .A2(new_n4321_), .B(new_n225_), .ZN(new_n4325_));
  NAND2_X1   g04083(.A1(\a[2] ), .A2(\a[40] ), .ZN(new_n4326_));
  NOR2_X1    g04084(.A1(new_n4325_), .A2(new_n4323_), .ZN(new_n4327_));
  INV_X1     g04085(.I(new_n4327_), .ZN(new_n4328_));
  NOR2_X1    g04086(.A1(new_n1916_), .A2(new_n3783_), .ZN(new_n4329_));
  AOI21_X1   g04087(.A1(\a[3] ), .A2(\a[16] ), .B(new_n4329_), .ZN(new_n4330_));
  INV_X1     g04088(.I(new_n4330_), .ZN(new_n4331_));
  OAI22_X1   g04089(.A1(new_n4328_), .A2(new_n4331_), .B1(new_n4325_), .B2(new_n4326_), .ZN(new_n4332_));
  NAND2_X1   g04090(.A1(\a[4] ), .A2(\a[28] ), .ZN(new_n4333_));
  NAND2_X1   g04091(.A1(\a[14] ), .A2(\a[38] ), .ZN(new_n4334_));
  NOR2_X1    g04092(.A1(new_n4333_), .A2(new_n4334_), .ZN(new_n4335_));
  NOR4_X1    g04093(.A1(new_n282_), .A2(new_n875_), .A3(new_n2098_), .A4(new_n3804_), .ZN(new_n4336_));
  NAND2_X1   g04094(.A1(new_n4336_), .A2(new_n4335_), .ZN(new_n4337_));
  AOI21_X1   g04095(.A1(new_n4337_), .A2(new_n2692_), .B(new_n1018_), .ZN(new_n4338_));
  NOR3_X1    g04096(.A1(new_n4338_), .A2(new_n875_), .A3(new_n2098_), .ZN(new_n4339_));
  OAI22_X1   g04097(.A1(new_n1018_), .A2(new_n2692_), .B1(new_n4333_), .B2(new_n4334_), .ZN(new_n4340_));
  INV_X1     g04098(.I(new_n4340_), .ZN(new_n4341_));
  AOI21_X1   g04099(.A1(\a[28] ), .A2(\a[38] ), .B(new_n1023_), .ZN(new_n4342_));
  NAND2_X1   g04100(.A1(new_n4341_), .A2(new_n4342_), .ZN(new_n4343_));
  INV_X1     g04101(.I(new_n4343_), .ZN(new_n4344_));
  INV_X1     g04102(.I(new_n3373_), .ZN(new_n4345_));
  NAND2_X1   g04103(.A1(new_n1441_), .A2(new_n4345_), .ZN(new_n4346_));
  NAND2_X1   g04104(.A1(new_n4199_), .A2(new_n4346_), .ZN(new_n4347_));
  NOR2_X1    g04105(.A1(new_n885_), .A2(new_n1999_), .ZN(new_n4348_));
  INV_X1     g04106(.I(new_n4348_), .ZN(new_n4349_));
  NOR4_X1    g04107(.A1(new_n4347_), .A2(new_n2331_), .A3(new_n2543_), .A4(new_n4349_), .ZN(new_n4350_));
  INV_X1     g04108(.I(new_n4350_), .ZN(new_n4351_));
  NOR3_X1    g04109(.A1(new_n4351_), .A2(new_n4339_), .A3(new_n4344_), .ZN(new_n4352_));
  NOR2_X1    g04110(.A1(new_n4339_), .A2(new_n4344_), .ZN(new_n4353_));
  NOR2_X1    g04111(.A1(new_n4353_), .A2(new_n4350_), .ZN(new_n4354_));
  NOR2_X1    g04112(.A1(new_n4354_), .A2(new_n4352_), .ZN(new_n4355_));
  NOR2_X1    g04113(.A1(new_n4355_), .A2(new_n4332_), .ZN(new_n4356_));
  XOR2_X1    g04114(.A1(new_n4353_), .A2(new_n4350_), .Z(new_n4357_));
  AOI21_X1   g04115(.A1(new_n4332_), .A2(new_n4357_), .B(new_n4356_), .ZN(new_n4358_));
  NOR2_X1    g04116(.A1(new_n2655_), .A2(new_n3393_), .ZN(new_n4359_));
  INV_X1     g04117(.I(new_n4359_), .ZN(new_n4360_));
  OAI22_X1   g04118(.A1(new_n478_), .A2(new_n4360_), .B1(new_n3967_), .B2(new_n879_), .ZN(new_n4361_));
  NOR2_X1    g04119(.A1(new_n268_), .A2(new_n3423_), .ZN(new_n4362_));
  NOR2_X1    g04120(.A1(new_n675_), .A2(new_n2655_), .ZN(new_n4363_));
  XNOR2_X1   g04121(.A1(new_n4362_), .A2(new_n4363_), .ZN(new_n4364_));
  NOR2_X1    g04122(.A1(new_n4364_), .A2(new_n4362_), .ZN(new_n4365_));
  OAI21_X1   g04123(.A1(new_n242_), .A2(new_n3393_), .B(new_n4364_), .ZN(new_n4366_));
  OAI21_X1   g04124(.A1(new_n4361_), .A2(new_n4365_), .B(new_n4366_), .ZN(new_n4367_));
  NOR2_X1    g04125(.A1(new_n2765_), .A2(new_n3371_), .ZN(new_n4368_));
  NAND2_X1   g04126(.A1(new_n3851_), .A2(new_n4368_), .ZN(new_n4369_));
  OAI21_X1   g04127(.A1(new_n391_), .A2(new_n525_), .B(new_n4369_), .ZN(new_n4370_));
  INV_X1     g04128(.I(new_n4370_), .ZN(new_n4371_));
  NOR2_X1    g04129(.A1(new_n2868_), .A2(new_n3371_), .ZN(new_n4372_));
  NOR4_X1    g04130(.A1(new_n4372_), .A2(new_n454_), .A3(new_n461_), .A4(new_n2765_), .ZN(new_n4373_));
  NAND2_X1   g04131(.A1(new_n4371_), .A2(new_n4373_), .ZN(new_n4374_));
  XNOR2_X1   g04132(.A1(new_n4367_), .A2(new_n4374_), .ZN(new_n4375_));
  NOR3_X1    g04133(.A1(new_n4375_), .A2(new_n4185_), .A3(new_n4187_), .ZN(new_n4376_));
  NOR2_X1    g04134(.A1(new_n4187_), .A2(new_n4185_), .ZN(new_n4377_));
  NOR2_X1    g04135(.A1(new_n4367_), .A2(new_n4374_), .ZN(new_n4378_));
  INV_X1     g04136(.I(new_n4378_), .ZN(new_n4379_));
  NAND2_X1   g04137(.A1(new_n4367_), .A2(new_n4374_), .ZN(new_n4380_));
  AOI21_X1   g04138(.A1(new_n4379_), .A2(new_n4380_), .B(new_n4377_), .ZN(new_n4381_));
  NOR2_X1    g04139(.A1(new_n4376_), .A2(new_n4381_), .ZN(new_n4382_));
  XOR2_X1    g04140(.A1(new_n4382_), .A2(new_n4358_), .Z(new_n4383_));
  INV_X1     g04141(.I(new_n4382_), .ZN(new_n4384_));
  NAND2_X1   g04142(.A1(new_n4384_), .A2(new_n4358_), .ZN(new_n4385_));
  INV_X1     g04143(.I(new_n4385_), .ZN(new_n4386_));
  NOR2_X1    g04144(.A1(new_n4384_), .A2(new_n4358_), .ZN(new_n4387_));
  OAI21_X1   g04145(.A1(new_n4386_), .A2(new_n4387_), .B(new_n4320_), .ZN(new_n4388_));
  OAI21_X1   g04146(.A1(new_n4320_), .A2(new_n4383_), .B(new_n4388_), .ZN(new_n4389_));
  OAI21_X1   g04147(.A1(new_n4232_), .A2(new_n4264_), .B(new_n4265_), .ZN(new_n4390_));
  INV_X1     g04148(.I(new_n4390_), .ZN(new_n4391_));
  OAI22_X1   g04149(.A1(new_n481_), .A2(new_n3967_), .B1(new_n4164_), .B2(new_n879_), .ZN(new_n4392_));
  INV_X1     g04150(.I(new_n4191_), .ZN(new_n4393_));
  OAI21_X1   g04151(.A1(new_n4192_), .A2(new_n4194_), .B(new_n4393_), .ZN(new_n4394_));
  NOR2_X1    g04152(.A1(new_n359_), .A2(new_n2868_), .ZN(new_n4395_));
  OAI21_X1   g04153(.A1(new_n2978_), .A2(new_n4173_), .B(new_n4395_), .ZN(new_n4396_));
  NAND2_X1   g04154(.A1(new_n4396_), .A2(new_n4174_), .ZN(new_n4397_));
  XOR2_X1    g04155(.A1(new_n4394_), .A2(new_n4397_), .Z(new_n4398_));
  INV_X1     g04156(.I(new_n4397_), .ZN(new_n4399_));
  NOR2_X1    g04157(.A1(new_n4394_), .A2(new_n4399_), .ZN(new_n4400_));
  NAND2_X1   g04158(.A1(new_n4394_), .A2(new_n4399_), .ZN(new_n4401_));
  INV_X1     g04159(.I(new_n4401_), .ZN(new_n4402_));
  OAI21_X1   g04160(.A1(new_n4402_), .A2(new_n4400_), .B(new_n4392_), .ZN(new_n4403_));
  OAI21_X1   g04161(.A1(new_n4392_), .A2(new_n4398_), .B(new_n4403_), .ZN(new_n4404_));
  NAND2_X1   g04162(.A1(new_n4180_), .A2(new_n4176_), .ZN(new_n4405_));
  OAI21_X1   g04163(.A1(new_n4170_), .A2(new_n4181_), .B(new_n4405_), .ZN(new_n4406_));
  NAND2_X1   g04164(.A1(new_n2328_), .A2(new_n3037_), .ZN(new_n4407_));
  NOR2_X1    g04165(.A1(new_n2328_), .A2(new_n3037_), .ZN(new_n4408_));
  NOR2_X1    g04166(.A1(\a[3] ), .A2(\a[38] ), .ZN(new_n4409_));
  AOI21_X1   g04167(.A1(new_n4407_), .A2(new_n4409_), .B(new_n4408_), .ZN(new_n4410_));
  INV_X1     g04168(.I(new_n4410_), .ZN(new_n4411_));
  AOI22_X1   g04169(.A1(new_n4199_), .A2(new_n4201_), .B1(new_n1441_), .B2(new_n2543_), .ZN(new_n4412_));
  NAND3_X1   g04170(.A1(new_n4142_), .A2(new_n1769_), .A3(new_n4015_), .ZN(new_n4413_));
  INV_X1     g04171(.I(\a[41] ), .ZN(new_n4414_));
  NOR2_X1    g04172(.A1(new_n3783_), .A2(new_n4414_), .ZN(new_n4415_));
  NAND2_X1   g04173(.A1(new_n4415_), .A2(new_n218_), .ZN(new_n4416_));
  NAND2_X1   g04174(.A1(new_n4413_), .A2(new_n4416_), .ZN(new_n4417_));
  XOR2_X1    g04175(.A1(new_n4417_), .A2(new_n4412_), .Z(new_n4418_));
  NOR2_X1    g04176(.A1(new_n4418_), .A2(new_n4411_), .ZN(new_n4419_));
  INV_X1     g04177(.I(new_n4412_), .ZN(new_n4420_));
  NOR2_X1    g04178(.A1(new_n4417_), .A2(new_n4420_), .ZN(new_n4421_));
  INV_X1     g04179(.I(new_n4421_), .ZN(new_n4422_));
  NAND2_X1   g04180(.A1(new_n4417_), .A2(new_n4420_), .ZN(new_n4423_));
  AOI21_X1   g04181(.A1(new_n4422_), .A2(new_n4423_), .B(new_n4410_), .ZN(new_n4424_));
  NOR2_X1    g04182(.A1(new_n4419_), .A2(new_n4424_), .ZN(new_n4425_));
  OR2_X2     g04183(.A1(new_n4406_), .A2(new_n4425_), .Z(new_n4426_));
  NAND2_X1   g04184(.A1(new_n4406_), .A2(new_n4425_), .ZN(new_n4427_));
  NAND2_X1   g04185(.A1(new_n4426_), .A2(new_n4427_), .ZN(new_n4428_));
  NAND2_X1   g04186(.A1(new_n4428_), .A2(new_n4404_), .ZN(new_n4429_));
  INV_X1     g04187(.I(new_n4404_), .ZN(new_n4430_));
  XOR2_X1    g04188(.A1(new_n4406_), .A2(new_n4425_), .Z(new_n4431_));
  NAND2_X1   g04189(.A1(new_n4431_), .A2(new_n4430_), .ZN(new_n4432_));
  NAND2_X1   g04190(.A1(new_n4429_), .A2(new_n4432_), .ZN(new_n4433_));
  OAI21_X1   g04191(.A1(new_n4251_), .A2(new_n4257_), .B(new_n4259_), .ZN(new_n4434_));
  INV_X1     g04192(.I(new_n4434_), .ZN(new_n4435_));
  NOR2_X1    g04193(.A1(new_n1478_), .A2(new_n4240_), .ZN(new_n4436_));
  INV_X1     g04194(.I(new_n1949_), .ZN(new_n4437_));
  NAND2_X1   g04195(.A1(\a[1] ), .A2(\a[41] ), .ZN(new_n4438_));
  INV_X1     g04196(.I(new_n4438_), .ZN(new_n4439_));
  NOR2_X1    g04197(.A1(new_n4437_), .A2(new_n4439_), .ZN(new_n4440_));
  NOR2_X1    g04198(.A1(new_n1949_), .A2(new_n4438_), .ZN(new_n4441_));
  OAI21_X1   g04199(.A1(new_n4440_), .A2(new_n4441_), .B(new_n4436_), .ZN(new_n4442_));
  XOR2_X1    g04200(.A1(new_n4442_), .A2(\a[0] ), .Z(new_n4443_));
  XOR2_X1    g04201(.A1(new_n4443_), .A2(\a[42] ), .Z(new_n4444_));
  NOR4_X1    g04202(.A1(new_n353_), .A2(new_n599_), .A3(new_n2499_), .A4(new_n3837_), .ZN(new_n4445_));
  NOR2_X1    g04203(.A1(new_n3175_), .A2(new_n1150_), .ZN(new_n4446_));
  NOR2_X1    g04204(.A1(new_n4446_), .A2(new_n4445_), .ZN(new_n4447_));
  INV_X1     g04205(.I(new_n4447_), .ZN(new_n4448_));
  NOR2_X1    g04206(.A1(new_n353_), .A2(new_n3837_), .ZN(new_n4449_));
  NOR2_X1    g04207(.A1(new_n566_), .A2(new_n2461_), .ZN(new_n4450_));
  XNOR2_X1   g04208(.A1(new_n4449_), .A2(new_n4450_), .ZN(new_n4451_));
  OAI21_X1   g04209(.A1(new_n353_), .A2(new_n3837_), .B(new_n4450_), .ZN(new_n4452_));
  NOR2_X1    g04210(.A1(new_n599_), .A2(new_n2499_), .ZN(new_n4453_));
  INV_X1     g04211(.I(new_n4453_), .ZN(new_n4454_));
  AOI22_X1   g04212(.A1(new_n4448_), .A2(new_n4452_), .B1(new_n4451_), .B2(new_n4454_), .ZN(new_n4455_));
  XOR2_X1    g04213(.A1(new_n4444_), .A2(new_n4455_), .Z(new_n4456_));
  INV_X1     g04214(.I(new_n4444_), .ZN(new_n4457_));
  NAND2_X1   g04215(.A1(new_n4457_), .A2(new_n4455_), .ZN(new_n4458_));
  INV_X1     g04216(.I(new_n4458_), .ZN(new_n4459_));
  NOR2_X1    g04217(.A1(new_n4457_), .A2(new_n4455_), .ZN(new_n4460_));
  OAI21_X1   g04218(.A1(new_n4459_), .A2(new_n4460_), .B(new_n4435_), .ZN(new_n4461_));
  OAI21_X1   g04219(.A1(new_n4456_), .A2(new_n4435_), .B(new_n4461_), .ZN(new_n4462_));
  XNOR2_X1   g04220(.A1(new_n4433_), .A2(new_n4462_), .ZN(new_n4463_));
  AND2_X2    g04221(.A1(new_n4433_), .A2(new_n4462_), .Z(new_n4464_));
  NOR2_X1    g04222(.A1(new_n4433_), .A2(new_n4462_), .ZN(new_n4465_));
  OAI21_X1   g04223(.A1(new_n4464_), .A2(new_n4465_), .B(new_n4391_), .ZN(new_n4466_));
  OAI21_X1   g04224(.A1(new_n4391_), .A2(new_n4463_), .B(new_n4466_), .ZN(new_n4467_));
  NAND2_X1   g04225(.A1(new_n4467_), .A2(new_n4389_), .ZN(new_n4468_));
  NOR2_X1    g04226(.A1(new_n4467_), .A2(new_n4389_), .ZN(new_n4469_));
  INV_X1     g04227(.I(new_n4469_), .ZN(new_n4470_));
  AOI21_X1   g04228(.A1(new_n4470_), .A2(new_n4468_), .B(new_n4318_), .ZN(new_n4471_));
  XNOR2_X1   g04229(.A1(new_n4467_), .A2(new_n4389_), .ZN(new_n4472_));
  NOR2_X1    g04230(.A1(new_n4472_), .A2(new_n4317_), .ZN(new_n4473_));
  NOR2_X1    g04231(.A1(new_n4473_), .A2(new_n4471_), .ZN(new_n4474_));
  NOR2_X1    g04232(.A1(new_n4474_), .A2(new_n4315_), .ZN(new_n4475_));
  INV_X1     g04233(.I(new_n4315_), .ZN(new_n4476_));
  INV_X1     g04234(.I(new_n4468_), .ZN(new_n4477_));
  OAI21_X1   g04235(.A1(new_n4477_), .A2(new_n4469_), .B(new_n4317_), .ZN(new_n4478_));
  OAI21_X1   g04236(.A1(new_n4317_), .A2(new_n4472_), .B(new_n4478_), .ZN(new_n4479_));
  NOR2_X1    g04237(.A1(new_n4479_), .A2(new_n4476_), .ZN(new_n4480_));
  OAI21_X1   g04238(.A1(new_n4475_), .A2(new_n4480_), .B(new_n4294_), .ZN(new_n4481_));
  NOR2_X1    g04239(.A1(new_n4474_), .A2(new_n4476_), .ZN(new_n4482_));
  NOR2_X1    g04240(.A1(new_n4479_), .A2(new_n4315_), .ZN(new_n4483_));
  OAI21_X1   g04241(.A1(new_n4482_), .A2(new_n4483_), .B(new_n4293_), .ZN(new_n4484_));
  NAND2_X1   g04242(.A1(new_n4481_), .A2(new_n4484_), .ZN(new_n4485_));
  XOR2_X1    g04243(.A1(new_n4485_), .A2(new_n4291_), .Z(new_n4486_));
  NAND2_X1   g04244(.A1(new_n4485_), .A2(new_n4290_), .ZN(new_n4487_));
  NAND3_X1   g04245(.A1(new_n4481_), .A2(new_n4484_), .A3(new_n4291_), .ZN(new_n4488_));
  NAND2_X1   g04246(.A1(new_n4487_), .A2(new_n4488_), .ZN(new_n4489_));
  NAND2_X1   g04247(.A1(new_n4288_), .A2(new_n4489_), .ZN(new_n4490_));
  OAI21_X1   g04248(.A1(new_n4288_), .A2(new_n4486_), .B(new_n4490_), .ZN(\asquared[43] ));
  OAI21_X1   g04249(.A1(new_n4287_), .A2(new_n4282_), .B(new_n4488_), .ZN(new_n4492_));
  NAND2_X1   g04250(.A1(new_n4492_), .A2(new_n4487_), .ZN(new_n4493_));
  NAND2_X1   g04251(.A1(new_n4474_), .A2(new_n4315_), .ZN(new_n4494_));
  AOI21_X1   g04252(.A1(new_n4294_), .A2(new_n4494_), .B(new_n4475_), .ZN(new_n4495_));
  INV_X1     g04253(.I(new_n4495_), .ZN(new_n4496_));
  OAI21_X1   g04254(.A1(new_n4296_), .A2(new_n4311_), .B(new_n4312_), .ZN(new_n4497_));
  INV_X1     g04255(.I(new_n4497_), .ZN(new_n4498_));
  NAND2_X1   g04256(.A1(new_n4307_), .A2(new_n4304_), .ZN(new_n4499_));
  NAND2_X1   g04257(.A1(new_n4499_), .A2(new_n4306_), .ZN(new_n4500_));
  INV_X1     g04258(.I(\a[43] ), .ZN(new_n4501_));
  NOR3_X1    g04259(.A1(new_n3954_), .A2(new_n282_), .A3(new_n4501_), .ZN(new_n4502_));
  NAND4_X1   g04260(.A1(new_n4502_), .A2(\a[40] ), .A3(new_n216_), .A4(\a[43] ), .ZN(new_n4503_));
  AOI21_X1   g04261(.A1(new_n4503_), .A2(new_n212_), .B(new_n4321_), .ZN(new_n4504_));
  NOR3_X1    g04262(.A1(new_n4504_), .A2(new_n282_), .A3(new_n3783_), .ZN(new_n4505_));
  NAND2_X1   g04263(.A1(\a[40] ), .A2(\a[43] ), .ZN(new_n4506_));
  OAI22_X1   g04264(.A1(new_n214_), .A2(new_n4506_), .B1(new_n212_), .B2(new_n4321_), .ZN(new_n4507_));
  INV_X1     g04265(.I(new_n4507_), .ZN(new_n4508_));
  AND3_X2    g04266(.A1(new_n4508_), .A2(new_n214_), .A3(new_n4506_), .Z(new_n4509_));
  NOR2_X1    g04267(.A1(new_n4505_), .A2(new_n4509_), .ZN(new_n4510_));
  INV_X1     g04268(.I(new_n4510_), .ZN(new_n4511_));
  AOI22_X1   g04269(.A1(new_n1447_), .A2(new_n2500_), .B1(new_n1718_), .B2(new_n2690_), .ZN(new_n4512_));
  NOR4_X1    g04270(.A1(new_n1719_), .A2(new_n2797_), .A3(new_n650_), .A4(new_n2499_), .ZN(new_n4513_));
  AND2_X2    g04271(.A1(new_n4512_), .A2(new_n4513_), .Z(new_n4514_));
  INV_X1     g04272(.I(new_n2679_), .ZN(new_n4515_));
  NAND2_X1   g04273(.A1(new_n2752_), .A2(new_n4515_), .ZN(new_n4516_));
  NAND2_X1   g04274(.A1(new_n4346_), .A2(new_n4516_), .ZN(new_n4517_));
  NAND2_X1   g04275(.A1(new_n2331_), .A2(new_n2277_), .ZN(new_n4518_));
  NAND2_X1   g04276(.A1(\a[18] ), .A2(\a[25] ), .ZN(new_n4519_));
  NAND2_X1   g04277(.A1(new_n1955_), .A2(new_n4519_), .ZN(new_n4520_));
  NAND4_X1   g04278(.A1(new_n4518_), .A2(\a[17] ), .A3(\a[26] ), .A4(new_n4520_), .ZN(new_n4521_));
  NOR2_X1    g04279(.A1(new_n4521_), .A2(new_n4517_), .ZN(new_n4522_));
  NAND2_X1   g04280(.A1(new_n4514_), .A2(new_n4522_), .ZN(new_n4523_));
  NOR2_X1    g04281(.A1(new_n4514_), .A2(new_n4522_), .ZN(new_n4524_));
  INV_X1     g04282(.I(new_n4524_), .ZN(new_n4525_));
  AOI21_X1   g04283(.A1(new_n4523_), .A2(new_n4525_), .B(new_n4511_), .ZN(new_n4526_));
  XNOR2_X1   g04284(.A1(new_n4514_), .A2(new_n4522_), .ZN(new_n4527_));
  NOR2_X1    g04285(.A1(new_n4527_), .A2(new_n4510_), .ZN(new_n4528_));
  NOR2_X1    g04286(.A1(new_n4526_), .A2(new_n4528_), .ZN(new_n4529_));
  INV_X1     g04287(.I(new_n3424_), .ZN(new_n4530_));
  NOR2_X1    g04288(.A1(new_n268_), .A2(new_n3393_), .ZN(new_n4531_));
  NOR2_X1    g04289(.A1(new_n4530_), .A2(new_n391_), .ZN(new_n4532_));
  NOR4_X1    g04290(.A1(new_n268_), .A2(new_n461_), .A3(new_n2868_), .A4(new_n3393_), .ZN(new_n4533_));
  NAND2_X1   g04291(.A1(new_n4532_), .A2(new_n4533_), .ZN(new_n4534_));
  AOI21_X1   g04292(.A1(new_n4534_), .A2(new_n3967_), .B(new_n392_), .ZN(new_n4535_));
  NOR2_X1    g04293(.A1(new_n4530_), .A2(new_n391_), .ZN(new_n4536_));
  NOR2_X1    g04294(.A1(new_n1711_), .A2(new_n2285_), .ZN(new_n4537_));
  INV_X1     g04295(.I(new_n1773_), .ZN(new_n4538_));
  NOR2_X1    g04296(.A1(new_n1215_), .A2(new_n2368_), .ZN(new_n4539_));
  NOR2_X1    g04297(.A1(new_n4539_), .A2(new_n4538_), .ZN(new_n4540_));
  NAND2_X1   g04298(.A1(new_n4540_), .A2(new_n4537_), .ZN(new_n4541_));
  NOR2_X1    g04299(.A1(new_n364_), .A2(new_n3371_), .ZN(new_n4542_));
  XNOR2_X1   g04300(.A1(new_n4541_), .A2(new_n4542_), .ZN(new_n4543_));
  INV_X1     g04301(.I(new_n4543_), .ZN(new_n4544_));
  NAND2_X1   g04302(.A1(\a[5] ), .A2(\a[38] ), .ZN(new_n4545_));
  NAND2_X1   g04303(.A1(\a[13] ), .A2(\a[30] ), .ZN(new_n4546_));
  NOR2_X1    g04304(.A1(new_n4545_), .A2(new_n4546_), .ZN(new_n4547_));
  XOR2_X1    g04305(.A1(new_n4547_), .A2(\a[2] ), .Z(new_n4548_));
  NAND2_X1   g04306(.A1(new_n4548_), .A2(new_n4414_), .ZN(new_n4549_));
  INV_X1     g04307(.I(new_n4549_), .ZN(new_n4550_));
  NOR2_X1    g04308(.A1(new_n4548_), .A2(new_n4414_), .ZN(new_n4551_));
  NOR2_X1    g04309(.A1(new_n4550_), .A2(new_n4551_), .ZN(new_n4552_));
  NOR2_X1    g04310(.A1(new_n4552_), .A2(new_n4544_), .ZN(new_n4553_));
  NOR3_X1    g04311(.A1(new_n4543_), .A2(new_n4550_), .A3(new_n4551_), .ZN(new_n4554_));
  OAI21_X1   g04312(.A1(new_n4553_), .A2(new_n4554_), .B(new_n4536_), .ZN(new_n4555_));
  INV_X1     g04313(.I(new_n4536_), .ZN(new_n4556_));
  XOR2_X1    g04314(.A1(new_n4552_), .A2(new_n4544_), .Z(new_n4557_));
  NAND2_X1   g04315(.A1(new_n4557_), .A2(new_n4556_), .ZN(new_n4558_));
  NAND2_X1   g04316(.A1(new_n4558_), .A2(new_n4555_), .ZN(new_n4559_));
  XOR2_X1    g04317(.A1(new_n4559_), .A2(new_n4529_), .Z(new_n4560_));
  INV_X1     g04318(.I(new_n4560_), .ZN(new_n4561_));
  OAI21_X1   g04319(.A1(new_n4526_), .A2(new_n4528_), .B(new_n4559_), .ZN(new_n4562_));
  NAND3_X1   g04320(.A1(new_n4558_), .A2(new_n4529_), .A3(new_n4555_), .ZN(new_n4563_));
  AOI21_X1   g04321(.A1(new_n4562_), .A2(new_n4563_), .B(new_n4500_), .ZN(new_n4564_));
  AOI21_X1   g04322(.A1(new_n4561_), .A2(new_n4500_), .B(new_n4564_), .ZN(new_n4565_));
  OAI21_X1   g04323(.A1(new_n4435_), .A2(new_n4460_), .B(new_n4458_), .ZN(new_n4566_));
  NAND2_X1   g04324(.A1(new_n4362_), .A2(new_n4363_), .ZN(new_n4567_));
  NAND2_X1   g04325(.A1(new_n4361_), .A2(new_n4567_), .ZN(new_n4568_));
  AOI22_X1   g04326(.A1(new_n4199_), .A2(new_n4346_), .B1(new_n2331_), .B2(new_n2543_), .ZN(new_n4569_));
  NAND2_X1   g04327(.A1(new_n4568_), .A2(new_n4569_), .ZN(new_n4570_));
  INV_X1     g04328(.I(new_n4568_), .ZN(new_n4571_));
  INV_X1     g04329(.I(new_n4569_), .ZN(new_n4572_));
  NAND2_X1   g04330(.A1(new_n4571_), .A2(new_n4572_), .ZN(new_n4573_));
  AOI21_X1   g04331(.A1(new_n4573_), .A2(new_n4570_), .B(new_n4340_), .ZN(new_n4574_));
  NOR2_X1    g04332(.A1(new_n4572_), .A2(new_n4568_), .ZN(new_n4575_));
  INV_X1     g04333(.I(new_n4575_), .ZN(new_n4576_));
  NAND2_X1   g04334(.A1(new_n4572_), .A2(new_n4568_), .ZN(new_n4577_));
  AOI21_X1   g04335(.A1(new_n4576_), .A2(new_n4577_), .B(new_n4341_), .ZN(new_n4578_));
  NOR2_X1    g04336(.A1(new_n4578_), .A2(new_n4574_), .ZN(new_n4579_));
  NAND2_X1   g04337(.A1(new_n4449_), .A2(new_n4450_), .ZN(new_n4580_));
  NAND2_X1   g04338(.A1(new_n4447_), .A2(new_n4580_), .ZN(new_n4581_));
  OR3_X2     g04339(.A1(new_n4440_), .A2(new_n4436_), .A3(new_n4441_), .Z(new_n4582_));
  NAND3_X1   g04340(.A1(new_n4582_), .A2(\a[0] ), .A3(\a[42] ), .ZN(new_n4583_));
  NAND2_X1   g04341(.A1(new_n4583_), .A2(new_n4442_), .ZN(new_n4584_));
  XOR2_X1    g04342(.A1(new_n4584_), .A2(new_n4581_), .Z(new_n4585_));
  NOR2_X1    g04343(.A1(new_n4585_), .A2(new_n4328_), .ZN(new_n4586_));
  NAND3_X1   g04344(.A1(new_n4584_), .A2(new_n4447_), .A3(new_n4580_), .ZN(new_n4587_));
  NAND3_X1   g04345(.A1(new_n4583_), .A2(new_n4442_), .A3(new_n4581_), .ZN(new_n4588_));
  AOI21_X1   g04346(.A1(new_n4587_), .A2(new_n4588_), .B(new_n4327_), .ZN(new_n4589_));
  NOR2_X1    g04347(.A1(new_n4586_), .A2(new_n4589_), .ZN(new_n4590_));
  XOR2_X1    g04348(.A1(new_n4590_), .A2(new_n4579_), .Z(new_n4591_));
  NAND2_X1   g04349(.A1(new_n4591_), .A2(new_n4566_), .ZN(new_n4592_));
  INV_X1     g04350(.I(new_n4566_), .ZN(new_n4593_));
  NOR2_X1    g04351(.A1(new_n4590_), .A2(new_n4579_), .ZN(new_n4594_));
  NAND2_X1   g04352(.A1(new_n4590_), .A2(new_n4579_), .ZN(new_n4595_));
  INV_X1     g04353(.I(new_n4595_), .ZN(new_n4596_));
  OAI21_X1   g04354(.A1(new_n4596_), .A2(new_n4594_), .B(new_n4593_), .ZN(new_n4597_));
  NAND2_X1   g04355(.A1(new_n4592_), .A2(new_n4597_), .ZN(new_n4598_));
  INV_X1     g04356(.I(new_n4400_), .ZN(new_n4599_));
  OAI21_X1   g04357(.A1(new_n4392_), .A2(new_n4402_), .B(new_n4599_), .ZN(new_n4600_));
  INV_X1     g04358(.I(new_n4600_), .ZN(new_n4601_));
  NAND4_X1   g04359(.A1(\a[6] ), .A2(\a[11] ), .A3(\a[32] ), .A4(\a[37] ), .ZN(new_n4602_));
  INV_X1     g04360(.I(new_n4602_), .ZN(new_n4603_));
  NOR3_X1    g04361(.A1(new_n1099_), .A2(new_n2655_), .A3(new_n3837_), .ZN(new_n4604_));
  NAND2_X1   g04362(.A1(new_n4603_), .A2(new_n4604_), .ZN(new_n4605_));
  AOI21_X1   g04363(.A1(new_n4605_), .A2(new_n651_), .B(new_n4184_), .ZN(new_n4606_));
  NAND2_X1   g04364(.A1(\a[12] ), .A2(\a[31] ), .ZN(new_n4607_));
  OAI21_X1   g04365(.A1(new_n4184_), .A2(new_n651_), .B(new_n4602_), .ZN(new_n4608_));
  AOI21_X1   g04366(.A1(\a[32] ), .A2(\a[37] ), .B(new_n880_), .ZN(new_n4609_));
  INV_X1     g04367(.I(new_n4609_), .ZN(new_n4610_));
  OAI22_X1   g04368(.A1(new_n4606_), .A2(new_n4607_), .B1(new_n4608_), .B2(new_n4610_), .ZN(new_n4611_));
  AOI21_X1   g04369(.A1(new_n4410_), .A2(new_n4423_), .B(new_n4421_), .ZN(new_n4612_));
  XNOR2_X1   g04370(.A1(new_n4612_), .A2(new_n4611_), .ZN(new_n4613_));
  NOR2_X1    g04371(.A1(new_n4613_), .A2(new_n4601_), .ZN(new_n4614_));
  NOR2_X1    g04372(.A1(new_n4612_), .A2(new_n4611_), .ZN(new_n4615_));
  NAND2_X1   g04373(.A1(new_n4612_), .A2(new_n4611_), .ZN(new_n4616_));
  INV_X1     g04374(.I(new_n4616_), .ZN(new_n4617_));
  NOR2_X1    g04375(.A1(new_n4617_), .A2(new_n4615_), .ZN(new_n4618_));
  NOR2_X1    g04376(.A1(new_n4618_), .A2(new_n4600_), .ZN(new_n4619_));
  NOR2_X1    g04377(.A1(new_n4619_), .A2(new_n4614_), .ZN(new_n4620_));
  INV_X1     g04378(.I(new_n4620_), .ZN(new_n4621_));
  NAND2_X1   g04379(.A1(new_n4426_), .A2(new_n4430_), .ZN(new_n4622_));
  AOI21_X1   g04380(.A1(new_n4427_), .A2(new_n4622_), .B(new_n4621_), .ZN(new_n4623_));
  NAND2_X1   g04381(.A1(new_n4622_), .A2(new_n4427_), .ZN(new_n4624_));
  NOR2_X1    g04382(.A1(new_n4624_), .A2(new_n4620_), .ZN(new_n4625_));
  OAI21_X1   g04383(.A1(new_n4623_), .A2(new_n4625_), .B(new_n4598_), .ZN(new_n4626_));
  XOR2_X1    g04384(.A1(new_n4624_), .A2(new_n4621_), .Z(new_n4627_));
  OAI21_X1   g04385(.A1(new_n4598_), .A2(new_n4627_), .B(new_n4626_), .ZN(new_n4628_));
  XOR2_X1    g04386(.A1(new_n4628_), .A2(new_n4565_), .Z(new_n4629_));
  NOR2_X1    g04387(.A1(new_n4629_), .A2(new_n4498_), .ZN(new_n4630_));
  INV_X1     g04388(.I(new_n4565_), .ZN(new_n4631_));
  NAND2_X1   g04389(.A1(new_n4628_), .A2(new_n4631_), .ZN(new_n4632_));
  OR2_X2     g04390(.A1(new_n4628_), .A2(new_n4631_), .Z(new_n4633_));
  AOI21_X1   g04391(.A1(new_n4633_), .A2(new_n4632_), .B(new_n4497_), .ZN(new_n4634_));
  NOR2_X1    g04392(.A1(new_n4630_), .A2(new_n4634_), .ZN(new_n4635_));
  AOI21_X1   g04393(.A1(new_n4317_), .A2(new_n4468_), .B(new_n4469_), .ZN(new_n4636_));
  NOR2_X1    g04394(.A1(new_n4464_), .A2(new_n4391_), .ZN(new_n4637_));
  NOR2_X1    g04395(.A1(new_n4637_), .A2(new_n4465_), .ZN(new_n4638_));
  NOR2_X1    g04396(.A1(new_n4386_), .A2(new_n4320_), .ZN(new_n4639_));
  NOR2_X1    g04397(.A1(new_n4639_), .A2(new_n4387_), .ZN(new_n4640_));
  NOR2_X1    g04398(.A1(new_n4332_), .A2(new_n4354_), .ZN(new_n4641_));
  NAND2_X1   g04399(.A1(new_n4380_), .A2(new_n4377_), .ZN(new_n4642_));
  NAND2_X1   g04400(.A1(new_n4642_), .A2(new_n4379_), .ZN(new_n4643_));
  INV_X1     g04401(.I(new_n4372_), .ZN(new_n4644_));
  OAI21_X1   g04402(.A1(new_n453_), .A2(new_n4644_), .B(new_n4370_), .ZN(new_n4645_));
  NAND2_X1   g04403(.A1(\a[1] ), .A2(\a[42] ), .ZN(new_n4646_));
  XOR2_X1    g04404(.A1(new_n4646_), .A2(\a[22] ), .Z(new_n4647_));
  XOR2_X1    g04405(.A1(new_n4647_), .A2(new_n4441_), .Z(new_n4648_));
  NOR2_X1    g04406(.A1(new_n4648_), .A2(new_n4645_), .ZN(new_n4649_));
  INV_X1     g04407(.I(new_n4441_), .ZN(new_n4650_));
  NOR2_X1    g04408(.A1(new_n4647_), .A2(new_n4650_), .ZN(new_n4651_));
  INV_X1     g04409(.I(new_n4651_), .ZN(new_n4652_));
  NAND2_X1   g04410(.A1(new_n4647_), .A2(new_n4650_), .ZN(new_n4653_));
  NAND2_X1   g04411(.A1(new_n4652_), .A2(new_n4653_), .ZN(new_n4654_));
  AOI21_X1   g04412(.A1(new_n4645_), .A2(new_n4654_), .B(new_n4649_), .ZN(new_n4655_));
  XOR2_X1    g04413(.A1(new_n4643_), .A2(new_n4655_), .Z(new_n4656_));
  OAI21_X1   g04414(.A1(new_n4352_), .A2(new_n4641_), .B(new_n4656_), .ZN(new_n4657_));
  NOR2_X1    g04415(.A1(new_n4641_), .A2(new_n4352_), .ZN(new_n4658_));
  NOR2_X1    g04416(.A1(new_n4643_), .A2(new_n4655_), .ZN(new_n4659_));
  NAND2_X1   g04417(.A1(new_n4643_), .A2(new_n4655_), .ZN(new_n4660_));
  INV_X1     g04418(.I(new_n4660_), .ZN(new_n4661_));
  OAI21_X1   g04419(.A1(new_n4661_), .A2(new_n4659_), .B(new_n4658_), .ZN(new_n4662_));
  NAND2_X1   g04420(.A1(new_n4657_), .A2(new_n4662_), .ZN(new_n4663_));
  XOR2_X1    g04421(.A1(new_n4640_), .A2(new_n4663_), .Z(new_n4664_));
  INV_X1     g04422(.I(new_n4664_), .ZN(new_n4665_));
  NOR2_X1    g04423(.A1(new_n4665_), .A2(new_n4638_), .ZN(new_n4666_));
  INV_X1     g04424(.I(new_n4640_), .ZN(new_n4667_));
  INV_X1     g04425(.I(new_n4663_), .ZN(new_n4668_));
  NOR2_X1    g04426(.A1(new_n4667_), .A2(new_n4668_), .ZN(new_n4669_));
  INV_X1     g04427(.I(new_n4669_), .ZN(new_n4670_));
  NAND2_X1   g04428(.A1(new_n4667_), .A2(new_n4668_), .ZN(new_n4671_));
  NAND2_X1   g04429(.A1(new_n4670_), .A2(new_n4671_), .ZN(new_n4672_));
  AOI21_X1   g04430(.A1(new_n4638_), .A2(new_n4672_), .B(new_n4666_), .ZN(new_n4673_));
  INV_X1     g04431(.I(new_n4673_), .ZN(new_n4674_));
  NAND2_X1   g04432(.A1(new_n4674_), .A2(new_n4636_), .ZN(new_n4675_));
  INV_X1     g04433(.I(new_n4636_), .ZN(new_n4676_));
  NAND2_X1   g04434(.A1(new_n4676_), .A2(new_n4673_), .ZN(new_n4677_));
  AOI21_X1   g04435(.A1(new_n4675_), .A2(new_n4677_), .B(new_n4635_), .ZN(new_n4678_));
  XOR2_X1    g04436(.A1(new_n4673_), .A2(new_n4636_), .Z(new_n4679_));
  NOR3_X1    g04437(.A1(new_n4679_), .A2(new_n4630_), .A3(new_n4634_), .ZN(new_n4680_));
  NOR2_X1    g04438(.A1(new_n4680_), .A2(new_n4678_), .ZN(new_n4681_));
  NOR2_X1    g04439(.A1(new_n4496_), .A2(new_n4681_), .ZN(new_n4682_));
  NOR3_X1    g04440(.A1(new_n4495_), .A2(new_n4678_), .A3(new_n4680_), .ZN(new_n4683_));
  NOR2_X1    g04441(.A1(new_n4682_), .A2(new_n4683_), .ZN(new_n4684_));
  XNOR2_X1   g04442(.A1(new_n4493_), .A2(new_n4684_), .ZN(\asquared[44] ));
  NOR2_X1    g04443(.A1(new_n4683_), .A2(new_n4485_), .ZN(new_n4686_));
  AOI21_X1   g04444(.A1(new_n4683_), .A2(new_n4485_), .B(new_n4290_), .ZN(new_n4687_));
  NOR2_X1    g04445(.A1(new_n4687_), .A2(new_n4686_), .ZN(new_n4688_));
  OAI21_X1   g04446(.A1(new_n4287_), .A2(new_n4282_), .B(new_n4688_), .ZN(new_n4689_));
  NAND2_X1   g04447(.A1(new_n4675_), .A2(new_n4635_), .ZN(new_n4690_));
  AND2_X2    g04448(.A1(new_n4690_), .A2(new_n4677_), .Z(new_n4691_));
  INV_X1     g04449(.I(new_n4691_), .ZN(new_n4692_));
  NAND2_X1   g04450(.A1(new_n4632_), .A2(new_n4497_), .ZN(new_n4693_));
  AND2_X2    g04451(.A1(new_n4693_), .A2(new_n4633_), .Z(new_n4694_));
  INV_X1     g04452(.I(new_n4694_), .ZN(new_n4695_));
  OAI21_X1   g04453(.A1(new_n4638_), .A2(new_n4669_), .B(new_n4671_), .ZN(new_n4696_));
  OAI21_X1   g04454(.A1(new_n4658_), .A2(new_n4659_), .B(new_n4660_), .ZN(new_n4697_));
  NAND2_X1   g04455(.A1(new_n2500_), .A2(new_n1143_), .ZN(new_n4698_));
  NOR2_X1    g04456(.A1(new_n200_), .A2(new_n4414_), .ZN(new_n4699_));
  XOR2_X1    g04457(.A1(new_n4698_), .A2(new_n4699_), .Z(new_n4700_));
  OAI21_X1   g04458(.A1(new_n1342_), .A2(new_n1536_), .B(new_n4516_), .ZN(new_n4701_));
  NOR2_X1    g04459(.A1(new_n1276_), .A2(new_n1916_), .ZN(new_n4702_));
  INV_X1     g04460(.I(new_n4702_), .ZN(new_n4703_));
  NOR4_X1    g04461(.A1(new_n4701_), .A2(new_n1798_), .A3(new_n2277_), .A4(new_n4703_), .ZN(new_n4704_));
  NAND2_X1   g04462(.A1(\a[33] ), .A2(\a[38] ), .ZN(new_n4705_));
  NAND2_X1   g04463(.A1(\a[37] ), .A2(\a[38] ), .ZN(new_n4706_));
  OAI22_X1   g04464(.A1(new_n478_), .A2(new_n879_), .B1(new_n4705_), .B2(new_n4706_), .ZN(new_n4707_));
  NAND4_X1   g04465(.A1(\a[7] ), .A2(\a[11] ), .A3(\a[33] ), .A4(\a[37] ), .ZN(new_n4708_));
  AOI21_X1   g04466(.A1(\a[33] ), .A2(\a[37] ), .B(new_n1009_), .ZN(new_n4709_));
  NAND4_X1   g04467(.A1(new_n4709_), .A2(new_n4708_), .A3(\a[6] ), .A4(\a[38] ), .ZN(new_n4710_));
  NOR2_X1    g04468(.A1(new_n4710_), .A2(new_n4707_), .ZN(new_n4711_));
  AND2_X2    g04469(.A1(new_n4704_), .A2(new_n4711_), .Z(new_n4712_));
  NOR2_X1    g04470(.A1(new_n4704_), .A2(new_n4711_), .ZN(new_n4713_));
  NOR2_X1    g04471(.A1(new_n4712_), .A2(new_n4713_), .ZN(new_n4714_));
  XOR2_X1    g04472(.A1(new_n4704_), .A2(new_n4711_), .Z(new_n4715_));
  NAND2_X1   g04473(.A1(new_n4715_), .A2(new_n4700_), .ZN(new_n4716_));
  OAI21_X1   g04474(.A1(new_n4700_), .A2(new_n4714_), .B(new_n4716_), .ZN(new_n4717_));
  NAND2_X1   g04475(.A1(\a[4] ), .A2(\a[40] ), .ZN(new_n4718_));
  NAND2_X1   g04476(.A1(\a[14] ), .A2(\a[30] ), .ZN(new_n4719_));
  XNOR2_X1   g04477(.A1(new_n4718_), .A2(new_n4719_), .ZN(new_n4720_));
  NAND2_X1   g04478(.A1(\a[16] ), .A2(\a[40] ), .ZN(new_n4721_));
  NOR2_X1    g04479(.A1(new_n4333_), .A2(new_n4721_), .ZN(new_n4722_));
  AOI21_X1   g04480(.A1(new_n1718_), .A2(new_n3354_), .B(new_n4722_), .ZN(new_n4723_));
  INV_X1     g04481(.I(new_n4719_), .ZN(new_n4724_));
  AOI21_X1   g04482(.A1(new_n4718_), .A2(new_n4724_), .B(new_n4723_), .ZN(new_n4725_));
  AOI21_X1   g04483(.A1(new_n2176_), .A2(new_n4720_), .B(new_n4725_), .ZN(new_n4726_));
  NOR2_X1    g04484(.A1(new_n3371_), .A2(new_n3393_), .ZN(new_n4727_));
  INV_X1     g04485(.I(new_n4727_), .ZN(new_n4728_));
  NOR2_X1    g04486(.A1(new_n3967_), .A2(new_n4728_), .ZN(new_n4729_));
  NOR2_X1    g04487(.A1(new_n4729_), .A2(new_n1720_), .ZN(new_n4730_));
  NOR2_X1    g04488(.A1(new_n359_), .A2(new_n3393_), .ZN(new_n4731_));
  NAND4_X1   g04489(.A1(new_n4730_), .A2(new_n525_), .A3(new_n3712_), .A4(new_n4731_), .ZN(new_n4732_));
  NAND2_X1   g04490(.A1(new_n3981_), .A2(new_n1220_), .ZN(new_n4733_));
  NAND2_X1   g04491(.A1(\a[5] ), .A2(\a[39] ), .ZN(new_n4734_));
  XNOR2_X1   g04492(.A1(new_n4733_), .A2(new_n4734_), .ZN(new_n4735_));
  NOR2_X1    g04493(.A1(new_n4732_), .A2(new_n4735_), .ZN(new_n4736_));
  NAND2_X1   g04494(.A1(new_n4732_), .A2(new_n4735_), .ZN(new_n4737_));
  INV_X1     g04495(.I(new_n4737_), .ZN(new_n4738_));
  OAI21_X1   g04496(.A1(new_n4738_), .A2(new_n4736_), .B(new_n4726_), .ZN(new_n4739_));
  XNOR2_X1   g04497(.A1(new_n4732_), .A2(new_n4735_), .ZN(new_n4740_));
  OAI21_X1   g04498(.A1(new_n4726_), .A2(new_n4740_), .B(new_n4739_), .ZN(new_n4741_));
  XNOR2_X1   g04499(.A1(new_n4717_), .A2(new_n4741_), .ZN(new_n4742_));
  INV_X1     g04500(.I(new_n4742_), .ZN(new_n4743_));
  NAND2_X1   g04501(.A1(new_n4717_), .A2(new_n4741_), .ZN(new_n4744_));
  NOR2_X1    g04502(.A1(new_n4717_), .A2(new_n4741_), .ZN(new_n4745_));
  INV_X1     g04503(.I(new_n4745_), .ZN(new_n4746_));
  AOI21_X1   g04504(.A1(new_n4746_), .A2(new_n4744_), .B(new_n4697_), .ZN(new_n4747_));
  AOI21_X1   g04505(.A1(new_n4697_), .A2(new_n4743_), .B(new_n4747_), .ZN(new_n4748_));
  INV_X1     g04506(.I(new_n4748_), .ZN(new_n4749_));
  NOR2_X1    g04507(.A1(new_n4617_), .A2(new_n4601_), .ZN(new_n4750_));
  NOR2_X1    g04508(.A1(new_n4535_), .A2(new_n4532_), .ZN(new_n4751_));
  INV_X1     g04509(.I(new_n4751_), .ZN(new_n4752_));
  INV_X1     g04510(.I(new_n4537_), .ZN(new_n4753_));
  NAND3_X1   g04511(.A1(new_n4753_), .A2(new_n364_), .A3(new_n3371_), .ZN(new_n4754_));
  NAND2_X1   g04512(.A1(new_n4754_), .A2(new_n4540_), .ZN(new_n4755_));
  NOR2_X1    g04513(.A1(new_n194_), .A2(new_n4501_), .ZN(new_n4756_));
  XOR2_X1    g04514(.A1(new_n4756_), .A2(new_n1706_), .Z(new_n4757_));
  XOR2_X1    g04515(.A1(new_n4755_), .A2(new_n4757_), .Z(new_n4758_));
  NOR2_X1    g04516(.A1(new_n4758_), .A2(new_n4752_), .ZN(new_n4759_));
  INV_X1     g04517(.I(new_n4755_), .ZN(new_n4760_));
  NOR2_X1    g04518(.A1(new_n4760_), .A2(new_n4757_), .ZN(new_n4761_));
  INV_X1     g04519(.I(new_n4761_), .ZN(new_n4762_));
  INV_X1     g04520(.I(new_n4757_), .ZN(new_n4763_));
  NOR2_X1    g04521(.A1(new_n4763_), .A2(new_n4755_), .ZN(new_n4764_));
  INV_X1     g04522(.I(new_n4764_), .ZN(new_n4765_));
  AOI21_X1   g04523(.A1(new_n4762_), .A2(new_n4765_), .B(new_n4751_), .ZN(new_n4766_));
  NOR2_X1    g04524(.A1(new_n4766_), .A2(new_n4759_), .ZN(new_n4767_));
  AOI21_X1   g04525(.A1(new_n1719_), .A2(new_n2797_), .B(new_n4512_), .ZN(new_n4768_));
  INV_X1     g04526(.I(\a[42] ), .ZN(new_n4769_));
  INV_X1     g04527(.I(\a[44] ), .ZN(new_n4770_));
  NOR2_X1    g04528(.A1(new_n4769_), .A2(new_n4770_), .ZN(new_n4771_));
  NOR2_X1    g04529(.A1(new_n1601_), .A2(new_n4769_), .ZN(new_n4772_));
  XOR2_X1    g04530(.A1(new_n4771_), .A2(new_n197_), .Z(new_n4773_));
  NOR2_X1    g04531(.A1(new_n4773_), .A2(new_n4608_), .ZN(new_n4774_));
  INV_X1     g04532(.I(new_n4774_), .ZN(new_n4775_));
  NAND2_X1   g04533(.A1(new_n4773_), .A2(new_n4608_), .ZN(new_n4776_));
  NAND2_X1   g04534(.A1(new_n4775_), .A2(new_n4776_), .ZN(new_n4777_));
  XNOR2_X1   g04535(.A1(new_n4773_), .A2(new_n4608_), .ZN(new_n4778_));
  NOR2_X1    g04536(.A1(new_n4778_), .A2(new_n4768_), .ZN(new_n4779_));
  AOI21_X1   g04537(.A1(new_n4768_), .A2(new_n4777_), .B(new_n4779_), .ZN(new_n4780_));
  XNOR2_X1   g04538(.A1(new_n4767_), .A2(new_n4780_), .ZN(new_n4781_));
  OAI21_X1   g04539(.A1(new_n4615_), .A2(new_n4750_), .B(new_n4781_), .ZN(new_n4782_));
  NOR2_X1    g04540(.A1(new_n4750_), .A2(new_n4615_), .ZN(new_n4783_));
  INV_X1     g04541(.I(new_n4780_), .ZN(new_n4784_));
  NAND2_X1   g04542(.A1(new_n4784_), .A2(new_n4767_), .ZN(new_n4785_));
  INV_X1     g04543(.I(new_n4785_), .ZN(new_n4786_));
  NOR2_X1    g04544(.A1(new_n4784_), .A2(new_n4767_), .ZN(new_n4787_));
  OAI21_X1   g04545(.A1(new_n4786_), .A2(new_n4787_), .B(new_n4783_), .ZN(new_n4788_));
  NAND2_X1   g04546(.A1(new_n4782_), .A2(new_n4788_), .ZN(new_n4789_));
  OAI21_X1   g04547(.A1(new_n4593_), .A2(new_n4594_), .B(new_n4595_), .ZN(new_n4790_));
  NAND2_X1   g04548(.A1(new_n4588_), .A2(new_n4327_), .ZN(new_n4791_));
  AND2_X2    g04549(.A1(new_n4791_), .A2(new_n4587_), .Z(new_n4792_));
  INV_X1     g04550(.I(new_n4792_), .ZN(new_n4793_));
  AOI21_X1   g04551(.A1(new_n4572_), .A2(new_n4568_), .B(new_n4340_), .ZN(new_n4794_));
  NOR2_X1    g04552(.A1(new_n4794_), .A2(new_n4575_), .ZN(new_n4795_));
  OAI21_X1   g04553(.A1(new_n4645_), .A2(new_n4651_), .B(new_n4653_), .ZN(new_n4796_));
  XNOR2_X1   g04554(.A1(new_n4795_), .A2(new_n4796_), .ZN(new_n4797_));
  INV_X1     g04555(.I(new_n4795_), .ZN(new_n4798_));
  NAND2_X1   g04556(.A1(new_n4798_), .A2(new_n4796_), .ZN(new_n4799_));
  INV_X1     g04557(.I(new_n4796_), .ZN(new_n4800_));
  NAND2_X1   g04558(.A1(new_n4800_), .A2(new_n4795_), .ZN(new_n4801_));
  AOI21_X1   g04559(.A1(new_n4799_), .A2(new_n4801_), .B(new_n4793_), .ZN(new_n4802_));
  AOI21_X1   g04560(.A1(new_n4793_), .A2(new_n4797_), .B(new_n4802_), .ZN(new_n4803_));
  NOR2_X1    g04561(.A1(new_n4790_), .A2(new_n4803_), .ZN(new_n4804_));
  INV_X1     g04562(.I(new_n4804_), .ZN(new_n4805_));
  NAND2_X1   g04563(.A1(new_n4790_), .A2(new_n4803_), .ZN(new_n4806_));
  NAND2_X1   g04564(.A1(new_n4805_), .A2(new_n4806_), .ZN(new_n4807_));
  NAND2_X1   g04565(.A1(new_n4807_), .A2(new_n4789_), .ZN(new_n4808_));
  XNOR2_X1   g04566(.A1(new_n4790_), .A2(new_n4803_), .ZN(new_n4809_));
  OAI21_X1   g04567(.A1(new_n4789_), .A2(new_n4809_), .B(new_n4808_), .ZN(new_n4810_));
  NAND2_X1   g04568(.A1(new_n4810_), .A2(new_n4749_), .ZN(new_n4811_));
  OR2_X2     g04569(.A1(new_n4810_), .A2(new_n4749_), .Z(new_n4812_));
  NAND2_X1   g04570(.A1(new_n4812_), .A2(new_n4811_), .ZN(new_n4813_));
  XOR2_X1    g04571(.A1(new_n4810_), .A2(new_n4748_), .Z(new_n4814_));
  NOR2_X1    g04572(.A1(new_n4814_), .A2(new_n4696_), .ZN(new_n4815_));
  AOI21_X1   g04573(.A1(new_n4696_), .A2(new_n4813_), .B(new_n4815_), .ZN(new_n4816_));
  NOR2_X1    g04574(.A1(new_n4598_), .A2(new_n4625_), .ZN(new_n4817_));
  NOR2_X1    g04575(.A1(new_n4817_), .A2(new_n4623_), .ZN(new_n4818_));
  NAND2_X1   g04576(.A1(new_n4500_), .A2(new_n4563_), .ZN(new_n4819_));
  NAND2_X1   g04577(.A1(new_n4819_), .A2(new_n4562_), .ZN(new_n4820_));
  INV_X1     g04578(.I(new_n4553_), .ZN(new_n4821_));
  OAI21_X1   g04579(.A1(new_n4556_), .A2(new_n4554_), .B(new_n4821_), .ZN(new_n4822_));
  OAI21_X1   g04580(.A1(new_n4511_), .A2(new_n4524_), .B(new_n4523_), .ZN(new_n4823_));
  AOI22_X1   g04581(.A1(new_n4346_), .A2(new_n4516_), .B1(new_n2331_), .B2(new_n2277_), .ZN(new_n4824_));
  AOI21_X1   g04582(.A1(new_n4545_), .A2(new_n4546_), .B(new_n4141_), .ZN(new_n4825_));
  NOR2_X1    g04583(.A1(new_n4825_), .A2(new_n4547_), .ZN(new_n4826_));
  INV_X1     g04584(.I(new_n4826_), .ZN(new_n4827_));
  XOR2_X1    g04585(.A1(new_n4824_), .A2(new_n4827_), .Z(new_n4828_));
  AND2_X2    g04586(.A1(new_n4824_), .A2(new_n4827_), .Z(new_n4829_));
  NOR2_X1    g04587(.A1(new_n4824_), .A2(new_n4827_), .ZN(new_n4830_));
  NOR2_X1    g04588(.A1(new_n4829_), .A2(new_n4830_), .ZN(new_n4831_));
  NOR2_X1    g04589(.A1(new_n4831_), .A2(new_n4508_), .ZN(new_n4832_));
  AOI21_X1   g04590(.A1(new_n4508_), .A2(new_n4828_), .B(new_n4832_), .ZN(new_n4833_));
  XOR2_X1    g04591(.A1(new_n4833_), .A2(new_n4823_), .Z(new_n4834_));
  NAND2_X1   g04592(.A1(new_n4834_), .A2(new_n4822_), .ZN(new_n4835_));
  OR2_X2     g04593(.A1(new_n4833_), .A2(new_n4823_), .Z(new_n4836_));
  NAND2_X1   g04594(.A1(new_n4833_), .A2(new_n4823_), .ZN(new_n4837_));
  AND2_X2    g04595(.A1(new_n4836_), .A2(new_n4837_), .Z(new_n4838_));
  OR2_X2     g04596(.A1(new_n4838_), .A2(new_n4822_), .Z(new_n4839_));
  NAND2_X1   g04597(.A1(new_n4839_), .A2(new_n4835_), .ZN(new_n4840_));
  XOR2_X1    g04598(.A1(new_n4840_), .A2(new_n4820_), .Z(new_n4841_));
  AOI21_X1   g04599(.A1(new_n4839_), .A2(new_n4835_), .B(new_n4820_), .ZN(new_n4842_));
  AOI21_X1   g04600(.A1(new_n4562_), .A2(new_n4819_), .B(new_n4840_), .ZN(new_n4843_));
  OAI21_X1   g04601(.A1(new_n4842_), .A2(new_n4843_), .B(new_n4818_), .ZN(new_n4844_));
  OAI21_X1   g04602(.A1(new_n4818_), .A2(new_n4841_), .B(new_n4844_), .ZN(new_n4845_));
  NAND2_X1   g04603(.A1(new_n4816_), .A2(new_n4845_), .ZN(new_n4846_));
  NOR2_X1    g04604(.A1(new_n4816_), .A2(new_n4845_), .ZN(new_n4847_));
  INV_X1     g04605(.I(new_n4847_), .ZN(new_n4848_));
  NAND2_X1   g04606(.A1(new_n4848_), .A2(new_n4846_), .ZN(new_n4849_));
  NAND2_X1   g04607(.A1(new_n4849_), .A2(new_n4695_), .ZN(new_n4850_));
  XOR2_X1    g04608(.A1(new_n4816_), .A2(new_n4845_), .Z(new_n4851_));
  NAND2_X1   g04609(.A1(new_n4851_), .A2(new_n4694_), .ZN(new_n4852_));
  NAND2_X1   g04610(.A1(new_n4850_), .A2(new_n4852_), .ZN(new_n4853_));
  NAND2_X1   g04611(.A1(new_n4853_), .A2(new_n4692_), .ZN(new_n4854_));
  XNOR2_X1   g04612(.A1(new_n4689_), .A2(new_n4854_), .ZN(new_n4855_));
  XNOR2_X1   g04613(.A1(new_n4855_), .A2(new_n4682_), .ZN(\asquared[45] ));
  NAND2_X1   g04614(.A1(new_n4682_), .A2(new_n4692_), .ZN(new_n4857_));
  OAI21_X1   g04615(.A1(new_n4682_), .A2(new_n4692_), .B(new_n4853_), .ZN(new_n4858_));
  OAI21_X1   g04616(.A1(new_n4689_), .A2(new_n4858_), .B(new_n4857_), .ZN(new_n4859_));
  INV_X1     g04617(.I(new_n4859_), .ZN(new_n4860_));
  NAND2_X1   g04618(.A1(new_n4846_), .A2(new_n4695_), .ZN(new_n4861_));
  NAND2_X1   g04619(.A1(new_n4861_), .A2(new_n4848_), .ZN(new_n4862_));
  INV_X1     g04620(.I(new_n4744_), .ZN(new_n4863_));
  AOI21_X1   g04621(.A1(new_n4697_), .A2(new_n4746_), .B(new_n4863_), .ZN(new_n4864_));
  OAI21_X1   g04622(.A1(new_n4789_), .A2(new_n4804_), .B(new_n4806_), .ZN(new_n4865_));
  NAND2_X1   g04623(.A1(new_n4793_), .A2(new_n4801_), .ZN(new_n4866_));
  NAND2_X1   g04624(.A1(new_n4866_), .A2(new_n4799_), .ZN(new_n4867_));
  NOR2_X1    g04625(.A1(new_n3371_), .A2(new_n3783_), .ZN(new_n4868_));
  INV_X1     g04626(.I(new_n4868_), .ZN(new_n4869_));
  NOR2_X1    g04627(.A1(new_n4869_), .A2(new_n879_), .ZN(new_n4870_));
  NAND4_X1   g04628(.A1(new_n4870_), .A2(\a[12] ), .A3(new_n3850_), .A4(\a[39] ), .ZN(new_n4871_));
  AOI21_X1   g04629(.A1(new_n4871_), .A2(new_n4644_), .B(new_n651_), .ZN(new_n4872_));
  NAND2_X1   g04630(.A1(\a[12] ), .A2(\a[33] ), .ZN(new_n4873_));
  NOR2_X1    g04631(.A1(new_n4872_), .A2(new_n4870_), .ZN(new_n4874_));
  INV_X1     g04632(.I(new_n4874_), .ZN(new_n4875_));
  NAND2_X1   g04633(.A1(new_n4869_), .A2(new_n879_), .ZN(new_n4876_));
  OAI22_X1   g04634(.A1(new_n4875_), .A2(new_n4876_), .B1(new_n4872_), .B2(new_n4873_), .ZN(new_n4877_));
  INV_X1     g04635(.I(new_n4877_), .ZN(new_n4878_));
  AOI22_X1   g04636(.A1(new_n1719_), .A2(new_n3354_), .B1(new_n2898_), .B2(new_n1143_), .ZN(new_n4879_));
  NOR2_X1    g04637(.A1(new_n875_), .A2(new_n2461_), .ZN(new_n4880_));
  NAND4_X1   g04638(.A1(new_n4879_), .A2(new_n1274_), .A3(new_n2689_), .A4(new_n4880_), .ZN(new_n4881_));
  NAND2_X1   g04639(.A1(new_n4756_), .A2(new_n1707_), .ZN(new_n4882_));
  AOI21_X1   g04640(.A1(\a[1] ), .A2(\a[44] ), .B(\a[23] ), .ZN(new_n4883_));
  NOR2_X1    g04641(.A1(new_n1684_), .A2(new_n4770_), .ZN(new_n4884_));
  NOR2_X1    g04642(.A1(new_n4884_), .A2(new_n4883_), .ZN(new_n4885_));
  NOR2_X1    g04643(.A1(new_n4885_), .A2(new_n4882_), .ZN(new_n4886_));
  XOR2_X1    g04644(.A1(new_n4886_), .A2(new_n200_), .Z(new_n4887_));
  XOR2_X1    g04645(.A1(new_n4887_), .A2(\a[42] ), .Z(new_n4888_));
  NOR2_X1    g04646(.A1(new_n4888_), .A2(new_n4881_), .ZN(new_n4889_));
  AND2_X2    g04647(.A1(new_n4888_), .A2(new_n4881_), .Z(new_n4890_));
  OAI21_X1   g04648(.A1(new_n4890_), .A2(new_n4889_), .B(new_n4878_), .ZN(new_n4891_));
  XNOR2_X1   g04649(.A1(new_n4888_), .A2(new_n4881_), .ZN(new_n4892_));
  OAI21_X1   g04650(.A1(new_n4892_), .A2(new_n4878_), .B(new_n4891_), .ZN(new_n4893_));
  NAND2_X1   g04651(.A1(new_n2500_), .A2(new_n1143_), .ZN(new_n4894_));
  NOR2_X1    g04652(.A1(new_n2500_), .A2(new_n1143_), .ZN(new_n4895_));
  NOR2_X1    g04653(.A1(\a[3] ), .A2(\a[41] ), .ZN(new_n4896_));
  AOI21_X1   g04654(.A1(new_n4894_), .A2(new_n4896_), .B(new_n4895_), .ZN(new_n4897_));
  OAI21_X1   g04655(.A1(new_n1715_), .A2(new_n2276_), .B(new_n4701_), .ZN(new_n4898_));
  AOI21_X1   g04656(.A1(new_n4772_), .A2(new_n218_), .B(new_n4771_), .ZN(new_n4899_));
  XNOR2_X1   g04657(.A1(new_n4898_), .A2(new_n4899_), .ZN(new_n4900_));
  INV_X1     g04658(.I(new_n4900_), .ZN(new_n4901_));
  NOR2_X1    g04659(.A1(new_n4898_), .A2(new_n4899_), .ZN(new_n4902_));
  INV_X1     g04660(.I(new_n4902_), .ZN(new_n4903_));
  NAND2_X1   g04661(.A1(new_n4898_), .A2(new_n4899_), .ZN(new_n4904_));
  AOI21_X1   g04662(.A1(new_n4903_), .A2(new_n4904_), .B(new_n4897_), .ZN(new_n4905_));
  AOI21_X1   g04663(.A1(new_n4901_), .A2(new_n4897_), .B(new_n4905_), .ZN(new_n4906_));
  XNOR2_X1   g04664(.A1(new_n4893_), .A2(new_n4906_), .ZN(new_n4907_));
  INV_X1     g04665(.I(new_n4907_), .ZN(new_n4908_));
  NOR2_X1    g04666(.A1(new_n4893_), .A2(new_n4906_), .ZN(new_n4909_));
  INV_X1     g04667(.I(new_n4909_), .ZN(new_n4910_));
  NAND2_X1   g04668(.A1(new_n4893_), .A2(new_n4906_), .ZN(new_n4911_));
  AOI21_X1   g04669(.A1(new_n4910_), .A2(new_n4911_), .B(new_n4867_), .ZN(new_n4912_));
  AOI21_X1   g04670(.A1(new_n4908_), .A2(new_n4867_), .B(new_n4912_), .ZN(new_n4913_));
  NOR2_X1    g04671(.A1(new_n4913_), .A2(new_n4865_), .ZN(new_n4914_));
  INV_X1     g04672(.I(new_n4914_), .ZN(new_n4915_));
  NAND2_X1   g04673(.A1(new_n4913_), .A2(new_n4865_), .ZN(new_n4916_));
  AOI21_X1   g04674(.A1(new_n4915_), .A2(new_n4916_), .B(new_n4864_), .ZN(new_n4917_));
  XOR2_X1    g04675(.A1(new_n4913_), .A2(new_n4865_), .Z(new_n4918_));
  AND2_X2    g04676(.A1(new_n4918_), .A2(new_n4864_), .Z(new_n4919_));
  NOR2_X1    g04677(.A1(new_n4919_), .A2(new_n4917_), .ZN(new_n4920_));
  NAND2_X1   g04678(.A1(new_n4811_), .A2(new_n4696_), .ZN(new_n4921_));
  NAND2_X1   g04679(.A1(new_n4921_), .A2(new_n4812_), .ZN(new_n4922_));
  NOR2_X1    g04680(.A1(new_n4818_), .A2(new_n4842_), .ZN(new_n4923_));
  NOR2_X1    g04681(.A1(new_n4923_), .A2(new_n4843_), .ZN(new_n4924_));
  OAI21_X1   g04682(.A1(new_n4783_), .A2(new_n4787_), .B(new_n4785_), .ZN(new_n4925_));
  INV_X1     g04683(.I(new_n4925_), .ZN(new_n4926_));
  AOI21_X1   g04684(.A1(new_n4762_), .A2(new_n4751_), .B(new_n4764_), .ZN(new_n4927_));
  INV_X1     g04685(.I(new_n4927_), .ZN(new_n4928_));
  NAND2_X1   g04686(.A1(new_n4776_), .A2(new_n4768_), .ZN(new_n4929_));
  NAND2_X1   g04687(.A1(new_n4929_), .A2(new_n4775_), .ZN(new_n4930_));
  NOR2_X1    g04688(.A1(new_n4830_), .A2(new_n4507_), .ZN(new_n4931_));
  NOR2_X1    g04689(.A1(new_n4931_), .A2(new_n4829_), .ZN(new_n4932_));
  XNOR2_X1   g04690(.A1(new_n4932_), .A2(new_n4930_), .ZN(new_n4933_));
  NAND2_X1   g04691(.A1(new_n4933_), .A2(new_n4928_), .ZN(new_n4934_));
  AOI21_X1   g04692(.A1(new_n4775_), .A2(new_n4929_), .B(new_n4932_), .ZN(new_n4935_));
  NOR3_X1    g04693(.A1(new_n4930_), .A2(new_n4829_), .A3(new_n4931_), .ZN(new_n4936_));
  OAI21_X1   g04694(.A1(new_n4935_), .A2(new_n4936_), .B(new_n4927_), .ZN(new_n4937_));
  NAND2_X1   g04695(.A1(new_n4934_), .A2(new_n4937_), .ZN(new_n4938_));
  INV_X1     g04696(.I(new_n4938_), .ZN(new_n4939_));
  NAND3_X1   g04697(.A1(new_n4724_), .A2(\a[4] ), .A3(\a[40] ), .ZN(new_n4940_));
  NAND2_X1   g04698(.A1(new_n4723_), .A2(new_n4940_), .ZN(new_n4941_));
  NAND2_X1   g04699(.A1(new_n3981_), .A2(new_n1220_), .ZN(new_n4942_));
  NOR2_X1    g04700(.A1(new_n3981_), .A2(new_n1220_), .ZN(new_n4943_));
  NOR2_X1    g04701(.A1(\a[5] ), .A2(\a[39] ), .ZN(new_n4944_));
  AOI21_X1   g04702(.A1(new_n4942_), .A2(new_n4944_), .B(new_n4943_), .ZN(new_n4945_));
  XNOR2_X1   g04703(.A1(new_n4941_), .A2(new_n4945_), .ZN(new_n4946_));
  NAND3_X1   g04704(.A1(new_n4946_), .A2(new_n4707_), .A3(new_n4708_), .ZN(new_n4947_));
  NAND2_X1   g04705(.A1(new_n4707_), .A2(new_n4708_), .ZN(new_n4948_));
  INV_X1     g04706(.I(new_n4945_), .ZN(new_n4949_));
  NOR2_X1    g04707(.A1(new_n4949_), .A2(new_n4941_), .ZN(new_n4950_));
  AOI21_X1   g04708(.A1(new_n4723_), .A2(new_n4940_), .B(new_n4945_), .ZN(new_n4951_));
  OAI21_X1   g04709(.A1(new_n4950_), .A2(new_n4951_), .B(new_n4948_), .ZN(new_n4952_));
  NAND2_X1   g04710(.A1(new_n4947_), .A2(new_n4952_), .ZN(new_n4953_));
  INV_X1     g04711(.I(new_n4953_), .ZN(new_n4954_));
  AOI21_X1   g04712(.A1(new_n4726_), .A2(new_n4737_), .B(new_n4736_), .ZN(new_n4955_));
  NOR2_X1    g04713(.A1(new_n4713_), .A2(new_n4700_), .ZN(new_n4956_));
  NOR2_X1    g04714(.A1(new_n4956_), .A2(new_n4712_), .ZN(new_n4957_));
  NOR2_X1    g04715(.A1(new_n4957_), .A2(new_n4955_), .ZN(new_n4958_));
  AND2_X2    g04716(.A1(new_n4957_), .A2(new_n4955_), .Z(new_n4959_));
  NOR2_X1    g04717(.A1(new_n4959_), .A2(new_n4958_), .ZN(new_n4960_));
  XOR2_X1    g04718(.A1(new_n4957_), .A2(new_n4955_), .Z(new_n4961_));
  NAND2_X1   g04719(.A1(new_n4961_), .A2(new_n4954_), .ZN(new_n4962_));
  OAI21_X1   g04720(.A1(new_n4954_), .A2(new_n4960_), .B(new_n4962_), .ZN(new_n4963_));
  XOR2_X1    g04721(.A1(new_n4963_), .A2(new_n4939_), .Z(new_n4964_));
  NOR2_X1    g04722(.A1(new_n4964_), .A2(new_n4926_), .ZN(new_n4965_));
  NAND2_X1   g04723(.A1(new_n4963_), .A2(new_n4938_), .ZN(new_n4966_));
  OR2_X2     g04724(.A1(new_n4963_), .A2(new_n4938_), .Z(new_n4967_));
  AOI21_X1   g04725(.A1(new_n4967_), .A2(new_n4966_), .B(new_n4925_), .ZN(new_n4968_));
  NOR2_X1    g04726(.A1(new_n4965_), .A2(new_n4968_), .ZN(new_n4969_));
  NAND2_X1   g04727(.A1(new_n4836_), .A2(new_n4822_), .ZN(new_n4970_));
  NAND2_X1   g04728(.A1(new_n4970_), .A2(new_n4837_), .ZN(new_n4971_));
  NOR2_X1    g04729(.A1(new_n353_), .A2(new_n599_), .ZN(new_n4972_));
  INV_X1     g04730(.I(new_n4972_), .ZN(new_n4973_));
  NOR2_X1    g04731(.A1(new_n2765_), .A2(new_n4240_), .ZN(new_n4974_));
  INV_X1     g04732(.I(new_n4974_), .ZN(new_n4975_));
  NOR2_X1    g04733(.A1(new_n4973_), .A2(new_n4975_), .ZN(new_n4976_));
  NOR4_X1    g04734(.A1(new_n353_), .A2(new_n650_), .A3(new_n2655_), .A4(new_n4240_), .ZN(new_n4977_));
  NAND2_X1   g04735(.A1(new_n4976_), .A2(new_n4977_), .ZN(new_n4978_));
  AOI21_X1   g04736(.A1(new_n4978_), .A2(new_n786_), .B(new_n4184_), .ZN(new_n4979_));
  NOR3_X1    g04737(.A1(new_n4979_), .A2(new_n650_), .A3(new_n2655_), .ZN(new_n4980_));
  OAI22_X1   g04738(.A1(new_n4973_), .A2(new_n4975_), .B1(new_n4184_), .B2(new_n786_), .ZN(new_n4981_));
  NOR3_X1    g04739(.A1(new_n4981_), .A2(new_n4972_), .A3(new_n4974_), .ZN(new_n4982_));
  NOR2_X1    g04740(.A1(new_n4980_), .A2(new_n4982_), .ZN(new_n4983_));
  AOI21_X1   g04741(.A1(new_n597_), .A2(new_n3487_), .B(new_n4730_), .ZN(new_n4984_));
  INV_X1     g04742(.I(new_n1536_), .ZN(new_n4985_));
  AOI22_X1   g04743(.A1(new_n2331_), .A2(new_n2890_), .B1(new_n2533_), .B2(new_n4985_), .ZN(new_n4986_));
  INV_X1     g04744(.I(new_n4986_), .ZN(new_n4987_));
  NOR2_X1    g04745(.A1(new_n1276_), .A2(new_n2098_), .ZN(new_n4988_));
  INV_X1     g04746(.I(new_n4988_), .ZN(new_n4989_));
  NOR4_X1    g04747(.A1(new_n4987_), .A2(new_n1798_), .A3(new_n2752_), .A4(new_n4989_), .ZN(new_n4990_));
  AND2_X2    g04748(.A1(new_n4984_), .A2(new_n4990_), .Z(new_n4991_));
  NOR2_X1    g04749(.A1(new_n4984_), .A2(new_n4990_), .ZN(new_n4992_));
  OAI21_X1   g04750(.A1(new_n4991_), .A2(new_n4992_), .B(new_n4983_), .ZN(new_n4993_));
  INV_X1     g04751(.I(new_n4983_), .ZN(new_n4994_));
  XOR2_X1    g04752(.A1(new_n4984_), .A2(new_n4990_), .Z(new_n4995_));
  NAND2_X1   g04753(.A1(new_n4994_), .A2(new_n4995_), .ZN(new_n4996_));
  NAND2_X1   g04754(.A1(new_n4996_), .A2(new_n4993_), .ZN(new_n4997_));
  INV_X1     g04755(.I(new_n4997_), .ZN(new_n4998_));
  INV_X1     g04756(.I(new_n260_), .ZN(new_n4999_));
  INV_X1     g04757(.I(new_n1142_), .ZN(new_n5000_));
  NAND3_X1   g04758(.A1(\a[41] ), .A2(\a[43] ), .A3(\a[45] ), .ZN(new_n5001_));
  NAND2_X1   g04759(.A1(new_n5000_), .A2(new_n5001_), .ZN(new_n5002_));
  NOR2_X1    g04760(.A1(new_n4414_), .A2(new_n4501_), .ZN(new_n5003_));
  INV_X1     g04761(.I(\a[45] ), .ZN(new_n5004_));
  NOR2_X1    g04762(.A1(new_n199_), .A2(new_n5004_), .ZN(new_n5005_));
  INV_X1     g04763(.I(new_n5005_), .ZN(new_n5006_));
  NOR4_X1    g04764(.A1(new_n5002_), .A2(new_n4999_), .A3(new_n5003_), .A4(new_n5006_), .ZN(new_n5007_));
  INV_X1     g04765(.I(new_n3805_), .ZN(new_n5008_));
  OAI21_X1   g04766(.A1(new_n5008_), .A2(new_n4706_), .B(new_n1779_), .ZN(new_n5009_));
  INV_X1     g04767(.I(new_n5009_), .ZN(new_n5010_));
  NOR4_X1    g04768(.A1(new_n3838_), .A2(new_n454_), .A3(new_n268_), .A4(new_n3804_), .ZN(new_n5011_));
  NAND2_X1   g04769(.A1(new_n5010_), .A2(new_n5011_), .ZN(new_n5012_));
  NOR2_X1    g04770(.A1(new_n1773_), .A2(new_n1956_), .ZN(new_n5013_));
  INV_X1     g04771(.I(new_n5013_), .ZN(new_n5014_));
  OAI21_X1   g04772(.A1(new_n1313_), .A2(new_n1691_), .B(new_n2285_), .ZN(new_n5015_));
  NOR2_X1    g04773(.A1(new_n5014_), .A2(new_n5015_), .ZN(new_n5016_));
  NOR2_X1    g04774(.A1(new_n461_), .A2(new_n3423_), .ZN(new_n5017_));
  XNOR2_X1   g04775(.A1(new_n5016_), .A2(new_n5017_), .ZN(new_n5018_));
  NOR2_X1    g04776(.A1(new_n5018_), .A2(new_n5012_), .ZN(new_n5019_));
  NAND2_X1   g04777(.A1(new_n5018_), .A2(new_n5012_), .ZN(new_n5020_));
  INV_X1     g04778(.I(new_n5020_), .ZN(new_n5021_));
  OAI21_X1   g04779(.A1(new_n5021_), .A2(new_n5019_), .B(new_n5007_), .ZN(new_n5022_));
  XNOR2_X1   g04780(.A1(new_n5018_), .A2(new_n5012_), .ZN(new_n5023_));
  OAI21_X1   g04781(.A1(new_n5007_), .A2(new_n5023_), .B(new_n5022_), .ZN(new_n5024_));
  INV_X1     g04782(.I(new_n5024_), .ZN(new_n5025_));
  NOR2_X1    g04783(.A1(new_n5025_), .A2(new_n4998_), .ZN(new_n5026_));
  NOR2_X1    g04784(.A1(new_n5024_), .A2(new_n4997_), .ZN(new_n5027_));
  OAI21_X1   g04785(.A1(new_n5026_), .A2(new_n5027_), .B(new_n4971_), .ZN(new_n5028_));
  XNOR2_X1   g04786(.A1(new_n5024_), .A2(new_n4997_), .ZN(new_n5029_));
  OAI21_X1   g04787(.A1(new_n4971_), .A2(new_n5029_), .B(new_n5028_), .ZN(new_n5030_));
  INV_X1     g04788(.I(new_n5030_), .ZN(new_n5031_));
  XOR2_X1    g04789(.A1(new_n4969_), .A2(new_n5031_), .Z(new_n5032_));
  NOR2_X1    g04790(.A1(new_n5032_), .A2(new_n4924_), .ZN(new_n5033_));
  INV_X1     g04791(.I(new_n4924_), .ZN(new_n5034_));
  NAND2_X1   g04792(.A1(new_n4969_), .A2(new_n5030_), .ZN(new_n5035_));
  OAI21_X1   g04793(.A1(new_n4965_), .A2(new_n4968_), .B(new_n5031_), .ZN(new_n5036_));
  AOI21_X1   g04794(.A1(new_n5035_), .A2(new_n5036_), .B(new_n5034_), .ZN(new_n5037_));
  NOR2_X1    g04795(.A1(new_n5037_), .A2(new_n5033_), .ZN(new_n5038_));
  NOR2_X1    g04796(.A1(new_n5038_), .A2(new_n4922_), .ZN(new_n5039_));
  AND2_X2    g04797(.A1(new_n5038_), .A2(new_n4922_), .Z(new_n5040_));
  NOR2_X1    g04798(.A1(new_n5040_), .A2(new_n5039_), .ZN(new_n5041_));
  XOR2_X1    g04799(.A1(new_n5038_), .A2(new_n4922_), .Z(new_n5042_));
  NAND2_X1   g04800(.A1(new_n5042_), .A2(new_n4920_), .ZN(new_n5043_));
  OAI21_X1   g04801(.A1(new_n4920_), .A2(new_n5041_), .B(new_n5043_), .ZN(new_n5044_));
  XNOR2_X1   g04802(.A1(new_n5044_), .A2(new_n4862_), .ZN(new_n5045_));
  NAND2_X1   g04803(.A1(new_n5044_), .A2(new_n4862_), .ZN(new_n5046_));
  NOR2_X1    g04804(.A1(new_n5044_), .A2(new_n4862_), .ZN(new_n5047_));
  INV_X1     g04805(.I(new_n5047_), .ZN(new_n5048_));
  NAND2_X1   g04806(.A1(new_n5048_), .A2(new_n5046_), .ZN(new_n5049_));
  NAND2_X1   g04807(.A1(new_n4860_), .A2(new_n5049_), .ZN(new_n5050_));
  OAI21_X1   g04808(.A1(new_n4860_), .A2(new_n5045_), .B(new_n5050_), .ZN(\asquared[46] ));
  OAI21_X1   g04809(.A1(new_n4860_), .A2(new_n5047_), .B(new_n5046_), .ZN(new_n5052_));
  NOR2_X1    g04810(.A1(new_n5039_), .A2(new_n4920_), .ZN(new_n5053_));
  NOR2_X1    g04811(.A1(new_n5053_), .A2(new_n5040_), .ZN(new_n5054_));
  NAND2_X1   g04812(.A1(new_n5034_), .A2(new_n5036_), .ZN(new_n5055_));
  NAND2_X1   g04813(.A1(new_n5055_), .A2(new_n5035_), .ZN(new_n5056_));
  NOR2_X1    g04814(.A1(new_n4963_), .A2(new_n4938_), .ZN(new_n5057_));
  AOI21_X1   g04815(.A1(new_n4925_), .A2(new_n4966_), .B(new_n5057_), .ZN(new_n5058_));
  INV_X1     g04816(.I(new_n4971_), .ZN(new_n5059_));
  INV_X1     g04817(.I(new_n5026_), .ZN(new_n5060_));
  OAI21_X1   g04818(.A1(new_n5059_), .A2(new_n5027_), .B(new_n5060_), .ZN(new_n5061_));
  NOR2_X1    g04819(.A1(new_n599_), .A2(new_n4240_), .ZN(new_n5062_));
  NAND2_X1   g04820(.A1(new_n3850_), .A2(new_n5062_), .ZN(new_n5063_));
  INV_X1     g04821(.I(new_n5063_), .ZN(new_n5064_));
  NOR4_X1    g04822(.A1(new_n242_), .A2(new_n650_), .A3(new_n2765_), .A4(new_n4240_), .ZN(new_n5065_));
  NAND2_X1   g04823(.A1(new_n5064_), .A2(new_n5065_), .ZN(new_n5066_));
  AOI21_X1   g04824(.A1(new_n5066_), .A2(new_n3852_), .B(new_n786_), .ZN(new_n5067_));
  NAND2_X1   g04825(.A1(\a[14] ), .A2(\a[32] ), .ZN(new_n5068_));
  NOR2_X1    g04826(.A1(new_n5067_), .A2(new_n5064_), .ZN(new_n5069_));
  INV_X1     g04827(.I(new_n5069_), .ZN(new_n5070_));
  AOI22_X1   g04828(.A1(\a[6] ), .A2(\a[13] ), .B1(\a[33] ), .B2(\a[40] ), .ZN(new_n5071_));
  INV_X1     g04829(.I(new_n5071_), .ZN(new_n5072_));
  OAI22_X1   g04830(.A1(new_n5070_), .A2(new_n5072_), .B1(new_n5067_), .B2(new_n5068_), .ZN(new_n5073_));
  INV_X1     g04831(.I(new_n5073_), .ZN(new_n5074_));
  NOR2_X1    g04832(.A1(new_n4951_), .A2(new_n4948_), .ZN(new_n5075_));
  NOR2_X1    g04833(.A1(new_n5075_), .A2(new_n4950_), .ZN(new_n5076_));
  NAND4_X1   g04834(.A1(\a[5] ), .A2(\a[15] ), .A3(\a[31] ), .A4(\a[41] ), .ZN(new_n5077_));
  NAND2_X1   g04835(.A1(\a[2] ), .A2(\a[44] ), .ZN(new_n5078_));
  XNOR2_X1   g04836(.A1(new_n5077_), .A2(new_n5078_), .ZN(new_n5079_));
  XOR2_X1    g04837(.A1(new_n5076_), .A2(new_n5079_), .Z(new_n5080_));
  NAND2_X1   g04838(.A1(new_n5080_), .A2(new_n5074_), .ZN(new_n5081_));
  NOR2_X1    g04839(.A1(new_n5076_), .A2(new_n5079_), .ZN(new_n5082_));
  NAND2_X1   g04840(.A1(new_n5076_), .A2(new_n5079_), .ZN(new_n5083_));
  INV_X1     g04841(.I(new_n5083_), .ZN(new_n5084_));
  OAI21_X1   g04842(.A1(new_n5084_), .A2(new_n5082_), .B(new_n5073_), .ZN(new_n5085_));
  NAND2_X1   g04843(.A1(new_n5081_), .A2(new_n5085_), .ZN(new_n5086_));
  NOR2_X1    g04844(.A1(new_n4927_), .A2(new_n4936_), .ZN(new_n5087_));
  NOR2_X1    g04845(.A1(new_n5087_), .A2(new_n4935_), .ZN(new_n5088_));
  INV_X1     g04846(.I(new_n5088_), .ZN(new_n5089_));
  AOI21_X1   g04847(.A1(new_n1275_), .A2(new_n2690_), .B(new_n4879_), .ZN(new_n5090_));
  AOI21_X1   g04848(.A1(new_n1798_), .A2(new_n2752_), .B(new_n4986_), .ZN(new_n5091_));
  XOR2_X1    g04849(.A1(new_n5090_), .A2(new_n5091_), .Z(new_n5092_));
  NAND2_X1   g04850(.A1(new_n5092_), .A2(new_n4874_), .ZN(new_n5093_));
  AND2_X2    g04851(.A1(new_n5090_), .A2(new_n5091_), .Z(new_n5094_));
  NOR2_X1    g04852(.A1(new_n5090_), .A2(new_n5091_), .ZN(new_n5095_));
  OAI21_X1   g04853(.A1(new_n5095_), .A2(new_n5094_), .B(new_n4875_), .ZN(new_n5096_));
  NAND2_X1   g04854(.A1(new_n5096_), .A2(new_n5093_), .ZN(new_n5097_));
  INV_X1     g04855(.I(new_n5097_), .ZN(new_n5098_));
  NOR2_X1    g04856(.A1(new_n5089_), .A2(new_n5098_), .ZN(new_n5099_));
  NOR2_X1    g04857(.A1(new_n5088_), .A2(new_n5097_), .ZN(new_n5100_));
  NOR2_X1    g04858(.A1(new_n5099_), .A2(new_n5100_), .ZN(new_n5101_));
  XNOR2_X1   g04859(.A1(new_n5088_), .A2(new_n5097_), .ZN(new_n5102_));
  MUX2_X1    g04860(.I0(new_n5102_), .I1(new_n5101_), .S(new_n5086_), .Z(new_n5103_));
  XNOR2_X1   g04861(.A1(new_n5103_), .A2(new_n5061_), .ZN(new_n5104_));
  NOR2_X1    g04862(.A1(new_n5103_), .A2(new_n5061_), .ZN(new_n5105_));
  NAND2_X1   g04863(.A1(new_n5103_), .A2(new_n5061_), .ZN(new_n5106_));
  INV_X1     g04864(.I(new_n5106_), .ZN(new_n5107_));
  OAI21_X1   g04865(.A1(new_n5107_), .A2(new_n5105_), .B(new_n5058_), .ZN(new_n5108_));
  OAI21_X1   g04866(.A1(new_n5058_), .A2(new_n5104_), .B(new_n5108_), .ZN(new_n5109_));
  XOR2_X1    g04867(.A1(new_n5056_), .A2(new_n5109_), .Z(new_n5110_));
  INV_X1     g04868(.I(new_n5109_), .ZN(new_n5111_));
  NOR2_X1    g04869(.A1(new_n5056_), .A2(new_n5111_), .ZN(new_n5112_));
  AOI21_X1   g04870(.A1(new_n5055_), .A2(new_n5035_), .B(new_n5109_), .ZN(new_n5113_));
  OAI21_X1   g04871(.A1(new_n5112_), .A2(new_n5113_), .B(new_n5054_), .ZN(new_n5114_));
  OAI21_X1   g04872(.A1(new_n5054_), .A2(new_n5110_), .B(new_n5114_), .ZN(new_n5115_));
  OAI21_X1   g04873(.A1(new_n4864_), .A2(new_n4914_), .B(new_n4916_), .ZN(new_n5116_));
  NOR2_X1    g04874(.A1(new_n4890_), .A2(new_n4877_), .ZN(new_n5117_));
  NOR2_X1    g04875(.A1(new_n5117_), .A2(new_n4889_), .ZN(new_n5118_));
  NOR2_X1    g04876(.A1(new_n4994_), .A2(new_n4992_), .ZN(new_n5119_));
  NOR2_X1    g04877(.A1(new_n5119_), .A2(new_n4991_), .ZN(new_n5120_));
  AND2_X2    g04878(.A1(new_n5020_), .A2(new_n5007_), .Z(new_n5121_));
  NOR2_X1    g04879(.A1(new_n5121_), .A2(new_n5019_), .ZN(new_n5122_));
  XNOR2_X1   g04880(.A1(new_n5120_), .A2(new_n5122_), .ZN(new_n5123_));
  NOR2_X1    g04881(.A1(new_n5123_), .A2(new_n5118_), .ZN(new_n5124_));
  INV_X1     g04882(.I(new_n5118_), .ZN(new_n5125_));
  NOR2_X1    g04883(.A1(new_n5120_), .A2(new_n5122_), .ZN(new_n5126_));
  INV_X1     g04884(.I(new_n5126_), .ZN(new_n5127_));
  NAND2_X1   g04885(.A1(new_n5120_), .A2(new_n5122_), .ZN(new_n5128_));
  AOI21_X1   g04886(.A1(new_n5127_), .A2(new_n5128_), .B(new_n5125_), .ZN(new_n5129_));
  NOR2_X1    g04887(.A1(new_n5129_), .A2(new_n5124_), .ZN(new_n5130_));
  NAND2_X1   g04888(.A1(new_n4910_), .A2(new_n4867_), .ZN(new_n5131_));
  NAND2_X1   g04889(.A1(new_n5131_), .A2(new_n4911_), .ZN(new_n5132_));
  AOI22_X1   g04890(.A1(new_n5000_), .A2(new_n5001_), .B1(new_n4999_), .B2(new_n5003_), .ZN(new_n5133_));
  AOI21_X1   g04891(.A1(new_n454_), .A2(new_n3838_), .B(new_n5010_), .ZN(new_n5134_));
  XNOR2_X1   g04892(.A1(new_n5134_), .A2(new_n4981_), .ZN(new_n5135_));
  INV_X1     g04893(.I(new_n5134_), .ZN(new_n5136_));
  NOR2_X1    g04894(.A1(new_n5136_), .A2(new_n4981_), .ZN(new_n5137_));
  INV_X1     g04895(.I(new_n5137_), .ZN(new_n5138_));
  NAND2_X1   g04896(.A1(new_n5136_), .A2(new_n4981_), .ZN(new_n5139_));
  AOI21_X1   g04897(.A1(new_n5138_), .A2(new_n5139_), .B(new_n5133_), .ZN(new_n5140_));
  AOI21_X1   g04898(.A1(new_n5135_), .A2(new_n5133_), .B(new_n5140_), .ZN(new_n5141_));
  AOI21_X1   g04899(.A1(new_n4897_), .A2(new_n4904_), .B(new_n4902_), .ZN(new_n5142_));
  INV_X1     g04900(.I(new_n5142_), .ZN(new_n5143_));
  NOR2_X1    g04901(.A1(\a[10] ), .A2(\a[35] ), .ZN(new_n5144_));
  AOI21_X1   g04902(.A1(new_n5014_), .A2(new_n5144_), .B(new_n5015_), .ZN(new_n5145_));
  INV_X1     g04903(.I(new_n4884_), .ZN(new_n5146_));
  NOR2_X1    g04904(.A1(new_n194_), .A2(new_n5004_), .ZN(new_n5147_));
  XOR2_X1    g04905(.A1(new_n5147_), .A2(new_n2384_), .Z(new_n5148_));
  XOR2_X1    g04906(.A1(new_n5148_), .A2(new_n5146_), .Z(new_n5149_));
  NAND2_X1   g04907(.A1(new_n5149_), .A2(new_n5145_), .ZN(new_n5150_));
  INV_X1     g04908(.I(new_n5145_), .ZN(new_n5151_));
  NOR2_X1    g04909(.A1(new_n5148_), .A2(new_n5146_), .ZN(new_n5152_));
  NAND2_X1   g04910(.A1(new_n5148_), .A2(new_n5146_), .ZN(new_n5153_));
  INV_X1     g04911(.I(new_n5153_), .ZN(new_n5154_));
  OAI21_X1   g04912(.A1(new_n5154_), .A2(new_n5152_), .B(new_n5151_), .ZN(new_n5155_));
  NAND2_X1   g04913(.A1(new_n5150_), .A2(new_n5155_), .ZN(new_n5156_));
  INV_X1     g04914(.I(new_n5156_), .ZN(new_n5157_));
  NOR2_X1    g04915(.A1(new_n5157_), .A2(new_n5143_), .ZN(new_n5158_));
  NOR2_X1    g04916(.A1(new_n5156_), .A2(new_n5142_), .ZN(new_n5159_));
  NOR2_X1    g04917(.A1(new_n5158_), .A2(new_n5159_), .ZN(new_n5160_));
  XOR2_X1    g04918(.A1(new_n5156_), .A2(new_n5143_), .Z(new_n5161_));
  MUX2_X1    g04919(.I0(new_n5160_), .I1(new_n5161_), .S(new_n5141_), .Z(new_n5162_));
  NOR2_X1    g04920(.A1(new_n5132_), .A2(new_n5162_), .ZN(new_n5163_));
  INV_X1     g04921(.I(new_n5163_), .ZN(new_n5164_));
  NAND2_X1   g04922(.A1(new_n5132_), .A2(new_n5162_), .ZN(new_n5165_));
  AOI21_X1   g04923(.A1(new_n5164_), .A2(new_n5165_), .B(new_n5130_), .ZN(new_n5166_));
  XOR2_X1    g04924(.A1(new_n5132_), .A2(new_n5162_), .Z(new_n5167_));
  NAND2_X1   g04925(.A1(new_n5167_), .A2(new_n5130_), .ZN(new_n5168_));
  INV_X1     g04926(.I(new_n5168_), .ZN(new_n5169_));
  NOR2_X1    g04927(.A1(new_n5169_), .A2(new_n5166_), .ZN(new_n5170_));
  NOR2_X1    g04928(.A1(new_n4959_), .A2(new_n4953_), .ZN(new_n5171_));
  NOR2_X1    g04929(.A1(new_n5171_), .A2(new_n4958_), .ZN(new_n5172_));
  NOR2_X1    g04930(.A1(new_n4769_), .A2(new_n4501_), .ZN(new_n5173_));
  INV_X1     g04931(.I(new_n5173_), .ZN(new_n5174_));
  INV_X1     g04932(.I(\a[46] ), .ZN(new_n5175_));
  NOR3_X1    g04933(.A1(new_n257_), .A2(new_n4769_), .A3(new_n5175_), .ZN(new_n5176_));
  NAND4_X1   g04934(.A1(new_n5176_), .A2(\a[43] ), .A3(\a[46] ), .A4(new_n216_), .ZN(new_n5177_));
  AOI21_X1   g04935(.A1(new_n5177_), .A2(new_n212_), .B(new_n5174_), .ZN(new_n5178_));
  NOR3_X1    g04936(.A1(new_n5178_), .A2(new_n200_), .A3(new_n4501_), .ZN(new_n5179_));
  NOR2_X1    g04937(.A1(new_n4769_), .A2(new_n5175_), .ZN(new_n5180_));
  NOR3_X1    g04938(.A1(new_n5178_), .A2(new_n3123_), .A3(new_n5180_), .ZN(new_n5181_));
  NOR2_X1    g04939(.A1(new_n5179_), .A2(new_n5181_), .ZN(new_n5182_));
  INV_X1     g04940(.I(new_n1236_), .ZN(new_n5183_));
  NOR2_X1    g04941(.A1(new_n3423_), .A2(new_n3837_), .ZN(new_n5184_));
  AOI22_X1   g04942(.A1(new_n597_), .A2(new_n5184_), .B1(new_n3838_), .B2(new_n5183_), .ZN(new_n5185_));
  NOR2_X1    g04943(.A1(new_n364_), .A2(new_n3837_), .ZN(new_n5186_));
  NAND4_X1   g04944(.A1(new_n5185_), .A2(new_n796_), .A3(new_n3967_), .A4(new_n5186_), .ZN(new_n5187_));
  AOI22_X1   g04945(.A1(new_n1769_), .A2(new_n2533_), .B1(new_n2890_), .B2(new_n1798_), .ZN(new_n5188_));
  INV_X1     g04946(.I(new_n5188_), .ZN(new_n5189_));
  NAND4_X1   g04947(.A1(new_n2753_), .A2(\a[19] ), .A3(\a[27] ), .A4(new_n1711_), .ZN(new_n5190_));
  NOR3_X1    g04948(.A1(new_n5187_), .A2(new_n5189_), .A3(new_n5190_), .ZN(new_n5191_));
  INV_X1     g04949(.I(new_n5187_), .ZN(new_n5192_));
  NOR2_X1    g04950(.A1(new_n5189_), .A2(new_n5190_), .ZN(new_n5193_));
  NOR2_X1    g04951(.A1(new_n5192_), .A2(new_n5193_), .ZN(new_n5194_));
  OAI21_X1   g04952(.A1(new_n5191_), .A2(new_n5194_), .B(new_n5182_), .ZN(new_n5195_));
  XOR2_X1    g04953(.A1(new_n5193_), .A2(new_n5187_), .Z(new_n5196_));
  OAI21_X1   g04954(.A1(new_n5182_), .A2(new_n5196_), .B(new_n5195_), .ZN(new_n5197_));
  NAND2_X1   g04955(.A1(new_n4885_), .A2(new_n4882_), .ZN(new_n5198_));
  NAND3_X1   g04956(.A1(new_n5198_), .A2(\a[3] ), .A3(\a[42] ), .ZN(new_n5199_));
  OAI21_X1   g04957(.A1(new_n4882_), .A2(new_n4885_), .B(new_n5199_), .ZN(new_n5200_));
  AOI22_X1   g04958(.A1(new_n4200_), .A2(new_n2898_), .B1(new_n3354_), .B2(new_n1275_), .ZN(new_n5201_));
  NOR4_X1    g04959(.A1(new_n1441_), .A2(new_n2690_), .A3(new_n800_), .A4(new_n2461_), .ZN(new_n5202_));
  NAND2_X1   g04960(.A1(new_n5201_), .A2(new_n5202_), .ZN(new_n5203_));
  INV_X1     g04961(.I(new_n3636_), .ZN(new_n5204_));
  NAND2_X1   g04962(.A1(\a[38] ), .A2(\a[39] ), .ZN(new_n5205_));
  XNOR2_X1   g04963(.A1(new_n392_), .A2(new_n5205_), .ZN(new_n5206_));
  XOR2_X1    g04964(.A1(new_n5203_), .A2(new_n5206_), .Z(new_n5207_));
  NOR2_X1    g04965(.A1(new_n5203_), .A2(new_n5206_), .ZN(new_n5208_));
  INV_X1     g04966(.I(new_n5208_), .ZN(new_n5209_));
  NAND2_X1   g04967(.A1(new_n5203_), .A2(new_n5206_), .ZN(new_n5210_));
  AOI21_X1   g04968(.A1(new_n5209_), .A2(new_n5210_), .B(new_n5200_), .ZN(new_n5211_));
  AOI21_X1   g04969(.A1(new_n5200_), .A2(new_n5207_), .B(new_n5211_), .ZN(new_n5212_));
  XNOR2_X1   g04970(.A1(new_n5197_), .A2(new_n5212_), .ZN(new_n5213_));
  NOR2_X1    g04971(.A1(new_n5213_), .A2(new_n5172_), .ZN(new_n5214_));
  INV_X1     g04972(.I(new_n5172_), .ZN(new_n5215_));
  OR2_X2     g04973(.A1(new_n5197_), .A2(new_n5212_), .Z(new_n5216_));
  NAND2_X1   g04974(.A1(new_n5197_), .A2(new_n5212_), .ZN(new_n5217_));
  AOI21_X1   g04975(.A1(new_n5216_), .A2(new_n5217_), .B(new_n5215_), .ZN(new_n5218_));
  NOR2_X1    g04976(.A1(new_n5218_), .A2(new_n5214_), .ZN(new_n5219_));
  XOR2_X1    g04977(.A1(new_n5170_), .A2(new_n5219_), .Z(new_n5220_));
  OAI22_X1   g04978(.A1(new_n5169_), .A2(new_n5166_), .B1(new_n5214_), .B2(new_n5218_), .ZN(new_n5221_));
  NAND2_X1   g04979(.A1(new_n5170_), .A2(new_n5219_), .ZN(new_n5222_));
  NAND2_X1   g04980(.A1(new_n5222_), .A2(new_n5221_), .ZN(new_n5223_));
  MUX2_X1    g04981(.I0(new_n5223_), .I1(new_n5220_), .S(new_n5116_), .Z(new_n5224_));
  XOR2_X1    g04982(.A1(new_n5115_), .A2(new_n5224_), .Z(new_n5225_));
  NAND2_X1   g04983(.A1(new_n5052_), .A2(new_n5225_), .ZN(new_n5226_));
  XOR2_X1    g04984(.A1(new_n5115_), .A2(new_n5224_), .Z(new_n5227_));
  OAI21_X1   g04985(.A1(new_n5052_), .A2(new_n5227_), .B(new_n5226_), .ZN(\asquared[47] ));
  NAND2_X1   g04986(.A1(new_n5115_), .A2(new_n5224_), .ZN(new_n5229_));
  NOR2_X1    g04987(.A1(new_n5115_), .A2(new_n5224_), .ZN(new_n5230_));
  NOR2_X1    g04988(.A1(new_n5230_), .A2(new_n5044_), .ZN(new_n5231_));
  AOI21_X1   g04989(.A1(new_n5230_), .A2(new_n5044_), .B(new_n4862_), .ZN(new_n5232_));
  NOR2_X1    g04990(.A1(new_n5232_), .A2(new_n5231_), .ZN(new_n5233_));
  NAND2_X1   g04991(.A1(new_n4859_), .A2(new_n5233_), .ZN(new_n5234_));
  NOR2_X1    g04992(.A1(new_n5054_), .A2(new_n5112_), .ZN(new_n5235_));
  NOR2_X1    g04993(.A1(new_n5235_), .A2(new_n5113_), .ZN(new_n5236_));
  OAI21_X1   g04994(.A1(new_n5058_), .A2(new_n5105_), .B(new_n5106_), .ZN(new_n5237_));
  NAND2_X1   g04995(.A1(new_n5164_), .A2(new_n5130_), .ZN(new_n5238_));
  NAND2_X1   g04996(.A1(new_n5238_), .A2(new_n5165_), .ZN(new_n5239_));
  AOI21_X1   g04997(.A1(new_n5074_), .A2(new_n5083_), .B(new_n5082_), .ZN(new_n5240_));
  NOR3_X1    g04998(.A1(new_n5194_), .A2(new_n5179_), .A3(new_n5181_), .ZN(new_n5241_));
  NOR2_X1    g04999(.A1(new_n5241_), .A2(new_n5191_), .ZN(new_n5242_));
  NOR2_X1    g05000(.A1(new_n5178_), .A2(new_n5176_), .ZN(new_n5243_));
  AOI21_X1   g05001(.A1(new_n2978_), .A2(new_n2752_), .B(new_n5188_), .ZN(new_n5244_));
  NOR2_X1    g05002(.A1(new_n2655_), .A2(new_n4414_), .ZN(new_n5245_));
  NOR2_X1    g05003(.A1(new_n353_), .A2(new_n875_), .ZN(new_n5246_));
  NOR4_X1    g05004(.A1(new_n353_), .A2(new_n875_), .A3(new_n2655_), .A4(new_n4414_), .ZN(new_n5247_));
  NAND2_X1   g05005(.A1(new_n201_), .A2(new_n4770_), .ZN(new_n5248_));
  OAI22_X1   g05006(.A1(new_n5247_), .A2(new_n5248_), .B1(new_n5245_), .B2(new_n5246_), .ZN(new_n5249_));
  XNOR2_X1   g05007(.A1(new_n5244_), .A2(new_n5249_), .ZN(new_n5250_));
  INV_X1     g05008(.I(new_n5244_), .ZN(new_n5251_));
  NOR2_X1    g05009(.A1(new_n5251_), .A2(new_n5249_), .ZN(new_n5252_));
  INV_X1     g05010(.I(new_n5252_), .ZN(new_n5253_));
  NAND2_X1   g05011(.A1(new_n5251_), .A2(new_n5249_), .ZN(new_n5254_));
  AOI21_X1   g05012(.A1(new_n5253_), .A2(new_n5254_), .B(new_n5243_), .ZN(new_n5255_));
  AOI21_X1   g05013(.A1(new_n5243_), .A2(new_n5250_), .B(new_n5255_), .ZN(new_n5256_));
  XOR2_X1    g05014(.A1(new_n5256_), .A2(new_n5242_), .Z(new_n5257_));
  NOR2_X1    g05015(.A1(new_n5257_), .A2(new_n5240_), .ZN(new_n5258_));
  INV_X1     g05016(.I(new_n5240_), .ZN(new_n5259_));
  INV_X1     g05017(.I(new_n5242_), .ZN(new_n5260_));
  NOR2_X1    g05018(.A1(new_n5256_), .A2(new_n5260_), .ZN(new_n5261_));
  INV_X1     g05019(.I(new_n5261_), .ZN(new_n5262_));
  NAND2_X1   g05020(.A1(new_n5256_), .A2(new_n5260_), .ZN(new_n5263_));
  AOI21_X1   g05021(.A1(new_n5262_), .A2(new_n5263_), .B(new_n5259_), .ZN(new_n5264_));
  NOR2_X1    g05022(.A1(new_n5258_), .A2(new_n5264_), .ZN(new_n5265_));
  INV_X1     g05023(.I(new_n5100_), .ZN(new_n5266_));
  OAI21_X1   g05024(.A1(new_n5086_), .A2(new_n5099_), .B(new_n5266_), .ZN(new_n5267_));
  NAND2_X1   g05025(.A1(new_n5215_), .A2(new_n5216_), .ZN(new_n5268_));
  NAND2_X1   g05026(.A1(new_n5268_), .A2(new_n5217_), .ZN(new_n5269_));
  NAND2_X1   g05027(.A1(new_n5269_), .A2(new_n5267_), .ZN(new_n5270_));
  NOR2_X1    g05028(.A1(new_n5269_), .A2(new_n5267_), .ZN(new_n5271_));
  INV_X1     g05029(.I(new_n5271_), .ZN(new_n5272_));
  AOI21_X1   g05030(.A1(new_n5272_), .A2(new_n5270_), .B(new_n5265_), .ZN(new_n5273_));
  INV_X1     g05031(.I(new_n5265_), .ZN(new_n5274_));
  XNOR2_X1   g05032(.A1(new_n5269_), .A2(new_n5267_), .ZN(new_n5275_));
  NOR2_X1    g05033(.A1(new_n5275_), .A2(new_n5274_), .ZN(new_n5276_));
  NOR2_X1    g05034(.A1(new_n5276_), .A2(new_n5273_), .ZN(new_n5277_));
  NOR2_X1    g05035(.A1(new_n5239_), .A2(new_n5277_), .ZN(new_n5278_));
  NAND2_X1   g05036(.A1(new_n5239_), .A2(new_n5277_), .ZN(new_n5279_));
  INV_X1     g05037(.I(new_n5279_), .ZN(new_n5280_));
  OAI21_X1   g05038(.A1(new_n5280_), .A2(new_n5278_), .B(new_n5237_), .ZN(new_n5281_));
  XNOR2_X1   g05039(.A1(new_n5239_), .A2(new_n5277_), .ZN(new_n5282_));
  OAI21_X1   g05040(.A1(new_n5237_), .A2(new_n5282_), .B(new_n5281_), .ZN(new_n5283_));
  INV_X1     g05041(.I(new_n5283_), .ZN(new_n5284_));
  NAND2_X1   g05042(.A1(new_n5221_), .A2(new_n5116_), .ZN(new_n5285_));
  NAND2_X1   g05043(.A1(new_n5285_), .A2(new_n5222_), .ZN(new_n5286_));
  AOI21_X1   g05044(.A1(new_n5125_), .A2(new_n5128_), .B(new_n5126_), .ZN(new_n5287_));
  NOR2_X1    g05045(.A1(new_n4875_), .A2(new_n5095_), .ZN(new_n5288_));
  NOR2_X1    g05046(.A1(new_n5288_), .A2(new_n5094_), .ZN(new_n5289_));
  OAI21_X1   g05047(.A1(new_n5151_), .A2(new_n5152_), .B(new_n5153_), .ZN(new_n5290_));
  NOR2_X1    g05048(.A1(new_n566_), .A2(new_n4240_), .ZN(new_n5291_));
  INV_X1     g05049(.I(new_n5291_), .ZN(new_n5292_));
  NOR3_X1    g05050(.A1(new_n5292_), .A2(new_n268_), .A3(new_n3423_), .ZN(new_n5293_));
  NOR4_X1    g05051(.A1(new_n268_), .A2(new_n566_), .A3(new_n3423_), .A4(new_n4240_), .ZN(new_n5297_));
  INV_X1     g05052(.I(new_n5297_), .ZN(new_n5298_));
  XOR2_X1    g05053(.A1(new_n5290_), .A2(new_n5298_), .Z(new_n5299_));
  NOR2_X1    g05054(.A1(new_n5299_), .A2(new_n5289_), .ZN(new_n5300_));
  INV_X1     g05055(.I(new_n5289_), .ZN(new_n5301_));
  INV_X1     g05056(.I(new_n5290_), .ZN(new_n5302_));
  NOR2_X1    g05057(.A1(new_n5302_), .A2(new_n5298_), .ZN(new_n5303_));
  NOR2_X1    g05058(.A1(new_n5290_), .A2(new_n5297_), .ZN(new_n5304_));
  NOR2_X1    g05059(.A1(new_n5303_), .A2(new_n5304_), .ZN(new_n5305_));
  NOR2_X1    g05060(.A1(new_n5301_), .A2(new_n5305_), .ZN(new_n5306_));
  NOR2_X1    g05061(.A1(new_n5306_), .A2(new_n5300_), .ZN(new_n5307_));
  INV_X1     g05062(.I(new_n5307_), .ZN(new_n5308_));
  INV_X1     g05063(.I(new_n5159_), .ZN(new_n5309_));
  OAI21_X1   g05064(.A1(new_n5143_), .A2(new_n5157_), .B(new_n5141_), .ZN(new_n5310_));
  NAND2_X1   g05065(.A1(new_n5310_), .A2(new_n5309_), .ZN(new_n5311_));
  XOR2_X1    g05066(.A1(new_n5311_), .A2(new_n5308_), .Z(new_n5312_));
  NOR2_X1    g05067(.A1(new_n5312_), .A2(new_n5287_), .ZN(new_n5313_));
  INV_X1     g05068(.I(new_n5287_), .ZN(new_n5314_));
  INV_X1     g05069(.I(new_n5311_), .ZN(new_n5315_));
  NOR2_X1    g05070(.A1(new_n5315_), .A2(new_n5308_), .ZN(new_n5316_));
  NOR2_X1    g05071(.A1(new_n5311_), .A2(new_n5307_), .ZN(new_n5317_));
  NOR2_X1    g05072(.A1(new_n5316_), .A2(new_n5317_), .ZN(new_n5318_));
  NOR2_X1    g05073(.A1(new_n5318_), .A2(new_n5314_), .ZN(new_n5319_));
  NOR2_X1    g05074(.A1(new_n5319_), .A2(new_n5313_), .ZN(new_n5320_));
  NOR2_X1    g05075(.A1(new_n4501_), .A2(new_n4770_), .ZN(new_n5321_));
  INV_X1     g05076(.I(new_n5321_), .ZN(new_n5322_));
  NAND2_X1   g05077(.A1(\a[15] ), .A2(\a[43] ), .ZN(new_n5323_));
  NOR3_X1    g05078(.A1(new_n5323_), .A2(new_n282_), .A3(new_n2765_), .ZN(new_n5324_));
  NAND4_X1   g05079(.A1(new_n5324_), .A2(\a[15] ), .A3(new_n3208_), .A4(\a[44] ), .ZN(new_n5325_));
  AOI21_X1   g05080(.A1(new_n5325_), .A2(new_n5322_), .B(new_n212_), .ZN(new_n5326_));
  NOR3_X1    g05081(.A1(new_n5326_), .A2(new_n200_), .A3(new_n4770_), .ZN(new_n5327_));
  NOR2_X1    g05082(.A1(new_n5326_), .A2(new_n5324_), .ZN(new_n5328_));
  AOI22_X1   g05083(.A1(\a[4] ), .A2(\a[15] ), .B1(\a[32] ), .B2(\a[43] ), .ZN(new_n5329_));
  AOI21_X1   g05084(.A1(new_n5328_), .A2(new_n5329_), .B(new_n5327_), .ZN(new_n5330_));
  AOI21_X1   g05085(.A1(new_n1441_), .A2(new_n2690_), .B(new_n5201_), .ZN(new_n5331_));
  INV_X1     g05086(.I(new_n5331_), .ZN(new_n5332_));
  NOR2_X1    g05087(.A1(new_n5070_), .A2(new_n5332_), .ZN(new_n5333_));
  NOR2_X1    g05088(.A1(new_n5069_), .A2(new_n5331_), .ZN(new_n5334_));
  OAI21_X1   g05089(.A1(new_n5333_), .A2(new_n5334_), .B(new_n5330_), .ZN(new_n5335_));
  XOR2_X1    g05090(.A1(new_n5069_), .A2(new_n5332_), .Z(new_n5336_));
  OAI21_X1   g05091(.A1(new_n5330_), .A2(new_n5336_), .B(new_n5335_), .ZN(new_n5337_));
  INV_X1     g05092(.I(new_n5337_), .ZN(new_n5338_));
  NOR2_X1    g05093(.A1(new_n3804_), .A2(new_n3783_), .ZN(new_n5339_));
  INV_X1     g05094(.I(new_n5339_), .ZN(new_n5340_));
  NOR2_X1    g05095(.A1(new_n675_), .A2(new_n3783_), .ZN(new_n5341_));
  NAND4_X1   g05096(.A1(new_n3805_), .A2(new_n4731_), .A3(new_n5341_), .A4(new_n5183_), .ZN(new_n5342_));
  AOI21_X1   g05097(.A1(new_n5342_), .A2(new_n5340_), .B(new_n453_), .ZN(new_n5343_));
  NOR2_X1    g05098(.A1(new_n5008_), .A2(new_n1236_), .ZN(new_n5345_));
  INV_X1     g05099(.I(new_n5345_), .ZN(new_n5346_));
  NOR2_X1    g05100(.A1(new_n2868_), .A2(new_n4414_), .ZN(new_n5347_));
  INV_X1     g05101(.I(new_n5347_), .ZN(new_n5348_));
  NOR2_X1    g05102(.A1(new_n1199_), .A2(new_n5348_), .ZN(new_n5349_));
  NOR2_X1    g05103(.A1(new_n4414_), .A2(new_n4769_), .ZN(new_n5350_));
  NOR2_X1    g05104(.A1(new_n1199_), .A2(new_n5348_), .ZN(new_n5354_));
  INV_X1     g05105(.I(new_n5354_), .ZN(new_n5355_));
  NOR2_X1    g05106(.A1(new_n2276_), .A2(new_n2285_), .ZN(new_n5356_));
  NOR2_X1    g05107(.A1(new_n1674_), .A2(new_n1999_), .ZN(new_n5357_));
  NOR2_X1    g05108(.A1(new_n5357_), .A2(new_n2543_), .ZN(new_n5358_));
  NAND2_X1   g05109(.A1(new_n5358_), .A2(new_n5356_), .ZN(new_n5359_));
  NOR2_X1    g05110(.A1(new_n461_), .A2(new_n3837_), .ZN(new_n5360_));
  XOR2_X1    g05111(.A1(new_n5359_), .A2(new_n5360_), .Z(new_n5361_));
  NOR2_X1    g05112(.A1(new_n5361_), .A2(new_n5355_), .ZN(new_n5362_));
  INV_X1     g05113(.I(new_n5361_), .ZN(new_n5363_));
  NOR2_X1    g05114(.A1(new_n5363_), .A2(new_n5354_), .ZN(new_n5364_));
  NOR2_X1    g05115(.A1(new_n5364_), .A2(new_n5362_), .ZN(new_n5365_));
  NOR2_X1    g05116(.A1(new_n5365_), .A2(new_n5346_), .ZN(new_n5366_));
  XOR2_X1    g05117(.A1(new_n5361_), .A2(new_n5354_), .Z(new_n5367_));
  NOR2_X1    g05118(.A1(new_n5367_), .A2(new_n5345_), .ZN(new_n5368_));
  NOR2_X1    g05119(.A1(new_n5366_), .A2(new_n5368_), .ZN(new_n5369_));
  NAND2_X1   g05120(.A1(\a[45] ), .A2(\a[47] ), .ZN(new_n5370_));
  XNOR2_X1   g05121(.A1(new_n197_), .A2(new_n5370_), .ZN(new_n5371_));
  INV_X1     g05122(.I(new_n5371_), .ZN(new_n5372_));
  AOI22_X1   g05123(.A1(new_n4200_), .A2(new_n3126_), .B1(new_n3733_), .B2(new_n1275_), .ZN(new_n5373_));
  INV_X1     g05124(.I(new_n5373_), .ZN(new_n5374_));
  NAND4_X1   g05125(.A1(new_n3175_), .A2(\a[16] ), .A3(\a[31] ), .A4(new_n1268_), .ZN(new_n5375_));
  AOI22_X1   g05126(.A1(new_n1769_), .A2(new_n2797_), .B1(new_n1798_), .B2(new_n3037_), .ZN(new_n5376_));
  INV_X1     g05127(.I(new_n5376_), .ZN(new_n5377_));
  NAND4_X1   g05128(.A1(new_n2534_), .A2(\a[19] ), .A3(\a[28] ), .A4(new_n1711_), .ZN(new_n5378_));
  NOR4_X1    g05129(.A1(new_n5374_), .A2(new_n5377_), .A3(new_n5375_), .A4(new_n5378_), .ZN(new_n5379_));
  NOR2_X1    g05130(.A1(new_n5374_), .A2(new_n5375_), .ZN(new_n5380_));
  NOR2_X1    g05131(.A1(new_n5377_), .A2(new_n5378_), .ZN(new_n5381_));
  NOR2_X1    g05132(.A1(new_n5380_), .A2(new_n5381_), .ZN(new_n5382_));
  OAI21_X1   g05133(.A1(new_n5382_), .A2(new_n5379_), .B(new_n5372_), .ZN(new_n5383_));
  XOR2_X1    g05134(.A1(new_n5380_), .A2(new_n5381_), .Z(new_n5384_));
  NAND2_X1   g05135(.A1(new_n5384_), .A2(new_n5371_), .ZN(new_n5385_));
  NAND2_X1   g05136(.A1(new_n5385_), .A2(new_n5383_), .ZN(new_n5386_));
  XOR2_X1    g05137(.A1(new_n5369_), .A2(new_n5386_), .Z(new_n5387_));
  NOR2_X1    g05138(.A1(new_n5387_), .A2(new_n5338_), .ZN(new_n5388_));
  INV_X1     g05139(.I(new_n5386_), .ZN(new_n5389_));
  NOR2_X1    g05140(.A1(new_n5369_), .A2(new_n5389_), .ZN(new_n5390_));
  INV_X1     g05141(.I(new_n5390_), .ZN(new_n5391_));
  NAND2_X1   g05142(.A1(new_n5369_), .A2(new_n5389_), .ZN(new_n5392_));
  AOI21_X1   g05143(.A1(new_n5391_), .A2(new_n5392_), .B(new_n5337_), .ZN(new_n5393_));
  NOR2_X1    g05144(.A1(new_n5388_), .A2(new_n5393_), .ZN(new_n5394_));
  INV_X1     g05145(.I(new_n5394_), .ZN(new_n5395_));
  AOI21_X1   g05146(.A1(new_n5200_), .A2(new_n5210_), .B(new_n5208_), .ZN(new_n5396_));
  AOI21_X1   g05147(.A1(new_n5133_), .A2(new_n5139_), .B(new_n5137_), .ZN(new_n5397_));
  AOI21_X1   g05148(.A1(new_n797_), .A2(new_n3966_), .B(new_n5185_), .ZN(new_n5398_));
  AOI21_X1   g05149(.A1(new_n609_), .A2(new_n5204_), .B(new_n5339_), .ZN(new_n5399_));
  INV_X1     g05150(.I(new_n5399_), .ZN(new_n5400_));
  NAND2_X1   g05151(.A1(\a[1] ), .A2(\a[46] ), .ZN(new_n5401_));
  XOR2_X1    g05152(.A1(new_n5401_), .A2(\a[24] ), .Z(new_n5402_));
  NOR2_X1    g05153(.A1(new_n5400_), .A2(new_n5402_), .ZN(new_n5403_));
  INV_X1     g05154(.I(new_n5402_), .ZN(new_n5404_));
  NOR2_X1    g05155(.A1(new_n5404_), .A2(new_n5399_), .ZN(new_n5405_));
  NOR2_X1    g05156(.A1(new_n5405_), .A2(new_n5403_), .ZN(new_n5406_));
  XOR2_X1    g05157(.A1(new_n5402_), .A2(new_n5399_), .Z(new_n5407_));
  MUX2_X1    g05158(.I0(new_n5407_), .I1(new_n5406_), .S(new_n5398_), .Z(new_n5408_));
  NOR2_X1    g05159(.A1(new_n5397_), .A2(new_n5408_), .ZN(new_n5409_));
  INV_X1     g05160(.I(new_n5409_), .ZN(new_n5410_));
  NAND2_X1   g05161(.A1(new_n5397_), .A2(new_n5408_), .ZN(new_n5411_));
  AOI21_X1   g05162(.A1(new_n5410_), .A2(new_n5411_), .B(new_n5396_), .ZN(new_n5412_));
  INV_X1     g05163(.I(new_n5396_), .ZN(new_n5413_));
  XNOR2_X1   g05164(.A1(new_n5397_), .A2(new_n5408_), .ZN(new_n5414_));
  NOR2_X1    g05165(.A1(new_n5414_), .A2(new_n5413_), .ZN(new_n5415_));
  NOR2_X1    g05166(.A1(new_n5415_), .A2(new_n5412_), .ZN(new_n5416_));
  NOR2_X1    g05167(.A1(new_n5395_), .A2(new_n5416_), .ZN(new_n5417_));
  INV_X1     g05168(.I(new_n5417_), .ZN(new_n5418_));
  NAND2_X1   g05169(.A1(new_n5395_), .A2(new_n5416_), .ZN(new_n5419_));
  AOI21_X1   g05170(.A1(new_n5419_), .A2(new_n5418_), .B(new_n5320_), .ZN(new_n5420_));
  XOR2_X1    g05171(.A1(new_n5394_), .A2(new_n5416_), .Z(new_n5421_));
  INV_X1     g05172(.I(new_n5421_), .ZN(new_n5422_));
  AOI21_X1   g05173(.A1(new_n5320_), .A2(new_n5422_), .B(new_n5420_), .ZN(new_n5423_));
  XNOR2_X1   g05174(.A1(new_n5286_), .A2(new_n5423_), .ZN(new_n5424_));
  NOR2_X1    g05175(.A1(new_n5424_), .A2(new_n5284_), .ZN(new_n5425_));
  NOR2_X1    g05176(.A1(new_n5286_), .A2(new_n5423_), .ZN(new_n5426_));
  INV_X1     g05177(.I(new_n5426_), .ZN(new_n5427_));
  NAND2_X1   g05178(.A1(new_n5286_), .A2(new_n5423_), .ZN(new_n5428_));
  AOI21_X1   g05179(.A1(new_n5427_), .A2(new_n5428_), .B(new_n5283_), .ZN(new_n5429_));
  NOR2_X1    g05180(.A1(new_n5425_), .A2(new_n5429_), .ZN(new_n5430_));
  NOR2_X1    g05181(.A1(new_n5430_), .A2(new_n5236_), .ZN(new_n5431_));
  XOR2_X1    g05182(.A1(new_n5234_), .A2(new_n5431_), .Z(new_n5432_));
  XOR2_X1    g05183(.A1(new_n5432_), .A2(new_n5229_), .Z(\asquared[48] ));
  INV_X1     g05184(.I(new_n5431_), .ZN(new_n5434_));
  AOI21_X1   g05185(.A1(new_n5236_), .A2(new_n5430_), .B(new_n5229_), .ZN(new_n5435_));
  NAND3_X1   g05186(.A1(new_n4859_), .A2(new_n5233_), .A3(new_n5435_), .ZN(new_n5436_));
  NAND2_X1   g05187(.A1(new_n5436_), .A2(new_n5434_), .ZN(new_n5437_));
  INV_X1     g05188(.I(new_n5278_), .ZN(new_n5438_));
  AOI21_X1   g05189(.A1(new_n5237_), .A2(new_n5438_), .B(new_n5280_), .ZN(new_n5439_));
  AOI21_X1   g05190(.A1(new_n5320_), .A2(new_n5419_), .B(new_n5417_), .ZN(new_n5440_));
  OAI21_X1   g05191(.A1(new_n5240_), .A2(new_n5261_), .B(new_n5263_), .ZN(new_n5441_));
  INV_X1     g05192(.I(new_n5441_), .ZN(new_n5442_));
  INV_X1     g05193(.I(new_n5334_), .ZN(new_n5443_));
  AOI21_X1   g05194(.A1(new_n5330_), .A2(new_n5443_), .B(new_n5333_), .ZN(new_n5444_));
  AOI21_X1   g05195(.A1(new_n5243_), .A2(new_n5254_), .B(new_n5252_), .ZN(new_n5445_));
  NAND2_X1   g05196(.A1(\a[1] ), .A2(\a[47] ), .ZN(new_n5446_));
  NAND2_X1   g05197(.A1(new_n1912_), .A2(new_n5446_), .ZN(new_n5447_));
  NOR2_X1    g05198(.A1(new_n1912_), .A2(new_n5446_), .ZN(new_n5448_));
  INV_X1     g05199(.I(new_n5448_), .ZN(new_n5449_));
  NAND2_X1   g05200(.A1(new_n5449_), .A2(new_n5447_), .ZN(new_n5450_));
  NOR2_X1    g05201(.A1(new_n1801_), .A2(new_n5175_), .ZN(new_n5451_));
  NAND2_X1   g05202(.A1(new_n5450_), .A2(new_n5451_), .ZN(new_n5452_));
  XOR2_X1    g05203(.A1(new_n5452_), .A2(\a[0] ), .Z(new_n5453_));
  XOR2_X1    g05204(.A1(new_n5453_), .A2(\a[48] ), .Z(new_n5454_));
  XNOR2_X1   g05205(.A1(new_n5454_), .A2(new_n5445_), .ZN(new_n5455_));
  NOR2_X1    g05206(.A1(new_n5454_), .A2(new_n5445_), .ZN(new_n5456_));
  NAND2_X1   g05207(.A1(new_n5454_), .A2(new_n5445_), .ZN(new_n5457_));
  INV_X1     g05208(.I(new_n5457_), .ZN(new_n5458_));
  OAI21_X1   g05209(.A1(new_n5458_), .A2(new_n5456_), .B(new_n5444_), .ZN(new_n5459_));
  OAI21_X1   g05210(.A1(new_n5444_), .A2(new_n5455_), .B(new_n5459_), .ZN(new_n5460_));
  AOI21_X1   g05211(.A1(new_n5413_), .A2(new_n5411_), .B(new_n5409_), .ZN(new_n5461_));
  XNOR2_X1   g05212(.A1(new_n5460_), .A2(new_n5461_), .ZN(new_n5462_));
  NOR2_X1    g05213(.A1(new_n5462_), .A2(new_n5442_), .ZN(new_n5463_));
  NOR2_X1    g05214(.A1(new_n5460_), .A2(new_n5461_), .ZN(new_n5464_));
  INV_X1     g05215(.I(new_n5464_), .ZN(new_n5465_));
  NAND2_X1   g05216(.A1(new_n5460_), .A2(new_n5461_), .ZN(new_n5466_));
  AOI21_X1   g05217(.A1(new_n5465_), .A2(new_n5466_), .B(new_n5441_), .ZN(new_n5467_));
  NOR2_X1    g05218(.A1(new_n5463_), .A2(new_n5467_), .ZN(new_n5468_));
  AOI21_X1   g05219(.A1(new_n5337_), .A2(new_n5392_), .B(new_n5390_), .ZN(new_n5469_));
  AOI21_X1   g05220(.A1(new_n5183_), .A2(new_n3805_), .B(new_n5343_), .ZN(new_n5470_));
  INV_X1     g05221(.I(new_n5470_), .ZN(new_n5471_));
  AOI21_X1   g05222(.A1(new_n608_), .A2(new_n5350_), .B(new_n5349_), .ZN(new_n5472_));
  AOI21_X1   g05223(.A1(new_n2978_), .A2(new_n2533_), .B(new_n5376_), .ZN(new_n5473_));
  XNOR2_X1   g05224(.A1(new_n5472_), .A2(new_n5473_), .ZN(new_n5474_));
  INV_X1     g05225(.I(new_n5472_), .ZN(new_n5475_));
  INV_X1     g05226(.I(new_n5473_), .ZN(new_n5476_));
  NOR2_X1    g05227(.A1(new_n5475_), .A2(new_n5476_), .ZN(new_n5477_));
  NOR2_X1    g05228(.A1(new_n5472_), .A2(new_n5473_), .ZN(new_n5478_));
  OAI21_X1   g05229(.A1(new_n5478_), .A2(new_n5477_), .B(new_n5471_), .ZN(new_n5479_));
  OAI21_X1   g05230(.A1(new_n5471_), .A2(new_n5474_), .B(new_n5479_), .ZN(new_n5480_));
  INV_X1     g05231(.I(new_n5362_), .ZN(new_n5481_));
  OAI21_X1   g05232(.A1(new_n5346_), .A2(new_n5364_), .B(new_n5481_), .ZN(new_n5482_));
  INV_X1     g05233(.I(new_n5482_), .ZN(new_n5483_));
  AOI21_X1   g05234(.A1(new_n1220_), .A2(new_n3487_), .B(new_n5293_), .ZN(new_n5484_));
  NAND2_X1   g05235(.A1(new_n461_), .A2(new_n3837_), .ZN(new_n5485_));
  OAI21_X1   g05236(.A1(new_n5356_), .A2(new_n5485_), .B(new_n5358_), .ZN(new_n5486_));
  NOR2_X1    g05237(.A1(new_n2765_), .A2(new_n5175_), .ZN(new_n5487_));
  NOR2_X1    g05238(.A1(new_n5004_), .A2(new_n5175_), .ZN(new_n5488_));
  AOI22_X1   g05239(.A1(new_n5487_), .A2(new_n5488_), .B1(new_n1025_), .B2(new_n232_), .ZN(new_n5489_));
  NAND2_X1   g05240(.A1(\a[3] ), .A2(\a[45] ), .ZN(new_n5490_));
  INV_X1     g05241(.I(new_n5490_), .ZN(new_n5491_));
  NAND2_X1   g05242(.A1(\a[16] ), .A2(\a[32] ), .ZN(new_n5492_));
  OAI21_X1   g05243(.A1(new_n5491_), .A2(new_n5492_), .B(new_n5489_), .ZN(new_n5493_));
  XNOR2_X1   g05244(.A1(new_n5490_), .A2(new_n5492_), .ZN(new_n5494_));
  OAI21_X1   g05245(.A1(new_n201_), .A2(new_n5175_), .B(new_n5494_), .ZN(new_n5495_));
  NAND2_X1   g05246(.A1(new_n5495_), .A2(new_n5493_), .ZN(new_n5496_));
  NOR2_X1    g05247(.A1(new_n5496_), .A2(new_n5486_), .ZN(new_n5497_));
  INV_X1     g05248(.I(new_n5497_), .ZN(new_n5498_));
  NAND2_X1   g05249(.A1(new_n5496_), .A2(new_n5486_), .ZN(new_n5499_));
  NAND2_X1   g05250(.A1(new_n5498_), .A2(new_n5499_), .ZN(new_n5500_));
  XNOR2_X1   g05251(.A1(new_n5496_), .A2(new_n5486_), .ZN(new_n5501_));
  NOR2_X1    g05252(.A1(new_n5501_), .A2(new_n5484_), .ZN(new_n5502_));
  AOI21_X1   g05253(.A1(new_n5484_), .A2(new_n5500_), .B(new_n5502_), .ZN(new_n5503_));
  NOR2_X1    g05254(.A1(new_n5503_), .A2(new_n5483_), .ZN(new_n5504_));
  INV_X1     g05255(.I(new_n5504_), .ZN(new_n5505_));
  NAND2_X1   g05256(.A1(new_n5503_), .A2(new_n5483_), .ZN(new_n5506_));
  NAND2_X1   g05257(.A1(new_n5505_), .A2(new_n5506_), .ZN(new_n5507_));
  XOR2_X1    g05258(.A1(new_n5503_), .A2(new_n5482_), .Z(new_n5508_));
  NOR2_X1    g05259(.A1(new_n5508_), .A2(new_n5480_), .ZN(new_n5509_));
  AOI21_X1   g05260(.A1(new_n5480_), .A2(new_n5507_), .B(new_n5509_), .ZN(new_n5510_));
  INV_X1     g05261(.I(\a[47] ), .ZN(new_n5511_));
  NOR2_X1    g05262(.A1(new_n5004_), .A2(new_n5511_), .ZN(new_n5512_));
  NOR3_X1    g05263(.A1(new_n2384_), .A2(new_n194_), .A3(new_n5004_), .ZN(new_n5513_));
  AOI21_X1   g05264(.A1(new_n5513_), .A2(new_n218_), .B(new_n5512_), .ZN(new_n5514_));
  AOI21_X1   g05265(.A1(new_n1441_), .A2(new_n2898_), .B(new_n5373_), .ZN(new_n5515_));
  XOR2_X1    g05266(.A1(new_n5515_), .A2(new_n5514_), .Z(new_n5516_));
  NOR3_X1    g05267(.A1(new_n5516_), .A2(new_n5324_), .A3(new_n5326_), .ZN(new_n5517_));
  INV_X1     g05268(.I(new_n5515_), .ZN(new_n5518_));
  NOR2_X1    g05269(.A1(new_n5518_), .A2(new_n5514_), .ZN(new_n5519_));
  INV_X1     g05270(.I(new_n5519_), .ZN(new_n5520_));
  NAND2_X1   g05271(.A1(new_n5518_), .A2(new_n5514_), .ZN(new_n5521_));
  AOI21_X1   g05272(.A1(new_n5520_), .A2(new_n5521_), .B(new_n5328_), .ZN(new_n5522_));
  NOR2_X1    g05273(.A1(new_n5517_), .A2(new_n5522_), .ZN(new_n5523_));
  INV_X1     g05274(.I(new_n5403_), .ZN(new_n5524_));
  AOI21_X1   g05275(.A1(new_n5524_), .A2(new_n5398_), .B(new_n5405_), .ZN(new_n5525_));
  NOR2_X1    g05276(.A1(new_n5382_), .A2(new_n5371_), .ZN(new_n5526_));
  NOR2_X1    g05277(.A1(new_n5526_), .A2(new_n5379_), .ZN(new_n5527_));
  NOR2_X1    g05278(.A1(new_n5527_), .A2(new_n5525_), .ZN(new_n5528_));
  INV_X1     g05279(.I(new_n5525_), .ZN(new_n5529_));
  NOR3_X1    g05280(.A1(new_n5529_), .A2(new_n5379_), .A3(new_n5526_), .ZN(new_n5530_));
  NOR2_X1    g05281(.A1(new_n5528_), .A2(new_n5530_), .ZN(new_n5531_));
  NOR2_X1    g05282(.A1(new_n5531_), .A2(new_n5523_), .ZN(new_n5532_));
  XOR2_X1    g05283(.A1(new_n5527_), .A2(new_n5529_), .Z(new_n5533_));
  INV_X1     g05284(.I(new_n5533_), .ZN(new_n5534_));
  AOI21_X1   g05285(.A1(new_n5523_), .A2(new_n5534_), .B(new_n5532_), .ZN(new_n5535_));
  XOR2_X1    g05286(.A1(new_n5510_), .A2(new_n5535_), .Z(new_n5536_));
  INV_X1     g05287(.I(new_n5536_), .ZN(new_n5537_));
  NOR2_X1    g05288(.A1(new_n5510_), .A2(new_n5535_), .ZN(new_n5538_));
  NAND2_X1   g05289(.A1(new_n5510_), .A2(new_n5535_), .ZN(new_n5539_));
  INV_X1     g05290(.I(new_n5539_), .ZN(new_n5540_));
  OAI21_X1   g05291(.A1(new_n5540_), .A2(new_n5538_), .B(new_n5469_), .ZN(new_n5541_));
  OAI21_X1   g05292(.A1(new_n5537_), .A2(new_n5469_), .B(new_n5541_), .ZN(new_n5542_));
  XOR2_X1    g05293(.A1(new_n5542_), .A2(new_n5468_), .Z(new_n5543_));
  NOR2_X1    g05294(.A1(new_n5543_), .A2(new_n5440_), .ZN(new_n5544_));
  INV_X1     g05295(.I(new_n5440_), .ZN(new_n5545_));
  INV_X1     g05296(.I(new_n5468_), .ZN(new_n5546_));
  NAND2_X1   g05297(.A1(new_n5542_), .A2(new_n5546_), .ZN(new_n5547_));
  NOR2_X1    g05298(.A1(new_n5542_), .A2(new_n5546_), .ZN(new_n5548_));
  INV_X1     g05299(.I(new_n5548_), .ZN(new_n5549_));
  AOI21_X1   g05300(.A1(new_n5549_), .A2(new_n5547_), .B(new_n5545_), .ZN(new_n5550_));
  NOR2_X1    g05301(.A1(new_n5544_), .A2(new_n5550_), .ZN(new_n5551_));
  OAI21_X1   g05302(.A1(new_n5274_), .A2(new_n5271_), .B(new_n5270_), .ZN(new_n5552_));
  NOR2_X1    g05303(.A1(new_n5317_), .A2(new_n5287_), .ZN(new_n5553_));
  NOR2_X1    g05304(.A1(new_n5553_), .A2(new_n5316_), .ZN(new_n5554_));
  INV_X1     g05305(.I(new_n5304_), .ZN(new_n5555_));
  AOI21_X1   g05306(.A1(new_n5301_), .A2(new_n5555_), .B(new_n5303_), .ZN(new_n5556_));
  NOR2_X1    g05307(.A1(new_n2868_), .A2(new_n4501_), .ZN(new_n5557_));
  NOR4_X1    g05308(.A1(new_n282_), .A2(new_n875_), .A3(new_n2868_), .A4(new_n4770_), .ZN(new_n5558_));
  NAND3_X1   g05309(.A1(new_n5558_), .A2(new_n5246_), .A3(new_n5557_), .ZN(new_n5559_));
  AOI21_X1   g05310(.A1(new_n5559_), .A2(new_n5322_), .B(new_n211_), .ZN(new_n5560_));
  NOR3_X1    g05311(.A1(new_n5560_), .A2(new_n282_), .A3(new_n4770_), .ZN(new_n5561_));
  INV_X1     g05312(.I(new_n5246_), .ZN(new_n5562_));
  INV_X1     g05313(.I(new_n5557_), .ZN(new_n5563_));
  OAI22_X1   g05314(.A1(new_n5562_), .A2(new_n5563_), .B1(new_n5322_), .B2(new_n211_), .ZN(new_n5564_));
  NOR3_X1    g05315(.A1(new_n5564_), .A2(new_n5246_), .A3(new_n5557_), .ZN(new_n5565_));
  NOR2_X1    g05316(.A1(new_n5561_), .A2(new_n5565_), .ZN(new_n5566_));
  AOI22_X1   g05317(.A1(new_n2978_), .A2(new_n3037_), .B1(new_n4437_), .B2(new_n2797_), .ZN(new_n5567_));
  INV_X1     g05318(.I(new_n5567_), .ZN(new_n5568_));
  NAND4_X1   g05319(.A1(new_n2534_), .A2(\a[20] ), .A3(\a[28] ), .A4(new_n1773_), .ZN(new_n5569_));
  AOI22_X1   g05320(.A1(new_n1441_), .A2(new_n3733_), .B1(new_n3126_), .B2(new_n4345_), .ZN(new_n5570_));
  INV_X1     g05321(.I(new_n5570_), .ZN(new_n5571_));
  NAND4_X1   g05322(.A1(new_n3175_), .A2(\a[17] ), .A3(\a[31] ), .A4(new_n1342_), .ZN(new_n5572_));
  NOR4_X1    g05323(.A1(new_n5571_), .A2(new_n5568_), .A3(new_n5569_), .A4(new_n5572_), .ZN(new_n5573_));
  NOR2_X1    g05324(.A1(new_n5568_), .A2(new_n5569_), .ZN(new_n5574_));
  NOR2_X1    g05325(.A1(new_n5571_), .A2(new_n5572_), .ZN(new_n5575_));
  NOR2_X1    g05326(.A1(new_n5575_), .A2(new_n5574_), .ZN(new_n5576_));
  OAI21_X1   g05327(.A1(new_n5573_), .A2(new_n5576_), .B(new_n5566_), .ZN(new_n5577_));
  XNOR2_X1   g05328(.A1(new_n5575_), .A2(new_n5574_), .ZN(new_n5578_));
  OAI21_X1   g05329(.A1(new_n5566_), .A2(new_n5578_), .B(new_n5577_), .ZN(new_n5579_));
  NAND2_X1   g05330(.A1(\a[6] ), .A2(\a[13] ), .ZN(new_n5580_));
  NAND2_X1   g05331(.A1(\a[35] ), .A2(\a[42] ), .ZN(new_n5581_));
  NOR2_X1    g05332(.A1(new_n5580_), .A2(new_n5581_), .ZN(new_n5582_));
  NOR4_X1    g05333(.A1(new_n242_), .A2(new_n650_), .A3(new_n3371_), .A4(new_n4769_), .ZN(new_n5583_));
  NAND2_X1   g05334(.A1(new_n5583_), .A2(new_n5582_), .ZN(new_n5584_));
  AOI21_X1   g05335(.A1(new_n5584_), .A2(new_n786_), .B(new_n3712_), .ZN(new_n5585_));
  NOR3_X1    g05336(.A1(new_n5585_), .A2(new_n650_), .A3(new_n3371_), .ZN(new_n5586_));
  OAI22_X1   g05337(.A1(new_n3712_), .A2(new_n786_), .B1(new_n5580_), .B2(new_n5581_), .ZN(new_n5587_));
  INV_X1     g05338(.I(new_n5587_), .ZN(new_n5588_));
  AND3_X2    g05339(.A1(new_n5588_), .A2(new_n5580_), .A3(new_n5581_), .Z(new_n5589_));
  NOR2_X1    g05340(.A1(new_n5589_), .A2(new_n5586_), .ZN(new_n5590_));
  NOR2_X1    g05341(.A1(new_n268_), .A2(new_n4414_), .ZN(new_n5591_));
  NOR2_X1    g05342(.A1(new_n4240_), .A2(new_n4414_), .ZN(new_n5592_));
  AOI22_X1   g05343(.A1(new_n3969_), .A2(new_n5591_), .B1(new_n5592_), .B2(new_n609_), .ZN(new_n5593_));
  INV_X1     g05344(.I(new_n5593_), .ZN(new_n5594_));
  INV_X1     g05345(.I(new_n4731_), .ZN(new_n5595_));
  NOR2_X1    g05346(.A1(new_n5595_), .A2(new_n5292_), .ZN(new_n5596_));
  INV_X1     g05347(.I(new_n5596_), .ZN(new_n5597_));
  AOI22_X1   g05348(.A1(\a[8] ), .A2(\a[12] ), .B1(\a[36] ), .B2(\a[40] ), .ZN(new_n5598_));
  NAND4_X1   g05349(.A1(new_n5597_), .A2(new_n5591_), .A3(new_n5594_), .A4(new_n5598_), .ZN(new_n5599_));
  INV_X1     g05350(.I(new_n4706_), .ZN(new_n5600_));
  NOR2_X1    g05351(.A1(new_n3837_), .A2(new_n3783_), .ZN(new_n5601_));
  AOI22_X1   g05352(.A1(new_n597_), .A2(new_n5601_), .B1(new_n5339_), .B2(new_n5183_), .ZN(new_n5602_));
  INV_X1     g05353(.I(new_n5602_), .ZN(new_n5603_));
  NOR2_X1    g05354(.A1(new_n364_), .A2(new_n3783_), .ZN(new_n5604_));
  INV_X1     g05355(.I(new_n5604_), .ZN(new_n5605_));
  NOR4_X1    g05356(.A1(new_n5603_), .A2(new_n797_), .A3(new_n5600_), .A4(new_n5605_), .ZN(new_n5606_));
  INV_X1     g05357(.I(new_n5606_), .ZN(new_n5607_));
  NOR2_X1    g05358(.A1(new_n5607_), .A2(new_n5599_), .ZN(new_n5608_));
  NAND2_X1   g05359(.A1(new_n5607_), .A2(new_n5599_), .ZN(new_n5609_));
  INV_X1     g05360(.I(new_n5609_), .ZN(new_n5610_));
  OAI21_X1   g05361(.A1(new_n5610_), .A2(new_n5608_), .B(new_n5590_), .ZN(new_n5611_));
  XOR2_X1    g05362(.A1(new_n5599_), .A2(new_n5606_), .Z(new_n5612_));
  OAI21_X1   g05363(.A1(new_n5590_), .A2(new_n5612_), .B(new_n5611_), .ZN(new_n5613_));
  XNOR2_X1   g05364(.A1(new_n5613_), .A2(new_n5579_), .ZN(new_n5614_));
  NOR2_X1    g05365(.A1(new_n5614_), .A2(new_n5556_), .ZN(new_n5615_));
  INV_X1     g05366(.I(new_n5556_), .ZN(new_n5616_));
  NAND2_X1   g05367(.A1(new_n5613_), .A2(new_n5579_), .ZN(new_n5617_));
  NOR2_X1    g05368(.A1(new_n5613_), .A2(new_n5579_), .ZN(new_n5618_));
  INV_X1     g05369(.I(new_n5618_), .ZN(new_n5619_));
  AOI21_X1   g05370(.A1(new_n5619_), .A2(new_n5617_), .B(new_n5616_), .ZN(new_n5620_));
  NOR2_X1    g05371(.A1(new_n5615_), .A2(new_n5620_), .ZN(new_n5621_));
  XOR2_X1    g05372(.A1(new_n5554_), .A2(new_n5621_), .Z(new_n5622_));
  INV_X1     g05373(.I(new_n5622_), .ZN(new_n5623_));
  INV_X1     g05374(.I(new_n5621_), .ZN(new_n5624_));
  NAND2_X1   g05375(.A1(new_n5554_), .A2(new_n5624_), .ZN(new_n5625_));
  NOR2_X1    g05376(.A1(new_n5554_), .A2(new_n5624_), .ZN(new_n5626_));
  INV_X1     g05377(.I(new_n5626_), .ZN(new_n5627_));
  AOI21_X1   g05378(.A1(new_n5627_), .A2(new_n5625_), .B(new_n5552_), .ZN(new_n5628_));
  AOI21_X1   g05379(.A1(new_n5623_), .A2(new_n5552_), .B(new_n5628_), .ZN(new_n5629_));
  XOR2_X1    g05380(.A1(new_n5551_), .A2(new_n5629_), .Z(new_n5630_));
  INV_X1     g05381(.I(new_n5630_), .ZN(new_n5631_));
  NOR2_X1    g05382(.A1(new_n5551_), .A2(new_n5629_), .ZN(new_n5632_));
  NAND2_X1   g05383(.A1(new_n5551_), .A2(new_n5629_), .ZN(new_n5633_));
  INV_X1     g05384(.I(new_n5633_), .ZN(new_n5634_));
  OAI21_X1   g05385(.A1(new_n5634_), .A2(new_n5632_), .B(new_n5439_), .ZN(new_n5635_));
  OAI21_X1   g05386(.A1(new_n5631_), .A2(new_n5439_), .B(new_n5635_), .ZN(new_n5636_));
  OAI21_X1   g05387(.A1(new_n5284_), .A2(new_n5426_), .B(new_n5428_), .ZN(new_n5637_));
  INV_X1     g05388(.I(new_n5637_), .ZN(new_n5638_));
  NOR2_X1    g05389(.A1(new_n5636_), .A2(new_n5638_), .ZN(new_n5639_));
  INV_X1     g05390(.I(new_n5639_), .ZN(new_n5640_));
  NAND2_X1   g05391(.A1(new_n5636_), .A2(new_n5638_), .ZN(new_n5641_));
  NAND2_X1   g05392(.A1(new_n5640_), .A2(new_n5641_), .ZN(new_n5642_));
  XOR2_X1    g05393(.A1(new_n5437_), .A2(new_n5642_), .Z(\asquared[49] ));
  OAI21_X1   g05394(.A1(new_n5437_), .A2(new_n5639_), .B(new_n5641_), .ZN(new_n5644_));
  AOI21_X1   g05395(.A1(new_n5545_), .A2(new_n5547_), .B(new_n5548_), .ZN(new_n5645_));
  AOI21_X1   g05396(.A1(new_n5552_), .A2(new_n5625_), .B(new_n5626_), .ZN(new_n5646_));
  INV_X1     g05397(.I(new_n5444_), .ZN(new_n5647_));
  AOI21_X1   g05398(.A1(new_n5647_), .A2(new_n5457_), .B(new_n5456_), .ZN(new_n5648_));
  INV_X1     g05399(.I(new_n5648_), .ZN(new_n5649_));
  NOR3_X1    g05400(.A1(new_n5576_), .A2(new_n5561_), .A3(new_n5565_), .ZN(new_n5650_));
  NOR2_X1    g05401(.A1(new_n5650_), .A2(new_n5573_), .ZN(new_n5651_));
  NOR2_X1    g05402(.A1(new_n5594_), .A2(new_n5596_), .ZN(new_n5652_));
  AOI21_X1   g05403(.A1(new_n2331_), .A2(new_n2898_), .B(new_n5570_), .ZN(new_n5653_));
  XOR2_X1    g05404(.A1(new_n5653_), .A2(new_n5588_), .Z(new_n5654_));
  INV_X1     g05405(.I(new_n5653_), .ZN(new_n5655_));
  NOR2_X1    g05406(.A1(new_n5655_), .A2(new_n5587_), .ZN(new_n5656_));
  NOR2_X1    g05407(.A1(new_n5653_), .A2(new_n5588_), .ZN(new_n5657_));
  NOR2_X1    g05408(.A1(new_n5656_), .A2(new_n5657_), .ZN(new_n5658_));
  NOR2_X1    g05409(.A1(new_n5658_), .A2(new_n5652_), .ZN(new_n5659_));
  AOI21_X1   g05410(.A1(new_n5652_), .A2(new_n5654_), .B(new_n5659_), .ZN(new_n5660_));
  XOR2_X1    g05411(.A1(new_n5660_), .A2(new_n5651_), .Z(new_n5661_));
  INV_X1     g05412(.I(new_n5661_), .ZN(new_n5662_));
  INV_X1     g05413(.I(new_n5651_), .ZN(new_n5663_));
  NOR2_X1    g05414(.A1(new_n5660_), .A2(new_n5663_), .ZN(new_n5664_));
  INV_X1     g05415(.I(new_n5664_), .ZN(new_n5665_));
  NAND2_X1   g05416(.A1(new_n5660_), .A2(new_n5663_), .ZN(new_n5666_));
  AOI21_X1   g05417(.A1(new_n5665_), .A2(new_n5666_), .B(new_n5649_), .ZN(new_n5667_));
  AOI21_X1   g05418(.A1(new_n5649_), .A2(new_n5662_), .B(new_n5667_), .ZN(new_n5668_));
  INV_X1     g05419(.I(new_n5668_), .ZN(new_n5669_));
  OAI21_X1   g05420(.A1(new_n5556_), .A2(new_n5618_), .B(new_n5617_), .ZN(new_n5670_));
  AOI21_X1   g05421(.A1(new_n4538_), .A2(new_n2533_), .B(new_n5567_), .ZN(new_n5671_));
  NOR2_X1    g05422(.A1(new_n5490_), .A2(new_n5492_), .ZN(new_n5672_));
  NOR2_X1    g05423(.A1(new_n5489_), .A2(new_n5672_), .ZN(new_n5673_));
  XNOR2_X1   g05424(.A1(new_n5671_), .A2(new_n5673_), .ZN(new_n5674_));
  NOR2_X1    g05425(.A1(new_n5674_), .A2(new_n5564_), .ZN(new_n5675_));
  INV_X1     g05426(.I(new_n5564_), .ZN(new_n5676_));
  NAND2_X1   g05427(.A1(new_n5671_), .A2(new_n5673_), .ZN(new_n5677_));
  NOR2_X1    g05428(.A1(new_n5671_), .A2(new_n5673_), .ZN(new_n5678_));
  INV_X1     g05429(.I(new_n5678_), .ZN(new_n5679_));
  AOI21_X1   g05430(.A1(new_n5679_), .A2(new_n5677_), .B(new_n5676_), .ZN(new_n5680_));
  NOR2_X1    g05431(.A1(new_n5675_), .A2(new_n5680_), .ZN(new_n5681_));
  AOI21_X1   g05432(.A1(new_n5590_), .A2(new_n5609_), .B(new_n5608_), .ZN(new_n5682_));
  AOI21_X1   g05433(.A1(new_n797_), .A2(new_n5600_), .B(new_n5602_), .ZN(new_n5683_));
  INV_X1     g05434(.I(new_n5683_), .ZN(new_n5684_));
  NAND2_X1   g05435(.A1(\a[1] ), .A2(\a[48] ), .ZN(new_n5685_));
  XOR2_X1    g05436(.A1(new_n5685_), .A2(\a[25] ), .Z(new_n5686_));
  XOR2_X1    g05437(.A1(new_n5686_), .A2(new_n5448_), .Z(new_n5687_));
  NOR2_X1    g05438(.A1(new_n5686_), .A2(new_n5449_), .ZN(new_n5688_));
  NAND2_X1   g05439(.A1(new_n5686_), .A2(new_n5449_), .ZN(new_n5689_));
  INV_X1     g05440(.I(new_n5689_), .ZN(new_n5690_));
  OAI21_X1   g05441(.A1(new_n5688_), .A2(new_n5690_), .B(new_n5684_), .ZN(new_n5691_));
  OAI21_X1   g05442(.A1(new_n5687_), .A2(new_n5684_), .B(new_n5691_), .ZN(new_n5692_));
  NAND2_X1   g05443(.A1(new_n5682_), .A2(new_n5692_), .ZN(new_n5693_));
  NOR2_X1    g05444(.A1(new_n5682_), .A2(new_n5692_), .ZN(new_n5694_));
  INV_X1     g05445(.I(new_n5694_), .ZN(new_n5695_));
  AOI21_X1   g05446(.A1(new_n5695_), .A2(new_n5693_), .B(new_n5681_), .ZN(new_n5696_));
  XNOR2_X1   g05447(.A1(new_n5682_), .A2(new_n5692_), .ZN(new_n5697_));
  INV_X1     g05448(.I(new_n5697_), .ZN(new_n5698_));
  AOI21_X1   g05449(.A1(new_n5698_), .A2(new_n5681_), .B(new_n5696_), .ZN(new_n5699_));
  NOR2_X1    g05450(.A1(new_n5699_), .A2(new_n5670_), .ZN(new_n5700_));
  NAND2_X1   g05451(.A1(new_n5699_), .A2(new_n5670_), .ZN(new_n5701_));
  INV_X1     g05452(.I(new_n5701_), .ZN(new_n5702_));
  OAI21_X1   g05453(.A1(new_n5700_), .A2(new_n5702_), .B(new_n5669_), .ZN(new_n5703_));
  XOR2_X1    g05454(.A1(new_n5699_), .A2(new_n5670_), .Z(new_n5704_));
  NAND2_X1   g05455(.A1(new_n5704_), .A2(new_n5668_), .ZN(new_n5705_));
  NAND2_X1   g05456(.A1(new_n5703_), .A2(new_n5705_), .ZN(new_n5706_));
  INV_X1     g05457(.I(new_n5477_), .ZN(new_n5707_));
  OAI21_X1   g05458(.A1(new_n5471_), .A2(new_n5478_), .B(new_n5707_), .ZN(new_n5708_));
  NAND2_X1   g05459(.A1(new_n5499_), .A2(new_n5484_), .ZN(new_n5709_));
  NAND2_X1   g05460(.A1(new_n5709_), .A2(new_n5498_), .ZN(new_n5710_));
  AOI21_X1   g05461(.A1(new_n5328_), .A2(new_n5521_), .B(new_n5519_), .ZN(new_n5711_));
  INV_X1     g05462(.I(new_n5711_), .ZN(new_n5712_));
  XOR2_X1    g05463(.A1(new_n5710_), .A2(new_n5712_), .Z(new_n5713_));
  NAND2_X1   g05464(.A1(new_n5710_), .A2(new_n5712_), .ZN(new_n5714_));
  NAND3_X1   g05465(.A1(new_n5711_), .A2(new_n5709_), .A3(new_n5498_), .ZN(new_n5715_));
  AOI21_X1   g05466(.A1(new_n5714_), .A2(new_n5715_), .B(new_n5708_), .ZN(new_n5716_));
  AOI21_X1   g05467(.A1(new_n5713_), .A2(new_n5708_), .B(new_n5716_), .ZN(new_n5717_));
  INV_X1     g05468(.I(new_n5480_), .ZN(new_n5718_));
  AOI21_X1   g05469(.A1(new_n5718_), .A2(new_n5506_), .B(new_n5504_), .ZN(new_n5719_));
  INV_X1     g05470(.I(new_n5530_), .ZN(new_n5720_));
  AOI21_X1   g05471(.A1(new_n5523_), .A2(new_n5720_), .B(new_n5528_), .ZN(new_n5721_));
  NOR2_X1    g05472(.A1(new_n5719_), .A2(new_n5721_), .ZN(new_n5722_));
  INV_X1     g05473(.I(new_n5722_), .ZN(new_n5723_));
  NAND2_X1   g05474(.A1(new_n5719_), .A2(new_n5721_), .ZN(new_n5724_));
  NAND2_X1   g05475(.A1(new_n5723_), .A2(new_n5724_), .ZN(new_n5725_));
  INV_X1     g05476(.I(new_n5725_), .ZN(new_n5726_));
  NOR2_X1    g05477(.A1(new_n5726_), .A2(new_n5717_), .ZN(new_n5727_));
  XNOR2_X1   g05478(.A1(new_n5719_), .A2(new_n5721_), .ZN(new_n5728_));
  INV_X1     g05479(.I(new_n5728_), .ZN(new_n5729_));
  AOI21_X1   g05480(.A1(new_n5717_), .A2(new_n5729_), .B(new_n5727_), .ZN(new_n5730_));
  XOR2_X1    g05481(.A1(new_n5730_), .A2(new_n5706_), .Z(new_n5731_));
  AOI21_X1   g05482(.A1(new_n5703_), .A2(new_n5705_), .B(new_n5730_), .ZN(new_n5732_));
  INV_X1     g05483(.I(new_n5730_), .ZN(new_n5733_));
  NOR2_X1    g05484(.A1(new_n5733_), .A2(new_n5706_), .ZN(new_n5734_));
  OAI21_X1   g05485(.A1(new_n5734_), .A2(new_n5732_), .B(new_n5646_), .ZN(new_n5735_));
  OAI21_X1   g05486(.A1(new_n5646_), .A2(new_n5731_), .B(new_n5735_), .ZN(new_n5736_));
  OAI21_X1   g05487(.A1(new_n5469_), .A2(new_n5538_), .B(new_n5539_), .ZN(new_n5737_));
  NAND2_X1   g05488(.A1(new_n5466_), .A2(new_n5441_), .ZN(new_n5738_));
  NAND2_X1   g05489(.A1(new_n5738_), .A2(new_n5465_), .ZN(new_n5739_));
  AOI22_X1   g05490(.A1(\a[44] ), .A2(new_n1011_), .B1(new_n3123_), .B2(\a[45] ), .ZN(new_n5740_));
  NOR2_X1    g05491(.A1(new_n5740_), .A2(\a[49] ), .ZN(new_n5741_));
  NOR2_X1    g05492(.A1(new_n4770_), .A2(new_n5004_), .ZN(new_n5742_));
  INV_X1     g05493(.I(new_n5742_), .ZN(new_n5743_));
  OR3_X2     g05494(.A1(new_n5741_), .A2(new_n211_), .A3(new_n5743_), .Z(new_n5744_));
  INV_X1     g05495(.I(\a[49] ), .ZN(new_n5745_));
  NOR2_X1    g05496(.A1(new_n199_), .A2(new_n5745_), .ZN(new_n5746_));
  AOI21_X1   g05497(.A1(\a[44] ), .A2(\a[45] ), .B(new_n229_), .ZN(new_n5747_));
  AOI21_X1   g05498(.A1(new_n5744_), .A2(new_n5746_), .B(new_n5747_), .ZN(new_n5748_));
  INV_X1     g05499(.I(new_n5748_), .ZN(new_n5749_));
  INV_X1     g05500(.I(\a[48] ), .ZN(new_n5750_));
  NOR2_X1    g05501(.A1(new_n199_), .A2(new_n5750_), .ZN(new_n5751_));
  OAI21_X1   g05502(.A1(new_n5450_), .A2(new_n5451_), .B(new_n5751_), .ZN(new_n5752_));
  NAND2_X1   g05503(.A1(new_n5752_), .A2(new_n5452_), .ZN(new_n5753_));
  NAND2_X1   g05504(.A1(new_n3979_), .A2(new_n4201_), .ZN(new_n5754_));
  NOR2_X1    g05505(.A1(new_n800_), .A2(new_n2868_), .ZN(new_n5755_));
  INV_X1     g05506(.I(new_n5755_), .ZN(new_n5756_));
  NOR4_X1    g05507(.A1(new_n5754_), .A2(new_n1441_), .A3(new_n3981_), .A4(new_n5756_), .ZN(new_n5757_));
  XNOR2_X1   g05508(.A1(new_n5753_), .A2(new_n5757_), .ZN(new_n5758_));
  NOR2_X1    g05509(.A1(new_n5758_), .A2(new_n5749_), .ZN(new_n5759_));
  INV_X1     g05510(.I(new_n5753_), .ZN(new_n5760_));
  INV_X1     g05511(.I(new_n5757_), .ZN(new_n5761_));
  NOR2_X1    g05512(.A1(new_n5760_), .A2(new_n5761_), .ZN(new_n5762_));
  NOR2_X1    g05513(.A1(new_n5753_), .A2(new_n5757_), .ZN(new_n5763_));
  NOR2_X1    g05514(.A1(new_n5762_), .A2(new_n5763_), .ZN(new_n5764_));
  NOR2_X1    g05515(.A1(new_n5764_), .A2(new_n5748_), .ZN(new_n5765_));
  NOR2_X1    g05516(.A1(new_n5765_), .A2(new_n5759_), .ZN(new_n5766_));
  NOR3_X1    g05517(.A1(new_n1199_), .A2(new_n3423_), .A3(new_n4501_), .ZN(new_n5767_));
  NOR3_X1    g05518(.A1(new_n1199_), .A2(new_n3423_), .A3(new_n4501_), .ZN(new_n5771_));
  INV_X1     g05519(.I(new_n5771_), .ZN(new_n5772_));
  NAND2_X1   g05520(.A1(new_n5350_), .A2(new_n609_), .ZN(new_n5773_));
  XNOR2_X1   g05521(.A1(new_n5773_), .A2(new_n3840_), .ZN(new_n5774_));
  NOR2_X1    g05522(.A1(new_n2368_), .A2(new_n1916_), .ZN(new_n5775_));
  NAND2_X1   g05523(.A1(new_n5775_), .A2(new_n2277_), .ZN(new_n5776_));
  XOR2_X1    g05524(.A1(new_n5776_), .A2(\a[11] ), .Z(new_n5777_));
  XOR2_X1    g05525(.A1(new_n5777_), .A2(\a[38] ), .Z(new_n5778_));
  NOR2_X1    g05526(.A1(new_n5778_), .A2(new_n5774_), .ZN(new_n5779_));
  INV_X1     g05527(.I(new_n5779_), .ZN(new_n5780_));
  NAND2_X1   g05528(.A1(new_n5778_), .A2(new_n5774_), .ZN(new_n5781_));
  AOI21_X1   g05529(.A1(new_n5780_), .A2(new_n5781_), .B(new_n5772_), .ZN(new_n5782_));
  XNOR2_X1   g05530(.A1(new_n5778_), .A2(new_n5774_), .ZN(new_n5783_));
  NOR2_X1    g05531(.A1(new_n5783_), .A2(new_n5771_), .ZN(new_n5784_));
  NOR2_X1    g05532(.A1(new_n5784_), .A2(new_n5782_), .ZN(new_n5785_));
  INV_X1     g05533(.I(new_n5601_), .ZN(new_n5786_));
  NOR2_X1    g05534(.A1(new_n5786_), .A2(new_n523_), .ZN(new_n5788_));
  NAND3_X1   g05535(.A1(new_n5788_), .A2(new_n5186_), .A3(new_n5291_), .ZN(new_n5789_));
  AOI21_X1   g05536(.A1(new_n5789_), .A2(new_n4321_), .B(new_n525_), .ZN(new_n5790_));
  NOR2_X1    g05537(.A1(new_n5786_), .A2(new_n523_), .ZN(new_n5791_));
  INV_X1     g05538(.I(new_n5791_), .ZN(new_n5792_));
  NAND2_X1   g05539(.A1(\a[46] ), .A2(\a[47] ), .ZN(new_n5793_));
  NOR2_X1    g05540(.A1(new_n225_), .A2(new_n5793_), .ZN(new_n5794_));
  XOR2_X1    g05541(.A1(new_n5794_), .A2(new_n2532_), .Z(new_n5795_));
  AOI22_X1   g05542(.A1(new_n1769_), .A2(new_n2898_), .B1(new_n3354_), .B2(new_n1798_), .ZN(new_n5796_));
  NOR4_X1    g05543(.A1(new_n2978_), .A2(new_n2690_), .A3(new_n1339_), .A4(new_n2461_), .ZN(new_n5797_));
  NAND2_X1   g05544(.A1(new_n5796_), .A2(new_n5797_), .ZN(new_n5798_));
  NOR2_X1    g05545(.A1(new_n5795_), .A2(new_n5798_), .ZN(new_n5799_));
  INV_X1     g05546(.I(new_n5799_), .ZN(new_n5800_));
  NAND2_X1   g05547(.A1(new_n5795_), .A2(new_n5798_), .ZN(new_n5801_));
  AOI21_X1   g05548(.A1(new_n5800_), .A2(new_n5801_), .B(new_n5792_), .ZN(new_n5802_));
  XNOR2_X1   g05549(.A1(new_n5795_), .A2(new_n5798_), .ZN(new_n5803_));
  NOR2_X1    g05550(.A1(new_n5803_), .A2(new_n5791_), .ZN(new_n5804_));
  NOR2_X1    g05551(.A1(new_n5804_), .A2(new_n5802_), .ZN(new_n5805_));
  NOR2_X1    g05552(.A1(new_n5785_), .A2(new_n5805_), .ZN(new_n5806_));
  INV_X1     g05553(.I(new_n5785_), .ZN(new_n5807_));
  INV_X1     g05554(.I(new_n5805_), .ZN(new_n5808_));
  NOR2_X1    g05555(.A1(new_n5807_), .A2(new_n5808_), .ZN(new_n5809_));
  NOR2_X1    g05556(.A1(new_n5809_), .A2(new_n5806_), .ZN(new_n5810_));
  NOR2_X1    g05557(.A1(new_n5810_), .A2(new_n5766_), .ZN(new_n5811_));
  INV_X1     g05558(.I(new_n5766_), .ZN(new_n5812_));
  XOR2_X1    g05559(.A1(new_n5785_), .A2(new_n5808_), .Z(new_n5813_));
  NOR2_X1    g05560(.A1(new_n5813_), .A2(new_n5812_), .ZN(new_n5814_));
  NOR2_X1    g05561(.A1(new_n5811_), .A2(new_n5814_), .ZN(new_n5815_));
  XNOR2_X1   g05562(.A1(new_n5815_), .A2(new_n5739_), .ZN(new_n5816_));
  INV_X1     g05563(.I(new_n5816_), .ZN(new_n5817_));
  NOR2_X1    g05564(.A1(new_n5815_), .A2(new_n5739_), .ZN(new_n5818_));
  INV_X1     g05565(.I(new_n5818_), .ZN(new_n5819_));
  NAND2_X1   g05566(.A1(new_n5815_), .A2(new_n5739_), .ZN(new_n5820_));
  AOI21_X1   g05567(.A1(new_n5819_), .A2(new_n5820_), .B(new_n5737_), .ZN(new_n5821_));
  AOI21_X1   g05568(.A1(new_n5817_), .A2(new_n5737_), .B(new_n5821_), .ZN(new_n5822_));
  XOR2_X1    g05569(.A1(new_n5736_), .A2(new_n5822_), .Z(new_n5823_));
  NOR2_X1    g05570(.A1(new_n5823_), .A2(new_n5645_), .ZN(new_n5824_));
  XNOR2_X1   g05571(.A1(new_n5736_), .A2(new_n5822_), .ZN(new_n5825_));
  INV_X1     g05572(.I(new_n5825_), .ZN(new_n5826_));
  AOI21_X1   g05573(.A1(new_n5645_), .A2(new_n5826_), .B(new_n5824_), .ZN(new_n5827_));
  OAI21_X1   g05574(.A1(new_n5439_), .A2(new_n5632_), .B(new_n5633_), .ZN(new_n5828_));
  XNOR2_X1   g05575(.A1(new_n5827_), .A2(new_n5828_), .ZN(new_n5829_));
  XNOR2_X1   g05576(.A1(new_n5827_), .A2(new_n5828_), .ZN(new_n5830_));
  NAND2_X1   g05577(.A1(new_n5644_), .A2(new_n5830_), .ZN(new_n5831_));
  OAI21_X1   g05578(.A1(new_n5644_), .A2(new_n5829_), .B(new_n5831_), .ZN(\asquared[50] ));
  NOR2_X1    g05579(.A1(new_n5827_), .A2(new_n5828_), .ZN(new_n5833_));
  NAND4_X1   g05580(.A1(new_n5636_), .A2(new_n5638_), .A3(new_n5827_), .A4(new_n5828_), .ZN(new_n5834_));
  NAND3_X1   g05581(.A1(new_n5436_), .A2(new_n5434_), .A3(new_n5834_), .ZN(new_n5835_));
  AND3_X2    g05582(.A1(new_n5835_), .A2(new_n5639_), .A3(new_n5833_), .Z(\asquared[51] ));
  NAND2_X1   g05583(.A1(new_n5724_), .A2(new_n5717_), .ZN(new_n5837_));
  NAND2_X1   g05584(.A1(new_n5837_), .A2(new_n5723_), .ZN(new_n5838_));
  INV_X1     g05585(.I(new_n5838_), .ZN(new_n5839_));
  NOR3_X1    g05586(.A1(new_n5562_), .A2(new_n3423_), .A3(new_n5004_), .ZN(new_n5840_));
  NOR2_X1    g05587(.A1(new_n800_), .A2(new_n5004_), .ZN(new_n5841_));
  NAND4_X1   g05588(.A1(new_n5840_), .A2(\a[5] ), .A3(\a[34] ), .A4(new_n5841_), .ZN(new_n5842_));
  AOI21_X1   g05589(.A1(new_n5842_), .A2(new_n3712_), .B(new_n1021_), .ZN(new_n5843_));
  NAND2_X1   g05590(.A1(\a[16] ), .A2(\a[34] ), .ZN(new_n5844_));
  NOR2_X1    g05591(.A1(new_n5843_), .A2(new_n5840_), .ZN(new_n5845_));
  INV_X1     g05592(.I(new_n5845_), .ZN(new_n5846_));
  NOR2_X1    g05593(.A1(new_n3423_), .A2(new_n5004_), .ZN(new_n5847_));
  NOR2_X1    g05594(.A1(new_n5246_), .A2(new_n5847_), .ZN(new_n5848_));
  INV_X1     g05595(.I(new_n5848_), .ZN(new_n5849_));
  OAI22_X1   g05596(.A1(new_n5846_), .A2(new_n5849_), .B1(new_n5843_), .B2(new_n5844_), .ZN(new_n5850_));
  NOR2_X1    g05597(.A1(new_n2368_), .A2(new_n2765_), .ZN(new_n5851_));
  INV_X1     g05598(.I(new_n5851_), .ZN(new_n5852_));
  NOR2_X1    g05599(.A1(new_n4989_), .A2(new_n5852_), .ZN(new_n5853_));
  NOR3_X1    g05600(.A1(new_n1676_), .A2(new_n2178_), .A3(new_n2765_), .ZN(new_n5854_));
  NAND2_X1   g05601(.A1(new_n5854_), .A2(new_n5853_), .ZN(new_n5855_));
  AOI21_X1   g05602(.A1(new_n5855_), .A2(new_n2692_), .B(new_n2285_), .ZN(new_n5856_));
  NOR3_X1    g05603(.A1(new_n5856_), .A2(new_n1674_), .A3(new_n2178_), .ZN(new_n5857_));
  NOR2_X1    g05604(.A1(new_n5856_), .A2(new_n5853_), .ZN(new_n5858_));
  INV_X1     g05605(.I(new_n5858_), .ZN(new_n5859_));
  OAI21_X1   g05606(.A1(new_n1276_), .A2(new_n2368_), .B(new_n3504_), .ZN(new_n5860_));
  NOR2_X1    g05607(.A1(new_n5859_), .A2(new_n5860_), .ZN(new_n5861_));
  NOR2_X1    g05608(.A1(new_n5861_), .A2(new_n5857_), .ZN(new_n5862_));
  OAI21_X1   g05609(.A1(new_n5684_), .A2(new_n5688_), .B(new_n5689_), .ZN(new_n5863_));
  INV_X1     g05610(.I(new_n5863_), .ZN(new_n5864_));
  XOR2_X1    g05611(.A1(new_n5862_), .A2(new_n5864_), .Z(new_n5865_));
  NOR3_X1    g05612(.A1(new_n5861_), .A2(new_n5857_), .A3(new_n5864_), .ZN(new_n5866_));
  NOR2_X1    g05613(.A1(new_n5862_), .A2(new_n5863_), .ZN(new_n5867_));
  OAI21_X1   g05614(.A1(new_n5867_), .A2(new_n5866_), .B(new_n5850_), .ZN(new_n5868_));
  OAI21_X1   g05615(.A1(new_n5865_), .A2(new_n5850_), .B(new_n5868_), .ZN(new_n5869_));
  NOR2_X1    g05616(.A1(new_n650_), .A2(new_n4501_), .ZN(new_n5870_));
  NOR3_X1    g05617(.A1(new_n1199_), .A2(new_n3393_), .A3(new_n4770_), .ZN(new_n5871_));
  NAND3_X1   g05618(.A1(new_n5871_), .A2(new_n4531_), .A3(new_n5870_), .ZN(new_n5872_));
  AOI21_X1   g05619(.A1(new_n5872_), .A2(new_n5322_), .B(new_n478_), .ZN(new_n5873_));
  NAND2_X1   g05620(.A1(\a[6] ), .A2(\a[44] ), .ZN(new_n5874_));
  NAND2_X1   g05621(.A1(new_n4531_), .A2(new_n5870_), .ZN(new_n5875_));
  OAI21_X1   g05622(.A1(new_n478_), .A2(new_n5322_), .B(new_n5875_), .ZN(new_n5876_));
  NAND2_X1   g05623(.A1(\a[36] ), .A2(\a[43] ), .ZN(new_n5877_));
  OAI21_X1   g05624(.A1(new_n268_), .A2(new_n650_), .B(new_n5877_), .ZN(new_n5878_));
  OAI22_X1   g05625(.A1(new_n5873_), .A2(new_n5874_), .B1(new_n5876_), .B2(new_n5878_), .ZN(new_n5879_));
  INV_X1     g05626(.I(new_n5879_), .ZN(new_n5880_));
  INV_X1     g05627(.I(new_n5350_), .ZN(new_n5881_));
  NOR2_X1    g05628(.A1(new_n3837_), .A2(new_n4414_), .ZN(new_n5882_));
  INV_X1     g05629(.I(new_n5882_), .ZN(new_n5883_));
  NOR2_X1    g05630(.A1(new_n5883_), .A2(new_n596_), .ZN(new_n5884_));
  NOR4_X1    g05631(.A1(new_n359_), .A2(new_n599_), .A3(new_n3837_), .A4(new_n4769_), .ZN(new_n5885_));
  NAND2_X1   g05632(.A1(new_n5884_), .A2(new_n5885_), .ZN(new_n5886_));
  AOI21_X1   g05633(.A1(new_n5886_), .A2(new_n5881_), .B(new_n453_), .ZN(new_n5887_));
  NOR3_X1    g05634(.A1(new_n5887_), .A2(new_n359_), .A3(new_n4769_), .ZN(new_n5888_));
  OAI22_X1   g05635(.A1(new_n453_), .A2(new_n5881_), .B1(new_n5883_), .B2(new_n596_), .ZN(new_n5889_));
  NAND2_X1   g05636(.A1(new_n5883_), .A2(new_n596_), .ZN(new_n5890_));
  NOR2_X1    g05637(.A1(new_n5889_), .A2(new_n5890_), .ZN(new_n5891_));
  NOR2_X1    g05638(.A1(new_n5888_), .A2(new_n5891_), .ZN(new_n5892_));
  INV_X1     g05639(.I(new_n5892_), .ZN(new_n5893_));
  AOI22_X1   g05640(.A1(new_n1479_), .A2(new_n5339_), .B1(new_n4241_), .B2(new_n3061_), .ZN(new_n5894_));
  NOR2_X1    g05641(.A1(new_n566_), .A2(new_n3804_), .ZN(new_n5895_));
  NAND4_X1   g05642(.A1(new_n5894_), .A2(new_n796_), .A3(new_n4321_), .A4(new_n5895_), .ZN(new_n5896_));
  NOR2_X1    g05643(.A1(new_n5893_), .A2(new_n5896_), .ZN(new_n5897_));
  INV_X1     g05644(.I(new_n5896_), .ZN(new_n5898_));
  NOR2_X1    g05645(.A1(new_n5892_), .A2(new_n5898_), .ZN(new_n5899_));
  OAI21_X1   g05646(.A1(new_n5897_), .A2(new_n5899_), .B(new_n5880_), .ZN(new_n5900_));
  XOR2_X1    g05647(.A1(new_n5892_), .A2(new_n5896_), .Z(new_n5901_));
  OAI21_X1   g05648(.A1(new_n5880_), .A2(new_n5901_), .B(new_n5900_), .ZN(new_n5902_));
  NAND2_X1   g05649(.A1(\a[48] ), .A2(\a[50] ), .ZN(new_n5903_));
  XNOR2_X1   g05650(.A1(new_n197_), .A2(new_n5903_), .ZN(new_n5904_));
  INV_X1     g05651(.I(new_n5904_), .ZN(new_n5905_));
  NAND2_X1   g05652(.A1(\a[3] ), .A2(\a[33] ), .ZN(new_n5906_));
  NAND2_X1   g05653(.A1(\a[17] ), .A2(\a[47] ), .ZN(new_n5907_));
  OAI22_X1   g05654(.A1(new_n212_), .A2(new_n5907_), .B1(new_n5906_), .B2(new_n5793_), .ZN(new_n5908_));
  NOR2_X1    g05655(.A1(new_n2868_), .A2(new_n5175_), .ZN(new_n5909_));
  INV_X1     g05656(.I(new_n5909_), .ZN(new_n5910_));
  NAND4_X1   g05657(.A1(new_n5910_), .A2(\a[3] ), .A3(\a[47] ), .A4(new_n1354_), .ZN(new_n5911_));
  AOI22_X1   g05658(.A1(new_n1769_), .A2(new_n3126_), .B1(new_n3733_), .B2(new_n1798_), .ZN(new_n5912_));
  INV_X1     g05659(.I(new_n5912_), .ZN(new_n5913_));
  NAND4_X1   g05660(.A1(new_n3175_), .A2(\a[19] ), .A3(\a[31] ), .A4(new_n1711_), .ZN(new_n5914_));
  NOR4_X1    g05661(.A1(new_n5913_), .A2(new_n5908_), .A3(new_n5911_), .A4(new_n5914_), .ZN(new_n5915_));
  NOR2_X1    g05662(.A1(new_n5911_), .A2(new_n5908_), .ZN(new_n5916_));
  NOR2_X1    g05663(.A1(new_n5913_), .A2(new_n5914_), .ZN(new_n5917_));
  NOR2_X1    g05664(.A1(new_n5917_), .A2(new_n5916_), .ZN(new_n5918_));
  OAI21_X1   g05665(.A1(new_n5918_), .A2(new_n5915_), .B(new_n5905_), .ZN(new_n5919_));
  XOR2_X1    g05666(.A1(new_n5917_), .A2(new_n5916_), .Z(new_n5920_));
  NAND2_X1   g05667(.A1(new_n5920_), .A2(new_n5904_), .ZN(new_n5921_));
  NAND2_X1   g05668(.A1(new_n5921_), .A2(new_n5919_), .ZN(new_n5922_));
  AND2_X2    g05669(.A1(new_n5902_), .A2(new_n5922_), .Z(new_n5923_));
  NOR2_X1    g05670(.A1(new_n5902_), .A2(new_n5922_), .ZN(new_n5924_));
  OAI21_X1   g05671(.A1(new_n5923_), .A2(new_n5924_), .B(new_n5869_), .ZN(new_n5925_));
  XNOR2_X1   g05672(.A1(new_n5902_), .A2(new_n5922_), .ZN(new_n5926_));
  OAI21_X1   g05673(.A1(new_n5869_), .A2(new_n5926_), .B(new_n5925_), .ZN(new_n5927_));
  NOR2_X1    g05674(.A1(new_n5839_), .A2(new_n5927_), .ZN(new_n5928_));
  OAI21_X1   g05675(.A1(new_n5669_), .A2(new_n5700_), .B(new_n5701_), .ZN(new_n5929_));
  NAND2_X1   g05676(.A1(new_n5839_), .A2(new_n5927_), .ZN(new_n5930_));
  AOI21_X1   g05677(.A1(new_n5929_), .A2(new_n5930_), .B(new_n5928_), .ZN(new_n5931_));
  NAND2_X1   g05678(.A1(new_n5781_), .A2(new_n5771_), .ZN(new_n5932_));
  NAND2_X1   g05679(.A1(new_n5350_), .A2(new_n609_), .ZN(new_n5933_));
  NOR2_X1    g05680(.A1(new_n5350_), .A2(new_n609_), .ZN(new_n5934_));
  NOR2_X1    g05681(.A1(\a[13] ), .A2(\a[36] ), .ZN(new_n5935_));
  AOI21_X1   g05682(.A1(new_n5933_), .A2(new_n5935_), .B(new_n5934_), .ZN(new_n5936_));
  INV_X1     g05683(.I(new_n5936_), .ZN(new_n5937_));
  AOI21_X1   g05684(.A1(new_n2978_), .A2(new_n2690_), .B(new_n5796_), .ZN(new_n5938_));
  OAI21_X1   g05685(.A1(new_n1268_), .A2(new_n4184_), .B(new_n5754_), .ZN(new_n5939_));
  XOR2_X1    g05686(.A1(new_n5939_), .A2(new_n5938_), .Z(new_n5940_));
  NOR2_X1    g05687(.A1(new_n5940_), .A2(new_n5937_), .ZN(new_n5941_));
  INV_X1     g05688(.I(new_n5938_), .ZN(new_n5942_));
  NOR2_X1    g05689(.A1(new_n5942_), .A2(new_n5939_), .ZN(new_n5943_));
  INV_X1     g05690(.I(new_n5943_), .ZN(new_n5944_));
  NAND2_X1   g05691(.A1(new_n5942_), .A2(new_n5939_), .ZN(new_n5945_));
  AOI21_X1   g05692(.A1(new_n5944_), .A2(new_n5945_), .B(new_n5936_), .ZN(new_n5946_));
  NOR2_X1    g05693(.A1(new_n5941_), .A2(new_n5946_), .ZN(new_n5947_));
  INV_X1     g05694(.I(new_n5947_), .ZN(new_n5948_));
  AOI21_X1   g05695(.A1(new_n5780_), .A2(new_n5932_), .B(new_n5948_), .ZN(new_n5949_));
  NAND2_X1   g05696(.A1(new_n5715_), .A2(new_n5708_), .ZN(new_n5950_));
  NAND2_X1   g05697(.A1(new_n5950_), .A2(new_n5714_), .ZN(new_n5951_));
  INV_X1     g05698(.I(new_n5951_), .ZN(new_n5952_));
  NAND2_X1   g05699(.A1(new_n5932_), .A2(new_n5780_), .ZN(new_n5953_));
  NOR2_X1    g05700(.A1(new_n5953_), .A2(new_n5947_), .ZN(new_n5954_));
  NOR2_X1    g05701(.A1(new_n5952_), .A2(new_n5954_), .ZN(new_n5955_));
  NOR2_X1    g05702(.A1(new_n5955_), .A2(new_n5949_), .ZN(new_n5956_));
  NAND2_X1   g05703(.A1(new_n5801_), .A2(new_n5791_), .ZN(new_n5957_));
  NAND2_X1   g05704(.A1(new_n5957_), .A2(new_n5800_), .ZN(new_n5958_));
  INV_X1     g05705(.I(new_n5958_), .ZN(new_n5959_));
  NOR2_X1    g05706(.A1(new_n5790_), .A2(new_n5788_), .ZN(new_n5960_));
  INV_X1     g05707(.I(new_n5960_), .ZN(new_n5961_));
  NOR2_X1    g05708(.A1(new_n675_), .A2(new_n3804_), .ZN(new_n5962_));
  OAI21_X1   g05709(.A1(new_n2277_), .A2(new_n5775_), .B(new_n5962_), .ZN(new_n5963_));
  NAND2_X1   g05710(.A1(new_n5963_), .A2(new_n5776_), .ZN(new_n5964_));
  NAND2_X1   g05711(.A1(\a[1] ), .A2(\a[49] ), .ZN(new_n5965_));
  XNOR2_X1   g05712(.A1(new_n2679_), .A2(new_n5965_), .ZN(new_n5966_));
  XNOR2_X1   g05713(.A1(new_n5964_), .A2(new_n5966_), .ZN(new_n5967_));
  NOR2_X1    g05714(.A1(new_n5964_), .A2(new_n5966_), .ZN(new_n5968_));
  NAND2_X1   g05715(.A1(new_n5964_), .A2(new_n5966_), .ZN(new_n5969_));
  INV_X1     g05716(.I(new_n5969_), .ZN(new_n5970_));
  OAI21_X1   g05717(.A1(new_n5968_), .A2(new_n5970_), .B(new_n5961_), .ZN(new_n5971_));
  OAI21_X1   g05718(.A1(new_n5961_), .A2(new_n5967_), .B(new_n5971_), .ZN(new_n5972_));
  NOR2_X1    g05719(.A1(new_n5972_), .A2(new_n5959_), .ZN(new_n5973_));
  INV_X1     g05720(.I(new_n5763_), .ZN(new_n5974_));
  AOI21_X1   g05721(.A1(new_n5748_), .A2(new_n5974_), .B(new_n5762_), .ZN(new_n5975_));
  INV_X1     g05722(.I(new_n5975_), .ZN(new_n5976_));
  NAND2_X1   g05723(.A1(new_n5972_), .A2(new_n5959_), .ZN(new_n5977_));
  AOI21_X1   g05724(.A1(new_n5976_), .A2(new_n5977_), .B(new_n5973_), .ZN(new_n5978_));
  NAND3_X1   g05725(.A1(new_n229_), .A2(\a[44] ), .A3(\a[45] ), .ZN(new_n5979_));
  INV_X1     g05726(.I(new_n5793_), .ZN(new_n5980_));
  NAND2_X1   g05727(.A1(new_n1674_), .A2(new_n2098_), .ZN(new_n5981_));
  AOI21_X1   g05728(.A1(new_n232_), .A2(new_n5980_), .B(new_n5981_), .ZN(new_n5982_));
  AOI21_X1   g05729(.A1(new_n225_), .A2(new_n5793_), .B(new_n5982_), .ZN(new_n5983_));
  NAND2_X1   g05730(.A1(new_n5983_), .A2(new_n5979_), .ZN(new_n5984_));
  INV_X1     g05731(.I(new_n5984_), .ZN(new_n5985_));
  AOI21_X1   g05732(.A1(new_n1447_), .A2(new_n3487_), .B(new_n5767_), .ZN(new_n5986_));
  NOR2_X1    g05733(.A1(new_n5983_), .A2(new_n5979_), .ZN(new_n5987_));
  INV_X1     g05734(.I(new_n5987_), .ZN(new_n5988_));
  AOI21_X1   g05735(.A1(new_n5986_), .A2(new_n5988_), .B(new_n5985_), .ZN(new_n5989_));
  INV_X1     g05736(.I(new_n5989_), .ZN(new_n5990_));
  OAI21_X1   g05737(.A1(new_n5961_), .A2(new_n5968_), .B(new_n5969_), .ZN(new_n5991_));
  NOR2_X1    g05738(.A1(new_n5918_), .A2(new_n5904_), .ZN(new_n5992_));
  NOR2_X1    g05739(.A1(new_n5992_), .A2(new_n5915_), .ZN(new_n5993_));
  XNOR2_X1   g05740(.A1(new_n5991_), .A2(new_n5993_), .ZN(new_n5994_));
  NAND2_X1   g05741(.A1(new_n5994_), .A2(new_n5990_), .ZN(new_n5995_));
  INV_X1     g05742(.I(new_n5991_), .ZN(new_n5996_));
  NOR2_X1    g05743(.A1(new_n5996_), .A2(new_n5993_), .ZN(new_n5997_));
  NAND2_X1   g05744(.A1(new_n5996_), .A2(new_n5993_), .ZN(new_n5998_));
  INV_X1     g05745(.I(new_n5998_), .ZN(new_n5999_));
  OAI21_X1   g05746(.A1(new_n5999_), .A2(new_n5997_), .B(new_n5989_), .ZN(new_n6000_));
  NAND2_X1   g05747(.A1(new_n6000_), .A2(new_n5995_), .ZN(new_n6001_));
  XNOR2_X1   g05748(.A1(new_n6001_), .A2(new_n5978_), .ZN(new_n6002_));
  AND2_X2    g05749(.A1(new_n6001_), .A2(new_n5978_), .Z(new_n6003_));
  NOR2_X1    g05750(.A1(new_n6001_), .A2(new_n5978_), .ZN(new_n6004_));
  OAI21_X1   g05751(.A1(new_n6003_), .A2(new_n6004_), .B(new_n5956_), .ZN(new_n6005_));
  OAI21_X1   g05752(.A1(new_n6002_), .A2(new_n5956_), .B(new_n6005_), .ZN(new_n6006_));
  NOR2_X1    g05753(.A1(new_n5869_), .A2(new_n5924_), .ZN(new_n6007_));
  NOR2_X1    g05754(.A1(new_n6007_), .A2(new_n5923_), .ZN(new_n6008_));
  NOR2_X1    g05755(.A1(new_n5867_), .A2(new_n5850_), .ZN(new_n6009_));
  NOR2_X1    g05756(.A1(new_n6009_), .A2(new_n5866_), .ZN(new_n6010_));
  OAI21_X1   g05757(.A1(new_n5564_), .A2(new_n5678_), .B(new_n5677_), .ZN(new_n6011_));
  INV_X1     g05758(.I(new_n6011_), .ZN(new_n6012_));
  INV_X1     g05759(.I(new_n5986_), .ZN(new_n6013_));
  XNOR2_X1   g05760(.A1(new_n5983_), .A2(new_n5979_), .ZN(new_n6014_));
  NOR2_X1    g05761(.A1(new_n6014_), .A2(new_n6013_), .ZN(new_n6015_));
  AOI21_X1   g05762(.A1(new_n5988_), .A2(new_n5984_), .B(new_n5986_), .ZN(new_n6016_));
  NOR3_X1    g05763(.A1(new_n6012_), .A2(new_n6015_), .A3(new_n6016_), .ZN(new_n6017_));
  INV_X1     g05764(.I(new_n5657_), .ZN(new_n6018_));
  AOI21_X1   g05765(.A1(new_n5652_), .A2(new_n6018_), .B(new_n5656_), .ZN(new_n6019_));
  NOR2_X1    g05766(.A1(new_n6015_), .A2(new_n6016_), .ZN(new_n6020_));
  NOR2_X1    g05767(.A1(new_n6020_), .A2(new_n6011_), .ZN(new_n6021_));
  NOR2_X1    g05768(.A1(new_n6021_), .A2(new_n6019_), .ZN(new_n6022_));
  NOR2_X1    g05769(.A1(new_n6022_), .A2(new_n6017_), .ZN(new_n6023_));
  INV_X1     g05770(.I(new_n4321_), .ZN(new_n6024_));
  AOI21_X1   g05771(.A1(new_n797_), .A2(new_n6024_), .B(new_n5894_), .ZN(new_n6025_));
  INV_X1     g05772(.I(new_n6025_), .ZN(new_n6026_));
  NOR2_X1    g05773(.A1(new_n5511_), .A2(new_n5745_), .ZN(new_n6027_));
  NOR2_X1    g05774(.A1(new_n5750_), .A2(new_n5745_), .ZN(new_n6028_));
  AOI21_X1   g05775(.A1(new_n6027_), .A2(new_n6028_), .B(new_n1271_), .ZN(new_n6029_));
  NOR2_X1    g05776(.A1(new_n5511_), .A2(new_n5750_), .ZN(new_n6030_));
  NOR4_X1    g05777(.A1(new_n6030_), .A2(new_n267_), .A3(new_n201_), .A4(new_n5745_), .ZN(new_n6031_));
  NAND2_X1   g05778(.A1(new_n6029_), .A2(new_n6031_), .ZN(new_n6032_));
  NOR2_X1    g05779(.A1(new_n6026_), .A2(new_n6032_), .ZN(new_n6033_));
  AOI21_X1   g05780(.A1(new_n6029_), .A2(new_n6031_), .B(new_n6025_), .ZN(new_n6034_));
  NOR2_X1    g05781(.A1(new_n6033_), .A2(new_n6034_), .ZN(new_n6035_));
  NOR2_X1    g05782(.A1(new_n6035_), .A2(new_n5846_), .ZN(new_n6036_));
  XOR2_X1    g05783(.A1(new_n6025_), .A2(new_n6032_), .Z(new_n6037_));
  NOR2_X1    g05784(.A1(new_n6037_), .A2(new_n5845_), .ZN(new_n6038_));
  NOR2_X1    g05785(.A1(new_n6036_), .A2(new_n6038_), .ZN(new_n6039_));
  XOR2_X1    g05786(.A1(new_n6023_), .A2(new_n6039_), .Z(new_n6040_));
  INV_X1     g05787(.I(new_n6040_), .ZN(new_n6041_));
  NOR2_X1    g05788(.A1(new_n6023_), .A2(new_n6039_), .ZN(new_n6042_));
  NOR4_X1    g05789(.A1(new_n6022_), .A2(new_n6017_), .A3(new_n6036_), .A4(new_n6038_), .ZN(new_n6043_));
  OAI21_X1   g05790(.A1(new_n6042_), .A2(new_n6043_), .B(new_n6010_), .ZN(new_n6044_));
  OAI21_X1   g05791(.A1(new_n6041_), .A2(new_n6010_), .B(new_n6044_), .ZN(new_n6045_));
  INV_X1     g05792(.I(new_n5897_), .ZN(new_n6046_));
  OAI21_X1   g05793(.A1(new_n5879_), .A2(new_n5899_), .B(new_n6046_), .ZN(new_n6047_));
  XNOR2_X1   g05794(.A1(new_n5876_), .A2(new_n5889_), .ZN(new_n6048_));
  NOR2_X1    g05795(.A1(new_n5859_), .A2(new_n6048_), .ZN(new_n6049_));
  NOR2_X1    g05796(.A1(new_n5876_), .A2(new_n5889_), .ZN(new_n6050_));
  INV_X1     g05797(.I(new_n6050_), .ZN(new_n6051_));
  NAND2_X1   g05798(.A1(new_n5876_), .A2(new_n5889_), .ZN(new_n6052_));
  AOI21_X1   g05799(.A1(new_n6051_), .A2(new_n6052_), .B(new_n5858_), .ZN(new_n6053_));
  NOR2_X1    g05800(.A1(new_n6049_), .A2(new_n6053_), .ZN(new_n6054_));
  INV_X1     g05801(.I(\a[50] ), .ZN(new_n6055_));
  NOR2_X1    g05802(.A1(new_n5750_), .A2(new_n6055_), .ZN(new_n6056_));
  NOR3_X1    g05803(.A1(new_n194_), .A2(new_n1999_), .A3(new_n5750_), .ZN(new_n6057_));
  AOI21_X1   g05804(.A1(new_n6057_), .A2(new_n218_), .B(new_n6056_), .ZN(new_n6058_));
  INV_X1     g05805(.I(new_n6058_), .ZN(new_n6059_));
  INV_X1     g05806(.I(new_n1354_), .ZN(new_n6060_));
  NAND2_X1   g05807(.A1(new_n5909_), .A2(new_n6060_), .ZN(new_n6061_));
  NAND2_X1   g05808(.A1(new_n6061_), .A2(new_n5908_), .ZN(new_n6062_));
  INV_X1     g05809(.I(new_n6062_), .ZN(new_n6063_));
  AOI21_X1   g05810(.A1(new_n2978_), .A2(new_n2898_), .B(new_n5912_), .ZN(new_n6064_));
  XOR2_X1    g05811(.A1(new_n6064_), .A2(new_n6063_), .Z(new_n6065_));
  NAND2_X1   g05812(.A1(new_n6065_), .A2(new_n6059_), .ZN(new_n6066_));
  AND2_X2    g05813(.A1(new_n6064_), .A2(new_n6063_), .Z(new_n6067_));
  NOR2_X1    g05814(.A1(new_n6064_), .A2(new_n6063_), .ZN(new_n6068_));
  OAI21_X1   g05815(.A1(new_n6067_), .A2(new_n6068_), .B(new_n6058_), .ZN(new_n6069_));
  NAND2_X1   g05816(.A1(new_n6066_), .A2(new_n6069_), .ZN(new_n6070_));
  XNOR2_X1   g05817(.A1(new_n6054_), .A2(new_n6070_), .ZN(new_n6071_));
  AND2_X2    g05818(.A1(new_n6071_), .A2(new_n6047_), .Z(new_n6072_));
  OAI21_X1   g05819(.A1(new_n6049_), .A2(new_n6053_), .B(new_n6070_), .ZN(new_n6073_));
  NAND3_X1   g05820(.A1(new_n6054_), .A2(new_n6066_), .A3(new_n6069_), .ZN(new_n6074_));
  AOI21_X1   g05821(.A1(new_n6074_), .A2(new_n6073_), .B(new_n6047_), .ZN(new_n6075_));
  NOR2_X1    g05822(.A1(new_n6072_), .A2(new_n6075_), .ZN(new_n6076_));
  XOR2_X1    g05823(.A1(new_n6045_), .A2(new_n6076_), .Z(new_n6077_));
  INV_X1     g05824(.I(new_n6076_), .ZN(new_n6078_));
  NAND2_X1   g05825(.A1(new_n6045_), .A2(new_n6078_), .ZN(new_n6079_));
  INV_X1     g05826(.I(new_n6079_), .ZN(new_n6080_));
  NOR2_X1    g05827(.A1(new_n6045_), .A2(new_n6078_), .ZN(new_n6081_));
  OAI21_X1   g05828(.A1(new_n6080_), .A2(new_n6081_), .B(new_n6008_), .ZN(new_n6082_));
  OAI21_X1   g05829(.A1(new_n6008_), .A2(new_n6077_), .B(new_n6082_), .ZN(new_n6083_));
  XNOR2_X1   g05830(.A1(new_n6083_), .A2(new_n6006_), .ZN(new_n6084_));
  NOR2_X1    g05831(.A1(new_n6084_), .A2(new_n5931_), .ZN(new_n6085_));
  INV_X1     g05832(.I(new_n5931_), .ZN(new_n6086_));
  NAND2_X1   g05833(.A1(new_n6083_), .A2(new_n6006_), .ZN(new_n6087_));
  OR2_X2     g05834(.A1(new_n6083_), .A2(new_n6006_), .Z(new_n6088_));
  AOI21_X1   g05835(.A1(new_n6088_), .A2(new_n6087_), .B(new_n6086_), .ZN(new_n6089_));
  NOR2_X1    g05836(.A1(new_n6085_), .A2(new_n6089_), .ZN(new_n6090_));
  OAI21_X1   g05837(.A1(new_n5648_), .A2(new_n5664_), .B(new_n5666_), .ZN(new_n6091_));
  INV_X1     g05838(.I(new_n6091_), .ZN(new_n6092_));
  NAND2_X1   g05839(.A1(new_n5693_), .A2(new_n5681_), .ZN(new_n6093_));
  NAND2_X1   g05840(.A1(new_n6093_), .A2(new_n5695_), .ZN(new_n6094_));
  XOR2_X1    g05841(.A1(new_n6020_), .A2(new_n6012_), .Z(new_n6095_));
  OAI21_X1   g05842(.A1(new_n6021_), .A2(new_n6017_), .B(new_n6019_), .ZN(new_n6096_));
  OAI21_X1   g05843(.A1(new_n6095_), .A2(new_n6019_), .B(new_n6096_), .ZN(new_n6097_));
  XOR2_X1    g05844(.A1(new_n6097_), .A2(new_n6094_), .Z(new_n6098_));
  NOR2_X1    g05845(.A1(new_n6098_), .A2(new_n6092_), .ZN(new_n6099_));
  INV_X1     g05846(.I(new_n6097_), .ZN(new_n6100_));
  NOR2_X1    g05847(.A1(new_n6100_), .A2(new_n6094_), .ZN(new_n6101_));
  INV_X1     g05848(.I(new_n6101_), .ZN(new_n6102_));
  NAND2_X1   g05849(.A1(new_n6100_), .A2(new_n6094_), .ZN(new_n6103_));
  AOI21_X1   g05850(.A1(new_n6102_), .A2(new_n6103_), .B(new_n6091_), .ZN(new_n6104_));
  NOR2_X1    g05851(.A1(new_n6104_), .A2(new_n6099_), .ZN(new_n6105_));
  INV_X1     g05852(.I(new_n6105_), .ZN(new_n6106_));
  XOR2_X1    g05853(.A1(new_n5972_), .A2(new_n5958_), .Z(new_n6107_));
  NOR2_X1    g05854(.A1(new_n6107_), .A2(new_n5975_), .ZN(new_n6108_));
  INV_X1     g05855(.I(new_n5973_), .ZN(new_n6109_));
  AOI21_X1   g05856(.A1(new_n6109_), .A2(new_n5977_), .B(new_n5976_), .ZN(new_n6110_));
  NOR2_X1    g05857(.A1(new_n6108_), .A2(new_n6110_), .ZN(new_n6111_));
  INV_X1     g05858(.I(new_n6111_), .ZN(new_n6112_));
  XOR2_X1    g05859(.A1(new_n5953_), .A2(new_n5948_), .Z(new_n6113_));
  OAI21_X1   g05860(.A1(new_n5949_), .A2(new_n5954_), .B(new_n5952_), .ZN(new_n6114_));
  OAI21_X1   g05861(.A1(new_n5952_), .A2(new_n6113_), .B(new_n6114_), .ZN(new_n6115_));
  INV_X1     g05862(.I(new_n5806_), .ZN(new_n6116_));
  OAI21_X1   g05863(.A1(new_n5812_), .A2(new_n5809_), .B(new_n6116_), .ZN(new_n6117_));
  INV_X1     g05864(.I(new_n6117_), .ZN(new_n6118_));
  NOR2_X1    g05865(.A1(new_n6118_), .A2(new_n6115_), .ZN(new_n6119_));
  INV_X1     g05866(.I(new_n6115_), .ZN(new_n6120_));
  NOR2_X1    g05867(.A1(new_n6120_), .A2(new_n6117_), .ZN(new_n6121_));
  OAI21_X1   g05868(.A1(new_n6119_), .A2(new_n6121_), .B(new_n6112_), .ZN(new_n6122_));
  XOR2_X1    g05869(.A1(new_n6117_), .A2(new_n6115_), .Z(new_n6123_));
  OAI21_X1   g05870(.A1(new_n6112_), .A2(new_n6123_), .B(new_n6122_), .ZN(new_n6124_));
  NOR2_X1    g05871(.A1(new_n6124_), .A2(new_n6106_), .ZN(new_n6125_));
  INV_X1     g05872(.I(new_n5820_), .ZN(new_n6126_));
  AOI21_X1   g05873(.A1(new_n5737_), .A2(new_n5819_), .B(new_n6126_), .ZN(new_n6127_));
  INV_X1     g05874(.I(new_n6127_), .ZN(new_n6128_));
  NAND2_X1   g05875(.A1(new_n6124_), .A2(new_n6106_), .ZN(new_n6129_));
  AOI21_X1   g05876(.A1(new_n6128_), .A2(new_n6129_), .B(new_n6125_), .ZN(new_n6130_));
  INV_X1     g05877(.I(new_n6130_), .ZN(new_n6131_));
  OAI21_X1   g05878(.A1(new_n6092_), .A2(new_n6101_), .B(new_n6103_), .ZN(new_n6132_));
  INV_X1     g05879(.I(new_n6132_), .ZN(new_n6133_));
  NOR2_X1    g05880(.A1(new_n6121_), .A2(new_n6112_), .ZN(new_n6134_));
  NOR2_X1    g05881(.A1(new_n6134_), .A2(new_n6119_), .ZN(new_n6135_));
  NOR2_X1    g05882(.A1(new_n599_), .A2(new_n4501_), .ZN(new_n6136_));
  INV_X1     g05883(.I(new_n6136_), .ZN(new_n6137_));
  NOR3_X1    g05884(.A1(new_n6137_), .A2(new_n359_), .A3(new_n3804_), .ZN(new_n6138_));
  NOR4_X1    g05885(.A1(new_n268_), .A2(new_n599_), .A3(new_n3804_), .A4(new_n4770_), .ZN(new_n6139_));
  NAND2_X1   g05886(.A1(new_n6138_), .A2(new_n6139_), .ZN(new_n6140_));
  AOI21_X1   g05887(.A1(new_n6140_), .A2(new_n5322_), .B(new_n392_), .ZN(new_n6141_));
  NOR3_X1    g05888(.A1(new_n6141_), .A2(new_n268_), .A3(new_n4770_), .ZN(new_n6142_));
  NOR2_X1    g05889(.A1(new_n6141_), .A2(new_n6138_), .ZN(new_n6143_));
  AOI22_X1   g05890(.A1(\a[8] ), .A2(\a[13] ), .B1(\a[38] ), .B2(\a[43] ), .ZN(new_n6144_));
  AOI21_X1   g05891(.A1(new_n6143_), .A2(new_n6144_), .B(new_n6142_), .ZN(new_n6145_));
  INV_X1     g05892(.I(new_n4415_), .ZN(new_n6146_));
  NOR2_X1    g05893(.A1(new_n364_), .A2(new_n4769_), .ZN(new_n6147_));
  NOR2_X1    g05894(.A1(new_n6146_), .A2(new_n523_), .ZN(new_n6148_));
  NAND4_X1   g05895(.A1(new_n6148_), .A2(\a[12] ), .A3(new_n6147_), .A4(\a[39] ), .ZN(new_n6149_));
  AOI21_X1   g05896(.A1(new_n6149_), .A2(new_n5881_), .B(new_n525_), .ZN(new_n6150_));
  NOR2_X1    g05897(.A1(new_n6146_), .A2(new_n523_), .ZN(new_n6151_));
  INV_X1     g05898(.I(new_n6151_), .ZN(new_n6152_));
  NOR2_X1    g05899(.A1(new_n2534_), .A2(new_n2276_), .ZN(new_n6153_));
  INV_X1     g05900(.I(new_n6153_), .ZN(new_n6154_));
  AOI21_X1   g05901(.A1(\a[24] ), .A2(\a[27] ), .B(new_n2752_), .ZN(new_n6155_));
  INV_X1     g05902(.I(new_n6155_), .ZN(new_n6156_));
  NOR2_X1    g05903(.A1(new_n6154_), .A2(new_n6156_), .ZN(new_n6157_));
  NOR2_X1    g05904(.A1(new_n675_), .A2(new_n4240_), .ZN(new_n6158_));
  XNOR2_X1   g05905(.A1(new_n6157_), .A2(new_n6158_), .ZN(new_n6159_));
  NOR2_X1    g05906(.A1(new_n6159_), .A2(new_n6152_), .ZN(new_n6160_));
  INV_X1     g05907(.I(new_n6159_), .ZN(new_n6161_));
  NOR2_X1    g05908(.A1(new_n6161_), .A2(new_n6151_), .ZN(new_n6162_));
  OAI21_X1   g05909(.A1(new_n6162_), .A2(new_n6160_), .B(new_n6145_), .ZN(new_n6163_));
  XOR2_X1    g05910(.A1(new_n6159_), .A2(new_n6151_), .Z(new_n6164_));
  OAI21_X1   g05911(.A1(new_n6164_), .A2(new_n6145_), .B(new_n6163_), .ZN(new_n6165_));
  AOI21_X1   g05912(.A1(new_n5936_), .A2(new_n5945_), .B(new_n5943_), .ZN(new_n6166_));
  NOR2_X1    g05913(.A1(new_n2679_), .A2(new_n5965_), .ZN(new_n6167_));
  NOR2_X1    g05914(.A1(new_n194_), .A2(new_n6055_), .ZN(new_n6168_));
  NAND3_X1   g05915(.A1(\a[1] ), .A2(\a[26] ), .A3(\a[50] ), .ZN(new_n6169_));
  OAI21_X1   g05916(.A1(new_n6168_), .A2(\a[26] ), .B(new_n6169_), .ZN(new_n6170_));
  NAND2_X1   g05917(.A1(new_n6170_), .A2(new_n6167_), .ZN(new_n6171_));
  XOR2_X1    g05918(.A1(new_n6171_), .A2(\a[0] ), .Z(new_n6172_));
  XOR2_X1    g05919(.A1(new_n6172_), .A2(\a[51] ), .Z(new_n6173_));
  NAND2_X1   g05920(.A1(new_n3981_), .A2(new_n1798_), .ZN(new_n6174_));
  NOR2_X1    g05921(.A1(new_n885_), .A2(new_n3371_), .ZN(new_n6175_));
  XOR2_X1    g05922(.A1(new_n6174_), .A2(new_n6175_), .Z(new_n6176_));
  XNOR2_X1   g05923(.A1(new_n6173_), .A2(new_n6176_), .ZN(new_n6177_));
  NOR2_X1    g05924(.A1(new_n6173_), .A2(new_n6176_), .ZN(new_n6178_));
  NAND2_X1   g05925(.A1(new_n6173_), .A2(new_n6176_), .ZN(new_n6179_));
  INV_X1     g05926(.I(new_n6179_), .ZN(new_n6180_));
  OAI21_X1   g05927(.A1(new_n6180_), .A2(new_n6178_), .B(new_n6166_), .ZN(new_n6181_));
  OAI21_X1   g05928(.A1(new_n6166_), .A2(new_n6177_), .B(new_n6181_), .ZN(new_n6182_));
  NOR2_X1    g05929(.A1(new_n875_), .A2(new_n3393_), .ZN(new_n6183_));
  NOR3_X1    g05930(.A1(new_n1199_), .A2(new_n3837_), .A3(new_n5004_), .ZN(new_n6184_));
  NAND4_X1   g05931(.A1(new_n6184_), .A2(\a[6] ), .A3(\a[45] ), .A4(new_n6183_), .ZN(new_n6185_));
  AOI21_X1   g05932(.A1(new_n6185_), .A2(new_n3839_), .B(new_n1018_), .ZN(new_n6186_));
  NOR3_X1    g05933(.A1(new_n1199_), .A2(new_n3837_), .A3(new_n5004_), .ZN(new_n6187_));
  AOI22_X1   g05934(.A1(new_n1531_), .A2(new_n3424_), .B1(new_n5909_), .B2(new_n4200_), .ZN(new_n6188_));
  NOR2_X1    g05935(.A1(new_n353_), .A2(new_n5175_), .ZN(new_n6189_));
  NOR2_X1    g05936(.A1(new_n800_), .A2(new_n3423_), .ZN(new_n6190_));
  XNOR2_X1   g05937(.A1(new_n6189_), .A2(new_n6190_), .ZN(new_n6191_));
  OAI21_X1   g05938(.A1(new_n6191_), .A2(new_n6189_), .B(new_n6188_), .ZN(new_n6192_));
  OAI21_X1   g05939(.A1(new_n1276_), .A2(new_n2868_), .B(new_n6191_), .ZN(new_n6193_));
  NAND2_X1   g05940(.A1(new_n6193_), .A2(new_n6192_), .ZN(new_n6194_));
  NOR2_X1    g05941(.A1(new_n1706_), .A2(new_n1773_), .ZN(new_n6195_));
  NOR2_X1    g05942(.A1(new_n3356_), .A2(new_n6195_), .ZN(new_n6196_));
  NOR4_X1    g05943(.A1(new_n2286_), .A2(new_n2690_), .A3(new_n1313_), .A4(new_n2461_), .ZN(new_n6197_));
  NAND2_X1   g05944(.A1(new_n6196_), .A2(new_n6197_), .ZN(new_n6198_));
  NOR2_X1    g05945(.A1(new_n6194_), .A2(new_n6198_), .ZN(new_n6199_));
  INV_X1     g05946(.I(new_n6198_), .ZN(new_n6200_));
  AOI21_X1   g05947(.A1(new_n6193_), .A2(new_n6192_), .B(new_n6200_), .ZN(new_n6201_));
  OAI21_X1   g05948(.A1(new_n6201_), .A2(new_n6199_), .B(new_n6187_), .ZN(new_n6202_));
  XOR2_X1    g05949(.A1(new_n6194_), .A2(new_n6200_), .Z(new_n6203_));
  OAI21_X1   g05950(.A1(new_n6203_), .A2(new_n6187_), .B(new_n6202_), .ZN(new_n6204_));
  XOR2_X1    g05951(.A1(new_n6182_), .A2(new_n6204_), .Z(new_n6205_));
  INV_X1     g05952(.I(new_n6205_), .ZN(new_n6206_));
  INV_X1     g05953(.I(new_n6204_), .ZN(new_n6207_));
  NOR2_X1    g05954(.A1(new_n6182_), .A2(new_n6207_), .ZN(new_n6208_));
  INV_X1     g05955(.I(new_n6208_), .ZN(new_n6209_));
  NAND2_X1   g05956(.A1(new_n6182_), .A2(new_n6207_), .ZN(new_n6210_));
  AOI21_X1   g05957(.A1(new_n6209_), .A2(new_n6210_), .B(new_n6165_), .ZN(new_n6211_));
  AOI21_X1   g05958(.A1(new_n6206_), .A2(new_n6165_), .B(new_n6211_), .ZN(new_n6212_));
  XOR2_X1    g05959(.A1(new_n6135_), .A2(new_n6212_), .Z(new_n6213_));
  NOR2_X1    g05960(.A1(new_n6213_), .A2(new_n6133_), .ZN(new_n6214_));
  INV_X1     g05961(.I(new_n6135_), .ZN(new_n6215_));
  NOR2_X1    g05962(.A1(new_n6215_), .A2(new_n6212_), .ZN(new_n6216_));
  INV_X1     g05963(.I(new_n6216_), .ZN(new_n6217_));
  NAND2_X1   g05964(.A1(new_n6215_), .A2(new_n6212_), .ZN(new_n6218_));
  AOI21_X1   g05965(.A1(new_n6217_), .A2(new_n6218_), .B(new_n6132_), .ZN(new_n6219_));
  NOR2_X1    g05966(.A1(new_n6219_), .A2(new_n6214_), .ZN(new_n6220_));
  NOR2_X1    g05967(.A1(new_n6220_), .A2(new_n6131_), .ZN(new_n6221_));
  INV_X1     g05968(.I(new_n6221_), .ZN(new_n6222_));
  NAND2_X1   g05969(.A1(new_n6220_), .A2(new_n6131_), .ZN(new_n6223_));
  AOI21_X1   g05970(.A1(new_n6222_), .A2(new_n6223_), .B(new_n6090_), .ZN(new_n6224_));
  INV_X1     g05971(.I(new_n6090_), .ZN(new_n6225_));
  XOR2_X1    g05972(.A1(new_n6220_), .A2(new_n6130_), .Z(new_n6226_));
  NOR2_X1    g05973(.A1(new_n6225_), .A2(new_n6226_), .ZN(new_n6227_));
  NOR2_X1    g05974(.A1(new_n6227_), .A2(new_n6224_), .ZN(new_n6228_));
  XNOR2_X1   g05975(.A1(new_n5927_), .A2(new_n5838_), .ZN(new_n6229_));
  NAND2_X1   g05976(.A1(new_n6229_), .A2(new_n5929_), .ZN(new_n6230_));
  INV_X1     g05977(.I(new_n5930_), .ZN(new_n6231_));
  NOR2_X1    g05978(.A1(new_n6231_), .A2(new_n5928_), .ZN(new_n6232_));
  OAI21_X1   g05979(.A1(new_n5929_), .A2(new_n6232_), .B(new_n6230_), .ZN(new_n6233_));
  XOR2_X1    g05980(.A1(new_n6124_), .A2(new_n6105_), .Z(new_n6234_));
  INV_X1     g05981(.I(new_n6129_), .ZN(new_n6235_));
  OAI21_X1   g05982(.A1(new_n6235_), .A2(new_n6125_), .B(new_n6127_), .ZN(new_n6236_));
  OAI21_X1   g05983(.A1(new_n6127_), .A2(new_n6234_), .B(new_n6236_), .ZN(new_n6237_));
  NOR2_X1    g05984(.A1(new_n6237_), .A2(new_n6233_), .ZN(new_n6238_));
  INV_X1     g05985(.I(new_n5734_), .ZN(new_n6239_));
  OAI21_X1   g05986(.A1(new_n5646_), .A2(new_n5732_), .B(new_n6239_), .ZN(new_n6240_));
  NAND2_X1   g05987(.A1(new_n6237_), .A2(new_n6233_), .ZN(new_n6241_));
  AOI21_X1   g05988(.A1(new_n6240_), .A2(new_n6241_), .B(new_n6238_), .ZN(new_n6242_));
  XNOR2_X1   g05989(.A1(new_n6228_), .A2(new_n6242_), .ZN(new_n6243_));
  NAND2_X1   g05990(.A1(\asquared[51] ), .A2(new_n6243_), .ZN(new_n6244_));
  XNOR2_X1   g05991(.A1(new_n6228_), .A2(new_n6242_), .ZN(new_n6245_));
  OAI21_X1   g05992(.A1(\asquared[51] ), .A2(new_n6245_), .B(new_n6244_), .ZN(\asquared[52] ));
  INV_X1     g05993(.I(new_n6228_), .ZN(new_n6247_));
  NOR2_X1    g05994(.A1(new_n6247_), .A2(new_n6242_), .ZN(new_n6248_));
  NAND2_X1   g05995(.A1(new_n6247_), .A2(new_n6242_), .ZN(new_n6249_));
  AOI21_X1   g05996(.A1(\asquared[51] ), .A2(new_n6249_), .B(new_n6248_), .ZN(new_n6250_));
  OAI21_X1   g05997(.A1(new_n6133_), .A2(new_n6216_), .B(new_n6218_), .ZN(new_n6251_));
  INV_X1     g05998(.I(new_n6042_), .ZN(new_n6252_));
  OAI21_X1   g05999(.A1(new_n6010_), .A2(new_n6043_), .B(new_n6252_), .ZN(new_n6253_));
  INV_X1     g06000(.I(new_n6162_), .ZN(new_n6254_));
  AOI21_X1   g06001(.A1(new_n6254_), .A2(new_n6145_), .B(new_n6160_), .ZN(new_n6255_));
  INV_X1     g06002(.I(new_n6034_), .ZN(new_n6256_));
  AOI21_X1   g06003(.A1(new_n6256_), .A2(new_n5845_), .B(new_n6033_), .ZN(new_n6257_));
  NOR2_X1    g06004(.A1(\a[11] ), .A2(\a[40] ), .ZN(new_n6258_));
  AOI21_X1   g06005(.A1(new_n6154_), .A2(new_n6258_), .B(new_n6156_), .ZN(new_n6259_));
  INV_X1     g06006(.I(\a[51] ), .ZN(new_n6260_));
  NOR2_X1    g06007(.A1(new_n194_), .A2(new_n6260_), .ZN(new_n6261_));
  XNOR2_X1   g06008(.A1(new_n2890_), .A2(new_n6261_), .ZN(new_n6262_));
  XOR2_X1    g06009(.A1(new_n6262_), .A2(new_n6169_), .Z(new_n6263_));
  NAND2_X1   g06010(.A1(new_n6263_), .A2(new_n6259_), .ZN(new_n6264_));
  INV_X1     g06011(.I(new_n6259_), .ZN(new_n6265_));
  NOR2_X1    g06012(.A1(new_n6262_), .A2(new_n6169_), .ZN(new_n6266_));
  NAND2_X1   g06013(.A1(new_n6262_), .A2(new_n6169_), .ZN(new_n6267_));
  INV_X1     g06014(.I(new_n6267_), .ZN(new_n6268_));
  OAI21_X1   g06015(.A1(new_n6268_), .A2(new_n6266_), .B(new_n6265_), .ZN(new_n6269_));
  NAND2_X1   g06016(.A1(new_n6264_), .A2(new_n6269_), .ZN(new_n6270_));
  XNOR2_X1   g06017(.A1(new_n6270_), .A2(new_n6257_), .ZN(new_n6271_));
  AND2_X2    g06018(.A1(new_n6270_), .A2(new_n6257_), .Z(new_n6272_));
  NOR2_X1    g06019(.A1(new_n6270_), .A2(new_n6257_), .ZN(new_n6273_));
  OAI21_X1   g06020(.A1(new_n6272_), .A2(new_n6273_), .B(new_n6255_), .ZN(new_n6274_));
  OAI21_X1   g06021(.A1(new_n6255_), .A2(new_n6271_), .B(new_n6274_), .ZN(new_n6275_));
  AOI21_X1   g06022(.A1(new_n5858_), .A2(new_n6052_), .B(new_n6050_), .ZN(new_n6276_));
  INV_X1     g06023(.I(new_n6276_), .ZN(new_n6277_));
  NOR2_X1    g06024(.A1(new_n6068_), .A2(new_n6058_), .ZN(new_n6278_));
  NOR2_X1    g06025(.A1(new_n6278_), .A2(new_n6067_), .ZN(new_n6279_));
  NOR2_X1    g06026(.A1(new_n5745_), .A2(new_n6055_), .ZN(new_n6280_));
  NAND2_X1   g06027(.A1(new_n6280_), .A2(new_n232_), .ZN(new_n6281_));
  NAND2_X1   g06028(.A1(\a[19] ), .A2(\a[33] ), .ZN(new_n6282_));
  XNOR2_X1   g06029(.A1(new_n6281_), .A2(new_n6282_), .ZN(new_n6283_));
  XOR2_X1    g06030(.A1(new_n6279_), .A2(new_n6283_), .Z(new_n6284_));
  NOR2_X1    g06031(.A1(new_n6279_), .A2(new_n6283_), .ZN(new_n6285_));
  INV_X1     g06032(.I(new_n6285_), .ZN(new_n6286_));
  NAND2_X1   g06033(.A1(new_n6279_), .A2(new_n6283_), .ZN(new_n6287_));
  AOI21_X1   g06034(.A1(new_n6286_), .A2(new_n6287_), .B(new_n6277_), .ZN(new_n6288_));
  AOI21_X1   g06035(.A1(new_n6277_), .A2(new_n6284_), .B(new_n6288_), .ZN(new_n6289_));
  XOR2_X1    g06036(.A1(new_n6275_), .A2(new_n6289_), .Z(new_n6290_));
  INV_X1     g06037(.I(new_n6290_), .ZN(new_n6291_));
  INV_X1     g06038(.I(new_n6275_), .ZN(new_n6292_));
  NOR2_X1    g06039(.A1(new_n6292_), .A2(new_n6289_), .ZN(new_n6293_));
  INV_X1     g06040(.I(new_n6293_), .ZN(new_n6294_));
  NAND2_X1   g06041(.A1(new_n6292_), .A2(new_n6289_), .ZN(new_n6295_));
  AOI21_X1   g06042(.A1(new_n6294_), .A2(new_n6295_), .B(new_n6253_), .ZN(new_n6296_));
  AOI21_X1   g06043(.A1(new_n6253_), .A2(new_n6291_), .B(new_n6296_), .ZN(new_n6297_));
  AOI21_X1   g06044(.A1(new_n5990_), .A2(new_n5998_), .B(new_n5997_), .ZN(new_n6298_));
  INV_X1     g06045(.I(new_n6298_), .ZN(new_n6299_));
  NOR2_X1    g06046(.A1(new_n6150_), .A2(new_n6148_), .ZN(new_n6300_));
  NOR2_X1    g06047(.A1(new_n3423_), .A2(new_n5750_), .ZN(new_n6301_));
  AOI21_X1   g06048(.A1(new_n3123_), .A2(new_n886_), .B(new_n6301_), .ZN(new_n6302_));
  NOR2_X1    g06049(.A1(\a[0] ), .A2(\a[52] ), .ZN(new_n6303_));
  NOR3_X1    g06050(.A1(new_n1354_), .A2(new_n3423_), .A3(new_n5750_), .ZN(new_n6304_));
  INV_X1     g06051(.I(new_n6304_), .ZN(new_n6305_));
  NOR3_X1    g06052(.A1(new_n6302_), .A2(new_n6303_), .A3(new_n6305_), .ZN(new_n6306_));
  NAND2_X1   g06053(.A1(new_n6302_), .A2(\a[52] ), .ZN(new_n6307_));
  NAND2_X1   g06054(.A1(new_n6307_), .A2(new_n6305_), .ZN(new_n6308_));
  NOR3_X1    g06055(.A1(new_n6308_), .A2(new_n6060_), .A3(new_n6301_), .ZN(new_n6309_));
  NOR2_X1    g06056(.A1(new_n6309_), .A2(new_n6306_), .ZN(new_n6310_));
  INV_X1     g06057(.I(new_n6310_), .ZN(new_n6311_));
  NOR2_X1    g06058(.A1(new_n199_), .A2(new_n6260_), .ZN(new_n6312_));
  OAI21_X1   g06059(.A1(new_n6170_), .A2(new_n6167_), .B(new_n6312_), .ZN(new_n6313_));
  NAND2_X1   g06060(.A1(new_n6313_), .A2(new_n6171_), .ZN(new_n6314_));
  INV_X1     g06061(.I(new_n6314_), .ZN(new_n6315_));
  NOR2_X1    g06062(.A1(new_n6311_), .A2(new_n6315_), .ZN(new_n6316_));
  NOR2_X1    g06063(.A1(new_n6310_), .A2(new_n6314_), .ZN(new_n6317_));
  NOR2_X1    g06064(.A1(new_n6316_), .A2(new_n6317_), .ZN(new_n6318_));
  XOR2_X1    g06065(.A1(new_n6310_), .A2(new_n6315_), .Z(new_n6319_));
  MUX2_X1    g06066(.I0(new_n6319_), .I1(new_n6318_), .S(new_n6300_), .Z(new_n6320_));
  NOR2_X1    g06067(.A1(new_n6180_), .A2(new_n6166_), .ZN(new_n6321_));
  NOR2_X1    g06068(.A1(new_n6321_), .A2(new_n6178_), .ZN(new_n6322_));
  XOR2_X1    g06069(.A1(new_n6322_), .A2(new_n6320_), .Z(new_n6323_));
  NAND2_X1   g06070(.A1(new_n6323_), .A2(new_n6299_), .ZN(new_n6324_));
  NOR2_X1    g06071(.A1(new_n6322_), .A2(new_n6320_), .ZN(new_n6325_));
  NAND2_X1   g06072(.A1(new_n6322_), .A2(new_n6320_), .ZN(new_n6326_));
  INV_X1     g06073(.I(new_n6326_), .ZN(new_n6327_));
  OAI21_X1   g06074(.A1(new_n6327_), .A2(new_n6325_), .B(new_n6298_), .ZN(new_n6328_));
  NAND2_X1   g06075(.A1(new_n6324_), .A2(new_n6328_), .ZN(new_n6329_));
  INV_X1     g06076(.I(new_n6329_), .ZN(new_n6330_));
  AOI21_X1   g06077(.A1(new_n6165_), .A2(new_n6210_), .B(new_n6208_), .ZN(new_n6331_));
  INV_X1     g06078(.I(new_n6188_), .ZN(new_n6332_));
  NAND2_X1   g06079(.A1(new_n6189_), .A2(new_n6190_), .ZN(new_n6333_));
  NAND2_X1   g06080(.A1(new_n6332_), .A2(new_n6333_), .ZN(new_n6334_));
  AOI21_X1   g06081(.A1(new_n2286_), .A2(new_n2690_), .B(new_n6196_), .ZN(new_n6335_));
  XOR2_X1    g06082(.A1(new_n6335_), .A2(new_n6334_), .Z(new_n6336_));
  INV_X1     g06083(.I(new_n6336_), .ZN(new_n6337_));
  INV_X1     g06084(.I(new_n6335_), .ZN(new_n6338_));
  NOR2_X1    g06085(.A1(new_n6338_), .A2(new_n6334_), .ZN(new_n6339_));
  INV_X1     g06086(.I(new_n6339_), .ZN(new_n6340_));
  NAND2_X1   g06087(.A1(new_n6338_), .A2(new_n6334_), .ZN(new_n6341_));
  AOI21_X1   g06088(.A1(new_n6340_), .A2(new_n6341_), .B(new_n6143_), .ZN(new_n6342_));
  AOI21_X1   g06089(.A1(new_n6337_), .A2(new_n6143_), .B(new_n6342_), .ZN(new_n6343_));
  NOR2_X1    g06090(.A1(new_n6186_), .A2(new_n6184_), .ZN(new_n6344_));
  NOR2_X1    g06091(.A1(new_n3981_), .A2(new_n1798_), .ZN(new_n6345_));
  NAND2_X1   g06092(.A1(new_n885_), .A2(new_n3371_), .ZN(new_n6346_));
  AOI21_X1   g06093(.A1(new_n1798_), .A2(new_n3981_), .B(new_n6346_), .ZN(new_n6347_));
  NOR2_X1    g06094(.A1(new_n6347_), .A2(new_n6345_), .ZN(new_n6348_));
  AOI21_X1   g06095(.A1(new_n267_), .A2(new_n6030_), .B(new_n6029_), .ZN(new_n6349_));
  XOR2_X1    g06096(.A1(new_n6349_), .A2(new_n6348_), .Z(new_n6350_));
  NAND2_X1   g06097(.A1(new_n6350_), .A2(new_n6344_), .ZN(new_n6351_));
  AND2_X2    g06098(.A1(new_n6349_), .A2(new_n6348_), .Z(new_n6352_));
  NOR2_X1    g06099(.A1(new_n6349_), .A2(new_n6348_), .ZN(new_n6353_));
  NOR2_X1    g06100(.A1(new_n6352_), .A2(new_n6353_), .ZN(new_n6354_));
  OAI21_X1   g06101(.A1(new_n6344_), .A2(new_n6354_), .B(new_n6351_), .ZN(new_n6355_));
  INV_X1     g06102(.I(new_n6201_), .ZN(new_n6356_));
  AOI21_X1   g06103(.A1(new_n6356_), .A2(new_n6187_), .B(new_n6199_), .ZN(new_n6357_));
  NOR2_X1    g06104(.A1(new_n6355_), .A2(new_n6357_), .ZN(new_n6358_));
  NAND2_X1   g06105(.A1(new_n6355_), .A2(new_n6357_), .ZN(new_n6359_));
  INV_X1     g06106(.I(new_n6359_), .ZN(new_n6360_));
  NOR2_X1    g06107(.A1(new_n6360_), .A2(new_n6358_), .ZN(new_n6361_));
  XNOR2_X1   g06108(.A1(new_n6355_), .A2(new_n6357_), .ZN(new_n6362_));
  INV_X1     g06109(.I(new_n6362_), .ZN(new_n6363_));
  NAND2_X1   g06110(.A1(new_n6363_), .A2(new_n6343_), .ZN(new_n6364_));
  OAI21_X1   g06111(.A1(new_n6343_), .A2(new_n6361_), .B(new_n6364_), .ZN(new_n6365_));
  XNOR2_X1   g06112(.A1(new_n6365_), .A2(new_n6331_), .ZN(new_n6366_));
  AND2_X2    g06113(.A1(new_n6365_), .A2(new_n6331_), .Z(new_n6367_));
  NOR2_X1    g06114(.A1(new_n6365_), .A2(new_n6331_), .ZN(new_n6368_));
  OAI21_X1   g06115(.A1(new_n6367_), .A2(new_n6368_), .B(new_n6330_), .ZN(new_n6369_));
  OAI21_X1   g06116(.A1(new_n6330_), .A2(new_n6366_), .B(new_n6369_), .ZN(new_n6370_));
  AND2_X2    g06117(.A1(new_n6370_), .A2(new_n6297_), .Z(new_n6371_));
  NOR2_X1    g06118(.A1(new_n6370_), .A2(new_n6297_), .ZN(new_n6372_));
  OAI21_X1   g06119(.A1(new_n6371_), .A2(new_n6372_), .B(new_n6251_), .ZN(new_n6373_));
  INV_X1     g06120(.I(new_n6251_), .ZN(new_n6374_));
  XOR2_X1    g06121(.A1(new_n6370_), .A2(new_n6297_), .Z(new_n6375_));
  NAND2_X1   g06122(.A1(new_n6375_), .A2(new_n6374_), .ZN(new_n6376_));
  NAND2_X1   g06123(.A1(new_n6376_), .A2(new_n6373_), .ZN(new_n6377_));
  NAND2_X1   g06124(.A1(new_n6087_), .A2(new_n6086_), .ZN(new_n6378_));
  NAND2_X1   g06125(.A1(new_n6378_), .A2(new_n6088_), .ZN(new_n6379_));
  OAI21_X1   g06126(.A1(new_n5923_), .A2(new_n6007_), .B(new_n6079_), .ZN(new_n6380_));
  OAI21_X1   g06127(.A1(new_n6045_), .A2(new_n6078_), .B(new_n6380_), .ZN(new_n6381_));
  NOR2_X1    g06128(.A1(new_n6003_), .A2(new_n5956_), .ZN(new_n6382_));
  NOR2_X1    g06129(.A1(new_n6382_), .A2(new_n6004_), .ZN(new_n6383_));
  NAND2_X1   g06130(.A1(new_n6047_), .A2(new_n6073_), .ZN(new_n6384_));
  NOR2_X1    g06131(.A1(new_n353_), .A2(new_n5511_), .ZN(new_n6385_));
  NOR3_X1    g06132(.A1(new_n798_), .A2(new_n3393_), .A3(new_n5175_), .ZN(new_n6386_));
  NAND4_X1   g06133(.A1(new_n6386_), .A2(\a[16] ), .A3(new_n6385_), .A4(\a[36] ), .ZN(new_n6387_));
  AOI21_X1   g06134(.A1(new_n6387_), .A2(new_n5793_), .B(new_n481_), .ZN(new_n6388_));
  NOR3_X1    g06135(.A1(new_n798_), .A2(new_n3393_), .A3(new_n5175_), .ZN(new_n6389_));
  NOR3_X1    g06136(.A1(new_n4240_), .A2(new_n4414_), .A3(new_n4769_), .ZN(new_n6390_));
  AOI21_X1   g06137(.A1(new_n1479_), .A2(new_n797_), .B(new_n6390_), .ZN(new_n6391_));
  INV_X1     g06138(.I(new_n6391_), .ZN(new_n6392_));
  NOR2_X1    g06139(.A1(new_n461_), .A2(new_n4769_), .ZN(new_n6393_));
  INV_X1     g06140(.I(new_n6393_), .ZN(new_n6394_));
  NOR4_X1    g06141(.A1(new_n6392_), .A2(new_n3061_), .A3(new_n5592_), .A4(new_n6394_), .ZN(new_n6395_));
  INV_X1     g06142(.I(new_n6395_), .ZN(new_n6396_));
  NAND2_X1   g06143(.A1(new_n5742_), .A2(new_n609_), .ZN(new_n6397_));
  NOR2_X1    g06144(.A1(new_n875_), .A2(new_n3837_), .ZN(new_n6398_));
  XOR2_X1    g06145(.A1(new_n6397_), .A2(new_n6398_), .Z(new_n6399_));
  NOR2_X1    g06146(.A1(new_n6396_), .A2(new_n6399_), .ZN(new_n6400_));
  INV_X1     g06147(.I(new_n6400_), .ZN(new_n6401_));
  NAND2_X1   g06148(.A1(new_n6396_), .A2(new_n6399_), .ZN(new_n6402_));
  NAND2_X1   g06149(.A1(new_n6401_), .A2(new_n6402_), .ZN(new_n6403_));
  XOR2_X1    g06150(.A1(new_n6395_), .A2(new_n6399_), .Z(new_n6404_));
  NOR2_X1    g06151(.A1(new_n6404_), .A2(new_n6389_), .ZN(new_n6405_));
  AOI21_X1   g06152(.A1(new_n6389_), .A2(new_n6403_), .B(new_n6405_), .ZN(new_n6406_));
  NOR2_X1    g06153(.A1(new_n4184_), .A2(new_n1711_), .ZN(new_n6407_));
  NOR2_X1    g06154(.A1(new_n4184_), .A2(new_n1711_), .ZN(new_n6411_));
  INV_X1     g06155(.I(new_n6411_), .ZN(new_n6412_));
  NOR2_X1    g06156(.A1(new_n5605_), .A2(new_n6137_), .ZN(new_n6413_));
  NOR4_X1    g06157(.A1(new_n364_), .A2(new_n599_), .A3(new_n3783_), .A4(new_n4501_), .ZN(new_n6419_));
  INV_X1     g06158(.I(new_n6419_), .ZN(new_n6420_));
  AOI22_X1   g06159(.A1(new_n2383_), .A2(new_n2898_), .B1(new_n3354_), .B2(new_n2286_), .ZN(new_n6421_));
  NOR4_X1    g06160(.A1(new_n2543_), .A2(new_n2690_), .A3(new_n1674_), .A4(new_n2461_), .ZN(new_n6422_));
  NAND2_X1   g06161(.A1(new_n6421_), .A2(new_n6422_), .ZN(new_n6423_));
  NOR2_X1    g06162(.A1(new_n6423_), .A2(new_n6420_), .ZN(new_n6424_));
  AOI21_X1   g06163(.A1(new_n6421_), .A2(new_n6422_), .B(new_n6419_), .ZN(new_n6425_));
  NOR2_X1    g06164(.A1(new_n6424_), .A2(new_n6425_), .ZN(new_n6426_));
  NOR2_X1    g06165(.A1(new_n6426_), .A2(new_n6412_), .ZN(new_n6427_));
  XOR2_X1    g06166(.A1(new_n6423_), .A2(new_n6419_), .Z(new_n6428_));
  NOR2_X1    g06167(.A1(new_n6428_), .A2(new_n6411_), .ZN(new_n6429_));
  NOR2_X1    g06168(.A1(new_n6429_), .A2(new_n6427_), .ZN(new_n6430_));
  XNOR2_X1   g06169(.A1(new_n6406_), .A2(new_n6430_), .ZN(new_n6431_));
  AOI21_X1   g06170(.A1(new_n6074_), .A2(new_n6384_), .B(new_n6431_), .ZN(new_n6432_));
  NAND2_X1   g06171(.A1(new_n6384_), .A2(new_n6074_), .ZN(new_n6433_));
  NOR2_X1    g06172(.A1(new_n6406_), .A2(new_n6430_), .ZN(new_n6434_));
  INV_X1     g06173(.I(new_n6434_), .ZN(new_n6435_));
  NAND2_X1   g06174(.A1(new_n6406_), .A2(new_n6430_), .ZN(new_n6436_));
  AOI21_X1   g06175(.A1(new_n6435_), .A2(new_n6436_), .B(new_n6433_), .ZN(new_n6437_));
  NOR2_X1    g06176(.A1(new_n6437_), .A2(new_n6432_), .ZN(new_n6438_));
  INV_X1     g06177(.I(new_n6438_), .ZN(new_n6439_));
  XOR2_X1    g06178(.A1(new_n6383_), .A2(new_n6439_), .Z(new_n6440_));
  NAND2_X1   g06179(.A1(new_n6381_), .A2(new_n6440_), .ZN(new_n6441_));
  INV_X1     g06180(.I(new_n6381_), .ZN(new_n6442_));
  NAND2_X1   g06181(.A1(new_n6383_), .A2(new_n6439_), .ZN(new_n6443_));
  INV_X1     g06182(.I(new_n6443_), .ZN(new_n6444_));
  NOR2_X1    g06183(.A1(new_n6383_), .A2(new_n6439_), .ZN(new_n6445_));
  OAI21_X1   g06184(.A1(new_n6444_), .A2(new_n6445_), .B(new_n6442_), .ZN(new_n6446_));
  NAND2_X1   g06185(.A1(new_n6446_), .A2(new_n6441_), .ZN(new_n6447_));
  XNOR2_X1   g06186(.A1(new_n6379_), .A2(new_n6447_), .ZN(new_n6448_));
  NAND3_X1   g06187(.A1(new_n6447_), .A2(new_n6088_), .A3(new_n6378_), .ZN(new_n6449_));
  NAND3_X1   g06188(.A1(new_n6379_), .A2(new_n6441_), .A3(new_n6446_), .ZN(new_n6450_));
  AOI21_X1   g06189(.A1(new_n6449_), .A2(new_n6450_), .B(new_n6377_), .ZN(new_n6451_));
  AOI21_X1   g06190(.A1(new_n6377_), .A2(new_n6448_), .B(new_n6451_), .ZN(new_n6452_));
  OAI21_X1   g06191(.A1(new_n6225_), .A2(new_n6221_), .B(new_n6223_), .ZN(new_n6453_));
  NAND2_X1   g06192(.A1(new_n6452_), .A2(new_n6453_), .ZN(new_n6454_));
  NOR2_X1    g06193(.A1(new_n6452_), .A2(new_n6453_), .ZN(new_n6455_));
  INV_X1     g06194(.I(new_n6455_), .ZN(new_n6456_));
  NAND2_X1   g06195(.A1(new_n6456_), .A2(new_n6454_), .ZN(new_n6457_));
  XNOR2_X1   g06196(.A1(new_n6250_), .A2(new_n6457_), .ZN(\asquared[53] ));
  NAND2_X1   g06197(.A1(new_n6454_), .A2(new_n6228_), .ZN(new_n6459_));
  OAI21_X1   g06198(.A1(new_n6454_), .A2(new_n6228_), .B(new_n6242_), .ZN(new_n6460_));
  AND2_X2    g06199(.A1(new_n6460_), .A2(new_n6459_), .Z(new_n6461_));
  NAND4_X1   g06200(.A1(new_n5835_), .A2(new_n5639_), .A3(new_n5833_), .A4(new_n6461_), .ZN(new_n6462_));
  INV_X1     g06201(.I(new_n6450_), .ZN(new_n6463_));
  AOI21_X1   g06202(.A1(new_n6377_), .A2(new_n6449_), .B(new_n6463_), .ZN(new_n6464_));
  INV_X1     g06203(.I(new_n6464_), .ZN(new_n6465_));
  NOR2_X1    g06204(.A1(new_n6374_), .A2(new_n6372_), .ZN(new_n6466_));
  NOR2_X1    g06205(.A1(new_n6466_), .A2(new_n6371_), .ZN(new_n6467_));
  INV_X1     g06206(.I(new_n6295_), .ZN(new_n6468_));
  AOI21_X1   g06207(.A1(new_n6253_), .A2(new_n6294_), .B(new_n6468_), .ZN(new_n6469_));
  INV_X1     g06208(.I(new_n6425_), .ZN(new_n6470_));
  AOI21_X1   g06209(.A1(new_n6470_), .A2(new_n6411_), .B(new_n6424_), .ZN(new_n6471_));
  INV_X1     g06210(.I(new_n6317_), .ZN(new_n6472_));
  AOI21_X1   g06211(.A1(new_n6300_), .A2(new_n6472_), .B(new_n6316_), .ZN(new_n6473_));
  NAND2_X1   g06212(.A1(new_n6280_), .A2(new_n232_), .ZN(new_n6474_));
  NOR2_X1    g06213(.A1(new_n6280_), .A2(new_n232_), .ZN(new_n6475_));
  NOR2_X1    g06214(.A1(\a[19] ), .A2(\a[33] ), .ZN(new_n6476_));
  AOI21_X1   g06215(.A1(new_n6474_), .A2(new_n6476_), .B(new_n6475_), .ZN(new_n6477_));
  AOI21_X1   g06216(.A1(new_n2543_), .A2(new_n2690_), .B(new_n6421_), .ZN(new_n6478_));
  XOR2_X1    g06217(.A1(new_n6308_), .A2(new_n6478_), .Z(new_n6479_));
  INV_X1     g06218(.I(new_n6479_), .ZN(new_n6480_));
  INV_X1     g06219(.I(new_n6478_), .ZN(new_n6481_));
  NOR2_X1    g06220(.A1(new_n6481_), .A2(new_n6308_), .ZN(new_n6482_));
  INV_X1     g06221(.I(new_n6482_), .ZN(new_n6483_));
  NAND2_X1   g06222(.A1(new_n6481_), .A2(new_n6308_), .ZN(new_n6484_));
  AOI21_X1   g06223(.A1(new_n6483_), .A2(new_n6484_), .B(new_n6477_), .ZN(new_n6485_));
  AOI21_X1   g06224(.A1(new_n6477_), .A2(new_n6480_), .B(new_n6485_), .ZN(new_n6486_));
  XOR2_X1    g06225(.A1(new_n6473_), .A2(new_n6486_), .Z(new_n6487_));
  NOR2_X1    g06226(.A1(new_n6487_), .A2(new_n6471_), .ZN(new_n6488_));
  INV_X1     g06227(.I(new_n6473_), .ZN(new_n6489_));
  NOR2_X1    g06228(.A1(new_n6489_), .A2(new_n6486_), .ZN(new_n6490_));
  INV_X1     g06229(.I(new_n6490_), .ZN(new_n6491_));
  NAND2_X1   g06230(.A1(new_n6489_), .A2(new_n6486_), .ZN(new_n6492_));
  NAND2_X1   g06231(.A1(new_n6491_), .A2(new_n6492_), .ZN(new_n6493_));
  AOI21_X1   g06232(.A1(new_n6471_), .A2(new_n6493_), .B(new_n6488_), .ZN(new_n6494_));
  AOI21_X1   g06233(.A1(new_n4985_), .A2(new_n4368_), .B(new_n6407_), .ZN(new_n6495_));
  NOR2_X1    g06234(.A1(new_n5742_), .A2(new_n609_), .ZN(new_n6496_));
  NAND2_X1   g06235(.A1(new_n875_), .A2(new_n3837_), .ZN(new_n6497_));
  AOI21_X1   g06236(.A1(new_n609_), .A2(new_n5742_), .B(new_n6497_), .ZN(new_n6498_));
  NOR2_X1    g06237(.A1(new_n6498_), .A2(new_n6496_), .ZN(new_n6499_));
  INV_X1     g06238(.I(new_n6499_), .ZN(new_n6500_));
  XOR2_X1    g06239(.A1(new_n6495_), .A2(new_n6500_), .Z(new_n6501_));
  NOR3_X1    g06240(.A1(new_n6501_), .A2(new_n6386_), .A3(new_n6388_), .ZN(new_n6502_));
  NOR2_X1    g06241(.A1(new_n6388_), .A2(new_n6386_), .ZN(new_n6503_));
  INV_X1     g06242(.I(new_n6495_), .ZN(new_n6504_));
  NOR2_X1    g06243(.A1(new_n6504_), .A2(new_n6500_), .ZN(new_n6505_));
  NOR2_X1    g06244(.A1(new_n6495_), .A2(new_n6499_), .ZN(new_n6506_));
  NOR2_X1    g06245(.A1(new_n6505_), .A2(new_n6506_), .ZN(new_n6507_));
  NOR2_X1    g06246(.A1(new_n6507_), .A2(new_n6503_), .ZN(new_n6508_));
  NOR2_X1    g06247(.A1(new_n6502_), .A2(new_n6508_), .ZN(new_n6509_));
  NAND2_X1   g06248(.A1(new_n6402_), .A2(new_n6389_), .ZN(new_n6510_));
  NAND2_X1   g06249(.A1(new_n6510_), .A2(new_n6401_), .ZN(new_n6511_));
  AOI21_X1   g06250(.A1(new_n787_), .A2(new_n5339_), .B(new_n6413_), .ZN(new_n6512_));
  AOI21_X1   g06251(.A1(new_n3061_), .A2(new_n5592_), .B(new_n6391_), .ZN(new_n6513_));
  NAND2_X1   g06252(.A1(\a[1] ), .A2(\a[52] ), .ZN(new_n6514_));
  XOR2_X1    g06253(.A1(new_n6514_), .A2(\a[27] ), .Z(new_n6515_));
  XOR2_X1    g06254(.A1(new_n6513_), .A2(new_n6515_), .Z(new_n6516_));
  NAND2_X1   g06255(.A1(new_n6516_), .A2(new_n6512_), .ZN(new_n6517_));
  INV_X1     g06256(.I(new_n6512_), .ZN(new_n6518_));
  NOR2_X1    g06257(.A1(new_n6513_), .A2(new_n6515_), .ZN(new_n6519_));
  AND2_X2    g06258(.A1(new_n6513_), .A2(new_n6515_), .Z(new_n6520_));
  OAI21_X1   g06259(.A1(new_n6520_), .A2(new_n6519_), .B(new_n6518_), .ZN(new_n6521_));
  NAND2_X1   g06260(.A1(new_n6517_), .A2(new_n6521_), .ZN(new_n6522_));
  XOR2_X1    g06261(.A1(new_n6511_), .A2(new_n6522_), .Z(new_n6523_));
  NOR2_X1    g06262(.A1(new_n6523_), .A2(new_n6509_), .ZN(new_n6524_));
  INV_X1     g06263(.I(new_n6509_), .ZN(new_n6525_));
  INV_X1     g06264(.I(new_n6522_), .ZN(new_n6526_));
  NOR2_X1    g06265(.A1(new_n6526_), .A2(new_n6511_), .ZN(new_n6527_));
  INV_X1     g06266(.I(new_n6527_), .ZN(new_n6528_));
  NAND2_X1   g06267(.A1(new_n6526_), .A2(new_n6511_), .ZN(new_n6529_));
  AOI21_X1   g06268(.A1(new_n6528_), .A2(new_n6529_), .B(new_n6525_), .ZN(new_n6530_));
  NOR2_X1    g06269(.A1(new_n6530_), .A2(new_n6524_), .ZN(new_n6531_));
  XOR2_X1    g06270(.A1(new_n6494_), .A2(new_n6531_), .Z(new_n6532_));
  INV_X1     g06271(.I(new_n6531_), .ZN(new_n6533_));
  NAND2_X1   g06272(.A1(new_n6494_), .A2(new_n6533_), .ZN(new_n6534_));
  NOR2_X1    g06273(.A1(new_n6494_), .A2(new_n6533_), .ZN(new_n6535_));
  INV_X1     g06274(.I(new_n6535_), .ZN(new_n6536_));
  NAND2_X1   g06275(.A1(new_n6536_), .A2(new_n6534_), .ZN(new_n6537_));
  NAND2_X1   g06276(.A1(new_n6469_), .A2(new_n6537_), .ZN(new_n6538_));
  OAI21_X1   g06277(.A1(new_n6469_), .A2(new_n6532_), .B(new_n6538_), .ZN(new_n6539_));
  AOI21_X1   g06278(.A1(new_n6433_), .A2(new_n6436_), .B(new_n6434_), .ZN(new_n6540_));
  AOI21_X1   g06279(.A1(new_n6299_), .A2(new_n6326_), .B(new_n6325_), .ZN(new_n6541_));
  AOI21_X1   g06280(.A1(new_n6143_), .A2(new_n6341_), .B(new_n6339_), .ZN(new_n6542_));
  INV_X1     g06281(.I(new_n6353_), .ZN(new_n6543_));
  AOI21_X1   g06282(.A1(new_n6344_), .A2(new_n6543_), .B(new_n6352_), .ZN(new_n6544_));
  OAI21_X1   g06283(.A1(new_n6265_), .A2(new_n6266_), .B(new_n6267_), .ZN(new_n6545_));
  XOR2_X1    g06284(.A1(new_n6544_), .A2(new_n6545_), .Z(new_n6546_));
  NOR2_X1    g06285(.A1(new_n6546_), .A2(new_n6542_), .ZN(new_n6547_));
  INV_X1     g06286(.I(new_n6542_), .ZN(new_n6548_));
  INV_X1     g06287(.I(new_n6545_), .ZN(new_n6549_));
  NOR2_X1    g06288(.A1(new_n6544_), .A2(new_n6549_), .ZN(new_n6550_));
  INV_X1     g06289(.I(new_n6550_), .ZN(new_n6551_));
  NAND2_X1   g06290(.A1(new_n6544_), .A2(new_n6549_), .ZN(new_n6552_));
  AOI21_X1   g06291(.A1(new_n6551_), .A2(new_n6552_), .B(new_n6548_), .ZN(new_n6553_));
  NOR2_X1    g06292(.A1(new_n6547_), .A2(new_n6553_), .ZN(new_n6554_));
  XOR2_X1    g06293(.A1(new_n6541_), .A2(new_n6554_), .Z(new_n6555_));
  NOR2_X1    g06294(.A1(new_n6555_), .A2(new_n6540_), .ZN(new_n6556_));
  INV_X1     g06295(.I(new_n6540_), .ZN(new_n6557_));
  INV_X1     g06296(.I(new_n6554_), .ZN(new_n6558_));
  NAND2_X1   g06297(.A1(new_n6541_), .A2(new_n6558_), .ZN(new_n6559_));
  NOR2_X1    g06298(.A1(new_n6541_), .A2(new_n6558_), .ZN(new_n6560_));
  INV_X1     g06299(.I(new_n6560_), .ZN(new_n6561_));
  AOI21_X1   g06300(.A1(new_n6561_), .A2(new_n6559_), .B(new_n6557_), .ZN(new_n6562_));
  OR2_X2     g06301(.A1(new_n6556_), .A2(new_n6562_), .Z(new_n6563_));
  INV_X1     g06302(.I(new_n6563_), .ZN(new_n6564_));
  INV_X1     g06303(.I(new_n6445_), .ZN(new_n6565_));
  OAI21_X1   g06304(.A1(new_n6442_), .A2(new_n6444_), .B(new_n6565_), .ZN(new_n6566_));
  NAND2_X1   g06305(.A1(new_n6566_), .A2(new_n6564_), .ZN(new_n6567_));
  INV_X1     g06306(.I(new_n6567_), .ZN(new_n6568_));
  NOR2_X1    g06307(.A1(new_n6566_), .A2(new_n6564_), .ZN(new_n6569_));
  OAI21_X1   g06308(.A1(new_n6568_), .A2(new_n6569_), .B(new_n6539_), .ZN(new_n6570_));
  XOR2_X1    g06309(.A1(new_n6566_), .A2(new_n6563_), .Z(new_n6571_));
  OAI21_X1   g06310(.A1(new_n6539_), .A2(new_n6571_), .B(new_n6570_), .ZN(new_n6572_));
  NOR2_X1    g06311(.A1(new_n6367_), .A2(new_n6329_), .ZN(new_n6573_));
  NOR2_X1    g06312(.A1(new_n6573_), .A2(new_n6368_), .ZN(new_n6574_));
  NOR2_X1    g06313(.A1(new_n6255_), .A2(new_n6272_), .ZN(new_n6575_));
  NOR2_X1    g06314(.A1(new_n6575_), .A2(new_n6273_), .ZN(new_n6576_));
  AOI21_X1   g06315(.A1(new_n6343_), .A2(new_n6359_), .B(new_n6358_), .ZN(new_n6577_));
  INV_X1     g06316(.I(new_n5003_), .ZN(new_n6578_));
  INV_X1     g06317(.I(new_n5592_), .ZN(new_n6579_));
  NOR2_X1    g06318(.A1(new_n6578_), .A2(new_n523_), .ZN(new_n6580_));
  NAND4_X1   g06319(.A1(new_n6580_), .A2(\a[10] ), .A3(new_n6136_), .A4(\a[40] ), .ZN(new_n6581_));
  AOI21_X1   g06320(.A1(new_n6581_), .A2(new_n6579_), .B(new_n1150_), .ZN(new_n6582_));
  NOR2_X1    g06321(.A1(new_n6578_), .A2(new_n523_), .ZN(new_n6583_));
  AOI22_X1   g06322(.A1(new_n2383_), .A2(new_n3126_), .B1(new_n3733_), .B2(new_n2286_), .ZN(new_n6584_));
  INV_X1     g06323(.I(new_n6584_), .ZN(new_n6585_));
  NOR4_X1    g06324(.A1(new_n6585_), .A2(new_n2543_), .A3(new_n2653_), .A4(new_n2898_), .ZN(new_n6586_));
  INV_X1     g06325(.I(new_n6586_), .ZN(new_n6587_));
  NOR2_X1    g06326(.A1(new_n2753_), .A2(new_n2692_), .ZN(new_n6588_));
  INV_X1     g06327(.I(new_n6588_), .ZN(new_n6589_));
  AOI21_X1   g06328(.A1(\a[25] ), .A2(\a[28] ), .B(new_n2533_), .ZN(new_n6590_));
  INV_X1     g06329(.I(new_n6590_), .ZN(new_n6591_));
  NOR2_X1    g06330(.A1(new_n6589_), .A2(new_n6591_), .ZN(new_n6592_));
  NAND2_X1   g06331(.A1(\a[11] ), .A2(\a[42] ), .ZN(new_n6593_));
  XOR2_X1    g06332(.A1(new_n6592_), .A2(new_n6593_), .Z(new_n6594_));
  NOR2_X1    g06333(.A1(new_n6594_), .A2(new_n6587_), .ZN(new_n6595_));
  INV_X1     g06334(.I(new_n6595_), .ZN(new_n6596_));
  NAND2_X1   g06335(.A1(new_n6594_), .A2(new_n6587_), .ZN(new_n6597_));
  NAND2_X1   g06336(.A1(new_n6596_), .A2(new_n6597_), .ZN(new_n6598_));
  XOR2_X1    g06337(.A1(new_n6594_), .A2(new_n6586_), .Z(new_n6599_));
  NOR2_X1    g06338(.A1(new_n6599_), .A2(new_n6583_), .ZN(new_n6600_));
  AOI21_X1   g06339(.A1(new_n6583_), .A2(new_n6598_), .B(new_n6600_), .ZN(new_n6601_));
  XNOR2_X1   g06340(.A1(new_n6601_), .A2(new_n6577_), .ZN(new_n6602_));
  NOR2_X1    g06341(.A1(new_n6602_), .A2(new_n6576_), .ZN(new_n6603_));
  INV_X1     g06342(.I(new_n6576_), .ZN(new_n6604_));
  NOR2_X1    g06343(.A1(new_n6601_), .A2(new_n6577_), .ZN(new_n6605_));
  INV_X1     g06344(.I(new_n6605_), .ZN(new_n6606_));
  NAND2_X1   g06345(.A1(new_n6601_), .A2(new_n6577_), .ZN(new_n6607_));
  AOI21_X1   g06346(.A1(new_n6606_), .A2(new_n6607_), .B(new_n6604_), .ZN(new_n6608_));
  NOR2_X1    g06347(.A1(new_n6603_), .A2(new_n6608_), .ZN(new_n6609_));
  AOI21_X1   g06348(.A1(new_n6277_), .A2(new_n6287_), .B(new_n6285_), .ZN(new_n6610_));
  NOR2_X1    g06349(.A1(new_n359_), .A2(new_n5004_), .ZN(new_n6611_));
  NAND3_X1   g06350(.A1(new_n6611_), .A2(\a[14] ), .A3(\a[39] ), .ZN(new_n6612_));
  OAI21_X1   g06351(.A1(new_n453_), .A2(new_n5743_), .B(new_n6612_), .ZN(new_n6613_));
  NOR2_X1    g06352(.A1(new_n650_), .A2(new_n4770_), .ZN(new_n6614_));
  INV_X1     g06353(.I(new_n6614_), .ZN(new_n6615_));
  NOR2_X1    g06354(.A1(new_n5605_), .A2(new_n6615_), .ZN(new_n6616_));
  INV_X1     g06355(.I(new_n6616_), .ZN(new_n6617_));
  AOI22_X1   g06356(.A1(\a[9] ), .A2(\a[14] ), .B1(\a[39] ), .B2(\a[44] ), .ZN(new_n6618_));
  NAND4_X1   g06357(.A1(new_n6617_), .A2(new_n6613_), .A3(new_n6611_), .A4(new_n6618_), .ZN(new_n6619_));
  NAND4_X1   g06358(.A1(\a[6] ), .A2(\a[7] ), .A3(\a[46] ), .A4(\a[47] ), .ZN(new_n6621_));
  NAND4_X1   g06359(.A1(\a[5] ), .A2(\a[16] ), .A3(\a[37] ), .A4(\a[48] ), .ZN(new_n6622_));
  NAND2_X1   g06360(.A1(\a[0] ), .A2(\a[53] ), .ZN(new_n6623_));
  XNOR2_X1   g06361(.A1(new_n6622_), .A2(new_n6623_), .ZN(new_n6624_));
  NOR2_X1    g06362(.A1(new_n6624_), .A2(new_n6621_), .ZN(new_n6625_));
  AND2_X2    g06363(.A1(new_n6624_), .A2(new_n6621_), .Z(new_n6626_));
  NOR2_X1    g06364(.A1(new_n6626_), .A2(new_n6625_), .ZN(new_n6627_));
  NOR2_X1    g06365(.A1(new_n6627_), .A2(new_n6619_), .ZN(new_n6628_));
  INV_X1     g06366(.I(new_n6619_), .ZN(new_n6629_));
  XNOR2_X1   g06367(.A1(new_n6624_), .A2(new_n6621_), .ZN(new_n6630_));
  NOR2_X1    g06368(.A1(new_n6630_), .A2(new_n6629_), .ZN(new_n6631_));
  NOR2_X1    g06369(.A1(new_n6628_), .A2(new_n6631_), .ZN(new_n6632_));
  NAND2_X1   g06370(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n6633_));
  XNOR2_X1   g06371(.A1(new_n225_), .A2(new_n6633_), .ZN(new_n6634_));
  NAND2_X1   g06372(.A1(new_n3966_), .A2(new_n1441_), .ZN(new_n6635_));
  NOR2_X1    g06373(.A1(new_n282_), .A2(new_n5745_), .ZN(new_n6636_));
  XOR2_X1    g06374(.A1(new_n6635_), .A2(new_n6636_), .Z(new_n6637_));
  NOR2_X1    g06375(.A1(new_n1710_), .A2(new_n1715_), .ZN(new_n6638_));
  AOI21_X1   g06376(.A1(new_n4368_), .A2(new_n4372_), .B(new_n6638_), .ZN(new_n6639_));
  NOR4_X1    g06377(.A1(new_n3851_), .A2(new_n2978_), .A3(new_n1339_), .A4(new_n3371_), .ZN(new_n6640_));
  NAND2_X1   g06378(.A1(new_n6639_), .A2(new_n6640_), .ZN(new_n6641_));
  NOR2_X1    g06379(.A1(new_n6637_), .A2(new_n6641_), .ZN(new_n6642_));
  INV_X1     g06380(.I(new_n6642_), .ZN(new_n6643_));
  NAND2_X1   g06381(.A1(new_n6637_), .A2(new_n6641_), .ZN(new_n6644_));
  AOI21_X1   g06382(.A1(new_n6643_), .A2(new_n6644_), .B(new_n6634_), .ZN(new_n6645_));
  INV_X1     g06383(.I(new_n6634_), .ZN(new_n6646_));
  XNOR2_X1   g06384(.A1(new_n6637_), .A2(new_n6641_), .ZN(new_n6647_));
  NOR2_X1    g06385(.A1(new_n6647_), .A2(new_n6646_), .ZN(new_n6648_));
  NOR2_X1    g06386(.A1(new_n6648_), .A2(new_n6645_), .ZN(new_n6649_));
  XNOR2_X1   g06387(.A1(new_n6649_), .A2(new_n6632_), .ZN(new_n6650_));
  NOR2_X1    g06388(.A1(new_n6650_), .A2(new_n6610_), .ZN(new_n6651_));
  INV_X1     g06389(.I(new_n6610_), .ZN(new_n6652_));
  NOR2_X1    g06390(.A1(new_n6649_), .A2(new_n6632_), .ZN(new_n6653_));
  INV_X1     g06391(.I(new_n6653_), .ZN(new_n6654_));
  NAND2_X1   g06392(.A1(new_n6649_), .A2(new_n6632_), .ZN(new_n6655_));
  AOI21_X1   g06393(.A1(new_n6654_), .A2(new_n6655_), .B(new_n6652_), .ZN(new_n6656_));
  NOR2_X1    g06394(.A1(new_n6651_), .A2(new_n6656_), .ZN(new_n6657_));
  XNOR2_X1   g06395(.A1(new_n6609_), .A2(new_n6657_), .ZN(new_n6658_));
  NOR2_X1    g06396(.A1(new_n6609_), .A2(new_n6657_), .ZN(new_n6659_));
  NAND2_X1   g06397(.A1(new_n6609_), .A2(new_n6657_), .ZN(new_n6660_));
  INV_X1     g06398(.I(new_n6660_), .ZN(new_n6661_));
  OAI21_X1   g06399(.A1(new_n6659_), .A2(new_n6661_), .B(new_n6574_), .ZN(new_n6662_));
  OAI21_X1   g06400(.A1(new_n6574_), .A2(new_n6658_), .B(new_n6662_), .ZN(new_n6663_));
  XNOR2_X1   g06401(.A1(new_n6572_), .A2(new_n6663_), .ZN(new_n6664_));
  NAND2_X1   g06402(.A1(new_n6572_), .A2(new_n6663_), .ZN(new_n6665_));
  NOR2_X1    g06403(.A1(new_n6572_), .A2(new_n6663_), .ZN(new_n6666_));
  INV_X1     g06404(.I(new_n6666_), .ZN(new_n6667_));
  NAND2_X1   g06405(.A1(new_n6667_), .A2(new_n6665_), .ZN(new_n6668_));
  NAND2_X1   g06406(.A1(new_n6668_), .A2(new_n6467_), .ZN(new_n6669_));
  OAI21_X1   g06407(.A1(new_n6467_), .A2(new_n6664_), .B(new_n6669_), .ZN(new_n6670_));
  NAND2_X1   g06408(.A1(new_n6670_), .A2(new_n6465_), .ZN(new_n6671_));
  XOR2_X1    g06409(.A1(new_n6462_), .A2(new_n6671_), .Z(new_n6672_));
  XOR2_X1    g06410(.A1(new_n6672_), .A2(new_n6455_), .Z(\asquared[54] ));
  OAI21_X1   g06411(.A1(new_n6670_), .A2(new_n6465_), .B(new_n6455_), .ZN(new_n6674_));
  OAI21_X1   g06412(.A1(new_n6462_), .A2(new_n6674_), .B(new_n6671_), .ZN(new_n6675_));
  INV_X1     g06413(.I(new_n6675_), .ZN(new_n6676_));
  INV_X1     g06414(.I(new_n6467_), .ZN(new_n6677_));
  AOI21_X1   g06415(.A1(new_n6677_), .A2(new_n6665_), .B(new_n6666_), .ZN(new_n6678_));
  OAI21_X1   g06416(.A1(new_n6469_), .A2(new_n6535_), .B(new_n6534_), .ZN(new_n6679_));
  NAND2_X1   g06417(.A1(new_n6559_), .A2(new_n6557_), .ZN(new_n6680_));
  NAND2_X1   g06418(.A1(new_n6680_), .A2(new_n6561_), .ZN(new_n6681_));
  INV_X1     g06419(.I(new_n6681_), .ZN(new_n6682_));
  OAI21_X1   g06420(.A1(new_n6525_), .A2(new_n6527_), .B(new_n6529_), .ZN(new_n6683_));
  OAI21_X1   g06421(.A1(new_n6471_), .A2(new_n6490_), .B(new_n6492_), .ZN(new_n6684_));
  INV_X1     g06422(.I(new_n6684_), .ZN(new_n6685_));
  NOR2_X1    g06423(.A1(new_n3852_), .A2(new_n1773_), .ZN(new_n6686_));
  NOR2_X1    g06424(.A1(new_n3852_), .A2(new_n1773_), .ZN(new_n6690_));
  INV_X1     g06425(.I(new_n6690_), .ZN(new_n6691_));
  INV_X1     g06426(.I(\a[52] ), .ZN(new_n6692_));
  NOR2_X1    g06427(.A1(new_n2256_), .A2(new_n6692_), .ZN(new_n6693_));
  INV_X1     g06428(.I(\a[53] ), .ZN(new_n6694_));
  NOR2_X1    g06429(.A1(new_n194_), .A2(new_n6694_), .ZN(new_n6695_));
  XOR2_X1    g06430(.A1(new_n6695_), .A2(new_n3036_), .Z(new_n6696_));
  NAND2_X1   g06431(.A1(new_n6696_), .A2(new_n6693_), .ZN(new_n6697_));
  XOR2_X1    g06432(.A1(new_n6697_), .A2(\a[0] ), .Z(new_n6698_));
  XOR2_X1    g06433(.A1(new_n6698_), .A2(\a[54] ), .Z(new_n6699_));
  NOR2_X1    g06434(.A1(new_n1912_), .A2(new_n1956_), .ZN(new_n6700_));
  AOI21_X1   g06435(.A1(new_n3126_), .A2(new_n3733_), .B(new_n6700_), .ZN(new_n6701_));
  INV_X1     g06436(.I(new_n6701_), .ZN(new_n6702_));
  NOR2_X1    g06437(.A1(new_n3175_), .A2(new_n2276_), .ZN(new_n6703_));
  NAND2_X1   g06438(.A1(\a[23] ), .A2(\a[31] ), .ZN(new_n6704_));
  AOI21_X1   g06439(.A1(\a[25] ), .A2(\a[29] ), .B(new_n2899_), .ZN(new_n6705_));
  NOR4_X1    g06440(.A1(new_n6702_), .A2(new_n6703_), .A3(new_n6704_), .A4(new_n6705_), .ZN(new_n6706_));
  INV_X1     g06441(.I(new_n6706_), .ZN(new_n6707_));
  NOR2_X1    g06442(.A1(new_n6699_), .A2(new_n6707_), .ZN(new_n6708_));
  INV_X1     g06443(.I(new_n6708_), .ZN(new_n6709_));
  NAND2_X1   g06444(.A1(new_n6699_), .A2(new_n6707_), .ZN(new_n6710_));
  AOI21_X1   g06445(.A1(new_n6709_), .A2(new_n6710_), .B(new_n6691_), .ZN(new_n6711_));
  XOR2_X1    g06446(.A1(new_n6699_), .A2(new_n6706_), .Z(new_n6712_));
  NOR2_X1    g06447(.A1(new_n6712_), .A2(new_n6690_), .ZN(new_n6713_));
  NOR2_X1    g06448(.A1(new_n6713_), .A2(new_n6711_), .ZN(new_n6714_));
  NOR2_X1    g06449(.A1(new_n6714_), .A2(new_n6685_), .ZN(new_n6715_));
  NOR3_X1    g06450(.A1(new_n6684_), .A2(new_n6713_), .A3(new_n6711_), .ZN(new_n6716_));
  NOR2_X1    g06451(.A1(new_n6715_), .A2(new_n6716_), .ZN(new_n6717_));
  XOR2_X1    g06452(.A1(new_n6714_), .A2(new_n6684_), .Z(new_n6718_));
  MUX2_X1    g06453(.I0(new_n6718_), .I1(new_n6717_), .S(new_n6683_), .Z(new_n6719_));
  NOR2_X1    g06454(.A1(new_n6719_), .A2(new_n6682_), .ZN(new_n6720_));
  INV_X1     g06455(.I(new_n6720_), .ZN(new_n6721_));
  NAND2_X1   g06456(.A1(new_n6719_), .A2(new_n6682_), .ZN(new_n6722_));
  NAND2_X1   g06457(.A1(new_n6721_), .A2(new_n6722_), .ZN(new_n6723_));
  XOR2_X1    g06458(.A1(new_n6719_), .A2(new_n6681_), .Z(new_n6724_));
  NOR2_X1    g06459(.A1(new_n6724_), .A2(new_n6679_), .ZN(new_n6725_));
  AOI21_X1   g06460(.A1(new_n6679_), .A2(new_n6723_), .B(new_n6725_), .ZN(new_n6726_));
  OAI21_X1   g06461(.A1(new_n6539_), .A2(new_n6569_), .B(new_n6567_), .ZN(new_n6727_));
  INV_X1     g06462(.I(new_n6727_), .ZN(new_n6728_));
  OAI21_X1   g06463(.A1(new_n6574_), .A2(new_n6659_), .B(new_n6660_), .ZN(new_n6729_));
  INV_X1     g06464(.I(new_n6729_), .ZN(new_n6730_));
  AOI21_X1   g06465(.A1(new_n6604_), .A2(new_n6607_), .B(new_n6605_), .ZN(new_n6731_));
  NOR2_X1    g06466(.A1(new_n1276_), .A2(new_n5745_), .ZN(new_n6732_));
  INV_X1     g06467(.I(new_n6732_), .ZN(new_n6733_));
  NOR3_X1    g06468(.A1(new_n6733_), .A2(new_n353_), .A3(new_n3393_), .ZN(new_n6734_));
  NOR2_X1    g06469(.A1(new_n1215_), .A2(new_n5745_), .ZN(new_n6735_));
  NAND4_X1   g06470(.A1(new_n6734_), .A2(\a[5] ), .A3(new_n6735_), .A4(\a[34] ), .ZN(new_n6736_));
  AOI21_X1   g06471(.A1(new_n6736_), .A2(new_n4728_), .B(new_n1536_), .ZN(new_n6737_));
  NOR3_X1    g06472(.A1(new_n6737_), .A2(new_n1215_), .A3(new_n3371_), .ZN(new_n6738_));
  NOR2_X1    g06473(.A1(new_n6737_), .A2(new_n6734_), .ZN(new_n6739_));
  NOR2_X1    g06474(.A1(new_n3393_), .A2(new_n5745_), .ZN(new_n6740_));
  NOR2_X1    g06475(.A1(new_n1531_), .A2(new_n6740_), .ZN(new_n6741_));
  AOI21_X1   g06476(.A1(new_n6739_), .A2(new_n6741_), .B(new_n6738_), .ZN(new_n6742_));
  NOR2_X1    g06477(.A1(new_n3804_), .A2(new_n5750_), .ZN(new_n6743_));
  INV_X1     g06478(.I(new_n6743_), .ZN(new_n6744_));
  NOR2_X1    g06479(.A1(new_n6744_), .A2(new_n798_), .ZN(new_n6745_));
  NOR2_X1    g06480(.A1(new_n6744_), .A2(new_n798_), .ZN(new_n6749_));
  INV_X1     g06481(.I(new_n6749_), .ZN(new_n6750_));
  AOI22_X1   g06482(.A1(new_n5003_), .A2(new_n5350_), .B1(new_n1220_), .B2(new_n1001_), .ZN(new_n6751_));
  NOR4_X1    g06483(.A1(new_n5173_), .A2(new_n3061_), .A3(new_n599_), .A4(new_n4414_), .ZN(new_n6752_));
  NAND2_X1   g06484(.A1(new_n6751_), .A2(new_n6752_), .ZN(new_n6753_));
  NOR2_X1    g06485(.A1(new_n6753_), .A2(new_n6750_), .ZN(new_n6754_));
  INV_X1     g06486(.I(new_n6754_), .ZN(new_n6755_));
  NAND2_X1   g06487(.A1(new_n6753_), .A2(new_n6750_), .ZN(new_n6756_));
  NAND2_X1   g06488(.A1(new_n6755_), .A2(new_n6756_), .ZN(new_n6757_));
  XOR2_X1    g06489(.A1(new_n6753_), .A2(new_n6749_), .Z(new_n6758_));
  NOR2_X1    g06490(.A1(new_n6742_), .A2(new_n6758_), .ZN(new_n6759_));
  AOI21_X1   g06491(.A1(new_n6742_), .A2(new_n6757_), .B(new_n6759_), .ZN(new_n6760_));
  INV_X1     g06492(.I(new_n6760_), .ZN(new_n6761_));
  NAND2_X1   g06493(.A1(new_n6548_), .A2(new_n6552_), .ZN(new_n6762_));
  NAND2_X1   g06494(.A1(new_n6762_), .A2(new_n6551_), .ZN(new_n6763_));
  NOR3_X1    g06495(.A1(new_n6615_), .A2(new_n461_), .A3(new_n4240_), .ZN(new_n6764_));
  NOR4_X1    g06496(.A1(new_n364_), .A2(new_n650_), .A3(new_n4240_), .A4(new_n5004_), .ZN(new_n6765_));
  NAND2_X1   g06497(.A1(new_n6764_), .A2(new_n6765_), .ZN(new_n6766_));
  NAND2_X1   g06498(.A1(new_n6766_), .A2(new_n5743_), .ZN(new_n6767_));
  NAND2_X1   g06499(.A1(\a[9] ), .A2(\a[45] ), .ZN(new_n6768_));
  AOI21_X1   g06500(.A1(new_n6767_), .A2(new_n597_), .B(new_n6768_), .ZN(new_n6769_));
  AOI21_X1   g06501(.A1(new_n597_), .A2(new_n5742_), .B(new_n6764_), .ZN(new_n6770_));
  INV_X1     g06502(.I(new_n6770_), .ZN(new_n6771_));
  NOR2_X1    g06503(.A1(new_n4240_), .A2(new_n4770_), .ZN(new_n6772_));
  NOR2_X1    g06504(.A1(new_n461_), .A2(new_n650_), .ZN(new_n6773_));
  NOR3_X1    g06505(.A1(new_n6771_), .A2(new_n6772_), .A3(new_n6773_), .ZN(new_n6774_));
  NOR2_X1    g06506(.A1(new_n6774_), .A2(new_n6769_), .ZN(new_n6775_));
  NOR2_X1    g06507(.A1(new_n6055_), .A2(new_n6692_), .ZN(new_n6776_));
  NOR2_X1    g06508(.A1(new_n6260_), .A2(new_n6692_), .ZN(new_n6777_));
  AOI21_X1   g06509(.A1(new_n6776_), .A2(new_n6777_), .B(new_n1271_), .ZN(new_n6778_));
  NOR2_X1    g06510(.A1(new_n6055_), .A2(new_n6260_), .ZN(new_n6779_));
  NOR4_X1    g06511(.A1(new_n6779_), .A2(new_n267_), .A3(new_n201_), .A4(new_n6692_), .ZN(new_n6780_));
  NAND2_X1   g06512(.A1(new_n6778_), .A2(new_n6780_), .ZN(new_n6781_));
  NOR2_X1    g06513(.A1(new_n875_), .A2(new_n3783_), .ZN(new_n6782_));
  NAND4_X1   g06514(.A1(\a[7] ), .A2(\a[8] ), .A3(\a[46] ), .A4(\a[47] ), .ZN(new_n6783_));
  OR2_X2     g06515(.A1(new_n6781_), .A2(new_n6783_), .Z(new_n6784_));
  NAND2_X1   g06516(.A1(new_n6781_), .A2(new_n6783_), .ZN(new_n6785_));
  NAND2_X1   g06517(.A1(new_n6784_), .A2(new_n6785_), .ZN(new_n6786_));
  NAND2_X1   g06518(.A1(new_n6775_), .A2(new_n6786_), .ZN(new_n6787_));
  XNOR2_X1   g06519(.A1(new_n6781_), .A2(new_n6783_), .ZN(new_n6788_));
  OAI21_X1   g06520(.A1(new_n6775_), .A2(new_n6788_), .B(new_n6787_), .ZN(new_n6789_));
  XOR2_X1    g06521(.A1(new_n6763_), .A2(new_n6789_), .Z(new_n6790_));
  NAND2_X1   g06522(.A1(new_n6763_), .A2(new_n6789_), .ZN(new_n6791_));
  NOR2_X1    g06523(.A1(new_n6763_), .A2(new_n6789_), .ZN(new_n6792_));
  INV_X1     g06524(.I(new_n6792_), .ZN(new_n6793_));
  AOI21_X1   g06525(.A1(new_n6793_), .A2(new_n6791_), .B(new_n6761_), .ZN(new_n6794_));
  AOI21_X1   g06526(.A1(new_n6761_), .A2(new_n6790_), .B(new_n6794_), .ZN(new_n6795_));
  NOR2_X1    g06527(.A1(new_n6582_), .A2(new_n6580_), .ZN(new_n6796_));
  NOR3_X1    g06528(.A1(new_n2891_), .A2(new_n194_), .A3(new_n6260_), .ZN(new_n6797_));
  AOI21_X1   g06529(.A1(new_n6797_), .A2(new_n232_), .B(new_n6779_), .ZN(new_n6798_));
  XOR2_X1    g06530(.A1(new_n6796_), .A2(new_n6798_), .Z(new_n6799_));
  NOR3_X1    g06531(.A1(new_n6799_), .A2(new_n6613_), .A3(new_n6616_), .ZN(new_n6800_));
  NOR2_X1    g06532(.A1(new_n6613_), .A2(new_n6616_), .ZN(new_n6801_));
  INV_X1     g06533(.I(new_n6796_), .ZN(new_n6802_));
  NOR2_X1    g06534(.A1(new_n6802_), .A2(new_n6798_), .ZN(new_n6803_));
  INV_X1     g06535(.I(new_n6803_), .ZN(new_n6804_));
  NAND2_X1   g06536(.A1(new_n6802_), .A2(new_n6798_), .ZN(new_n6805_));
  AOI21_X1   g06537(.A1(new_n6804_), .A2(new_n6805_), .B(new_n6801_), .ZN(new_n6806_));
  NOR2_X1    g06538(.A1(new_n6806_), .A2(new_n6800_), .ZN(new_n6807_));
  NAND2_X1   g06539(.A1(new_n6597_), .A2(new_n6583_), .ZN(new_n6808_));
  NAND2_X1   g06540(.A1(new_n6808_), .A2(new_n6596_), .ZN(new_n6809_));
  NAND2_X1   g06541(.A1(new_n6644_), .A2(new_n6646_), .ZN(new_n6810_));
  NAND2_X1   g06542(.A1(new_n6810_), .A2(new_n6643_), .ZN(new_n6811_));
  NAND2_X1   g06543(.A1(new_n6809_), .A2(new_n6811_), .ZN(new_n6812_));
  INV_X1     g06544(.I(new_n6811_), .ZN(new_n6813_));
  NAND3_X1   g06545(.A1(new_n6808_), .A2(new_n6596_), .A3(new_n6813_), .ZN(new_n6814_));
  AOI21_X1   g06546(.A1(new_n6812_), .A2(new_n6814_), .B(new_n6807_), .ZN(new_n6815_));
  XOR2_X1    g06547(.A1(new_n6809_), .A2(new_n6811_), .Z(new_n6816_));
  AOI21_X1   g06548(.A1(new_n6816_), .A2(new_n6807_), .B(new_n6815_), .ZN(new_n6817_));
  NOR2_X1    g06549(.A1(new_n6795_), .A2(new_n6817_), .ZN(new_n6818_));
  INV_X1     g06550(.I(new_n6818_), .ZN(new_n6819_));
  NAND2_X1   g06551(.A1(new_n6795_), .A2(new_n6817_), .ZN(new_n6820_));
  AOI21_X1   g06552(.A1(new_n6819_), .A2(new_n6820_), .B(new_n6731_), .ZN(new_n6821_));
  INV_X1     g06553(.I(new_n6731_), .ZN(new_n6822_));
  XNOR2_X1   g06554(.A1(new_n6795_), .A2(new_n6817_), .ZN(new_n6823_));
  NOR2_X1    g06555(.A1(new_n6823_), .A2(new_n6822_), .ZN(new_n6824_));
  NOR2_X1    g06556(.A1(new_n6824_), .A2(new_n6821_), .ZN(new_n6825_));
  INV_X1     g06557(.I(new_n6825_), .ZN(new_n6826_));
  AOI21_X1   g06558(.A1(new_n6652_), .A2(new_n6655_), .B(new_n6653_), .ZN(new_n6827_));
  INV_X1     g06559(.I(new_n6506_), .ZN(new_n6828_));
  AOI21_X1   g06560(.A1(new_n6503_), .A2(new_n6828_), .B(new_n6505_), .ZN(new_n6829_));
  NOR2_X1    g06561(.A1(new_n6519_), .A2(new_n6518_), .ZN(new_n6830_));
  NOR2_X1    g06562(.A1(new_n6830_), .A2(new_n6520_), .ZN(new_n6831_));
  NAND2_X1   g06563(.A1(new_n6484_), .A2(new_n6477_), .ZN(new_n6832_));
  NAND2_X1   g06564(.A1(new_n6832_), .A2(new_n6483_), .ZN(new_n6833_));
  XOR2_X1    g06565(.A1(new_n6833_), .A2(new_n6831_), .Z(new_n6834_));
  INV_X1     g06566(.I(new_n6833_), .ZN(new_n6835_));
  NOR2_X1    g06567(.A1(new_n6835_), .A2(new_n6831_), .ZN(new_n6836_));
  NAND2_X1   g06568(.A1(new_n6835_), .A2(new_n6831_), .ZN(new_n6837_));
  INV_X1     g06569(.I(new_n6837_), .ZN(new_n6838_));
  OAI21_X1   g06570(.A1(new_n6838_), .A2(new_n6836_), .B(new_n6829_), .ZN(new_n6839_));
  OAI21_X1   g06571(.A1(new_n6829_), .A2(new_n6834_), .B(new_n6839_), .ZN(new_n6840_));
  NOR2_X1    g06572(.A1(new_n6626_), .A2(new_n6619_), .ZN(new_n6841_));
  NOR2_X1    g06573(.A1(new_n6841_), .A2(new_n6625_), .ZN(new_n6842_));
  NOR4_X1    g06574(.A1(new_n242_), .A2(new_n268_), .A3(new_n5175_), .A4(new_n5511_), .ZN(new_n6843_));
  NOR4_X1    g06575(.A1(new_n353_), .A2(new_n800_), .A3(new_n3837_), .A4(new_n5750_), .ZN(new_n6844_));
  NOR2_X1    g06576(.A1(new_n3837_), .A2(new_n5750_), .ZN(new_n6845_));
  NAND2_X1   g06577(.A1(new_n199_), .A2(new_n6694_), .ZN(new_n6846_));
  OAI22_X1   g06578(.A1(new_n6844_), .A2(new_n6846_), .B1(new_n1344_), .B2(new_n6845_), .ZN(new_n6847_));
  NOR2_X1    g06579(.A1(\a[11] ), .A2(\a[42] ), .ZN(new_n6848_));
  AOI21_X1   g06580(.A1(new_n6589_), .A2(new_n6848_), .B(new_n6591_), .ZN(new_n6849_));
  XNOR2_X1   g06581(.A1(new_n6849_), .A2(new_n6847_), .ZN(new_n6850_));
  NAND2_X1   g06582(.A1(new_n6850_), .A2(new_n6843_), .ZN(new_n6851_));
  INV_X1     g06583(.I(new_n6843_), .ZN(new_n6852_));
  INV_X1     g06584(.I(new_n6849_), .ZN(new_n6853_));
  NOR2_X1    g06585(.A1(new_n6853_), .A2(new_n6847_), .ZN(new_n6854_));
  NAND2_X1   g06586(.A1(new_n6853_), .A2(new_n6847_), .ZN(new_n6855_));
  INV_X1     g06587(.I(new_n6855_), .ZN(new_n6856_));
  OAI21_X1   g06588(.A1(new_n6856_), .A2(new_n6854_), .B(new_n6852_), .ZN(new_n6857_));
  NAND2_X1   g06589(.A1(new_n6857_), .A2(new_n6851_), .ZN(new_n6858_));
  NAND2_X1   g06590(.A1(new_n3966_), .A2(new_n1441_), .ZN(new_n6859_));
  NOR2_X1    g06591(.A1(new_n3966_), .A2(new_n1441_), .ZN(new_n6860_));
  NOR2_X1    g06592(.A1(\a[4] ), .A2(\a[49] ), .ZN(new_n6861_));
  AOI21_X1   g06593(.A1(new_n6859_), .A2(new_n6861_), .B(new_n6860_), .ZN(new_n6862_));
  AOI21_X1   g06594(.A1(new_n2978_), .A2(new_n3851_), .B(new_n6639_), .ZN(new_n6863_));
  AOI21_X1   g06595(.A1(new_n2543_), .A2(new_n2898_), .B(new_n6584_), .ZN(new_n6864_));
  XOR2_X1    g06596(.A1(new_n6863_), .A2(new_n6864_), .Z(new_n6865_));
  NAND2_X1   g06597(.A1(new_n6865_), .A2(new_n6862_), .ZN(new_n6866_));
  INV_X1     g06598(.I(new_n6862_), .ZN(new_n6867_));
  AND2_X2    g06599(.A1(new_n6863_), .A2(new_n6864_), .Z(new_n6868_));
  NOR2_X1    g06600(.A1(new_n6863_), .A2(new_n6864_), .ZN(new_n6869_));
  OAI21_X1   g06601(.A1(new_n6868_), .A2(new_n6869_), .B(new_n6867_), .ZN(new_n6870_));
  NAND2_X1   g06602(.A1(new_n6866_), .A2(new_n6870_), .ZN(new_n6871_));
  XNOR2_X1   g06603(.A1(new_n6858_), .A2(new_n6871_), .ZN(new_n6872_));
  AOI22_X1   g06604(.A1(new_n6857_), .A2(new_n6851_), .B1(new_n6866_), .B2(new_n6870_), .ZN(new_n6873_));
  NOR2_X1    g06605(.A1(new_n6858_), .A2(new_n6871_), .ZN(new_n6874_));
  OAI21_X1   g06606(.A1(new_n6874_), .A2(new_n6873_), .B(new_n6842_), .ZN(new_n6875_));
  OAI21_X1   g06607(.A1(new_n6872_), .A2(new_n6842_), .B(new_n6875_), .ZN(new_n6876_));
  XNOR2_X1   g06608(.A1(new_n6876_), .A2(new_n6840_), .ZN(new_n6877_));
  NOR2_X1    g06609(.A1(new_n6877_), .A2(new_n6827_), .ZN(new_n6878_));
  INV_X1     g06610(.I(new_n6827_), .ZN(new_n6879_));
  NAND2_X1   g06611(.A1(new_n6876_), .A2(new_n6840_), .ZN(new_n6880_));
  NOR2_X1    g06612(.A1(new_n6876_), .A2(new_n6840_), .ZN(new_n6881_));
  INV_X1     g06613(.I(new_n6881_), .ZN(new_n6882_));
  AOI21_X1   g06614(.A1(new_n6882_), .A2(new_n6880_), .B(new_n6879_), .ZN(new_n6883_));
  NOR2_X1    g06615(.A1(new_n6878_), .A2(new_n6883_), .ZN(new_n6884_));
  NOR2_X1    g06616(.A1(new_n6826_), .A2(new_n6884_), .ZN(new_n6885_));
  INV_X1     g06617(.I(new_n6885_), .ZN(new_n6886_));
  NAND2_X1   g06618(.A1(new_n6826_), .A2(new_n6884_), .ZN(new_n6887_));
  AOI21_X1   g06619(.A1(new_n6886_), .A2(new_n6887_), .B(new_n6730_), .ZN(new_n6888_));
  XOR2_X1    g06620(.A1(new_n6825_), .A2(new_n6884_), .Z(new_n6889_));
  NOR2_X1    g06621(.A1(new_n6889_), .A2(new_n6729_), .ZN(new_n6890_));
  NOR2_X1    g06622(.A1(new_n6888_), .A2(new_n6890_), .ZN(new_n6891_));
  NOR2_X1    g06623(.A1(new_n6891_), .A2(new_n6728_), .ZN(new_n6892_));
  NOR3_X1    g06624(.A1(new_n6727_), .A2(new_n6888_), .A3(new_n6890_), .ZN(new_n6893_));
  NOR2_X1    g06625(.A1(new_n6892_), .A2(new_n6893_), .ZN(new_n6894_));
  XOR2_X1    g06626(.A1(new_n6891_), .A2(new_n6728_), .Z(new_n6895_));
  NAND2_X1   g06627(.A1(new_n6895_), .A2(new_n6726_), .ZN(new_n6896_));
  OAI21_X1   g06628(.A1(new_n6726_), .A2(new_n6894_), .B(new_n6896_), .ZN(new_n6897_));
  XOR2_X1    g06629(.A1(new_n6897_), .A2(new_n6678_), .Z(new_n6898_));
  INV_X1     g06630(.I(new_n6678_), .ZN(new_n6899_));
  NAND2_X1   g06631(.A1(new_n6897_), .A2(new_n6899_), .ZN(new_n6900_));
  NOR2_X1    g06632(.A1(new_n6897_), .A2(new_n6899_), .ZN(new_n6901_));
  INV_X1     g06633(.I(new_n6901_), .ZN(new_n6902_));
  NAND2_X1   g06634(.A1(new_n6902_), .A2(new_n6900_), .ZN(new_n6903_));
  NAND2_X1   g06635(.A1(new_n6676_), .A2(new_n6903_), .ZN(new_n6904_));
  OAI21_X1   g06636(.A1(new_n6676_), .A2(new_n6898_), .B(new_n6904_), .ZN(\asquared[55] ));
  OAI21_X1   g06637(.A1(new_n6676_), .A2(new_n6901_), .B(new_n6900_), .ZN(new_n6906_));
  NOR2_X1    g06638(.A1(new_n6893_), .A2(new_n6726_), .ZN(new_n6907_));
  NOR2_X1    g06639(.A1(new_n6907_), .A2(new_n6892_), .ZN(new_n6908_));
  AOI21_X1   g06640(.A1(new_n6679_), .A2(new_n6722_), .B(new_n6720_), .ZN(new_n6909_));
  OAI21_X1   g06641(.A1(new_n6760_), .A2(new_n6792_), .B(new_n6791_), .ZN(new_n6910_));
  AOI21_X1   g06642(.A1(new_n6801_), .A2(new_n6805_), .B(new_n6803_), .ZN(new_n6911_));
  AOI21_X1   g06643(.A1(new_n6843_), .A2(new_n6855_), .B(new_n6854_), .ZN(new_n6912_));
  AOI21_X1   g06644(.A1(new_n3061_), .A2(new_n5173_), .B(new_n6751_), .ZN(new_n6913_));
  NAND2_X1   g06645(.A1(new_n6695_), .A2(new_n3037_), .ZN(new_n6914_));
  NAND2_X1   g06646(.A1(\a[1] ), .A2(\a[54] ), .ZN(new_n6915_));
  XOR2_X1    g06647(.A1(new_n6915_), .A2(\a[28] ), .Z(new_n6916_));
  NOR2_X1    g06648(.A1(new_n6916_), .A2(new_n6914_), .ZN(new_n6917_));
  NAND2_X1   g06649(.A1(new_n6916_), .A2(new_n6914_), .ZN(new_n6918_));
  INV_X1     g06650(.I(new_n6918_), .ZN(new_n6919_));
  OAI21_X1   g06651(.A1(new_n6919_), .A2(new_n6917_), .B(new_n6913_), .ZN(new_n6920_));
  INV_X1     g06652(.I(new_n6913_), .ZN(new_n6921_));
  XOR2_X1    g06653(.A1(new_n6916_), .A2(new_n6914_), .Z(new_n6922_));
  NAND2_X1   g06654(.A1(new_n6922_), .A2(new_n6921_), .ZN(new_n6923_));
  NAND2_X1   g06655(.A1(new_n6923_), .A2(new_n6920_), .ZN(new_n6924_));
  INV_X1     g06656(.I(new_n6924_), .ZN(new_n6925_));
  NOR2_X1    g06657(.A1(new_n6912_), .A2(new_n6925_), .ZN(new_n6926_));
  INV_X1     g06658(.I(new_n6926_), .ZN(new_n6927_));
  NAND2_X1   g06659(.A1(new_n6912_), .A2(new_n6925_), .ZN(new_n6928_));
  AOI21_X1   g06660(.A1(new_n6927_), .A2(new_n6928_), .B(new_n6911_), .ZN(new_n6929_));
  INV_X1     g06661(.I(new_n6911_), .ZN(new_n6930_));
  XOR2_X1    g06662(.A1(new_n6912_), .A2(new_n6924_), .Z(new_n6931_));
  NOR2_X1    g06663(.A1(new_n6931_), .A2(new_n6930_), .ZN(new_n6932_));
  INV_X1     g06664(.I(new_n6739_), .ZN(new_n6933_));
  AOI21_X1   g06665(.A1(new_n267_), .A2(new_n6779_), .B(new_n6778_), .ZN(new_n6934_));
  XNOR2_X1   g06666(.A1(new_n6770_), .A2(new_n6934_), .ZN(new_n6935_));
  AND2_X2    g06667(.A1(new_n6770_), .A2(new_n6934_), .Z(new_n6936_));
  NOR2_X1    g06668(.A1(new_n6770_), .A2(new_n6934_), .ZN(new_n6937_));
  OAI21_X1   g06669(.A1(new_n6936_), .A2(new_n6937_), .B(new_n6933_), .ZN(new_n6938_));
  OAI21_X1   g06670(.A1(new_n6935_), .A2(new_n6933_), .B(new_n6938_), .ZN(new_n6939_));
  INV_X1     g06671(.I(new_n6939_), .ZN(new_n6940_));
  NAND2_X1   g06672(.A1(new_n6710_), .A2(new_n6690_), .ZN(new_n6941_));
  NAND2_X1   g06673(.A1(new_n6941_), .A2(new_n6709_), .ZN(new_n6942_));
  NOR4_X1    g06674(.A1(new_n268_), .A2(new_n359_), .A3(new_n5175_), .A4(new_n5511_), .ZN(new_n6943_));
  INV_X1     g06675(.I(new_n6943_), .ZN(new_n6944_));
  INV_X1     g06676(.I(\a[54] ), .ZN(new_n6945_));
  NOR2_X1    g06677(.A1(new_n199_), .A2(new_n6945_), .ZN(new_n6946_));
  OAI21_X1   g06678(.A1(new_n6696_), .A2(new_n6693_), .B(new_n6946_), .ZN(new_n6947_));
  NAND2_X1   g06679(.A1(new_n6947_), .A2(new_n6697_), .ZN(new_n6948_));
  INV_X1     g06680(.I(new_n6948_), .ZN(new_n6949_));
  NAND2_X1   g06681(.A1(new_n3838_), .A2(new_n2331_), .ZN(new_n6950_));
  NAND2_X1   g06682(.A1(\a[5] ), .A2(\a[50] ), .ZN(new_n6951_));
  XNOR2_X1   g06683(.A1(new_n6950_), .A2(new_n6951_), .ZN(new_n6952_));
  NOR2_X1    g06684(.A1(new_n6949_), .A2(new_n6952_), .ZN(new_n6953_));
  INV_X1     g06685(.I(new_n6952_), .ZN(new_n6954_));
  NOR2_X1    g06686(.A1(new_n6948_), .A2(new_n6954_), .ZN(new_n6955_));
  NOR2_X1    g06687(.A1(new_n6953_), .A2(new_n6955_), .ZN(new_n6956_));
  NOR2_X1    g06688(.A1(new_n6956_), .A2(new_n6944_), .ZN(new_n6957_));
  XOR2_X1    g06689(.A1(new_n6948_), .A2(new_n6952_), .Z(new_n6958_));
  NOR2_X1    g06690(.A1(new_n6958_), .A2(new_n6943_), .ZN(new_n6959_));
  NOR2_X1    g06691(.A1(new_n6957_), .A2(new_n6959_), .ZN(new_n6960_));
  XOR2_X1    g06692(.A1(new_n6942_), .A2(new_n6960_), .Z(new_n6961_));
  AOI21_X1   g06693(.A1(new_n6941_), .A2(new_n6709_), .B(new_n6960_), .ZN(new_n6962_));
  NOR3_X1    g06694(.A1(new_n6942_), .A2(new_n6957_), .A3(new_n6959_), .ZN(new_n6963_));
  OAI21_X1   g06695(.A1(new_n6963_), .A2(new_n6962_), .B(new_n6940_), .ZN(new_n6964_));
  OAI21_X1   g06696(.A1(new_n6961_), .A2(new_n6940_), .B(new_n6964_), .ZN(new_n6965_));
  OAI21_X1   g06697(.A1(new_n6929_), .A2(new_n6932_), .B(new_n6965_), .ZN(new_n6966_));
  NOR2_X1    g06698(.A1(new_n6932_), .A2(new_n6929_), .ZN(new_n6967_));
  INV_X1     g06699(.I(new_n6965_), .ZN(new_n6968_));
  NAND2_X1   g06700(.A1(new_n6968_), .A2(new_n6967_), .ZN(new_n6969_));
  NAND2_X1   g06701(.A1(new_n6969_), .A2(new_n6966_), .ZN(new_n6970_));
  XOR2_X1    g06702(.A1(new_n6965_), .A2(new_n6967_), .Z(new_n6971_));
  NOR2_X1    g06703(.A1(new_n6971_), .A2(new_n6910_), .ZN(new_n6972_));
  AOI21_X1   g06704(.A1(new_n6910_), .A2(new_n6970_), .B(new_n6972_), .ZN(new_n6973_));
  INV_X1     g06705(.I(new_n6716_), .ZN(new_n6974_));
  AOI21_X1   g06706(.A1(new_n6974_), .A2(new_n6683_), .B(new_n6715_), .ZN(new_n6975_));
  AOI21_X1   g06707(.A1(new_n6742_), .A2(new_n6756_), .B(new_n6754_), .ZN(new_n6976_));
  NAND2_X1   g06708(.A1(new_n6775_), .A2(new_n6785_), .ZN(new_n6977_));
  NAND2_X1   g06709(.A1(new_n6977_), .A2(new_n6784_), .ZN(new_n6978_));
  AOI21_X1   g06710(.A1(new_n1769_), .A2(new_n3424_), .B(new_n6686_), .ZN(new_n6979_));
  AOI21_X1   g06711(.A1(new_n1275_), .A2(new_n5600_), .B(new_n6745_), .ZN(new_n6980_));
  NOR2_X1    g06712(.A1(new_n6701_), .A2(new_n6703_), .ZN(new_n6981_));
  XNOR2_X1   g06713(.A1(new_n6980_), .A2(new_n6981_), .ZN(new_n6982_));
  INV_X1     g06714(.I(new_n6980_), .ZN(new_n6983_));
  INV_X1     g06715(.I(new_n6981_), .ZN(new_n6984_));
  NOR2_X1    g06716(.A1(new_n6983_), .A2(new_n6984_), .ZN(new_n6985_));
  NOR2_X1    g06717(.A1(new_n6980_), .A2(new_n6981_), .ZN(new_n6986_));
  NOR2_X1    g06718(.A1(new_n6985_), .A2(new_n6986_), .ZN(new_n6987_));
  MUX2_X1    g06719(.I0(new_n6987_), .I1(new_n6982_), .S(new_n6979_), .Z(new_n6988_));
  XNOR2_X1   g06720(.A1(new_n6978_), .A2(new_n6988_), .ZN(new_n6989_));
  NOR2_X1    g06721(.A1(new_n6978_), .A2(new_n6988_), .ZN(new_n6990_));
  NAND2_X1   g06722(.A1(new_n6978_), .A2(new_n6988_), .ZN(new_n6991_));
  INV_X1     g06723(.I(new_n6991_), .ZN(new_n6992_));
  OAI21_X1   g06724(.A1(new_n6992_), .A2(new_n6990_), .B(new_n6976_), .ZN(new_n6993_));
  OAI21_X1   g06725(.A1(new_n6976_), .A2(new_n6989_), .B(new_n6993_), .ZN(new_n6994_));
  INV_X1     g06726(.I(new_n6994_), .ZN(new_n6995_));
  NOR2_X1    g06727(.A1(new_n6838_), .A2(new_n6829_), .ZN(new_n6996_));
  NOR2_X1    g06728(.A1(new_n6996_), .A2(new_n6836_), .ZN(new_n6997_));
  INV_X1     g06729(.I(new_n6997_), .ZN(new_n6998_));
  INV_X1     g06730(.I(\a[55] ), .ZN(new_n6999_));
  NOR2_X1    g06731(.A1(new_n6260_), .A2(new_n6694_), .ZN(new_n7000_));
  INV_X1     g06732(.I(new_n7000_), .ZN(new_n7001_));
  NOR3_X1    g06733(.A1(new_n1142_), .A2(\a[55] ), .A3(new_n7000_), .ZN(new_n7002_));
  NOR3_X1    g06734(.A1(new_n7002_), .A2(new_n260_), .A3(new_n7001_), .ZN(new_n7003_));
  NOR3_X1    g06735(.A1(new_n7003_), .A2(new_n199_), .A3(new_n6999_), .ZN(new_n7004_));
  NAND2_X1   g06736(.A1(new_n7000_), .A2(new_n4999_), .ZN(new_n7005_));
  NOR2_X1    g06737(.A1(new_n7000_), .A2(new_n4999_), .ZN(new_n7006_));
  AOI21_X1   g06738(.A1(new_n7005_), .A2(new_n7006_), .B(new_n7004_), .ZN(new_n7007_));
  NOR2_X1    g06739(.A1(new_n4530_), .A2(new_n3712_), .ZN(new_n7008_));
  NOR2_X1    g06740(.A1(new_n1711_), .A2(new_n1949_), .ZN(new_n7009_));
  NOR2_X1    g06741(.A1(new_n7008_), .A2(new_n7009_), .ZN(new_n7010_));
  NOR4_X1    g06742(.A1(new_n4372_), .A2(new_n4538_), .A3(new_n1215_), .A4(new_n3423_), .ZN(new_n7011_));
  NAND2_X1   g06743(.A1(new_n7010_), .A2(new_n7011_), .ZN(new_n7012_));
  AOI22_X1   g06744(.A1(new_n1913_), .A2(new_n3981_), .B1(new_n2766_), .B2(new_n2543_), .ZN(new_n7013_));
  INV_X1     g06745(.I(new_n7013_), .ZN(new_n7014_));
  NOR4_X1    g06746(.A1(new_n7014_), .A2(new_n2277_), .A3(new_n3126_), .A4(new_n5852_), .ZN(new_n7015_));
  INV_X1     g06747(.I(new_n7015_), .ZN(new_n7016_));
  NOR2_X1    g06748(.A1(new_n7016_), .A2(new_n7012_), .ZN(new_n7017_));
  INV_X1     g06749(.I(new_n7012_), .ZN(new_n7018_));
  NOR2_X1    g06750(.A1(new_n7018_), .A2(new_n7015_), .ZN(new_n7019_));
  OAI21_X1   g06751(.A1(new_n7017_), .A2(new_n7019_), .B(new_n7007_), .ZN(new_n7020_));
  XOR2_X1    g06752(.A1(new_n7015_), .A2(new_n7012_), .Z(new_n7021_));
  OAI21_X1   g06753(.A1(new_n7007_), .A2(new_n7021_), .B(new_n7020_), .ZN(new_n7022_));
  INV_X1     g06754(.I(new_n4771_), .ZN(new_n7023_));
  NOR2_X1    g06755(.A1(new_n461_), .A2(new_n5004_), .ZN(new_n7024_));
  NOR2_X1    g06756(.A1(new_n7023_), .A2(new_n870_), .ZN(new_n7025_));
  NAND4_X1   g06757(.A1(new_n7025_), .A2(\a[13] ), .A3(new_n6393_), .A4(\a[45] ), .ZN(new_n7026_));
  AOI21_X1   g06758(.A1(new_n7026_), .A2(new_n5743_), .B(new_n796_), .ZN(new_n7027_));
  NOR2_X1    g06759(.A1(new_n7023_), .A2(new_n870_), .ZN(new_n7028_));
  NAND2_X1   g06760(.A1(new_n6030_), .A2(new_n609_), .ZN(new_n7029_));
  XNOR2_X1   g06761(.A1(new_n7029_), .A2(new_n4322_), .ZN(new_n7030_));
  NOR2_X1    g06762(.A1(new_n1916_), .A2(new_n2499_), .ZN(new_n7031_));
  INV_X1     g06763(.I(new_n7031_), .ZN(new_n7032_));
  NOR2_X1    g06764(.A1(new_n7032_), .A2(new_n2692_), .ZN(new_n7033_));
  XOR2_X1    g06765(.A1(new_n7033_), .A2(new_n566_), .Z(new_n7034_));
  XOR2_X1    g06766(.A1(new_n7034_), .A2(\a[43] ), .Z(new_n7035_));
  NOR2_X1    g06767(.A1(new_n7035_), .A2(new_n7030_), .ZN(new_n7036_));
  INV_X1     g06768(.I(new_n7030_), .ZN(new_n7037_));
  INV_X1     g06769(.I(new_n7035_), .ZN(new_n7038_));
  NOR2_X1    g06770(.A1(new_n7038_), .A2(new_n7037_), .ZN(new_n7039_));
  OAI21_X1   g06771(.A1(new_n7039_), .A2(new_n7036_), .B(new_n7028_), .ZN(new_n7040_));
  XOR2_X1    g06772(.A1(new_n7035_), .A2(new_n7037_), .Z(new_n7041_));
  OAI21_X1   g06773(.A1(new_n7028_), .A2(new_n7041_), .B(new_n7040_), .ZN(new_n7042_));
  XOR2_X1    g06774(.A1(new_n7042_), .A2(new_n7022_), .Z(new_n7043_));
  NAND2_X1   g06775(.A1(new_n7042_), .A2(new_n7022_), .ZN(new_n7044_));
  OR2_X2     g06776(.A1(new_n7042_), .A2(new_n7022_), .Z(new_n7045_));
  AOI21_X1   g06777(.A1(new_n7045_), .A2(new_n7044_), .B(new_n6998_), .ZN(new_n7046_));
  AOI21_X1   g06778(.A1(new_n6998_), .A2(new_n7043_), .B(new_n7046_), .ZN(new_n7047_));
  NOR2_X1    g06779(.A1(new_n7047_), .A2(new_n6995_), .ZN(new_n7048_));
  INV_X1     g06780(.I(new_n7048_), .ZN(new_n7049_));
  NAND2_X1   g06781(.A1(new_n7047_), .A2(new_n6995_), .ZN(new_n7050_));
  AOI21_X1   g06782(.A1(new_n7049_), .A2(new_n7050_), .B(new_n6975_), .ZN(new_n7051_));
  XOR2_X1    g06783(.A1(new_n7047_), .A2(new_n6995_), .Z(new_n7052_));
  AOI21_X1   g06784(.A1(new_n6975_), .A2(new_n7052_), .B(new_n7051_), .ZN(new_n7053_));
  XNOR2_X1   g06785(.A1(new_n6973_), .A2(new_n7053_), .ZN(new_n7054_));
  NOR2_X1    g06786(.A1(new_n6973_), .A2(new_n7053_), .ZN(new_n7055_));
  INV_X1     g06787(.I(new_n7055_), .ZN(new_n7056_));
  NAND2_X1   g06788(.A1(new_n6973_), .A2(new_n7053_), .ZN(new_n7057_));
  NAND2_X1   g06789(.A1(new_n7056_), .A2(new_n7057_), .ZN(new_n7058_));
  NAND2_X1   g06790(.A1(new_n7058_), .A2(new_n6909_), .ZN(new_n7059_));
  OAI21_X1   g06791(.A1(new_n6909_), .A2(new_n7054_), .B(new_n7059_), .ZN(new_n7060_));
  OAI21_X1   g06792(.A1(new_n6730_), .A2(new_n6885_), .B(new_n6887_), .ZN(new_n7061_));
  OAI21_X1   g06793(.A1(new_n6731_), .A2(new_n6818_), .B(new_n6820_), .ZN(new_n7062_));
  INV_X1     g06794(.I(new_n7062_), .ZN(new_n7063_));
  NAND2_X1   g06795(.A1(new_n6880_), .A2(new_n6879_), .ZN(new_n7064_));
  NAND2_X1   g06796(.A1(new_n7064_), .A2(new_n6882_), .ZN(new_n7065_));
  NOR2_X1    g06797(.A1(new_n6873_), .A2(new_n6842_), .ZN(new_n7066_));
  NAND2_X1   g06798(.A1(new_n6807_), .A2(new_n6814_), .ZN(new_n7067_));
  NAND2_X1   g06799(.A1(new_n7067_), .A2(new_n6812_), .ZN(new_n7068_));
  NOR2_X1    g06800(.A1(new_n364_), .A2(new_n4414_), .ZN(new_n7069_));
  NAND2_X1   g06801(.A1(\a[14] ), .A2(\a[15] ), .ZN(new_n7070_));
  NOR2_X1    g06802(.A1(new_n6579_), .A2(new_n7070_), .ZN(new_n7071_));
  NAND2_X1   g06803(.A1(\a[15] ), .A2(\a[40] ), .ZN(new_n7072_));
  NOR2_X1    g06804(.A1(new_n650_), .A2(new_n5175_), .ZN(new_n7073_));
  AOI21_X1   g06805(.A1(new_n7069_), .A2(new_n7073_), .B(new_n7071_), .ZN(new_n7074_));
  INV_X1     g06806(.I(new_n7074_), .ZN(new_n7075_));
  AOI22_X1   g06807(.A1(\a[9] ), .A2(\a[14] ), .B1(\a[41] ), .B2(\a[46] ), .ZN(new_n7076_));
  INV_X1     g06808(.I(new_n7076_), .ZN(new_n7077_));
  OAI22_X1   g06809(.A1(new_n7075_), .A2(new_n7077_), .B1(new_n7071_), .B2(new_n7072_), .ZN(new_n7078_));
  NOR2_X1    g06810(.A1(new_n6869_), .A2(new_n6867_), .ZN(new_n7079_));
  NOR2_X1    g06811(.A1(new_n7079_), .A2(new_n6868_), .ZN(new_n7080_));
  NAND4_X1   g06812(.A1(\a[6] ), .A2(\a[17] ), .A3(\a[38] ), .A4(\a[49] ), .ZN(new_n7081_));
  NAND2_X1   g06813(.A1(\a[3] ), .A2(\a[52] ), .ZN(new_n7082_));
  XNOR2_X1   g06814(.A1(new_n7081_), .A2(new_n7082_), .ZN(new_n7083_));
  XNOR2_X1   g06815(.A1(new_n7080_), .A2(new_n7083_), .ZN(new_n7084_));
  NOR2_X1    g06816(.A1(new_n7084_), .A2(new_n7078_), .ZN(new_n7085_));
  INV_X1     g06817(.I(new_n7078_), .ZN(new_n7086_));
  NOR2_X1    g06818(.A1(new_n7080_), .A2(new_n7083_), .ZN(new_n7087_));
  INV_X1     g06819(.I(new_n7087_), .ZN(new_n7088_));
  NAND2_X1   g06820(.A1(new_n7080_), .A2(new_n7083_), .ZN(new_n7089_));
  AOI21_X1   g06821(.A1(new_n7088_), .A2(new_n7089_), .B(new_n7086_), .ZN(new_n7090_));
  NOR2_X1    g06822(.A1(new_n7085_), .A2(new_n7090_), .ZN(new_n7091_));
  XOR2_X1    g06823(.A1(new_n7068_), .A2(new_n7091_), .Z(new_n7092_));
  OAI21_X1   g06824(.A1(new_n6874_), .A2(new_n7066_), .B(new_n7092_), .ZN(new_n7093_));
  NOR2_X1    g06825(.A1(new_n7066_), .A2(new_n6874_), .ZN(new_n7094_));
  NOR2_X1    g06826(.A1(new_n7068_), .A2(new_n7091_), .ZN(new_n7095_));
  NAND2_X1   g06827(.A1(new_n7068_), .A2(new_n7091_), .ZN(new_n7096_));
  INV_X1     g06828(.I(new_n7096_), .ZN(new_n7097_));
  OAI21_X1   g06829(.A1(new_n7097_), .A2(new_n7095_), .B(new_n7094_), .ZN(new_n7098_));
  NAND2_X1   g06830(.A1(new_n7093_), .A2(new_n7098_), .ZN(new_n7099_));
  INV_X1     g06831(.I(new_n7099_), .ZN(new_n7100_));
  NOR2_X1    g06832(.A1(new_n7100_), .A2(new_n7065_), .ZN(new_n7101_));
  INV_X1     g06833(.I(new_n7101_), .ZN(new_n7102_));
  NAND2_X1   g06834(.A1(new_n7100_), .A2(new_n7065_), .ZN(new_n7103_));
  AOI21_X1   g06835(.A1(new_n7102_), .A2(new_n7103_), .B(new_n7063_), .ZN(new_n7104_));
  XOR2_X1    g06836(.A1(new_n7099_), .A2(new_n7065_), .Z(new_n7105_));
  NOR2_X1    g06837(.A1(new_n7105_), .A2(new_n7062_), .ZN(new_n7106_));
  NOR2_X1    g06838(.A1(new_n7104_), .A2(new_n7106_), .ZN(new_n7107_));
  INV_X1     g06839(.I(new_n7107_), .ZN(new_n7108_));
  AND2_X2    g06840(.A1(new_n7061_), .A2(new_n7108_), .Z(new_n7109_));
  NOR2_X1    g06841(.A1(new_n7061_), .A2(new_n7108_), .ZN(new_n7110_));
  OAI21_X1   g06842(.A1(new_n7109_), .A2(new_n7110_), .B(new_n7060_), .ZN(new_n7111_));
  XOR2_X1    g06843(.A1(new_n7061_), .A2(new_n7107_), .Z(new_n7112_));
  OAI21_X1   g06844(.A1(new_n7060_), .A2(new_n7112_), .B(new_n7111_), .ZN(new_n7113_));
  NAND2_X1   g06845(.A1(new_n7113_), .A2(new_n6908_), .ZN(new_n7114_));
  NOR2_X1    g06846(.A1(new_n7113_), .A2(new_n6908_), .ZN(new_n7115_));
  INV_X1     g06847(.I(new_n7115_), .ZN(new_n7116_));
  NAND2_X1   g06848(.A1(new_n7116_), .A2(new_n7114_), .ZN(new_n7117_));
  XOR2_X1    g06849(.A1(new_n6906_), .A2(new_n7117_), .Z(\asquared[56] ));
  NOR2_X1    g06850(.A1(new_n7115_), .A2(new_n6897_), .ZN(new_n7119_));
  AOI21_X1   g06851(.A1(new_n7115_), .A2(new_n6897_), .B(new_n6899_), .ZN(new_n7120_));
  NOR2_X1    g06852(.A1(new_n7120_), .A2(new_n7119_), .ZN(new_n7121_));
  NAND2_X1   g06853(.A1(new_n6675_), .A2(new_n7121_), .ZN(new_n7122_));
  NOR2_X1    g06854(.A1(new_n7060_), .A2(new_n7110_), .ZN(new_n7123_));
  NOR2_X1    g06855(.A1(new_n7123_), .A2(new_n7109_), .ZN(new_n7124_));
  OAI21_X1   g06856(.A1(new_n7063_), .A2(new_n7101_), .B(new_n7103_), .ZN(new_n7125_));
  INV_X1     g06857(.I(new_n7125_), .ZN(new_n7126_));
  NAND4_X1   g06858(.A1(new_n4539_), .A2(\a[33] ), .A3(\a[34] ), .A4(\a[36] ), .ZN(new_n7127_));
  INV_X1     g06859(.I(new_n7127_), .ZN(new_n7128_));
  NOR3_X1    g06860(.A1(new_n4728_), .A2(new_n1949_), .A3(new_n2285_), .ZN(new_n7129_));
  NOR2_X1    g06861(.A1(new_n7128_), .A2(new_n7129_), .ZN(new_n7130_));
  NOR2_X1    g06862(.A1(new_n2368_), .A2(new_n2868_), .ZN(new_n7131_));
  INV_X1     g06863(.I(new_n7130_), .ZN(new_n7132_));
  AOI21_X1   g06864(.A1(new_n2286_), .A2(new_n4372_), .B(new_n7132_), .ZN(new_n7133_));
  AOI21_X1   g06865(.A1(new_n7133_), .A2(new_n7131_), .B(\a[34] ), .ZN(new_n7134_));
  OR2_X2     g06866(.A1(new_n7134_), .A2(new_n1674_), .Z(new_n7135_));
  NOR2_X1    g06867(.A1(\a[20] ), .A2(\a[36] ), .ZN(new_n7136_));
  AOI21_X1   g06868(.A1(new_n7135_), .A2(new_n7136_), .B(new_n7130_), .ZN(new_n7137_));
  INV_X1     g06869(.I(new_n7137_), .ZN(new_n7138_));
  INV_X1     g06870(.I(new_n7073_), .ZN(new_n7139_));
  NOR2_X1    g06871(.A1(new_n6394_), .A2(new_n7139_), .ZN(new_n7140_));
  INV_X1     g06872(.I(new_n6147_), .ZN(new_n7141_));
  NOR3_X1    g06873(.A1(new_n7141_), .A2(new_n650_), .A3(new_n5511_), .ZN(new_n7142_));
  NAND2_X1   g06874(.A1(new_n7142_), .A2(new_n7140_), .ZN(new_n7143_));
  AOI21_X1   g06875(.A1(new_n7143_), .A2(new_n5793_), .B(new_n525_), .ZN(new_n7144_));
  NOR3_X1    g06876(.A1(new_n7144_), .A2(new_n364_), .A3(new_n5511_), .ZN(new_n7145_));
  NOR2_X1    g06877(.A1(new_n7144_), .A2(new_n7140_), .ZN(new_n7146_));
  INV_X1     g06878(.I(new_n7146_), .ZN(new_n7147_));
  NOR3_X1    g06879(.A1(new_n7147_), .A2(new_n5180_), .A3(new_n6773_), .ZN(new_n7148_));
  INV_X1     g06880(.I(new_n2749_), .ZN(new_n7149_));
  OAI21_X1   g06881(.A1(new_n3849_), .A2(new_n4184_), .B(new_n7149_), .ZN(new_n7150_));
  NOR2_X1    g06882(.A1(new_n1691_), .A2(new_n2765_), .ZN(new_n7151_));
  INV_X1     g06883(.I(new_n7151_), .ZN(new_n7152_));
  NOR4_X1    g06884(.A1(new_n7150_), .A2(new_n2752_), .A3(new_n3126_), .A4(new_n7152_), .ZN(new_n7153_));
  INV_X1     g06885(.I(new_n7153_), .ZN(new_n7154_));
  NOR3_X1    g06886(.A1(new_n7148_), .A2(new_n7145_), .A3(new_n7154_), .ZN(new_n7155_));
  NOR2_X1    g06887(.A1(new_n7148_), .A2(new_n7145_), .ZN(new_n7156_));
  NOR2_X1    g06888(.A1(new_n7156_), .A2(new_n7153_), .ZN(new_n7157_));
  NOR2_X1    g06889(.A1(new_n7157_), .A2(new_n7155_), .ZN(new_n7158_));
  NOR2_X1    g06890(.A1(new_n7138_), .A2(new_n7158_), .ZN(new_n7159_));
  XOR2_X1    g06891(.A1(new_n7156_), .A2(new_n7154_), .Z(new_n7160_));
  INV_X1     g06892(.I(new_n7160_), .ZN(new_n7161_));
  AOI21_X1   g06893(.A1(new_n7161_), .A2(new_n7138_), .B(new_n7159_), .ZN(new_n7162_));
  NAND2_X1   g06894(.A1(\a[15] ), .A2(\a[48] ), .ZN(new_n7163_));
  NOR3_X1    g06895(.A1(new_n7163_), .A2(new_n359_), .A3(new_n4414_), .ZN(new_n7164_));
  INV_X1     g06896(.I(new_n1722_), .ZN(new_n7165_));
  NOR3_X1    g06897(.A1(new_n7165_), .A2(new_n4240_), .A3(new_n5750_), .ZN(new_n7166_));
  NAND2_X1   g06898(.A1(new_n7166_), .A2(new_n7164_), .ZN(new_n7167_));
  AOI21_X1   g06899(.A1(new_n7167_), .A2(new_n6579_), .B(new_n1021_), .ZN(new_n7168_));
  NOR2_X1    g06900(.A1(new_n7168_), .A2(new_n7164_), .ZN(new_n7169_));
  INV_X1     g06901(.I(new_n7169_), .ZN(new_n7170_));
  NAND2_X1   g06902(.A1(\a[41] ), .A2(\a[48] ), .ZN(new_n7171_));
  OAI21_X1   g06903(.A1(new_n359_), .A2(new_n875_), .B(new_n7171_), .ZN(new_n7172_));
  OAI22_X1   g06904(.A1(new_n7170_), .A2(new_n7172_), .B1(new_n4721_), .B2(new_n7168_), .ZN(new_n7173_));
  NAND2_X1   g06905(.A1(\a[17] ), .A2(\a[50] ), .ZN(new_n7174_));
  NOR3_X1    g06906(.A1(new_n7174_), .A2(new_n242_), .A3(new_n3783_), .ZN(new_n7175_));
  AOI21_X1   g06907(.A1(new_n479_), .A2(new_n6280_), .B(new_n7175_), .ZN(new_n7176_));
  NOR2_X1    g06908(.A1(new_n268_), .A2(new_n5745_), .ZN(new_n7177_));
  NOR2_X1    g06909(.A1(new_n885_), .A2(new_n3783_), .ZN(new_n7178_));
  XNOR2_X1   g06910(.A1(new_n7177_), .A2(new_n7178_), .ZN(new_n7179_));
  NOR2_X1    g06911(.A1(new_n7179_), .A2(new_n7177_), .ZN(new_n7180_));
  NOR2_X1    g06912(.A1(new_n7176_), .A2(new_n7180_), .ZN(new_n7181_));
  OAI21_X1   g06913(.A1(new_n242_), .A2(new_n6055_), .B(new_n7179_), .ZN(new_n7182_));
  INV_X1     g06914(.I(new_n7182_), .ZN(new_n7183_));
  NOR2_X1    g06915(.A1(new_n7183_), .A2(new_n7181_), .ZN(new_n7184_));
  INV_X1     g06916(.I(new_n7184_), .ZN(new_n7185_));
  NOR2_X1    g06917(.A1(new_n4501_), .A2(new_n5004_), .ZN(new_n7186_));
  INV_X1     g06918(.I(new_n7186_), .ZN(new_n7187_));
  NOR2_X1    g06919(.A1(new_n7187_), .A2(new_n5743_), .ZN(new_n7188_));
  NOR2_X1    g06920(.A1(new_n7188_), .A2(new_n2668_), .ZN(new_n7189_));
  NOR2_X1    g06921(.A1(new_n5322_), .A2(new_n1150_), .ZN(new_n7190_));
  AOI21_X1   g06922(.A1(\a[12] ), .A2(\a[44] ), .B(new_n6136_), .ZN(new_n7191_));
  NOR4_X1    g06923(.A1(new_n7190_), .A2(new_n675_), .A3(new_n7191_), .A4(new_n5004_), .ZN(new_n7192_));
  NAND2_X1   g06924(.A1(new_n7192_), .A2(new_n7189_), .ZN(new_n7193_));
  NOR2_X1    g06925(.A1(new_n7185_), .A2(new_n7193_), .ZN(new_n7194_));
  INV_X1     g06926(.I(new_n7194_), .ZN(new_n7195_));
  NAND2_X1   g06927(.A1(new_n7185_), .A2(new_n7193_), .ZN(new_n7196_));
  AOI21_X1   g06928(.A1(new_n7195_), .A2(new_n7196_), .B(new_n7173_), .ZN(new_n7197_));
  XNOR2_X1   g06929(.A1(new_n7184_), .A2(new_n7193_), .ZN(new_n7198_));
  AOI21_X1   g06930(.A1(new_n7173_), .A2(new_n7198_), .B(new_n7197_), .ZN(new_n7199_));
  NAND2_X1   g06931(.A1(new_n6030_), .A2(new_n609_), .ZN(new_n7200_));
  NOR2_X1    g06932(.A1(new_n6030_), .A2(new_n609_), .ZN(new_n7201_));
  NOR2_X1    g06933(.A1(\a[16] ), .A2(\a[39] ), .ZN(new_n7202_));
  AOI21_X1   g06934(.A1(new_n7200_), .A2(new_n7202_), .B(new_n7201_), .ZN(new_n7203_));
  NOR2_X1    g06935(.A1(new_n6692_), .A2(new_n6694_), .ZN(new_n7204_));
  NOR2_X1    g06936(.A1(new_n3837_), .A2(new_n6694_), .ZN(new_n7205_));
  AOI22_X1   g06937(.A1(new_n1340_), .A2(new_n7204_), .B1(new_n7205_), .B2(new_n267_), .ZN(new_n7206_));
  INV_X1     g06938(.I(new_n7206_), .ZN(new_n7207_));
  NOR2_X1    g06939(.A1(new_n282_), .A2(new_n6692_), .ZN(new_n7208_));
  NOR2_X1    g06940(.A1(new_n1339_), .A2(new_n3837_), .ZN(new_n7209_));
  XNOR2_X1   g06941(.A1(new_n7208_), .A2(new_n7209_), .ZN(new_n7210_));
  NOR2_X1    g06942(.A1(new_n7210_), .A2(new_n7208_), .ZN(new_n7211_));
  NOR2_X1    g06943(.A1(new_n7207_), .A2(new_n7211_), .ZN(new_n7212_));
  OAI21_X1   g06944(.A1(new_n200_), .A2(new_n6694_), .B(new_n7210_), .ZN(new_n7213_));
  INV_X1     g06945(.I(new_n7213_), .ZN(new_n7214_));
  NOR2_X1    g06946(.A1(new_n7214_), .A2(new_n7212_), .ZN(new_n7215_));
  INV_X1     g06947(.I(\a[56] ), .ZN(new_n7216_));
  NOR2_X1    g06948(.A1(new_n201_), .A2(new_n7216_), .ZN(new_n7217_));
  XNOR2_X1   g06949(.A1(new_n6946_), .A2(new_n7217_), .ZN(new_n7218_));
  NOR2_X1    g06950(.A1(new_n2178_), .A2(new_n6945_), .ZN(new_n7219_));
  NAND2_X1   g06951(.A1(new_n7219_), .A2(\a[1] ), .ZN(new_n7220_));
  INV_X1     g06952(.I(new_n7220_), .ZN(new_n7221_));
  XOR2_X1    g06953(.A1(new_n7218_), .A2(new_n7221_), .Z(new_n7222_));
  NOR2_X1    g06954(.A1(new_n7215_), .A2(new_n7222_), .ZN(new_n7223_));
  AND2_X2    g06955(.A1(new_n7215_), .A2(new_n7222_), .Z(new_n7224_));
  OAI21_X1   g06956(.A1(new_n7224_), .A2(new_n7223_), .B(new_n7203_), .ZN(new_n7225_));
  INV_X1     g06957(.I(new_n7203_), .ZN(new_n7226_));
  XOR2_X1    g06958(.A1(new_n7215_), .A2(new_n7222_), .Z(new_n7227_));
  NAND2_X1   g06959(.A1(new_n7227_), .A2(new_n7226_), .ZN(new_n7228_));
  NAND2_X1   g06960(.A1(new_n7228_), .A2(new_n7225_), .ZN(new_n7229_));
  XOR2_X1    g06961(.A1(new_n7199_), .A2(new_n7229_), .Z(new_n7230_));
  INV_X1     g06962(.I(new_n7229_), .ZN(new_n7231_));
  NOR2_X1    g06963(.A1(new_n7199_), .A2(new_n7231_), .ZN(new_n7232_));
  NAND2_X1   g06964(.A1(new_n7199_), .A2(new_n7231_), .ZN(new_n7233_));
  INV_X1     g06965(.I(new_n7233_), .ZN(new_n7234_));
  OAI21_X1   g06966(.A1(new_n7234_), .A2(new_n7232_), .B(new_n7162_), .ZN(new_n7235_));
  OAI21_X1   g06967(.A1(new_n7162_), .A2(new_n7230_), .B(new_n7235_), .ZN(new_n7236_));
  OAI21_X1   g06968(.A1(new_n7094_), .A2(new_n7095_), .B(new_n7096_), .ZN(new_n7237_));
  INV_X1     g06969(.I(new_n7039_), .ZN(new_n7238_));
  AOI21_X1   g06970(.A1(new_n7238_), .A2(new_n7028_), .B(new_n7036_), .ZN(new_n7239_));
  INV_X1     g06971(.I(new_n7239_), .ZN(new_n7240_));
  NOR2_X1    g06972(.A1(new_n7027_), .A2(new_n7025_), .ZN(new_n7241_));
  NOR2_X1    g06973(.A1(new_n566_), .A2(new_n4501_), .ZN(new_n7242_));
  OAI21_X1   g06974(.A1(new_n2797_), .A2(new_n7031_), .B(new_n7242_), .ZN(new_n7243_));
  OAI21_X1   g06975(.A1(new_n2692_), .A2(new_n7032_), .B(new_n7243_), .ZN(new_n7244_));
  NOR2_X1    g06976(.A1(new_n194_), .A2(new_n6999_), .ZN(new_n7245_));
  XNOR2_X1   g06977(.A1(new_n2500_), .A2(new_n7245_), .ZN(new_n7246_));
  XOR2_X1    g06978(.A1(new_n7244_), .A2(new_n7246_), .Z(new_n7247_));
  NAND2_X1   g06979(.A1(new_n7247_), .A2(new_n7241_), .ZN(new_n7248_));
  INV_X1     g06980(.I(new_n7241_), .ZN(new_n7249_));
  NOR2_X1    g06981(.A1(new_n7244_), .A2(new_n7246_), .ZN(new_n7250_));
  NAND2_X1   g06982(.A1(new_n7244_), .A2(new_n7246_), .ZN(new_n7251_));
  INV_X1     g06983(.I(new_n7251_), .ZN(new_n7252_));
  OAI21_X1   g06984(.A1(new_n7250_), .A2(new_n7252_), .B(new_n7249_), .ZN(new_n7253_));
  NAND2_X1   g06985(.A1(new_n7253_), .A2(new_n7248_), .ZN(new_n7254_));
  NAND4_X1   g06986(.A1(\a[6] ), .A2(\a[17] ), .A3(\a[38] ), .A4(\a[49] ), .ZN(new_n7255_));
  AOI22_X1   g06987(.A1(\a[6] ), .A2(\a[17] ), .B1(\a[38] ), .B2(\a[49] ), .ZN(new_n7256_));
  NOR2_X1    g06988(.A1(\a[3] ), .A2(\a[52] ), .ZN(new_n7257_));
  AOI21_X1   g06989(.A1(new_n7255_), .A2(new_n7257_), .B(new_n7256_), .ZN(new_n7258_));
  AOI21_X1   g06990(.A1(new_n4538_), .A2(new_n4372_), .B(new_n7010_), .ZN(new_n7259_));
  AOI21_X1   g06991(.A1(new_n2277_), .A2(new_n3126_), .B(new_n7013_), .ZN(new_n7260_));
  INV_X1     g06992(.I(new_n7260_), .ZN(new_n7261_));
  XOR2_X1    g06993(.A1(new_n7259_), .A2(new_n7261_), .Z(new_n7262_));
  INV_X1     g06994(.I(new_n7259_), .ZN(new_n7263_));
  NOR2_X1    g06995(.A1(new_n7263_), .A2(new_n7261_), .ZN(new_n7264_));
  NOR2_X1    g06996(.A1(new_n7259_), .A2(new_n7260_), .ZN(new_n7265_));
  NOR2_X1    g06997(.A1(new_n7264_), .A2(new_n7265_), .ZN(new_n7266_));
  MUX2_X1    g06998(.I0(new_n7266_), .I1(new_n7262_), .S(new_n7258_), .Z(new_n7267_));
  XNOR2_X1   g06999(.A1(new_n7267_), .A2(new_n7254_), .ZN(new_n7268_));
  NAND2_X1   g07000(.A1(new_n7268_), .A2(new_n7240_), .ZN(new_n7269_));
  INV_X1     g07001(.I(new_n7254_), .ZN(new_n7270_));
  NOR2_X1    g07002(.A1(new_n7270_), .A2(new_n7267_), .ZN(new_n7271_));
  NAND2_X1   g07003(.A1(new_n7270_), .A2(new_n7267_), .ZN(new_n7272_));
  INV_X1     g07004(.I(new_n7272_), .ZN(new_n7273_));
  OAI21_X1   g07005(.A1(new_n7273_), .A2(new_n7271_), .B(new_n7239_), .ZN(new_n7274_));
  NAND2_X1   g07006(.A1(new_n7269_), .A2(new_n7274_), .ZN(new_n7275_));
  XNOR2_X1   g07007(.A1(new_n7237_), .A2(new_n7275_), .ZN(new_n7276_));
  INV_X1     g07008(.I(new_n7275_), .ZN(new_n7277_));
  NOR2_X1    g07009(.A1(new_n7277_), .A2(new_n7237_), .ZN(new_n7278_));
  INV_X1     g07010(.I(new_n7278_), .ZN(new_n7279_));
  NAND2_X1   g07011(.A1(new_n7277_), .A2(new_n7237_), .ZN(new_n7280_));
  AOI21_X1   g07012(.A1(new_n7279_), .A2(new_n7280_), .B(new_n7236_), .ZN(new_n7281_));
  AOI21_X1   g07013(.A1(new_n7236_), .A2(new_n7276_), .B(new_n7281_), .ZN(new_n7282_));
  AOI21_X1   g07014(.A1(new_n6930_), .A2(new_n6928_), .B(new_n6926_), .ZN(new_n7283_));
  NOR2_X1    g07015(.A1(new_n3838_), .A2(new_n2331_), .ZN(new_n7284_));
  NAND2_X1   g07016(.A1(new_n353_), .A2(new_n6055_), .ZN(new_n7285_));
  AOI21_X1   g07017(.A1(new_n2331_), .A2(new_n3838_), .B(new_n7285_), .ZN(new_n7286_));
  NOR2_X1    g07018(.A1(new_n7286_), .A2(new_n7284_), .ZN(new_n7287_));
  XOR2_X1    g07019(.A1(new_n7074_), .A2(new_n7287_), .Z(new_n7288_));
  NAND2_X1   g07020(.A1(new_n7288_), .A2(new_n7005_), .ZN(new_n7289_));
  INV_X1     g07021(.I(new_n7005_), .ZN(new_n7290_));
  NOR3_X1    g07022(.A1(new_n7075_), .A2(new_n7284_), .A3(new_n7286_), .ZN(new_n7291_));
  NOR2_X1    g07023(.A1(new_n7074_), .A2(new_n7287_), .ZN(new_n7292_));
  OAI21_X1   g07024(.A1(new_n7291_), .A2(new_n7292_), .B(new_n7290_), .ZN(new_n7293_));
  NAND2_X1   g07025(.A1(new_n7289_), .A2(new_n7293_), .ZN(new_n7294_));
  NAND2_X1   g07026(.A1(new_n7089_), .A2(new_n7086_), .ZN(new_n7295_));
  NAND2_X1   g07027(.A1(new_n7295_), .A2(new_n7088_), .ZN(new_n7296_));
  XOR2_X1    g07028(.A1(new_n7296_), .A2(new_n7294_), .Z(new_n7297_));
  NOR2_X1    g07029(.A1(new_n7297_), .A2(new_n7283_), .ZN(new_n7298_));
  INV_X1     g07030(.I(new_n7283_), .ZN(new_n7299_));
  INV_X1     g07031(.I(new_n7296_), .ZN(new_n7300_));
  NOR2_X1    g07032(.A1(new_n7300_), .A2(new_n7294_), .ZN(new_n7301_));
  INV_X1     g07033(.I(new_n7301_), .ZN(new_n7302_));
  NAND2_X1   g07034(.A1(new_n7300_), .A2(new_n7294_), .ZN(new_n7303_));
  AOI21_X1   g07035(.A1(new_n7302_), .A2(new_n7303_), .B(new_n7299_), .ZN(new_n7304_));
  NOR2_X1    g07036(.A1(new_n7304_), .A2(new_n7298_), .ZN(new_n7305_));
  INV_X1     g07037(.I(new_n7305_), .ZN(new_n7306_));
  INV_X1     g07038(.I(new_n7019_), .ZN(new_n7307_));
  AOI21_X1   g07039(.A1(new_n7307_), .A2(new_n7007_), .B(new_n7017_), .ZN(new_n7308_));
  INV_X1     g07040(.I(new_n6986_), .ZN(new_n7309_));
  AOI21_X1   g07041(.A1(new_n6979_), .A2(new_n7309_), .B(new_n6985_), .ZN(new_n7310_));
  NOR2_X1    g07042(.A1(new_n6955_), .A2(new_n6944_), .ZN(new_n7311_));
  NOR2_X1    g07043(.A1(new_n7311_), .A2(new_n6953_), .ZN(new_n7312_));
  XNOR2_X1   g07044(.A1(new_n7312_), .A2(new_n7310_), .ZN(new_n7313_));
  NOR2_X1    g07045(.A1(new_n7313_), .A2(new_n7308_), .ZN(new_n7314_));
  INV_X1     g07046(.I(new_n7308_), .ZN(new_n7315_));
  NOR2_X1    g07047(.A1(new_n7312_), .A2(new_n7310_), .ZN(new_n7316_));
  INV_X1     g07048(.I(new_n7316_), .ZN(new_n7317_));
  NAND2_X1   g07049(.A1(new_n7312_), .A2(new_n7310_), .ZN(new_n7318_));
  AOI21_X1   g07050(.A1(new_n7317_), .A2(new_n7318_), .B(new_n7315_), .ZN(new_n7319_));
  NOR2_X1    g07051(.A1(new_n7314_), .A2(new_n7319_), .ZN(new_n7320_));
  NAND2_X1   g07052(.A1(new_n7045_), .A2(new_n6998_), .ZN(new_n7321_));
  NAND2_X1   g07053(.A1(new_n7321_), .A2(new_n7044_), .ZN(new_n7322_));
  AND2_X2    g07054(.A1(new_n7322_), .A2(new_n7320_), .Z(new_n7323_));
  NOR2_X1    g07055(.A1(new_n7322_), .A2(new_n7320_), .ZN(new_n7324_));
  OAI21_X1   g07056(.A1(new_n7323_), .A2(new_n7324_), .B(new_n7306_), .ZN(new_n7325_));
  XOR2_X1    g07057(.A1(new_n7322_), .A2(new_n7320_), .Z(new_n7326_));
  NAND2_X1   g07058(.A1(new_n7326_), .A2(new_n7305_), .ZN(new_n7327_));
  NAND2_X1   g07059(.A1(new_n7327_), .A2(new_n7325_), .ZN(new_n7328_));
  AND2_X2    g07060(.A1(new_n7328_), .A2(new_n7282_), .Z(new_n7329_));
  NOR2_X1    g07061(.A1(new_n7328_), .A2(new_n7282_), .ZN(new_n7330_));
  NOR2_X1    g07062(.A1(new_n7329_), .A2(new_n7330_), .ZN(new_n7331_));
  NOR2_X1    g07063(.A1(new_n7331_), .A2(new_n7126_), .ZN(new_n7332_));
  XNOR2_X1   g07064(.A1(new_n7328_), .A2(new_n7282_), .ZN(new_n7333_));
  NOR2_X1    g07065(.A1(new_n7333_), .A2(new_n7125_), .ZN(new_n7334_));
  NOR2_X1    g07066(.A1(new_n7332_), .A2(new_n7334_), .ZN(new_n7335_));
  INV_X1     g07067(.I(new_n7335_), .ZN(new_n7336_));
  INV_X1     g07068(.I(new_n6909_), .ZN(new_n7337_));
  NAND2_X1   g07069(.A1(new_n7057_), .A2(new_n7337_), .ZN(new_n7338_));
  NAND2_X1   g07070(.A1(new_n7338_), .A2(new_n7056_), .ZN(new_n7339_));
  OAI21_X1   g07071(.A1(new_n6976_), .A2(new_n6990_), .B(new_n6991_), .ZN(new_n7340_));
  NOR2_X1    g07072(.A1(new_n6963_), .A2(new_n6939_), .ZN(new_n7341_));
  NOR2_X1    g07073(.A1(new_n7341_), .A2(new_n6962_), .ZN(new_n7342_));
  NOR2_X1    g07074(.A1(new_n6933_), .A2(new_n6937_), .ZN(new_n7343_));
  NOR2_X1    g07075(.A1(new_n7343_), .A2(new_n6936_), .ZN(new_n7344_));
  OAI21_X1   g07076(.A1(new_n6921_), .A2(new_n6917_), .B(new_n6918_), .ZN(new_n7345_));
  NAND2_X1   g07077(.A1(\a[38] ), .A2(\a[51] ), .ZN(new_n7346_));
  NOR2_X1    g07078(.A1(new_n1532_), .A2(new_n7346_), .ZN(new_n7347_));
  NAND2_X1   g07079(.A1(\a[21] ), .A2(\a[35] ), .ZN(new_n7348_));
  XOR2_X1    g07080(.A1(new_n7347_), .A2(new_n7348_), .Z(new_n7349_));
  XOR2_X1    g07081(.A1(new_n7345_), .A2(new_n7349_), .Z(new_n7350_));
  INV_X1     g07082(.I(new_n7345_), .ZN(new_n7351_));
  NOR2_X1    g07083(.A1(new_n7351_), .A2(new_n7349_), .ZN(new_n7352_));
  NAND2_X1   g07084(.A1(new_n7351_), .A2(new_n7349_), .ZN(new_n7353_));
  INV_X1     g07085(.I(new_n7353_), .ZN(new_n7354_));
  OAI21_X1   g07086(.A1(new_n7352_), .A2(new_n7354_), .B(new_n7344_), .ZN(new_n7355_));
  OAI21_X1   g07087(.A1(new_n7344_), .A2(new_n7350_), .B(new_n7355_), .ZN(new_n7356_));
  XNOR2_X1   g07088(.A1(new_n7342_), .A2(new_n7356_), .ZN(new_n7357_));
  INV_X1     g07089(.I(new_n7357_), .ZN(new_n7358_));
  NAND2_X1   g07090(.A1(new_n7342_), .A2(new_n7356_), .ZN(new_n7359_));
  NOR2_X1    g07091(.A1(new_n7342_), .A2(new_n7356_), .ZN(new_n7360_));
  INV_X1     g07092(.I(new_n7360_), .ZN(new_n7361_));
  AOI21_X1   g07093(.A1(new_n7361_), .A2(new_n7359_), .B(new_n7340_), .ZN(new_n7362_));
  AOI21_X1   g07094(.A1(new_n7358_), .A2(new_n7340_), .B(new_n7362_), .ZN(new_n7363_));
  NAND2_X1   g07095(.A1(new_n6969_), .A2(new_n6910_), .ZN(new_n7364_));
  NAND2_X1   g07096(.A1(new_n7364_), .A2(new_n6966_), .ZN(new_n7365_));
  OAI21_X1   g07097(.A1(new_n6975_), .A2(new_n7048_), .B(new_n7050_), .ZN(new_n7366_));
  NAND2_X1   g07098(.A1(new_n7365_), .A2(new_n7366_), .ZN(new_n7367_));
  NOR2_X1    g07099(.A1(new_n7365_), .A2(new_n7366_), .ZN(new_n7368_));
  INV_X1     g07100(.I(new_n7368_), .ZN(new_n7369_));
  AOI21_X1   g07101(.A1(new_n7369_), .A2(new_n7367_), .B(new_n7363_), .ZN(new_n7370_));
  INV_X1     g07102(.I(new_n7363_), .ZN(new_n7371_));
  XNOR2_X1   g07103(.A1(new_n7365_), .A2(new_n7366_), .ZN(new_n7372_));
  NOR2_X1    g07104(.A1(new_n7372_), .A2(new_n7371_), .ZN(new_n7373_));
  NOR2_X1    g07105(.A1(new_n7373_), .A2(new_n7370_), .ZN(new_n7374_));
  XOR2_X1    g07106(.A1(new_n7374_), .A2(new_n7339_), .Z(new_n7375_));
  NOR2_X1    g07107(.A1(new_n7374_), .A2(new_n7339_), .ZN(new_n7376_));
  INV_X1     g07108(.I(new_n7376_), .ZN(new_n7377_));
  NAND2_X1   g07109(.A1(new_n7374_), .A2(new_n7339_), .ZN(new_n7378_));
  AOI21_X1   g07110(.A1(new_n7377_), .A2(new_n7378_), .B(new_n7336_), .ZN(new_n7379_));
  AOI21_X1   g07111(.A1(new_n7336_), .A2(new_n7375_), .B(new_n7379_), .ZN(new_n7380_));
  NOR2_X1    g07112(.A1(new_n7380_), .A2(new_n7124_), .ZN(new_n7381_));
  XOR2_X1    g07113(.A1(new_n7122_), .A2(new_n7381_), .Z(new_n7382_));
  XOR2_X1    g07114(.A1(new_n7382_), .A2(new_n7114_), .Z(\asquared[57] ));
  INV_X1     g07115(.I(new_n7381_), .ZN(new_n7384_));
  AOI21_X1   g07116(.A1(new_n7124_), .A2(new_n7380_), .B(new_n7114_), .ZN(new_n7385_));
  NAND3_X1   g07117(.A1(new_n6675_), .A2(new_n7121_), .A3(new_n7385_), .ZN(new_n7386_));
  NAND2_X1   g07118(.A1(new_n7386_), .A2(new_n7384_), .ZN(new_n7387_));
  OAI21_X1   g07119(.A1(new_n7335_), .A2(new_n7376_), .B(new_n7378_), .ZN(new_n7388_));
  INV_X1     g07120(.I(new_n7329_), .ZN(new_n7389_));
  AOI21_X1   g07121(.A1(new_n7389_), .A2(new_n7125_), .B(new_n7330_), .ZN(new_n7390_));
  OAI21_X1   g07122(.A1(new_n7371_), .A2(new_n7368_), .B(new_n7367_), .ZN(new_n7391_));
  INV_X1     g07123(.I(new_n7391_), .ZN(new_n7392_));
  NOR2_X1    g07124(.A1(new_n7138_), .A2(new_n7157_), .ZN(new_n7393_));
  NOR2_X1    g07125(.A1(new_n7393_), .A2(new_n7155_), .ZN(new_n7394_));
  OAI21_X1   g07126(.A1(new_n7249_), .A2(new_n7250_), .B(new_n7251_), .ZN(new_n7395_));
  NOR2_X1    g07127(.A1(new_n7223_), .A2(new_n7226_), .ZN(new_n7396_));
  NOR2_X1    g07128(.A1(new_n7396_), .A2(new_n7224_), .ZN(new_n7397_));
  XOR2_X1    g07129(.A1(new_n7397_), .A2(new_n7395_), .Z(new_n7398_));
  NOR2_X1    g07130(.A1(new_n7394_), .A2(new_n7398_), .ZN(new_n7399_));
  INV_X1     g07131(.I(new_n7395_), .ZN(new_n7400_));
  NOR2_X1    g07132(.A1(new_n7397_), .A2(new_n7400_), .ZN(new_n7401_));
  INV_X1     g07133(.I(new_n7401_), .ZN(new_n7402_));
  NAND2_X1   g07134(.A1(new_n7397_), .A2(new_n7400_), .ZN(new_n7403_));
  NAND2_X1   g07135(.A1(new_n7402_), .A2(new_n7403_), .ZN(new_n7404_));
  AOI21_X1   g07136(.A1(new_n7394_), .A2(new_n7404_), .B(new_n7399_), .ZN(new_n7405_));
  NOR2_X1    g07137(.A1(new_n7234_), .A2(new_n7162_), .ZN(new_n7406_));
  INV_X1     g07138(.I(new_n7173_), .ZN(new_n7407_));
  AOI21_X1   g07139(.A1(new_n7407_), .A2(new_n7196_), .B(new_n7194_), .ZN(new_n7408_));
  INV_X1     g07140(.I(new_n7408_), .ZN(new_n7409_));
  NAND2_X1   g07141(.A1(new_n7177_), .A2(new_n7178_), .ZN(new_n7410_));
  AND2_X2    g07142(.A1(new_n7176_), .A2(new_n7410_), .Z(new_n7411_));
  OAI21_X1   g07143(.A1(new_n2753_), .A2(new_n3127_), .B(new_n7150_), .ZN(new_n7412_));
  XOR2_X1    g07144(.A1(new_n7169_), .A2(new_n7412_), .Z(new_n7413_));
  INV_X1     g07145(.I(new_n7413_), .ZN(new_n7414_));
  NOR2_X1    g07146(.A1(new_n7170_), .A2(new_n7412_), .ZN(new_n7415_));
  INV_X1     g07147(.I(new_n7415_), .ZN(new_n7416_));
  NAND2_X1   g07148(.A1(new_n7170_), .A2(new_n7412_), .ZN(new_n7417_));
  AOI21_X1   g07149(.A1(new_n7416_), .A2(new_n7417_), .B(new_n7411_), .ZN(new_n7418_));
  AOI21_X1   g07150(.A1(new_n7411_), .A2(new_n7414_), .B(new_n7418_), .ZN(new_n7419_));
  AOI21_X1   g07151(.A1(new_n7208_), .A2(new_n7209_), .B(new_n7206_), .ZN(new_n7420_));
  NOR2_X1    g07152(.A1(new_n6945_), .A2(new_n7216_), .ZN(new_n7421_));
  INV_X1     g07153(.I(new_n7421_), .ZN(new_n7422_));
  OAI22_X1   g07154(.A1(new_n7218_), .A2(new_n7220_), .B1(new_n197_), .B2(new_n7422_), .ZN(new_n7423_));
  XOR2_X1    g07155(.A1(new_n7423_), .A2(new_n7420_), .Z(new_n7424_));
  INV_X1     g07156(.I(new_n7424_), .ZN(new_n7425_));
  INV_X1     g07157(.I(new_n7420_), .ZN(new_n7426_));
  NOR2_X1    g07158(.A1(new_n7423_), .A2(new_n7426_), .ZN(new_n7427_));
  INV_X1     g07159(.I(new_n7427_), .ZN(new_n7428_));
  NAND2_X1   g07160(.A1(new_n7423_), .A2(new_n7426_), .ZN(new_n7429_));
  AOI21_X1   g07161(.A1(new_n7428_), .A2(new_n7429_), .B(new_n7133_), .ZN(new_n7430_));
  AOI21_X1   g07162(.A1(new_n7425_), .A2(new_n7133_), .B(new_n7430_), .ZN(new_n7431_));
  XOR2_X1    g07163(.A1(new_n7419_), .A2(new_n7431_), .Z(new_n7432_));
  NAND2_X1   g07164(.A1(new_n7432_), .A2(new_n7409_), .ZN(new_n7433_));
  NOR2_X1    g07165(.A1(new_n7419_), .A2(new_n7431_), .ZN(new_n7434_));
  NAND2_X1   g07166(.A1(new_n7419_), .A2(new_n7431_), .ZN(new_n7435_));
  INV_X1     g07167(.I(new_n7435_), .ZN(new_n7436_));
  OAI21_X1   g07168(.A1(new_n7436_), .A2(new_n7434_), .B(new_n7408_), .ZN(new_n7437_));
  NAND2_X1   g07169(.A1(new_n7433_), .A2(new_n7437_), .ZN(new_n7438_));
  INV_X1     g07170(.I(new_n7438_), .ZN(new_n7439_));
  NOR3_X1    g07171(.A1(new_n7439_), .A2(new_n7232_), .A3(new_n7406_), .ZN(new_n7440_));
  NOR2_X1    g07172(.A1(new_n7406_), .A2(new_n7232_), .ZN(new_n7441_));
  NOR2_X1    g07173(.A1(new_n7441_), .A2(new_n7438_), .ZN(new_n7442_));
  NOR2_X1    g07174(.A1(new_n7440_), .A2(new_n7442_), .ZN(new_n7443_));
  NOR2_X1    g07175(.A1(new_n7443_), .A2(new_n7405_), .ZN(new_n7444_));
  XOR2_X1    g07176(.A1(new_n7441_), .A2(new_n7438_), .Z(new_n7445_));
  AOI21_X1   g07177(.A1(new_n7405_), .A2(new_n7445_), .B(new_n7444_), .ZN(new_n7446_));
  INV_X1     g07178(.I(new_n7446_), .ZN(new_n7447_));
  NAND2_X1   g07179(.A1(new_n7359_), .A2(new_n7340_), .ZN(new_n7448_));
  NAND2_X1   g07180(.A1(new_n7448_), .A2(new_n7361_), .ZN(new_n7449_));
  AOI21_X1   g07181(.A1(new_n7315_), .A2(new_n7318_), .B(new_n7316_), .ZN(new_n7450_));
  INV_X1     g07182(.I(new_n7450_), .ZN(new_n7451_));
  NOR2_X1    g07183(.A1(new_n4770_), .A2(new_n5175_), .ZN(new_n7452_));
  INV_X1     g07184(.I(new_n7452_), .ZN(new_n7453_));
  NOR2_X1    g07185(.A1(new_n7453_), .A2(new_n870_), .ZN(new_n7454_));
  NAND4_X1   g07186(.A1(new_n7454_), .A2(\a[11] ), .A3(new_n7073_), .A4(\a[43] ), .ZN(new_n7455_));
  AOI21_X1   g07187(.A1(new_n7455_), .A2(new_n5322_), .B(new_n786_), .ZN(new_n7456_));
  NOR3_X1    g07188(.A1(new_n870_), .A2(new_n4770_), .A3(new_n5175_), .ZN(new_n7457_));
  NOR2_X1    g07189(.A1(new_n885_), .A2(new_n6260_), .ZN(new_n7458_));
  INV_X1     g07190(.I(new_n7458_), .ZN(new_n7459_));
  NOR3_X1    g07191(.A1(new_n7459_), .A2(new_n242_), .A3(new_n4240_), .ZN(new_n7460_));
  NOR2_X1    g07192(.A1(new_n3783_), .A2(new_n6260_), .ZN(new_n7461_));
  INV_X1     g07193(.I(new_n7461_), .ZN(new_n7462_));
  NOR4_X1    g07194(.A1(new_n242_), .A2(new_n885_), .A3(new_n4240_), .A4(new_n6260_), .ZN(new_n7466_));
  INV_X1     g07195(.I(new_n7466_), .ZN(new_n7467_));
  NOR2_X1    g07196(.A1(new_n3175_), .A2(new_n2692_), .ZN(new_n7468_));
  INV_X1     g07197(.I(new_n7468_), .ZN(new_n7469_));
  NAND2_X1   g07198(.A1(\a[27] ), .A2(\a[30] ), .ZN(new_n7470_));
  NAND2_X1   g07199(.A1(new_n2689_), .A2(new_n7470_), .ZN(new_n7471_));
  NOR2_X1    g07200(.A1(new_n7469_), .A2(new_n7471_), .ZN(new_n7472_));
  NOR2_X1    g07201(.A1(new_n566_), .A2(new_n5004_), .ZN(new_n7473_));
  XNOR2_X1   g07202(.A1(new_n7472_), .A2(new_n7473_), .ZN(new_n7474_));
  NOR2_X1    g07203(.A1(new_n7474_), .A2(new_n7467_), .ZN(new_n7475_));
  INV_X1     g07204(.I(new_n7475_), .ZN(new_n7476_));
  NAND2_X1   g07205(.A1(new_n7474_), .A2(new_n7467_), .ZN(new_n7477_));
  NAND2_X1   g07206(.A1(new_n7476_), .A2(new_n7477_), .ZN(new_n7478_));
  XOR2_X1    g07207(.A1(new_n7474_), .A2(new_n7466_), .Z(new_n7479_));
  NOR2_X1    g07208(.A1(new_n7479_), .A2(new_n7457_), .ZN(new_n7480_));
  AOI21_X1   g07209(.A1(new_n7457_), .A2(new_n7478_), .B(new_n7480_), .ZN(new_n7481_));
  NOR2_X1    g07210(.A1(new_n6694_), .A2(new_n6945_), .ZN(new_n7482_));
  NOR2_X1    g07211(.A1(new_n6945_), .A2(new_n6999_), .ZN(new_n7483_));
  AOI22_X1   g07212(.A1(new_n267_), .A2(new_n7483_), .B1(new_n7482_), .B2(new_n232_), .ZN(new_n7484_));
  NOR2_X1    g07213(.A1(new_n6694_), .A2(new_n6999_), .ZN(new_n7485_));
  INV_X1     g07214(.I(new_n7485_), .ZN(new_n7486_));
  NOR2_X1    g07215(.A1(new_n200_), .A2(new_n6945_), .ZN(new_n7487_));
  NAND4_X1   g07216(.A1(new_n7484_), .A2(new_n260_), .A3(new_n7486_), .A4(new_n7487_), .ZN(new_n7488_));
  NAND2_X1   g07217(.A1(new_n1798_), .A2(new_n5600_), .ZN(new_n7489_));
  NAND2_X1   g07218(.A1(\a[5] ), .A2(\a[52] ), .ZN(new_n7490_));
  XNOR2_X1   g07219(.A1(new_n7489_), .A2(new_n7490_), .ZN(new_n7491_));
  NAND2_X1   g07220(.A1(new_n6030_), .A2(new_n597_), .ZN(new_n7492_));
  NAND2_X1   g07221(.A1(\a[15] ), .A2(\a[42] ), .ZN(new_n7493_));
  XNOR2_X1   g07222(.A1(new_n7492_), .A2(new_n7493_), .ZN(new_n7494_));
  NOR2_X1    g07223(.A1(new_n7494_), .A2(new_n7491_), .ZN(new_n7495_));
  AND2_X2    g07224(.A1(new_n7491_), .A2(new_n7494_), .Z(new_n7496_));
  NOR2_X1    g07225(.A1(new_n7496_), .A2(new_n7495_), .ZN(new_n7497_));
  XOR2_X1    g07226(.A1(new_n7494_), .A2(new_n7491_), .Z(new_n7498_));
  NAND2_X1   g07227(.A1(new_n7498_), .A2(new_n7488_), .ZN(new_n7499_));
  OAI21_X1   g07228(.A1(new_n7488_), .A2(new_n7497_), .B(new_n7499_), .ZN(new_n7500_));
  INV_X1     g07229(.I(new_n7500_), .ZN(new_n7501_));
  XOR2_X1    g07230(.A1(new_n7481_), .A2(new_n7501_), .Z(new_n7502_));
  NAND2_X1   g07231(.A1(new_n7502_), .A2(new_n7451_), .ZN(new_n7503_));
  NOR2_X1    g07232(.A1(new_n7481_), .A2(new_n7501_), .ZN(new_n7504_));
  NAND2_X1   g07233(.A1(new_n7481_), .A2(new_n7501_), .ZN(new_n7505_));
  INV_X1     g07234(.I(new_n7505_), .ZN(new_n7506_));
  OAI21_X1   g07235(.A1(new_n7506_), .A2(new_n7504_), .B(new_n7450_), .ZN(new_n7507_));
  NAND2_X1   g07236(.A1(new_n7503_), .A2(new_n7507_), .ZN(new_n7508_));
  INV_X1     g07237(.I(new_n7508_), .ZN(new_n7509_));
  NOR2_X1    g07238(.A1(new_n7344_), .A2(new_n7354_), .ZN(new_n7510_));
  NOR2_X1    g07239(.A1(new_n7510_), .A2(new_n7352_), .ZN(new_n7511_));
  INV_X1     g07240(.I(new_n6280_), .ZN(new_n7512_));
  NOR2_X1    g07241(.A1(new_n800_), .A2(new_n5745_), .ZN(new_n7513_));
  INV_X1     g07242(.I(new_n7513_), .ZN(new_n7514_));
  NOR3_X1    g07243(.A1(new_n7514_), .A2(new_n359_), .A3(new_n4414_), .ZN(new_n7515_));
  INV_X1     g07244(.I(new_n5591_), .ZN(new_n7516_));
  NOR3_X1    g07245(.A1(new_n7516_), .A2(new_n800_), .A3(new_n6055_), .ZN(new_n7517_));
  NAND2_X1   g07246(.A1(new_n7515_), .A2(new_n7517_), .ZN(new_n7518_));
  AOI21_X1   g07247(.A1(new_n7518_), .A2(new_n7512_), .B(new_n392_), .ZN(new_n7519_));
  NOR3_X1    g07248(.A1(new_n7519_), .A2(new_n268_), .A3(new_n6055_), .ZN(new_n7520_));
  INV_X1     g07249(.I(new_n7520_), .ZN(new_n7521_));
  NOR2_X1    g07250(.A1(new_n7519_), .A2(new_n7515_), .ZN(new_n7522_));
  NAND2_X1   g07251(.A1(\a[41] ), .A2(\a[49] ), .ZN(new_n7523_));
  NAND3_X1   g07252(.A1(new_n7522_), .A2(new_n7165_), .A3(new_n7523_), .ZN(new_n7524_));
  AND2_X2    g07253(.A1(new_n7524_), .A2(new_n7521_), .Z(new_n7525_));
  INV_X1     g07254(.I(new_n7525_), .ZN(new_n7526_));
  OAI22_X1   g07255(.A1(new_n1706_), .A2(new_n1773_), .B1(new_n3967_), .B2(new_n4728_), .ZN(new_n7527_));
  NAND4_X1   g07256(.A1(new_n3712_), .A2(\a[21] ), .A3(\a[36] ), .A4(new_n2285_), .ZN(new_n7528_));
  NOR2_X1    g07257(.A1(new_n7527_), .A2(new_n7528_), .ZN(new_n7529_));
  INV_X1     g07258(.I(new_n7529_), .ZN(new_n7530_));
  NAND2_X1   g07259(.A1(new_n7149_), .A2(new_n3979_), .ZN(new_n7531_));
  NAND4_X1   g07260(.A1(new_n2753_), .A2(new_n4184_), .A3(\a[24] ), .A4(\a[33] ), .ZN(new_n7532_));
  NOR2_X1    g07261(.A1(new_n7531_), .A2(new_n7532_), .ZN(new_n7533_));
  INV_X1     g07262(.I(new_n7533_), .ZN(new_n7534_));
  NOR2_X1    g07263(.A1(new_n7530_), .A2(new_n7534_), .ZN(new_n7535_));
  NOR2_X1    g07264(.A1(new_n7529_), .A2(new_n7533_), .ZN(new_n7536_));
  NOR2_X1    g07265(.A1(new_n7535_), .A2(new_n7536_), .ZN(new_n7537_));
  NOR2_X1    g07266(.A1(new_n7526_), .A2(new_n7537_), .ZN(new_n7538_));
  XNOR2_X1   g07267(.A1(new_n7529_), .A2(new_n7533_), .ZN(new_n7539_));
  NOR2_X1    g07268(.A1(new_n7525_), .A2(new_n7539_), .ZN(new_n7540_));
  NOR2_X1    g07269(.A1(new_n7538_), .A2(new_n7540_), .ZN(new_n7541_));
  NOR2_X1    g07270(.A1(new_n7189_), .A2(new_n7190_), .ZN(new_n7542_));
  NAND2_X1   g07271(.A1(new_n1532_), .A2(new_n7346_), .ZN(new_n7543_));
  INV_X1     g07272(.I(new_n7543_), .ZN(new_n7544_));
  NOR2_X1    g07273(.A1(new_n1532_), .A2(new_n7346_), .ZN(new_n7545_));
  NOR3_X1    g07274(.A1(new_n7545_), .A2(\a[21] ), .A3(\a[35] ), .ZN(new_n7546_));
  NOR2_X1    g07275(.A1(new_n7546_), .A2(new_n7544_), .ZN(new_n7547_));
  XOR2_X1    g07276(.A1(new_n7547_), .A2(new_n7542_), .Z(new_n7548_));
  NAND2_X1   g07277(.A1(new_n7548_), .A2(new_n7146_), .ZN(new_n7549_));
  NOR4_X1    g07278(.A1(new_n7546_), .A2(new_n7189_), .A3(new_n7190_), .A4(new_n7544_), .ZN(new_n7550_));
  NOR2_X1    g07279(.A1(new_n7547_), .A2(new_n7542_), .ZN(new_n7551_));
  OAI21_X1   g07280(.A1(new_n7550_), .A2(new_n7551_), .B(new_n7147_), .ZN(new_n7552_));
  NAND2_X1   g07281(.A1(new_n7549_), .A2(new_n7552_), .ZN(new_n7553_));
  INV_X1     g07282(.I(new_n7553_), .ZN(new_n7554_));
  XOR2_X1    g07283(.A1(new_n7541_), .A2(new_n7554_), .Z(new_n7555_));
  NOR2_X1    g07284(.A1(new_n7555_), .A2(new_n7511_), .ZN(new_n7556_));
  INV_X1     g07285(.I(new_n7511_), .ZN(new_n7557_));
  NOR3_X1    g07286(.A1(new_n7538_), .A2(new_n7540_), .A3(new_n7554_), .ZN(new_n7558_));
  NOR2_X1    g07287(.A1(new_n7541_), .A2(new_n7553_), .ZN(new_n7559_));
  NOR2_X1    g07288(.A1(new_n7559_), .A2(new_n7558_), .ZN(new_n7560_));
  NOR2_X1    g07289(.A1(new_n7560_), .A2(new_n7557_), .ZN(new_n7561_));
  NOR2_X1    g07290(.A1(new_n7556_), .A2(new_n7561_), .ZN(new_n7562_));
  NOR2_X1    g07291(.A1(new_n7509_), .A2(new_n7562_), .ZN(new_n7563_));
  INV_X1     g07292(.I(new_n7563_), .ZN(new_n7564_));
  NAND2_X1   g07293(.A1(new_n7509_), .A2(new_n7562_), .ZN(new_n7565_));
  NAND2_X1   g07294(.A1(new_n7564_), .A2(new_n7565_), .ZN(new_n7566_));
  XOR2_X1    g07295(.A1(new_n7508_), .A2(new_n7562_), .Z(new_n7567_));
  NOR2_X1    g07296(.A1(new_n7567_), .A2(new_n7449_), .ZN(new_n7568_));
  AOI21_X1   g07297(.A1(new_n7449_), .A2(new_n7566_), .B(new_n7568_), .ZN(new_n7569_));
  NOR2_X1    g07298(.A1(new_n7447_), .A2(new_n7569_), .ZN(new_n7570_));
  INV_X1     g07299(.I(new_n7570_), .ZN(new_n7571_));
  NAND2_X1   g07300(.A1(new_n7447_), .A2(new_n7569_), .ZN(new_n7572_));
  AOI21_X1   g07301(.A1(new_n7571_), .A2(new_n7572_), .B(new_n7392_), .ZN(new_n7573_));
  XNOR2_X1   g07302(.A1(new_n7569_), .A2(new_n7446_), .ZN(new_n7574_));
  AOI21_X1   g07303(.A1(new_n7392_), .A2(new_n7574_), .B(new_n7573_), .ZN(new_n7575_));
  OAI21_X1   g07304(.A1(new_n7236_), .A2(new_n7278_), .B(new_n7280_), .ZN(new_n7576_));
  NOR2_X1    g07305(.A1(new_n7324_), .A2(new_n7306_), .ZN(new_n7577_));
  NOR2_X1    g07306(.A1(new_n7577_), .A2(new_n7323_), .ZN(new_n7578_));
  AOI21_X1   g07307(.A1(new_n7299_), .A2(new_n7303_), .B(new_n7301_), .ZN(new_n7579_));
  INV_X1     g07308(.I(new_n7579_), .ZN(new_n7580_));
  OAI21_X1   g07309(.A1(new_n7239_), .A2(new_n7271_), .B(new_n7272_), .ZN(new_n7581_));
  NOR2_X1    g07310(.A1(new_n7292_), .A2(new_n7290_), .ZN(new_n7582_));
  NOR2_X1    g07311(.A1(new_n7582_), .A2(new_n7291_), .ZN(new_n7583_));
  INV_X1     g07312(.I(new_n7265_), .ZN(new_n7584_));
  AOI21_X1   g07313(.A1(new_n7258_), .A2(new_n7584_), .B(new_n7264_), .ZN(new_n7585_));
  NAND2_X1   g07314(.A1(new_n2500_), .A2(new_n7245_), .ZN(new_n7586_));
  NAND2_X1   g07315(.A1(\a[1] ), .A2(\a[56] ), .ZN(new_n7587_));
  NOR2_X1    g07316(.A1(new_n2499_), .A2(new_n7216_), .ZN(new_n7588_));
  AOI22_X1   g07317(.A1(new_n7588_), .A2(\a[1] ), .B1(new_n2499_), .B2(new_n7587_), .ZN(new_n7589_));
  NOR2_X1    g07318(.A1(new_n7589_), .A2(new_n7586_), .ZN(new_n7590_));
  XOR2_X1    g07319(.A1(new_n7590_), .A2(new_n199_), .Z(new_n7591_));
  XOR2_X1    g07320(.A1(new_n7591_), .A2(\a[57] ), .Z(new_n7592_));
  XNOR2_X1   g07321(.A1(new_n7585_), .A2(new_n7592_), .ZN(new_n7593_));
  NOR2_X1    g07322(.A1(new_n7593_), .A2(new_n7583_), .ZN(new_n7594_));
  INV_X1     g07323(.I(new_n7583_), .ZN(new_n7595_));
  NOR2_X1    g07324(.A1(new_n7585_), .A2(new_n7592_), .ZN(new_n7596_));
  INV_X1     g07325(.I(new_n7596_), .ZN(new_n7597_));
  NAND2_X1   g07326(.A1(new_n7585_), .A2(new_n7592_), .ZN(new_n7598_));
  AOI21_X1   g07327(.A1(new_n7597_), .A2(new_n7598_), .B(new_n7595_), .ZN(new_n7599_));
  NOR2_X1    g07328(.A1(new_n7594_), .A2(new_n7599_), .ZN(new_n7600_));
  XOR2_X1    g07329(.A1(new_n7600_), .A2(new_n7581_), .Z(new_n7601_));
  NAND2_X1   g07330(.A1(new_n7601_), .A2(new_n7580_), .ZN(new_n7602_));
  NOR2_X1    g07331(.A1(new_n7600_), .A2(new_n7581_), .ZN(new_n7603_));
  NAND2_X1   g07332(.A1(new_n7600_), .A2(new_n7581_), .ZN(new_n7604_));
  INV_X1     g07333(.I(new_n7604_), .ZN(new_n7605_));
  OAI21_X1   g07334(.A1(new_n7605_), .A2(new_n7603_), .B(new_n7579_), .ZN(new_n7606_));
  NAND2_X1   g07335(.A1(new_n7602_), .A2(new_n7606_), .ZN(new_n7607_));
  INV_X1     g07336(.I(new_n7607_), .ZN(new_n7608_));
  XOR2_X1    g07337(.A1(new_n7578_), .A2(new_n7608_), .Z(new_n7609_));
  INV_X1     g07338(.I(new_n7578_), .ZN(new_n7610_));
  NOR2_X1    g07339(.A1(new_n7610_), .A2(new_n7608_), .ZN(new_n7611_));
  NOR2_X1    g07340(.A1(new_n7578_), .A2(new_n7607_), .ZN(new_n7612_));
  NOR2_X1    g07341(.A1(new_n7611_), .A2(new_n7612_), .ZN(new_n7613_));
  MUX2_X1    g07342(.I0(new_n7613_), .I1(new_n7609_), .S(new_n7576_), .Z(new_n7614_));
  XOR2_X1    g07343(.A1(new_n7575_), .A2(new_n7614_), .Z(new_n7615_));
  NOR2_X1    g07344(.A1(new_n7615_), .A2(new_n7390_), .ZN(new_n7616_));
  INV_X1     g07345(.I(new_n7390_), .ZN(new_n7617_));
  INV_X1     g07346(.I(new_n7575_), .ZN(new_n7618_));
  NOR2_X1    g07347(.A1(new_n7618_), .A2(new_n7614_), .ZN(new_n7619_));
  INV_X1     g07348(.I(new_n7619_), .ZN(new_n7620_));
  NAND2_X1   g07349(.A1(new_n7618_), .A2(new_n7614_), .ZN(new_n7621_));
  AOI21_X1   g07350(.A1(new_n7620_), .A2(new_n7621_), .B(new_n7617_), .ZN(new_n7622_));
  NOR2_X1    g07351(.A1(new_n7622_), .A2(new_n7616_), .ZN(new_n7623_));
  XOR2_X1    g07352(.A1(new_n7623_), .A2(new_n7388_), .Z(new_n7624_));
  NAND2_X1   g07353(.A1(new_n7387_), .A2(new_n7624_), .ZN(new_n7625_));
  INV_X1     g07354(.I(new_n7388_), .ZN(new_n7626_));
  OAI21_X1   g07355(.A1(new_n7622_), .A2(new_n7616_), .B(new_n7626_), .ZN(new_n7627_));
  NAND2_X1   g07356(.A1(new_n7623_), .A2(new_n7388_), .ZN(new_n7628_));
  AND2_X2    g07357(.A1(new_n7628_), .A2(new_n7627_), .Z(new_n7629_));
  OAI21_X1   g07358(.A1(new_n7387_), .A2(new_n7629_), .B(new_n7625_), .ZN(\asquared[58] ));
  NAND2_X1   g07359(.A1(new_n7387_), .A2(new_n7627_), .ZN(new_n7631_));
  NAND2_X1   g07360(.A1(new_n7631_), .A2(new_n7628_), .ZN(new_n7632_));
  OAI21_X1   g07361(.A1(new_n7390_), .A2(new_n7619_), .B(new_n7621_), .ZN(new_n7633_));
  INV_X1     g07362(.I(new_n7611_), .ZN(new_n7634_));
  AOI21_X1   g07363(.A1(new_n7634_), .A2(new_n7576_), .B(new_n7612_), .ZN(new_n7635_));
  INV_X1     g07364(.I(new_n7394_), .ZN(new_n7636_));
  AOI21_X1   g07365(.A1(new_n7636_), .A2(new_n7403_), .B(new_n7401_), .ZN(new_n7637_));
  INV_X1     g07366(.I(new_n1029_), .ZN(new_n7638_));
  NOR2_X1    g07367(.A1(new_n4769_), .A2(new_n5745_), .ZN(new_n7639_));
  INV_X1     g07368(.I(new_n7639_), .ZN(new_n7640_));
  NOR2_X1    g07369(.A1(new_n7640_), .A2(new_n7638_), .ZN(new_n7641_));
  NOR2_X1    g07370(.A1(new_n7640_), .A2(new_n7638_), .ZN(new_n7646_));
  INV_X1     g07371(.I(\a[58] ), .ZN(new_n7647_));
  NOR2_X1    g07372(.A1(new_n7216_), .A2(new_n7647_), .ZN(new_n7648_));
  AOI22_X1   g07373(.A1(new_n7421_), .A2(new_n7648_), .B1(new_n218_), .B2(new_n4999_), .ZN(new_n7649_));
  INV_X1     g07374(.I(new_n7217_), .ZN(new_n7650_));
  NAND3_X1   g07375(.A1(new_n6946_), .A2(\a[4] ), .A3(\a[58] ), .ZN(new_n7651_));
  INV_X1     g07376(.I(new_n7651_), .ZN(new_n7652_));
  NOR2_X1    g07377(.A1(new_n6945_), .A2(new_n7647_), .ZN(new_n7653_));
  NOR4_X1    g07378(.A1(new_n7652_), .A2(new_n3123_), .A3(new_n7650_), .A4(new_n7653_), .ZN(new_n7654_));
  NAND2_X1   g07379(.A1(new_n7654_), .A2(new_n7649_), .ZN(new_n7655_));
  NAND2_X1   g07380(.A1(new_n2978_), .A2(new_n5600_), .ZN(new_n7656_));
  NAND2_X1   g07381(.A1(\a[5] ), .A2(\a[53] ), .ZN(new_n7657_));
  XNOR2_X1   g07382(.A1(new_n7656_), .A2(new_n7657_), .ZN(new_n7658_));
  NOR2_X1    g07383(.A1(new_n7655_), .A2(new_n7658_), .ZN(new_n7659_));
  INV_X1     g07384(.I(new_n7655_), .ZN(new_n7660_));
  INV_X1     g07385(.I(new_n7658_), .ZN(new_n7661_));
  NOR2_X1    g07386(.A1(new_n7660_), .A2(new_n7661_), .ZN(new_n7662_));
  OAI21_X1   g07387(.A1(new_n7662_), .A2(new_n7659_), .B(new_n7646_), .ZN(new_n7663_));
  XNOR2_X1   g07388(.A1(new_n7655_), .A2(new_n7658_), .ZN(new_n7664_));
  OAI21_X1   g07389(.A1(new_n7646_), .A2(new_n7664_), .B(new_n7663_), .ZN(new_n7665_));
  NAND2_X1   g07390(.A1(new_n6779_), .A2(new_n609_), .ZN(new_n7666_));
  NAND2_X1   g07391(.A1(\a[18] ), .A2(\a[40] ), .ZN(new_n7667_));
  XNOR2_X1   g07392(.A1(new_n7666_), .A2(new_n7667_), .ZN(new_n7668_));
  INV_X1     g07393(.I(new_n7668_), .ZN(new_n7669_));
  AOI22_X1   g07394(.A1(new_n2383_), .A2(new_n3966_), .B1(new_n4727_), .B2(new_n2286_), .ZN(new_n7670_));
  NOR2_X1    g07395(.A1(new_n1674_), .A2(new_n3393_), .ZN(new_n7671_));
  NAND4_X1   g07396(.A1(new_n7670_), .A2(new_n1956_), .A3(new_n3712_), .A4(new_n7671_), .ZN(new_n7672_));
  AOI22_X1   g07397(.A1(new_n2752_), .A2(new_n2869_), .B1(new_n2890_), .B2(new_n3851_), .ZN(new_n7673_));
  NOR2_X1    g07398(.A1(new_n2534_), .A2(new_n4184_), .ZN(new_n7674_));
  INV_X1     g07399(.I(new_n7674_), .ZN(new_n7675_));
  OAI21_X1   g07400(.A1(new_n2098_), .A2(new_n2655_), .B(new_n3500_), .ZN(new_n7676_));
  NAND4_X1   g07401(.A1(new_n7675_), .A2(new_n3474_), .A3(new_n7673_), .A4(new_n7676_), .ZN(new_n7677_));
  NOR2_X1    g07402(.A1(new_n7677_), .A2(new_n7672_), .ZN(new_n7678_));
  AND2_X2    g07403(.A1(new_n7677_), .A2(new_n7672_), .Z(new_n7679_));
  OAI21_X1   g07404(.A1(new_n7679_), .A2(new_n7678_), .B(new_n7669_), .ZN(new_n7680_));
  XNOR2_X1   g07405(.A1(new_n7677_), .A2(new_n7672_), .ZN(new_n7681_));
  OAI21_X1   g07406(.A1(new_n7669_), .A2(new_n7681_), .B(new_n7680_), .ZN(new_n7682_));
  XNOR2_X1   g07407(.A1(new_n7665_), .A2(new_n7682_), .ZN(new_n7683_));
  NOR2_X1    g07408(.A1(new_n7637_), .A2(new_n7683_), .ZN(new_n7684_));
  INV_X1     g07409(.I(new_n7637_), .ZN(new_n7685_));
  NAND2_X1   g07410(.A1(new_n7665_), .A2(new_n7682_), .ZN(new_n7686_));
  NOR2_X1    g07411(.A1(new_n7665_), .A2(new_n7682_), .ZN(new_n7687_));
  INV_X1     g07412(.I(new_n7687_), .ZN(new_n7688_));
  AOI21_X1   g07413(.A1(new_n7686_), .A2(new_n7688_), .B(new_n7685_), .ZN(new_n7689_));
  NOR2_X1    g07414(.A1(new_n7689_), .A2(new_n7684_), .ZN(new_n7690_));
  OAI21_X1   g07415(.A1(new_n7579_), .A2(new_n7603_), .B(new_n7604_), .ZN(new_n7691_));
  AOI21_X1   g07416(.A1(new_n7595_), .A2(new_n7598_), .B(new_n7596_), .ZN(new_n7692_));
  INV_X1     g07417(.I(new_n6030_), .ZN(new_n7693_));
  NOR3_X1    g07418(.A1(new_n868_), .A2(new_n4501_), .A3(new_n5511_), .ZN(new_n7694_));
  NOR3_X1    g07419(.A1(new_n7163_), .A2(new_n461_), .A3(new_n4501_), .ZN(new_n7695_));
  NAND2_X1   g07420(.A1(new_n7694_), .A2(new_n7695_), .ZN(new_n7696_));
  AOI21_X1   g07421(.A1(new_n7696_), .A2(new_n7693_), .B(new_n796_), .ZN(new_n7697_));
  NOR3_X1    g07422(.A1(new_n7697_), .A2(new_n461_), .A3(new_n5750_), .ZN(new_n7698_));
  NOR2_X1    g07423(.A1(new_n675_), .A2(new_n5511_), .ZN(new_n7699_));
  INV_X1     g07424(.I(new_n7699_), .ZN(new_n7700_));
  NOR2_X1    g07425(.A1(new_n7697_), .A2(new_n7694_), .ZN(new_n7701_));
  INV_X1     g07426(.I(new_n7701_), .ZN(new_n7702_));
  AOI21_X1   g07427(.A1(new_n5323_), .A2(new_n7700_), .B(new_n7702_), .ZN(new_n7703_));
  NOR2_X1    g07428(.A1(new_n653_), .A2(new_n786_), .ZN(new_n7704_));
  AOI21_X1   g07429(.A1(new_n5742_), .A2(new_n7452_), .B(new_n7704_), .ZN(new_n7705_));
  INV_X1     g07430(.I(new_n7705_), .ZN(new_n7706_));
  NOR4_X1    g07431(.A1(new_n7706_), .A2(new_n1220_), .A3(new_n5488_), .A4(new_n6615_), .ZN(new_n7707_));
  INV_X1     g07432(.I(new_n7707_), .ZN(new_n7708_));
  NOR2_X1    g07433(.A1(new_n242_), .A2(new_n6692_), .ZN(new_n7709_));
  INV_X1     g07434(.I(new_n7709_), .ZN(new_n7710_));
  NOR2_X1    g07435(.A1(new_n1339_), .A2(new_n3783_), .ZN(new_n7711_));
  INV_X1     g07436(.I(new_n7711_), .ZN(new_n7712_));
  NOR2_X1    g07437(.A1(new_n7710_), .A2(new_n7712_), .ZN(new_n7713_));
  XOR2_X1    g07438(.A1(new_n7713_), .A2(new_n200_), .Z(new_n7714_));
  XOR2_X1    g07439(.A1(new_n7714_), .A2(\a[55] ), .Z(new_n7715_));
  NOR2_X1    g07440(.A1(new_n7715_), .A2(new_n7708_), .ZN(new_n7716_));
  AND2_X2    g07441(.A1(new_n7715_), .A2(new_n7708_), .Z(new_n7717_));
  NOR2_X1    g07442(.A1(new_n7717_), .A2(new_n7716_), .ZN(new_n7718_));
  NOR3_X1    g07443(.A1(new_n7718_), .A2(new_n7698_), .A3(new_n7703_), .ZN(new_n7719_));
  NOR2_X1    g07444(.A1(new_n7703_), .A2(new_n7698_), .ZN(new_n7720_));
  XOR2_X1    g07445(.A1(new_n7715_), .A2(new_n7707_), .Z(new_n7721_));
  NOR2_X1    g07446(.A1(new_n7721_), .A2(new_n7720_), .ZN(new_n7722_));
  NOR2_X1    g07447(.A1(new_n7719_), .A2(new_n7722_), .ZN(new_n7723_));
  NOR2_X1    g07448(.A1(new_n242_), .A2(new_n1276_), .ZN(new_n7724_));
  AOI21_X1   g07449(.A1(new_n1441_), .A2(new_n6024_), .B(new_n7460_), .ZN(new_n7725_));
  NAND2_X1   g07450(.A1(new_n7589_), .A2(new_n7586_), .ZN(new_n7726_));
  INV_X1     g07451(.I(\a[57] ), .ZN(new_n7727_));
  NOR2_X1    g07452(.A1(new_n199_), .A2(new_n7727_), .ZN(new_n7728_));
  AOI21_X1   g07453(.A1(new_n7726_), .A2(new_n7728_), .B(new_n7590_), .ZN(new_n7729_));
  XOR2_X1    g07454(.A1(new_n7729_), .A2(new_n7725_), .Z(new_n7730_));
  INV_X1     g07455(.I(new_n7730_), .ZN(new_n7731_));
  INV_X1     g07456(.I(new_n7725_), .ZN(new_n7732_));
  NOR2_X1    g07457(.A1(new_n7732_), .A2(new_n7729_), .ZN(new_n7733_));
  INV_X1     g07458(.I(new_n7733_), .ZN(new_n7734_));
  NAND2_X1   g07459(.A1(new_n7732_), .A2(new_n7729_), .ZN(new_n7735_));
  AOI21_X1   g07460(.A1(new_n7734_), .A2(new_n7735_), .B(new_n7522_), .ZN(new_n7736_));
  AOI21_X1   g07461(.A1(new_n7731_), .A2(new_n7522_), .B(new_n7736_), .ZN(new_n7737_));
  XOR2_X1    g07462(.A1(new_n7723_), .A2(new_n7737_), .Z(new_n7738_));
  NOR2_X1    g07463(.A1(new_n7738_), .A2(new_n7692_), .ZN(new_n7739_));
  INV_X1     g07464(.I(new_n7723_), .ZN(new_n7740_));
  NOR2_X1    g07465(.A1(new_n7740_), .A2(new_n7737_), .ZN(new_n7741_));
  INV_X1     g07466(.I(new_n7741_), .ZN(new_n7742_));
  NAND2_X1   g07467(.A1(new_n7740_), .A2(new_n7737_), .ZN(new_n7743_));
  NAND2_X1   g07468(.A1(new_n7742_), .A2(new_n7743_), .ZN(new_n7744_));
  AOI21_X1   g07469(.A1(new_n7692_), .A2(new_n7744_), .B(new_n7739_), .ZN(new_n7745_));
  XNOR2_X1   g07470(.A1(new_n7745_), .A2(new_n7691_), .ZN(new_n7746_));
  NOR2_X1    g07471(.A1(new_n7746_), .A2(new_n7690_), .ZN(new_n7747_));
  INV_X1     g07472(.I(new_n7690_), .ZN(new_n7748_));
  NOR2_X1    g07473(.A1(new_n7745_), .A2(new_n7691_), .ZN(new_n7749_));
  INV_X1     g07474(.I(new_n7749_), .ZN(new_n7750_));
  NAND2_X1   g07475(.A1(new_n7745_), .A2(new_n7691_), .ZN(new_n7751_));
  AOI21_X1   g07476(.A1(new_n7750_), .A2(new_n7751_), .B(new_n7748_), .ZN(new_n7752_));
  NOR2_X1    g07477(.A1(new_n7747_), .A2(new_n7752_), .ZN(new_n7753_));
  INV_X1     g07478(.I(new_n7753_), .ZN(new_n7754_));
  AOI21_X1   g07479(.A1(new_n7451_), .A2(new_n7505_), .B(new_n7504_), .ZN(new_n7755_));
  INV_X1     g07480(.I(new_n7536_), .ZN(new_n7756_));
  AOI21_X1   g07481(.A1(new_n7525_), .A2(new_n7756_), .B(new_n7535_), .ZN(new_n7757_));
  INV_X1     g07482(.I(new_n7757_), .ZN(new_n7758_));
  NOR2_X1    g07483(.A1(new_n7456_), .A2(new_n7454_), .ZN(new_n7759_));
  AOI21_X1   g07484(.A1(new_n4999_), .A2(new_n7485_), .B(new_n7484_), .ZN(new_n7760_));
  NAND2_X1   g07485(.A1(new_n1798_), .A2(new_n5600_), .ZN(new_n7761_));
  NOR2_X1    g07486(.A1(new_n1798_), .A2(new_n5600_), .ZN(new_n7762_));
  NOR2_X1    g07487(.A1(\a[5] ), .A2(\a[52] ), .ZN(new_n7763_));
  AOI21_X1   g07488(.A1(new_n7761_), .A2(new_n7763_), .B(new_n7762_), .ZN(new_n7764_));
  XOR2_X1    g07489(.A1(new_n7760_), .A2(new_n7764_), .Z(new_n7765_));
  NAND2_X1   g07490(.A1(new_n7765_), .A2(new_n7759_), .ZN(new_n7766_));
  INV_X1     g07491(.I(new_n7759_), .ZN(new_n7767_));
  AND2_X2    g07492(.A1(new_n7760_), .A2(new_n7764_), .Z(new_n7768_));
  NOR2_X1    g07493(.A1(new_n7760_), .A2(new_n7764_), .ZN(new_n7769_));
  OAI21_X1   g07494(.A1(new_n7768_), .A2(new_n7769_), .B(new_n7767_), .ZN(new_n7770_));
  NAND2_X1   g07495(.A1(new_n7770_), .A2(new_n7766_), .ZN(new_n7771_));
  OAI21_X1   g07496(.A1(new_n2285_), .A2(new_n3712_), .B(new_n7527_), .ZN(new_n7772_));
  OAI21_X1   g07497(.A1(new_n2753_), .A2(new_n4184_), .B(new_n7531_), .ZN(new_n7773_));
  NOR2_X1    g07498(.A1(new_n6030_), .A2(new_n597_), .ZN(new_n7774_));
  NAND2_X1   g07499(.A1(new_n875_), .A2(new_n4769_), .ZN(new_n7775_));
  AOI21_X1   g07500(.A1(new_n597_), .A2(new_n6030_), .B(new_n7775_), .ZN(new_n7776_));
  NOR2_X1    g07501(.A1(new_n7776_), .A2(new_n7774_), .ZN(new_n7777_));
  XOR2_X1    g07502(.A1(new_n7773_), .A2(new_n7777_), .Z(new_n7778_));
  NOR2_X1    g07503(.A1(new_n7778_), .A2(new_n7772_), .ZN(new_n7779_));
  INV_X1     g07504(.I(new_n7772_), .ZN(new_n7780_));
  INV_X1     g07505(.I(new_n7777_), .ZN(new_n7781_));
  NOR2_X1    g07506(.A1(new_n7773_), .A2(new_n7781_), .ZN(new_n7782_));
  INV_X1     g07507(.I(new_n7782_), .ZN(new_n7783_));
  NAND2_X1   g07508(.A1(new_n7773_), .A2(new_n7781_), .ZN(new_n7784_));
  AOI21_X1   g07509(.A1(new_n7783_), .A2(new_n7784_), .B(new_n7780_), .ZN(new_n7785_));
  NOR2_X1    g07510(.A1(new_n7779_), .A2(new_n7785_), .ZN(new_n7786_));
  XNOR2_X1   g07511(.A1(new_n7771_), .A2(new_n7786_), .ZN(new_n7787_));
  NAND2_X1   g07512(.A1(new_n7787_), .A2(new_n7758_), .ZN(new_n7788_));
  INV_X1     g07513(.I(new_n7771_), .ZN(new_n7789_));
  NOR2_X1    g07514(.A1(new_n7789_), .A2(new_n7786_), .ZN(new_n7790_));
  NAND2_X1   g07515(.A1(new_n7789_), .A2(new_n7786_), .ZN(new_n7791_));
  INV_X1     g07516(.I(new_n7791_), .ZN(new_n7792_));
  OAI21_X1   g07517(.A1(new_n7792_), .A2(new_n7790_), .B(new_n7757_), .ZN(new_n7793_));
  NAND2_X1   g07518(.A1(new_n7793_), .A2(new_n7788_), .ZN(new_n7794_));
  AOI21_X1   g07519(.A1(new_n7457_), .A2(new_n7477_), .B(new_n7475_), .ZN(new_n7795_));
  NOR2_X1    g07520(.A1(new_n7496_), .A2(new_n7488_), .ZN(new_n7796_));
  NOR2_X1    g07521(.A1(new_n7796_), .A2(new_n7495_), .ZN(new_n7797_));
  NOR2_X1    g07522(.A1(\a[12] ), .A2(\a[45] ), .ZN(new_n7798_));
  AOI21_X1   g07523(.A1(new_n7469_), .A2(new_n7798_), .B(new_n7471_), .ZN(new_n7799_));
  NOR2_X1    g07524(.A1(new_n194_), .A2(new_n7727_), .ZN(new_n7800_));
  XOR2_X1    g07525(.A1(new_n7800_), .A2(new_n3355_), .Z(new_n7801_));
  NOR2_X1    g07526(.A1(new_n2462_), .A2(new_n7216_), .ZN(new_n7802_));
  INV_X1     g07527(.I(new_n7802_), .ZN(new_n7803_));
  XOR2_X1    g07528(.A1(new_n7801_), .A2(new_n7803_), .Z(new_n7804_));
  NAND2_X1   g07529(.A1(new_n7804_), .A2(new_n7799_), .ZN(new_n7805_));
  INV_X1     g07530(.I(new_n7799_), .ZN(new_n7806_));
  NOR2_X1    g07531(.A1(new_n7801_), .A2(new_n7803_), .ZN(new_n7807_));
  NAND2_X1   g07532(.A1(new_n7801_), .A2(new_n7803_), .ZN(new_n7808_));
  INV_X1     g07533(.I(new_n7808_), .ZN(new_n7809_));
  OAI21_X1   g07534(.A1(new_n7809_), .A2(new_n7807_), .B(new_n7806_), .ZN(new_n7810_));
  NAND2_X1   g07535(.A1(new_n7805_), .A2(new_n7810_), .ZN(new_n7811_));
  XNOR2_X1   g07536(.A1(new_n7811_), .A2(new_n7797_), .ZN(new_n7812_));
  AND2_X2    g07537(.A1(new_n7811_), .A2(new_n7797_), .Z(new_n7813_));
  NOR2_X1    g07538(.A1(new_n7811_), .A2(new_n7797_), .ZN(new_n7814_));
  OAI21_X1   g07539(.A1(new_n7813_), .A2(new_n7814_), .B(new_n7795_), .ZN(new_n7815_));
  OAI21_X1   g07540(.A1(new_n7795_), .A2(new_n7812_), .B(new_n7815_), .ZN(new_n7816_));
  INV_X1     g07541(.I(new_n7816_), .ZN(new_n7817_));
  XOR2_X1    g07542(.A1(new_n7794_), .A2(new_n7817_), .Z(new_n7818_));
  NOR2_X1    g07543(.A1(new_n7818_), .A2(new_n7755_), .ZN(new_n7819_));
  INV_X1     g07544(.I(new_n7755_), .ZN(new_n7820_));
  AOI21_X1   g07545(.A1(new_n7788_), .A2(new_n7793_), .B(new_n7817_), .ZN(new_n7821_));
  NOR2_X1    g07546(.A1(new_n7794_), .A2(new_n7816_), .ZN(new_n7822_));
  NOR2_X1    g07547(.A1(new_n7821_), .A2(new_n7822_), .ZN(new_n7823_));
  NOR2_X1    g07548(.A1(new_n7823_), .A2(new_n7820_), .ZN(new_n7824_));
  NOR2_X1    g07549(.A1(new_n7819_), .A2(new_n7824_), .ZN(new_n7825_));
  NOR2_X1    g07550(.A1(new_n7754_), .A2(new_n7825_), .ZN(new_n7826_));
  INV_X1     g07551(.I(new_n7826_), .ZN(new_n7827_));
  NAND2_X1   g07552(.A1(new_n7754_), .A2(new_n7825_), .ZN(new_n7828_));
  AOI21_X1   g07553(.A1(new_n7827_), .A2(new_n7828_), .B(new_n7635_), .ZN(new_n7829_));
  INV_X1     g07554(.I(new_n7635_), .ZN(new_n7830_));
  XOR2_X1    g07555(.A1(new_n7753_), .A2(new_n7825_), .Z(new_n7831_));
  NOR2_X1    g07556(.A1(new_n7831_), .A2(new_n7830_), .ZN(new_n7832_));
  NOR2_X1    g07557(.A1(new_n7829_), .A2(new_n7832_), .ZN(new_n7833_));
  NAND2_X1   g07558(.A1(new_n7572_), .A2(new_n7391_), .ZN(new_n7834_));
  NAND2_X1   g07559(.A1(new_n7834_), .A2(new_n7571_), .ZN(new_n7835_));
  INV_X1     g07560(.I(new_n7440_), .ZN(new_n7836_));
  AOI21_X1   g07561(.A1(new_n7836_), .A2(new_n7405_), .B(new_n7442_), .ZN(new_n7837_));
  INV_X1     g07562(.I(new_n7449_), .ZN(new_n7838_));
  OAI21_X1   g07563(.A1(new_n7838_), .A2(new_n7563_), .B(new_n7565_), .ZN(new_n7839_));
  INV_X1     g07564(.I(new_n7558_), .ZN(new_n7840_));
  AOI21_X1   g07565(.A1(new_n7840_), .A2(new_n7557_), .B(new_n7559_), .ZN(new_n7841_));
  OAI21_X1   g07566(.A1(new_n7408_), .A2(new_n7434_), .B(new_n7435_), .ZN(new_n7842_));
  NOR2_X1    g07567(.A1(new_n7147_), .A2(new_n7551_), .ZN(new_n7843_));
  NOR2_X1    g07568(.A1(new_n7843_), .A2(new_n7550_), .ZN(new_n7844_));
  NAND2_X1   g07569(.A1(new_n7133_), .A2(new_n7429_), .ZN(new_n7845_));
  NAND2_X1   g07570(.A1(new_n7845_), .A2(new_n7428_), .ZN(new_n7846_));
  AOI21_X1   g07571(.A1(new_n7411_), .A2(new_n7417_), .B(new_n7415_), .ZN(new_n7847_));
  XOR2_X1    g07572(.A1(new_n7847_), .A2(new_n7846_), .Z(new_n7848_));
  NOR2_X1    g07573(.A1(new_n7848_), .A2(new_n7844_), .ZN(new_n7849_));
  INV_X1     g07574(.I(new_n7844_), .ZN(new_n7850_));
  INV_X1     g07575(.I(new_n7846_), .ZN(new_n7851_));
  NOR2_X1    g07576(.A1(new_n7847_), .A2(new_n7851_), .ZN(new_n7852_));
  INV_X1     g07577(.I(new_n7852_), .ZN(new_n7853_));
  NAND2_X1   g07578(.A1(new_n7847_), .A2(new_n7851_), .ZN(new_n7854_));
  AOI21_X1   g07579(.A1(new_n7853_), .A2(new_n7854_), .B(new_n7850_), .ZN(new_n7855_));
  NOR2_X1    g07580(.A1(new_n7849_), .A2(new_n7855_), .ZN(new_n7856_));
  XNOR2_X1   g07581(.A1(new_n7856_), .A2(new_n7842_), .ZN(new_n7857_));
  NOR2_X1    g07582(.A1(new_n7857_), .A2(new_n7841_), .ZN(new_n7858_));
  INV_X1     g07583(.I(new_n7841_), .ZN(new_n7859_));
  NOR2_X1    g07584(.A1(new_n7856_), .A2(new_n7842_), .ZN(new_n7860_));
  INV_X1     g07585(.I(new_n7860_), .ZN(new_n7861_));
  NAND2_X1   g07586(.A1(new_n7856_), .A2(new_n7842_), .ZN(new_n7862_));
  AOI21_X1   g07587(.A1(new_n7861_), .A2(new_n7862_), .B(new_n7859_), .ZN(new_n7863_));
  NOR2_X1    g07588(.A1(new_n7858_), .A2(new_n7863_), .ZN(new_n7864_));
  XNOR2_X1   g07589(.A1(new_n7839_), .A2(new_n7864_), .ZN(new_n7865_));
  NOR2_X1    g07590(.A1(new_n7839_), .A2(new_n7864_), .ZN(new_n7866_));
  NAND2_X1   g07591(.A1(new_n7839_), .A2(new_n7864_), .ZN(new_n7867_));
  INV_X1     g07592(.I(new_n7867_), .ZN(new_n7868_));
  OAI21_X1   g07593(.A1(new_n7868_), .A2(new_n7866_), .B(new_n7837_), .ZN(new_n7869_));
  OAI21_X1   g07594(.A1(new_n7837_), .A2(new_n7865_), .B(new_n7869_), .ZN(new_n7870_));
  XOR2_X1    g07595(.A1(new_n7835_), .A2(new_n7870_), .Z(new_n7871_));
  NOR2_X1    g07596(.A1(new_n7871_), .A2(new_n7833_), .ZN(new_n7872_));
  INV_X1     g07597(.I(new_n7870_), .ZN(new_n7873_));
  NOR2_X1    g07598(.A1(new_n7873_), .A2(new_n7835_), .ZN(new_n7874_));
  INV_X1     g07599(.I(new_n7874_), .ZN(new_n7875_));
  NAND2_X1   g07600(.A1(new_n7873_), .A2(new_n7835_), .ZN(new_n7876_));
  NAND2_X1   g07601(.A1(new_n7875_), .A2(new_n7876_), .ZN(new_n7877_));
  AOI21_X1   g07602(.A1(new_n7833_), .A2(new_n7877_), .B(new_n7872_), .ZN(new_n7878_));
  NOR2_X1    g07603(.A1(new_n7878_), .A2(new_n7633_), .ZN(new_n7879_));
  INV_X1     g07604(.I(new_n7879_), .ZN(new_n7880_));
  NAND2_X1   g07605(.A1(new_n7878_), .A2(new_n7633_), .ZN(new_n7881_));
  NAND2_X1   g07606(.A1(new_n7880_), .A2(new_n7881_), .ZN(new_n7882_));
  XOR2_X1    g07607(.A1(new_n7632_), .A2(new_n7882_), .Z(\asquared[59] ));
  NAND2_X1   g07608(.A1(new_n7623_), .A2(new_n7881_), .ZN(new_n7884_));
  OAI21_X1   g07609(.A1(new_n7623_), .A2(new_n7881_), .B(new_n7626_), .ZN(new_n7885_));
  NAND2_X1   g07610(.A1(new_n7885_), .A2(new_n7884_), .ZN(new_n7886_));
  AOI21_X1   g07611(.A1(new_n7386_), .A2(new_n7384_), .B(new_n7886_), .ZN(new_n7887_));
  OAI21_X1   g07612(.A1(new_n7635_), .A2(new_n7826_), .B(new_n7828_), .ZN(new_n7888_));
  INV_X1     g07613(.I(new_n7888_), .ZN(new_n7889_));
  OAI21_X1   g07614(.A1(new_n7748_), .A2(new_n7749_), .B(new_n7751_), .ZN(new_n7890_));
  INV_X1     g07615(.I(new_n7821_), .ZN(new_n7891_));
  AOI21_X1   g07616(.A1(new_n7891_), .A2(new_n7820_), .B(new_n7822_), .ZN(new_n7892_));
  OAI21_X1   g07617(.A1(new_n7692_), .A2(new_n7741_), .B(new_n7743_), .ZN(new_n7893_));
  INV_X1     g07618(.I(new_n7893_), .ZN(new_n7894_));
  OAI21_X1   g07619(.A1(new_n7757_), .A2(new_n7790_), .B(new_n7791_), .ZN(new_n7895_));
  AOI21_X1   g07620(.A1(new_n7522_), .A2(new_n7735_), .B(new_n7733_), .ZN(new_n7896_));
  NOR2_X1    g07621(.A1(new_n7767_), .A2(new_n7769_), .ZN(new_n7897_));
  NOR2_X1    g07622(.A1(new_n7897_), .A2(new_n7768_), .ZN(new_n7898_));
  NAND2_X1   g07623(.A1(new_n7780_), .A2(new_n7784_), .ZN(new_n7899_));
  NAND2_X1   g07624(.A1(new_n7899_), .A2(new_n7783_), .ZN(new_n7900_));
  XOR2_X1    g07625(.A1(new_n7898_), .A2(new_n7900_), .Z(new_n7901_));
  INV_X1     g07626(.I(new_n7900_), .ZN(new_n7902_));
  NOR2_X1    g07627(.A1(new_n7898_), .A2(new_n7902_), .ZN(new_n7903_));
  NAND2_X1   g07628(.A1(new_n7898_), .A2(new_n7902_), .ZN(new_n7904_));
  INV_X1     g07629(.I(new_n7904_), .ZN(new_n7905_));
  OAI21_X1   g07630(.A1(new_n7905_), .A2(new_n7903_), .B(new_n7896_), .ZN(new_n7906_));
  OAI21_X1   g07631(.A1(new_n7896_), .A2(new_n7901_), .B(new_n7906_), .ZN(new_n7907_));
  XOR2_X1    g07632(.A1(new_n7907_), .A2(new_n7895_), .Z(new_n7908_));
  NOR2_X1    g07633(.A1(new_n7894_), .A2(new_n7908_), .ZN(new_n7909_));
  INV_X1     g07634(.I(new_n7907_), .ZN(new_n7910_));
  NOR2_X1    g07635(.A1(new_n7910_), .A2(new_n7895_), .ZN(new_n7911_));
  INV_X1     g07636(.I(new_n7911_), .ZN(new_n7912_));
  NAND2_X1   g07637(.A1(new_n7910_), .A2(new_n7895_), .ZN(new_n7913_));
  AOI21_X1   g07638(.A1(new_n7912_), .A2(new_n7913_), .B(new_n7893_), .ZN(new_n7914_));
  NOR2_X1    g07639(.A1(new_n7909_), .A2(new_n7914_), .ZN(new_n7915_));
  XOR2_X1    g07640(.A1(new_n7915_), .A2(new_n7892_), .Z(new_n7916_));
  INV_X1     g07641(.I(new_n7916_), .ZN(new_n7917_));
  INV_X1     g07642(.I(new_n7892_), .ZN(new_n7918_));
  NOR2_X1    g07643(.A1(new_n7915_), .A2(new_n7918_), .ZN(new_n7919_));
  INV_X1     g07644(.I(new_n7919_), .ZN(new_n7920_));
  NAND2_X1   g07645(.A1(new_n7915_), .A2(new_n7918_), .ZN(new_n7921_));
  AOI21_X1   g07646(.A1(new_n7920_), .A2(new_n7921_), .B(new_n7890_), .ZN(new_n7922_));
  AOI21_X1   g07647(.A1(new_n7917_), .A2(new_n7890_), .B(new_n7922_), .ZN(new_n7923_));
  OAI21_X1   g07648(.A1(new_n7837_), .A2(new_n7866_), .B(new_n7867_), .ZN(new_n7924_));
  INV_X1     g07649(.I(new_n7924_), .ZN(new_n7925_));
  OAI21_X1   g07650(.A1(new_n7637_), .A2(new_n7687_), .B(new_n7686_), .ZN(new_n7926_));
  INV_X1     g07651(.I(new_n7926_), .ZN(new_n7927_));
  INV_X1     g07652(.I(new_n7717_), .ZN(new_n7928_));
  AOI21_X1   g07653(.A1(new_n7928_), .A2(new_n7720_), .B(new_n7716_), .ZN(new_n7929_));
  INV_X1     g07654(.I(new_n7659_), .ZN(new_n7930_));
  OAI21_X1   g07655(.A1(new_n7660_), .A2(new_n7661_), .B(new_n7646_), .ZN(new_n7931_));
  NAND2_X1   g07656(.A1(new_n7931_), .A2(new_n7930_), .ZN(new_n7932_));
  NOR2_X1    g07657(.A1(new_n7679_), .A2(new_n7668_), .ZN(new_n7933_));
  NOR2_X1    g07658(.A1(new_n7933_), .A2(new_n7678_), .ZN(new_n7934_));
  XOR2_X1    g07659(.A1(new_n7934_), .A2(new_n7932_), .Z(new_n7935_));
  NOR2_X1    g07660(.A1(new_n7929_), .A2(new_n7935_), .ZN(new_n7936_));
  INV_X1     g07661(.I(new_n7932_), .ZN(new_n7937_));
  NOR2_X1    g07662(.A1(new_n7937_), .A2(new_n7934_), .ZN(new_n7938_));
  INV_X1     g07663(.I(new_n7938_), .ZN(new_n7939_));
  NAND2_X1   g07664(.A1(new_n7937_), .A2(new_n7934_), .ZN(new_n7940_));
  NAND2_X1   g07665(.A1(new_n7939_), .A2(new_n7940_), .ZN(new_n7941_));
  AOI21_X1   g07666(.A1(new_n7929_), .A2(new_n7941_), .B(new_n7936_), .ZN(new_n7942_));
  AOI21_X1   g07667(.A1(new_n1275_), .A2(new_n5350_), .B(new_n7641_), .ZN(new_n7943_));
  INV_X1     g07668(.I(new_n7943_), .ZN(new_n7944_));
  NOR2_X1    g07669(.A1(new_n7652_), .A2(new_n7649_), .ZN(new_n7945_));
  NOR2_X1    g07670(.A1(new_n200_), .A2(new_n6999_), .ZN(new_n7946_));
  OAI21_X1   g07671(.A1(new_n7709_), .A2(new_n7711_), .B(new_n7946_), .ZN(new_n7947_));
  OAI21_X1   g07672(.A1(new_n7710_), .A2(new_n7712_), .B(new_n7947_), .ZN(new_n7948_));
  XNOR2_X1   g07673(.A1(new_n7945_), .A2(new_n7948_), .ZN(new_n7949_));
  NOR2_X1    g07674(.A1(new_n7949_), .A2(new_n7944_), .ZN(new_n7950_));
  INV_X1     g07675(.I(new_n7945_), .ZN(new_n7951_));
  INV_X1     g07676(.I(new_n7948_), .ZN(new_n7952_));
  NOR2_X1    g07677(.A1(new_n7951_), .A2(new_n7952_), .ZN(new_n7953_));
  NOR2_X1    g07678(.A1(new_n7945_), .A2(new_n7948_), .ZN(new_n7954_));
  NOR2_X1    g07679(.A1(new_n7953_), .A2(new_n7954_), .ZN(new_n7955_));
  NOR2_X1    g07680(.A1(new_n7955_), .A2(new_n7943_), .ZN(new_n7956_));
  NOR2_X1    g07681(.A1(new_n7956_), .A2(new_n7950_), .ZN(new_n7957_));
  INV_X1     g07682(.I(new_n7957_), .ZN(new_n7958_));
  AOI21_X1   g07683(.A1(new_n1220_), .A2(new_n5488_), .B(new_n7705_), .ZN(new_n7959_));
  NAND2_X1   g07684(.A1(\a[1] ), .A2(\a[58] ), .ZN(new_n7960_));
  XOR2_X1    g07685(.A1(new_n7960_), .A2(\a[30] ), .Z(new_n7961_));
  XNOR2_X1   g07686(.A1(new_n7959_), .A2(new_n7961_), .ZN(new_n7962_));
  NOR2_X1    g07687(.A1(new_n7962_), .A2(new_n7702_), .ZN(new_n7963_));
  NOR2_X1    g07688(.A1(new_n7959_), .A2(new_n7961_), .ZN(new_n7964_));
  INV_X1     g07689(.I(new_n7964_), .ZN(new_n7965_));
  NAND2_X1   g07690(.A1(new_n7959_), .A2(new_n7961_), .ZN(new_n7966_));
  AOI21_X1   g07691(.A1(new_n7965_), .A2(new_n7966_), .B(new_n7701_), .ZN(new_n7967_));
  NOR2_X1    g07692(.A1(new_n7963_), .A2(new_n7967_), .ZN(new_n7968_));
  NAND2_X1   g07693(.A1(new_n2978_), .A2(new_n5600_), .ZN(new_n7969_));
  NOR2_X1    g07694(.A1(new_n2978_), .A2(new_n5600_), .ZN(new_n7970_));
  NOR2_X1    g07695(.A1(\a[5] ), .A2(\a[53] ), .ZN(new_n7971_));
  AOI21_X1   g07696(.A1(new_n7969_), .A2(new_n7971_), .B(new_n7970_), .ZN(new_n7972_));
  INV_X1     g07697(.I(new_n7972_), .ZN(new_n7973_));
  NAND2_X1   g07698(.A1(new_n6779_), .A2(new_n609_), .ZN(new_n7974_));
  NOR2_X1    g07699(.A1(new_n6779_), .A2(new_n609_), .ZN(new_n7975_));
  NOR2_X1    g07700(.A1(\a[18] ), .A2(\a[40] ), .ZN(new_n7976_));
  AOI21_X1   g07701(.A1(new_n7974_), .A2(new_n7976_), .B(new_n7975_), .ZN(new_n7977_));
  AOI21_X1   g07702(.A1(new_n2543_), .A2(new_n3487_), .B(new_n7670_), .ZN(new_n7978_));
  XNOR2_X1   g07703(.A1(new_n7978_), .A2(new_n7977_), .ZN(new_n7979_));
  NOR2_X1    g07704(.A1(new_n7979_), .A2(new_n7973_), .ZN(new_n7980_));
  INV_X1     g07705(.I(new_n7977_), .ZN(new_n7981_));
  INV_X1     g07706(.I(new_n7978_), .ZN(new_n7982_));
  NOR2_X1    g07707(.A1(new_n7982_), .A2(new_n7981_), .ZN(new_n7983_));
  NOR2_X1    g07708(.A1(new_n7978_), .A2(new_n7977_), .ZN(new_n7984_));
  NOR2_X1    g07709(.A1(new_n7983_), .A2(new_n7984_), .ZN(new_n7985_));
  NOR2_X1    g07710(.A1(new_n7985_), .A2(new_n7972_), .ZN(new_n7986_));
  NOR2_X1    g07711(.A1(new_n7986_), .A2(new_n7980_), .ZN(new_n7987_));
  NOR2_X1    g07712(.A1(new_n7987_), .A2(new_n7968_), .ZN(new_n7988_));
  NOR4_X1    g07713(.A1(new_n7986_), .A2(new_n7980_), .A3(new_n7963_), .A4(new_n7967_), .ZN(new_n7989_));
  OAI21_X1   g07714(.A1(new_n7988_), .A2(new_n7989_), .B(new_n7958_), .ZN(new_n7990_));
  XOR2_X1    g07715(.A1(new_n7987_), .A2(new_n7968_), .Z(new_n7991_));
  NAND2_X1   g07716(.A1(new_n7991_), .A2(new_n7957_), .ZN(new_n7992_));
  NAND2_X1   g07717(.A1(new_n7992_), .A2(new_n7990_), .ZN(new_n7993_));
  XOR2_X1    g07718(.A1(new_n7942_), .A2(new_n7993_), .Z(new_n7994_));
  INV_X1     g07719(.I(new_n7993_), .ZN(new_n7995_));
  NOR2_X1    g07720(.A1(new_n7995_), .A2(new_n7942_), .ZN(new_n7996_));
  NAND2_X1   g07721(.A1(new_n7995_), .A2(new_n7942_), .ZN(new_n7997_));
  INV_X1     g07722(.I(new_n7997_), .ZN(new_n7998_));
  OAI21_X1   g07723(.A1(new_n7996_), .A2(new_n7998_), .B(new_n7927_), .ZN(new_n7999_));
  OAI21_X1   g07724(.A1(new_n7927_), .A2(new_n7994_), .B(new_n7999_), .ZN(new_n8000_));
  OAI21_X1   g07725(.A1(new_n7841_), .A2(new_n7860_), .B(new_n7862_), .ZN(new_n8001_));
  INV_X1     g07726(.I(new_n8001_), .ZN(new_n8002_));
  NOR2_X1    g07727(.A1(new_n7813_), .A2(new_n7795_), .ZN(new_n8003_));
  NOR2_X1    g07728(.A1(new_n8003_), .A2(new_n7814_), .ZN(new_n8004_));
  INV_X1     g07729(.I(new_n7483_), .ZN(new_n8005_));
  NOR2_X1    g07730(.A1(new_n4240_), .A2(new_n6945_), .ZN(new_n8006_));
  INV_X1     g07731(.I(new_n8006_), .ZN(new_n8007_));
  NOR3_X1    g07732(.A1(new_n8007_), .A2(new_n353_), .A3(new_n1339_), .ZN(new_n8008_));
  NOR3_X1    g07733(.A1(new_n4718_), .A2(new_n1339_), .A3(new_n6999_), .ZN(new_n8009_));
  NAND2_X1   g07734(.A1(new_n8008_), .A2(new_n8009_), .ZN(new_n8010_));
  AOI21_X1   g07735(.A1(new_n8010_), .A2(new_n8005_), .B(new_n211_), .ZN(new_n8011_));
  NOR3_X1    g07736(.A1(new_n8011_), .A2(new_n282_), .A3(new_n6999_), .ZN(new_n8012_));
  NOR2_X1    g07737(.A1(new_n353_), .A2(new_n1339_), .ZN(new_n8013_));
  NOR3_X1    g07738(.A1(new_n8011_), .A2(new_n8013_), .A3(new_n8006_), .ZN(new_n8014_));
  NOR2_X1    g07739(.A1(new_n8012_), .A2(new_n8014_), .ZN(new_n8015_));
  INV_X1     g07740(.I(new_n8015_), .ZN(new_n8016_));
  NOR2_X1    g07741(.A1(new_n7674_), .A2(new_n7673_), .ZN(new_n8017_));
  NAND2_X1   g07742(.A1(\a[56] ), .A2(\a[57] ), .ZN(new_n8018_));
  XNOR2_X1   g07743(.A1(new_n225_), .A2(new_n8018_), .ZN(new_n8019_));
  XOR2_X1    g07744(.A1(new_n8017_), .A2(new_n8019_), .Z(new_n8020_));
  NOR3_X1    g07745(.A1(new_n8019_), .A2(new_n7673_), .A3(new_n7674_), .ZN(new_n8021_));
  INV_X1     g07746(.I(new_n8019_), .ZN(new_n8022_));
  NOR2_X1    g07747(.A1(new_n8017_), .A2(new_n8022_), .ZN(new_n8023_));
  OAI21_X1   g07748(.A1(new_n8021_), .A2(new_n8023_), .B(new_n8016_), .ZN(new_n8024_));
  OAI21_X1   g07749(.A1(new_n8016_), .A2(new_n8020_), .B(new_n8024_), .ZN(new_n8025_));
  INV_X1     g07750(.I(new_n5512_), .ZN(new_n8026_));
  NOR3_X1    g07751(.A1(new_n1812_), .A2(new_n5004_), .A3(new_n5750_), .ZN(new_n8027_));
  NAND3_X1   g07752(.A1(new_n8027_), .A2(new_n654_), .A3(new_n5512_), .ZN(new_n8028_));
  AOI21_X1   g07753(.A1(new_n8028_), .A2(new_n7693_), .B(new_n651_), .ZN(new_n8029_));
  NOR2_X1    g07754(.A1(new_n8026_), .A2(new_n653_), .ZN(new_n8031_));
  NAND2_X1   g07755(.A1(new_n5173_), .A2(new_n1275_), .ZN(new_n8032_));
  NAND2_X1   g07756(.A1(\a[8] ), .A2(\a[51] ), .ZN(new_n8033_));
  XNOR2_X1   g07757(.A1(new_n8032_), .A2(new_n8033_), .ZN(new_n8034_));
  NOR2_X1    g07758(.A1(new_n599_), .A2(new_n5175_), .ZN(new_n8035_));
  INV_X1     g07759(.I(new_n8035_), .ZN(new_n8036_));
  NOR2_X1    g07760(.A1(new_n8036_), .A2(new_n3175_), .ZN(new_n8037_));
  XOR2_X1    g07761(.A1(new_n8037_), .A2(new_n2178_), .Z(new_n8038_));
  XOR2_X1    g07762(.A1(new_n8038_), .A2(\a[31] ), .Z(new_n8039_));
  NOR2_X1    g07763(.A1(new_n8039_), .A2(new_n8034_), .ZN(new_n8040_));
  AND2_X2    g07764(.A1(new_n8039_), .A2(new_n8034_), .Z(new_n8041_));
  OAI21_X1   g07765(.A1(new_n8041_), .A2(new_n8040_), .B(new_n8031_), .ZN(new_n8042_));
  INV_X1     g07766(.I(new_n8031_), .ZN(new_n8043_));
  XOR2_X1    g07767(.A1(new_n8039_), .A2(new_n8034_), .Z(new_n8044_));
  NAND2_X1   g07768(.A1(new_n8044_), .A2(new_n8043_), .ZN(new_n8045_));
  NAND2_X1   g07769(.A1(new_n8045_), .A2(new_n8042_), .ZN(new_n8046_));
  XOR2_X1    g07770(.A1(new_n8046_), .A2(new_n8025_), .Z(new_n8047_));
  NOR2_X1    g07771(.A1(new_n8047_), .A2(new_n8004_), .ZN(new_n8048_));
  INV_X1     g07772(.I(new_n8004_), .ZN(new_n8049_));
  INV_X1     g07773(.I(new_n8046_), .ZN(new_n8050_));
  NOR2_X1    g07774(.A1(new_n8050_), .A2(new_n8025_), .ZN(new_n8051_));
  INV_X1     g07775(.I(new_n8051_), .ZN(new_n8052_));
  NAND2_X1   g07776(.A1(new_n8050_), .A2(new_n8025_), .ZN(new_n8053_));
  AOI21_X1   g07777(.A1(new_n8052_), .A2(new_n8053_), .B(new_n8049_), .ZN(new_n8054_));
  NOR2_X1    g07778(.A1(new_n8054_), .A2(new_n8048_), .ZN(new_n8055_));
  INV_X1     g07779(.I(new_n7204_), .ZN(new_n8056_));
  NOR2_X1    g07780(.A1(new_n1276_), .A2(new_n6692_), .ZN(new_n8057_));
  INV_X1     g07781(.I(new_n8057_), .ZN(new_n8058_));
  NOR2_X1    g07782(.A1(new_n7516_), .A2(new_n8058_), .ZN(new_n8059_));
  NAND4_X1   g07783(.A1(new_n8059_), .A2(\a[41] ), .A3(\a[53] ), .A4(new_n7724_), .ZN(new_n8060_));
  AOI21_X1   g07784(.A1(new_n8060_), .A2(new_n8056_), .B(new_n478_), .ZN(new_n8061_));
  NAND2_X1   g07785(.A1(\a[6] ), .A2(\a[53] ), .ZN(new_n8062_));
  NOR2_X1    g07786(.A1(new_n8061_), .A2(new_n8059_), .ZN(new_n8063_));
  INV_X1     g07787(.I(new_n8063_), .ZN(new_n8064_));
  OAI21_X1   g07788(.A1(new_n4414_), .A2(new_n6692_), .B(new_n1004_), .ZN(new_n8065_));
  OAI22_X1   g07789(.A1(new_n8064_), .A2(new_n8065_), .B1(new_n8061_), .B2(new_n8062_), .ZN(new_n8066_));
  NOR3_X1    g07790(.A1(new_n1785_), .A2(new_n4770_), .A3(new_n5745_), .ZN(new_n8067_));
  NOR4_X1    g07791(.A1(new_n364_), .A2(new_n875_), .A3(new_n4770_), .A4(new_n6055_), .ZN(new_n8068_));
  NAND2_X1   g07792(.A1(new_n8068_), .A2(new_n8067_), .ZN(new_n8069_));
  AOI21_X1   g07793(.A1(new_n8069_), .A2(new_n7512_), .B(new_n525_), .ZN(new_n8070_));
  NOR3_X1    g07794(.A1(new_n8070_), .A2(new_n364_), .A3(new_n6055_), .ZN(new_n8071_));
  NOR2_X1    g07795(.A1(new_n4770_), .A2(new_n5745_), .ZN(new_n8072_));
  NOR3_X1    g07796(.A1(new_n8070_), .A2(new_n1786_), .A3(new_n8072_), .ZN(new_n8073_));
  NOR2_X1    g07797(.A1(new_n8071_), .A2(new_n8073_), .ZN(new_n8074_));
  OAI21_X1   g07798(.A1(new_n7806_), .A2(new_n7807_), .B(new_n7808_), .ZN(new_n8075_));
  XNOR2_X1   g07799(.A1(new_n8075_), .A2(new_n8074_), .ZN(new_n8076_));
  AND2_X2    g07800(.A1(new_n8075_), .A2(new_n8074_), .Z(new_n8077_));
  NOR2_X1    g07801(.A1(new_n8075_), .A2(new_n8074_), .ZN(new_n8078_));
  OAI21_X1   g07802(.A1(new_n8077_), .A2(new_n8078_), .B(new_n8066_), .ZN(new_n8079_));
  OAI21_X1   g07803(.A1(new_n8066_), .A2(new_n8076_), .B(new_n8079_), .ZN(new_n8080_));
  INV_X1     g07804(.I(new_n8080_), .ZN(new_n8081_));
  NAND2_X1   g07805(.A1(new_n7854_), .A2(new_n7850_), .ZN(new_n8082_));
  NAND2_X1   g07806(.A1(new_n8082_), .A2(new_n7853_), .ZN(new_n8083_));
  INV_X1     g07807(.I(new_n8083_), .ZN(new_n8084_));
  INV_X1     g07808(.I(\a[59] ), .ZN(new_n8085_));
  NOR2_X1    g07809(.A1(new_n2765_), .A2(new_n8085_), .ZN(new_n8086_));
  INV_X1     g07810(.I(new_n8086_), .ZN(new_n8087_));
  NOR2_X1    g07811(.A1(new_n8087_), .A2(new_n2281_), .ZN(new_n8088_));
  NAND4_X1   g07812(.A1(new_n8088_), .A2(\a[33] ), .A3(\a[59] ), .A4(new_n2057_), .ZN(new_n8089_));
  AOI21_X1   g07813(.A1(new_n8089_), .A2(new_n2534_), .B(new_n3852_), .ZN(new_n8090_));
  NOR3_X1    g07814(.A1(new_n8090_), .A2(new_n1916_), .A3(new_n2868_), .ZN(new_n8091_));
  NOR2_X1    g07815(.A1(new_n8090_), .A2(new_n8088_), .ZN(new_n8092_));
  AND3_X2    g07816(.A1(new_n8092_), .A2(new_n2281_), .A3(new_n8087_), .Z(new_n8093_));
  NOR2_X1    g07817(.A1(new_n8093_), .A2(new_n8091_), .ZN(new_n8094_));
  AOI22_X1   g07818(.A1(new_n2978_), .A2(new_n5601_), .B1(new_n5339_), .B2(new_n4437_), .ZN(new_n8095_));
  NOR4_X1    g07819(.A1(new_n4538_), .A2(new_n5600_), .A3(new_n1215_), .A4(new_n3783_), .ZN(new_n8096_));
  AND2_X2    g07820(.A1(new_n8095_), .A2(new_n8096_), .Z(new_n8097_));
  NOR2_X1    g07821(.A1(new_n4729_), .A2(new_n6700_), .ZN(new_n8098_));
  NOR4_X1    g07822(.A1(new_n3487_), .A2(new_n2277_), .A3(new_n2368_), .A4(new_n3393_), .ZN(new_n8099_));
  NAND2_X1   g07823(.A1(new_n8098_), .A2(new_n8099_), .ZN(new_n8100_));
  INV_X1     g07824(.I(new_n8100_), .ZN(new_n8101_));
  NAND2_X1   g07825(.A1(new_n8101_), .A2(new_n8097_), .ZN(new_n8102_));
  INV_X1     g07826(.I(new_n8102_), .ZN(new_n8103_));
  NOR2_X1    g07827(.A1(new_n8101_), .A2(new_n8097_), .ZN(new_n8104_));
  OAI21_X1   g07828(.A1(new_n8103_), .A2(new_n8104_), .B(new_n8094_), .ZN(new_n8105_));
  XOR2_X1    g07829(.A1(new_n8100_), .A2(new_n8097_), .Z(new_n8106_));
  OAI21_X1   g07830(.A1(new_n8094_), .A2(new_n8106_), .B(new_n8105_), .ZN(new_n8107_));
  INV_X1     g07831(.I(new_n8107_), .ZN(new_n8108_));
  NOR2_X1    g07832(.A1(new_n8084_), .A2(new_n8108_), .ZN(new_n8109_));
  NOR2_X1    g07833(.A1(new_n8083_), .A2(new_n8107_), .ZN(new_n8110_));
  NOR2_X1    g07834(.A1(new_n8109_), .A2(new_n8110_), .ZN(new_n8111_));
  NOR2_X1    g07835(.A1(new_n8111_), .A2(new_n8081_), .ZN(new_n8112_));
  XNOR2_X1   g07836(.A1(new_n8083_), .A2(new_n8107_), .ZN(new_n8113_));
  NOR2_X1    g07837(.A1(new_n8113_), .A2(new_n8080_), .ZN(new_n8114_));
  NOR2_X1    g07838(.A1(new_n8112_), .A2(new_n8114_), .ZN(new_n8115_));
  NOR2_X1    g07839(.A1(new_n8115_), .A2(new_n8055_), .ZN(new_n8116_));
  INV_X1     g07840(.I(new_n8116_), .ZN(new_n8117_));
  NAND2_X1   g07841(.A1(new_n8115_), .A2(new_n8055_), .ZN(new_n8118_));
  AOI21_X1   g07842(.A1(new_n8117_), .A2(new_n8118_), .B(new_n8002_), .ZN(new_n8119_));
  XOR2_X1    g07843(.A1(new_n8115_), .A2(new_n8055_), .Z(new_n8120_));
  AOI21_X1   g07844(.A1(new_n8002_), .A2(new_n8120_), .B(new_n8119_), .ZN(new_n8121_));
  XNOR2_X1   g07845(.A1(new_n8121_), .A2(new_n8000_), .ZN(new_n8122_));
  NOR2_X1    g07846(.A1(new_n8121_), .A2(new_n8000_), .ZN(new_n8123_));
  INV_X1     g07847(.I(new_n8123_), .ZN(new_n8124_));
  NAND2_X1   g07848(.A1(new_n8121_), .A2(new_n8000_), .ZN(new_n8125_));
  NAND2_X1   g07849(.A1(new_n8124_), .A2(new_n8125_), .ZN(new_n8126_));
  NAND2_X1   g07850(.A1(new_n8126_), .A2(new_n7925_), .ZN(new_n8127_));
  OAI21_X1   g07851(.A1(new_n7925_), .A2(new_n8122_), .B(new_n8127_), .ZN(new_n8128_));
  XOR2_X1    g07852(.A1(new_n8128_), .A2(new_n7923_), .Z(new_n8129_));
  NOR2_X1    g07853(.A1(new_n8129_), .A2(new_n7889_), .ZN(new_n8130_));
  INV_X1     g07854(.I(new_n8128_), .ZN(new_n8131_));
  NOR2_X1    g07855(.A1(new_n8131_), .A2(new_n7923_), .ZN(new_n8132_));
  INV_X1     g07856(.I(new_n8132_), .ZN(new_n8133_));
  NAND2_X1   g07857(.A1(new_n8131_), .A2(new_n7923_), .ZN(new_n8134_));
  AOI21_X1   g07858(.A1(new_n8133_), .A2(new_n8134_), .B(new_n7888_), .ZN(new_n8135_));
  NOR2_X1    g07859(.A1(new_n8135_), .A2(new_n8130_), .ZN(new_n8136_));
  OAI21_X1   g07860(.A1(new_n7833_), .A2(new_n7874_), .B(new_n7876_), .ZN(new_n8137_));
  INV_X1     g07861(.I(new_n8137_), .ZN(new_n8138_));
  NOR2_X1    g07862(.A1(new_n8136_), .A2(new_n8138_), .ZN(new_n8139_));
  XOR2_X1    g07863(.A1(new_n7887_), .A2(new_n8139_), .Z(new_n8140_));
  XOR2_X1    g07864(.A1(new_n8140_), .A2(new_n7879_), .Z(\asquared[60] ));
  NOR2_X1    g07865(.A1(new_n7880_), .A2(new_n8136_), .ZN(new_n8142_));
  AOI21_X1   g07866(.A1(new_n7880_), .A2(new_n8136_), .B(new_n8138_), .ZN(new_n8143_));
  AOI21_X1   g07867(.A1(new_n7887_), .A2(new_n8143_), .B(new_n8142_), .ZN(new_n8144_));
  INV_X1     g07868(.I(new_n7921_), .ZN(new_n8145_));
  AOI21_X1   g07869(.A1(new_n7890_), .A2(new_n7920_), .B(new_n8145_), .ZN(new_n8146_));
  OAI21_X1   g07870(.A1(new_n7894_), .A2(new_n7911_), .B(new_n7913_), .ZN(new_n8147_));
  INV_X1     g07871(.I(new_n8147_), .ZN(new_n8148_));
  NOR2_X1    g07872(.A1(new_n7988_), .A2(new_n7958_), .ZN(new_n8149_));
  NOR2_X1    g07873(.A1(new_n8149_), .A2(new_n7989_), .ZN(new_n8150_));
  OAI21_X1   g07874(.A1(new_n7702_), .A2(new_n7964_), .B(new_n7966_), .ZN(new_n8151_));
  INV_X1     g07875(.I(new_n8151_), .ZN(new_n8152_));
  NOR2_X1    g07876(.A1(new_n2625_), .A2(new_n7647_), .ZN(new_n8153_));
  INV_X1     g07877(.I(new_n8153_), .ZN(new_n8154_));
  NOR2_X1    g07878(.A1(new_n194_), .A2(new_n8085_), .ZN(new_n8155_));
  XNOR2_X1   g07879(.A1(new_n8155_), .A2(new_n3734_), .ZN(new_n8156_));
  NOR2_X1    g07880(.A1(new_n8156_), .A2(new_n8154_), .ZN(new_n8157_));
  XOR2_X1    g07881(.A1(new_n8157_), .A2(new_n199_), .Z(new_n8158_));
  XOR2_X1    g07882(.A1(new_n8158_), .A2(\a[60] ), .Z(new_n8159_));
  AOI22_X1   g07883(.A1(new_n3851_), .A2(new_n4190_), .B1(new_n7131_), .B2(new_n2797_), .ZN(new_n8160_));
  INV_X1     g07884(.I(new_n8160_), .ZN(new_n8161_));
  NOR2_X1    g07885(.A1(new_n2178_), .A2(new_n2765_), .ZN(new_n8162_));
  NOR2_X1    g07886(.A1(new_n2368_), .A2(new_n3837_), .ZN(new_n8163_));
  XNOR2_X1   g07887(.A1(new_n8162_), .A2(new_n8163_), .ZN(new_n8164_));
  INV_X1     g07888(.I(new_n8164_), .ZN(new_n8165_));
  NOR2_X1    g07889(.A1(new_n8164_), .A2(new_n8162_), .ZN(new_n8166_));
  NOR2_X1    g07890(.A1(new_n2098_), .A2(new_n2868_), .ZN(new_n8167_));
  OAI22_X1   g07891(.A1(new_n8166_), .A2(new_n8161_), .B1(new_n8165_), .B2(new_n8167_), .ZN(new_n8168_));
  XNOR2_X1   g07892(.A1(new_n8159_), .A2(new_n8168_), .ZN(new_n8169_));
  NOR2_X1    g07893(.A1(new_n8169_), .A2(new_n8152_), .ZN(new_n8170_));
  NOR2_X1    g07894(.A1(new_n8159_), .A2(new_n8168_), .ZN(new_n8171_));
  INV_X1     g07895(.I(new_n8171_), .ZN(new_n8172_));
  NAND2_X1   g07896(.A1(new_n8159_), .A2(new_n8168_), .ZN(new_n8173_));
  AOI21_X1   g07897(.A1(new_n8172_), .A2(new_n8173_), .B(new_n8151_), .ZN(new_n8174_));
  NOR2_X1    g07898(.A1(new_n8170_), .A2(new_n8174_), .ZN(new_n8175_));
  NOR2_X1    g07899(.A1(new_n4769_), .A2(new_n6694_), .ZN(new_n8177_));
  NAND2_X1   g07900(.A1(\a[7] ), .A2(\a[8] ), .ZN(new_n8178_));
  NOR2_X1    g07901(.A1(new_n8056_), .A2(new_n8178_), .ZN(new_n8179_));
  NAND2_X1   g07902(.A1(\a[7] ), .A2(\a[53] ), .ZN(new_n8180_));
  INV_X1     g07903(.I(new_n1918_), .ZN(new_n8181_));
  NOR3_X1    g07904(.A1(new_n8181_), .A2(new_n4769_), .A3(new_n6692_), .ZN(new_n8182_));
  NOR2_X1    g07905(.A1(new_n8182_), .A2(new_n8179_), .ZN(new_n8183_));
  INV_X1     g07906(.I(new_n8183_), .ZN(new_n8184_));
  OAI21_X1   g07907(.A1(new_n4769_), .A2(new_n6692_), .B(new_n8181_), .ZN(new_n8185_));
  OAI22_X1   g07908(.A1(new_n8184_), .A2(new_n8185_), .B1(new_n8179_), .B2(new_n8180_), .ZN(new_n8186_));
  NOR2_X1    g07909(.A1(new_n4414_), .A2(new_n6999_), .ZN(new_n8187_));
  AOI22_X1   g07910(.A1(new_n8013_), .A2(new_n8187_), .B1(new_n7483_), .B2(new_n608_), .ZN(new_n8188_));
  NOR2_X1    g07911(.A1(new_n242_), .A2(new_n6945_), .ZN(new_n8189_));
  INV_X1     g07912(.I(new_n8189_), .ZN(new_n8190_));
  NOR2_X1    g07913(.A1(new_n1339_), .A2(new_n4414_), .ZN(new_n8191_));
  AOI21_X1   g07914(.A1(new_n8190_), .A2(new_n8191_), .B(new_n8188_), .ZN(new_n8192_));
  INV_X1     g07915(.I(new_n8192_), .ZN(new_n8193_));
  XNOR2_X1   g07916(.A1(new_n8189_), .A2(new_n8191_), .ZN(new_n8194_));
  OAI21_X1   g07917(.A1(new_n353_), .A2(new_n6999_), .B(new_n8194_), .ZN(new_n8195_));
  AND2_X2    g07918(.A1(new_n8195_), .A2(new_n8193_), .Z(new_n8196_));
  INV_X1     g07919(.I(new_n8196_), .ZN(new_n8197_));
  NOR2_X1    g07920(.A1(new_n5175_), .A2(new_n5750_), .ZN(new_n8198_));
  INV_X1     g07921(.I(new_n8198_), .ZN(new_n8199_));
  NOR2_X1    g07922(.A1(new_n8199_), .A2(new_n5793_), .ZN(new_n8200_));
  NOR2_X1    g07923(.A1(new_n8200_), .A2(new_n7704_), .ZN(new_n8201_));
  INV_X1     g07924(.I(new_n8201_), .ZN(new_n8202_));
  NOR4_X1    g07925(.A1(new_n8202_), .A2(new_n1220_), .A3(new_n6030_), .A4(new_n7139_), .ZN(new_n8203_));
  INV_X1     g07926(.I(new_n8203_), .ZN(new_n8204_));
  NOR2_X1    g07927(.A1(new_n8197_), .A2(new_n8204_), .ZN(new_n8205_));
  NOR2_X1    g07928(.A1(new_n8196_), .A2(new_n8203_), .ZN(new_n8206_));
  NOR2_X1    g07929(.A1(new_n8205_), .A2(new_n8206_), .ZN(new_n8207_));
  NOR2_X1    g07930(.A1(new_n8207_), .A2(new_n8186_), .ZN(new_n8208_));
  INV_X1     g07931(.I(new_n8186_), .ZN(new_n8209_));
  XOR2_X1    g07932(.A1(new_n8196_), .A2(new_n8204_), .Z(new_n8210_));
  NOR2_X1    g07933(.A1(new_n8210_), .A2(new_n8209_), .ZN(new_n8211_));
  NOR2_X1    g07934(.A1(new_n8208_), .A2(new_n8211_), .ZN(new_n8212_));
  XOR2_X1    g07935(.A1(new_n8175_), .A2(new_n8212_), .Z(new_n8213_));
  NOR3_X1    g07936(.A1(new_n8170_), .A2(new_n8174_), .A3(new_n8212_), .ZN(new_n8214_));
  NOR3_X1    g07937(.A1(new_n8175_), .A2(new_n8208_), .A3(new_n8211_), .ZN(new_n8215_));
  OAI21_X1   g07938(.A1(new_n8215_), .A2(new_n8214_), .B(new_n8150_), .ZN(new_n8216_));
  OAI21_X1   g07939(.A1(new_n8213_), .A2(new_n8150_), .B(new_n8216_), .ZN(new_n8217_));
  NOR2_X1    g07940(.A1(new_n7905_), .A2(new_n7896_), .ZN(new_n8218_));
  NOR2_X1    g07941(.A1(new_n8218_), .A2(new_n7903_), .ZN(new_n8219_));
  AOI21_X1   g07942(.A1(new_n654_), .A2(new_n5512_), .B(new_n8029_), .ZN(new_n8220_));
  INV_X1     g07943(.I(new_n8220_), .ZN(new_n8221_));
  NOR3_X1    g07944(.A1(new_n7638_), .A2(new_n4770_), .A3(new_n6260_), .ZN(new_n8222_));
  NOR3_X1    g07945(.A1(new_n7638_), .A2(new_n4770_), .A3(new_n6260_), .ZN(new_n8226_));
  NOR2_X1    g07946(.A1(new_n5004_), .A2(new_n5745_), .ZN(new_n8227_));
  INV_X1     g07947(.I(new_n8227_), .ZN(new_n8228_));
  NOR2_X1    g07948(.A1(new_n8228_), .A2(new_n868_), .ZN(new_n8229_));
  NAND4_X1   g07949(.A1(new_n8229_), .A2(\a[45] ), .A3(new_n1786_), .A4(\a[50] ), .ZN(new_n8230_));
  AOI21_X1   g07950(.A1(new_n8230_), .A2(new_n7512_), .B(new_n796_), .ZN(new_n8231_));
  NOR2_X1    g07951(.A1(new_n8228_), .A2(new_n868_), .ZN(new_n8233_));
  XNOR2_X1   g07952(.A1(new_n8226_), .A2(new_n8233_), .ZN(new_n8234_));
  NOR2_X1    g07953(.A1(new_n8221_), .A2(new_n8234_), .ZN(new_n8235_));
  INV_X1     g07954(.I(new_n8226_), .ZN(new_n8236_));
  INV_X1     g07955(.I(new_n8233_), .ZN(new_n8237_));
  NOR2_X1    g07956(.A1(new_n8236_), .A2(new_n8237_), .ZN(new_n8238_));
  NOR2_X1    g07957(.A1(new_n8226_), .A2(new_n8233_), .ZN(new_n8239_));
  OR2_X2     g07958(.A1(new_n8238_), .A2(new_n8239_), .Z(new_n8240_));
  AOI21_X1   g07959(.A1(new_n8221_), .A2(new_n8240_), .B(new_n8235_), .ZN(new_n8241_));
  NOR2_X1    g07960(.A1(new_n7216_), .A2(new_n7727_), .ZN(new_n8242_));
  INV_X1     g07961(.I(new_n8242_), .ZN(new_n8243_));
  INV_X1     g07962(.I(new_n7648_), .ZN(new_n8244_));
  NOR2_X1    g07963(.A1(new_n7727_), .A2(new_n7647_), .ZN(new_n8245_));
  INV_X1     g07964(.I(new_n8245_), .ZN(new_n8246_));
  NOR2_X1    g07965(.A1(new_n8244_), .A2(new_n8246_), .ZN(new_n8247_));
  NOR2_X1    g07966(.A1(new_n8247_), .A2(new_n1271_), .ZN(new_n8248_));
  NOR2_X1    g07967(.A1(new_n201_), .A2(new_n7647_), .ZN(new_n8249_));
  NAND4_X1   g07968(.A1(new_n8248_), .A2(new_n212_), .A3(new_n8243_), .A4(new_n8249_), .ZN(new_n8250_));
  INV_X1     g07969(.I(new_n4241_), .ZN(new_n8251_));
  NOR2_X1    g07970(.A1(new_n8251_), .A2(new_n4321_), .ZN(new_n8252_));
  NOR2_X1    g07971(.A1(new_n8252_), .A2(new_n7009_), .ZN(new_n8253_));
  NOR4_X1    g07972(.A1(new_n5339_), .A2(new_n4538_), .A3(new_n1215_), .A4(new_n4240_), .ZN(new_n8254_));
  NAND2_X1   g07973(.A1(new_n8253_), .A2(new_n8254_), .ZN(new_n8255_));
  AOI22_X1   g07974(.A1(new_n2277_), .A2(new_n4727_), .B1(new_n3966_), .B2(new_n4515_), .ZN(new_n8256_));
  NOR4_X1    g07975(.A1(new_n2752_), .A2(new_n3487_), .A3(new_n1691_), .A4(new_n3393_), .ZN(new_n8257_));
  NAND2_X1   g07976(.A1(new_n8256_), .A2(new_n8257_), .ZN(new_n8258_));
  NOR2_X1    g07977(.A1(new_n8255_), .A2(new_n8258_), .ZN(new_n8259_));
  INV_X1     g07978(.I(new_n8258_), .ZN(new_n8260_));
  AOI21_X1   g07979(.A1(new_n8253_), .A2(new_n8254_), .B(new_n8260_), .ZN(new_n8261_));
  NOR2_X1    g07980(.A1(new_n8261_), .A2(new_n8259_), .ZN(new_n8262_));
  NOR2_X1    g07981(.A1(new_n8262_), .A2(new_n8250_), .ZN(new_n8263_));
  INV_X1     g07982(.I(new_n8250_), .ZN(new_n8264_));
  XOR2_X1    g07983(.A1(new_n8255_), .A2(new_n8260_), .Z(new_n8265_));
  NOR2_X1    g07984(.A1(new_n8265_), .A2(new_n8264_), .ZN(new_n8266_));
  NOR2_X1    g07985(.A1(new_n8266_), .A2(new_n8263_), .ZN(new_n8267_));
  XOR2_X1    g07986(.A1(new_n8267_), .A2(new_n8241_), .Z(new_n8268_));
  INV_X1     g07987(.I(new_n8241_), .ZN(new_n8269_));
  NOR2_X1    g07988(.A1(new_n8267_), .A2(new_n8269_), .ZN(new_n8270_));
  NAND2_X1   g07989(.A1(new_n8267_), .A2(new_n8269_), .ZN(new_n8271_));
  INV_X1     g07990(.I(new_n8271_), .ZN(new_n8272_));
  OAI21_X1   g07991(.A1(new_n8270_), .A2(new_n8272_), .B(new_n8219_), .ZN(new_n8273_));
  OAI21_X1   g07992(.A1(new_n8219_), .A2(new_n8268_), .B(new_n8273_), .ZN(new_n8274_));
  NAND2_X1   g07993(.A1(new_n8217_), .A2(new_n8274_), .ZN(new_n8275_));
  NOR2_X1    g07994(.A1(new_n8217_), .A2(new_n8274_), .ZN(new_n8276_));
  INV_X1     g07995(.I(new_n8276_), .ZN(new_n8277_));
  AOI21_X1   g07996(.A1(new_n8277_), .A2(new_n8275_), .B(new_n8148_), .ZN(new_n8278_));
  XNOR2_X1   g07997(.A1(new_n8217_), .A2(new_n8274_), .ZN(new_n8279_));
  NOR2_X1    g07998(.A1(new_n8279_), .A2(new_n8147_), .ZN(new_n8280_));
  NOR2_X1    g07999(.A1(new_n8280_), .A2(new_n8278_), .ZN(new_n8281_));
  AOI21_X1   g08000(.A1(new_n8049_), .A2(new_n8053_), .B(new_n8051_), .ZN(new_n8282_));
  INV_X1     g08001(.I(new_n8282_), .ZN(new_n8283_));
  NOR2_X1    g08002(.A1(new_n8066_), .A2(new_n8078_), .ZN(new_n8284_));
  NOR2_X1    g08003(.A1(new_n8284_), .A2(new_n8077_), .ZN(new_n8285_));
  NOR2_X1    g08004(.A1(new_n8011_), .A2(new_n8008_), .ZN(new_n8286_));
  AOI21_X1   g08005(.A1(new_n4538_), .A2(new_n5600_), .B(new_n8095_), .ZN(new_n8287_));
  AOI21_X1   g08006(.A1(new_n2277_), .A2(new_n3487_), .B(new_n8098_), .ZN(new_n8288_));
  XOR2_X1    g08007(.A1(new_n8288_), .A2(new_n8287_), .Z(new_n8289_));
  NAND2_X1   g08008(.A1(new_n8289_), .A2(new_n8286_), .ZN(new_n8290_));
  INV_X1     g08009(.I(new_n8286_), .ZN(new_n8291_));
  AND2_X2    g08010(.A1(new_n8288_), .A2(new_n8287_), .Z(new_n8292_));
  NOR2_X1    g08011(.A1(new_n8288_), .A2(new_n8287_), .ZN(new_n8293_));
  OAI21_X1   g08012(.A1(new_n8292_), .A2(new_n8293_), .B(new_n8291_), .ZN(new_n8294_));
  NAND2_X1   g08013(.A1(new_n8290_), .A2(new_n8294_), .ZN(new_n8295_));
  NOR2_X1    g08014(.A1(new_n8070_), .A2(new_n8067_), .ZN(new_n8296_));
  NOR3_X1    g08015(.A1(new_n3355_), .A2(new_n194_), .A3(new_n7727_), .ZN(new_n8297_));
  AOI21_X1   g08016(.A1(new_n8297_), .A2(new_n232_), .B(new_n8242_), .ZN(new_n8298_));
  XOR2_X1    g08017(.A1(new_n8092_), .A2(new_n8298_), .Z(new_n8299_));
  INV_X1     g08018(.I(new_n8299_), .ZN(new_n8300_));
  INV_X1     g08019(.I(new_n8092_), .ZN(new_n8301_));
  NOR2_X1    g08020(.A1(new_n8301_), .A2(new_n8298_), .ZN(new_n8302_));
  INV_X1     g08021(.I(new_n8302_), .ZN(new_n8303_));
  NAND2_X1   g08022(.A1(new_n8301_), .A2(new_n8298_), .ZN(new_n8304_));
  AOI21_X1   g08023(.A1(new_n8303_), .A2(new_n8304_), .B(new_n8296_), .ZN(new_n8305_));
  AOI21_X1   g08024(.A1(new_n8296_), .A2(new_n8300_), .B(new_n8305_), .ZN(new_n8306_));
  XOR2_X1    g08025(.A1(new_n8306_), .A2(new_n8295_), .Z(new_n8307_));
  INV_X1     g08026(.I(new_n8295_), .ZN(new_n8308_));
  NOR2_X1    g08027(.A1(new_n8306_), .A2(new_n8308_), .ZN(new_n8309_));
  NAND2_X1   g08028(.A1(new_n8306_), .A2(new_n8308_), .ZN(new_n8310_));
  INV_X1     g08029(.I(new_n8310_), .ZN(new_n8311_));
  OAI21_X1   g08030(.A1(new_n8311_), .A2(new_n8309_), .B(new_n8285_), .ZN(new_n8312_));
  OAI21_X1   g08031(.A1(new_n8285_), .A2(new_n8307_), .B(new_n8312_), .ZN(new_n8313_));
  NAND2_X1   g08032(.A1(new_n5173_), .A2(new_n1275_), .ZN(new_n8314_));
  NOR2_X1    g08033(.A1(new_n5173_), .A2(new_n1275_), .ZN(new_n8315_));
  NOR2_X1    g08034(.A1(\a[8] ), .A2(\a[51] ), .ZN(new_n8316_));
  AOI21_X1   g08035(.A1(new_n8314_), .A2(new_n8316_), .B(new_n8315_), .ZN(new_n8317_));
  NOR2_X1    g08036(.A1(new_n2178_), .A2(new_n2655_), .ZN(new_n8318_));
  OAI21_X1   g08037(.A1(new_n2898_), .A2(new_n8035_), .B(new_n8318_), .ZN(new_n8319_));
  OAI21_X1   g08038(.A1(new_n3175_), .A2(new_n8036_), .B(new_n8319_), .ZN(new_n8320_));
  XNOR2_X1   g08039(.A1(new_n8320_), .A2(new_n8317_), .ZN(new_n8321_));
  NOR2_X1    g08040(.A1(new_n8064_), .A2(new_n8321_), .ZN(new_n8322_));
  INV_X1     g08041(.I(new_n8317_), .ZN(new_n8323_));
  INV_X1     g08042(.I(new_n8320_), .ZN(new_n8324_));
  NOR2_X1    g08043(.A1(new_n8324_), .A2(new_n8323_), .ZN(new_n8325_));
  NOR2_X1    g08044(.A1(new_n8320_), .A2(new_n8317_), .ZN(new_n8326_));
  NOR2_X1    g08045(.A1(new_n8325_), .A2(new_n8326_), .ZN(new_n8327_));
  NOR2_X1    g08046(.A1(new_n8327_), .A2(new_n8063_), .ZN(new_n8328_));
  NOR2_X1    g08047(.A1(new_n8322_), .A2(new_n8328_), .ZN(new_n8329_));
  INV_X1     g08048(.I(new_n8094_), .ZN(new_n8330_));
  OAI21_X1   g08049(.A1(new_n8330_), .A2(new_n8104_), .B(new_n8102_), .ZN(new_n8331_));
  INV_X1     g08050(.I(new_n8331_), .ZN(new_n8332_));
  NOR2_X1    g08051(.A1(new_n8041_), .A2(new_n8043_), .ZN(new_n8333_));
  NOR2_X1    g08052(.A1(new_n8333_), .A2(new_n8040_), .ZN(new_n8334_));
  NOR2_X1    g08053(.A1(new_n8332_), .A2(new_n8334_), .ZN(new_n8335_));
  INV_X1     g08054(.I(new_n8335_), .ZN(new_n8336_));
  NAND2_X1   g08055(.A1(new_n8332_), .A2(new_n8334_), .ZN(new_n8337_));
  AOI21_X1   g08056(.A1(new_n8336_), .A2(new_n8337_), .B(new_n8329_), .ZN(new_n8338_));
  XOR2_X1    g08057(.A1(new_n8334_), .A2(new_n8331_), .Z(new_n8339_));
  INV_X1     g08058(.I(new_n8339_), .ZN(new_n8340_));
  AOI21_X1   g08059(.A1(new_n8340_), .A2(new_n8329_), .B(new_n8338_), .ZN(new_n8341_));
  XNOR2_X1   g08060(.A1(new_n8341_), .A2(new_n8313_), .ZN(new_n8342_));
  NAND2_X1   g08061(.A1(new_n8342_), .A2(new_n8283_), .ZN(new_n8343_));
  INV_X1     g08062(.I(new_n8313_), .ZN(new_n8344_));
  NOR2_X1    g08063(.A1(new_n8344_), .A2(new_n8341_), .ZN(new_n8345_));
  NAND2_X1   g08064(.A1(new_n8344_), .A2(new_n8341_), .ZN(new_n8346_));
  INV_X1     g08065(.I(new_n8346_), .ZN(new_n8347_));
  OAI21_X1   g08066(.A1(new_n8347_), .A2(new_n8345_), .B(new_n8282_), .ZN(new_n8348_));
  NAND2_X1   g08067(.A1(new_n8343_), .A2(new_n8348_), .ZN(new_n8349_));
  INV_X1     g08068(.I(new_n8349_), .ZN(new_n8350_));
  XOR2_X1    g08069(.A1(new_n8281_), .A2(new_n8350_), .Z(new_n8351_));
  NOR2_X1    g08070(.A1(new_n8351_), .A2(new_n8146_), .ZN(new_n8352_));
  INV_X1     g08071(.I(new_n8146_), .ZN(new_n8353_));
  NOR3_X1    g08072(.A1(new_n8280_), .A2(new_n8278_), .A3(new_n8350_), .ZN(new_n8354_));
  NOR2_X1    g08073(.A1(new_n8281_), .A2(new_n8349_), .ZN(new_n8355_));
  NOR2_X1    g08074(.A1(new_n8355_), .A2(new_n8354_), .ZN(new_n8356_));
  NOR2_X1    g08075(.A1(new_n8356_), .A2(new_n8353_), .ZN(new_n8357_));
  NOR2_X1    g08076(.A1(new_n8352_), .A2(new_n8357_), .ZN(new_n8358_));
  NAND2_X1   g08077(.A1(new_n7924_), .A2(new_n8125_), .ZN(new_n8359_));
  NAND2_X1   g08078(.A1(new_n8359_), .A2(new_n8124_), .ZN(new_n8360_));
  OAI21_X1   g08079(.A1(new_n7927_), .A2(new_n7996_), .B(new_n7997_), .ZN(new_n8361_));
  INV_X1     g08080(.I(new_n8361_), .ZN(new_n8362_));
  OAI21_X1   g08081(.A1(new_n8002_), .A2(new_n8116_), .B(new_n8118_), .ZN(new_n8363_));
  NOR2_X1    g08082(.A1(new_n8016_), .A2(new_n8023_), .ZN(new_n8364_));
  NOR2_X1    g08083(.A1(new_n8364_), .A2(new_n8021_), .ZN(new_n8365_));
  NOR2_X1    g08084(.A1(new_n7944_), .A2(new_n7954_), .ZN(new_n8366_));
  NOR2_X1    g08085(.A1(new_n8366_), .A2(new_n7953_), .ZN(new_n8367_));
  NOR2_X1    g08086(.A1(new_n7984_), .A2(new_n7973_), .ZN(new_n8368_));
  NOR2_X1    g08087(.A1(new_n8368_), .A2(new_n7983_), .ZN(new_n8369_));
  XNOR2_X1   g08088(.A1(new_n8367_), .A2(new_n8369_), .ZN(new_n8370_));
  NOR2_X1    g08089(.A1(new_n8367_), .A2(new_n8369_), .ZN(new_n8371_));
  NAND2_X1   g08090(.A1(new_n8367_), .A2(new_n8369_), .ZN(new_n8372_));
  INV_X1     g08091(.I(new_n8372_), .ZN(new_n8373_));
  OAI21_X1   g08092(.A1(new_n8371_), .A2(new_n8373_), .B(new_n8365_), .ZN(new_n8374_));
  OAI21_X1   g08093(.A1(new_n8370_), .A2(new_n8365_), .B(new_n8374_), .ZN(new_n8375_));
  INV_X1     g08094(.I(new_n8375_), .ZN(new_n8376_));
  INV_X1     g08095(.I(new_n7929_), .ZN(new_n8377_));
  AOI21_X1   g08096(.A1(new_n8377_), .A2(new_n7940_), .B(new_n7938_), .ZN(new_n8378_));
  NOR2_X1    g08097(.A1(new_n8110_), .A2(new_n8080_), .ZN(new_n8379_));
  NOR2_X1    g08098(.A1(new_n8379_), .A2(new_n8109_), .ZN(new_n8380_));
  NOR2_X1    g08099(.A1(new_n8380_), .A2(new_n8378_), .ZN(new_n8381_));
  INV_X1     g08100(.I(new_n8381_), .ZN(new_n8382_));
  NAND2_X1   g08101(.A1(new_n8380_), .A2(new_n8378_), .ZN(new_n8383_));
  AOI21_X1   g08102(.A1(new_n8382_), .A2(new_n8383_), .B(new_n8376_), .ZN(new_n8384_));
  XNOR2_X1   g08103(.A1(new_n8380_), .A2(new_n8378_), .ZN(new_n8385_));
  NOR2_X1    g08104(.A1(new_n8385_), .A2(new_n8375_), .ZN(new_n8386_));
  NOR2_X1    g08105(.A1(new_n8386_), .A2(new_n8384_), .ZN(new_n8387_));
  XNOR2_X1   g08106(.A1(new_n8387_), .A2(new_n8363_), .ZN(new_n8388_));
  NOR2_X1    g08107(.A1(new_n8388_), .A2(new_n8362_), .ZN(new_n8389_));
  NOR2_X1    g08108(.A1(new_n8387_), .A2(new_n8363_), .ZN(new_n8390_));
  INV_X1     g08109(.I(new_n8390_), .ZN(new_n8391_));
  NAND2_X1   g08110(.A1(new_n8387_), .A2(new_n8363_), .ZN(new_n8392_));
  AOI21_X1   g08111(.A1(new_n8391_), .A2(new_n8392_), .B(new_n8361_), .ZN(new_n8393_));
  NOR2_X1    g08112(.A1(new_n8389_), .A2(new_n8393_), .ZN(new_n8394_));
  NOR2_X1    g08113(.A1(new_n8360_), .A2(new_n8394_), .ZN(new_n8395_));
  INV_X1     g08114(.I(new_n8395_), .ZN(new_n8396_));
  NAND2_X1   g08115(.A1(new_n8360_), .A2(new_n8394_), .ZN(new_n8397_));
  AOI21_X1   g08116(.A1(new_n8396_), .A2(new_n8397_), .B(new_n8358_), .ZN(new_n8398_));
  INV_X1     g08117(.I(new_n8358_), .ZN(new_n8399_));
  XNOR2_X1   g08118(.A1(new_n8360_), .A2(new_n8394_), .ZN(new_n8400_));
  NOR2_X1    g08119(.A1(new_n8399_), .A2(new_n8400_), .ZN(new_n8401_));
  NOR2_X1    g08120(.A1(new_n8401_), .A2(new_n8398_), .ZN(new_n8402_));
  OAI21_X1   g08121(.A1(new_n7889_), .A2(new_n8132_), .B(new_n8134_), .ZN(new_n8403_));
  XNOR2_X1   g08122(.A1(new_n8402_), .A2(new_n8403_), .ZN(new_n8404_));
  NAND2_X1   g08123(.A1(new_n8402_), .A2(new_n8403_), .ZN(new_n8405_));
  OR2_X2     g08124(.A1(new_n8402_), .A2(new_n8403_), .Z(new_n8406_));
  NAND2_X1   g08125(.A1(new_n8406_), .A2(new_n8405_), .ZN(new_n8407_));
  NAND2_X1   g08126(.A1(new_n8144_), .A2(new_n8407_), .ZN(new_n8408_));
  OAI21_X1   g08127(.A1(new_n8144_), .A2(new_n8404_), .B(new_n8408_), .ZN(\asquared[61] ));
  NOR2_X1    g08128(.A1(new_n8402_), .A2(new_n8403_), .ZN(new_n8410_));
  OAI21_X1   g08129(.A1(new_n8144_), .A2(new_n8410_), .B(new_n8405_), .ZN(new_n8411_));
  OAI21_X1   g08130(.A1(new_n8399_), .A2(new_n8395_), .B(new_n8397_), .ZN(new_n8412_));
  INV_X1     g08131(.I(new_n8354_), .ZN(new_n8413_));
  AOI21_X1   g08132(.A1(new_n8413_), .A2(new_n8353_), .B(new_n8355_), .ZN(new_n8414_));
  OAI21_X1   g08133(.A1(new_n8362_), .A2(new_n8390_), .B(new_n8392_), .ZN(new_n8415_));
  INV_X1     g08134(.I(new_n8415_), .ZN(new_n8416_));
  OAI21_X1   g08135(.A1(new_n8282_), .A2(new_n8345_), .B(new_n8346_), .ZN(new_n8417_));
  INV_X1     g08136(.I(new_n8417_), .ZN(new_n8418_));
  NAND2_X1   g08137(.A1(new_n8383_), .A2(new_n8376_), .ZN(new_n8419_));
  NAND2_X1   g08138(.A1(new_n8419_), .A2(new_n8382_), .ZN(new_n8420_));
  NOR2_X1    g08139(.A1(new_n8365_), .A2(new_n8373_), .ZN(new_n8421_));
  NOR2_X1    g08140(.A1(new_n8421_), .A2(new_n8371_), .ZN(new_n8422_));
  INV_X1     g08141(.I(new_n8422_), .ZN(new_n8423_));
  INV_X1     g08142(.I(new_n5488_), .ZN(new_n8424_));
  NAND3_X1   g08143(.A1(new_n1786_), .A2(\a[46] ), .A3(\a[51] ), .ZN(new_n8425_));
  INV_X1     g08144(.I(new_n8425_), .ZN(new_n8426_));
  NAND4_X1   g08145(.A1(new_n8426_), .A2(\a[10] ), .A3(\a[51] ), .A4(new_n5841_), .ZN(new_n8427_));
  AOI21_X1   g08146(.A1(new_n8427_), .A2(new_n8424_), .B(new_n1021_), .ZN(new_n8428_));
  NOR3_X1    g08147(.A1(new_n1785_), .A2(new_n5175_), .A3(new_n6260_), .ZN(new_n8429_));
  NOR2_X1    g08148(.A1(new_n650_), .A2(new_n6055_), .ZN(new_n8430_));
  AOI22_X1   g08149(.A1(new_n6280_), .A2(new_n7699_), .B1(new_n8430_), .B2(new_n3061_), .ZN(new_n8431_));
  NOR4_X1    g08150(.A1(new_n6027_), .A2(new_n654_), .A3(new_n675_), .A4(new_n6055_), .ZN(new_n8432_));
  NAND2_X1   g08151(.A1(new_n8431_), .A2(new_n8432_), .ZN(new_n8433_));
  NOR2_X1    g08152(.A1(new_n3175_), .A2(new_n4184_), .ZN(new_n8434_));
  INV_X1     g08153(.I(new_n8434_), .ZN(new_n8435_));
  AOI21_X1   g08154(.A1(\a[29] ), .A2(\a[32] ), .B(new_n3126_), .ZN(new_n8436_));
  INV_X1     g08155(.I(new_n8436_), .ZN(new_n8437_));
  NOR2_X1    g08156(.A1(new_n8435_), .A2(new_n8437_), .ZN(new_n8438_));
  NAND2_X1   g08157(.A1(\a[13] ), .A2(\a[48] ), .ZN(new_n8439_));
  XOR2_X1    g08158(.A1(new_n8438_), .A2(new_n8439_), .Z(new_n8440_));
  NOR2_X1    g08159(.A1(new_n8440_), .A2(new_n8433_), .ZN(new_n8441_));
  INV_X1     g08160(.I(new_n8441_), .ZN(new_n8442_));
  NAND2_X1   g08161(.A1(new_n8440_), .A2(new_n8433_), .ZN(new_n8443_));
  NAND2_X1   g08162(.A1(new_n8442_), .A2(new_n8443_), .ZN(new_n8444_));
  XNOR2_X1   g08163(.A1(new_n8440_), .A2(new_n8433_), .ZN(new_n8445_));
  NOR2_X1    g08164(.A1(new_n8445_), .A2(new_n8429_), .ZN(new_n8446_));
  AOI21_X1   g08165(.A1(new_n8429_), .A2(new_n8444_), .B(new_n8446_), .ZN(new_n8447_));
  NOR2_X1    g08166(.A1(new_n3839_), .A2(new_n2276_), .ZN(new_n8448_));
  NOR2_X1    g08167(.A1(new_n3839_), .A2(new_n2276_), .ZN(new_n8452_));
  INV_X1     g08168(.I(\a[61] ), .ZN(new_n8453_));
  NOR2_X1    g08169(.A1(new_n7216_), .A2(new_n8453_), .ZN(new_n8454_));
  NOR2_X1    g08170(.A1(new_n8085_), .A2(new_n8453_), .ZN(new_n8455_));
  AOI22_X1   g08171(.A1(new_n218_), .A2(new_n8455_), .B1(new_n8454_), .B2(new_n1011_), .ZN(new_n8456_));
  NOR3_X1    g08172(.A1(new_n7650_), .A2(new_n353_), .A3(new_n8085_), .ZN(new_n8457_));
  INV_X1     g08173(.I(new_n8457_), .ZN(new_n8458_));
  NOR2_X1    g08174(.A1(new_n199_), .A2(new_n8453_), .ZN(new_n8459_));
  NOR2_X1    g08175(.A1(new_n7216_), .A2(new_n8085_), .ZN(new_n8460_));
  INV_X1     g08176(.I(new_n8460_), .ZN(new_n8461_));
  NAND4_X1   g08177(.A1(new_n8458_), .A2(new_n233_), .A3(new_n8459_), .A4(new_n8461_), .ZN(new_n8462_));
  NOR2_X1    g08178(.A1(new_n8462_), .A2(new_n8456_), .ZN(new_n8463_));
  INV_X1     g08179(.I(new_n8463_), .ZN(new_n8464_));
  NAND2_X1   g08180(.A1(new_n5592_), .A2(new_n2978_), .ZN(new_n8465_));
  NAND2_X1   g08181(.A1(\a[6] ), .A2(\a[55] ), .ZN(new_n8466_));
  XNOR2_X1   g08182(.A1(new_n8465_), .A2(new_n8466_), .ZN(new_n8467_));
  NOR2_X1    g08183(.A1(new_n8464_), .A2(new_n8467_), .ZN(new_n8468_));
  INV_X1     g08184(.I(new_n8467_), .ZN(new_n8469_));
  NOR2_X1    g08185(.A1(new_n8463_), .A2(new_n8469_), .ZN(new_n8470_));
  NOR2_X1    g08186(.A1(new_n8468_), .A2(new_n8470_), .ZN(new_n8471_));
  XOR2_X1    g08187(.A1(new_n8463_), .A2(new_n8467_), .Z(new_n8472_));
  MUX2_X1    g08188(.I0(new_n8472_), .I1(new_n8471_), .S(new_n8452_), .Z(new_n8473_));
  XOR2_X1    g08189(.A1(new_n8447_), .A2(new_n8473_), .Z(new_n8474_));
  NOR2_X1    g08190(.A1(new_n8447_), .A2(new_n8473_), .ZN(new_n8475_));
  INV_X1     g08191(.I(new_n8475_), .ZN(new_n8476_));
  NAND2_X1   g08192(.A1(new_n8447_), .A2(new_n8473_), .ZN(new_n8477_));
  AOI21_X1   g08193(.A1(new_n8476_), .A2(new_n8477_), .B(new_n8423_), .ZN(new_n8478_));
  AOI21_X1   g08194(.A1(new_n8474_), .A2(new_n8423_), .B(new_n8478_), .ZN(new_n8479_));
  XNOR2_X1   g08195(.A1(new_n8420_), .A2(new_n8479_), .ZN(new_n8480_));
  NOR2_X1    g08196(.A1(new_n8480_), .A2(new_n8418_), .ZN(new_n8481_));
  NOR2_X1    g08197(.A1(new_n8420_), .A2(new_n8479_), .ZN(new_n8482_));
  INV_X1     g08198(.I(new_n8482_), .ZN(new_n8483_));
  NAND2_X1   g08199(.A1(new_n8420_), .A2(new_n8479_), .ZN(new_n8484_));
  AOI21_X1   g08200(.A1(new_n8483_), .A2(new_n8484_), .B(new_n8417_), .ZN(new_n8485_));
  NOR2_X1    g08201(.A1(new_n8481_), .A2(new_n8485_), .ZN(new_n8486_));
  NOR2_X1    g08202(.A1(new_n8215_), .A2(new_n8150_), .ZN(new_n8487_));
  NOR2_X1    g08203(.A1(new_n8487_), .A2(new_n8214_), .ZN(new_n8488_));
  AOI21_X1   g08204(.A1(new_n8151_), .A2(new_n8173_), .B(new_n8171_), .ZN(new_n8489_));
  AOI21_X1   g08205(.A1(new_n1275_), .A2(new_n5321_), .B(new_n8222_), .ZN(new_n8490_));
  INV_X1     g08206(.I(new_n8490_), .ZN(new_n8491_));
  NAND2_X1   g08207(.A1(\a[0] ), .A2(\a[60] ), .ZN(new_n8492_));
  AOI21_X1   g08208(.A1(new_n8156_), .A2(new_n8154_), .B(new_n8492_), .ZN(new_n8493_));
  NOR2_X1    g08209(.A1(new_n8493_), .A2(new_n8157_), .ZN(new_n8494_));
  XOR2_X1    g08210(.A1(new_n8494_), .A2(new_n8183_), .Z(new_n8495_));
  NOR2_X1    g08211(.A1(new_n8495_), .A2(new_n8491_), .ZN(new_n8496_));
  NOR2_X1    g08212(.A1(new_n8494_), .A2(new_n8184_), .ZN(new_n8497_));
  INV_X1     g08213(.I(new_n8497_), .ZN(new_n8498_));
  NAND2_X1   g08214(.A1(new_n8494_), .A2(new_n8184_), .ZN(new_n8499_));
  AOI21_X1   g08215(.A1(new_n8498_), .A2(new_n8499_), .B(new_n8490_), .ZN(new_n8500_));
  NOR2_X1    g08216(.A1(new_n8496_), .A2(new_n8500_), .ZN(new_n8501_));
  NOR2_X1    g08217(.A1(new_n8206_), .A2(new_n8186_), .ZN(new_n8502_));
  NOR2_X1    g08218(.A1(new_n8502_), .A2(new_n8205_), .ZN(new_n8503_));
  XOR2_X1    g08219(.A1(new_n8501_), .A2(new_n8503_), .Z(new_n8504_));
  NOR2_X1    g08220(.A1(new_n8504_), .A2(new_n8489_), .ZN(new_n8505_));
  INV_X1     g08221(.I(new_n8501_), .ZN(new_n8506_));
  NOR2_X1    g08222(.A1(new_n8506_), .A2(new_n8503_), .ZN(new_n8507_));
  INV_X1     g08223(.I(new_n8507_), .ZN(new_n8508_));
  NAND2_X1   g08224(.A1(new_n8506_), .A2(new_n8503_), .ZN(new_n8509_));
  NAND2_X1   g08225(.A1(new_n8508_), .A2(new_n8509_), .ZN(new_n8510_));
  AOI21_X1   g08226(.A1(new_n8489_), .A2(new_n8510_), .B(new_n8505_), .ZN(new_n8511_));
  INV_X1     g08227(.I(new_n8191_), .ZN(new_n8512_));
  OAI21_X1   g08228(.A1(new_n8190_), .A2(new_n8512_), .B(new_n8188_), .ZN(new_n8513_));
  NOR2_X1    g08229(.A1(new_n8231_), .A2(new_n8229_), .ZN(new_n8514_));
  AOI21_X1   g08230(.A1(new_n267_), .A2(new_n8242_), .B(new_n8248_), .ZN(new_n8515_));
  INV_X1     g08231(.I(new_n8515_), .ZN(new_n8516_));
  XOR2_X1    g08232(.A1(new_n8514_), .A2(new_n8516_), .Z(new_n8517_));
  NOR2_X1    g08233(.A1(new_n8517_), .A2(new_n8513_), .ZN(new_n8518_));
  INV_X1     g08234(.I(new_n8513_), .ZN(new_n8519_));
  INV_X1     g08235(.I(new_n8514_), .ZN(new_n8520_));
  NOR2_X1    g08236(.A1(new_n8520_), .A2(new_n8516_), .ZN(new_n8521_));
  NOR2_X1    g08237(.A1(new_n8514_), .A2(new_n8515_), .ZN(new_n8522_));
  NOR2_X1    g08238(.A1(new_n8521_), .A2(new_n8522_), .ZN(new_n8523_));
  NOR2_X1    g08239(.A1(new_n8523_), .A2(new_n8519_), .ZN(new_n8524_));
  NOR2_X1    g08240(.A1(new_n8524_), .A2(new_n8518_), .ZN(new_n8525_));
  INV_X1     g08241(.I(new_n8261_), .ZN(new_n8526_));
  AOI21_X1   g08242(.A1(new_n8526_), .A2(new_n8264_), .B(new_n8259_), .ZN(new_n8527_));
  INV_X1     g08243(.I(new_n8527_), .ZN(new_n8528_));
  AOI21_X1   g08244(.A1(new_n8162_), .A2(new_n8163_), .B(new_n8160_), .ZN(new_n8529_));
  AOI21_X1   g08245(.A1(new_n4538_), .A2(new_n5339_), .B(new_n8253_), .ZN(new_n8530_));
  AOI21_X1   g08246(.A1(new_n2752_), .A2(new_n3487_), .B(new_n8256_), .ZN(new_n8531_));
  XOR2_X1    g08247(.A1(new_n8530_), .A2(new_n8531_), .Z(new_n8532_));
  NAND2_X1   g08248(.A1(new_n8532_), .A2(new_n8529_), .ZN(new_n8533_));
  INV_X1     g08249(.I(new_n8529_), .ZN(new_n8534_));
  AND2_X2    g08250(.A1(new_n8530_), .A2(new_n8531_), .Z(new_n8535_));
  NOR2_X1    g08251(.A1(new_n8530_), .A2(new_n8531_), .ZN(new_n8536_));
  OAI21_X1   g08252(.A1(new_n8535_), .A2(new_n8536_), .B(new_n8534_), .ZN(new_n8537_));
  AOI21_X1   g08253(.A1(new_n8533_), .A2(new_n8537_), .B(new_n8528_), .ZN(new_n8538_));
  NAND2_X1   g08254(.A1(new_n8533_), .A2(new_n8537_), .ZN(new_n8539_));
  NOR2_X1    g08255(.A1(new_n8539_), .A2(new_n8527_), .ZN(new_n8540_));
  NOR2_X1    g08256(.A1(new_n8540_), .A2(new_n8538_), .ZN(new_n8541_));
  NOR2_X1    g08257(.A1(new_n8541_), .A2(new_n8525_), .ZN(new_n8542_));
  XOR2_X1    g08258(.A1(new_n8539_), .A2(new_n8528_), .Z(new_n8543_));
  INV_X1     g08259(.I(new_n8543_), .ZN(new_n8544_));
  AOI21_X1   g08260(.A1(new_n8544_), .A2(new_n8525_), .B(new_n8542_), .ZN(new_n8545_));
  NOR2_X1    g08261(.A1(new_n8511_), .A2(new_n8545_), .ZN(new_n8546_));
  INV_X1     g08262(.I(new_n8546_), .ZN(new_n8547_));
  NAND2_X1   g08263(.A1(new_n8511_), .A2(new_n8545_), .ZN(new_n8548_));
  AOI21_X1   g08264(.A1(new_n8547_), .A2(new_n8548_), .B(new_n8488_), .ZN(new_n8549_));
  XNOR2_X1   g08265(.A1(new_n8511_), .A2(new_n8545_), .ZN(new_n8550_));
  NOR3_X1    g08266(.A1(new_n8550_), .A2(new_n8214_), .A3(new_n8487_), .ZN(new_n8551_));
  NOR2_X1    g08267(.A1(new_n8551_), .A2(new_n8549_), .ZN(new_n8552_));
  XOR2_X1    g08268(.A1(new_n8486_), .A2(new_n8552_), .Z(new_n8553_));
  NOR3_X1    g08269(.A1(new_n8481_), .A2(new_n8485_), .A3(new_n8552_), .ZN(new_n8554_));
  NOR3_X1    g08270(.A1(new_n8486_), .A2(new_n8549_), .A3(new_n8551_), .ZN(new_n8555_));
  OAI21_X1   g08271(.A1(new_n8555_), .A2(new_n8554_), .B(new_n8416_), .ZN(new_n8556_));
  OAI21_X1   g08272(.A1(new_n8553_), .A2(new_n8416_), .B(new_n8556_), .ZN(new_n8557_));
  AOI21_X1   g08273(.A1(new_n8147_), .A2(new_n8275_), .B(new_n8276_), .ZN(new_n8558_));
  OAI21_X1   g08274(.A1(new_n8285_), .A2(new_n8309_), .B(new_n8310_), .ZN(new_n8559_));
  INV_X1     g08275(.I(new_n8559_), .ZN(new_n8560_));
  NAND2_X1   g08276(.A1(new_n8337_), .A2(new_n8329_), .ZN(new_n8561_));
  NAND2_X1   g08277(.A1(new_n8561_), .A2(new_n8336_), .ZN(new_n8562_));
  INV_X1     g08278(.I(new_n8562_), .ZN(new_n8563_));
  NOR2_X1    g08279(.A1(new_n4770_), .A2(new_n6692_), .ZN(new_n8564_));
  INV_X1     g08280(.I(new_n8564_), .ZN(new_n8565_));
  NOR2_X1    g08281(.A1(new_n8565_), .A2(new_n1965_), .ZN(new_n8566_));
  NOR2_X1    g08282(.A1(new_n8565_), .A2(new_n1965_), .ZN(new_n8570_));
  NAND2_X1   g08283(.A1(new_n7482_), .A2(new_n609_), .ZN(new_n8571_));
  NOR2_X1    g08284(.A1(new_n1339_), .A2(new_n4769_), .ZN(new_n8572_));
  XOR2_X1    g08285(.A1(new_n8571_), .A2(new_n8572_), .Z(new_n8573_));
  NOR2_X1    g08286(.A1(new_n2534_), .A2(new_n3036_), .ZN(new_n8574_));
  NOR2_X1    g08287(.A1(new_n7008_), .A2(new_n8574_), .ZN(new_n8575_));
  NOR4_X1    g08288(.A1(new_n4372_), .A2(new_n2797_), .A3(new_n1916_), .A4(new_n3423_), .ZN(new_n8576_));
  NAND2_X1   g08289(.A1(new_n8575_), .A2(new_n8576_), .ZN(new_n8577_));
  OR2_X2     g08290(.A1(new_n8577_), .A2(new_n8573_), .Z(new_n8578_));
  NAND2_X1   g08291(.A1(new_n8577_), .A2(new_n8573_), .ZN(new_n8579_));
  NAND2_X1   g08292(.A1(new_n8578_), .A2(new_n8579_), .ZN(new_n8580_));
  XNOR2_X1   g08293(.A1(new_n8577_), .A2(new_n8573_), .ZN(new_n8581_));
  NOR2_X1    g08294(.A1(new_n8581_), .A2(new_n8570_), .ZN(new_n8582_));
  AOI21_X1   g08295(.A1(new_n8570_), .A2(new_n8580_), .B(new_n8582_), .ZN(new_n8583_));
  NOR2_X1    g08296(.A1(new_n8563_), .A2(new_n8583_), .ZN(new_n8584_));
  INV_X1     g08297(.I(new_n8583_), .ZN(new_n8585_));
  NOR2_X1    g08298(.A1(new_n8562_), .A2(new_n8585_), .ZN(new_n8586_));
  NOR2_X1    g08299(.A1(new_n8584_), .A2(new_n8586_), .ZN(new_n8587_));
  NOR2_X1    g08300(.A1(new_n8587_), .A2(new_n8560_), .ZN(new_n8588_));
  XOR2_X1    g08301(.A1(new_n8562_), .A2(new_n8583_), .Z(new_n8589_));
  NOR2_X1    g08302(.A1(new_n8589_), .A2(new_n8559_), .ZN(new_n8590_));
  NOR2_X1    g08303(.A1(new_n8588_), .A2(new_n8590_), .ZN(new_n8591_));
  NOR2_X1    g08304(.A1(new_n8219_), .A2(new_n8272_), .ZN(new_n8592_));
  AOI21_X1   g08305(.A1(new_n8296_), .A2(new_n8304_), .B(new_n8302_), .ZN(new_n8593_));
  INV_X1     g08306(.I(new_n8326_), .ZN(new_n8594_));
  AOI21_X1   g08307(.A1(new_n8063_), .A2(new_n8594_), .B(new_n8325_), .ZN(new_n8595_));
  NAND2_X1   g08308(.A1(new_n8245_), .A2(new_n267_), .ZN(new_n8596_));
  NAND2_X1   g08309(.A1(\a[23] ), .A2(\a[38] ), .ZN(new_n8597_));
  XNOR2_X1   g08310(.A1(new_n8596_), .A2(new_n8597_), .ZN(new_n8598_));
  NOR2_X1    g08311(.A1(new_n8595_), .A2(new_n8598_), .ZN(new_n8599_));
  AND2_X2    g08312(.A1(new_n8595_), .A2(new_n8598_), .Z(new_n8600_));
  NOR2_X1    g08313(.A1(new_n8600_), .A2(new_n8599_), .ZN(new_n8601_));
  NOR2_X1    g08314(.A1(new_n8601_), .A2(new_n8593_), .ZN(new_n8602_));
  INV_X1     g08315(.I(new_n8593_), .ZN(new_n8603_));
  XNOR2_X1   g08316(.A1(new_n8595_), .A2(new_n8598_), .ZN(new_n8604_));
  NOR2_X1    g08317(.A1(new_n8603_), .A2(new_n8604_), .ZN(new_n8605_));
  NOR2_X1    g08318(.A1(new_n8605_), .A2(new_n8602_), .ZN(new_n8606_));
  INV_X1     g08319(.I(new_n8606_), .ZN(new_n8607_));
  INV_X1     g08320(.I(new_n8239_), .ZN(new_n8608_));
  AOI21_X1   g08321(.A1(new_n8220_), .A2(new_n8608_), .B(new_n8238_), .ZN(new_n8609_));
  NOR2_X1    g08322(.A1(new_n8291_), .A2(new_n8293_), .ZN(new_n8610_));
  NOR2_X1    g08323(.A1(new_n8610_), .A2(new_n8292_), .ZN(new_n8611_));
  AOI21_X1   g08324(.A1(new_n1220_), .A2(new_n6030_), .B(new_n8201_), .ZN(new_n8612_));
  NAND2_X1   g08325(.A1(new_n3733_), .A2(new_n8155_), .ZN(new_n8613_));
  NAND2_X1   g08326(.A1(\a[1] ), .A2(\a[60] ), .ZN(new_n8614_));
  XOR2_X1    g08327(.A1(new_n8614_), .A2(\a[31] ), .Z(new_n8615_));
  XOR2_X1    g08328(.A1(new_n8615_), .A2(new_n8613_), .Z(new_n8616_));
  NAND2_X1   g08329(.A1(new_n8612_), .A2(new_n8616_), .ZN(new_n8617_));
  INV_X1     g08330(.I(new_n8612_), .ZN(new_n8618_));
  NOR2_X1    g08331(.A1(new_n8615_), .A2(new_n8613_), .ZN(new_n8619_));
  NAND2_X1   g08332(.A1(new_n8615_), .A2(new_n8613_), .ZN(new_n8620_));
  INV_X1     g08333(.I(new_n8620_), .ZN(new_n8621_));
  OAI21_X1   g08334(.A1(new_n8619_), .A2(new_n8621_), .B(new_n8618_), .ZN(new_n8622_));
  NAND2_X1   g08335(.A1(new_n8622_), .A2(new_n8617_), .ZN(new_n8623_));
  XNOR2_X1   g08336(.A1(new_n8611_), .A2(new_n8623_), .ZN(new_n8624_));
  NOR2_X1    g08337(.A1(new_n8624_), .A2(new_n8609_), .ZN(new_n8625_));
  INV_X1     g08338(.I(new_n8609_), .ZN(new_n8626_));
  AND2_X2    g08339(.A1(new_n8611_), .A2(new_n8623_), .Z(new_n8627_));
  NOR2_X1    g08340(.A1(new_n8611_), .A2(new_n8623_), .ZN(new_n8628_));
  NOR2_X1    g08341(.A1(new_n8627_), .A2(new_n8628_), .ZN(new_n8629_));
  NOR2_X1    g08342(.A1(new_n8629_), .A2(new_n8626_), .ZN(new_n8630_));
  NOR2_X1    g08343(.A1(new_n8630_), .A2(new_n8625_), .ZN(new_n8631_));
  XOR2_X1    g08344(.A1(new_n8631_), .A2(new_n8607_), .Z(new_n8632_));
  OAI21_X1   g08345(.A1(new_n8270_), .A2(new_n8592_), .B(new_n8632_), .ZN(new_n8633_));
  NOR2_X1    g08346(.A1(new_n8592_), .A2(new_n8270_), .ZN(new_n8634_));
  NOR2_X1    g08347(.A1(new_n8631_), .A2(new_n8607_), .ZN(new_n8635_));
  NAND2_X1   g08348(.A1(new_n8631_), .A2(new_n8607_), .ZN(new_n8636_));
  INV_X1     g08349(.I(new_n8636_), .ZN(new_n8637_));
  OAI21_X1   g08350(.A1(new_n8637_), .A2(new_n8635_), .B(new_n8634_), .ZN(new_n8638_));
  NAND2_X1   g08351(.A1(new_n8633_), .A2(new_n8638_), .ZN(new_n8639_));
  INV_X1     g08352(.I(new_n8639_), .ZN(new_n8640_));
  XOR2_X1    g08353(.A1(new_n8591_), .A2(new_n8640_), .Z(new_n8641_));
  INV_X1     g08354(.I(new_n8591_), .ZN(new_n8642_));
  NOR2_X1    g08355(.A1(new_n8642_), .A2(new_n8640_), .ZN(new_n8643_));
  NOR2_X1    g08356(.A1(new_n8591_), .A2(new_n8639_), .ZN(new_n8644_));
  NOR2_X1    g08357(.A1(new_n8643_), .A2(new_n8644_), .ZN(new_n8645_));
  MUX2_X1    g08358(.I0(new_n8641_), .I1(new_n8645_), .S(new_n8558_), .Z(new_n8646_));
  XOR2_X1    g08359(.A1(new_n8557_), .A2(new_n8646_), .Z(new_n8647_));
  NOR2_X1    g08360(.A1(new_n8647_), .A2(new_n8414_), .ZN(new_n8648_));
  XNOR2_X1   g08361(.A1(new_n8557_), .A2(new_n8646_), .ZN(new_n8649_));
  INV_X1     g08362(.I(new_n8649_), .ZN(new_n8650_));
  AOI21_X1   g08363(.A1(new_n8414_), .A2(new_n8650_), .B(new_n8648_), .ZN(new_n8651_));
  XOR2_X1    g08364(.A1(new_n8651_), .A2(new_n8412_), .Z(new_n8652_));
  NAND2_X1   g08365(.A1(new_n8411_), .A2(new_n8652_), .ZN(new_n8653_));
  NOR2_X1    g08366(.A1(new_n8651_), .A2(new_n8412_), .ZN(new_n8654_));
  NAND2_X1   g08367(.A1(new_n8651_), .A2(new_n8412_), .ZN(new_n8655_));
  INV_X1     g08368(.I(new_n8655_), .ZN(new_n8656_));
  NOR2_X1    g08369(.A1(new_n8656_), .A2(new_n8654_), .ZN(new_n8657_));
  OAI21_X1   g08370(.A1(new_n8411_), .A2(new_n8657_), .B(new_n8653_), .ZN(\asquared[62] ));
  INV_X1     g08371(.I(new_n8654_), .ZN(new_n8659_));
  NOR2_X1    g08372(.A1(new_n8655_), .A2(new_n8402_), .ZN(new_n8660_));
  NOR2_X1    g08373(.A1(new_n8660_), .A2(new_n8403_), .ZN(new_n8661_));
  AOI21_X1   g08374(.A1(new_n8402_), .A2(new_n8655_), .B(new_n8661_), .ZN(new_n8662_));
  INV_X1     g08375(.I(new_n8662_), .ZN(new_n8663_));
  NOR3_X1    g08376(.A1(new_n8144_), .A2(new_n8659_), .A3(new_n8663_), .ZN(\asquared[63] ));
  INV_X1     g08377(.I(new_n8644_), .ZN(new_n8665_));
  OAI21_X1   g08378(.A1(new_n8558_), .A2(new_n8643_), .B(new_n8665_), .ZN(new_n8666_));
  INV_X1     g08379(.I(new_n8666_), .ZN(new_n8667_));
  AOI21_X1   g08380(.A1(new_n8423_), .A2(new_n8477_), .B(new_n8475_), .ZN(new_n8668_));
  INV_X1     g08381(.I(new_n8600_), .ZN(new_n8669_));
  AOI21_X1   g08382(.A1(new_n8603_), .A2(new_n8669_), .B(new_n8599_), .ZN(new_n8670_));
  AOI21_X1   g08383(.A1(new_n1441_), .A2(new_n5321_), .B(new_n8566_), .ZN(new_n8671_));
  NOR2_X1    g08384(.A1(new_n8428_), .A2(new_n8426_), .ZN(new_n8672_));
  INV_X1     g08385(.I(new_n8672_), .ZN(new_n8673_));
  NOR2_X1    g08386(.A1(new_n7727_), .A2(new_n8085_), .ZN(new_n8674_));
  INV_X1     g08387(.I(new_n8674_), .ZN(new_n8675_));
  NOR2_X1    g08388(.A1(new_n7647_), .A2(new_n8085_), .ZN(new_n8676_));
  INV_X1     g08389(.I(new_n8676_), .ZN(new_n8677_));
  NOR2_X1    g08390(.A1(new_n8675_), .A2(new_n8677_), .ZN(new_n8678_));
  NOR2_X1    g08391(.A1(new_n8678_), .A2(new_n1713_), .ZN(new_n8679_));
  NOR4_X1    g08392(.A1(new_n8245_), .A2(new_n229_), .A3(new_n200_), .A4(new_n8085_), .ZN(new_n8680_));
  NAND2_X1   g08393(.A1(new_n8679_), .A2(new_n8680_), .ZN(new_n8681_));
  NOR2_X1    g08394(.A1(new_n8673_), .A2(new_n8681_), .ZN(new_n8682_));
  AOI21_X1   g08395(.A1(new_n8679_), .A2(new_n8680_), .B(new_n8672_), .ZN(new_n8683_));
  NOR2_X1    g08396(.A1(new_n8682_), .A2(new_n8683_), .ZN(new_n8684_));
  XOR2_X1    g08397(.A1(new_n8672_), .A2(new_n8681_), .Z(new_n8685_));
  MUX2_X1    g08398(.I0(new_n8685_), .I1(new_n8684_), .S(new_n8671_), .Z(new_n8686_));
  NAND2_X1   g08399(.A1(new_n8579_), .A2(new_n8570_), .ZN(new_n8687_));
  NAND2_X1   g08400(.A1(new_n8687_), .A2(new_n8578_), .ZN(new_n8688_));
  XOR2_X1    g08401(.A1(new_n8686_), .A2(new_n8688_), .Z(new_n8689_));
  NOR2_X1    g08402(.A1(new_n8689_), .A2(new_n8670_), .ZN(new_n8690_));
  INV_X1     g08403(.I(new_n8670_), .ZN(new_n8691_));
  INV_X1     g08404(.I(new_n8688_), .ZN(new_n8692_));
  NOR2_X1    g08405(.A1(new_n8686_), .A2(new_n8692_), .ZN(new_n8693_));
  INV_X1     g08406(.I(new_n8693_), .ZN(new_n8694_));
  NAND2_X1   g08407(.A1(new_n8686_), .A2(new_n8692_), .ZN(new_n8695_));
  AOI21_X1   g08408(.A1(new_n8694_), .A2(new_n8695_), .B(new_n8691_), .ZN(new_n8696_));
  NOR2_X1    g08409(.A1(new_n8690_), .A2(new_n8696_), .ZN(new_n8697_));
  AOI21_X1   g08410(.A1(new_n8490_), .A2(new_n8499_), .B(new_n8497_), .ZN(new_n8698_));
  INV_X1     g08411(.I(new_n8698_), .ZN(new_n8699_));
  OAI21_X1   g08412(.A1(new_n8618_), .A2(new_n8619_), .B(new_n8620_), .ZN(new_n8700_));
  INV_X1     g08413(.I(new_n8700_), .ZN(new_n8701_));
  NOR2_X1    g08414(.A1(new_n8536_), .A2(new_n8534_), .ZN(new_n8702_));
  NOR2_X1    g08415(.A1(new_n8702_), .A2(new_n8535_), .ZN(new_n8703_));
  XOR2_X1    g08416(.A1(new_n8703_), .A2(new_n8701_), .Z(new_n8704_));
  NAND2_X1   g08417(.A1(new_n8704_), .A2(new_n8699_), .ZN(new_n8705_));
  NOR2_X1    g08418(.A1(new_n8703_), .A2(new_n8701_), .ZN(new_n8706_));
  NAND2_X1   g08419(.A1(new_n8703_), .A2(new_n8701_), .ZN(new_n8707_));
  INV_X1     g08420(.I(new_n8707_), .ZN(new_n8708_));
  OAI21_X1   g08421(.A1(new_n8708_), .A2(new_n8706_), .B(new_n8698_), .ZN(new_n8709_));
  NAND2_X1   g08422(.A1(new_n8705_), .A2(new_n8709_), .ZN(new_n8710_));
  XOR2_X1    g08423(.A1(new_n8697_), .A2(new_n8710_), .Z(new_n8711_));
  NOR2_X1    g08424(.A1(new_n8711_), .A2(new_n8668_), .ZN(new_n8712_));
  INV_X1     g08425(.I(new_n8668_), .ZN(new_n8713_));
  INV_X1     g08426(.I(new_n8710_), .ZN(new_n8714_));
  NOR2_X1    g08427(.A1(new_n8697_), .A2(new_n8714_), .ZN(new_n8715_));
  INV_X1     g08428(.I(new_n8715_), .ZN(new_n8716_));
  NAND2_X1   g08429(.A1(new_n8697_), .A2(new_n8714_), .ZN(new_n8717_));
  AOI21_X1   g08430(.A1(new_n8716_), .A2(new_n8717_), .B(new_n8713_), .ZN(new_n8718_));
  NOR2_X1    g08431(.A1(new_n8712_), .A2(new_n8718_), .ZN(new_n8719_));
  OAI21_X1   g08432(.A1(new_n8488_), .A2(new_n8546_), .B(new_n8548_), .ZN(new_n8720_));
  INV_X1     g08433(.I(new_n8720_), .ZN(new_n8721_));
  OAI21_X1   g08434(.A1(new_n8634_), .A2(new_n8635_), .B(new_n8636_), .ZN(new_n8722_));
  NOR2_X1    g08435(.A1(new_n885_), .A2(new_n6692_), .ZN(new_n8723_));
  NAND2_X1   g08436(.A1(\a[9] ), .A2(\a[10] ), .ZN(new_n8725_));
  NOR2_X1    g08437(.A1(new_n8056_), .A2(new_n8725_), .ZN(new_n8726_));
  INV_X1     g08438(.I(new_n8726_), .ZN(new_n8727_));
  NOR2_X1    g08439(.A1(new_n364_), .A2(new_n6694_), .ZN(new_n8728_));
  NAND2_X1   g08440(.A1(new_n7024_), .A2(new_n8723_), .ZN(new_n8729_));
  NAND2_X1   g08441(.A1(new_n8727_), .A2(new_n8729_), .ZN(new_n8730_));
  INV_X1     g08442(.I(new_n8730_), .ZN(new_n8731_));
  AOI21_X1   g08443(.A1(\a[45] ), .A2(\a[52] ), .B(new_n2062_), .ZN(new_n8732_));
  AOI22_X1   g08444(.A1(new_n8731_), .A2(new_n8732_), .B1(new_n8727_), .B2(new_n8728_), .ZN(new_n8733_));
  INV_X1     g08445(.I(new_n8733_), .ZN(new_n8734_));
  NAND2_X1   g08446(.A1(new_n2752_), .A2(new_n3838_), .ZN(new_n8735_));
  NAND2_X1   g08447(.A1(\a[21] ), .A2(\a[41] ), .ZN(new_n8736_));
  XNOR2_X1   g08448(.A1(new_n8735_), .A2(new_n8736_), .ZN(new_n8737_));
  NAND2_X1   g08449(.A1(\a[60] ), .A2(\a[62] ), .ZN(new_n8738_));
  XNOR2_X1   g08450(.A1(new_n197_), .A2(new_n8738_), .ZN(new_n8739_));
  NOR2_X1    g08451(.A1(new_n8737_), .A2(new_n8739_), .ZN(new_n8740_));
  INV_X1     g08452(.I(new_n8740_), .ZN(new_n8741_));
  AND2_X2    g08453(.A1(new_n8737_), .A2(new_n8739_), .Z(new_n8742_));
  INV_X1     g08454(.I(new_n8742_), .ZN(new_n8743_));
  AOI21_X1   g08455(.A1(new_n8743_), .A2(new_n8741_), .B(new_n8734_), .ZN(new_n8744_));
  XNOR2_X1   g08456(.A1(new_n8737_), .A2(new_n8739_), .ZN(new_n8745_));
  NOR2_X1    g08457(.A1(new_n8745_), .A2(new_n8733_), .ZN(new_n8746_));
  NOR2_X1    g08458(.A1(new_n8744_), .A2(new_n8746_), .ZN(new_n8747_));
  INV_X1     g08459(.I(new_n8747_), .ZN(new_n8748_));
  NAND2_X1   g08460(.A1(\a[46] ), .A2(\a[47] ), .ZN(new_n8749_));
  NOR3_X1    g08461(.A1(new_n868_), .A2(new_n5511_), .A3(new_n6260_), .ZN(new_n8751_));
  AOI22_X1   g08462(.A1(new_n654_), .A2(new_n6280_), .B1(new_n6056_), .B2(new_n1220_), .ZN(new_n8752_));
  NOR4_X1    g08463(.A1(new_n6028_), .A2(new_n787_), .A3(new_n566_), .A4(new_n6055_), .ZN(new_n8753_));
  NAND2_X1   g08464(.A1(new_n8752_), .A2(new_n8753_), .ZN(new_n8754_));
  NOR2_X1    g08465(.A1(new_n6999_), .A2(new_n7216_), .ZN(new_n8755_));
  NAND2_X1   g08466(.A1(new_n8755_), .A2(new_n479_), .ZN(new_n8756_));
  NOR2_X1    g08467(.A1(new_n1215_), .A2(new_n4769_), .ZN(new_n8757_));
  XOR2_X1    g08468(.A1(new_n8756_), .A2(new_n8757_), .Z(new_n8758_));
  NOR2_X1    g08469(.A1(new_n8758_), .A2(new_n8754_), .ZN(new_n8759_));
  NAND2_X1   g08470(.A1(new_n8758_), .A2(new_n8754_), .ZN(new_n8760_));
  INV_X1     g08471(.I(new_n8760_), .ZN(new_n8761_));
  OAI21_X1   g08472(.A1(new_n8761_), .A2(new_n8759_), .B(new_n8751_), .ZN(new_n8762_));
  INV_X1     g08473(.I(new_n8751_), .ZN(new_n8763_));
  XOR2_X1    g08474(.A1(new_n8758_), .A2(new_n8754_), .Z(new_n8764_));
  NAND2_X1   g08475(.A1(new_n8764_), .A2(new_n8763_), .ZN(new_n8765_));
  NAND2_X1   g08476(.A1(new_n8765_), .A2(new_n8762_), .ZN(new_n8766_));
  NOR2_X1    g08477(.A1(new_n4501_), .A2(new_n6945_), .ZN(new_n8767_));
  AOI22_X1   g08478(.A1(new_n2060_), .A2(new_n8767_), .B1(new_n5321_), .B2(new_n2331_), .ZN(new_n8768_));
  INV_X1     g08479(.I(new_n8768_), .ZN(new_n8769_));
  NOR3_X1    g08480(.A1(new_n8181_), .A2(new_n4770_), .A3(new_n6945_), .ZN(new_n8770_));
  NAND2_X1   g08481(.A1(\a[19] ), .A2(\a[43] ), .ZN(new_n8771_));
  AOI21_X1   g08482(.A1(\a[44] ), .A2(\a[54] ), .B(new_n1918_), .ZN(new_n8772_));
  NAND4_X1   g08483(.A1(new_n8769_), .A2(new_n8770_), .A3(new_n8771_), .A4(new_n8772_), .ZN(new_n8773_));
  INV_X1     g08484(.I(new_n8773_), .ZN(new_n8774_));
  AOI22_X1   g08485(.A1(new_n2500_), .A2(new_n3487_), .B1(new_n3424_), .B2(new_n2797_), .ZN(new_n8775_));
  NOR4_X1    g08486(.A1(new_n4372_), .A2(new_n2690_), .A3(new_n2098_), .A4(new_n3423_), .ZN(new_n8776_));
  NAND2_X1   g08487(.A1(new_n8775_), .A2(new_n8776_), .ZN(new_n8777_));
  NOR2_X1    g08488(.A1(new_n2384_), .A2(new_n2285_), .ZN(new_n8778_));
  NOR2_X1    g08489(.A1(new_n8252_), .A2(new_n8778_), .ZN(new_n8779_));
  NOR4_X1    g08490(.A1(new_n5339_), .A2(new_n2543_), .A3(new_n1674_), .A4(new_n4240_), .ZN(new_n8780_));
  NAND2_X1   g08491(.A1(new_n8779_), .A2(new_n8780_), .ZN(new_n8781_));
  NOR2_X1    g08492(.A1(new_n8781_), .A2(new_n8777_), .ZN(new_n8782_));
  AOI22_X1   g08493(.A1(new_n8779_), .A2(new_n8780_), .B1(new_n8775_), .B2(new_n8776_), .ZN(new_n8783_));
  OAI21_X1   g08494(.A1(new_n8782_), .A2(new_n8783_), .B(new_n8774_), .ZN(new_n8784_));
  XOR2_X1    g08495(.A1(new_n8781_), .A2(new_n8777_), .Z(new_n8785_));
  NAND2_X1   g08496(.A1(new_n8785_), .A2(new_n8773_), .ZN(new_n8786_));
  NAND2_X1   g08497(.A1(new_n8786_), .A2(new_n8784_), .ZN(new_n8787_));
  XOR2_X1    g08498(.A1(new_n8787_), .A2(new_n8766_), .Z(new_n8788_));
  INV_X1     g08499(.I(new_n8766_), .ZN(new_n8789_));
  INV_X1     g08500(.I(new_n8787_), .ZN(new_n8790_));
  NOR2_X1    g08501(.A1(new_n8790_), .A2(new_n8789_), .ZN(new_n8791_));
  NOR2_X1    g08502(.A1(new_n8787_), .A2(new_n8766_), .ZN(new_n8792_));
  NOR2_X1    g08503(.A1(new_n8791_), .A2(new_n8792_), .ZN(new_n8793_));
  NOR2_X1    g08504(.A1(new_n8793_), .A2(new_n8748_), .ZN(new_n8794_));
  AOI21_X1   g08505(.A1(new_n8748_), .A2(new_n8788_), .B(new_n8794_), .ZN(new_n8795_));
  NOR2_X1    g08506(.A1(new_n8722_), .A2(new_n8795_), .ZN(new_n8796_));
  INV_X1     g08507(.I(new_n8796_), .ZN(new_n8797_));
  NAND2_X1   g08508(.A1(new_n8722_), .A2(new_n8795_), .ZN(new_n8798_));
  AOI21_X1   g08509(.A1(new_n8797_), .A2(new_n8798_), .B(new_n8721_), .ZN(new_n8799_));
  XOR2_X1    g08510(.A1(new_n8722_), .A2(new_n8795_), .Z(new_n8800_));
  AOI21_X1   g08511(.A1(new_n8721_), .A2(new_n8800_), .B(new_n8799_), .ZN(new_n8801_));
  XOR2_X1    g08512(.A1(new_n8801_), .A2(new_n8719_), .Z(new_n8802_));
  NOR2_X1    g08513(.A1(new_n8802_), .A2(new_n8667_), .ZN(new_n8803_));
  INV_X1     g08514(.I(new_n8719_), .ZN(new_n8804_));
  NOR2_X1    g08515(.A1(new_n8801_), .A2(new_n8804_), .ZN(new_n8805_));
  INV_X1     g08516(.I(new_n8805_), .ZN(new_n8806_));
  NAND2_X1   g08517(.A1(new_n8801_), .A2(new_n8804_), .ZN(new_n8807_));
  AOI21_X1   g08518(.A1(new_n8806_), .A2(new_n8807_), .B(new_n8666_), .ZN(new_n8808_));
  INV_X1     g08519(.I(new_n8586_), .ZN(new_n8809_));
  AOI21_X1   g08520(.A1(new_n8559_), .A2(new_n8809_), .B(new_n8584_), .ZN(new_n8810_));
  INV_X1     g08521(.I(new_n8522_), .ZN(new_n8811_));
  AOI21_X1   g08522(.A1(new_n8519_), .A2(new_n8811_), .B(new_n8521_), .ZN(new_n8812_));
  INV_X1     g08523(.I(new_n8470_), .ZN(new_n8813_));
  AOI21_X1   g08524(.A1(new_n8452_), .A2(new_n8813_), .B(new_n8468_), .ZN(new_n8814_));
  NAND2_X1   g08525(.A1(new_n8443_), .A2(new_n8429_), .ZN(new_n8815_));
  NAND2_X1   g08526(.A1(new_n8815_), .A2(new_n8442_), .ZN(new_n8816_));
  XOR2_X1    g08527(.A1(new_n8816_), .A2(new_n8814_), .Z(new_n8817_));
  AOI21_X1   g08528(.A1(new_n8815_), .A2(new_n8442_), .B(new_n8814_), .ZN(new_n8818_));
  INV_X1     g08529(.I(new_n8814_), .ZN(new_n8819_));
  NOR2_X1    g08530(.A1(new_n8816_), .A2(new_n8819_), .ZN(new_n8820_));
  OAI21_X1   g08531(.A1(new_n8820_), .A2(new_n8818_), .B(new_n8812_), .ZN(new_n8821_));
  OAI21_X1   g08532(.A1(new_n8812_), .A2(new_n8817_), .B(new_n8821_), .ZN(new_n8822_));
  AOI21_X1   g08533(.A1(new_n2383_), .A2(new_n5601_), .B(new_n8448_), .ZN(new_n8823_));
  INV_X1     g08534(.I(new_n8823_), .ZN(new_n8824_));
  AOI21_X1   g08535(.A1(new_n2797_), .A2(new_n4372_), .B(new_n8575_), .ZN(new_n8825_));
  NOR2_X1    g08536(.A1(new_n8245_), .A2(new_n267_), .ZN(new_n8826_));
  NAND2_X1   g08537(.A1(new_n2368_), .A2(new_n3804_), .ZN(new_n8827_));
  AOI21_X1   g08538(.A1(new_n267_), .A2(new_n8245_), .B(new_n8827_), .ZN(new_n8828_));
  NOR2_X1    g08539(.A1(new_n8828_), .A2(new_n8826_), .ZN(new_n8829_));
  INV_X1     g08540(.I(new_n8829_), .ZN(new_n8830_));
  XOR2_X1    g08541(.A1(new_n8825_), .A2(new_n8830_), .Z(new_n8831_));
  NOR2_X1    g08542(.A1(new_n8831_), .A2(new_n8824_), .ZN(new_n8832_));
  INV_X1     g08543(.I(new_n8825_), .ZN(new_n8833_));
  NOR2_X1    g08544(.A1(new_n8833_), .A2(new_n8830_), .ZN(new_n8834_));
  NOR2_X1    g08545(.A1(new_n8825_), .A2(new_n8829_), .ZN(new_n8835_));
  NOR2_X1    g08546(.A1(new_n8834_), .A2(new_n8835_), .ZN(new_n8836_));
  NOR2_X1    g08547(.A1(new_n8836_), .A2(new_n8823_), .ZN(new_n8837_));
  NOR2_X1    g08548(.A1(new_n8837_), .A2(new_n8832_), .ZN(new_n8838_));
  INV_X1     g08549(.I(new_n8838_), .ZN(new_n8839_));
  NAND2_X1   g08550(.A1(new_n7482_), .A2(new_n609_), .ZN(new_n8840_));
  NOR2_X1    g08551(.A1(new_n7482_), .A2(new_n609_), .ZN(new_n8841_));
  NOR2_X1    g08552(.A1(\a[19] ), .A2(\a[42] ), .ZN(new_n8842_));
  AOI21_X1   g08553(.A1(new_n8840_), .A2(new_n8842_), .B(new_n8841_), .ZN(new_n8843_));
  NAND2_X1   g08554(.A1(new_n8458_), .A2(new_n8456_), .ZN(new_n8844_));
  NAND2_X1   g08555(.A1(new_n5592_), .A2(new_n2978_), .ZN(new_n8845_));
  NOR2_X1    g08556(.A1(new_n5592_), .A2(new_n2978_), .ZN(new_n8846_));
  NOR2_X1    g08557(.A1(\a[6] ), .A2(\a[55] ), .ZN(new_n8847_));
  AOI21_X1   g08558(.A1(new_n8845_), .A2(new_n8847_), .B(new_n8846_), .ZN(new_n8848_));
  INV_X1     g08559(.I(new_n8848_), .ZN(new_n8849_));
  XOR2_X1    g08560(.A1(new_n8844_), .A2(new_n8849_), .Z(new_n8850_));
  NAND2_X1   g08561(.A1(new_n8850_), .A2(new_n8843_), .ZN(new_n8851_));
  INV_X1     g08562(.I(new_n8843_), .ZN(new_n8852_));
  NOR2_X1    g08563(.A1(new_n8844_), .A2(new_n8849_), .ZN(new_n8853_));
  NAND2_X1   g08564(.A1(new_n8844_), .A2(new_n8849_), .ZN(new_n8854_));
  INV_X1     g08565(.I(new_n8854_), .ZN(new_n8855_));
  OAI21_X1   g08566(.A1(new_n8855_), .A2(new_n8853_), .B(new_n8852_), .ZN(new_n8856_));
  NAND2_X1   g08567(.A1(new_n8851_), .A2(new_n8856_), .ZN(new_n8857_));
  AOI21_X1   g08568(.A1(new_n654_), .A2(new_n6027_), .B(new_n8431_), .ZN(new_n8858_));
  NOR2_X1    g08569(.A1(\a[13] ), .A2(\a[48] ), .ZN(new_n8859_));
  AOI21_X1   g08570(.A1(new_n8435_), .A2(new_n8859_), .B(new_n8437_), .ZN(new_n8860_));
  NAND2_X1   g08571(.A1(\a[1] ), .A2(\a[61] ), .ZN(new_n8861_));
  XOR2_X1    g08572(.A1(new_n2766_), .A2(new_n8861_), .Z(new_n8862_));
  XNOR2_X1   g08573(.A1(new_n8860_), .A2(new_n8862_), .ZN(new_n8863_));
  INV_X1     g08574(.I(new_n8863_), .ZN(new_n8864_));
  NOR2_X1    g08575(.A1(new_n8860_), .A2(new_n8862_), .ZN(new_n8865_));
  INV_X1     g08576(.I(new_n8865_), .ZN(new_n8866_));
  NAND2_X1   g08577(.A1(new_n8860_), .A2(new_n8862_), .ZN(new_n8867_));
  AOI21_X1   g08578(.A1(new_n8866_), .A2(new_n8867_), .B(new_n8858_), .ZN(new_n8868_));
  AOI21_X1   g08579(.A1(new_n8864_), .A2(new_n8858_), .B(new_n8868_), .ZN(new_n8869_));
  XNOR2_X1   g08580(.A1(new_n8869_), .A2(new_n8857_), .ZN(new_n8870_));
  NAND2_X1   g08581(.A1(new_n8870_), .A2(new_n8839_), .ZN(new_n8871_));
  INV_X1     g08582(.I(new_n8857_), .ZN(new_n8872_));
  NOR2_X1    g08583(.A1(new_n8872_), .A2(new_n8869_), .ZN(new_n8873_));
  NAND2_X1   g08584(.A1(new_n8872_), .A2(new_n8869_), .ZN(new_n8874_));
  INV_X1     g08585(.I(new_n8874_), .ZN(new_n8875_));
  OAI21_X1   g08586(.A1(new_n8875_), .A2(new_n8873_), .B(new_n8838_), .ZN(new_n8876_));
  NAND2_X1   g08587(.A1(new_n8871_), .A2(new_n8876_), .ZN(new_n8877_));
  XOR2_X1    g08588(.A1(new_n8877_), .A2(new_n8822_), .Z(new_n8878_));
  NOR2_X1    g08589(.A1(new_n8810_), .A2(new_n8878_), .ZN(new_n8879_));
  INV_X1     g08590(.I(new_n8810_), .ZN(new_n8880_));
  INV_X1     g08591(.I(new_n8877_), .ZN(new_n8881_));
  NOR2_X1    g08592(.A1(new_n8881_), .A2(new_n8822_), .ZN(new_n8882_));
  INV_X1     g08593(.I(new_n8882_), .ZN(new_n8883_));
  NAND2_X1   g08594(.A1(new_n8881_), .A2(new_n8822_), .ZN(new_n8884_));
  AOI21_X1   g08595(.A1(new_n8883_), .A2(new_n8884_), .B(new_n8880_), .ZN(new_n8885_));
  NOR2_X1    g08596(.A1(new_n8885_), .A2(new_n8879_), .ZN(new_n8886_));
  OAI21_X1   g08597(.A1(new_n8418_), .A2(new_n8482_), .B(new_n8484_), .ZN(new_n8887_));
  INV_X1     g08598(.I(new_n8489_), .ZN(new_n8888_));
  AOI21_X1   g08599(.A1(new_n8888_), .A2(new_n8509_), .B(new_n8507_), .ZN(new_n8889_));
  INV_X1     g08600(.I(new_n8889_), .ZN(new_n8890_));
  INV_X1     g08601(.I(new_n8538_), .ZN(new_n8891_));
  AOI21_X1   g08602(.A1(new_n8525_), .A2(new_n8891_), .B(new_n8540_), .ZN(new_n8892_));
  NOR2_X1    g08603(.A1(new_n8627_), .A2(new_n8609_), .ZN(new_n8893_));
  NOR2_X1    g08604(.A1(new_n8893_), .A2(new_n8628_), .ZN(new_n8894_));
  XOR2_X1    g08605(.A1(new_n8894_), .A2(new_n8892_), .Z(new_n8895_));
  NOR2_X1    g08606(.A1(new_n8894_), .A2(new_n8892_), .ZN(new_n8896_));
  INV_X1     g08607(.I(new_n8896_), .ZN(new_n8897_));
  NAND2_X1   g08608(.A1(new_n8894_), .A2(new_n8892_), .ZN(new_n8898_));
  AOI21_X1   g08609(.A1(new_n8898_), .A2(new_n8897_), .B(new_n8890_), .ZN(new_n8899_));
  AOI21_X1   g08610(.A1(new_n8890_), .A2(new_n8895_), .B(new_n8899_), .ZN(new_n8900_));
  NOR2_X1    g08611(.A1(new_n8887_), .A2(new_n8900_), .ZN(new_n8901_));
  INV_X1     g08612(.I(new_n8901_), .ZN(new_n8902_));
  NAND2_X1   g08613(.A1(new_n8887_), .A2(new_n8900_), .ZN(new_n8903_));
  AOI21_X1   g08614(.A1(new_n8902_), .A2(new_n8903_), .B(new_n8886_), .ZN(new_n8904_));
  INV_X1     g08615(.I(new_n8886_), .ZN(new_n8905_));
  XNOR2_X1   g08616(.A1(new_n8887_), .A2(new_n8900_), .ZN(new_n8906_));
  NOR2_X1    g08617(.A1(new_n8906_), .A2(new_n8905_), .ZN(new_n8907_));
  NOR4_X1    g08618(.A1(new_n8803_), .A2(new_n8808_), .A3(new_n8904_), .A4(new_n8907_), .ZN(new_n8908_));
  NOR2_X1    g08619(.A1(new_n8555_), .A2(new_n8416_), .ZN(new_n8909_));
  NOR2_X1    g08620(.A1(new_n8909_), .A2(new_n8554_), .ZN(new_n8910_));
  NOR2_X1    g08621(.A1(new_n8803_), .A2(new_n8808_), .ZN(new_n8911_));
  NOR2_X1    g08622(.A1(new_n8907_), .A2(new_n8904_), .ZN(new_n8912_));
  NOR2_X1    g08623(.A1(new_n8911_), .A2(new_n8912_), .ZN(new_n8913_));
  NOR2_X1    g08624(.A1(new_n8913_), .A2(new_n8910_), .ZN(new_n8914_));
  NOR2_X1    g08625(.A1(new_n8914_), .A2(new_n8908_), .ZN(new_n8915_));
  INV_X1     g08626(.I(new_n8915_), .ZN(new_n8916_));
  AOI21_X1   g08627(.A1(new_n8666_), .A2(new_n8807_), .B(new_n8805_), .ZN(new_n8917_));
  OAI21_X1   g08628(.A1(new_n8905_), .A2(new_n8901_), .B(new_n8903_), .ZN(new_n8918_));
  INV_X1     g08629(.I(new_n8918_), .ZN(new_n8919_));
  NAND2_X1   g08630(.A1(new_n8880_), .A2(new_n8884_), .ZN(new_n8920_));
  NAND2_X1   g08631(.A1(new_n8920_), .A2(new_n8883_), .ZN(new_n8921_));
  INV_X1     g08632(.I(new_n8921_), .ZN(new_n8922_));
  OAI21_X1   g08633(.A1(new_n8668_), .A2(new_n8715_), .B(new_n8717_), .ZN(new_n8923_));
  NOR2_X1    g08634(.A1(new_n5511_), .A2(new_n6692_), .ZN(new_n8924_));
  INV_X1     g08635(.I(new_n8924_), .ZN(new_n8925_));
  NOR2_X1    g08636(.A1(new_n8925_), .A2(new_n2066_), .ZN(new_n8926_));
  NOR2_X1    g08637(.A1(new_n800_), .A2(new_n6694_), .ZN(new_n8927_));
  NAND4_X1   g08638(.A1(new_n8926_), .A2(\a[10] ), .A3(new_n8927_), .A4(\a[47] ), .ZN(new_n8928_));
  AOI21_X1   g08639(.A1(new_n8928_), .A2(new_n8056_), .B(new_n796_), .ZN(new_n8929_));
  NOR3_X1    g08640(.A1(new_n8929_), .A2(new_n461_), .A3(new_n6694_), .ZN(new_n8930_));
  NOR3_X1    g08641(.A1(new_n8929_), .A2(new_n2252_), .A3(new_n8924_), .ZN(new_n8931_));
  NOR2_X1    g08642(.A1(new_n8930_), .A2(new_n8931_), .ZN(new_n8932_));
  NOR2_X1    g08643(.A1(new_n5175_), .A2(new_n6945_), .ZN(new_n8933_));
  INV_X1     g08644(.I(new_n8933_), .ZN(new_n8934_));
  NOR2_X1    g08645(.A1(new_n8934_), .A2(new_n1965_), .ZN(new_n8935_));
  NOR2_X1    g08646(.A1(new_n8934_), .A2(new_n1965_), .ZN(new_n8939_));
  INV_X1     g08647(.I(new_n8939_), .ZN(new_n8940_));
  INV_X1     g08648(.I(new_n6779_), .ZN(new_n8941_));
  NOR2_X1    g08649(.A1(new_n8941_), .A2(new_n1150_), .ZN(new_n8942_));
  NOR2_X1    g08650(.A1(new_n8941_), .A2(new_n1150_), .ZN(new_n8946_));
  INV_X1     g08651(.I(new_n8946_), .ZN(new_n8947_));
  NOR2_X1    g08652(.A1(new_n8940_), .A2(new_n8947_), .ZN(new_n8948_));
  NOR2_X1    g08653(.A1(new_n8939_), .A2(new_n8946_), .ZN(new_n8949_));
  OAI21_X1   g08654(.A1(new_n8948_), .A2(new_n8949_), .B(new_n8932_), .ZN(new_n8950_));
  XNOR2_X1   g08655(.A1(new_n8939_), .A2(new_n8946_), .ZN(new_n8951_));
  OAI21_X1   g08656(.A1(new_n8932_), .A2(new_n8951_), .B(new_n8950_), .ZN(new_n8952_));
  INV_X1     g08657(.I(new_n8755_), .ZN(new_n8953_));
  INV_X1     g08658(.I(new_n2060_), .ZN(new_n8954_));
  NOR2_X1    g08659(.A1(new_n4770_), .A2(new_n6999_), .ZN(new_n8955_));
  INV_X1     g08660(.I(new_n8955_), .ZN(new_n8956_));
  NOR2_X1    g08661(.A1(new_n8954_), .A2(new_n8956_), .ZN(new_n8957_));
  NOR3_X1    g08662(.A1(new_n1961_), .A2(new_n4770_), .A3(new_n7216_), .ZN(new_n8958_));
  NAND2_X1   g08663(.A1(new_n8957_), .A2(new_n8958_), .ZN(new_n8959_));
  AOI21_X1   g08664(.A1(new_n8959_), .A2(new_n8953_), .B(new_n392_), .ZN(new_n8960_));
  NAND2_X1   g08665(.A1(\a[7] ), .A2(\a[56] ), .ZN(new_n8961_));
  NOR2_X1    g08666(.A1(new_n8960_), .A2(new_n8957_), .ZN(new_n8962_));
  INV_X1     g08667(.I(new_n8962_), .ZN(new_n8963_));
  NAND2_X1   g08668(.A1(new_n8954_), .A2(new_n8956_), .ZN(new_n8964_));
  OAI22_X1   g08669(.A1(new_n8963_), .A2(new_n8964_), .B1(new_n8960_), .B2(new_n8961_), .ZN(new_n8965_));
  NOR2_X1    g08670(.A1(new_n1215_), .A2(new_n4501_), .ZN(new_n8966_));
  INV_X1     g08671(.I(new_n8966_), .ZN(new_n8967_));
  NOR2_X1    g08672(.A1(new_n2368_), .A2(new_n4240_), .ZN(new_n8968_));
  INV_X1     g08673(.I(new_n8968_), .ZN(new_n8969_));
  NOR2_X1    g08674(.A1(new_n8967_), .A2(new_n8969_), .ZN(new_n8970_));
  XOR2_X1    g08675(.A1(new_n8970_), .A2(new_n242_), .Z(new_n8971_));
  XOR2_X1    g08676(.A1(new_n8971_), .A2(\a[57] ), .Z(new_n8972_));
  NOR2_X1    g08677(.A1(new_n2461_), .A2(new_n2868_), .ZN(new_n8973_));
  INV_X1     g08678(.I(new_n8973_), .ZN(new_n8974_));
  NOR2_X1    g08679(.A1(new_n8974_), .A2(new_n4184_), .ZN(new_n8975_));
  XOR2_X1    g08680(.A1(new_n8975_), .A2(new_n650_), .Z(new_n8976_));
  XOR2_X1    g08681(.A1(new_n8976_), .A2(\a[49] ), .Z(new_n8977_));
  NOR2_X1    g08682(.A1(new_n8972_), .A2(new_n8977_), .ZN(new_n8978_));
  AND2_X2    g08683(.A1(new_n8972_), .A2(new_n8977_), .Z(new_n8979_));
  NOR2_X1    g08684(.A1(new_n8979_), .A2(new_n8978_), .ZN(new_n8980_));
  NOR2_X1    g08685(.A1(new_n8980_), .A2(new_n8965_), .ZN(new_n8981_));
  INV_X1     g08686(.I(new_n8965_), .ZN(new_n8982_));
  XNOR2_X1   g08687(.A1(new_n8972_), .A2(new_n8977_), .ZN(new_n8983_));
  NOR2_X1    g08688(.A1(new_n8983_), .A2(new_n8982_), .ZN(new_n8984_));
  NOR2_X1    g08689(.A1(new_n8981_), .A2(new_n8984_), .ZN(new_n8985_));
  NOR3_X1    g08690(.A1(new_n868_), .A2(new_n5511_), .A3(new_n6260_), .ZN(new_n8986_));
  NOR2_X1    g08691(.A1(new_n1021_), .A2(new_n8749_), .ZN(new_n8987_));
  NOR2_X1    g08692(.A1(new_n8986_), .A2(new_n8987_), .ZN(new_n8988_));
  INV_X1     g08693(.I(new_n8455_), .ZN(new_n8989_));
  INV_X1     g08694(.I(\a[60] ), .ZN(new_n8990_));
  NOR2_X1    g08695(.A1(new_n8990_), .A2(new_n8453_), .ZN(new_n8991_));
  INV_X1     g08696(.I(new_n8991_), .ZN(new_n8992_));
  NOR2_X1    g08697(.A1(new_n8989_), .A2(new_n8992_), .ZN(new_n8993_));
  NOR2_X1    g08698(.A1(new_n8993_), .A2(new_n1271_), .ZN(new_n8994_));
  INV_X1     g08699(.I(new_n8994_), .ZN(new_n8995_));
  NOR2_X1    g08700(.A1(new_n8085_), .A2(new_n8990_), .ZN(new_n8996_));
  NOR2_X1    g08701(.A1(new_n201_), .A2(new_n8453_), .ZN(new_n8997_));
  INV_X1     g08702(.I(new_n8997_), .ZN(new_n8998_));
  NOR4_X1    g08703(.A1(new_n8995_), .A2(new_n267_), .A3(new_n8996_), .A4(new_n8998_), .ZN(new_n8999_));
  NAND2_X1   g08704(.A1(new_n5350_), .A2(new_n4538_), .ZN(new_n9000_));
  NOR2_X1    g08705(.A1(new_n353_), .A2(new_n7647_), .ZN(new_n9001_));
  XOR2_X1    g08706(.A1(new_n9000_), .A2(new_n9001_), .Z(new_n9002_));
  XNOR2_X1   g08707(.A1(new_n8999_), .A2(new_n9002_), .ZN(new_n9003_));
  INV_X1     g08708(.I(new_n8999_), .ZN(new_n9004_));
  NOR2_X1    g08709(.A1(new_n9004_), .A2(new_n9002_), .ZN(new_n9005_));
  INV_X1     g08710(.I(new_n9005_), .ZN(new_n9006_));
  NAND2_X1   g08711(.A1(new_n9004_), .A2(new_n9002_), .ZN(new_n9007_));
  AOI21_X1   g08712(.A1(new_n9006_), .A2(new_n9007_), .B(new_n8988_), .ZN(new_n9008_));
  AOI21_X1   g08713(.A1(new_n8988_), .A2(new_n9003_), .B(new_n9008_), .ZN(new_n9009_));
  XNOR2_X1   g08714(.A1(new_n8985_), .A2(new_n9009_), .ZN(new_n9010_));
  INV_X1     g08715(.I(new_n8985_), .ZN(new_n9011_));
  NOR2_X1    g08716(.A1(new_n9011_), .A2(new_n9009_), .ZN(new_n9012_));
  INV_X1     g08717(.I(new_n9012_), .ZN(new_n9013_));
  NAND2_X1   g08718(.A1(new_n9011_), .A2(new_n9009_), .ZN(new_n9014_));
  AOI21_X1   g08719(.A1(new_n9013_), .A2(new_n9014_), .B(new_n8952_), .ZN(new_n9015_));
  AOI21_X1   g08720(.A1(new_n8952_), .A2(new_n9010_), .B(new_n9015_), .ZN(new_n9016_));
  NOR2_X1    g08721(.A1(new_n9016_), .A2(new_n8923_), .ZN(new_n9017_));
  INV_X1     g08722(.I(new_n9017_), .ZN(new_n9018_));
  NAND2_X1   g08723(.A1(new_n9016_), .A2(new_n8923_), .ZN(new_n9019_));
  AOI21_X1   g08724(.A1(new_n9018_), .A2(new_n9019_), .B(new_n8922_), .ZN(new_n9020_));
  XNOR2_X1   g08725(.A1(new_n9016_), .A2(new_n8923_), .ZN(new_n9021_));
  NOR2_X1    g08726(.A1(new_n8921_), .A2(new_n9021_), .ZN(new_n9022_));
  NOR2_X1    g08727(.A1(new_n9020_), .A2(new_n9022_), .ZN(new_n9023_));
  INV_X1     g08728(.I(new_n9023_), .ZN(new_n9024_));
  AOI21_X1   g08729(.A1(new_n8890_), .A2(new_n8898_), .B(new_n8896_), .ZN(new_n9025_));
  AOI21_X1   g08730(.A1(new_n8699_), .A2(new_n8707_), .B(new_n8706_), .ZN(new_n9026_));
  AOI21_X1   g08731(.A1(new_n8743_), .A2(new_n8733_), .B(new_n8740_), .ZN(new_n9027_));
  NOR2_X1    g08732(.A1(new_n3849_), .A2(new_n8861_), .ZN(new_n9028_));
  INV_X1     g08733(.I(\a[62] ), .ZN(new_n9029_));
  OAI21_X1   g08734(.A1(new_n194_), .A2(new_n9029_), .B(new_n2765_), .ZN(new_n9030_));
  NOR2_X1    g08735(.A1(new_n2765_), .A2(new_n9029_), .ZN(new_n9031_));
  NAND2_X1   g08736(.A1(new_n9031_), .A2(\a[1] ), .ZN(new_n9032_));
  NAND2_X1   g08737(.A1(new_n9032_), .A2(new_n9030_), .ZN(new_n9033_));
  NAND2_X1   g08738(.A1(new_n9033_), .A2(new_n9028_), .ZN(new_n9034_));
  XOR2_X1    g08739(.A1(new_n9034_), .A2(\a[0] ), .Z(new_n9035_));
  XOR2_X1    g08740(.A1(new_n9035_), .A2(\a[63] ), .Z(new_n9036_));
  AOI22_X1   g08741(.A1(new_n2277_), .A2(new_n5601_), .B1(new_n5339_), .B2(new_n4515_), .ZN(new_n9037_));
  INV_X1     g08742(.I(new_n9037_), .ZN(new_n9038_));
  NAND4_X1   g08743(.A1(new_n2753_), .A2(new_n4706_), .A3(\a[24] ), .A4(\a[39] ), .ZN(new_n9039_));
  NOR2_X1    g08744(.A1(new_n9038_), .A2(new_n9039_), .ZN(new_n9040_));
  INV_X1     g08745(.I(new_n9040_), .ZN(new_n9041_));
  NOR2_X1    g08746(.A1(new_n3174_), .A2(new_n2692_), .ZN(new_n9042_));
  NOR2_X1    g08747(.A1(new_n4729_), .A2(new_n9042_), .ZN(new_n9043_));
  NOR4_X1    g08748(.A1(new_n3487_), .A2(new_n2690_), .A3(new_n2098_), .A4(new_n3393_), .ZN(new_n9044_));
  NAND2_X1   g08749(.A1(new_n9043_), .A2(new_n9044_), .ZN(new_n9045_));
  NOR2_X1    g08750(.A1(new_n9041_), .A2(new_n9045_), .ZN(new_n9046_));
  AOI21_X1   g08751(.A1(new_n9043_), .A2(new_n9044_), .B(new_n9040_), .ZN(new_n9047_));
  NOR2_X1    g08752(.A1(new_n9046_), .A2(new_n9047_), .ZN(new_n9048_));
  NOR2_X1    g08753(.A1(new_n9036_), .A2(new_n9048_), .ZN(new_n9049_));
  INV_X1     g08754(.I(new_n9036_), .ZN(new_n9050_));
  XOR2_X1    g08755(.A1(new_n9045_), .A2(new_n9040_), .Z(new_n9051_));
  NOR2_X1    g08756(.A1(new_n9050_), .A2(new_n9051_), .ZN(new_n9052_));
  NOR2_X1    g08757(.A1(new_n9052_), .A2(new_n9049_), .ZN(new_n9053_));
  NOR2_X1    g08758(.A1(new_n9053_), .A2(new_n9027_), .ZN(new_n9054_));
  INV_X1     g08759(.I(new_n9054_), .ZN(new_n9055_));
  NAND2_X1   g08760(.A1(new_n9053_), .A2(new_n9027_), .ZN(new_n9056_));
  AOI21_X1   g08761(.A1(new_n9055_), .A2(new_n9056_), .B(new_n9026_), .ZN(new_n9057_));
  INV_X1     g08762(.I(new_n9026_), .ZN(new_n9058_));
  XNOR2_X1   g08763(.A1(new_n9053_), .A2(new_n9027_), .ZN(new_n9059_));
  NOR2_X1    g08764(.A1(new_n9059_), .A2(new_n9058_), .ZN(new_n9060_));
  NOR2_X1    g08765(.A1(new_n9060_), .A2(new_n9057_), .ZN(new_n9061_));
  AOI21_X1   g08766(.A1(new_n8751_), .A2(new_n8760_), .B(new_n8759_), .ZN(new_n9062_));
  AOI21_X1   g08767(.A1(new_n2690_), .A2(new_n4372_), .B(new_n8775_), .ZN(new_n9063_));
  XOR2_X1    g08768(.A1(new_n8730_), .A2(new_n9063_), .Z(new_n9064_));
  NOR3_X1    g08769(.A1(new_n9064_), .A2(new_n8769_), .A3(new_n8770_), .ZN(new_n9065_));
  NOR2_X1    g08770(.A1(new_n8769_), .A2(new_n8770_), .ZN(new_n9066_));
  INV_X1     g08771(.I(new_n9063_), .ZN(new_n9067_));
  NOR2_X1    g08772(.A1(new_n9067_), .A2(new_n8730_), .ZN(new_n9068_));
  NOR2_X1    g08773(.A1(new_n8731_), .A2(new_n9063_), .ZN(new_n9069_));
  NOR2_X1    g08774(.A1(new_n9069_), .A2(new_n9068_), .ZN(new_n9070_));
  NOR2_X1    g08775(.A1(new_n9070_), .A2(new_n9066_), .ZN(new_n9071_));
  NOR2_X1    g08776(.A1(new_n9071_), .A2(new_n9065_), .ZN(new_n9072_));
  NOR2_X1    g08777(.A1(new_n8783_), .A2(new_n8773_), .ZN(new_n9073_));
  NOR2_X1    g08778(.A1(new_n9073_), .A2(new_n8782_), .ZN(new_n9074_));
  XOR2_X1    g08779(.A1(new_n9072_), .A2(new_n9074_), .Z(new_n9075_));
  NOR2_X1    g08780(.A1(new_n9075_), .A2(new_n9062_), .ZN(new_n9076_));
  INV_X1     g08781(.I(new_n9062_), .ZN(new_n9077_));
  INV_X1     g08782(.I(new_n9072_), .ZN(new_n9078_));
  NOR2_X1    g08783(.A1(new_n9078_), .A2(new_n9074_), .ZN(new_n9079_));
  INV_X1     g08784(.I(new_n9079_), .ZN(new_n9080_));
  NAND2_X1   g08785(.A1(new_n9078_), .A2(new_n9074_), .ZN(new_n9081_));
  AOI21_X1   g08786(.A1(new_n9080_), .A2(new_n9081_), .B(new_n9077_), .ZN(new_n9082_));
  NOR2_X1    g08787(.A1(new_n9082_), .A2(new_n9076_), .ZN(new_n9083_));
  XOR2_X1    g08788(.A1(new_n9061_), .A2(new_n9083_), .Z(new_n9084_));
  NOR2_X1    g08789(.A1(new_n9084_), .A2(new_n9025_), .ZN(new_n9085_));
  INV_X1     g08790(.I(new_n9025_), .ZN(new_n9086_));
  INV_X1     g08791(.I(new_n9083_), .ZN(new_n9087_));
  NAND2_X1   g08792(.A1(new_n9061_), .A2(new_n9087_), .ZN(new_n9088_));
  NOR2_X1    g08793(.A1(new_n9061_), .A2(new_n9087_), .ZN(new_n9089_));
  INV_X1     g08794(.I(new_n9089_), .ZN(new_n9090_));
  AOI21_X1   g08795(.A1(new_n9090_), .A2(new_n9088_), .B(new_n9086_), .ZN(new_n9091_));
  NOR2_X1    g08796(.A1(new_n9085_), .A2(new_n9091_), .ZN(new_n9092_));
  NOR2_X1    g08797(.A1(new_n9024_), .A2(new_n9092_), .ZN(new_n9093_));
  INV_X1     g08798(.I(new_n9093_), .ZN(new_n9094_));
  NAND2_X1   g08799(.A1(new_n9024_), .A2(new_n9092_), .ZN(new_n9095_));
  AOI21_X1   g08800(.A1(new_n9094_), .A2(new_n9095_), .B(new_n8919_), .ZN(new_n9096_));
  XOR2_X1    g08801(.A1(new_n9023_), .A2(new_n9092_), .Z(new_n9097_));
  NOR2_X1    g08802(.A1(new_n9097_), .A2(new_n8918_), .ZN(new_n9098_));
  NOR2_X1    g08803(.A1(new_n9096_), .A2(new_n9098_), .ZN(new_n9099_));
  OAI21_X1   g08804(.A1(new_n8721_), .A2(new_n8796_), .B(new_n8798_), .ZN(new_n9100_));
  AOI21_X1   g08805(.A1(new_n8691_), .A2(new_n8695_), .B(new_n8693_), .ZN(new_n9101_));
  OAI21_X1   g08806(.A1(new_n8839_), .A2(new_n8873_), .B(new_n8874_), .ZN(new_n9102_));
  NOR2_X1    g08807(.A1(new_n8820_), .A2(new_n8812_), .ZN(new_n9103_));
  NOR2_X1    g08808(.A1(new_n9103_), .A2(new_n8818_), .ZN(new_n9104_));
  XOR2_X1    g08809(.A1(new_n9104_), .A2(new_n9102_), .Z(new_n9105_));
  NOR2_X1    g08810(.A1(new_n9105_), .A2(new_n9101_), .ZN(new_n9106_));
  INV_X1     g08811(.I(new_n9101_), .ZN(new_n9107_));
  INV_X1     g08812(.I(new_n9102_), .ZN(new_n9108_));
  NOR2_X1    g08813(.A1(new_n9104_), .A2(new_n9108_), .ZN(new_n9109_));
  INV_X1     g08814(.I(new_n9109_), .ZN(new_n9110_));
  NAND2_X1   g08815(.A1(new_n9104_), .A2(new_n9108_), .ZN(new_n9111_));
  AOI21_X1   g08816(.A1(new_n9110_), .A2(new_n9111_), .B(new_n9107_), .ZN(new_n9112_));
  NOR2_X1    g08817(.A1(new_n9106_), .A2(new_n9112_), .ZN(new_n9113_));
  INV_X1     g08818(.I(new_n8683_), .ZN(new_n9114_));
  AOI21_X1   g08819(.A1(new_n9114_), .A2(new_n8671_), .B(new_n8682_), .ZN(new_n9115_));
  NOR2_X1    g08820(.A1(new_n8835_), .A2(new_n8824_), .ZN(new_n9116_));
  NOR2_X1    g08821(.A1(new_n9116_), .A2(new_n8834_), .ZN(new_n9117_));
  NAND2_X1   g08822(.A1(new_n8866_), .A2(new_n8858_), .ZN(new_n9118_));
  NAND2_X1   g08823(.A1(new_n9118_), .A2(new_n8867_), .ZN(new_n9119_));
  XOR2_X1    g08824(.A1(new_n9119_), .A2(new_n9117_), .Z(new_n9120_));
  NOR2_X1    g08825(.A1(new_n9120_), .A2(new_n9115_), .ZN(new_n9121_));
  INV_X1     g08826(.I(new_n9115_), .ZN(new_n9122_));
  INV_X1     g08827(.I(new_n9119_), .ZN(new_n9123_));
  NOR2_X1    g08828(.A1(new_n9123_), .A2(new_n9117_), .ZN(new_n9124_));
  INV_X1     g08829(.I(new_n9124_), .ZN(new_n9125_));
  NAND2_X1   g08830(.A1(new_n9123_), .A2(new_n9117_), .ZN(new_n9126_));
  AOI21_X1   g08831(.A1(new_n9125_), .A2(new_n9126_), .B(new_n9122_), .ZN(new_n9127_));
  NOR2_X1    g08832(.A1(new_n9127_), .A2(new_n9121_), .ZN(new_n9128_));
  INV_X1     g08833(.I(new_n8792_), .ZN(new_n9129_));
  AOI21_X1   g08834(.A1(new_n8748_), .A2(new_n9129_), .B(new_n8791_), .ZN(new_n9130_));
  INV_X1     g08835(.I(new_n9130_), .ZN(new_n9131_));
  AOI21_X1   g08836(.A1(new_n2543_), .A2(new_n5339_), .B(new_n8779_), .ZN(new_n9132_));
  INV_X1     g08837(.I(new_n9132_), .ZN(new_n9133_));
  AOI21_X1   g08838(.A1(new_n787_), .A2(new_n6028_), .B(new_n8752_), .ZN(new_n9134_));
  NAND2_X1   g08839(.A1(new_n8755_), .A2(new_n479_), .ZN(new_n9135_));
  NOR2_X1    g08840(.A1(new_n8755_), .A2(new_n479_), .ZN(new_n9136_));
  NOR2_X1    g08841(.A1(\a[20] ), .A2(\a[42] ), .ZN(new_n9137_));
  AOI21_X1   g08842(.A1(new_n9135_), .A2(new_n9137_), .B(new_n9136_), .ZN(new_n9138_));
  XNOR2_X1   g08843(.A1(new_n9134_), .A2(new_n9138_), .ZN(new_n9139_));
  NOR2_X1    g08844(.A1(new_n9139_), .A2(new_n9133_), .ZN(new_n9140_));
  INV_X1     g08845(.I(new_n9134_), .ZN(new_n9141_));
  INV_X1     g08846(.I(new_n9138_), .ZN(new_n9142_));
  NOR2_X1    g08847(.A1(new_n9141_), .A2(new_n9142_), .ZN(new_n9143_));
  NOR2_X1    g08848(.A1(new_n9134_), .A2(new_n9138_), .ZN(new_n9144_));
  NOR2_X1    g08849(.A1(new_n9143_), .A2(new_n9144_), .ZN(new_n9145_));
  NOR2_X1    g08850(.A1(new_n9145_), .A2(new_n9132_), .ZN(new_n9146_));
  NOR2_X1    g08851(.A1(new_n9146_), .A2(new_n9140_), .ZN(new_n9147_));
  AOI21_X1   g08852(.A1(new_n229_), .A2(new_n8245_), .B(new_n8679_), .ZN(new_n9148_));
  INV_X1     g08853(.I(new_n9148_), .ZN(new_n9149_));
  NOR2_X1    g08854(.A1(\a[21] ), .A2(\a[41] ), .ZN(new_n9150_));
  OAI21_X1   g08855(.A1(new_n2753_), .A2(new_n3839_), .B(new_n9150_), .ZN(new_n9151_));
  OAI21_X1   g08856(.A1(new_n2752_), .A2(new_n3838_), .B(new_n9151_), .ZN(new_n9152_));
  NOR2_X1    g08857(.A1(new_n8990_), .A2(new_n9029_), .ZN(new_n9153_));
  NOR3_X1    g08858(.A1(new_n194_), .A2(new_n2655_), .A3(new_n8990_), .ZN(new_n9154_));
  AOI21_X1   g08859(.A1(new_n9154_), .A2(new_n218_), .B(new_n9153_), .ZN(new_n9155_));
  XNOR2_X1   g08860(.A1(new_n9152_), .A2(new_n9155_), .ZN(new_n9156_));
  NOR2_X1    g08861(.A1(new_n9156_), .A2(new_n9149_), .ZN(new_n9157_));
  NOR2_X1    g08862(.A1(new_n9152_), .A2(new_n9155_), .ZN(new_n9158_));
  INV_X1     g08863(.I(new_n9158_), .ZN(new_n9159_));
  NAND2_X1   g08864(.A1(new_n9152_), .A2(new_n9155_), .ZN(new_n9160_));
  AOI21_X1   g08865(.A1(new_n9159_), .A2(new_n9160_), .B(new_n9148_), .ZN(new_n9161_));
  NOR2_X1    g08866(.A1(new_n9157_), .A2(new_n9161_), .ZN(new_n9162_));
  INV_X1     g08867(.I(new_n9162_), .ZN(new_n9163_));
  AOI21_X1   g08868(.A1(new_n8843_), .A2(new_n8854_), .B(new_n8853_), .ZN(new_n9164_));
  NOR2_X1    g08869(.A1(new_n9163_), .A2(new_n9164_), .ZN(new_n9165_));
  INV_X1     g08870(.I(new_n9164_), .ZN(new_n9166_));
  NOR2_X1    g08871(.A1(new_n9162_), .A2(new_n9166_), .ZN(new_n9167_));
  NOR2_X1    g08872(.A1(new_n9165_), .A2(new_n9167_), .ZN(new_n9168_));
  NOR2_X1    g08873(.A1(new_n9168_), .A2(new_n9147_), .ZN(new_n9169_));
  XOR2_X1    g08874(.A1(new_n9162_), .A2(new_n9164_), .Z(new_n9170_));
  NOR3_X1    g08875(.A1(new_n9170_), .A2(new_n9140_), .A3(new_n9146_), .ZN(new_n9171_));
  NOR2_X1    g08876(.A1(new_n9169_), .A2(new_n9171_), .ZN(new_n9172_));
  NOR2_X1    g08877(.A1(new_n9172_), .A2(new_n9131_), .ZN(new_n9173_));
  INV_X1     g08878(.I(new_n9172_), .ZN(new_n9174_));
  NOR2_X1    g08879(.A1(new_n9174_), .A2(new_n9130_), .ZN(new_n9175_));
  NOR2_X1    g08880(.A1(new_n9175_), .A2(new_n9173_), .ZN(new_n9176_));
  NOR2_X1    g08881(.A1(new_n9176_), .A2(new_n9128_), .ZN(new_n9177_));
  XOR2_X1    g08882(.A1(new_n9172_), .A2(new_n9130_), .Z(new_n9178_));
  INV_X1     g08883(.I(new_n9178_), .ZN(new_n9179_));
  AOI21_X1   g08884(.A1(new_n9128_), .A2(new_n9179_), .B(new_n9177_), .ZN(new_n9180_));
  NOR2_X1    g08885(.A1(new_n9180_), .A2(new_n9113_), .ZN(new_n9181_));
  NAND2_X1   g08886(.A1(new_n9180_), .A2(new_n9113_), .ZN(new_n9182_));
  INV_X1     g08887(.I(new_n9182_), .ZN(new_n9183_));
  OAI21_X1   g08888(.A1(new_n9181_), .A2(new_n9183_), .B(new_n9100_), .ZN(new_n9184_));
  XNOR2_X1   g08889(.A1(new_n9180_), .A2(new_n9113_), .ZN(new_n9185_));
  OAI21_X1   g08890(.A1(new_n9100_), .A2(new_n9185_), .B(new_n9184_), .ZN(new_n9186_));
  XOR2_X1    g08891(.A1(new_n9099_), .A2(new_n9186_), .Z(new_n9187_));
  NOR2_X1    g08892(.A1(new_n9187_), .A2(new_n8917_), .ZN(new_n9188_));
  INV_X1     g08893(.I(new_n8917_), .ZN(new_n9189_));
  INV_X1     g08894(.I(new_n9186_), .ZN(new_n9190_));
  NOR2_X1    g08895(.A1(new_n9099_), .A2(new_n9190_), .ZN(new_n9191_));
  INV_X1     g08896(.I(new_n9191_), .ZN(new_n9192_));
  NAND2_X1   g08897(.A1(new_n9099_), .A2(new_n9190_), .ZN(new_n9193_));
  AOI21_X1   g08898(.A1(new_n9192_), .A2(new_n9193_), .B(new_n9189_), .ZN(new_n9194_));
  NOR2_X1    g08899(.A1(new_n9188_), .A2(new_n9194_), .ZN(new_n9195_));
  XOR2_X1    g08900(.A1(new_n9195_), .A2(new_n8916_), .Z(new_n9196_));
  NAND2_X1   g08901(.A1(\asquared[63] ), .A2(new_n9196_), .ZN(new_n9197_));
  NOR2_X1    g08902(.A1(new_n9195_), .A2(new_n8916_), .ZN(new_n9198_));
  INV_X1     g08903(.I(new_n9195_), .ZN(new_n9199_));
  NOR2_X1    g08904(.A1(new_n9199_), .A2(new_n8915_), .ZN(new_n9200_));
  NOR2_X1    g08905(.A1(new_n9200_), .A2(new_n9198_), .ZN(new_n9201_));
  OAI21_X1   g08906(.A1(\asquared[63] ), .A2(new_n9201_), .B(new_n9197_), .ZN(\asquared[64] ));
  INV_X1     g08907(.I(new_n9198_), .ZN(new_n9203_));
  AOI21_X1   g08908(.A1(\asquared[63] ), .A2(new_n9203_), .B(new_n9200_), .ZN(new_n9204_));
  OAI21_X1   g08909(.A1(new_n8919_), .A2(new_n9093_), .B(new_n9095_), .ZN(new_n9205_));
  INV_X1     g08910(.I(new_n9205_), .ZN(new_n9206_));
  OAI21_X1   g08911(.A1(new_n8922_), .A2(new_n9017_), .B(new_n9019_), .ZN(new_n9207_));
  INV_X1     g08912(.I(new_n9207_), .ZN(new_n9208_));
  AOI21_X1   g08913(.A1(new_n9086_), .A2(new_n9088_), .B(new_n9089_), .ZN(new_n9209_));
  INV_X1     g08914(.I(new_n9209_), .ZN(new_n9210_));
  INV_X1     g08915(.I(new_n8952_), .ZN(new_n9211_));
  OAI21_X1   g08916(.A1(new_n9211_), .A2(new_n9012_), .B(new_n9014_), .ZN(new_n9212_));
  INV_X1     g08917(.I(new_n9212_), .ZN(new_n9213_));
  NAND2_X1   g08918(.A1(new_n9056_), .A2(new_n9058_), .ZN(new_n9214_));
  NAND2_X1   g08919(.A1(new_n9214_), .A2(new_n9055_), .ZN(new_n9215_));
  AOI21_X1   g08920(.A1(new_n1441_), .A2(new_n5488_), .B(new_n8935_), .ZN(new_n9216_));
  INV_X1     g08921(.I(new_n9216_), .ZN(new_n9217_));
  AOI21_X1   g08922(.A1(new_n2690_), .A2(new_n3487_), .B(new_n9043_), .ZN(new_n9218_));
  NOR2_X1    g08923(.A1(new_n242_), .A2(new_n7727_), .ZN(new_n9219_));
  OAI21_X1   g08924(.A1(new_n8966_), .A2(new_n8968_), .B(new_n9219_), .ZN(new_n9220_));
  OAI21_X1   g08925(.A1(new_n8967_), .A2(new_n8969_), .B(new_n9220_), .ZN(new_n9221_));
  INV_X1     g08926(.I(new_n9221_), .ZN(new_n9222_));
  XOR2_X1    g08927(.A1(new_n9218_), .A2(new_n9222_), .Z(new_n9223_));
  NOR2_X1    g08928(.A1(new_n9223_), .A2(new_n9217_), .ZN(new_n9224_));
  INV_X1     g08929(.I(new_n9218_), .ZN(new_n9225_));
  NOR2_X1    g08930(.A1(new_n9225_), .A2(new_n9222_), .ZN(new_n9226_));
  NOR2_X1    g08931(.A1(new_n9218_), .A2(new_n9221_), .ZN(new_n9227_));
  NOR2_X1    g08932(.A1(new_n9226_), .A2(new_n9227_), .ZN(new_n9228_));
  NOR2_X1    g08933(.A1(new_n9228_), .A2(new_n9216_), .ZN(new_n9229_));
  NOR2_X1    g08934(.A1(new_n9229_), .A2(new_n9224_), .ZN(new_n9230_));
  INV_X1     g08935(.I(new_n9230_), .ZN(new_n9231_));
  AOI21_X1   g08936(.A1(new_n267_), .A2(new_n8996_), .B(new_n8994_), .ZN(new_n9232_));
  NOR2_X1    g08937(.A1(new_n5350_), .A2(new_n4538_), .ZN(new_n9233_));
  NAND2_X1   g08938(.A1(new_n353_), .A2(new_n7647_), .ZN(new_n9234_));
  AOI21_X1   g08939(.A1(new_n4538_), .A2(new_n5350_), .B(new_n9234_), .ZN(new_n9235_));
  NOR2_X1    g08940(.A1(new_n9235_), .A2(new_n9233_), .ZN(new_n9236_));
  INV_X1     g08941(.I(new_n9236_), .ZN(new_n9237_));
  XOR2_X1    g08942(.A1(new_n9232_), .A2(new_n9237_), .Z(new_n9238_));
  NOR2_X1    g08943(.A1(new_n9238_), .A2(new_n8963_), .ZN(new_n9239_));
  INV_X1     g08944(.I(new_n9232_), .ZN(new_n9240_));
  NOR2_X1    g08945(.A1(new_n9240_), .A2(new_n9237_), .ZN(new_n9241_));
  NOR2_X1    g08946(.A1(new_n9232_), .A2(new_n9236_), .ZN(new_n9242_));
  NOR2_X1    g08947(.A1(new_n9241_), .A2(new_n9242_), .ZN(new_n9243_));
  NOR2_X1    g08948(.A1(new_n9243_), .A2(new_n8962_), .ZN(new_n9244_));
  INV_X1     g08949(.I(new_n9047_), .ZN(new_n9245_));
  AOI21_X1   g08950(.A1(new_n9050_), .A2(new_n9245_), .B(new_n9046_), .ZN(new_n9246_));
  NOR3_X1    g08951(.A1(new_n9246_), .A2(new_n9239_), .A3(new_n9244_), .ZN(new_n9247_));
  NOR2_X1    g08952(.A1(new_n9244_), .A2(new_n9239_), .ZN(new_n9248_));
  INV_X1     g08953(.I(new_n9246_), .ZN(new_n9249_));
  NOR2_X1    g08954(.A1(new_n9249_), .A2(new_n9248_), .ZN(new_n9250_));
  OAI21_X1   g08955(.A1(new_n9250_), .A2(new_n9247_), .B(new_n9231_), .ZN(new_n9251_));
  XNOR2_X1   g08956(.A1(new_n9246_), .A2(new_n9248_), .ZN(new_n9252_));
  NAND2_X1   g08957(.A1(new_n9252_), .A2(new_n9230_), .ZN(new_n9253_));
  NAND2_X1   g08958(.A1(new_n9253_), .A2(new_n9251_), .ZN(new_n9254_));
  XOR2_X1    g08959(.A1(new_n9254_), .A2(new_n9215_), .Z(new_n9255_));
  NOR2_X1    g08960(.A1(new_n9255_), .A2(new_n9213_), .ZN(new_n9256_));
  INV_X1     g08961(.I(new_n9254_), .ZN(new_n9257_));
  NOR2_X1    g08962(.A1(new_n9257_), .A2(new_n9215_), .ZN(new_n9258_));
  INV_X1     g08963(.I(new_n9258_), .ZN(new_n9259_));
  NAND2_X1   g08964(.A1(new_n9257_), .A2(new_n9215_), .ZN(new_n9260_));
  AOI21_X1   g08965(.A1(new_n9259_), .A2(new_n9260_), .B(new_n9212_), .ZN(new_n9261_));
  NOR2_X1    g08966(.A1(new_n9261_), .A2(new_n9256_), .ZN(new_n9262_));
  NOR2_X1    g08967(.A1(new_n9262_), .A2(new_n9210_), .ZN(new_n9263_));
  INV_X1     g08968(.I(new_n9262_), .ZN(new_n9264_));
  NOR2_X1    g08969(.A1(new_n9264_), .A2(new_n9209_), .ZN(new_n9265_));
  NOR2_X1    g08970(.A1(new_n9265_), .A2(new_n9263_), .ZN(new_n9266_));
  NOR2_X1    g08971(.A1(new_n9208_), .A2(new_n9266_), .ZN(new_n9267_));
  XOR2_X1    g08972(.A1(new_n9262_), .A2(new_n9209_), .Z(new_n9268_));
  NOR2_X1    g08973(.A1(new_n9207_), .A2(new_n9268_), .ZN(new_n9269_));
  NOR2_X1    g08974(.A1(new_n9267_), .A2(new_n9269_), .ZN(new_n9270_));
  INV_X1     g08975(.I(new_n9181_), .ZN(new_n9271_));
  AOI21_X1   g08976(.A1(new_n9100_), .A2(new_n9271_), .B(new_n9183_), .ZN(new_n9272_));
  AOI21_X1   g08977(.A1(new_n9107_), .A2(new_n9111_), .B(new_n9109_), .ZN(new_n9273_));
  INV_X1     g08978(.I(new_n8979_), .ZN(new_n9274_));
  AOI21_X1   g08979(.A1(new_n9274_), .A2(new_n8982_), .B(new_n8978_), .ZN(new_n9275_));
  OAI21_X1   g08980(.A1(new_n8939_), .A2(new_n8946_), .B(new_n8932_), .ZN(new_n9276_));
  OAI21_X1   g08981(.A1(new_n8940_), .A2(new_n8947_), .B(new_n9276_), .ZN(new_n9277_));
  NOR2_X1    g08982(.A1(new_n8929_), .A2(new_n8926_), .ZN(new_n9278_));
  AOI21_X1   g08983(.A1(new_n2328_), .A2(new_n6056_), .B(new_n8942_), .ZN(new_n9279_));
  AOI21_X1   g08984(.A1(new_n2752_), .A2(new_n5600_), .B(new_n9037_), .ZN(new_n9280_));
  XOR2_X1    g08985(.A1(new_n9279_), .A2(new_n9280_), .Z(new_n9281_));
  AND2_X2    g08986(.A1(new_n9279_), .A2(new_n9280_), .Z(new_n9282_));
  NOR2_X1    g08987(.A1(new_n9279_), .A2(new_n9280_), .ZN(new_n9283_));
  NOR2_X1    g08988(.A1(new_n9282_), .A2(new_n9283_), .ZN(new_n9284_));
  NOR2_X1    g08989(.A1(new_n9284_), .A2(new_n9278_), .ZN(new_n9285_));
  AOI21_X1   g08990(.A1(new_n9278_), .A2(new_n9281_), .B(new_n9285_), .ZN(new_n9286_));
  XNOR2_X1   g08991(.A1(new_n9277_), .A2(new_n9286_), .ZN(new_n9287_));
  NOR2_X1    g08992(.A1(new_n9287_), .A2(new_n9275_), .ZN(new_n9288_));
  INV_X1     g08993(.I(new_n9275_), .ZN(new_n9289_));
  NOR2_X1    g08994(.A1(new_n9277_), .A2(new_n9286_), .ZN(new_n9290_));
  INV_X1     g08995(.I(new_n9290_), .ZN(new_n9291_));
  NAND2_X1   g08996(.A1(new_n9277_), .A2(new_n9286_), .ZN(new_n9292_));
  AOI21_X1   g08997(.A1(new_n9291_), .A2(new_n9292_), .B(new_n9289_), .ZN(new_n9293_));
  NOR2_X1    g08998(.A1(new_n9288_), .A2(new_n9293_), .ZN(new_n9294_));
  AOI21_X1   g08999(.A1(new_n9122_), .A2(new_n9126_), .B(new_n9124_), .ZN(new_n9295_));
  NOR2_X1    g09000(.A1(new_n5745_), .A2(new_n6945_), .ZN(new_n9296_));
  INV_X1     g09001(.I(new_n9296_), .ZN(new_n9297_));
  NOR2_X1    g09002(.A1(new_n9297_), .A2(new_n1785_), .ZN(new_n9298_));
  NOR2_X1    g09003(.A1(new_n5745_), .A2(new_n6999_), .ZN(new_n9299_));
  NAND4_X1   g09004(.A1(new_n9298_), .A2(\a[9] ), .A3(new_n9299_), .A4(\a[15] ), .ZN(new_n9300_));
  AOI21_X1   g09005(.A1(new_n9300_), .A2(new_n8005_), .B(new_n525_), .ZN(new_n9301_));
  NAND2_X1   g09006(.A1(\a[9] ), .A2(\a[55] ), .ZN(new_n9302_));
  NOR2_X1    g09007(.A1(new_n9301_), .A2(new_n9298_), .ZN(new_n9303_));
  INV_X1     g09008(.I(new_n9303_), .ZN(new_n9304_));
  NAND2_X1   g09009(.A1(new_n9297_), .A2(new_n1785_), .ZN(new_n9305_));
  OAI22_X1   g09010(.A1(new_n9304_), .A2(new_n9305_), .B1(new_n9301_), .B2(new_n9302_), .ZN(new_n9306_));
  NOR2_X1    g09011(.A1(new_n650_), .A2(new_n5745_), .ZN(new_n9307_));
  OAI21_X1   g09012(.A1(new_n3981_), .A2(new_n8973_), .B(new_n9307_), .ZN(new_n9308_));
  OAI21_X1   g09013(.A1(new_n4184_), .A2(new_n8974_), .B(new_n9308_), .ZN(new_n9309_));
  INV_X1     g09014(.I(\a[63] ), .ZN(new_n9310_));
  NOR3_X1    g09015(.A1(new_n194_), .A2(new_n9310_), .A3(\a[62] ), .ZN(new_n9311_));
  AOI21_X1   g09016(.A1(\a[1] ), .A2(\a[63] ), .B(new_n9029_), .ZN(new_n9312_));
  OAI21_X1   g09017(.A1(new_n9312_), .A2(new_n9311_), .B(\a[32] ), .ZN(new_n9313_));
  XNOR2_X1   g09018(.A1(new_n9309_), .A2(new_n9313_), .ZN(new_n9314_));
  AOI22_X1   g09019(.A1(new_n1220_), .A2(new_n7000_), .B1(new_n6777_), .B2(new_n1001_), .ZN(new_n9315_));
  NOR2_X1    g09020(.A1(new_n599_), .A2(new_n6260_), .ZN(new_n9316_));
  NAND4_X1   g09021(.A1(new_n9315_), .A2(new_n651_), .A3(new_n8056_), .A4(new_n9316_), .ZN(new_n9317_));
  NOR2_X1    g09022(.A1(new_n9314_), .A2(new_n9317_), .ZN(new_n9318_));
  AND2_X2    g09023(.A1(new_n9314_), .A2(new_n9317_), .Z(new_n9319_));
  NOR2_X1    g09024(.A1(new_n9319_), .A2(new_n9318_), .ZN(new_n9320_));
  NOR2_X1    g09025(.A1(new_n9320_), .A2(new_n9306_), .ZN(new_n9321_));
  INV_X1     g09026(.I(new_n9306_), .ZN(new_n9322_));
  XNOR2_X1   g09027(.A1(new_n9314_), .A2(new_n9317_), .ZN(new_n9323_));
  NOR2_X1    g09028(.A1(new_n9322_), .A2(new_n9323_), .ZN(new_n9324_));
  NOR2_X1    g09029(.A1(new_n9324_), .A2(new_n9321_), .ZN(new_n9325_));
  AOI21_X1   g09030(.A1(new_n8988_), .A2(new_n9007_), .B(new_n9005_), .ZN(new_n9326_));
  NOR2_X1    g09031(.A1(new_n9325_), .A2(new_n9326_), .ZN(new_n9327_));
  INV_X1     g09032(.I(new_n9326_), .ZN(new_n9328_));
  NOR3_X1    g09033(.A1(new_n9321_), .A2(new_n9324_), .A3(new_n9328_), .ZN(new_n9329_));
  NOR2_X1    g09034(.A1(new_n9327_), .A2(new_n9329_), .ZN(new_n9330_));
  NOR2_X1    g09035(.A1(new_n9330_), .A2(new_n9295_), .ZN(new_n9331_));
  INV_X1     g09036(.I(new_n9295_), .ZN(new_n9332_));
  XOR2_X1    g09037(.A1(new_n9325_), .A2(new_n9328_), .Z(new_n9333_));
  NOR2_X1    g09038(.A1(new_n9333_), .A2(new_n9332_), .ZN(new_n9334_));
  NOR2_X1    g09039(.A1(new_n9334_), .A2(new_n9331_), .ZN(new_n9335_));
  XOR2_X1    g09040(.A1(new_n9335_), .A2(new_n9294_), .Z(new_n9336_));
  NOR2_X1    g09041(.A1(new_n9336_), .A2(new_n9273_), .ZN(new_n9337_));
  INV_X1     g09042(.I(new_n9273_), .ZN(new_n9338_));
  INV_X1     g09043(.I(new_n9294_), .ZN(new_n9339_));
  NOR2_X1    g09044(.A1(new_n9339_), .A2(new_n9335_), .ZN(new_n9340_));
  INV_X1     g09045(.I(new_n9340_), .ZN(new_n9341_));
  NAND2_X1   g09046(.A1(new_n9339_), .A2(new_n9335_), .ZN(new_n9342_));
  AOI21_X1   g09047(.A1(new_n9341_), .A2(new_n9342_), .B(new_n9338_), .ZN(new_n9343_));
  NOR2_X1    g09048(.A1(new_n9337_), .A2(new_n9343_), .ZN(new_n9344_));
  INV_X1     g09049(.I(new_n9173_), .ZN(new_n9345_));
  AOI21_X1   g09050(.A1(new_n9345_), .A2(new_n9128_), .B(new_n9175_), .ZN(new_n9346_));
  NOR2_X1    g09051(.A1(new_n885_), .A2(new_n7727_), .ZN(new_n9347_));
  INV_X1     g09052(.I(new_n9347_), .ZN(new_n9348_));
  NOR3_X1    g09053(.A1(new_n9348_), .A2(new_n268_), .A3(new_n5511_), .ZN(new_n9349_));
  NOR4_X1    g09054(.A1(new_n242_), .A2(new_n885_), .A3(new_n5511_), .A4(new_n7647_), .ZN(new_n9350_));
  NAND2_X1   g09055(.A1(new_n9349_), .A2(new_n9350_), .ZN(new_n9351_));
  AOI21_X1   g09056(.A1(new_n9351_), .A2(new_n8246_), .B(new_n478_), .ZN(new_n9352_));
  NOR3_X1    g09057(.A1(new_n9352_), .A2(new_n242_), .A3(new_n7647_), .ZN(new_n9353_));
  OAI21_X1   g09058(.A1(new_n268_), .A2(new_n7727_), .B(new_n5907_), .ZN(new_n9354_));
  NOR2_X1    g09059(.A1(new_n9352_), .A2(new_n9349_), .ZN(new_n9355_));
  AOI21_X1   g09060(.A1(new_n9354_), .A2(new_n9355_), .B(new_n9353_), .ZN(new_n9356_));
  NOR2_X1    g09061(.A1(new_n7023_), .A2(new_n5322_), .ZN(new_n9357_));
  NOR2_X1    g09062(.A1(new_n9357_), .A2(new_n7009_), .ZN(new_n9358_));
  NOR4_X1    g09063(.A1(new_n5173_), .A2(new_n4538_), .A3(new_n1215_), .A4(new_n4770_), .ZN(new_n9359_));
  NAND2_X1   g09064(.A1(new_n9358_), .A2(new_n9359_), .ZN(new_n9360_));
  AOI22_X1   g09065(.A1(new_n1913_), .A2(new_n5592_), .B1(new_n4415_), .B2(new_n2543_), .ZN(new_n9361_));
  INV_X1     g09066(.I(new_n9361_), .ZN(new_n9362_));
  NAND4_X1   g09067(.A1(new_n2276_), .A2(new_n4321_), .A3(\a[23] ), .A4(\a[41] ), .ZN(new_n9363_));
  NOR3_X1    g09068(.A1(new_n9360_), .A2(new_n9362_), .A3(new_n9363_), .ZN(new_n9364_));
  INV_X1     g09069(.I(new_n9360_), .ZN(new_n9365_));
  NOR2_X1    g09070(.A1(new_n9362_), .A2(new_n9363_), .ZN(new_n9366_));
  NOR2_X1    g09071(.A1(new_n9365_), .A2(new_n9366_), .ZN(new_n9367_));
  OAI21_X1   g09072(.A1(new_n9364_), .A2(new_n9367_), .B(new_n9356_), .ZN(new_n9368_));
  XOR2_X1    g09073(.A1(new_n9360_), .A2(new_n9366_), .Z(new_n9369_));
  OAI21_X1   g09074(.A1(new_n9356_), .A2(new_n9369_), .B(new_n9368_), .ZN(new_n9370_));
  NAND3_X1   g09075(.A1(new_n1722_), .A2(\a[48] ), .A3(\a[56] ), .ZN(new_n9371_));
  NAND2_X1   g09076(.A1(\a[26] ), .A2(\a[38] ), .ZN(new_n9372_));
  XNOR2_X1   g09077(.A1(new_n9371_), .A2(new_n9372_), .ZN(new_n9373_));
  INV_X1     g09078(.I(new_n4190_), .ZN(new_n9374_));
  INV_X1     g09079(.I(new_n5184_), .ZN(new_n9375_));
  OAI22_X1   g09080(.A1(new_n3839_), .A2(new_n9375_), .B1(new_n3174_), .B2(new_n2692_), .ZN(new_n9376_));
  NOR4_X1    g09081(.A1(new_n9376_), .A2(new_n2690_), .A3(new_n3966_), .A4(new_n9374_), .ZN(new_n9377_));
  INV_X1     g09082(.I(new_n9377_), .ZN(new_n9378_));
  INV_X1     g09083(.I(new_n8430_), .ZN(new_n9379_));
  NAND2_X1   g09084(.A1(new_n2870_), .A2(new_n4041_), .ZN(new_n9380_));
  AOI21_X1   g09085(.A1(new_n9380_), .A2(new_n9379_), .B(new_n4644_), .ZN(new_n9381_));
  AND2_X2    g09086(.A1(new_n9381_), .A2(new_n3127_), .Z(new_n9382_));
  NOR2_X1    g09087(.A1(new_n9381_), .A2(new_n3127_), .ZN(new_n9383_));
  NOR2_X1    g09088(.A1(new_n9382_), .A2(new_n9383_), .ZN(new_n9384_));
  NOR2_X1    g09089(.A1(new_n9384_), .A2(new_n9378_), .ZN(new_n9385_));
  NOR3_X1    g09090(.A1(new_n9382_), .A2(new_n9377_), .A3(new_n9383_), .ZN(new_n9386_));
  NOR2_X1    g09091(.A1(new_n9385_), .A2(new_n9386_), .ZN(new_n9387_));
  XOR2_X1    g09092(.A1(new_n9384_), .A2(new_n9378_), .Z(new_n9388_));
  NAND2_X1   g09093(.A1(new_n9388_), .A2(new_n9373_), .ZN(new_n9389_));
  OAI21_X1   g09094(.A1(new_n9373_), .A2(new_n9387_), .B(new_n9389_), .ZN(new_n9390_));
  NOR2_X1    g09095(.A1(new_n199_), .A2(new_n9310_), .ZN(new_n9391_));
  OAI21_X1   g09096(.A1(new_n9033_), .A2(new_n9028_), .B(new_n9391_), .ZN(new_n9392_));
  NAND2_X1   g09097(.A1(new_n9392_), .A2(new_n9034_), .ZN(new_n9393_));
  NOR3_X1    g09098(.A1(new_n8990_), .A2(new_n8453_), .A3(new_n9029_), .ZN(new_n9394_));
  NOR2_X1    g09099(.A1(new_n1271_), .A2(new_n9394_), .ZN(new_n9395_));
  NOR4_X1    g09100(.A1(new_n8991_), .A2(new_n267_), .A3(new_n201_), .A4(new_n9029_), .ZN(new_n9396_));
  NAND2_X1   g09101(.A1(new_n9396_), .A2(new_n9395_), .ZN(new_n9397_));
  NOR2_X1    g09102(.A1(new_n353_), .A2(new_n8085_), .ZN(new_n9398_));
  XOR2_X1    g09103(.A1(new_n5488_), .A2(new_n1342_), .Z(new_n9399_));
  XNOR2_X1   g09104(.A1(new_n9397_), .A2(new_n9399_), .ZN(new_n9400_));
  INV_X1     g09105(.I(new_n9400_), .ZN(new_n9401_));
  NOR2_X1    g09106(.A1(new_n9397_), .A2(new_n9399_), .ZN(new_n9402_));
  INV_X1     g09107(.I(new_n9402_), .ZN(new_n9403_));
  NAND2_X1   g09108(.A1(new_n9397_), .A2(new_n9399_), .ZN(new_n9404_));
  AOI21_X1   g09109(.A1(new_n9403_), .A2(new_n9404_), .B(new_n9393_), .ZN(new_n9405_));
  AOI21_X1   g09110(.A1(new_n9401_), .A2(new_n9393_), .B(new_n9405_), .ZN(new_n9406_));
  XOR2_X1    g09111(.A1(new_n9390_), .A2(new_n9406_), .Z(new_n9407_));
  OR2_X2     g09112(.A1(new_n9390_), .A2(new_n9406_), .Z(new_n9408_));
  NAND2_X1   g09113(.A1(new_n9390_), .A2(new_n9406_), .ZN(new_n9409_));
  NAND2_X1   g09114(.A1(new_n9408_), .A2(new_n9409_), .ZN(new_n9410_));
  MUX2_X1    g09115(.I0(new_n9410_), .I1(new_n9407_), .S(new_n9370_), .Z(new_n9411_));
  AOI21_X1   g09116(.A1(new_n9077_), .A2(new_n9081_), .B(new_n9079_), .ZN(new_n9412_));
  INV_X1     g09117(.I(new_n9144_), .ZN(new_n9413_));
  AOI21_X1   g09118(.A1(new_n9132_), .A2(new_n9413_), .B(new_n9143_), .ZN(new_n9414_));
  INV_X1     g09119(.I(new_n9069_), .ZN(new_n9415_));
  AOI21_X1   g09120(.A1(new_n9415_), .A2(new_n9066_), .B(new_n9068_), .ZN(new_n9416_));
  NAND2_X1   g09121(.A1(new_n9160_), .A2(new_n9148_), .ZN(new_n9417_));
  NAND2_X1   g09122(.A1(new_n9417_), .A2(new_n9159_), .ZN(new_n9418_));
  XOR2_X1    g09123(.A1(new_n9416_), .A2(new_n9418_), .Z(new_n9419_));
  INV_X1     g09124(.I(new_n9418_), .ZN(new_n9420_));
  NOR2_X1    g09125(.A1(new_n9420_), .A2(new_n9416_), .ZN(new_n9421_));
  NAND2_X1   g09126(.A1(new_n9420_), .A2(new_n9416_), .ZN(new_n9422_));
  INV_X1     g09127(.I(new_n9422_), .ZN(new_n9423_));
  OAI21_X1   g09128(.A1(new_n9423_), .A2(new_n9421_), .B(new_n9414_), .ZN(new_n9424_));
  OAI21_X1   g09129(.A1(new_n9414_), .A2(new_n9419_), .B(new_n9424_), .ZN(new_n9425_));
  INV_X1     g09130(.I(new_n9167_), .ZN(new_n9426_));
  AOI21_X1   g09131(.A1(new_n9147_), .A2(new_n9426_), .B(new_n9165_), .ZN(new_n9427_));
  XNOR2_X1   g09132(.A1(new_n9425_), .A2(new_n9427_), .ZN(new_n9428_));
  NOR2_X1    g09133(.A1(new_n9425_), .A2(new_n9427_), .ZN(new_n9429_));
  AND2_X2    g09134(.A1(new_n9425_), .A2(new_n9427_), .Z(new_n9430_));
  OAI21_X1   g09135(.A1(new_n9430_), .A2(new_n9429_), .B(new_n9412_), .ZN(new_n9431_));
  OAI21_X1   g09136(.A1(new_n9412_), .A2(new_n9428_), .B(new_n9431_), .ZN(new_n9432_));
  NAND2_X1   g09137(.A1(new_n9432_), .A2(new_n9411_), .ZN(new_n9433_));
  NOR2_X1    g09138(.A1(new_n9432_), .A2(new_n9411_), .ZN(new_n9434_));
  INV_X1     g09139(.I(new_n9434_), .ZN(new_n9435_));
  AOI21_X1   g09140(.A1(new_n9435_), .A2(new_n9433_), .B(new_n9346_), .ZN(new_n9436_));
  XNOR2_X1   g09141(.A1(new_n9432_), .A2(new_n9411_), .ZN(new_n9437_));
  INV_X1     g09142(.I(new_n9437_), .ZN(new_n9438_));
  AOI21_X1   g09143(.A1(new_n9438_), .A2(new_n9346_), .B(new_n9436_), .ZN(new_n9439_));
  XOR2_X1    g09144(.A1(new_n9439_), .A2(new_n9344_), .Z(new_n9440_));
  NOR2_X1    g09145(.A1(new_n9440_), .A2(new_n9272_), .ZN(new_n9441_));
  INV_X1     g09146(.I(new_n9272_), .ZN(new_n9442_));
  INV_X1     g09147(.I(new_n9344_), .ZN(new_n9443_));
  NOR2_X1    g09148(.A1(new_n9439_), .A2(new_n9443_), .ZN(new_n9444_));
  INV_X1     g09149(.I(new_n9444_), .ZN(new_n9445_));
  NAND2_X1   g09150(.A1(new_n9439_), .A2(new_n9443_), .ZN(new_n9446_));
  AOI21_X1   g09151(.A1(new_n9445_), .A2(new_n9446_), .B(new_n9442_), .ZN(new_n9447_));
  NOR2_X1    g09152(.A1(new_n9441_), .A2(new_n9447_), .ZN(new_n9448_));
  XOR2_X1    g09153(.A1(new_n9448_), .A2(new_n9270_), .Z(new_n9449_));
  NOR2_X1    g09154(.A1(new_n9449_), .A2(new_n9206_), .ZN(new_n9450_));
  INV_X1     g09155(.I(new_n9270_), .ZN(new_n9451_));
  NOR2_X1    g09156(.A1(new_n9451_), .A2(new_n9448_), .ZN(new_n9452_));
  INV_X1     g09157(.I(new_n9452_), .ZN(new_n9453_));
  NAND2_X1   g09158(.A1(new_n9451_), .A2(new_n9448_), .ZN(new_n9454_));
  AOI21_X1   g09159(.A1(new_n9453_), .A2(new_n9454_), .B(new_n9205_), .ZN(new_n9455_));
  NOR2_X1    g09160(.A1(new_n9450_), .A2(new_n9455_), .ZN(new_n9456_));
  INV_X1     g09161(.I(new_n9456_), .ZN(new_n9457_));
  AOI21_X1   g09162(.A1(new_n9189_), .A2(new_n9193_), .B(new_n9191_), .ZN(new_n9458_));
  NOR2_X1    g09163(.A1(new_n9457_), .A2(new_n9458_), .ZN(new_n9459_));
  NAND2_X1   g09164(.A1(new_n9457_), .A2(new_n9458_), .ZN(new_n9460_));
  INV_X1     g09165(.I(new_n9460_), .ZN(new_n9461_));
  NOR2_X1    g09166(.A1(new_n9461_), .A2(new_n9459_), .ZN(new_n9462_));
  XOR2_X1    g09167(.A1(new_n9204_), .A2(new_n9462_), .Z(\asquared[65] ));
  NOR2_X1    g09168(.A1(new_n9199_), .A2(new_n9459_), .ZN(new_n9464_));
  AOI21_X1   g09169(.A1(new_n9199_), .A2(new_n9459_), .B(new_n8916_), .ZN(new_n9465_));
  NOR2_X1    g09170(.A1(new_n9465_), .A2(new_n9464_), .ZN(new_n9466_));
  INV_X1     g09171(.I(new_n9466_), .ZN(new_n9467_));
  NOR4_X1    g09172(.A1(new_n8144_), .A2(new_n8659_), .A3(new_n8663_), .A4(new_n9467_), .ZN(new_n9468_));
  INV_X1     g09173(.I(new_n9263_), .ZN(new_n9469_));
  AOI21_X1   g09174(.A1(new_n9207_), .A2(new_n9469_), .B(new_n9265_), .ZN(new_n9470_));
  OAI21_X1   g09175(.A1(new_n9213_), .A2(new_n9258_), .B(new_n9260_), .ZN(new_n9471_));
  OAI21_X1   g09176(.A1(new_n9275_), .A2(new_n9290_), .B(new_n9292_), .ZN(new_n9472_));
  INV_X1     g09177(.I(new_n9472_), .ZN(new_n9473_));
  NOR3_X1    g09178(.A1(new_n9283_), .A2(new_n8926_), .A3(new_n8929_), .ZN(new_n9474_));
  NOR2_X1    g09179(.A1(new_n9474_), .A2(new_n9282_), .ZN(new_n9475_));
  INV_X1     g09180(.I(new_n9227_), .ZN(new_n9476_));
  AOI21_X1   g09181(.A1(new_n9216_), .A2(new_n9476_), .B(new_n9226_), .ZN(new_n9477_));
  NOR2_X1    g09182(.A1(new_n8963_), .A2(new_n9242_), .ZN(new_n9478_));
  NOR2_X1    g09183(.A1(new_n9478_), .A2(new_n9241_), .ZN(new_n9479_));
  XNOR2_X1   g09184(.A1(new_n9479_), .A2(new_n9477_), .ZN(new_n9480_));
  NOR2_X1    g09185(.A1(new_n9480_), .A2(new_n9475_), .ZN(new_n9481_));
  INV_X1     g09186(.I(new_n9475_), .ZN(new_n9482_));
  NOR2_X1    g09187(.A1(new_n9479_), .A2(new_n9477_), .ZN(new_n9483_));
  INV_X1     g09188(.I(new_n9483_), .ZN(new_n9484_));
  NAND2_X1   g09189(.A1(new_n9479_), .A2(new_n9477_), .ZN(new_n9485_));
  AOI21_X1   g09190(.A1(new_n9484_), .A2(new_n9485_), .B(new_n9482_), .ZN(new_n9486_));
  NOR2_X1    g09191(.A1(new_n9481_), .A2(new_n9486_), .ZN(new_n9487_));
  NOR2_X1    g09192(.A1(new_n9250_), .A2(new_n9231_), .ZN(new_n9488_));
  NOR2_X1    g09193(.A1(new_n9488_), .A2(new_n9247_), .ZN(new_n9489_));
  XOR2_X1    g09194(.A1(new_n9489_), .A2(new_n9487_), .Z(new_n9490_));
  NOR2_X1    g09195(.A1(new_n9490_), .A2(new_n9473_), .ZN(new_n9491_));
  INV_X1     g09196(.I(new_n9487_), .ZN(new_n9492_));
  NOR2_X1    g09197(.A1(new_n9489_), .A2(new_n9492_), .ZN(new_n9493_));
  INV_X1     g09198(.I(new_n9493_), .ZN(new_n9494_));
  NAND2_X1   g09199(.A1(new_n9489_), .A2(new_n9492_), .ZN(new_n9495_));
  AOI21_X1   g09200(.A1(new_n9494_), .A2(new_n9495_), .B(new_n9472_), .ZN(new_n9496_));
  NOR2_X1    g09201(.A1(new_n9491_), .A2(new_n9496_), .ZN(new_n9497_));
  INV_X1     g09202(.I(new_n9497_), .ZN(new_n9498_));
  NOR2_X1    g09203(.A1(new_n1215_), .A2(new_n6999_), .ZN(new_n9499_));
  NAND2_X1   g09204(.A1(new_n7024_), .A2(new_n9499_), .ZN(new_n9500_));
  INV_X1     g09205(.I(new_n9500_), .ZN(new_n9501_));
  NOR2_X1    g09206(.A1(new_n1215_), .A2(new_n7216_), .ZN(new_n9502_));
  NAND4_X1   g09207(.A1(new_n9501_), .A2(\a[9] ), .A3(\a[45] ), .A4(new_n9502_), .ZN(new_n9503_));
  AOI21_X1   g09208(.A1(new_n9503_), .A2(new_n8953_), .B(new_n525_), .ZN(new_n9504_));
  NOR3_X1    g09209(.A1(new_n9504_), .A2(new_n364_), .A3(new_n7216_), .ZN(new_n9505_));
  NOR2_X1    g09210(.A1(new_n9504_), .A2(new_n9501_), .ZN(new_n9506_));
  NOR2_X1    g09211(.A1(new_n5004_), .A2(new_n6999_), .ZN(new_n9507_));
  NOR2_X1    g09212(.A1(new_n2548_), .A2(new_n9507_), .ZN(new_n9508_));
  AOI21_X1   g09213(.A1(new_n9506_), .A2(new_n9508_), .B(new_n9505_), .ZN(new_n9509_));
  NOR2_X1    g09214(.A1(new_n6700_), .A2(new_n6390_), .ZN(new_n9510_));
  NOR4_X1    g09215(.A1(new_n5592_), .A2(new_n2277_), .A3(new_n2368_), .A4(new_n4769_), .ZN(new_n9511_));
  NAND2_X1   g09216(.A1(new_n9511_), .A2(new_n9510_), .ZN(new_n9512_));
  AOI22_X1   g09217(.A1(new_n2533_), .A2(new_n5601_), .B1(new_n5339_), .B2(new_n3037_), .ZN(new_n9513_));
  NAND4_X1   g09218(.A1(new_n9513_), .A2(new_n2692_), .A3(new_n4329_), .A4(new_n4706_), .ZN(new_n9514_));
  NOR2_X1    g09219(.A1(new_n9514_), .A2(new_n9512_), .ZN(new_n9515_));
  INV_X1     g09220(.I(new_n9512_), .ZN(new_n9516_));
  INV_X1     g09221(.I(new_n9514_), .ZN(new_n9517_));
  NOR2_X1    g09222(.A1(new_n9517_), .A2(new_n9516_), .ZN(new_n9518_));
  OAI21_X1   g09223(.A1(new_n9515_), .A2(new_n9518_), .B(new_n9509_), .ZN(new_n9519_));
  XNOR2_X1   g09224(.A1(new_n9514_), .A2(new_n9512_), .ZN(new_n9520_));
  OAI21_X1   g09225(.A1(new_n9509_), .A2(new_n9520_), .B(new_n9519_), .ZN(new_n9521_));
  INV_X1     g09226(.I(new_n9521_), .ZN(new_n9522_));
  NOR2_X1    g09227(.A1(new_n3852_), .A2(new_n3712_), .ZN(new_n9523_));
  AOI21_X1   g09228(.A1(new_n3126_), .A2(new_n4163_), .B(new_n9523_), .ZN(new_n9524_));
  NOR2_X1    g09229(.A1(new_n4644_), .A2(new_n4184_), .ZN(new_n9525_));
  AOI21_X1   g09230(.A1(\a[31] ), .A2(\a[34] ), .B(new_n3851_), .ZN(new_n9526_));
  NOR3_X1    g09231(.A1(new_n9525_), .A2(new_n4164_), .A3(new_n9526_), .ZN(new_n9527_));
  AND2_X2    g09232(.A1(new_n9524_), .A2(new_n9527_), .Z(new_n9528_));
  NOR2_X1    g09233(.A1(new_n1339_), .A2(new_n5175_), .ZN(new_n9529_));
  INV_X1     g09234(.I(new_n9529_), .ZN(new_n9530_));
  NOR2_X1    g09235(.A1(new_n2499_), .A2(new_n3393_), .ZN(new_n9531_));
  INV_X1     g09236(.I(new_n9531_), .ZN(new_n9532_));
  NOR2_X1    g09237(.A1(new_n9530_), .A2(new_n9532_), .ZN(new_n9533_));
  XOR2_X1    g09238(.A1(new_n9533_), .A2(new_n675_), .Z(new_n9534_));
  XOR2_X1    g09239(.A1(new_n9534_), .A2(\a[54] ), .Z(new_n9535_));
  NOR2_X1    g09240(.A1(new_n885_), .A2(new_n5750_), .ZN(new_n9536_));
  NAND2_X1   g09241(.A1(new_n9536_), .A2(\a[33] ), .ZN(new_n9537_));
  XOR2_X1    g09242(.A1(new_n9537_), .A2(\a[3] ), .Z(new_n9538_));
  XOR2_X1    g09243(.A1(new_n9538_), .A2(\a[62] ), .Z(new_n9539_));
  NOR2_X1    g09244(.A1(new_n9535_), .A2(new_n9539_), .ZN(new_n9540_));
  NAND2_X1   g09245(.A1(new_n9535_), .A2(new_n9539_), .ZN(new_n9541_));
  INV_X1     g09246(.I(new_n9541_), .ZN(new_n9542_));
  OAI21_X1   g09247(.A1(new_n9542_), .A2(new_n9540_), .B(new_n9528_), .ZN(new_n9543_));
  XNOR2_X1   g09248(.A1(new_n9535_), .A2(new_n9539_), .ZN(new_n9544_));
  OAI21_X1   g09249(.A1(new_n9528_), .A2(new_n9544_), .B(new_n9543_), .ZN(new_n9545_));
  NAND2_X1   g09250(.A1(new_n5321_), .A2(new_n4538_), .ZN(new_n9546_));
  NAND2_X1   g09251(.A1(\a[8] ), .A2(\a[57] ), .ZN(new_n9547_));
  XNOR2_X1   g09252(.A1(new_n9546_), .A2(new_n9547_), .ZN(new_n9548_));
  NOR2_X1    g09253(.A1(new_n9029_), .A2(new_n9310_), .ZN(new_n9549_));
  INV_X1     g09254(.I(new_n9549_), .ZN(new_n9550_));
  NAND2_X1   g09255(.A1(new_n9309_), .A2(new_n2972_), .ZN(new_n9551_));
  OAI21_X1   g09256(.A1(new_n9313_), .A2(new_n9550_), .B(new_n9551_), .ZN(new_n9552_));
  INV_X1     g09257(.I(new_n8996_), .ZN(new_n9553_));
  NOR2_X1    g09258(.A1(new_n7647_), .A2(new_n8990_), .ZN(new_n9554_));
  INV_X1     g09259(.I(new_n9554_), .ZN(new_n9555_));
  NOR2_X1    g09260(.A1(new_n9553_), .A2(new_n9555_), .ZN(new_n9556_));
  AOI21_X1   g09261(.A1(new_n608_), .A2(new_n1151_), .B(new_n9556_), .ZN(new_n9557_));
  NOR4_X1    g09262(.A1(new_n8676_), .A2(new_n479_), .A3(new_n353_), .A4(new_n8990_), .ZN(new_n9558_));
  AND2_X2    g09263(.A1(new_n9557_), .A2(new_n9558_), .Z(new_n9559_));
  XNOR2_X1   g09264(.A1(new_n9552_), .A2(new_n9559_), .ZN(new_n9560_));
  NOR2_X1    g09265(.A1(new_n9560_), .A2(new_n9548_), .ZN(new_n9561_));
  INV_X1     g09266(.I(new_n9548_), .ZN(new_n9562_));
  INV_X1     g09267(.I(new_n9552_), .ZN(new_n9563_));
  INV_X1     g09268(.I(new_n9559_), .ZN(new_n9564_));
  NOR2_X1    g09269(.A1(new_n9563_), .A2(new_n9564_), .ZN(new_n9565_));
  NOR2_X1    g09270(.A1(new_n9552_), .A2(new_n9559_), .ZN(new_n9566_));
  NOR2_X1    g09271(.A1(new_n9565_), .A2(new_n9566_), .ZN(new_n9567_));
  NOR2_X1    g09272(.A1(new_n9567_), .A2(new_n9562_), .ZN(new_n9568_));
  NOR2_X1    g09273(.A1(new_n9568_), .A2(new_n9561_), .ZN(new_n9569_));
  NOR2_X1    g09274(.A1(new_n9545_), .A2(new_n9569_), .ZN(new_n9570_));
  INV_X1     g09275(.I(new_n9570_), .ZN(new_n9571_));
  NAND2_X1   g09276(.A1(new_n9545_), .A2(new_n9569_), .ZN(new_n9572_));
  AOI21_X1   g09277(.A1(new_n9571_), .A2(new_n9572_), .B(new_n9522_), .ZN(new_n9573_));
  XNOR2_X1   g09278(.A1(new_n9545_), .A2(new_n9569_), .ZN(new_n9574_));
  NOR2_X1    g09279(.A1(new_n9574_), .A2(new_n9521_), .ZN(new_n9575_));
  NOR2_X1    g09280(.A1(new_n9573_), .A2(new_n9575_), .ZN(new_n9576_));
  NOR2_X1    g09281(.A1(new_n9498_), .A2(new_n9576_), .ZN(new_n9577_));
  INV_X1     g09282(.I(new_n9577_), .ZN(new_n9578_));
  NAND2_X1   g09283(.A1(new_n9498_), .A2(new_n9576_), .ZN(new_n9579_));
  NAND2_X1   g09284(.A1(new_n9578_), .A2(new_n9579_), .ZN(new_n9580_));
  XOR2_X1    g09285(.A1(new_n9497_), .A2(new_n9576_), .Z(new_n9581_));
  NOR2_X1    g09286(.A1(new_n9581_), .A2(new_n9471_), .ZN(new_n9582_));
  AOI21_X1   g09287(.A1(new_n9471_), .A2(new_n9580_), .B(new_n9582_), .ZN(new_n9583_));
  INV_X1     g09288(.I(new_n9367_), .ZN(new_n9584_));
  AOI21_X1   g09289(.A1(new_n9356_), .A2(new_n9584_), .B(new_n9364_), .ZN(new_n9585_));
  AOI21_X1   g09290(.A1(new_n4538_), .A2(new_n5173_), .B(new_n9358_), .ZN(new_n9586_));
  INV_X1     g09291(.I(new_n9586_), .ZN(new_n9587_));
  OAI21_X1   g09292(.A1(new_n2689_), .A2(new_n3967_), .B(new_n9376_), .ZN(new_n9588_));
  AOI21_X1   g09293(.A1(new_n3061_), .A2(new_n7204_), .B(new_n9315_), .ZN(new_n9589_));
  XOR2_X1    g09294(.A1(new_n9588_), .A2(new_n9589_), .Z(new_n9590_));
  NOR2_X1    g09295(.A1(new_n9590_), .A2(new_n9587_), .ZN(new_n9591_));
  INV_X1     g09296(.I(new_n9589_), .ZN(new_n9592_));
  NOR2_X1    g09297(.A1(new_n9592_), .A2(new_n9588_), .ZN(new_n9593_));
  INV_X1     g09298(.I(new_n9593_), .ZN(new_n9594_));
  NAND2_X1   g09299(.A1(new_n9592_), .A2(new_n9588_), .ZN(new_n9595_));
  AOI21_X1   g09300(.A1(new_n9594_), .A2(new_n9595_), .B(new_n9586_), .ZN(new_n9596_));
  NOR2_X1    g09301(.A1(new_n9591_), .A2(new_n9596_), .ZN(new_n9597_));
  NOR2_X1    g09302(.A1(new_n9386_), .A2(new_n9373_), .ZN(new_n9598_));
  NOR2_X1    g09303(.A1(new_n9598_), .A2(new_n9385_), .ZN(new_n9599_));
  XOR2_X1    g09304(.A1(new_n9597_), .A2(new_n9599_), .Z(new_n9600_));
  NOR2_X1    g09305(.A1(new_n9600_), .A2(new_n9585_), .ZN(new_n9601_));
  INV_X1     g09306(.I(new_n9585_), .ZN(new_n9602_));
  INV_X1     g09307(.I(new_n9597_), .ZN(new_n9603_));
  NOR2_X1    g09308(.A1(new_n9603_), .A2(new_n9599_), .ZN(new_n9604_));
  INV_X1     g09309(.I(new_n9604_), .ZN(new_n9605_));
  NAND2_X1   g09310(.A1(new_n9603_), .A2(new_n9599_), .ZN(new_n9606_));
  AOI21_X1   g09311(.A1(new_n9605_), .A2(new_n9606_), .B(new_n9602_), .ZN(new_n9607_));
  NOR2_X1    g09312(.A1(new_n9607_), .A2(new_n9601_), .ZN(new_n9608_));
  NOR2_X1    g09313(.A1(new_n9430_), .A2(new_n9412_), .ZN(new_n9609_));
  NOR2_X1    g09314(.A1(new_n9609_), .A2(new_n9429_), .ZN(new_n9610_));
  INV_X1     g09315(.I(new_n9414_), .ZN(new_n9611_));
  AOI21_X1   g09316(.A1(new_n9611_), .A2(new_n9422_), .B(new_n9421_), .ZN(new_n9612_));
  OAI22_X1   g09317(.A1(new_n9380_), .A2(new_n3127_), .B1(new_n4644_), .B2(new_n9379_), .ZN(new_n9613_));
  NAND2_X1   g09318(.A1(\a[4] ), .A2(\a[63] ), .ZN(new_n9614_));
  XOR2_X1    g09319(.A1(new_n8997_), .A2(new_n9614_), .Z(new_n9615_));
  INV_X1     g09320(.I(new_n9615_), .ZN(new_n9616_));
  NAND2_X1   g09321(.A1(new_n9613_), .A2(new_n9616_), .ZN(new_n9617_));
  NOR2_X1    g09322(.A1(new_n9613_), .A2(new_n9616_), .ZN(new_n9618_));
  INV_X1     g09323(.I(new_n9618_), .ZN(new_n9619_));
  AND2_X2    g09324(.A1(new_n9619_), .A2(new_n9617_), .Z(new_n9620_));
  NOR2_X1    g09325(.A1(new_n8925_), .A2(new_n1002_), .ZN(new_n9621_));
  NOR4_X1    g09326(.A1(new_n566_), .A2(new_n1276_), .A3(new_n5511_), .A4(new_n6694_), .ZN(new_n9622_));
  NAND2_X1   g09327(.A1(new_n9621_), .A2(new_n9622_), .ZN(new_n9623_));
  AOI21_X1   g09328(.A1(new_n9623_), .A2(new_n1150_), .B(new_n8056_), .ZN(new_n9624_));
  NOR3_X1    g09329(.A1(new_n9624_), .A2(new_n566_), .A3(new_n6694_), .ZN(new_n9625_));
  NOR3_X1    g09330(.A1(new_n9624_), .A2(new_n1012_), .A3(new_n8924_), .ZN(new_n9626_));
  NOR2_X1    g09331(.A1(new_n9625_), .A2(new_n9626_), .ZN(new_n9627_));
  INV_X1     g09332(.I(new_n9627_), .ZN(new_n9628_));
  NOR2_X1    g09333(.A1(new_n5745_), .A2(new_n6260_), .ZN(new_n9629_));
  AOI22_X1   g09334(.A1(new_n1718_), .A2(new_n6280_), .B1(new_n9629_), .B2(new_n1719_), .ZN(new_n9630_));
  INV_X1     g09335(.I(new_n9630_), .ZN(new_n9631_));
  NOR4_X1    g09336(.A1(new_n9631_), .A2(new_n1447_), .A3(new_n6779_), .A4(new_n7514_), .ZN(new_n9632_));
  INV_X1     g09337(.I(new_n9632_), .ZN(new_n9633_));
  NOR2_X1    g09338(.A1(new_n9628_), .A2(new_n9633_), .ZN(new_n9634_));
  NOR2_X1    g09339(.A1(new_n9627_), .A2(new_n9632_), .ZN(new_n9635_));
  NOR2_X1    g09340(.A1(new_n9634_), .A2(new_n9635_), .ZN(new_n9636_));
  NOR2_X1    g09341(.A1(new_n9636_), .A2(new_n9620_), .ZN(new_n9637_));
  INV_X1     g09342(.I(new_n9620_), .ZN(new_n9638_));
  XOR2_X1    g09343(.A1(new_n9627_), .A2(new_n9633_), .Z(new_n9639_));
  NOR2_X1    g09344(.A1(new_n9639_), .A2(new_n9638_), .ZN(new_n9640_));
  NOR2_X1    g09345(.A1(new_n9637_), .A2(new_n9640_), .ZN(new_n9641_));
  AOI21_X1   g09346(.A1(new_n9393_), .A2(new_n9404_), .B(new_n9402_), .ZN(new_n9642_));
  NOR2_X1    g09347(.A1(new_n9641_), .A2(new_n9642_), .ZN(new_n9643_));
  INV_X1     g09348(.I(new_n9642_), .ZN(new_n9644_));
  NOR3_X1    g09349(.A1(new_n9637_), .A2(new_n9640_), .A3(new_n9644_), .ZN(new_n9645_));
  NOR2_X1    g09350(.A1(new_n9643_), .A2(new_n9645_), .ZN(new_n9646_));
  NOR2_X1    g09351(.A1(new_n9646_), .A2(new_n9612_), .ZN(new_n9647_));
  INV_X1     g09352(.I(new_n9612_), .ZN(new_n9648_));
  XOR2_X1    g09353(.A1(new_n9641_), .A2(new_n9644_), .Z(new_n9649_));
  NOR2_X1    g09354(.A1(new_n9649_), .A2(new_n9648_), .ZN(new_n9650_));
  NOR2_X1    g09355(.A1(new_n9650_), .A2(new_n9647_), .ZN(new_n9651_));
  XNOR2_X1   g09356(.A1(new_n9610_), .A2(new_n9651_), .ZN(new_n9652_));
  NOR2_X1    g09357(.A1(new_n9652_), .A2(new_n9608_), .ZN(new_n9653_));
  NOR2_X1    g09358(.A1(new_n9610_), .A2(new_n9651_), .ZN(new_n9654_));
  INV_X1     g09359(.I(new_n9654_), .ZN(new_n9655_));
  NAND2_X1   g09360(.A1(new_n9610_), .A2(new_n9651_), .ZN(new_n9656_));
  NAND2_X1   g09361(.A1(new_n9655_), .A2(new_n9656_), .ZN(new_n9657_));
  AOI21_X1   g09362(.A1(new_n9608_), .A2(new_n9657_), .B(new_n9653_), .ZN(new_n9658_));
  NOR2_X1    g09363(.A1(new_n9583_), .A2(new_n9658_), .ZN(new_n9659_));
  INV_X1     g09364(.I(new_n9659_), .ZN(new_n9660_));
  NAND2_X1   g09365(.A1(new_n9583_), .A2(new_n9658_), .ZN(new_n9661_));
  AOI21_X1   g09366(.A1(new_n9660_), .A2(new_n9661_), .B(new_n9470_), .ZN(new_n9662_));
  INV_X1     g09367(.I(new_n9470_), .ZN(new_n9663_));
  XNOR2_X1   g09368(.A1(new_n9583_), .A2(new_n9658_), .ZN(new_n9664_));
  NOR2_X1    g09369(.A1(new_n9664_), .A2(new_n9663_), .ZN(new_n9665_));
  NOR2_X1    g09370(.A1(new_n9665_), .A2(new_n9662_), .ZN(new_n9666_));
  NAND2_X1   g09371(.A1(new_n9442_), .A2(new_n9446_), .ZN(new_n9667_));
  NAND2_X1   g09372(.A1(new_n9667_), .A2(new_n9445_), .ZN(new_n9668_));
  AOI21_X1   g09373(.A1(new_n9338_), .A2(new_n9342_), .B(new_n9340_), .ZN(new_n9669_));
  AOI21_X1   g09374(.A1(new_n9432_), .A2(new_n9411_), .B(new_n9346_), .ZN(new_n9670_));
  NOR2_X1    g09375(.A1(new_n9670_), .A2(new_n9434_), .ZN(new_n9671_));
  NAND2_X1   g09376(.A1(new_n9408_), .A2(new_n9370_), .ZN(new_n9672_));
  NAND2_X1   g09377(.A1(new_n9672_), .A2(new_n9409_), .ZN(new_n9673_));
  INV_X1     g09378(.I(new_n9329_), .ZN(new_n9674_));
  AOI21_X1   g09379(.A1(new_n9332_), .A2(new_n9674_), .B(new_n9327_), .ZN(new_n9675_));
  INV_X1     g09380(.I(new_n9675_), .ZN(new_n9676_));
  INV_X1     g09381(.I(new_n9319_), .ZN(new_n9677_));
  AOI21_X1   g09382(.A1(new_n9322_), .A2(new_n9677_), .B(new_n9318_), .ZN(new_n9678_));
  INV_X1     g09383(.I(new_n9678_), .ZN(new_n9679_));
  INV_X1     g09384(.I(new_n9355_), .ZN(new_n9680_));
  AOI21_X1   g09385(.A1(new_n2277_), .A2(new_n6024_), .B(new_n9361_), .ZN(new_n9681_));
  INV_X1     g09386(.I(new_n9681_), .ZN(new_n9682_));
  XOR2_X1    g09387(.A1(new_n9303_), .A2(new_n9682_), .Z(new_n9683_));
  NOR2_X1    g09388(.A1(new_n9304_), .A2(new_n9682_), .ZN(new_n9684_));
  NOR2_X1    g09389(.A1(new_n9303_), .A2(new_n9681_), .ZN(new_n9685_));
  OAI21_X1   g09390(.A1(new_n9684_), .A2(new_n9685_), .B(new_n9680_), .ZN(new_n9686_));
  OAI21_X1   g09391(.A1(new_n9680_), .A2(new_n9683_), .B(new_n9686_), .ZN(new_n9687_));
  NAND3_X1   g09392(.A1(new_n1722_), .A2(\a[48] ), .A3(\a[56] ), .ZN(new_n9688_));
  AOI21_X1   g09393(.A1(\a[48] ), .A2(\a[56] ), .B(new_n1722_), .ZN(new_n9689_));
  NOR2_X1    g09394(.A1(\a[26] ), .A2(\a[38] ), .ZN(new_n9690_));
  AOI21_X1   g09395(.A1(new_n9688_), .A2(new_n9690_), .B(new_n9689_), .ZN(new_n9691_));
  AOI21_X1   g09396(.A1(new_n267_), .A2(new_n8991_), .B(new_n9395_), .ZN(new_n9692_));
  AOI21_X1   g09397(.A1(new_n2331_), .A2(new_n9398_), .B(new_n5488_), .ZN(new_n9693_));
  XOR2_X1    g09398(.A1(new_n9692_), .A2(new_n9693_), .Z(new_n9694_));
  INV_X1     g09399(.I(new_n9694_), .ZN(new_n9695_));
  INV_X1     g09400(.I(new_n9692_), .ZN(new_n9696_));
  NOR2_X1    g09401(.A1(new_n9696_), .A2(new_n9693_), .ZN(new_n9697_));
  INV_X1     g09402(.I(new_n9697_), .ZN(new_n9698_));
  NAND2_X1   g09403(.A1(new_n9696_), .A2(new_n9693_), .ZN(new_n9699_));
  AOI21_X1   g09404(.A1(new_n9698_), .A2(new_n9699_), .B(new_n9691_), .ZN(new_n9700_));
  AOI21_X1   g09405(.A1(new_n9691_), .A2(new_n9695_), .B(new_n9700_), .ZN(new_n9701_));
  XNOR2_X1   g09406(.A1(new_n9687_), .A2(new_n9701_), .ZN(new_n9702_));
  NAND2_X1   g09407(.A1(new_n9702_), .A2(new_n9679_), .ZN(new_n9703_));
  INV_X1     g09408(.I(new_n9687_), .ZN(new_n9704_));
  NOR2_X1    g09409(.A1(new_n9704_), .A2(new_n9701_), .ZN(new_n9705_));
  NAND2_X1   g09410(.A1(new_n9704_), .A2(new_n9701_), .ZN(new_n9706_));
  INV_X1     g09411(.I(new_n9706_), .ZN(new_n9707_));
  OAI21_X1   g09412(.A1(new_n9707_), .A2(new_n9705_), .B(new_n9678_), .ZN(new_n9708_));
  NAND2_X1   g09413(.A1(new_n9708_), .A2(new_n9703_), .ZN(new_n9709_));
  XOR2_X1    g09414(.A1(new_n9709_), .A2(new_n9676_), .Z(new_n9710_));
  AOI21_X1   g09415(.A1(new_n9703_), .A2(new_n9708_), .B(new_n9676_), .ZN(new_n9711_));
  NOR2_X1    g09416(.A1(new_n9709_), .A2(new_n9675_), .ZN(new_n9712_));
  NOR2_X1    g09417(.A1(new_n9712_), .A2(new_n9711_), .ZN(new_n9713_));
  MUX2_X1    g09418(.I0(new_n9713_), .I1(new_n9710_), .S(new_n9673_), .Z(new_n9714_));
  XOR2_X1    g09419(.A1(new_n9714_), .A2(new_n9671_), .Z(new_n9715_));
  NOR2_X1    g09420(.A1(new_n9715_), .A2(new_n9669_), .ZN(new_n9716_));
  INV_X1     g09421(.I(new_n9671_), .ZN(new_n9717_));
  NOR2_X1    g09422(.A1(new_n9717_), .A2(new_n9714_), .ZN(new_n9718_));
  INV_X1     g09423(.I(new_n9718_), .ZN(new_n9719_));
  NAND2_X1   g09424(.A1(new_n9717_), .A2(new_n9714_), .ZN(new_n9720_));
  NAND2_X1   g09425(.A1(new_n9719_), .A2(new_n9720_), .ZN(new_n9721_));
  AOI21_X1   g09426(.A1(new_n9669_), .A2(new_n9721_), .B(new_n9716_), .ZN(new_n9722_));
  XNOR2_X1   g09427(.A1(new_n9668_), .A2(new_n9722_), .ZN(new_n9723_));
  NOR2_X1    g09428(.A1(new_n9666_), .A2(new_n9723_), .ZN(new_n9724_));
  NOR2_X1    g09429(.A1(new_n9668_), .A2(new_n9722_), .ZN(new_n9725_));
  NAND2_X1   g09430(.A1(new_n9668_), .A2(new_n9722_), .ZN(new_n9726_));
  INV_X1     g09431(.I(new_n9726_), .ZN(new_n9727_));
  NOR2_X1    g09432(.A1(new_n9727_), .A2(new_n9725_), .ZN(new_n9728_));
  INV_X1     g09433(.I(new_n9728_), .ZN(new_n9729_));
  AOI21_X1   g09434(.A1(new_n9666_), .A2(new_n9729_), .B(new_n9724_), .ZN(new_n9730_));
  INV_X1     g09435(.I(new_n9730_), .ZN(new_n9731_));
  OAI21_X1   g09436(.A1(new_n9206_), .A2(new_n9452_), .B(new_n9454_), .ZN(new_n9732_));
  NAND2_X1   g09437(.A1(new_n9731_), .A2(new_n9732_), .ZN(new_n9733_));
  XOR2_X1    g09438(.A1(new_n9468_), .A2(new_n9733_), .Z(new_n9734_));
  XOR2_X1    g09439(.A1(new_n9734_), .A2(new_n9460_), .Z(\asquared[66] ));
  NOR2_X1    g09440(.A1(new_n9460_), .A2(new_n9730_), .ZN(new_n9736_));
  OAI21_X1   g09441(.A1(new_n9461_), .A2(new_n9731_), .B(new_n9732_), .ZN(new_n9737_));
  INV_X1     g09442(.I(new_n9737_), .ZN(new_n9738_));
  AOI21_X1   g09443(.A1(new_n9468_), .A2(new_n9738_), .B(new_n9736_), .ZN(new_n9739_));
  OAI21_X1   g09444(.A1(new_n9666_), .A2(new_n9725_), .B(new_n9726_), .ZN(new_n9740_));
  INV_X1     g09445(.I(new_n9740_), .ZN(new_n9741_));
  AOI21_X1   g09446(.A1(new_n9663_), .A2(new_n9661_), .B(new_n9659_), .ZN(new_n9742_));
  INV_X1     g09447(.I(new_n9742_), .ZN(new_n9743_));
  OAI21_X1   g09448(.A1(new_n9669_), .A2(new_n9718_), .B(new_n9720_), .ZN(new_n9744_));
  INV_X1     g09449(.I(new_n9744_), .ZN(new_n9745_));
  NAND2_X1   g09450(.A1(new_n9579_), .A2(new_n9471_), .ZN(new_n9746_));
  NAND2_X1   g09451(.A1(new_n9746_), .A2(new_n9578_), .ZN(new_n9747_));
  INV_X1     g09452(.I(new_n9711_), .ZN(new_n9748_));
  AOI21_X1   g09453(.A1(new_n9748_), .A2(new_n9673_), .B(new_n9712_), .ZN(new_n9749_));
  OAI21_X1   g09454(.A1(new_n9678_), .A2(new_n9705_), .B(new_n9706_), .ZN(new_n9750_));
  INV_X1     g09455(.I(new_n9750_), .ZN(new_n9751_));
  NAND2_X1   g09456(.A1(new_n9606_), .A2(new_n9602_), .ZN(new_n9752_));
  NAND2_X1   g09457(.A1(new_n9752_), .A2(new_n9605_), .ZN(new_n9753_));
  NOR2_X1    g09458(.A1(new_n9685_), .A2(new_n9680_), .ZN(new_n9754_));
  NOR2_X1    g09459(.A1(new_n9754_), .A2(new_n9684_), .ZN(new_n9755_));
  NAND2_X1   g09460(.A1(new_n9699_), .A2(new_n9691_), .ZN(new_n9756_));
  NAND2_X1   g09461(.A1(new_n9756_), .A2(new_n9698_), .ZN(new_n9757_));
  NAND2_X1   g09462(.A1(new_n9595_), .A2(new_n9586_), .ZN(new_n9758_));
  NAND2_X1   g09463(.A1(new_n9758_), .A2(new_n9594_), .ZN(new_n9759_));
  XNOR2_X1   g09464(.A1(new_n9759_), .A2(new_n9757_), .ZN(new_n9760_));
  AOI22_X1   g09465(.A1(new_n9758_), .A2(new_n9594_), .B1(new_n9756_), .B2(new_n9698_), .ZN(new_n9761_));
  NOR2_X1    g09466(.A1(new_n9759_), .A2(new_n9757_), .ZN(new_n9762_));
  OAI21_X1   g09467(.A1(new_n9761_), .A2(new_n9762_), .B(new_n9755_), .ZN(new_n9763_));
  OAI21_X1   g09468(.A1(new_n9755_), .A2(new_n9760_), .B(new_n9763_), .ZN(new_n9764_));
  XOR2_X1    g09469(.A1(new_n9753_), .A2(new_n9764_), .Z(new_n9765_));
  NOR2_X1    g09470(.A1(new_n9765_), .A2(new_n9751_), .ZN(new_n9766_));
  INV_X1     g09471(.I(new_n9764_), .ZN(new_n9767_));
  NOR2_X1    g09472(.A1(new_n9753_), .A2(new_n9767_), .ZN(new_n9768_));
  INV_X1     g09473(.I(new_n9768_), .ZN(new_n9769_));
  NAND2_X1   g09474(.A1(new_n9753_), .A2(new_n9767_), .ZN(new_n9770_));
  AOI21_X1   g09475(.A1(new_n9769_), .A2(new_n9770_), .B(new_n9750_), .ZN(new_n9771_));
  NOR2_X1    g09476(.A1(new_n9766_), .A2(new_n9771_), .ZN(new_n9772_));
  NOR4_X1    g09477(.A1(new_n566_), .A2(new_n1339_), .A3(new_n5511_), .A4(new_n6945_), .ZN(new_n9773_));
  NOR3_X1    g09478(.A1(new_n7700_), .A2(new_n1339_), .A3(new_n6999_), .ZN(new_n9774_));
  NAND2_X1   g09479(.A1(new_n9774_), .A2(new_n9773_), .ZN(new_n9775_));
  AOI21_X1   g09480(.A1(new_n9775_), .A2(new_n8005_), .B(new_n651_), .ZN(new_n9776_));
  NOR3_X1    g09481(.A1(new_n9776_), .A2(new_n675_), .A3(new_n6999_), .ZN(new_n9777_));
  NOR2_X1    g09482(.A1(new_n9776_), .A2(new_n9773_), .ZN(new_n9778_));
  AOI22_X1   g09483(.A1(\a[12] ), .A2(\a[19] ), .B1(\a[47] ), .B2(\a[54] ), .ZN(new_n9779_));
  AOI21_X1   g09484(.A1(new_n9778_), .A2(new_n9779_), .B(new_n9777_), .ZN(new_n9780_));
  NOR2_X1    g09485(.A1(new_n8453_), .A2(new_n9310_), .ZN(new_n9781_));
  AOI22_X1   g09486(.A1(new_n267_), .A2(new_n9781_), .B1(new_n9549_), .B2(new_n317_), .ZN(new_n9782_));
  INV_X1     g09487(.I(new_n9782_), .ZN(new_n9783_));
  NOR2_X1    g09488(.A1(new_n8453_), .A2(new_n9029_), .ZN(new_n9784_));
  INV_X1     g09489(.I(new_n9784_), .ZN(new_n9785_));
  NAND4_X1   g09490(.A1(new_n9785_), .A2(\a[3] ), .A3(\a[63] ), .A4(new_n211_), .ZN(new_n9786_));
  AOI21_X1   g09491(.A1(new_n5339_), .A2(new_n5601_), .B(new_n9042_), .ZN(new_n9787_));
  NOR4_X1    g09492(.A1(new_n2690_), .A2(new_n5600_), .A3(new_n2098_), .A4(new_n3783_), .ZN(new_n9788_));
  NAND2_X1   g09493(.A1(new_n9787_), .A2(new_n9788_), .ZN(new_n9789_));
  NOR3_X1    g09494(.A1(new_n9789_), .A2(new_n9783_), .A3(new_n9786_), .ZN(new_n9790_));
  NOR2_X1    g09495(.A1(new_n9783_), .A2(new_n9786_), .ZN(new_n9791_));
  INV_X1     g09496(.I(new_n9789_), .ZN(new_n9792_));
  NOR2_X1    g09497(.A1(new_n9792_), .A2(new_n9791_), .ZN(new_n9793_));
  OAI21_X1   g09498(.A1(new_n9790_), .A2(new_n9793_), .B(new_n9780_), .ZN(new_n9794_));
  XOR2_X1    g09499(.A1(new_n9789_), .A2(new_n9791_), .Z(new_n9795_));
  OAI21_X1   g09500(.A1(new_n9780_), .A2(new_n9795_), .B(new_n9794_), .ZN(new_n9796_));
  NAND2_X1   g09501(.A1(\a[23] ), .A2(\a[43] ), .ZN(new_n9797_));
  NOR2_X1    g09502(.A1(new_n1691_), .A2(new_n7727_), .ZN(new_n9798_));
  INV_X1     g09503(.I(new_n9798_), .ZN(new_n9799_));
  NOR2_X1    g09504(.A1(new_n7141_), .A2(new_n9799_), .ZN(new_n9800_));
  NOR4_X1    g09505(.A1(new_n364_), .A2(new_n1691_), .A3(new_n4769_), .A4(new_n7727_), .ZN(new_n9805_));
  INV_X1     g09506(.I(new_n9805_), .ZN(new_n9806_));
  AOI22_X1   g09507(.A1(new_n2978_), .A2(new_n7452_), .B1(new_n5488_), .B2(new_n4437_), .ZN(new_n9807_));
  NOR4_X1    g09508(.A1(new_n5742_), .A2(new_n4538_), .A3(new_n1215_), .A4(new_n5175_), .ZN(new_n9808_));
  NAND2_X1   g09509(.A1(new_n9807_), .A2(new_n9808_), .ZN(new_n9809_));
  NAND2_X1   g09510(.A1(new_n2752_), .A2(new_n5592_), .ZN(new_n9810_));
  NOR2_X1    g09511(.A1(new_n461_), .A2(new_n7216_), .ZN(new_n9811_));
  XOR2_X1    g09512(.A1(new_n9810_), .A2(new_n9811_), .Z(new_n9812_));
  NOR2_X1    g09513(.A1(new_n9812_), .A2(new_n9809_), .ZN(new_n9813_));
  INV_X1     g09514(.I(new_n9813_), .ZN(new_n9814_));
  NAND2_X1   g09515(.A1(new_n9812_), .A2(new_n9809_), .ZN(new_n9815_));
  AOI21_X1   g09516(.A1(new_n9814_), .A2(new_n9815_), .B(new_n9806_), .ZN(new_n9816_));
  XNOR2_X1   g09517(.A1(new_n9812_), .A2(new_n9809_), .ZN(new_n9817_));
  NOR2_X1    g09518(.A1(new_n9817_), .A2(new_n9805_), .ZN(new_n9818_));
  NOR2_X1    g09519(.A1(new_n9818_), .A2(new_n9816_), .ZN(new_n9819_));
  NAND2_X1   g09520(.A1(new_n7000_), .A2(new_n2328_), .ZN(new_n9820_));
  NAND2_X1   g09521(.A1(\a[18] ), .A2(\a[48] ), .ZN(new_n9821_));
  XNOR2_X1   g09522(.A1(new_n9820_), .A2(new_n9821_), .ZN(new_n9822_));
  NAND2_X1   g09523(.A1(new_n3126_), .A2(new_n3966_), .ZN(new_n9823_));
  NAND2_X1   g09524(.A1(\a[14] ), .A2(\a[52] ), .ZN(new_n9824_));
  XNOR2_X1   g09525(.A1(new_n9823_), .A2(new_n9824_), .ZN(new_n9825_));
  NAND2_X1   g09526(.A1(\a[49] ), .A2(\a[50] ), .ZN(new_n9826_));
  XNOR2_X1   g09527(.A1(new_n1274_), .A2(new_n9826_), .ZN(new_n9827_));
  NOR2_X1    g09528(.A1(new_n9825_), .A2(new_n9827_), .ZN(new_n9828_));
  AND2_X2    g09529(.A1(new_n9825_), .A2(new_n9827_), .Z(new_n9829_));
  NOR2_X1    g09530(.A1(new_n9829_), .A2(new_n9828_), .ZN(new_n9830_));
  NOR2_X1    g09531(.A1(new_n9830_), .A2(new_n9822_), .ZN(new_n9831_));
  INV_X1     g09532(.I(new_n9822_), .ZN(new_n9832_));
  XNOR2_X1   g09533(.A1(new_n9825_), .A2(new_n9827_), .ZN(new_n9833_));
  NOR2_X1    g09534(.A1(new_n9833_), .A2(new_n9832_), .ZN(new_n9834_));
  NOR2_X1    g09535(.A1(new_n9831_), .A2(new_n9834_), .ZN(new_n9835_));
  XOR2_X1    g09536(.A1(new_n9835_), .A2(new_n9819_), .Z(new_n9836_));
  AND2_X2    g09537(.A1(new_n9836_), .A2(new_n9796_), .Z(new_n9837_));
  OAI22_X1   g09538(.A1(new_n9831_), .A2(new_n9834_), .B1(new_n9818_), .B2(new_n9816_), .ZN(new_n9838_));
  NAND2_X1   g09539(.A1(new_n9835_), .A2(new_n9819_), .ZN(new_n9839_));
  AOI21_X1   g09540(.A1(new_n9838_), .A2(new_n9839_), .B(new_n9796_), .ZN(new_n9840_));
  NOR2_X1    g09541(.A1(new_n9837_), .A2(new_n9840_), .ZN(new_n9841_));
  XNOR2_X1   g09542(.A1(new_n9772_), .A2(new_n9841_), .ZN(new_n9842_));
  NOR2_X1    g09543(.A1(new_n9842_), .A2(new_n9749_), .ZN(new_n9843_));
  NOR2_X1    g09544(.A1(new_n9772_), .A2(new_n9841_), .ZN(new_n9844_));
  INV_X1     g09545(.I(new_n9844_), .ZN(new_n9845_));
  NAND2_X1   g09546(.A1(new_n9772_), .A2(new_n9841_), .ZN(new_n9846_));
  NAND2_X1   g09547(.A1(new_n9845_), .A2(new_n9846_), .ZN(new_n9847_));
  AOI21_X1   g09548(.A1(new_n9749_), .A2(new_n9847_), .B(new_n9843_), .ZN(new_n9848_));
  XNOR2_X1   g09549(.A1(new_n9747_), .A2(new_n9848_), .ZN(new_n9849_));
  NOR2_X1    g09550(.A1(new_n9849_), .A2(new_n9745_), .ZN(new_n9850_));
  NOR2_X1    g09551(.A1(new_n9747_), .A2(new_n9848_), .ZN(new_n9851_));
  INV_X1     g09552(.I(new_n9851_), .ZN(new_n9852_));
  NAND2_X1   g09553(.A1(new_n9747_), .A2(new_n9848_), .ZN(new_n9853_));
  AOI21_X1   g09554(.A1(new_n9852_), .A2(new_n9853_), .B(new_n9744_), .ZN(new_n9854_));
  NOR2_X1    g09555(.A1(new_n9850_), .A2(new_n9854_), .ZN(new_n9855_));
  INV_X1     g09556(.I(new_n9855_), .ZN(new_n9856_));
  NAND2_X1   g09557(.A1(new_n9495_), .A2(new_n9472_), .ZN(new_n9857_));
  NAND2_X1   g09558(.A1(new_n9857_), .A2(new_n9494_), .ZN(new_n9858_));
  AOI21_X1   g09559(.A1(new_n9482_), .A2(new_n9485_), .B(new_n9483_), .ZN(new_n9859_));
  INV_X1     g09560(.I(new_n9859_), .ZN(new_n9860_));
  INV_X1     g09561(.I(new_n9781_), .ZN(new_n9861_));
  NOR2_X1    g09562(.A1(new_n9861_), .A2(new_n260_), .ZN(new_n9862_));
  AOI21_X1   g09563(.A1(new_n2797_), .A2(new_n5600_), .B(new_n9513_), .ZN(new_n9863_));
  NOR2_X1    g09564(.A1(new_n9556_), .A2(new_n3039_), .ZN(new_n9864_));
  NOR4_X1    g09565(.A1(new_n8676_), .A2(new_n609_), .A3(new_n242_), .A4(new_n8990_), .ZN(new_n9865_));
  AND2_X2    g09566(.A1(new_n9864_), .A2(new_n9865_), .Z(new_n9866_));
  NAND2_X1   g09567(.A1(new_n9866_), .A2(new_n9863_), .ZN(new_n9867_));
  XOR2_X1    g09568(.A1(new_n9867_), .A2(new_n9618_), .Z(new_n9868_));
  XOR2_X1    g09569(.A1(new_n9868_), .A2(new_n9862_), .Z(new_n9869_));
  INV_X1     g09570(.I(new_n9635_), .ZN(new_n9870_));
  AOI21_X1   g09571(.A1(new_n9638_), .A2(new_n9870_), .B(new_n9634_), .ZN(new_n9871_));
  XOR2_X1    g09572(.A1(new_n9869_), .A2(new_n9871_), .Z(new_n9872_));
  NOR2_X1    g09573(.A1(new_n9869_), .A2(new_n9871_), .ZN(new_n9873_));
  INV_X1     g09574(.I(new_n9873_), .ZN(new_n9874_));
  NAND2_X1   g09575(.A1(new_n9869_), .A2(new_n9871_), .ZN(new_n9875_));
  AOI21_X1   g09576(.A1(new_n9874_), .A2(new_n9875_), .B(new_n9860_), .ZN(new_n9876_));
  AOI21_X1   g09577(.A1(new_n9860_), .A2(new_n9872_), .B(new_n9876_), .ZN(new_n9877_));
  AOI21_X1   g09578(.A1(new_n1447_), .A2(new_n6779_), .B(new_n9630_), .ZN(new_n9878_));
  NOR2_X1    g09579(.A1(new_n9524_), .A2(new_n9525_), .ZN(new_n9879_));
  NOR2_X1    g09580(.A1(new_n200_), .A2(new_n9029_), .ZN(new_n9880_));
  OAI21_X1   g09581(.A1(\a[33] ), .A2(new_n9536_), .B(new_n9880_), .ZN(new_n9881_));
  NAND2_X1   g09582(.A1(new_n9881_), .A2(new_n9537_), .ZN(new_n9882_));
  INV_X1     g09583(.I(new_n9882_), .ZN(new_n9883_));
  XOR2_X1    g09584(.A1(new_n9879_), .A2(new_n9883_), .Z(new_n9884_));
  INV_X1     g09585(.I(new_n9884_), .ZN(new_n9885_));
  NOR3_X1    g09586(.A1(new_n9524_), .A2(new_n9883_), .A3(new_n9525_), .ZN(new_n9886_));
  INV_X1     g09587(.I(new_n9886_), .ZN(new_n9887_));
  NOR2_X1    g09588(.A1(new_n9879_), .A2(new_n9882_), .ZN(new_n9888_));
  INV_X1     g09589(.I(new_n9888_), .ZN(new_n9889_));
  AOI21_X1   g09590(.A1(new_n9889_), .A2(new_n9887_), .B(new_n9878_), .ZN(new_n9890_));
  AOI21_X1   g09591(.A1(new_n9885_), .A2(new_n9878_), .B(new_n9890_), .ZN(new_n9891_));
  NAND2_X1   g09592(.A1(new_n5321_), .A2(new_n4538_), .ZN(new_n9892_));
  NOR2_X1    g09593(.A1(new_n5321_), .A2(new_n4538_), .ZN(new_n9893_));
  NOR2_X1    g09594(.A1(\a[8] ), .A2(\a[57] ), .ZN(new_n9894_));
  AOI21_X1   g09595(.A1(new_n9892_), .A2(new_n9894_), .B(new_n9893_), .ZN(new_n9895_));
  INV_X1     g09596(.I(new_n9895_), .ZN(new_n9896_));
  AOI21_X1   g09597(.A1(new_n479_), .A2(new_n8676_), .B(new_n9557_), .ZN(new_n9897_));
  NOR2_X1    g09598(.A1(new_n675_), .A2(new_n6945_), .ZN(new_n9898_));
  OAI21_X1   g09599(.A1(new_n9529_), .A2(new_n9531_), .B(new_n9898_), .ZN(new_n9899_));
  OAI21_X1   g09600(.A1(new_n9530_), .A2(new_n9532_), .B(new_n9899_), .ZN(new_n9900_));
  INV_X1     g09601(.I(new_n9900_), .ZN(new_n9901_));
  XOR2_X1    g09602(.A1(new_n9897_), .A2(new_n9901_), .Z(new_n9902_));
  NOR2_X1    g09603(.A1(new_n9902_), .A2(new_n9896_), .ZN(new_n9903_));
  AND2_X2    g09604(.A1(new_n9897_), .A2(new_n9900_), .Z(new_n9904_));
  NOR2_X1    g09605(.A1(new_n9897_), .A2(new_n9900_), .ZN(new_n9905_));
  NOR2_X1    g09606(.A1(new_n9904_), .A2(new_n9905_), .ZN(new_n9906_));
  NOR2_X1    g09607(.A1(new_n9906_), .A2(new_n9895_), .ZN(new_n9907_));
  NOR2_X1    g09608(.A1(new_n9907_), .A2(new_n9903_), .ZN(new_n9908_));
  INV_X1     g09609(.I(new_n9908_), .ZN(new_n9909_));
  AND2_X2    g09610(.A1(new_n9541_), .A2(new_n9528_), .Z(new_n9910_));
  NOR2_X1    g09611(.A1(new_n9910_), .A2(new_n9540_), .ZN(new_n9911_));
  NOR2_X1    g09612(.A1(new_n9911_), .A2(new_n9909_), .ZN(new_n9912_));
  NOR3_X1    g09613(.A1(new_n9910_), .A2(new_n9908_), .A3(new_n9540_), .ZN(new_n9913_));
  NOR2_X1    g09614(.A1(new_n9912_), .A2(new_n9913_), .ZN(new_n9914_));
  NOR2_X1    g09615(.A1(new_n9914_), .A2(new_n9891_), .ZN(new_n9915_));
  XOR2_X1    g09616(.A1(new_n9911_), .A2(new_n9908_), .Z(new_n9916_));
  INV_X1     g09617(.I(new_n9916_), .ZN(new_n9917_));
  AOI21_X1   g09618(.A1(new_n9891_), .A2(new_n9917_), .B(new_n9915_), .ZN(new_n9918_));
  XOR2_X1    g09619(.A1(new_n9918_), .A2(new_n9877_), .Z(new_n9919_));
  NOR2_X1    g09620(.A1(new_n9918_), .A2(new_n9877_), .ZN(new_n9920_));
  INV_X1     g09621(.I(new_n9920_), .ZN(new_n9921_));
  NAND2_X1   g09622(.A1(new_n9918_), .A2(new_n9877_), .ZN(new_n9922_));
  AOI21_X1   g09623(.A1(new_n9921_), .A2(new_n9922_), .B(new_n9858_), .ZN(new_n9923_));
  AOI21_X1   g09624(.A1(new_n9858_), .A2(new_n9919_), .B(new_n9923_), .ZN(new_n9924_));
  NAND2_X1   g09625(.A1(new_n9656_), .A2(new_n9608_), .ZN(new_n9925_));
  NAND2_X1   g09626(.A1(new_n9925_), .A2(new_n9655_), .ZN(new_n9926_));
  INV_X1     g09627(.I(new_n9518_), .ZN(new_n9927_));
  AOI21_X1   g09628(.A1(new_n9509_), .A2(new_n9927_), .B(new_n9515_), .ZN(new_n9928_));
  NOR2_X1    g09629(.A1(new_n9624_), .A2(new_n9621_), .ZN(new_n9929_));
  AOI21_X1   g09630(.A1(new_n2277_), .A2(new_n5592_), .B(new_n9510_), .ZN(new_n9930_));
  XOR2_X1    g09631(.A1(new_n9929_), .A2(new_n9930_), .Z(new_n9931_));
  INV_X1     g09632(.I(new_n9930_), .ZN(new_n9932_));
  NOR3_X1    g09633(.A1(new_n9624_), .A2(new_n9932_), .A3(new_n9621_), .ZN(new_n9933_));
  NOR2_X1    g09634(.A1(new_n9929_), .A2(new_n9930_), .ZN(new_n9934_));
  NOR2_X1    g09635(.A1(new_n9934_), .A2(new_n9933_), .ZN(new_n9935_));
  NOR2_X1    g09636(.A1(new_n9935_), .A2(new_n9506_), .ZN(new_n9936_));
  AOI21_X1   g09637(.A1(new_n9506_), .A2(new_n9931_), .B(new_n9936_), .ZN(new_n9937_));
  INV_X1     g09638(.I(new_n9566_), .ZN(new_n9938_));
  AOI21_X1   g09639(.A1(new_n9562_), .A2(new_n9938_), .B(new_n9565_), .ZN(new_n9939_));
  XOR2_X1    g09640(.A1(new_n9937_), .A2(new_n9939_), .Z(new_n9940_));
  NOR2_X1    g09641(.A1(new_n9940_), .A2(new_n9928_), .ZN(new_n9941_));
  XOR2_X1    g09642(.A1(new_n9937_), .A2(new_n9939_), .Z(new_n9942_));
  AOI21_X1   g09643(.A1(new_n9928_), .A2(new_n9942_), .B(new_n9941_), .ZN(new_n9943_));
  INV_X1     g09644(.I(new_n9943_), .ZN(new_n9944_));
  OAI21_X1   g09645(.A1(new_n9522_), .A2(new_n9570_), .B(new_n9572_), .ZN(new_n9945_));
  INV_X1     g09646(.I(new_n9945_), .ZN(new_n9946_));
  NOR2_X1    g09647(.A1(new_n9645_), .A2(new_n9612_), .ZN(new_n9947_));
  NOR2_X1    g09648(.A1(new_n9947_), .A2(new_n9643_), .ZN(new_n9948_));
  NOR2_X1    g09649(.A1(new_n9946_), .A2(new_n9948_), .ZN(new_n9949_));
  NAND2_X1   g09650(.A1(new_n9946_), .A2(new_n9948_), .ZN(new_n9950_));
  INV_X1     g09651(.I(new_n9950_), .ZN(new_n9951_));
  OAI21_X1   g09652(.A1(new_n9951_), .A2(new_n9949_), .B(new_n9944_), .ZN(new_n9952_));
  XNOR2_X1   g09653(.A1(new_n9945_), .A2(new_n9948_), .ZN(new_n9953_));
  NAND2_X1   g09654(.A1(new_n9953_), .A2(new_n9943_), .ZN(new_n9954_));
  NAND2_X1   g09655(.A1(new_n9952_), .A2(new_n9954_), .ZN(new_n9955_));
  XOR2_X1    g09656(.A1(new_n9926_), .A2(new_n9955_), .Z(new_n9956_));
  NOR2_X1    g09657(.A1(new_n9956_), .A2(new_n9924_), .ZN(new_n9957_));
  NAND3_X1   g09658(.A1(new_n9955_), .A2(new_n9655_), .A3(new_n9925_), .ZN(new_n9958_));
  NAND3_X1   g09659(.A1(new_n9926_), .A2(new_n9952_), .A3(new_n9954_), .ZN(new_n9959_));
  NAND2_X1   g09660(.A1(new_n9959_), .A2(new_n9958_), .ZN(new_n9960_));
  AOI21_X1   g09661(.A1(new_n9924_), .A2(new_n9960_), .B(new_n9957_), .ZN(new_n9961_));
  NOR2_X1    g09662(.A1(new_n9856_), .A2(new_n9961_), .ZN(new_n9962_));
  INV_X1     g09663(.I(new_n9961_), .ZN(new_n9963_));
  NOR2_X1    g09664(.A1(new_n9855_), .A2(new_n9963_), .ZN(new_n9964_));
  OAI21_X1   g09665(.A1(new_n9962_), .A2(new_n9964_), .B(new_n9743_), .ZN(new_n9965_));
  XOR2_X1    g09666(.A1(new_n9855_), .A2(new_n9961_), .Z(new_n9966_));
  OAI21_X1   g09667(.A1(new_n9743_), .A2(new_n9966_), .B(new_n9965_), .ZN(new_n9967_));
  XOR2_X1    g09668(.A1(new_n9967_), .A2(new_n9741_), .Z(new_n9968_));
  NAND2_X1   g09669(.A1(new_n9967_), .A2(new_n9740_), .ZN(new_n9969_));
  INV_X1     g09670(.I(new_n9967_), .ZN(new_n9970_));
  NAND2_X1   g09671(.A1(new_n9970_), .A2(new_n9741_), .ZN(new_n9971_));
  NAND2_X1   g09672(.A1(new_n9971_), .A2(new_n9969_), .ZN(new_n9972_));
  NAND2_X1   g09673(.A1(new_n9739_), .A2(new_n9972_), .ZN(new_n9973_));
  OAI21_X1   g09674(.A1(new_n9739_), .A2(new_n9968_), .B(new_n9973_), .ZN(\asquared[67] ));
  NOR2_X1    g09675(.A1(new_n9967_), .A2(new_n9740_), .ZN(new_n9975_));
  OAI21_X1   g09676(.A1(new_n9739_), .A2(new_n9975_), .B(new_n9969_), .ZN(new_n9976_));
  INV_X1     g09677(.I(new_n9962_), .ZN(new_n9977_));
  OAI21_X1   g09678(.A1(new_n9742_), .A2(new_n9964_), .B(new_n9977_), .ZN(new_n9978_));
  AOI21_X1   g09679(.A1(new_n9943_), .A2(new_n9950_), .B(new_n9949_), .ZN(new_n9979_));
  INV_X1     g09680(.I(new_n9939_), .ZN(new_n9980_));
  NAND2_X1   g09681(.A1(new_n9937_), .A2(new_n9980_), .ZN(new_n9981_));
  NOR2_X1    g09682(.A1(new_n9937_), .A2(new_n9980_), .ZN(new_n9982_));
  OAI21_X1   g09683(.A1(new_n9928_), .A2(new_n9982_), .B(new_n9981_), .ZN(new_n9983_));
  NOR3_X1    g09684(.A1(new_n9934_), .A2(new_n9501_), .A3(new_n9504_), .ZN(new_n9984_));
  NOR2_X1    g09685(.A1(new_n9984_), .A2(new_n9933_), .ZN(new_n9985_));
  INV_X1     g09686(.I(new_n9904_), .ZN(new_n9986_));
  OAI21_X1   g09687(.A1(new_n9896_), .A2(new_n9905_), .B(new_n9986_), .ZN(new_n9987_));
  NAND2_X1   g09688(.A1(new_n9889_), .A2(new_n9878_), .ZN(new_n9988_));
  NAND2_X1   g09689(.A1(new_n9988_), .A2(new_n9887_), .ZN(new_n9989_));
  XNOR2_X1   g09690(.A1(new_n9987_), .A2(new_n9989_), .ZN(new_n9990_));
  NOR2_X1    g09691(.A1(new_n9990_), .A2(new_n9985_), .ZN(new_n9991_));
  INV_X1     g09692(.I(new_n9985_), .ZN(new_n9992_));
  NAND2_X1   g09693(.A1(new_n9987_), .A2(new_n9989_), .ZN(new_n9993_));
  NOR2_X1    g09694(.A1(new_n9987_), .A2(new_n9989_), .ZN(new_n9994_));
  INV_X1     g09695(.I(new_n9994_), .ZN(new_n9995_));
  AOI21_X1   g09696(.A1(new_n9995_), .A2(new_n9993_), .B(new_n9992_), .ZN(new_n9996_));
  NOR2_X1    g09697(.A1(new_n9991_), .A2(new_n9996_), .ZN(new_n9997_));
  INV_X1     g09698(.I(new_n9913_), .ZN(new_n9998_));
  AOI21_X1   g09699(.A1(new_n9998_), .A2(new_n9891_), .B(new_n9912_), .ZN(new_n9999_));
  XOR2_X1    g09700(.A1(new_n9997_), .A2(new_n9999_), .Z(new_n10000_));
  INV_X1     g09701(.I(new_n10000_), .ZN(new_n10001_));
  INV_X1     g09702(.I(new_n9997_), .ZN(new_n10002_));
  NOR2_X1    g09703(.A1(new_n10002_), .A2(new_n9999_), .ZN(new_n10003_));
  INV_X1     g09704(.I(new_n10003_), .ZN(new_n10004_));
  NAND2_X1   g09705(.A1(new_n10002_), .A2(new_n9999_), .ZN(new_n10005_));
  AOI21_X1   g09706(.A1(new_n10004_), .A2(new_n10005_), .B(new_n9983_), .ZN(new_n10006_));
  AOI21_X1   g09707(.A1(new_n10001_), .A2(new_n9983_), .B(new_n10006_), .ZN(new_n10007_));
  NOR2_X1    g09708(.A1(new_n5750_), .A2(new_n6694_), .ZN(new_n10008_));
  NAND2_X1   g09709(.A1(new_n2684_), .A2(new_n1339_), .ZN(new_n10009_));
  AOI21_X1   g09710(.A1(new_n6056_), .A2(new_n10008_), .B(new_n10009_), .ZN(new_n10010_));
  NAND2_X1   g09711(.A1(\a[14] ), .A2(\a[53] ), .ZN(new_n10011_));
  NAND2_X1   g09712(.A1(\a[19] ), .A2(\a[48] ), .ZN(new_n10012_));
  NOR4_X1    g09713(.A1(new_n10010_), .A2(new_n7174_), .A3(new_n10011_), .A4(new_n10012_), .ZN(new_n10013_));
  NAND2_X1   g09714(.A1(\a[21] ), .A2(\a[42] ), .ZN(new_n10014_));
  NOR3_X1    g09715(.A1(new_n10014_), .A2(new_n1999_), .A3(new_n5175_), .ZN(new_n10015_));
  AOI21_X1   g09716(.A1(new_n2752_), .A2(new_n5350_), .B(new_n10015_), .ZN(new_n10016_));
  NOR2_X1    g09717(.A1(new_n1313_), .A2(new_n5175_), .ZN(new_n10017_));
  NOR2_X1    g09718(.A1(new_n1916_), .A2(new_n4414_), .ZN(new_n10018_));
  XNOR2_X1   g09719(.A1(new_n10017_), .A2(new_n10018_), .ZN(new_n10019_));
  NOR2_X1    g09720(.A1(new_n10019_), .A2(new_n10017_), .ZN(new_n10020_));
  NOR2_X1    g09721(.A1(new_n10016_), .A2(new_n10020_), .ZN(new_n10021_));
  OAI21_X1   g09722(.A1(new_n1999_), .A2(new_n4769_), .B(new_n10019_), .ZN(new_n10022_));
  INV_X1     g09723(.I(new_n10022_), .ZN(new_n10023_));
  NOR2_X1    g09724(.A1(new_n10023_), .A2(new_n10021_), .ZN(new_n10024_));
  INV_X1     g09725(.I(new_n10024_), .ZN(new_n10025_));
  NAND2_X1   g09726(.A1(new_n2797_), .A2(new_n6024_), .ZN(new_n10026_));
  XNOR2_X1   g09727(.A1(new_n10026_), .A2(new_n9614_), .ZN(new_n10027_));
  NOR2_X1    g09728(.A1(new_n10025_), .A2(new_n10027_), .ZN(new_n10028_));
  INV_X1     g09729(.I(new_n10027_), .ZN(new_n10029_));
  NOR2_X1    g09730(.A1(new_n10024_), .A2(new_n10029_), .ZN(new_n10030_));
  OAI21_X1   g09731(.A1(new_n10028_), .A2(new_n10030_), .B(new_n10013_), .ZN(new_n10031_));
  XOR2_X1    g09732(.A1(new_n10024_), .A2(new_n10027_), .Z(new_n10032_));
  OAI21_X1   g09733(.A1(new_n10032_), .A2(new_n10013_), .B(new_n10031_), .ZN(new_n10033_));
  INV_X1     g09734(.I(new_n6777_), .ZN(new_n10034_));
  NAND3_X1   g09735(.A1(new_n4880_), .A2(\a[37] ), .A3(\a[52] ), .ZN(new_n10035_));
  OAI21_X1   g09736(.A1(new_n1021_), .A2(new_n10034_), .B(new_n10035_), .ZN(new_n10036_));
  NOR2_X1    g09737(.A1(new_n800_), .A2(new_n6260_), .ZN(new_n10037_));
  NOR2_X1    g09738(.A1(new_n2461_), .A2(new_n3837_), .ZN(new_n10038_));
  XNOR2_X1   g09739(.A1(new_n10037_), .A2(new_n10038_), .ZN(new_n10039_));
  OAI21_X1   g09740(.A1(new_n10039_), .A2(new_n10037_), .B(new_n10036_), .ZN(new_n10040_));
  OAI21_X1   g09741(.A1(new_n875_), .A2(new_n6692_), .B(new_n10039_), .ZN(new_n10041_));
  NAND2_X1   g09742(.A1(new_n10041_), .A2(new_n10040_), .ZN(new_n10042_));
  AOI22_X1   g09743(.A1(new_n1778_), .A2(new_n8996_), .B1(new_n9554_), .B2(new_n609_), .ZN(new_n10043_));
  INV_X1     g09744(.I(new_n10043_), .ZN(new_n10044_));
  NOR2_X1    g09745(.A1(new_n268_), .A2(new_n8990_), .ZN(new_n10045_));
  INV_X1     g09746(.I(new_n10045_), .ZN(new_n10046_));
  NOR4_X1    g09747(.A1(new_n10044_), .A2(new_n454_), .A3(new_n8676_), .A4(new_n10046_), .ZN(new_n10047_));
  INV_X1     g09748(.I(new_n10047_), .ZN(new_n10048_));
  NOR2_X1    g09749(.A1(new_n7188_), .A2(new_n8778_), .ZN(new_n10049_));
  NOR4_X1    g09750(.A1(new_n5321_), .A2(new_n2543_), .A3(new_n1674_), .A4(new_n5004_), .ZN(new_n10050_));
  NAND2_X1   g09751(.A1(new_n10049_), .A2(new_n10050_), .ZN(new_n10051_));
  NOR2_X1    g09752(.A1(new_n10048_), .A2(new_n10051_), .ZN(new_n10052_));
  AOI21_X1   g09753(.A1(new_n10049_), .A2(new_n10050_), .B(new_n10047_), .ZN(new_n10053_));
  NOR2_X1    g09754(.A1(new_n10052_), .A2(new_n10053_), .ZN(new_n10054_));
  NOR2_X1    g09755(.A1(new_n10054_), .A2(new_n10042_), .ZN(new_n10055_));
  INV_X1     g09756(.I(new_n10042_), .ZN(new_n10056_));
  XOR2_X1    g09757(.A1(new_n10051_), .A2(new_n10047_), .Z(new_n10057_));
  NOR2_X1    g09758(.A1(new_n10057_), .A2(new_n10056_), .ZN(new_n10058_));
  NOR2_X1    g09759(.A1(new_n10055_), .A2(new_n10058_), .ZN(new_n10059_));
  AOI21_X1   g09760(.A1(new_n3966_), .A2(new_n4359_), .B(new_n9525_), .ZN(new_n10060_));
  AOI21_X1   g09761(.A1(\a[32] ), .A2(\a[35] ), .B(new_n4372_), .ZN(new_n10061_));
  NOR3_X1    g09762(.A1(new_n9523_), .A2(new_n4360_), .A3(new_n10061_), .ZN(new_n10062_));
  AND2_X2    g09763(.A1(new_n10060_), .A2(new_n10062_), .Z(new_n10063_));
  NAND2_X1   g09764(.A1(new_n7483_), .A2(new_n1220_), .ZN(new_n10064_));
  NAND2_X1   g09765(.A1(\a[29] ), .A2(\a[38] ), .ZN(new_n10065_));
  XNOR2_X1   g09766(.A1(new_n10064_), .A2(new_n10065_), .ZN(new_n10066_));
  NOR2_X1    g09767(.A1(new_n6733_), .A2(new_n3371_), .ZN(new_n10067_));
  XOR2_X1    g09768(.A1(new_n10067_), .A2(new_n353_), .Z(new_n10068_));
  NOR2_X1    g09769(.A1(new_n10068_), .A2(\a[62] ), .ZN(new_n10069_));
  NAND2_X1   g09770(.A1(new_n10068_), .A2(\a[62] ), .ZN(new_n10070_));
  INV_X1     g09771(.I(new_n10070_), .ZN(new_n10071_));
  NOR2_X1    g09772(.A1(new_n10071_), .A2(new_n10069_), .ZN(new_n10072_));
  NOR2_X1    g09773(.A1(new_n10072_), .A2(new_n10066_), .ZN(new_n10073_));
  INV_X1     g09774(.I(new_n10073_), .ZN(new_n10074_));
  INV_X1     g09775(.I(new_n10066_), .ZN(new_n10075_));
  NOR3_X1    g09776(.A1(new_n10071_), .A2(new_n10075_), .A3(new_n10069_), .ZN(new_n10076_));
  INV_X1     g09777(.I(new_n10076_), .ZN(new_n10077_));
  NAND2_X1   g09778(.A1(new_n10074_), .A2(new_n10077_), .ZN(new_n10078_));
  XOR2_X1    g09779(.A1(new_n10072_), .A2(new_n10075_), .Z(new_n10079_));
  NOR2_X1    g09780(.A1(new_n10079_), .A2(new_n10063_), .ZN(new_n10080_));
  AOI21_X1   g09781(.A1(new_n10063_), .A2(new_n10078_), .B(new_n10080_), .ZN(new_n10081_));
  XOR2_X1    g09782(.A1(new_n10081_), .A2(new_n10059_), .Z(new_n10082_));
  AND2_X2    g09783(.A1(new_n10082_), .A2(new_n10033_), .Z(new_n10083_));
  NOR2_X1    g09784(.A1(new_n10081_), .A2(new_n10059_), .ZN(new_n10084_));
  INV_X1     g09785(.I(new_n10084_), .ZN(new_n10085_));
  NAND2_X1   g09786(.A1(new_n10081_), .A2(new_n10059_), .ZN(new_n10086_));
  AOI21_X1   g09787(.A1(new_n10085_), .A2(new_n10086_), .B(new_n10033_), .ZN(new_n10087_));
  NOR2_X1    g09788(.A1(new_n10083_), .A2(new_n10087_), .ZN(new_n10088_));
  XNOR2_X1   g09789(.A1(new_n10007_), .A2(new_n10088_), .ZN(new_n10089_));
  NOR2_X1    g09790(.A1(new_n10089_), .A2(new_n9979_), .ZN(new_n10090_));
  INV_X1     g09791(.I(new_n9979_), .ZN(new_n10091_));
  NOR2_X1    g09792(.A1(new_n10007_), .A2(new_n10088_), .ZN(new_n10092_));
  INV_X1     g09793(.I(new_n10092_), .ZN(new_n10093_));
  NAND2_X1   g09794(.A1(new_n10007_), .A2(new_n10088_), .ZN(new_n10094_));
  AOI21_X1   g09795(.A1(new_n10093_), .A2(new_n10094_), .B(new_n10091_), .ZN(new_n10095_));
  NOR2_X1    g09796(.A1(new_n10090_), .A2(new_n10095_), .ZN(new_n10096_));
  NAND2_X1   g09797(.A1(new_n9924_), .A2(new_n9958_), .ZN(new_n10097_));
  NAND2_X1   g09798(.A1(new_n10097_), .A2(new_n9959_), .ZN(new_n10098_));
  OAI21_X1   g09799(.A1(new_n9749_), .A2(new_n9844_), .B(new_n9846_), .ZN(new_n10099_));
  INV_X1     g09800(.I(new_n10099_), .ZN(new_n10100_));
  XOR2_X1    g09801(.A1(new_n10098_), .A2(new_n10100_), .Z(new_n10101_));
  OAI21_X1   g09802(.A1(new_n9745_), .A2(new_n9851_), .B(new_n9853_), .ZN(new_n10102_));
  NAND2_X1   g09803(.A1(new_n9921_), .A2(new_n9858_), .ZN(new_n10103_));
  AND2_X2    g09804(.A1(new_n10103_), .A2(new_n9922_), .Z(new_n10104_));
  OAI21_X1   g09805(.A1(new_n9751_), .A2(new_n9768_), .B(new_n9770_), .ZN(new_n10105_));
  INV_X1     g09806(.I(new_n9793_), .ZN(new_n10106_));
  AOI21_X1   g09807(.A1(new_n9780_), .A2(new_n10106_), .B(new_n9790_), .ZN(new_n10107_));
  NAND2_X1   g09808(.A1(new_n9815_), .A2(new_n9805_), .ZN(new_n10108_));
  NAND2_X1   g09809(.A1(new_n10108_), .A2(new_n9814_), .ZN(new_n10109_));
  INV_X1     g09810(.I(new_n9863_), .ZN(new_n10110_));
  NAND2_X1   g09811(.A1(new_n9866_), .A2(new_n9862_), .ZN(new_n10111_));
  AOI21_X1   g09812(.A1(new_n9619_), .A2(new_n10110_), .B(new_n10111_), .ZN(new_n10112_));
  AOI21_X1   g09813(.A1(new_n9618_), .A2(new_n9863_), .B(new_n10112_), .ZN(new_n10113_));
  XOR2_X1    g09814(.A1(new_n10113_), .A2(new_n10109_), .Z(new_n10114_));
  NOR2_X1    g09815(.A1(new_n10114_), .A2(new_n10107_), .ZN(new_n10115_));
  INV_X1     g09816(.I(new_n10107_), .ZN(new_n10116_));
  INV_X1     g09817(.I(new_n10109_), .ZN(new_n10117_));
  NOR2_X1    g09818(.A1(new_n10113_), .A2(new_n10117_), .ZN(new_n10118_));
  INV_X1     g09819(.I(new_n10118_), .ZN(new_n10119_));
  NAND2_X1   g09820(.A1(new_n10113_), .A2(new_n10117_), .ZN(new_n10120_));
  AOI21_X1   g09821(.A1(new_n10119_), .A2(new_n10120_), .B(new_n10116_), .ZN(new_n10121_));
  NOR2_X1    g09822(.A1(new_n10115_), .A2(new_n10121_), .ZN(new_n10122_));
  AOI21_X1   g09823(.A1(new_n2543_), .A2(new_n5173_), .B(new_n9800_), .ZN(new_n10123_));
  AOI21_X1   g09824(.A1(new_n4538_), .A2(new_n5742_), .B(new_n9807_), .ZN(new_n10124_));
  NAND2_X1   g09825(.A1(new_n2752_), .A2(new_n5592_), .ZN(new_n10125_));
  NOR2_X1    g09826(.A1(new_n2752_), .A2(new_n5592_), .ZN(new_n10126_));
  NOR2_X1    g09827(.A1(\a[10] ), .A2(\a[56] ), .ZN(new_n10127_));
  AOI21_X1   g09828(.A1(new_n10125_), .A2(new_n10127_), .B(new_n10126_), .ZN(new_n10128_));
  XNOR2_X1   g09829(.A1(new_n10124_), .A2(new_n10128_), .ZN(new_n10129_));
  INV_X1     g09830(.I(new_n10129_), .ZN(new_n10130_));
  INV_X1     g09831(.I(new_n10124_), .ZN(new_n10131_));
  INV_X1     g09832(.I(new_n10128_), .ZN(new_n10132_));
  NOR2_X1    g09833(.A1(new_n10131_), .A2(new_n10132_), .ZN(new_n10133_));
  NOR2_X1    g09834(.A1(new_n10124_), .A2(new_n10128_), .ZN(new_n10134_));
  NOR2_X1    g09835(.A1(new_n10133_), .A2(new_n10134_), .ZN(new_n10135_));
  NOR2_X1    g09836(.A1(new_n10135_), .A2(new_n10123_), .ZN(new_n10136_));
  AOI21_X1   g09837(.A1(new_n10130_), .A2(new_n10123_), .B(new_n10136_), .ZN(new_n10137_));
  INV_X1     g09838(.I(new_n10137_), .ZN(new_n10138_));
  AOI21_X1   g09839(.A1(new_n609_), .A2(new_n8676_), .B(new_n9864_), .ZN(new_n10139_));
  INV_X1     g09840(.I(new_n10139_), .ZN(new_n10140_));
  AOI21_X1   g09841(.A1(new_n229_), .A2(new_n9784_), .B(new_n9782_), .ZN(new_n10141_));
  INV_X1     g09842(.I(new_n10141_), .ZN(new_n10142_));
  AOI21_X1   g09843(.A1(new_n2690_), .A2(new_n5600_), .B(new_n9787_), .ZN(new_n10143_));
  XOR2_X1    g09844(.A1(new_n10143_), .A2(new_n10142_), .Z(new_n10144_));
  NOR2_X1    g09845(.A1(new_n10144_), .A2(new_n10140_), .ZN(new_n10145_));
  INV_X1     g09846(.I(new_n10143_), .ZN(new_n10146_));
  NOR2_X1    g09847(.A1(new_n10146_), .A2(new_n10142_), .ZN(new_n10147_));
  NOR2_X1    g09848(.A1(new_n10143_), .A2(new_n10141_), .ZN(new_n10148_));
  NOR2_X1    g09849(.A1(new_n10147_), .A2(new_n10148_), .ZN(new_n10149_));
  NOR2_X1    g09850(.A1(new_n10149_), .A2(new_n10139_), .ZN(new_n10150_));
  NOR2_X1    g09851(.A1(new_n10150_), .A2(new_n10145_), .ZN(new_n10151_));
  NOR2_X1    g09852(.A1(\a[14] ), .A2(\a[52] ), .ZN(new_n10152_));
  OAI21_X1   g09853(.A1(new_n3127_), .A2(new_n3967_), .B(new_n10152_), .ZN(new_n10153_));
  OAI21_X1   g09854(.A1(new_n3126_), .A2(new_n3966_), .B(new_n10153_), .ZN(new_n10154_));
  AOI21_X1   g09855(.A1(new_n1275_), .A2(new_n4368_), .B(new_n6280_), .ZN(new_n10155_));
  NOR2_X1    g09856(.A1(new_n10154_), .A2(new_n10155_), .ZN(new_n10156_));
  XOR2_X1    g09857(.A1(new_n10156_), .A2(new_n242_), .Z(new_n10157_));
  XOR2_X1    g09858(.A1(new_n10157_), .A2(\a[61] ), .Z(new_n10158_));
  NOR2_X1    g09859(.A1(new_n10158_), .A2(new_n10151_), .ZN(new_n10159_));
  INV_X1     g09860(.I(new_n10151_), .ZN(new_n10160_));
  INV_X1     g09861(.I(new_n10158_), .ZN(new_n10161_));
  NOR2_X1    g09862(.A1(new_n10161_), .A2(new_n10160_), .ZN(new_n10162_));
  OAI21_X1   g09863(.A1(new_n10162_), .A2(new_n10159_), .B(new_n10138_), .ZN(new_n10163_));
  XOR2_X1    g09864(.A1(new_n10158_), .A2(new_n10151_), .Z(new_n10164_));
  NAND2_X1   g09865(.A1(new_n10164_), .A2(new_n10137_), .ZN(new_n10165_));
  NAND2_X1   g09866(.A1(new_n10165_), .A2(new_n10163_), .ZN(new_n10166_));
  XOR2_X1    g09867(.A1(new_n10166_), .A2(new_n10122_), .Z(new_n10167_));
  INV_X1     g09868(.I(new_n10167_), .ZN(new_n10168_));
  OAI21_X1   g09869(.A1(new_n10115_), .A2(new_n10121_), .B(new_n10166_), .ZN(new_n10169_));
  NAND3_X1   g09870(.A1(new_n10165_), .A2(new_n10122_), .A3(new_n10163_), .ZN(new_n10170_));
  AOI21_X1   g09871(.A1(new_n10169_), .A2(new_n10170_), .B(new_n10105_), .ZN(new_n10171_));
  AOI21_X1   g09872(.A1(new_n10105_), .A2(new_n10168_), .B(new_n10171_), .ZN(new_n10172_));
  NOR2_X1    g09873(.A1(new_n9755_), .A2(new_n9762_), .ZN(new_n10173_));
  NOR2_X1    g09874(.A1(new_n10173_), .A2(new_n9761_), .ZN(new_n10174_));
  INV_X1     g09875(.I(new_n9502_), .ZN(new_n10175_));
  NOR2_X1    g09876(.A1(new_n7700_), .A2(new_n10175_), .ZN(new_n10176_));
  NOR4_X1    g09877(.A1(new_n675_), .A2(new_n1215_), .A3(new_n5511_), .A4(new_n7216_), .ZN(new_n10181_));
  INV_X1     g09878(.I(new_n10181_), .ZN(new_n10182_));
  NOR2_X1    g09879(.A1(new_n7000_), .A2(new_n2328_), .ZN(new_n10183_));
  NAND2_X1   g09880(.A1(new_n1276_), .A2(new_n5750_), .ZN(new_n10184_));
  AOI21_X1   g09881(.A1(new_n2328_), .A2(new_n7000_), .B(new_n10184_), .ZN(new_n10185_));
  NOR2_X1    g09882(.A1(new_n10185_), .A2(new_n10183_), .ZN(new_n10186_));
  INV_X1     g09883(.I(new_n10186_), .ZN(new_n10187_));
  NOR2_X1    g09884(.A1(new_n10187_), .A2(new_n10182_), .ZN(new_n10188_));
  NOR2_X1    g09885(.A1(new_n10186_), .A2(new_n10181_), .ZN(new_n10189_));
  NOR2_X1    g09886(.A1(new_n10188_), .A2(new_n10189_), .ZN(new_n10190_));
  NOR3_X1    g09887(.A1(new_n10190_), .A2(new_n9773_), .A3(new_n9776_), .ZN(new_n10191_));
  XOR2_X1    g09888(.A1(new_n10186_), .A2(new_n10182_), .Z(new_n10192_));
  NOR2_X1    g09889(.A1(new_n9778_), .A2(new_n10192_), .ZN(new_n10193_));
  NOR2_X1    g09890(.A1(new_n10191_), .A2(new_n10193_), .ZN(new_n10194_));
  INV_X1     g09891(.I(new_n9829_), .ZN(new_n10195_));
  AOI21_X1   g09892(.A1(new_n10195_), .A2(new_n9832_), .B(new_n9828_), .ZN(new_n10196_));
  XNOR2_X1   g09893(.A1(new_n10196_), .A2(new_n10194_), .ZN(new_n10197_));
  NOR2_X1    g09894(.A1(new_n10174_), .A2(new_n10197_), .ZN(new_n10198_));
  OR2_X2     g09895(.A1(new_n10196_), .A2(new_n10194_), .Z(new_n10199_));
  NAND2_X1   g09896(.A1(new_n10196_), .A2(new_n10194_), .ZN(new_n10200_));
  NAND2_X1   g09897(.A1(new_n10199_), .A2(new_n10200_), .ZN(new_n10201_));
  AOI21_X1   g09898(.A1(new_n10174_), .A2(new_n10201_), .B(new_n10198_), .ZN(new_n10202_));
  NAND2_X1   g09899(.A1(new_n9796_), .A2(new_n9839_), .ZN(new_n10203_));
  NAND2_X1   g09900(.A1(new_n10203_), .A2(new_n9838_), .ZN(new_n10204_));
  INV_X1     g09901(.I(new_n10204_), .ZN(new_n10205_));
  NAND2_X1   g09902(.A1(new_n9875_), .A2(new_n9860_), .ZN(new_n10206_));
  NAND2_X1   g09903(.A1(new_n10206_), .A2(new_n9874_), .ZN(new_n10207_));
  INV_X1     g09904(.I(new_n10207_), .ZN(new_n10208_));
  NOR2_X1    g09905(.A1(new_n10208_), .A2(new_n10205_), .ZN(new_n10209_));
  NOR2_X1    g09906(.A1(new_n10207_), .A2(new_n10204_), .ZN(new_n10210_));
  NOR2_X1    g09907(.A1(new_n10209_), .A2(new_n10210_), .ZN(new_n10211_));
  NOR2_X1    g09908(.A1(new_n10211_), .A2(new_n10202_), .ZN(new_n10212_));
  XOR2_X1    g09909(.A1(new_n10207_), .A2(new_n10205_), .Z(new_n10213_));
  INV_X1     g09910(.I(new_n10213_), .ZN(new_n10214_));
  AOI21_X1   g09911(.A1(new_n10202_), .A2(new_n10214_), .B(new_n10212_), .ZN(new_n10215_));
  XNOR2_X1   g09912(.A1(new_n10215_), .A2(new_n10172_), .ZN(new_n10216_));
  NOR2_X1    g09913(.A1(new_n10216_), .A2(new_n10104_), .ZN(new_n10217_));
  NOR2_X1    g09914(.A1(new_n10215_), .A2(new_n10172_), .ZN(new_n10218_));
  INV_X1     g09915(.I(new_n10218_), .ZN(new_n10219_));
  NAND2_X1   g09916(.A1(new_n10215_), .A2(new_n10172_), .ZN(new_n10220_));
  NAND2_X1   g09917(.A1(new_n10219_), .A2(new_n10220_), .ZN(new_n10221_));
  AOI21_X1   g09918(.A1(new_n10104_), .A2(new_n10221_), .B(new_n10217_), .ZN(new_n10222_));
  XNOR2_X1   g09919(.A1(new_n10102_), .A2(new_n10222_), .ZN(new_n10223_));
  XOR2_X1    g09920(.A1(new_n10223_), .A2(new_n10101_), .Z(new_n10224_));
  XOR2_X1    g09921(.A1(new_n10224_), .A2(new_n10096_), .Z(new_n10225_));
  NOR2_X1    g09922(.A1(new_n10225_), .A2(new_n9978_), .ZN(new_n10226_));
  INV_X1     g09923(.I(new_n10226_), .ZN(new_n10227_));
  NAND2_X1   g09924(.A1(new_n10225_), .A2(new_n9978_), .ZN(new_n10228_));
  NAND2_X1   g09925(.A1(new_n10227_), .A2(new_n10228_), .ZN(new_n10229_));
  XOR2_X1    g09926(.A1(new_n9976_), .A2(new_n10229_), .Z(\asquared[68] ));
  OAI21_X1   g09927(.A1(new_n10228_), .A2(new_n9970_), .B(new_n9741_), .ZN(new_n10231_));
  INV_X1     g09928(.I(new_n10231_), .ZN(new_n10232_));
  AOI21_X1   g09929(.A1(new_n9970_), .A2(new_n10228_), .B(new_n10232_), .ZN(new_n10233_));
  INV_X1     g09930(.I(new_n10233_), .ZN(new_n10234_));
  NOR2_X1    g09931(.A1(new_n9739_), .A2(new_n10234_), .ZN(new_n10235_));
  NOR3_X1    g09932(.A1(new_n10090_), .A2(new_n10095_), .A3(new_n10100_), .ZN(new_n10236_));
  NOR2_X1    g09933(.A1(new_n10096_), .A2(new_n10099_), .ZN(new_n10237_));
  INV_X1     g09934(.I(new_n10237_), .ZN(new_n10238_));
  AOI21_X1   g09935(.A1(new_n10238_), .A2(new_n10098_), .B(new_n10236_), .ZN(new_n10239_));
  OAI21_X1   g09936(.A1(new_n10104_), .A2(new_n10218_), .B(new_n10220_), .ZN(new_n10240_));
  INV_X1     g09937(.I(new_n10240_), .ZN(new_n10241_));
  OAI21_X1   g09938(.A1(new_n9979_), .A2(new_n10092_), .B(new_n10094_), .ZN(new_n10242_));
  INV_X1     g09939(.I(new_n10210_), .ZN(new_n10243_));
  AOI21_X1   g09940(.A1(new_n10202_), .A2(new_n10243_), .B(new_n10209_), .ZN(new_n10244_));
  AOI21_X1   g09941(.A1(new_n10116_), .A2(new_n10120_), .B(new_n10118_), .ZN(new_n10245_));
  OAI21_X1   g09942(.A1(new_n10173_), .A2(new_n9761_), .B(new_n10200_), .ZN(new_n10246_));
  NAND2_X1   g09943(.A1(new_n10246_), .A2(new_n10199_), .ZN(new_n10247_));
  INV_X1     g09944(.I(new_n10162_), .ZN(new_n10248_));
  OAI21_X1   g09945(.A1(new_n10138_), .A2(new_n10159_), .B(new_n10248_), .ZN(new_n10249_));
  XNOR2_X1   g09946(.A1(new_n10249_), .A2(new_n10247_), .ZN(new_n10250_));
  NAND2_X1   g09947(.A1(new_n10249_), .A2(new_n10247_), .ZN(new_n10251_));
  INV_X1     g09948(.I(new_n10251_), .ZN(new_n10252_));
  NOR2_X1    g09949(.A1(new_n10249_), .A2(new_n10247_), .ZN(new_n10253_));
  OAI21_X1   g09950(.A1(new_n10252_), .A2(new_n10253_), .B(new_n10245_), .ZN(new_n10254_));
  OAI21_X1   g09951(.A1(new_n10245_), .A2(new_n10250_), .B(new_n10254_), .ZN(new_n10255_));
  NOR2_X1    g09952(.A1(new_n8678_), .A2(new_n2393_), .ZN(new_n10256_));
  NOR4_X1    g09953(.A1(new_n8245_), .A2(new_n797_), .A3(new_n364_), .A4(new_n8085_), .ZN(new_n10257_));
  NAND2_X1   g09954(.A1(new_n10256_), .A2(new_n10257_), .ZN(new_n10258_));
  INV_X1     g09955(.I(new_n10258_), .ZN(new_n10259_));
  AOI22_X1   g09956(.A1(new_n2500_), .A2(new_n5592_), .B1(new_n4415_), .B2(new_n2797_), .ZN(new_n10260_));
  NOR4_X1    g09957(.A1(new_n2690_), .A2(new_n6024_), .A3(new_n2098_), .A4(new_n4414_), .ZN(new_n10261_));
  NAND2_X1   g09958(.A1(new_n10260_), .A2(new_n10261_), .ZN(new_n10262_));
  NAND2_X1   g09959(.A1(new_n9549_), .A2(new_n608_), .ZN(new_n10263_));
  NOR2_X1    g09960(.A1(new_n1313_), .A2(new_n5511_), .ZN(new_n10264_));
  XOR2_X1    g09961(.A1(new_n10263_), .A2(new_n10264_), .Z(new_n10265_));
  NOR2_X1    g09962(.A1(new_n10265_), .A2(new_n10262_), .ZN(new_n10266_));
  INV_X1     g09963(.I(new_n10266_), .ZN(new_n10267_));
  NAND2_X1   g09964(.A1(new_n10265_), .A2(new_n10262_), .ZN(new_n10268_));
  NAND2_X1   g09965(.A1(new_n10267_), .A2(new_n10268_), .ZN(new_n10269_));
  XNOR2_X1   g09966(.A1(new_n10265_), .A2(new_n10262_), .ZN(new_n10270_));
  NOR2_X1    g09967(.A1(new_n10270_), .A2(new_n10259_), .ZN(new_n10271_));
  AOI21_X1   g09968(.A1(new_n10259_), .A2(new_n10269_), .B(new_n10271_), .ZN(new_n10272_));
  AOI22_X1   g09969(.A1(new_n3126_), .A2(new_n3805_), .B1(new_n2766_), .B2(new_n5600_), .ZN(new_n10273_));
  NOR2_X1    g09970(.A1(new_n2461_), .A2(new_n3804_), .ZN(new_n10274_));
  NAND4_X1   g09971(.A1(new_n10273_), .A2(new_n3839_), .A3(new_n4184_), .A4(new_n10274_), .ZN(new_n10275_));
  NAND4_X1   g09972(.A1(\a[12] ), .A2(\a[13] ), .A3(\a[55] ), .A4(\a[56] ), .ZN(new_n10276_));
  NAND2_X1   g09973(.A1(\a[49] ), .A2(\a[50] ), .ZN(new_n10277_));
  NOR2_X1    g09974(.A1(new_n2331_), .A2(new_n10277_), .ZN(new_n10278_));
  NAND2_X1   g09975(.A1(new_n2331_), .A2(new_n10277_), .ZN(new_n10279_));
  INV_X1     g09976(.I(new_n10279_), .ZN(new_n10280_));
  NOR2_X1    g09977(.A1(new_n10280_), .A2(new_n10278_), .ZN(new_n10281_));
  NOR2_X1    g09978(.A1(new_n10281_), .A2(new_n10276_), .ZN(new_n10282_));
  AND2_X2    g09979(.A1(new_n10281_), .A2(new_n10276_), .Z(new_n10283_));
  NOR2_X1    g09980(.A1(new_n10283_), .A2(new_n10282_), .ZN(new_n10284_));
  XOR2_X1    g09981(.A1(new_n10281_), .A2(new_n10276_), .Z(new_n10285_));
  NAND2_X1   g09982(.A1(new_n10285_), .A2(new_n10275_), .ZN(new_n10286_));
  OAI21_X1   g09983(.A1(new_n10275_), .A2(new_n10284_), .B(new_n10286_), .ZN(new_n10287_));
  INV_X1     g09984(.I(new_n7482_), .ZN(new_n10288_));
  NOR2_X1    g09985(.A1(new_n6692_), .A2(new_n6945_), .ZN(new_n10289_));
  INV_X1     g09986(.I(new_n10289_), .ZN(new_n10290_));
  NOR2_X1    g09987(.A1(new_n10288_), .A2(new_n10290_), .ZN(new_n10291_));
  NOR2_X1    g09988(.A1(new_n10291_), .A2(new_n1019_), .ZN(new_n10292_));
  NOR2_X1    g09989(.A1(new_n650_), .A2(new_n6945_), .ZN(new_n10293_));
  NAND4_X1   g09990(.A1(new_n10292_), .A2(new_n1021_), .A3(new_n8056_), .A4(new_n10293_), .ZN(new_n10294_));
  NAND2_X1   g09991(.A1(new_n5488_), .A2(new_n2286_), .ZN(new_n10295_));
  NOR2_X1    g09992(.A1(new_n1215_), .A2(new_n5750_), .ZN(new_n10296_));
  XOR2_X1    g09993(.A1(new_n10295_), .A2(new_n10296_), .Z(new_n10297_));
  NOR2_X1    g09994(.A1(new_n9357_), .A2(new_n2749_), .ZN(new_n10298_));
  NOR4_X1    g09995(.A1(new_n2752_), .A2(new_n5173_), .A3(new_n1691_), .A4(new_n4770_), .ZN(new_n10299_));
  NAND2_X1   g09996(.A1(new_n10298_), .A2(new_n10299_), .ZN(new_n10300_));
  NOR2_X1    g09997(.A1(new_n10300_), .A2(new_n10297_), .ZN(new_n10301_));
  INV_X1     g09998(.I(new_n10301_), .ZN(new_n10302_));
  NAND2_X1   g09999(.A1(new_n10300_), .A2(new_n10297_), .ZN(new_n10303_));
  AOI21_X1   g10000(.A1(new_n10302_), .A2(new_n10303_), .B(new_n10294_), .ZN(new_n10304_));
  INV_X1     g10001(.I(new_n10294_), .ZN(new_n10305_));
  XNOR2_X1   g10002(.A1(new_n10300_), .A2(new_n10297_), .ZN(new_n10306_));
  NOR2_X1    g10003(.A1(new_n10306_), .A2(new_n10305_), .ZN(new_n10307_));
  NOR2_X1    g10004(.A1(new_n10307_), .A2(new_n10304_), .ZN(new_n10308_));
  XOR2_X1    g10005(.A1(new_n10308_), .A2(new_n10287_), .Z(new_n10309_));
  INV_X1     g10006(.I(new_n10287_), .ZN(new_n10310_));
  NOR2_X1    g10007(.A1(new_n10308_), .A2(new_n10310_), .ZN(new_n10311_));
  NAND2_X1   g10008(.A1(new_n10308_), .A2(new_n10310_), .ZN(new_n10312_));
  INV_X1     g10009(.I(new_n10312_), .ZN(new_n10313_));
  OAI21_X1   g10010(.A1(new_n10313_), .A2(new_n10311_), .B(new_n10272_), .ZN(new_n10314_));
  OAI21_X1   g10011(.A1(new_n10272_), .A2(new_n10309_), .B(new_n10314_), .ZN(new_n10315_));
  XNOR2_X1   g10012(.A1(new_n10255_), .A2(new_n10315_), .ZN(new_n10316_));
  NOR2_X1    g10013(.A1(new_n10316_), .A2(new_n10244_), .ZN(new_n10317_));
  INV_X1     g10014(.I(new_n10244_), .ZN(new_n10318_));
  NAND2_X1   g10015(.A1(new_n10255_), .A2(new_n10315_), .ZN(new_n10319_));
  NOR2_X1    g10016(.A1(new_n10255_), .A2(new_n10315_), .ZN(new_n10320_));
  INV_X1     g10017(.I(new_n10320_), .ZN(new_n10321_));
  AOI21_X1   g10018(.A1(new_n10321_), .A2(new_n10319_), .B(new_n10318_), .ZN(new_n10322_));
  NOR2_X1    g10019(.A1(new_n10317_), .A2(new_n10322_), .ZN(new_n10323_));
  XNOR2_X1   g10020(.A1(new_n10323_), .A2(new_n10242_), .ZN(new_n10324_));
  NOR2_X1    g10021(.A1(new_n10323_), .A2(new_n10242_), .ZN(new_n10325_));
  NAND2_X1   g10022(.A1(new_n10323_), .A2(new_n10242_), .ZN(new_n10326_));
  INV_X1     g10023(.I(new_n10326_), .ZN(new_n10327_));
  OAI21_X1   g10024(.A1(new_n10327_), .A2(new_n10325_), .B(new_n10241_), .ZN(new_n10328_));
  OAI21_X1   g10025(.A1(new_n10241_), .A2(new_n10324_), .B(new_n10328_), .ZN(new_n10329_));
  NAND2_X1   g10026(.A1(new_n10005_), .A2(new_n9983_), .ZN(new_n10330_));
  NAND2_X1   g10027(.A1(new_n10330_), .A2(new_n10004_), .ZN(new_n10331_));
  INV_X1     g10028(.I(new_n10331_), .ZN(new_n10332_));
  OAI21_X1   g10029(.A1(new_n9985_), .A2(new_n9994_), .B(new_n9993_), .ZN(new_n10333_));
  INV_X1     g10030(.I(new_n10333_), .ZN(new_n10334_));
  AOI21_X1   g10031(.A1(new_n797_), .A2(new_n8242_), .B(new_n10176_), .ZN(new_n10335_));
  INV_X1     g10032(.I(new_n10335_), .ZN(new_n10336_));
  AOI21_X1   g10033(.A1(new_n454_), .A2(new_n8676_), .B(new_n10043_), .ZN(new_n10337_));
  AOI21_X1   g10034(.A1(new_n2543_), .A2(new_n5321_), .B(new_n10049_), .ZN(new_n10338_));
  XNOR2_X1   g10035(.A1(new_n10338_), .A2(new_n10337_), .ZN(new_n10339_));
  AND2_X2    g10036(.A1(new_n10338_), .A2(new_n10337_), .Z(new_n10340_));
  NOR2_X1    g10037(.A1(new_n10338_), .A2(new_n10337_), .ZN(new_n10341_));
  OAI21_X1   g10038(.A1(new_n10340_), .A2(new_n10341_), .B(new_n10336_), .ZN(new_n10342_));
  OAI21_X1   g10039(.A1(new_n10336_), .A2(new_n10339_), .B(new_n10342_), .ZN(new_n10343_));
  AOI21_X1   g10040(.A1(new_n10037_), .A2(new_n10038_), .B(new_n10036_), .ZN(new_n10344_));
  INV_X1     g10041(.I(new_n10344_), .ZN(new_n10345_));
  NAND2_X1   g10042(.A1(new_n2797_), .A2(new_n6024_), .ZN(new_n10346_));
  NOR2_X1    g10043(.A1(new_n2797_), .A2(new_n6024_), .ZN(new_n10347_));
  NOR2_X1    g10044(.A1(\a[4] ), .A2(\a[63] ), .ZN(new_n10348_));
  AOI21_X1   g10045(.A1(new_n10346_), .A2(new_n10348_), .B(new_n10347_), .ZN(new_n10349_));
  INV_X1     g10046(.I(new_n10349_), .ZN(new_n10350_));
  NOR2_X1    g10047(.A1(new_n10060_), .A2(new_n9523_), .ZN(new_n10351_));
  XOR2_X1    g10048(.A1(new_n10351_), .A2(new_n10350_), .Z(new_n10352_));
  NOR3_X1    g10049(.A1(new_n10350_), .A2(new_n10060_), .A3(new_n9523_), .ZN(new_n10353_));
  NOR2_X1    g10050(.A1(new_n10351_), .A2(new_n10349_), .ZN(new_n10354_));
  OAI21_X1   g10051(.A1(new_n10354_), .A2(new_n10353_), .B(new_n10345_), .ZN(new_n10355_));
  OAI21_X1   g10052(.A1(new_n10352_), .A2(new_n10345_), .B(new_n10355_), .ZN(new_n10356_));
  XNOR2_X1   g10053(.A1(new_n10343_), .A2(new_n10356_), .ZN(new_n10357_));
  NOR2_X1    g10054(.A1(new_n10334_), .A2(new_n10357_), .ZN(new_n10358_));
  NAND2_X1   g10055(.A1(new_n10343_), .A2(new_n10356_), .ZN(new_n10359_));
  NOR2_X1    g10056(.A1(new_n10343_), .A2(new_n10356_), .ZN(new_n10360_));
  INV_X1     g10057(.I(new_n10360_), .ZN(new_n10361_));
  AOI21_X1   g10058(.A1(new_n10361_), .A2(new_n10359_), .B(new_n10333_), .ZN(new_n10362_));
  NOR2_X1    g10059(.A1(new_n10358_), .A2(new_n10362_), .ZN(new_n10363_));
  NOR3_X1    g10060(.A1(new_n7174_), .A2(new_n650_), .A3(new_n6694_), .ZN(new_n10364_));
  NAND2_X1   g10061(.A1(new_n10017_), .A2(new_n10018_), .ZN(new_n10365_));
  AND2_X2    g10062(.A1(new_n10016_), .A2(new_n10365_), .Z(new_n10366_));
  NAND2_X1   g10063(.A1(new_n7483_), .A2(new_n1220_), .ZN(new_n10367_));
  NOR2_X1    g10064(.A1(new_n7483_), .A2(new_n1220_), .ZN(new_n10368_));
  NOR2_X1    g10065(.A1(\a[29] ), .A2(\a[38] ), .ZN(new_n10369_));
  AOI21_X1   g10066(.A1(new_n10367_), .A2(new_n10369_), .B(new_n10368_), .ZN(new_n10370_));
  INV_X1     g10067(.I(new_n10370_), .ZN(new_n10371_));
  XOR2_X1    g10068(.A1(new_n10366_), .A2(new_n10371_), .Z(new_n10372_));
  NOR2_X1    g10069(.A1(new_n10372_), .A2(new_n10364_), .ZN(new_n10373_));
  INV_X1     g10070(.I(new_n10364_), .ZN(new_n10374_));
  INV_X1     g10071(.I(new_n10366_), .ZN(new_n10375_));
  NOR2_X1    g10072(.A1(new_n10375_), .A2(new_n10371_), .ZN(new_n10376_));
  NOR2_X1    g10073(.A1(new_n10366_), .A2(new_n10370_), .ZN(new_n10377_));
  NOR2_X1    g10074(.A1(new_n10376_), .A2(new_n10377_), .ZN(new_n10378_));
  NOR2_X1    g10075(.A1(new_n10378_), .A2(new_n10374_), .ZN(new_n10379_));
  NOR2_X1    g10076(.A1(new_n10379_), .A2(new_n10373_), .ZN(new_n10380_));
  OAI21_X1   g10077(.A1(new_n10024_), .A2(new_n10029_), .B(new_n10013_), .ZN(new_n10381_));
  OAI21_X1   g10078(.A1(new_n10025_), .A2(new_n10027_), .B(new_n10381_), .ZN(new_n10382_));
  INV_X1     g10079(.I(new_n10382_), .ZN(new_n10383_));
  NAND2_X1   g10080(.A1(new_n10077_), .A2(new_n10063_), .ZN(new_n10384_));
  NAND2_X1   g10081(.A1(new_n10384_), .A2(new_n10074_), .ZN(new_n10385_));
  INV_X1     g10082(.I(new_n10385_), .ZN(new_n10386_));
  NOR2_X1    g10083(.A1(new_n10386_), .A2(new_n10383_), .ZN(new_n10387_));
  NOR2_X1    g10084(.A1(new_n10385_), .A2(new_n10382_), .ZN(new_n10388_));
  NOR2_X1    g10085(.A1(new_n10387_), .A2(new_n10388_), .ZN(new_n10389_));
  NOR2_X1    g10086(.A1(new_n10389_), .A2(new_n10380_), .ZN(new_n10390_));
  XOR2_X1    g10087(.A1(new_n10385_), .A2(new_n10383_), .Z(new_n10391_));
  INV_X1     g10088(.I(new_n10391_), .ZN(new_n10392_));
  AOI21_X1   g10089(.A1(new_n10380_), .A2(new_n10392_), .B(new_n10390_), .ZN(new_n10393_));
  XNOR2_X1   g10090(.A1(new_n10393_), .A2(new_n10363_), .ZN(new_n10394_));
  NOR2_X1    g10091(.A1(new_n10332_), .A2(new_n10394_), .ZN(new_n10395_));
  NOR2_X1    g10092(.A1(new_n10393_), .A2(new_n10363_), .ZN(new_n10396_));
  INV_X1     g10093(.I(new_n10396_), .ZN(new_n10397_));
  NAND2_X1   g10094(.A1(new_n10393_), .A2(new_n10363_), .ZN(new_n10398_));
  AOI21_X1   g10095(.A1(new_n10397_), .A2(new_n10398_), .B(new_n10331_), .ZN(new_n10399_));
  NOR2_X1    g10096(.A1(new_n10395_), .A2(new_n10399_), .ZN(new_n10400_));
  NAND2_X1   g10097(.A1(new_n10169_), .A2(new_n10105_), .ZN(new_n10401_));
  NAND2_X1   g10098(.A1(new_n10401_), .A2(new_n10170_), .ZN(new_n10402_));
  AOI21_X1   g10099(.A1(new_n10033_), .A2(new_n10086_), .B(new_n10084_), .ZN(new_n10403_));
  INV_X1     g10100(.I(new_n10403_), .ZN(new_n10404_));
  INV_X1     g10101(.I(new_n10189_), .ZN(new_n10405_));
  AOI21_X1   g10102(.A1(new_n9778_), .A2(new_n10405_), .B(new_n10188_), .ZN(new_n10406_));
  INV_X1     g10103(.I(new_n10134_), .ZN(new_n10407_));
  AOI21_X1   g10104(.A1(new_n10123_), .A2(new_n10407_), .B(new_n10133_), .ZN(new_n10408_));
  NOR2_X1    g10105(.A1(new_n10053_), .A2(new_n10042_), .ZN(new_n10409_));
  NOR2_X1    g10106(.A1(new_n10409_), .A2(new_n10052_), .ZN(new_n10410_));
  XNOR2_X1   g10107(.A1(new_n10410_), .A2(new_n10408_), .ZN(new_n10411_));
  NOR2_X1    g10108(.A1(new_n10411_), .A2(new_n10406_), .ZN(new_n10412_));
  INV_X1     g10109(.I(new_n10406_), .ZN(new_n10413_));
  NOR2_X1    g10110(.A1(new_n10410_), .A2(new_n10408_), .ZN(new_n10414_));
  INV_X1     g10111(.I(new_n10414_), .ZN(new_n10415_));
  NAND2_X1   g10112(.A1(new_n10410_), .A2(new_n10408_), .ZN(new_n10416_));
  AOI21_X1   g10113(.A1(new_n10415_), .A2(new_n10416_), .B(new_n10413_), .ZN(new_n10417_));
  NOR2_X1    g10114(.A1(new_n10412_), .A2(new_n10417_), .ZN(new_n10418_));
  NOR2_X1    g10115(.A1(new_n359_), .A2(new_n8453_), .ZN(new_n10419_));
  XNOR2_X1   g10116(.A1(new_n10045_), .A2(new_n10419_), .ZN(new_n10420_));
  INV_X1     g10117(.I(new_n10420_), .ZN(new_n10421_));
  INV_X1     g10118(.I(new_n10148_), .ZN(new_n10422_));
  AOI21_X1   g10119(.A1(new_n10139_), .A2(new_n10422_), .B(new_n10147_), .ZN(new_n10423_));
  NAND2_X1   g10120(.A1(new_n10154_), .A2(new_n10155_), .ZN(new_n10424_));
  NOR2_X1    g10121(.A1(new_n242_), .A2(new_n8453_), .ZN(new_n10425_));
  AOI21_X1   g10122(.A1(new_n10424_), .A2(new_n10425_), .B(new_n10156_), .ZN(new_n10426_));
  NAND2_X1   g10123(.A1(new_n6733_), .A2(new_n3371_), .ZN(new_n10427_));
  NOR2_X1    g10124(.A1(new_n353_), .A2(new_n9029_), .ZN(new_n10428_));
  AOI21_X1   g10125(.A1(new_n10427_), .A2(new_n10428_), .B(new_n10067_), .ZN(new_n10429_));
  INV_X1     g10126(.I(new_n10429_), .ZN(new_n10430_));
  XOR2_X1    g10127(.A1(new_n10426_), .A2(new_n10430_), .Z(new_n10431_));
  XNOR2_X1   g10128(.A1(new_n10431_), .A2(new_n10423_), .ZN(new_n10432_));
  XOR2_X1    g10129(.A1(new_n10432_), .A2(new_n10421_), .Z(new_n10433_));
  XOR2_X1    g10130(.A1(new_n10433_), .A2(new_n10418_), .Z(new_n10434_));
  NAND2_X1   g10131(.A1(new_n10434_), .A2(new_n10404_), .ZN(new_n10435_));
  NOR2_X1    g10132(.A1(new_n10433_), .A2(new_n10418_), .ZN(new_n10436_));
  INV_X1     g10133(.I(new_n10436_), .ZN(new_n10437_));
  NAND2_X1   g10134(.A1(new_n10433_), .A2(new_n10418_), .ZN(new_n10438_));
  NAND2_X1   g10135(.A1(new_n10437_), .A2(new_n10438_), .ZN(new_n10439_));
  NAND2_X1   g10136(.A1(new_n10439_), .A2(new_n10403_), .ZN(new_n10440_));
  NAND2_X1   g10137(.A1(new_n10440_), .A2(new_n10435_), .ZN(new_n10441_));
  XOR2_X1    g10138(.A1(new_n10441_), .A2(new_n10402_), .Z(new_n10442_));
  NOR2_X1    g10139(.A1(new_n10442_), .A2(new_n10400_), .ZN(new_n10443_));
  INV_X1     g10140(.I(new_n10441_), .ZN(new_n10444_));
  NOR2_X1    g10141(.A1(new_n10444_), .A2(new_n10402_), .ZN(new_n10445_));
  INV_X1     g10142(.I(new_n10445_), .ZN(new_n10446_));
  NAND2_X1   g10143(.A1(new_n10444_), .A2(new_n10402_), .ZN(new_n10447_));
  NAND2_X1   g10144(.A1(new_n10446_), .A2(new_n10447_), .ZN(new_n10448_));
  AOI21_X1   g10145(.A1(new_n10400_), .A2(new_n10448_), .B(new_n10443_), .ZN(new_n10449_));
  OR2_X2     g10146(.A1(new_n10329_), .A2(new_n10449_), .Z(new_n10450_));
  NAND2_X1   g10147(.A1(new_n10329_), .A2(new_n10449_), .ZN(new_n10451_));
  AOI21_X1   g10148(.A1(new_n10450_), .A2(new_n10451_), .B(new_n10239_), .ZN(new_n10452_));
  XOR2_X1    g10149(.A1(new_n10329_), .A2(new_n10449_), .Z(new_n10453_));
  AOI21_X1   g10150(.A1(new_n10239_), .A2(new_n10453_), .B(new_n10452_), .ZN(new_n10454_));
  INV_X1     g10151(.I(new_n10222_), .ZN(new_n10455_));
  NAND2_X1   g10152(.A1(new_n10455_), .A2(new_n10102_), .ZN(new_n10456_));
  NOR2_X1    g10153(.A1(new_n10455_), .A2(new_n10102_), .ZN(new_n10457_));
  XNOR2_X1   g10154(.A1(new_n10101_), .A2(new_n10096_), .ZN(new_n10458_));
  OAI21_X1   g10155(.A1(new_n10458_), .A2(new_n10457_), .B(new_n10456_), .ZN(new_n10459_));
  INV_X1     g10156(.I(new_n10459_), .ZN(new_n10460_));
  NOR2_X1    g10157(.A1(new_n10454_), .A2(new_n10460_), .ZN(new_n10461_));
  XOR2_X1    g10158(.A1(new_n10235_), .A2(new_n10461_), .Z(new_n10462_));
  XOR2_X1    g10159(.A1(new_n10462_), .A2(new_n10226_), .Z(\asquared[69] ));
  NOR2_X1    g10160(.A1(new_n10227_), .A2(new_n10454_), .ZN(new_n10464_));
  AOI21_X1   g10161(.A1(new_n10227_), .A2(new_n10454_), .B(new_n10460_), .ZN(new_n10465_));
  INV_X1     g10162(.I(new_n10465_), .ZN(new_n10466_));
  NOR3_X1    g10163(.A1(new_n9739_), .A2(new_n10234_), .A3(new_n10466_), .ZN(new_n10467_));
  NOR2_X1    g10164(.A1(new_n10467_), .A2(new_n10464_), .ZN(new_n10468_));
  OAI21_X1   g10165(.A1(new_n10241_), .A2(new_n10325_), .B(new_n10326_), .ZN(new_n10469_));
  INV_X1     g10166(.I(new_n10469_), .ZN(new_n10470_));
  NAND2_X1   g10167(.A1(new_n10446_), .A2(new_n10400_), .ZN(new_n10471_));
  AND2_X2    g10168(.A1(new_n10471_), .A2(new_n10447_), .Z(new_n10472_));
  NAND2_X1   g10169(.A1(new_n10319_), .A2(new_n10318_), .ZN(new_n10473_));
  NAND2_X1   g10170(.A1(new_n10473_), .A2(new_n10321_), .ZN(new_n10474_));
  INV_X1     g10171(.I(new_n10388_), .ZN(new_n10475_));
  AOI21_X1   g10172(.A1(new_n10380_), .A2(new_n10475_), .B(new_n10387_), .ZN(new_n10476_));
  NOR2_X1    g10173(.A1(new_n10341_), .A2(new_n10336_), .ZN(new_n10477_));
  NOR2_X1    g10174(.A1(new_n10477_), .A2(new_n10340_), .ZN(new_n10478_));
  AOI22_X1   g10175(.A1(new_n2331_), .A2(new_n6776_), .B1(new_n6779_), .B2(new_n4345_), .ZN(new_n10479_));
  INV_X1     g10176(.I(new_n10479_), .ZN(new_n10480_));
  NAND4_X1   g10177(.A1(new_n10034_), .A2(\a[19] ), .A3(\a[50] ), .A4(new_n1268_), .ZN(new_n10481_));
  NOR2_X1    g10178(.A1(new_n10480_), .A2(new_n10481_), .ZN(new_n10482_));
  NOR2_X1    g10179(.A1(new_n6146_), .A2(new_n6579_), .ZN(new_n10483_));
  NOR2_X1    g10180(.A1(new_n3355_), .A2(new_n2689_), .ZN(new_n10484_));
  NOR2_X1    g10181(.A1(new_n10483_), .A2(new_n10484_), .ZN(new_n10485_));
  NOR4_X1    g10182(.A1(new_n2898_), .A2(new_n6024_), .A3(new_n2178_), .A4(new_n4414_), .ZN(new_n10486_));
  NAND2_X1   g10183(.A1(new_n10485_), .A2(new_n10486_), .ZN(new_n10487_));
  XOR2_X1    g10184(.A1(new_n10487_), .A2(new_n10482_), .Z(new_n10488_));
  NOR2_X1    g10185(.A1(new_n10478_), .A2(new_n10488_), .ZN(new_n10489_));
  INV_X1     g10186(.I(new_n10478_), .ZN(new_n10490_));
  INV_X1     g10187(.I(new_n10482_), .ZN(new_n10491_));
  NOR2_X1    g10188(.A1(new_n10491_), .A2(new_n10487_), .ZN(new_n10492_));
  INV_X1     g10189(.I(new_n10492_), .ZN(new_n10493_));
  NAND2_X1   g10190(.A1(new_n10491_), .A2(new_n10487_), .ZN(new_n10494_));
  AOI21_X1   g10191(.A1(new_n10493_), .A2(new_n10494_), .B(new_n10490_), .ZN(new_n10495_));
  NOR2_X1    g10192(.A1(new_n10495_), .A2(new_n10489_), .ZN(new_n10496_));
  INV_X1     g10193(.I(new_n10496_), .ZN(new_n10497_));
  NOR2_X1    g10194(.A1(new_n1215_), .A2(new_n6945_), .ZN(new_n10498_));
  NOR2_X1    g10195(.A1(new_n875_), .A2(new_n5745_), .ZN(new_n10499_));
  AOI22_X1   g10196(.A1(new_n10498_), .A2(new_n10499_), .B1(new_n7482_), .B2(new_n1719_), .ZN(new_n10500_));
  INV_X1     g10197(.I(new_n10500_), .ZN(new_n10501_));
  XNOR2_X1   g10198(.A1(new_n6735_), .A2(new_n8927_), .ZN(new_n10502_));
  OAI21_X1   g10199(.A1(new_n10502_), .A2(new_n6735_), .B(new_n10501_), .ZN(new_n10503_));
  OAI21_X1   g10200(.A1(new_n875_), .A2(new_n6945_), .B(new_n10502_), .ZN(new_n10504_));
  NAND2_X1   g10201(.A1(new_n10504_), .A2(new_n10503_), .ZN(new_n10505_));
  AOI22_X1   g10202(.A1(new_n3805_), .A2(new_n3981_), .B1(new_n2869_), .B2(new_n5600_), .ZN(new_n10506_));
  NOR4_X1    g10203(.A1(new_n3851_), .A2(new_n3838_), .A3(new_n2655_), .A4(new_n3804_), .ZN(new_n10507_));
  NAND2_X1   g10204(.A1(new_n10506_), .A2(new_n10507_), .ZN(new_n10508_));
  NAND2_X1   g10205(.A1(\a[34] ), .A2(\a[62] ), .ZN(new_n10509_));
  XOR2_X1    g10206(.A1(new_n4362_), .A2(new_n10509_), .Z(new_n10510_));
  NOR2_X1    g10207(.A1(new_n10508_), .A2(new_n10510_), .ZN(new_n10511_));
  AND2_X2    g10208(.A1(new_n10508_), .A2(new_n10510_), .Z(new_n10512_));
  NOR2_X1    g10209(.A1(new_n10512_), .A2(new_n10511_), .ZN(new_n10513_));
  NOR2_X1    g10210(.A1(new_n10513_), .A2(new_n10505_), .ZN(new_n10514_));
  INV_X1     g10211(.I(new_n10505_), .ZN(new_n10515_));
  XNOR2_X1   g10212(.A1(new_n10508_), .A2(new_n10510_), .ZN(new_n10516_));
  NOR2_X1    g10213(.A1(new_n10515_), .A2(new_n10516_), .ZN(new_n10517_));
  NOR2_X1    g10214(.A1(new_n10517_), .A2(new_n10514_), .ZN(new_n10518_));
  NOR2_X1    g10215(.A1(new_n10497_), .A2(new_n10518_), .ZN(new_n10519_));
  NOR3_X1    g10216(.A1(new_n10496_), .A2(new_n10514_), .A3(new_n10517_), .ZN(new_n10520_));
  NOR2_X1    g10217(.A1(new_n10519_), .A2(new_n10520_), .ZN(new_n10521_));
  NOR2_X1    g10218(.A1(new_n10521_), .A2(new_n10476_), .ZN(new_n10522_));
  INV_X1     g10219(.I(new_n10476_), .ZN(new_n10523_));
  XOR2_X1    g10220(.A1(new_n10496_), .A2(new_n10518_), .Z(new_n10524_));
  NOR2_X1    g10221(.A1(new_n10523_), .A2(new_n10524_), .ZN(new_n10525_));
  NOR2_X1    g10222(.A1(new_n10525_), .A2(new_n10522_), .ZN(new_n10526_));
  OAI21_X1   g10223(.A1(new_n10403_), .A2(new_n10436_), .B(new_n10438_), .ZN(new_n10527_));
  NAND2_X1   g10224(.A1(new_n10416_), .A2(new_n10413_), .ZN(new_n10528_));
  NAND2_X1   g10225(.A1(new_n10528_), .A2(new_n10415_), .ZN(new_n10529_));
  INV_X1     g10226(.I(new_n391_), .ZN(new_n10530_));
  AOI22_X1   g10227(.A1(new_n10530_), .A2(new_n8991_), .B1(new_n8455_), .B2(new_n454_), .ZN(new_n10531_));
  NAND4_X1   g10228(.A1(new_n10531_), .A2(new_n525_), .A3(new_n9553_), .A4(new_n10419_), .ZN(new_n10532_));
  NOR2_X1    g10229(.A1(new_n8424_), .A2(new_n7453_), .ZN(new_n10533_));
  NOR2_X1    g10230(.A1(new_n10533_), .A2(new_n6700_), .ZN(new_n10534_));
  NOR4_X1    g10231(.A1(new_n5742_), .A2(new_n2277_), .A3(new_n2368_), .A4(new_n5175_), .ZN(new_n10535_));
  NAND2_X1   g10232(.A1(new_n10534_), .A2(new_n10535_), .ZN(new_n10536_));
  NAND2_X1   g10233(.A1(new_n2533_), .A2(new_n5173_), .ZN(new_n10537_));
  NOR2_X1    g10234(.A1(new_n242_), .A2(new_n9310_), .ZN(new_n10538_));
  XOR2_X1    g10235(.A1(new_n10537_), .A2(new_n10538_), .Z(new_n10539_));
  NOR2_X1    g10236(.A1(new_n10536_), .A2(new_n10539_), .ZN(new_n10540_));
  INV_X1     g10237(.I(new_n10540_), .ZN(new_n10541_));
  NAND2_X1   g10238(.A1(new_n10536_), .A2(new_n10539_), .ZN(new_n10542_));
  AOI21_X1   g10239(.A1(new_n10541_), .A2(new_n10542_), .B(new_n10532_), .ZN(new_n10543_));
  INV_X1     g10240(.I(new_n10532_), .ZN(new_n10544_));
  XNOR2_X1   g10241(.A1(new_n10536_), .A2(new_n10539_), .ZN(new_n10545_));
  NOR2_X1    g10242(.A1(new_n10545_), .A2(new_n10544_), .ZN(new_n10546_));
  NOR2_X1    g10243(.A1(new_n10546_), .A2(new_n10543_), .ZN(new_n10547_));
  INV_X1     g10244(.I(new_n10547_), .ZN(new_n10548_));
  NOR2_X1    g10245(.A1(new_n8247_), .A2(new_n2668_), .ZN(new_n10549_));
  NOR2_X1    g10246(.A1(new_n675_), .A2(new_n7647_), .ZN(new_n10550_));
  NAND4_X1   g10247(.A1(new_n10549_), .A2(new_n1150_), .A3(new_n8243_), .A4(new_n10550_), .ZN(new_n10551_));
  AOI22_X1   g10248(.A1(new_n10430_), .A2(new_n609_), .B1(new_n8991_), .B2(new_n10421_), .ZN(new_n10552_));
  NAND2_X1   g10249(.A1(new_n6030_), .A2(new_n4538_), .ZN(new_n10553_));
  NAND2_X1   g10250(.A1(\a[14] ), .A2(\a[55] ), .ZN(new_n10554_));
  XNOR2_X1   g10251(.A1(new_n10553_), .A2(new_n10554_), .ZN(new_n10555_));
  XNOR2_X1   g10252(.A1(new_n10552_), .A2(new_n10555_), .ZN(new_n10556_));
  NOR2_X1    g10253(.A1(new_n10556_), .A2(new_n10551_), .ZN(new_n10557_));
  INV_X1     g10254(.I(new_n10551_), .ZN(new_n10558_));
  NOR2_X1    g10255(.A1(new_n10552_), .A2(new_n10555_), .ZN(new_n10559_));
  INV_X1     g10256(.I(new_n10559_), .ZN(new_n10560_));
  NAND2_X1   g10257(.A1(new_n10552_), .A2(new_n10555_), .ZN(new_n10561_));
  AOI21_X1   g10258(.A1(new_n10560_), .A2(new_n10561_), .B(new_n10558_), .ZN(new_n10562_));
  NOR2_X1    g10259(.A1(new_n10557_), .A2(new_n10562_), .ZN(new_n10563_));
  XOR2_X1    g10260(.A1(new_n10563_), .A2(new_n10548_), .Z(new_n10564_));
  NAND2_X1   g10261(.A1(new_n10564_), .A2(new_n10529_), .ZN(new_n10565_));
  INV_X1     g10262(.I(new_n10529_), .ZN(new_n10566_));
  NOR2_X1    g10263(.A1(new_n10563_), .A2(new_n10548_), .ZN(new_n10567_));
  NAND2_X1   g10264(.A1(new_n10563_), .A2(new_n10548_), .ZN(new_n10568_));
  INV_X1     g10265(.I(new_n10568_), .ZN(new_n10569_));
  OAI21_X1   g10266(.A1(new_n10569_), .A2(new_n10567_), .B(new_n10566_), .ZN(new_n10570_));
  NAND2_X1   g10267(.A1(new_n10565_), .A2(new_n10570_), .ZN(new_n10571_));
  INV_X1     g10268(.I(new_n10571_), .ZN(new_n10572_));
  NOR2_X1    g10269(.A1(new_n10527_), .A2(new_n10572_), .ZN(new_n10573_));
  INV_X1     g10270(.I(new_n10573_), .ZN(new_n10574_));
  NAND2_X1   g10271(.A1(new_n10527_), .A2(new_n10572_), .ZN(new_n10575_));
  AOI21_X1   g10272(.A1(new_n10574_), .A2(new_n10575_), .B(new_n10526_), .ZN(new_n10576_));
  XOR2_X1    g10273(.A1(new_n10527_), .A2(new_n10571_), .Z(new_n10577_));
  INV_X1     g10274(.I(new_n10577_), .ZN(new_n10578_));
  AOI21_X1   g10275(.A1(new_n10578_), .A2(new_n10526_), .B(new_n10576_), .ZN(new_n10579_));
  XOR2_X1    g10276(.A1(new_n10474_), .A2(new_n10579_), .Z(new_n10580_));
  NOR2_X1    g10277(.A1(new_n10472_), .A2(new_n10580_), .ZN(new_n10581_));
  INV_X1     g10278(.I(new_n10474_), .ZN(new_n10582_));
  NOR2_X1    g10279(.A1(new_n10582_), .A2(new_n10579_), .ZN(new_n10583_));
  INV_X1     g10280(.I(new_n10583_), .ZN(new_n10584_));
  NAND2_X1   g10281(.A1(new_n10582_), .A2(new_n10579_), .ZN(new_n10585_));
  NAND2_X1   g10282(.A1(new_n10584_), .A2(new_n10585_), .ZN(new_n10586_));
  AOI21_X1   g10283(.A1(new_n10472_), .A2(new_n10586_), .B(new_n10581_), .ZN(new_n10587_));
  OAI21_X1   g10284(.A1(new_n10332_), .A2(new_n10396_), .B(new_n10398_), .ZN(new_n10588_));
  INV_X1     g10285(.I(new_n10588_), .ZN(new_n10589_));
  OAI21_X1   g10286(.A1(new_n10245_), .A2(new_n10253_), .B(new_n10251_), .ZN(new_n10590_));
  NOR2_X1    g10287(.A1(new_n10423_), .A2(new_n10426_), .ZN(new_n10591_));
  XNOR2_X1   g10288(.A1(new_n10429_), .A2(new_n10420_), .ZN(new_n10592_));
  AOI21_X1   g10289(.A1(new_n10423_), .A2(new_n10426_), .B(new_n10592_), .ZN(new_n10593_));
  NOR2_X1    g10290(.A1(new_n10593_), .A2(new_n10591_), .ZN(new_n10594_));
  NOR2_X1    g10291(.A1(new_n10283_), .A2(new_n10275_), .ZN(new_n10595_));
  NOR2_X1    g10292(.A1(new_n10595_), .A2(new_n10282_), .ZN(new_n10596_));
  NAND2_X1   g10293(.A1(new_n10305_), .A2(new_n10303_), .ZN(new_n10597_));
  NAND2_X1   g10294(.A1(new_n10597_), .A2(new_n10302_), .ZN(new_n10598_));
  XOR2_X1    g10295(.A1(new_n10598_), .A2(new_n10596_), .Z(new_n10599_));
  INV_X1     g10296(.I(new_n10598_), .ZN(new_n10600_));
  NOR2_X1    g10297(.A1(new_n10600_), .A2(new_n10596_), .ZN(new_n10601_));
  NAND2_X1   g10298(.A1(new_n10600_), .A2(new_n10596_), .ZN(new_n10602_));
  INV_X1     g10299(.I(new_n10602_), .ZN(new_n10603_));
  OAI21_X1   g10300(.A1(new_n10603_), .A2(new_n10601_), .B(new_n10594_), .ZN(new_n10604_));
  OAI21_X1   g10301(.A1(new_n10594_), .A2(new_n10599_), .B(new_n10604_), .ZN(new_n10605_));
  AOI21_X1   g10302(.A1(new_n797_), .A2(new_n8245_), .B(new_n10256_), .ZN(new_n10606_));
  NOR2_X1    g10303(.A1(new_n9549_), .A2(new_n608_), .ZN(new_n10607_));
  NAND2_X1   g10304(.A1(new_n1313_), .A2(new_n5511_), .ZN(new_n10608_));
  AOI21_X1   g10305(.A1(new_n608_), .A2(new_n9549_), .B(new_n10608_), .ZN(new_n10609_));
  NOR2_X1    g10306(.A1(new_n10609_), .A2(new_n10607_), .ZN(new_n10610_));
  NOR2_X1    g10307(.A1(new_n5488_), .A2(new_n2286_), .ZN(new_n10611_));
  NAND2_X1   g10308(.A1(new_n1215_), .A2(new_n5750_), .ZN(new_n10612_));
  AOI21_X1   g10309(.A1(new_n2286_), .A2(new_n5488_), .B(new_n10612_), .ZN(new_n10613_));
  NOR2_X1    g10310(.A1(new_n10613_), .A2(new_n10611_), .ZN(new_n10614_));
  XNOR2_X1   g10311(.A1(new_n10610_), .A2(new_n10614_), .ZN(new_n10615_));
  INV_X1     g10312(.I(new_n10615_), .ZN(new_n10616_));
  NOR4_X1    g10313(.A1(new_n10609_), .A2(new_n10613_), .A3(new_n10607_), .A4(new_n10611_), .ZN(new_n10617_));
  INV_X1     g10314(.I(new_n10617_), .ZN(new_n10618_));
  NOR2_X1    g10315(.A1(new_n10610_), .A2(new_n10614_), .ZN(new_n10619_));
  INV_X1     g10316(.I(new_n10619_), .ZN(new_n10620_));
  AOI21_X1   g10317(.A1(new_n10618_), .A2(new_n10620_), .B(new_n10606_), .ZN(new_n10621_));
  AOI21_X1   g10318(.A1(new_n10616_), .A2(new_n10606_), .B(new_n10621_), .ZN(new_n10622_));
  AOI21_X1   g10319(.A1(new_n3838_), .A2(new_n3981_), .B(new_n10273_), .ZN(new_n10623_));
  INV_X1     g10320(.I(new_n10623_), .ZN(new_n10624_));
  AOI21_X1   g10321(.A1(new_n1719_), .A2(new_n7204_), .B(new_n10292_), .ZN(new_n10625_));
  AOI21_X1   g10322(.A1(new_n2331_), .A2(new_n3424_), .B(new_n6280_), .ZN(new_n10626_));
  XOR2_X1    g10323(.A1(new_n10625_), .A2(new_n10626_), .Z(new_n10627_));
  INV_X1     g10324(.I(new_n10626_), .ZN(new_n10628_));
  AND2_X2    g10325(.A1(new_n10625_), .A2(new_n10628_), .Z(new_n10629_));
  NOR2_X1    g10326(.A1(new_n10625_), .A2(new_n10628_), .ZN(new_n10630_));
  OAI21_X1   g10327(.A1(new_n10629_), .A2(new_n10630_), .B(new_n10624_), .ZN(new_n10631_));
  OAI21_X1   g10328(.A1(new_n10624_), .A2(new_n10627_), .B(new_n10631_), .ZN(new_n10632_));
  NAND2_X1   g10329(.A1(new_n10259_), .A2(new_n10268_), .ZN(new_n10633_));
  NAND2_X1   g10330(.A1(new_n10633_), .A2(new_n10267_), .ZN(new_n10634_));
  INV_X1     g10331(.I(new_n10634_), .ZN(new_n10635_));
  NOR2_X1    g10332(.A1(new_n10632_), .A2(new_n10635_), .ZN(new_n10636_));
  INV_X1     g10333(.I(new_n10636_), .ZN(new_n10637_));
  NAND2_X1   g10334(.A1(new_n10632_), .A2(new_n10635_), .ZN(new_n10638_));
  NAND2_X1   g10335(.A1(new_n10637_), .A2(new_n10638_), .ZN(new_n10639_));
  XOR2_X1    g10336(.A1(new_n10632_), .A2(new_n10635_), .Z(new_n10640_));
  MUX2_X1    g10337(.I0(new_n10639_), .I1(new_n10640_), .S(new_n10622_), .Z(new_n10641_));
  XNOR2_X1   g10338(.A1(new_n10641_), .A2(new_n10605_), .ZN(new_n10642_));
  INV_X1     g10339(.I(new_n10642_), .ZN(new_n10643_));
  NAND2_X1   g10340(.A1(new_n10641_), .A2(new_n10605_), .ZN(new_n10644_));
  NOR2_X1    g10341(.A1(new_n10641_), .A2(new_n10605_), .ZN(new_n10645_));
  INV_X1     g10342(.I(new_n10645_), .ZN(new_n10646_));
  AOI21_X1   g10343(.A1(new_n10646_), .A2(new_n10644_), .B(new_n10590_), .ZN(new_n10647_));
  AOI21_X1   g10344(.A1(new_n10643_), .A2(new_n10590_), .B(new_n10647_), .ZN(new_n10648_));
  AOI21_X1   g10345(.A1(new_n10333_), .A2(new_n10359_), .B(new_n10360_), .ZN(new_n10649_));
  NOR2_X1    g10346(.A1(new_n10354_), .A2(new_n10345_), .ZN(new_n10650_));
  NOR2_X1    g10347(.A1(new_n10650_), .A2(new_n10353_), .ZN(new_n10651_));
  NOR2_X1    g10348(.A1(new_n10377_), .A2(new_n10364_), .ZN(new_n10652_));
  NOR2_X1    g10349(.A1(new_n10652_), .A2(new_n10376_), .ZN(new_n10653_));
  AOI21_X1   g10350(.A1(new_n2690_), .A2(new_n6024_), .B(new_n10260_), .ZN(new_n10654_));
  NOR4_X1    g10351(.A1(new_n566_), .A2(new_n599_), .A3(new_n6999_), .A4(new_n7216_), .ZN(new_n10655_));
  INV_X1     g10352(.I(new_n10655_), .ZN(new_n10656_));
  AOI21_X1   g10353(.A1(new_n2752_), .A2(new_n5173_), .B(new_n10298_), .ZN(new_n10657_));
  XOR2_X1    g10354(.A1(new_n10657_), .A2(new_n10656_), .Z(new_n10658_));
  INV_X1     g10355(.I(new_n10657_), .ZN(new_n10659_));
  NOR2_X1    g10356(.A1(new_n10659_), .A2(new_n10656_), .ZN(new_n10660_));
  NOR2_X1    g10357(.A1(new_n10657_), .A2(new_n10655_), .ZN(new_n10661_));
  NOR2_X1    g10358(.A1(new_n10660_), .A2(new_n10661_), .ZN(new_n10662_));
  MUX2_X1    g10359(.I0(new_n10662_), .I1(new_n10658_), .S(new_n10654_), .Z(new_n10663_));
  XOR2_X1    g10360(.A1(new_n10663_), .A2(new_n10653_), .Z(new_n10664_));
  INV_X1     g10361(.I(new_n10653_), .ZN(new_n10665_));
  NOR2_X1    g10362(.A1(new_n10663_), .A2(new_n10665_), .ZN(new_n10666_));
  NAND2_X1   g10363(.A1(new_n10663_), .A2(new_n10665_), .ZN(new_n10667_));
  INV_X1     g10364(.I(new_n10667_), .ZN(new_n10668_));
  OAI21_X1   g10365(.A1(new_n10668_), .A2(new_n10666_), .B(new_n10651_), .ZN(new_n10669_));
  OAI21_X1   g10366(.A1(new_n10651_), .A2(new_n10664_), .B(new_n10669_), .ZN(new_n10670_));
  NOR2_X1    g10367(.A1(new_n10313_), .A2(new_n10272_), .ZN(new_n10671_));
  NOR2_X1    g10368(.A1(new_n10671_), .A2(new_n10311_), .ZN(new_n10672_));
  XNOR2_X1   g10369(.A1(new_n10670_), .A2(new_n10672_), .ZN(new_n10673_));
  NOR2_X1    g10370(.A1(new_n10673_), .A2(new_n10649_), .ZN(new_n10674_));
  INV_X1     g10371(.I(new_n10649_), .ZN(new_n10675_));
  NOR2_X1    g10372(.A1(new_n10670_), .A2(new_n10672_), .ZN(new_n10676_));
  INV_X1     g10373(.I(new_n10676_), .ZN(new_n10677_));
  NAND2_X1   g10374(.A1(new_n10670_), .A2(new_n10672_), .ZN(new_n10678_));
  AOI21_X1   g10375(.A1(new_n10677_), .A2(new_n10678_), .B(new_n10675_), .ZN(new_n10679_));
  NOR2_X1    g10376(.A1(new_n10674_), .A2(new_n10679_), .ZN(new_n10680_));
  XNOR2_X1   g10377(.A1(new_n10648_), .A2(new_n10680_), .ZN(new_n10681_));
  NOR2_X1    g10378(.A1(new_n10681_), .A2(new_n10589_), .ZN(new_n10682_));
  NOR2_X1    g10379(.A1(new_n10648_), .A2(new_n10680_), .ZN(new_n10683_));
  INV_X1     g10380(.I(new_n10683_), .ZN(new_n10684_));
  NAND2_X1   g10381(.A1(new_n10648_), .A2(new_n10680_), .ZN(new_n10685_));
  AOI21_X1   g10382(.A1(new_n10684_), .A2(new_n10685_), .B(new_n10588_), .ZN(new_n10686_));
  NOR2_X1    g10383(.A1(new_n10682_), .A2(new_n10686_), .ZN(new_n10687_));
  NOR2_X1    g10384(.A1(new_n10587_), .A2(new_n10687_), .ZN(new_n10688_));
  INV_X1     g10385(.I(new_n10688_), .ZN(new_n10689_));
  NAND2_X1   g10386(.A1(new_n10587_), .A2(new_n10687_), .ZN(new_n10690_));
  AOI21_X1   g10387(.A1(new_n10689_), .A2(new_n10690_), .B(new_n10470_), .ZN(new_n10691_));
  XOR2_X1    g10388(.A1(new_n10587_), .A2(new_n10687_), .Z(new_n10692_));
  AOI21_X1   g10389(.A1(new_n10470_), .A2(new_n10692_), .B(new_n10691_), .ZN(new_n10693_));
  INV_X1     g10390(.I(new_n10239_), .ZN(new_n10694_));
  NAND2_X1   g10391(.A1(new_n10451_), .A2(new_n10694_), .ZN(new_n10695_));
  NAND2_X1   g10392(.A1(new_n10695_), .A2(new_n10450_), .ZN(new_n10696_));
  XOR2_X1    g10393(.A1(new_n10693_), .A2(new_n10696_), .Z(new_n10697_));
  INV_X1     g10394(.I(new_n10696_), .ZN(new_n10698_));
  OR2_X2     g10395(.A1(new_n10698_), .A2(new_n10693_), .Z(new_n10699_));
  NAND2_X1   g10396(.A1(new_n10698_), .A2(new_n10693_), .ZN(new_n10700_));
  NAND2_X1   g10397(.A1(new_n10699_), .A2(new_n10700_), .ZN(new_n10701_));
  NAND2_X1   g10398(.A1(new_n10468_), .A2(new_n10701_), .ZN(new_n10702_));
  OAI21_X1   g10399(.A1(new_n10468_), .A2(new_n10697_), .B(new_n10702_), .ZN(\asquared[70] ));
  OAI21_X1   g10400(.A1(new_n10467_), .A2(new_n10464_), .B(new_n10700_), .ZN(new_n10704_));
  NAND2_X1   g10401(.A1(new_n10704_), .A2(new_n10699_), .ZN(new_n10705_));
  OAI21_X1   g10402(.A1(new_n10589_), .A2(new_n10683_), .B(new_n10685_), .ZN(new_n10706_));
  INV_X1     g10403(.I(new_n10706_), .ZN(new_n10707_));
  NAND2_X1   g10404(.A1(new_n10678_), .A2(new_n10675_), .ZN(new_n10708_));
  NOR2_X1    g10405(.A1(new_n8036_), .A2(new_n9799_), .ZN(new_n10709_));
  NOR4_X1    g10406(.A1(new_n566_), .A2(new_n1691_), .A3(new_n5175_), .A4(new_n7647_), .ZN(new_n10710_));
  NAND2_X1   g10407(.A1(new_n10709_), .A2(new_n10710_), .ZN(new_n10711_));
  AOI21_X1   g10408(.A1(new_n10711_), .A2(new_n8246_), .B(new_n1150_), .ZN(new_n10712_));
  NAND2_X1   g10409(.A1(\a[12] ), .A2(\a[58] ), .ZN(new_n10713_));
  NOR2_X1    g10410(.A1(new_n10712_), .A2(new_n10709_), .ZN(new_n10714_));
  INV_X1     g10411(.I(new_n10714_), .ZN(new_n10715_));
  OAI22_X1   g10412(.A1(new_n599_), .A2(new_n1691_), .B1(new_n5175_), .B2(new_n7727_), .ZN(new_n10716_));
  OAI22_X1   g10413(.A1(new_n10715_), .A2(new_n10716_), .B1(new_n10712_), .B2(new_n10713_), .ZN(new_n10717_));
  INV_X1     g10414(.I(new_n10717_), .ZN(new_n10718_));
  OAI21_X1   g10415(.A1(new_n8989_), .A2(new_n8992_), .B(new_n2394_), .ZN(new_n10719_));
  NAND4_X1   g10416(.A1(new_n9553_), .A2(\a[9] ), .A3(\a[61] ), .A4(new_n796_), .ZN(new_n10720_));
  NOR2_X1    g10417(.A1(new_n10719_), .A2(new_n10720_), .ZN(new_n10721_));
  NOR2_X1    g10418(.A1(new_n8056_), .A2(new_n10290_), .ZN(new_n10722_));
  NOR2_X1    g10419(.A1(new_n10722_), .A2(new_n1269_), .ZN(new_n10723_));
  INV_X1     g10420(.I(new_n10723_), .ZN(new_n10724_));
  NOR4_X1    g10421(.A1(new_n10724_), .A2(new_n1275_), .A3(new_n7482_), .A4(new_n8058_), .ZN(new_n10725_));
  AND2_X2    g10422(.A1(new_n10725_), .A2(new_n10721_), .Z(new_n10726_));
  NOR2_X1    g10423(.A1(new_n10725_), .A2(new_n10721_), .ZN(new_n10727_));
  OAI21_X1   g10424(.A1(new_n10726_), .A2(new_n10727_), .B(new_n10718_), .ZN(new_n10728_));
  XNOR2_X1   g10425(.A1(new_n10725_), .A2(new_n10721_), .ZN(new_n10729_));
  OAI21_X1   g10426(.A1(new_n10718_), .A2(new_n10729_), .B(new_n10728_), .ZN(new_n10730_));
  INV_X1     g10427(.I(new_n10730_), .ZN(new_n10731_));
  AOI22_X1   g10428(.A1(new_n3805_), .A2(new_n4368_), .B1(new_n3851_), .B2(new_n5600_), .ZN(new_n10732_));
  OAI21_X1   g10429(.A1(new_n3839_), .A2(new_n4644_), .B(new_n10732_), .ZN(new_n10733_));
  INV_X1     g10430(.I(new_n10733_), .ZN(new_n10734_));
  AOI21_X1   g10431(.A1(new_n10734_), .A2(new_n4727_), .B(\a[37] ), .ZN(new_n10735_));
  NOR2_X1    g10432(.A1(\a[32] ), .A2(\a[38] ), .ZN(new_n10736_));
  OAI21_X1   g10433(.A1(new_n10735_), .A2(new_n2868_), .B(new_n10736_), .ZN(new_n10737_));
  AOI21_X1   g10434(.A1(new_n3838_), .A2(new_n4372_), .B(new_n10732_), .ZN(new_n10738_));
  NAND2_X1   g10435(.A1(new_n10737_), .A2(new_n10738_), .ZN(new_n10739_));
  AOI21_X1   g10436(.A1(new_n6735_), .A2(new_n8927_), .B(new_n10501_), .ZN(new_n10740_));
  AOI21_X1   g10437(.A1(new_n1441_), .A2(new_n6777_), .B(new_n10479_), .ZN(new_n10741_));
  AND2_X2    g10438(.A1(new_n10740_), .A2(new_n10741_), .Z(new_n10742_));
  NOR2_X1    g10439(.A1(new_n10740_), .A2(new_n10741_), .ZN(new_n10743_));
  NOR2_X1    g10440(.A1(new_n10742_), .A2(new_n10743_), .ZN(new_n10744_));
  NOR2_X1    g10441(.A1(new_n10739_), .A2(new_n10744_), .ZN(new_n10745_));
  XNOR2_X1   g10442(.A1(new_n10740_), .A2(new_n10741_), .ZN(new_n10746_));
  INV_X1     g10443(.I(new_n10746_), .ZN(new_n10747_));
  AOI21_X1   g10444(.A1(new_n10739_), .A2(new_n10747_), .B(new_n10745_), .ZN(new_n10748_));
  OAI21_X1   g10445(.A1(new_n10651_), .A2(new_n10666_), .B(new_n10667_), .ZN(new_n10749_));
  XOR2_X1    g10446(.A1(new_n10749_), .A2(new_n10748_), .Z(new_n10750_));
  INV_X1     g10447(.I(new_n10749_), .ZN(new_n10751_));
  NOR2_X1    g10448(.A1(new_n10751_), .A2(new_n10748_), .ZN(new_n10752_));
  NAND2_X1   g10449(.A1(new_n10751_), .A2(new_n10748_), .ZN(new_n10753_));
  INV_X1     g10450(.I(new_n10753_), .ZN(new_n10754_));
  OAI21_X1   g10451(.A1(new_n10754_), .A2(new_n10752_), .B(new_n10731_), .ZN(new_n10755_));
  OAI21_X1   g10452(.A1(new_n10731_), .A2(new_n10750_), .B(new_n10755_), .ZN(new_n10756_));
  NAND2_X1   g10453(.A1(new_n10638_), .A2(new_n10622_), .ZN(new_n10757_));
  NAND2_X1   g10454(.A1(new_n10757_), .A2(new_n10637_), .ZN(new_n10758_));
  NOR2_X1    g10455(.A1(new_n10630_), .A2(new_n10624_), .ZN(new_n10759_));
  NOR2_X1    g10456(.A1(new_n10759_), .A2(new_n10629_), .ZN(new_n10760_));
  NOR2_X1    g10457(.A1(new_n3175_), .A2(new_n3734_), .ZN(new_n10761_));
  NOR2_X1    g10458(.A1(new_n10483_), .A2(new_n10761_), .ZN(new_n10762_));
  NOR2_X1    g10459(.A1(new_n2499_), .A2(new_n4414_), .ZN(new_n10763_));
  NAND4_X1   g10460(.A1(new_n10762_), .A2(new_n3127_), .A3(new_n4321_), .A4(new_n10763_), .ZN(new_n10764_));
  NOR2_X1    g10461(.A1(new_n2368_), .A2(new_n5511_), .ZN(new_n10765_));
  INV_X1     g10462(.I(new_n10765_), .ZN(new_n10766_));
  NOR2_X1    g10463(.A1(new_n2178_), .A2(new_n4769_), .ZN(new_n10767_));
  INV_X1     g10464(.I(new_n10767_), .ZN(new_n10768_));
  NOR2_X1    g10465(.A1(new_n10766_), .A2(new_n10768_), .ZN(new_n10769_));
  XOR2_X1    g10466(.A1(new_n10769_), .A2(new_n268_), .Z(new_n10770_));
  XOR2_X1    g10467(.A1(new_n10770_), .A2(\a[63] ), .Z(new_n10771_));
  XNOR2_X1   g10468(.A1(new_n10771_), .A2(new_n10764_), .ZN(new_n10772_));
  NOR2_X1    g10469(.A1(new_n10772_), .A2(new_n10760_), .ZN(new_n10773_));
  INV_X1     g10470(.I(new_n10760_), .ZN(new_n10774_));
  NOR2_X1    g10471(.A1(new_n10771_), .A2(new_n10764_), .ZN(new_n10775_));
  INV_X1     g10472(.I(new_n10775_), .ZN(new_n10776_));
  NAND2_X1   g10473(.A1(new_n10771_), .A2(new_n10764_), .ZN(new_n10777_));
  AOI21_X1   g10474(.A1(new_n10776_), .A2(new_n10777_), .B(new_n10774_), .ZN(new_n10778_));
  NAND2_X1   g10475(.A1(new_n8755_), .A2(new_n1447_), .ZN(new_n10779_));
  NOR2_X1    g10476(.A1(new_n1674_), .A2(new_n5750_), .ZN(new_n10780_));
  XOR2_X1    g10477(.A1(new_n10779_), .A2(new_n10780_), .Z(new_n10781_));
  AOI21_X1   g10478(.A1(new_n2752_), .A2(new_n2890_), .B(new_n7188_), .ZN(new_n10782_));
  NOR4_X1    g10479(.A1(new_n2533_), .A2(new_n5321_), .A3(new_n1999_), .A4(new_n5004_), .ZN(new_n10783_));
  NAND2_X1   g10480(.A1(new_n10782_), .A2(new_n10783_), .ZN(new_n10784_));
  INV_X1     g10481(.I(new_n9629_), .ZN(new_n10785_));
  NOR2_X1    g10482(.A1(new_n7512_), .A2(new_n10785_), .ZN(new_n10786_));
  NOR2_X1    g10483(.A1(new_n10786_), .A2(new_n1712_), .ZN(new_n10787_));
  NOR4_X1    g10484(.A1(new_n6779_), .A2(new_n1798_), .A3(new_n1313_), .A4(new_n5745_), .ZN(new_n10788_));
  NAND2_X1   g10485(.A1(new_n10787_), .A2(new_n10788_), .ZN(new_n10789_));
  NOR2_X1    g10486(.A1(new_n10784_), .A2(new_n10789_), .ZN(new_n10790_));
  INV_X1     g10487(.I(new_n10784_), .ZN(new_n10791_));
  INV_X1     g10488(.I(new_n10789_), .ZN(new_n10792_));
  NOR2_X1    g10489(.A1(new_n10791_), .A2(new_n10792_), .ZN(new_n10793_));
  NOR2_X1    g10490(.A1(new_n10793_), .A2(new_n10790_), .ZN(new_n10794_));
  NOR2_X1    g10491(.A1(new_n10794_), .A2(new_n10781_), .ZN(new_n10795_));
  XOR2_X1    g10492(.A1(new_n10784_), .A2(new_n10789_), .Z(new_n10796_));
  AOI21_X1   g10493(.A1(new_n10796_), .A2(new_n10781_), .B(new_n10795_), .ZN(new_n10797_));
  NOR3_X1    g10494(.A1(new_n10773_), .A2(new_n10778_), .A3(new_n10797_), .ZN(new_n10798_));
  NOR2_X1    g10495(.A1(new_n10773_), .A2(new_n10778_), .ZN(new_n10799_));
  INV_X1     g10496(.I(new_n10797_), .ZN(new_n10800_));
  NOR2_X1    g10497(.A1(new_n10799_), .A2(new_n10800_), .ZN(new_n10801_));
  OAI21_X1   g10498(.A1(new_n10801_), .A2(new_n10798_), .B(new_n10758_), .ZN(new_n10802_));
  INV_X1     g10499(.I(new_n10758_), .ZN(new_n10803_));
  XOR2_X1    g10500(.A1(new_n10799_), .A2(new_n10800_), .Z(new_n10804_));
  NAND2_X1   g10501(.A1(new_n10804_), .A2(new_n10803_), .ZN(new_n10805_));
  NAND2_X1   g10502(.A1(new_n10805_), .A2(new_n10802_), .ZN(new_n10806_));
  INV_X1     g10503(.I(new_n10806_), .ZN(new_n10807_));
  NOR2_X1    g10504(.A1(new_n10807_), .A2(new_n10756_), .ZN(new_n10808_));
  INV_X1     g10505(.I(new_n10808_), .ZN(new_n10809_));
  NAND2_X1   g10506(.A1(new_n10807_), .A2(new_n10756_), .ZN(new_n10810_));
  AOI22_X1   g10507(.A1(new_n10809_), .A2(new_n10810_), .B1(new_n10677_), .B2(new_n10708_), .ZN(new_n10811_));
  NAND2_X1   g10508(.A1(new_n10708_), .A2(new_n10677_), .ZN(new_n10812_));
  XOR2_X1    g10509(.A1(new_n10756_), .A2(new_n10806_), .Z(new_n10813_));
  NOR2_X1    g10510(.A1(new_n10813_), .A2(new_n10812_), .ZN(new_n10814_));
  INV_X1     g10511(.I(new_n10520_), .ZN(new_n10815_));
  AOI21_X1   g10512(.A1(new_n10523_), .A2(new_n10815_), .B(new_n10519_), .ZN(new_n10816_));
  AOI21_X1   g10513(.A1(new_n10490_), .A2(new_n10494_), .B(new_n10492_), .ZN(new_n10817_));
  AOI21_X1   g10514(.A1(new_n2898_), .A2(new_n6024_), .B(new_n10485_), .ZN(new_n10818_));
  INV_X1     g10515(.I(new_n10818_), .ZN(new_n10819_));
  AOI21_X1   g10516(.A1(new_n2277_), .A2(new_n5742_), .B(new_n10534_), .ZN(new_n10820_));
  NOR2_X1    g10517(.A1(new_n2533_), .A2(new_n5173_), .ZN(new_n10821_));
  NAND2_X1   g10518(.A1(new_n242_), .A2(new_n9310_), .ZN(new_n10822_));
  AOI21_X1   g10519(.A1(new_n2533_), .A2(new_n5173_), .B(new_n10822_), .ZN(new_n10823_));
  NOR2_X1    g10520(.A1(new_n10823_), .A2(new_n10821_), .ZN(new_n10824_));
  INV_X1     g10521(.I(new_n10824_), .ZN(new_n10825_));
  XOR2_X1    g10522(.A1(new_n10820_), .A2(new_n10825_), .Z(new_n10826_));
  NOR2_X1    g10523(.A1(new_n10826_), .A2(new_n10819_), .ZN(new_n10827_));
  INV_X1     g10524(.I(new_n10820_), .ZN(new_n10828_));
  NOR2_X1    g10525(.A1(new_n10828_), .A2(new_n10825_), .ZN(new_n10829_));
  NOR2_X1    g10526(.A1(new_n10820_), .A2(new_n10824_), .ZN(new_n10830_));
  NOR2_X1    g10527(.A1(new_n10829_), .A2(new_n10830_), .ZN(new_n10831_));
  NOR2_X1    g10528(.A1(new_n10831_), .A2(new_n10818_), .ZN(new_n10832_));
  NOR2_X1    g10529(.A1(new_n10832_), .A2(new_n10827_), .ZN(new_n10833_));
  AOI21_X1   g10530(.A1(new_n3851_), .A2(new_n3838_), .B(new_n10506_), .ZN(new_n10834_));
  INV_X1     g10531(.I(new_n10834_), .ZN(new_n10835_));
  AOI21_X1   g10532(.A1(\a[62] ), .A2(new_n4362_), .B(new_n3487_), .ZN(new_n10836_));
  INV_X1     g10533(.I(new_n10836_), .ZN(new_n10837_));
  NOR2_X1    g10534(.A1(new_n10835_), .A2(new_n10837_), .ZN(new_n10838_));
  XOR2_X1    g10535(.A1(new_n10838_), .A2(new_n359_), .Z(new_n10839_));
  XOR2_X1    g10536(.A1(new_n10839_), .A2(\a[62] ), .Z(new_n10840_));
  XOR2_X1    g10537(.A1(new_n10840_), .A2(new_n10833_), .Z(new_n10841_));
  NOR2_X1    g10538(.A1(new_n10841_), .A2(new_n10817_), .ZN(new_n10842_));
  INV_X1     g10539(.I(new_n10817_), .ZN(new_n10843_));
  INV_X1     g10540(.I(new_n10833_), .ZN(new_n10844_));
  NOR2_X1    g10541(.A1(new_n10840_), .A2(new_n10844_), .ZN(new_n10845_));
  INV_X1     g10542(.I(new_n10845_), .ZN(new_n10846_));
  NAND2_X1   g10543(.A1(new_n10840_), .A2(new_n10844_), .ZN(new_n10847_));
  AOI21_X1   g10544(.A1(new_n10846_), .A2(new_n10847_), .B(new_n10843_), .ZN(new_n10848_));
  NOR2_X1    g10545(.A1(new_n10842_), .A2(new_n10848_), .ZN(new_n10849_));
  INV_X1     g10546(.I(new_n10512_), .ZN(new_n10850_));
  AOI21_X1   g10547(.A1(new_n10515_), .A2(new_n10850_), .B(new_n10511_), .ZN(new_n10851_));
  NAND2_X1   g10548(.A1(new_n10542_), .A2(new_n10544_), .ZN(new_n10852_));
  NAND2_X1   g10549(.A1(new_n10852_), .A2(new_n10541_), .ZN(new_n10853_));
  INV_X1     g10550(.I(new_n10853_), .ZN(new_n10854_));
  NAND2_X1   g10551(.A1(new_n10561_), .A2(new_n10558_), .ZN(new_n10855_));
  NAND2_X1   g10552(.A1(new_n10855_), .A2(new_n10560_), .ZN(new_n10856_));
  XOR2_X1    g10553(.A1(new_n10856_), .A2(new_n10854_), .Z(new_n10857_));
  NOR2_X1    g10554(.A1(new_n10857_), .A2(new_n10851_), .ZN(new_n10858_));
  INV_X1     g10555(.I(new_n10851_), .ZN(new_n10859_));
  INV_X1     g10556(.I(new_n10856_), .ZN(new_n10860_));
  NOR2_X1    g10557(.A1(new_n10860_), .A2(new_n10854_), .ZN(new_n10861_));
  NOR2_X1    g10558(.A1(new_n10856_), .A2(new_n10853_), .ZN(new_n10862_));
  NOR2_X1    g10559(.A1(new_n10861_), .A2(new_n10862_), .ZN(new_n10863_));
  NOR2_X1    g10560(.A1(new_n10863_), .A2(new_n10859_), .ZN(new_n10864_));
  NOR2_X1    g10561(.A1(new_n10864_), .A2(new_n10858_), .ZN(new_n10865_));
  XNOR2_X1   g10562(.A1(new_n10849_), .A2(new_n10865_), .ZN(new_n10866_));
  NOR2_X1    g10563(.A1(new_n10866_), .A2(new_n10816_), .ZN(new_n10867_));
  INV_X1     g10564(.I(new_n10816_), .ZN(new_n10868_));
  NOR2_X1    g10565(.A1(new_n10849_), .A2(new_n10865_), .ZN(new_n10869_));
  INV_X1     g10566(.I(new_n10869_), .ZN(new_n10870_));
  NAND2_X1   g10567(.A1(new_n10849_), .A2(new_n10865_), .ZN(new_n10871_));
  AOI21_X1   g10568(.A1(new_n10870_), .A2(new_n10871_), .B(new_n10868_), .ZN(new_n10872_));
  NOR2_X1    g10569(.A1(new_n10867_), .A2(new_n10872_), .ZN(new_n10873_));
  NOR3_X1    g10570(.A1(new_n10814_), .A2(new_n10811_), .A3(new_n10873_), .ZN(new_n10874_));
  NOR2_X1    g10571(.A1(new_n10814_), .A2(new_n10811_), .ZN(new_n10875_));
  INV_X1     g10572(.I(new_n10873_), .ZN(new_n10876_));
  NOR2_X1    g10573(.A1(new_n10875_), .A2(new_n10876_), .ZN(new_n10877_));
  NOR2_X1    g10574(.A1(new_n10877_), .A2(new_n10874_), .ZN(new_n10878_));
  NOR2_X1    g10575(.A1(new_n10878_), .A2(new_n10707_), .ZN(new_n10879_));
  XOR2_X1    g10576(.A1(new_n10875_), .A2(new_n10873_), .Z(new_n10880_));
  NOR2_X1    g10577(.A1(new_n10880_), .A2(new_n10706_), .ZN(new_n10881_));
  NOR2_X1    g10578(.A1(new_n10881_), .A2(new_n10879_), .ZN(new_n10882_));
  INV_X1     g10579(.I(new_n10585_), .ZN(new_n10883_));
  OAI21_X1   g10580(.A1(new_n10472_), .A2(new_n10883_), .B(new_n10584_), .ZN(new_n10884_));
  AOI21_X1   g10581(.A1(new_n10590_), .A2(new_n10644_), .B(new_n10645_), .ZN(new_n10885_));
  OAI21_X1   g10582(.A1(new_n10566_), .A2(new_n10567_), .B(new_n10568_), .ZN(new_n10886_));
  NOR2_X1    g10583(.A1(new_n10594_), .A2(new_n10603_), .ZN(new_n10887_));
  NOR2_X1    g10584(.A1(new_n10887_), .A2(new_n10601_), .ZN(new_n10888_));
  AOI21_X1   g10585(.A1(new_n597_), .A2(new_n8996_), .B(new_n10531_), .ZN(new_n10889_));
  AOI21_X1   g10586(.A1(new_n1220_), .A2(new_n8242_), .B(new_n10549_), .ZN(new_n10890_));
  NOR2_X1    g10587(.A1(new_n6030_), .A2(new_n4538_), .ZN(new_n10891_));
  NAND2_X1   g10588(.A1(new_n650_), .A2(new_n6999_), .ZN(new_n10892_));
  AOI21_X1   g10589(.A1(new_n4538_), .A2(new_n6030_), .B(new_n10892_), .ZN(new_n10893_));
  NOR2_X1    g10590(.A1(new_n10893_), .A2(new_n10891_), .ZN(new_n10894_));
  XOR2_X1    g10591(.A1(new_n10890_), .A2(new_n10894_), .Z(new_n10895_));
  NAND2_X1   g10592(.A1(new_n10895_), .A2(new_n10889_), .ZN(new_n10896_));
  INV_X1     g10593(.I(new_n10889_), .ZN(new_n10897_));
  AND2_X2    g10594(.A1(new_n10890_), .A2(new_n10894_), .Z(new_n10898_));
  NOR2_X1    g10595(.A1(new_n10890_), .A2(new_n10894_), .ZN(new_n10899_));
  OAI21_X1   g10596(.A1(new_n10898_), .A2(new_n10899_), .B(new_n10897_), .ZN(new_n10900_));
  NAND2_X1   g10597(.A1(new_n10896_), .A2(new_n10900_), .ZN(new_n10901_));
  NAND2_X1   g10598(.A1(new_n10606_), .A2(new_n10620_), .ZN(new_n10902_));
  INV_X1     g10599(.I(new_n10661_), .ZN(new_n10903_));
  AOI21_X1   g10600(.A1(new_n10654_), .A2(new_n10903_), .B(new_n10660_), .ZN(new_n10904_));
  AOI21_X1   g10601(.A1(new_n10618_), .A2(new_n10902_), .B(new_n10904_), .ZN(new_n10905_));
  NAND2_X1   g10602(.A1(new_n10902_), .A2(new_n10618_), .ZN(new_n10906_));
  INV_X1     g10603(.I(new_n10904_), .ZN(new_n10907_));
  NOR2_X1    g10604(.A1(new_n10907_), .A2(new_n10906_), .ZN(new_n10908_));
  OAI21_X1   g10605(.A1(new_n10908_), .A2(new_n10905_), .B(new_n10901_), .ZN(new_n10909_));
  XNOR2_X1   g10606(.A1(new_n10904_), .A2(new_n10906_), .ZN(new_n10910_));
  NAND3_X1   g10607(.A1(new_n10910_), .A2(new_n10896_), .A3(new_n10900_), .ZN(new_n10911_));
  NAND2_X1   g10608(.A1(new_n10911_), .A2(new_n10909_), .ZN(new_n10912_));
  AND2_X2    g10609(.A1(new_n10912_), .A2(new_n10888_), .Z(new_n10913_));
  NOR2_X1    g10610(.A1(new_n10912_), .A2(new_n10888_), .ZN(new_n10914_));
  NOR2_X1    g10611(.A1(new_n10913_), .A2(new_n10914_), .ZN(new_n10915_));
  XNOR2_X1   g10612(.A1(new_n10912_), .A2(new_n10888_), .ZN(new_n10916_));
  MUX2_X1    g10613(.I0(new_n10916_), .I1(new_n10915_), .S(new_n10886_), .Z(new_n10917_));
  OAI21_X1   g10614(.A1(new_n10526_), .A2(new_n10573_), .B(new_n10575_), .ZN(new_n10918_));
  XOR2_X1    g10615(.A1(new_n10918_), .A2(new_n10917_), .Z(new_n10919_));
  NOR2_X1    g10616(.A1(new_n10919_), .A2(new_n10885_), .ZN(new_n10920_));
  INV_X1     g10617(.I(new_n10885_), .ZN(new_n10921_));
  INV_X1     g10618(.I(new_n10918_), .ZN(new_n10922_));
  NOR2_X1    g10619(.A1(new_n10922_), .A2(new_n10917_), .ZN(new_n10923_));
  INV_X1     g10620(.I(new_n10923_), .ZN(new_n10924_));
  NAND2_X1   g10621(.A1(new_n10922_), .A2(new_n10917_), .ZN(new_n10925_));
  AOI21_X1   g10622(.A1(new_n10924_), .A2(new_n10925_), .B(new_n10921_), .ZN(new_n10926_));
  NOR2_X1    g10623(.A1(new_n10926_), .A2(new_n10920_), .ZN(new_n10927_));
  XNOR2_X1   g10624(.A1(new_n10884_), .A2(new_n10927_), .ZN(new_n10928_));
  NOR2_X1    g10625(.A1(new_n10884_), .A2(new_n10927_), .ZN(new_n10929_));
  NAND2_X1   g10626(.A1(new_n10884_), .A2(new_n10927_), .ZN(new_n10930_));
  INV_X1     g10627(.I(new_n10930_), .ZN(new_n10931_));
  OAI21_X1   g10628(.A1(new_n10931_), .A2(new_n10929_), .B(new_n10882_), .ZN(new_n10932_));
  OAI21_X1   g10629(.A1(new_n10882_), .A2(new_n10928_), .B(new_n10932_), .ZN(new_n10933_));
  INV_X1     g10630(.I(new_n10933_), .ZN(new_n10934_));
  OAI21_X1   g10631(.A1(new_n10470_), .A2(new_n10688_), .B(new_n10690_), .ZN(new_n10935_));
  NAND2_X1   g10632(.A1(new_n10934_), .A2(new_n10935_), .ZN(new_n10936_));
  NOR2_X1    g10633(.A1(new_n10934_), .A2(new_n10935_), .ZN(new_n10937_));
  INV_X1     g10634(.I(new_n10937_), .ZN(new_n10938_));
  NAND2_X1   g10635(.A1(new_n10938_), .A2(new_n10936_), .ZN(new_n10939_));
  XOR2_X1    g10636(.A1(new_n10705_), .A2(new_n10939_), .Z(\asquared[71] ));
  NAND2_X1   g10637(.A1(new_n10936_), .A2(new_n10698_), .ZN(new_n10941_));
  OAI21_X1   g10638(.A1(new_n10936_), .A2(new_n10698_), .B(new_n10693_), .ZN(new_n10942_));
  AND2_X2    g10639(.A1(new_n10942_), .A2(new_n10941_), .Z(new_n10943_));
  OAI21_X1   g10640(.A1(new_n10467_), .A2(new_n10464_), .B(new_n10943_), .ZN(new_n10944_));
  OAI21_X1   g10641(.A1(new_n10882_), .A2(new_n10929_), .B(new_n10930_), .ZN(new_n10945_));
  INV_X1     g10642(.I(new_n10945_), .ZN(new_n10946_));
  INV_X1     g10643(.I(new_n10874_), .ZN(new_n10947_));
  AOI21_X1   g10644(.A1(new_n10947_), .A2(new_n10706_), .B(new_n10877_), .ZN(new_n10948_));
  AOI21_X1   g10645(.A1(new_n10921_), .A2(new_n10925_), .B(new_n10923_), .ZN(new_n10949_));
  INV_X1     g10646(.I(new_n10913_), .ZN(new_n10950_));
  AOI21_X1   g10647(.A1(new_n10950_), .A2(new_n10886_), .B(new_n10914_), .ZN(new_n10951_));
  INV_X1     g10648(.I(new_n10862_), .ZN(new_n10952_));
  AOI21_X1   g10649(.A1(new_n10859_), .A2(new_n10952_), .B(new_n10861_), .ZN(new_n10953_));
  AOI21_X1   g10650(.A1(new_n1798_), .A2(new_n6779_), .B(new_n10787_), .ZN(new_n10954_));
  NOR2_X1    g10651(.A1(new_n599_), .A2(new_n8085_), .ZN(new_n10955_));
  XNOR2_X1   g10652(.A1(new_n10955_), .A2(new_n10713_), .ZN(new_n10956_));
  XOR2_X1    g10653(.A1(new_n10954_), .A2(new_n10956_), .Z(new_n10957_));
  NOR2_X1    g10654(.A1(new_n6999_), .A2(new_n7727_), .ZN(new_n10958_));
  INV_X1     g10655(.I(new_n10958_), .ZN(new_n10959_));
  OAI21_X1   g10656(.A1(new_n8243_), .A2(new_n10959_), .B(new_n3383_), .ZN(new_n10960_));
  NAND4_X1   g10657(.A1(new_n8953_), .A2(\a[14] ), .A3(\a[57] ), .A4(new_n1021_), .ZN(new_n10961_));
  NOR2_X1    g10658(.A1(new_n10960_), .A2(new_n10961_), .ZN(new_n10962_));
  INV_X1     g10659(.I(new_n10962_), .ZN(new_n10963_));
  AOI21_X1   g10660(.A1(new_n5512_), .A2(new_n5980_), .B(new_n2749_), .ZN(new_n10964_));
  INV_X1     g10661(.I(new_n10964_), .ZN(new_n10965_));
  NAND4_X1   g10662(.A1(new_n2753_), .A2(new_n8424_), .A3(\a[24] ), .A4(\a[47] ), .ZN(new_n10966_));
  NOR2_X1    g10663(.A1(new_n10965_), .A2(new_n10966_), .ZN(new_n10967_));
  INV_X1     g10664(.I(new_n10967_), .ZN(new_n10968_));
  NOR2_X1    g10665(.A1(new_n10968_), .A2(new_n10963_), .ZN(new_n10969_));
  NOR2_X1    g10666(.A1(new_n10967_), .A2(new_n10962_), .ZN(new_n10970_));
  NOR2_X1    g10667(.A1(new_n10969_), .A2(new_n10970_), .ZN(new_n10971_));
  NOR2_X1    g10668(.A1(new_n10957_), .A2(new_n10971_), .ZN(new_n10972_));
  INV_X1     g10669(.I(new_n10957_), .ZN(new_n10973_));
  XNOR2_X1   g10670(.A1(new_n10967_), .A2(new_n10962_), .ZN(new_n10974_));
  NOR2_X1    g10671(.A1(new_n10973_), .A2(new_n10974_), .ZN(new_n10975_));
  NOR2_X1    g10672(.A1(new_n10975_), .A2(new_n10972_), .ZN(new_n10976_));
  AOI22_X1   g10673(.A1(new_n2500_), .A2(new_n5321_), .B1(new_n4771_), .B2(new_n2797_), .ZN(new_n10977_));
  NOR2_X1    g10674(.A1(new_n2098_), .A2(new_n4770_), .ZN(new_n10978_));
  NAND4_X1   g10675(.A1(new_n10977_), .A2(new_n2689_), .A3(new_n5174_), .A4(new_n10978_), .ZN(new_n10979_));
  AOI22_X1   g10676(.A1(new_n2766_), .A2(new_n5592_), .B1(new_n3126_), .B2(new_n4415_), .ZN(new_n10980_));
  NOR4_X1    g10677(.A1(new_n3981_), .A2(new_n6024_), .A3(new_n2461_), .A4(new_n4414_), .ZN(new_n10981_));
  NAND2_X1   g10678(.A1(new_n10980_), .A2(new_n10981_), .ZN(new_n10982_));
  NAND2_X1   g10679(.A1(new_n7482_), .A2(new_n1441_), .ZN(new_n10983_));
  NOR2_X1    g10680(.A1(new_n2368_), .A2(new_n5750_), .ZN(new_n10984_));
  XOR2_X1    g10681(.A1(new_n10983_), .A2(new_n10984_), .Z(new_n10985_));
  OR2_X2     g10682(.A1(new_n10985_), .A2(new_n10982_), .Z(new_n10986_));
  NAND2_X1   g10683(.A1(new_n10985_), .A2(new_n10982_), .ZN(new_n10987_));
  AOI21_X1   g10684(.A1(new_n10986_), .A2(new_n10987_), .B(new_n10979_), .ZN(new_n10988_));
  INV_X1     g10685(.I(new_n10979_), .ZN(new_n10989_));
  XNOR2_X1   g10686(.A1(new_n10985_), .A2(new_n10982_), .ZN(new_n10990_));
  NOR2_X1    g10687(.A1(new_n10990_), .A2(new_n10989_), .ZN(new_n10991_));
  NOR2_X1    g10688(.A1(new_n10991_), .A2(new_n10988_), .ZN(new_n10992_));
  XNOR2_X1   g10689(.A1(new_n10976_), .A2(new_n10992_), .ZN(new_n10993_));
  NOR2_X1    g10690(.A1(new_n10976_), .A2(new_n10992_), .ZN(new_n10994_));
  NAND2_X1   g10691(.A1(new_n10976_), .A2(new_n10992_), .ZN(new_n10995_));
  INV_X1     g10692(.I(new_n10995_), .ZN(new_n10996_));
  OAI21_X1   g10693(.A1(new_n10994_), .A2(new_n10996_), .B(new_n10953_), .ZN(new_n10997_));
  OAI21_X1   g10694(.A1(new_n10953_), .A2(new_n10993_), .B(new_n10997_), .ZN(new_n10998_));
  NOR2_X1    g10695(.A1(new_n10908_), .A2(new_n10901_), .ZN(new_n10999_));
  NOR2_X1    g10696(.A1(new_n10999_), .A2(new_n10905_), .ZN(new_n11000_));
  INV_X1     g10697(.I(new_n6776_), .ZN(new_n11001_));
  NOR2_X1    g10698(.A1(new_n8941_), .A2(new_n11001_), .ZN(new_n11002_));
  NOR2_X1    g10699(.A1(new_n11002_), .A2(new_n1712_), .ZN(new_n11003_));
  NOR2_X1    g10700(.A1(new_n1313_), .A2(new_n6055_), .ZN(new_n11004_));
  NAND4_X1   g10701(.A1(new_n11003_), .A2(new_n1715_), .A3(new_n10034_), .A4(new_n11004_), .ZN(new_n11005_));
  NAND4_X1   g10702(.A1(\a[33] ), .A2(\a[34] ), .A3(\a[37] ), .A4(\a[38] ), .ZN(new_n11006_));
  NAND2_X1   g10703(.A1(\a[22] ), .A2(\a[49] ), .ZN(new_n11007_));
  NOR2_X1    g10704(.A1(new_n11007_), .A2(new_n3393_), .ZN(new_n11008_));
  XOR2_X1    g10705(.A1(new_n11008_), .A2(new_n364_), .Z(new_n11009_));
  XOR2_X1    g10706(.A1(new_n11009_), .A2(\a[62] ), .Z(new_n11010_));
  OR2_X2     g10707(.A1(new_n11010_), .A2(new_n11006_), .Z(new_n11011_));
  NAND2_X1   g10708(.A1(new_n11010_), .A2(new_n11006_), .ZN(new_n11012_));
  AOI21_X1   g10709(.A1(new_n11011_), .A2(new_n11012_), .B(new_n11005_), .ZN(new_n11013_));
  XOR2_X1    g10710(.A1(new_n11010_), .A2(new_n11006_), .Z(new_n11014_));
  AOI21_X1   g10711(.A1(new_n11005_), .A2(new_n11014_), .B(new_n11013_), .ZN(new_n11015_));
  AOI21_X1   g10712(.A1(new_n1275_), .A2(new_n7482_), .B(new_n10723_), .ZN(new_n11016_));
  INV_X1     g10713(.I(new_n1101_), .ZN(new_n11017_));
  NOR2_X1    g10714(.A1(new_n8990_), .A2(new_n9310_), .ZN(new_n11018_));
  AOI22_X1   g10715(.A1(new_n797_), .A2(new_n11018_), .B1(new_n8991_), .B2(new_n11017_), .ZN(new_n11019_));
  NOR4_X1    g10716(.A1(new_n9781_), .A2(new_n10530_), .A3(new_n675_), .A4(new_n8990_), .ZN(new_n11020_));
  NAND2_X1   g10717(.A1(new_n11019_), .A2(new_n11020_), .ZN(new_n11021_));
  NOR2_X1    g10718(.A1(new_n10733_), .A2(new_n11021_), .ZN(new_n11022_));
  AOI21_X1   g10719(.A1(new_n11019_), .A2(new_n11020_), .B(new_n10734_), .ZN(new_n11023_));
  NOR2_X1    g10720(.A1(new_n11023_), .A2(new_n11022_), .ZN(new_n11024_));
  XNOR2_X1   g10721(.A1(new_n10733_), .A2(new_n11021_), .ZN(new_n11025_));
  MUX2_X1    g10722(.I0(new_n11025_), .I1(new_n11024_), .S(new_n11016_), .Z(new_n11026_));
  XNOR2_X1   g10723(.A1(new_n11015_), .A2(new_n11026_), .ZN(new_n11027_));
  NOR2_X1    g10724(.A1(new_n11015_), .A2(new_n11026_), .ZN(new_n11028_));
  INV_X1     g10725(.I(new_n11028_), .ZN(new_n11029_));
  NAND2_X1   g10726(.A1(new_n11015_), .A2(new_n11026_), .ZN(new_n11030_));
  NAND2_X1   g10727(.A1(new_n11029_), .A2(new_n11030_), .ZN(new_n11031_));
  NAND2_X1   g10728(.A1(new_n11031_), .A2(new_n11000_), .ZN(new_n11032_));
  OAI21_X1   g10729(.A1(new_n11000_), .A2(new_n11027_), .B(new_n11032_), .ZN(new_n11033_));
  XNOR2_X1   g10730(.A1(new_n11033_), .A2(new_n10998_), .ZN(new_n11034_));
  NOR2_X1    g10731(.A1(new_n11034_), .A2(new_n10951_), .ZN(new_n11035_));
  INV_X1     g10732(.I(new_n10951_), .ZN(new_n11036_));
  NAND2_X1   g10733(.A1(new_n11033_), .A2(new_n10998_), .ZN(new_n11037_));
  NOR2_X1    g10734(.A1(new_n11033_), .A2(new_n10998_), .ZN(new_n11038_));
  INV_X1     g10735(.I(new_n11038_), .ZN(new_n11039_));
  AOI21_X1   g10736(.A1(new_n11039_), .A2(new_n11037_), .B(new_n11036_), .ZN(new_n11040_));
  NOR2_X1    g10737(.A1(new_n11040_), .A2(new_n11035_), .ZN(new_n11041_));
  NOR2_X1    g10738(.A1(new_n10717_), .A2(new_n10727_), .ZN(new_n11042_));
  NOR2_X1    g10739(.A1(new_n11042_), .A2(new_n10726_), .ZN(new_n11043_));
  NOR2_X1    g10740(.A1(new_n10899_), .A2(new_n10897_), .ZN(new_n11044_));
  NOR2_X1    g10741(.A1(new_n11044_), .A2(new_n10898_), .ZN(new_n11045_));
  INV_X1     g10742(.I(new_n10790_), .ZN(new_n11046_));
  OAI21_X1   g10743(.A1(new_n10781_), .A2(new_n10793_), .B(new_n11046_), .ZN(new_n11047_));
  XOR2_X1    g10744(.A1(new_n11047_), .A2(new_n11045_), .Z(new_n11048_));
  NOR2_X1    g10745(.A1(new_n11048_), .A2(new_n11043_), .ZN(new_n11049_));
  INV_X1     g10746(.I(new_n11043_), .ZN(new_n11050_));
  INV_X1     g10747(.I(new_n11047_), .ZN(new_n11051_));
  NOR2_X1    g10748(.A1(new_n11051_), .A2(new_n11045_), .ZN(new_n11052_));
  INV_X1     g10749(.I(new_n11052_), .ZN(new_n11053_));
  NAND2_X1   g10750(.A1(new_n11051_), .A2(new_n11045_), .ZN(new_n11054_));
  AOI21_X1   g10751(.A1(new_n11053_), .A2(new_n11054_), .B(new_n11050_), .ZN(new_n11055_));
  NOR2_X1    g10752(.A1(new_n11055_), .A2(new_n11049_), .ZN(new_n11056_));
  NOR2_X1    g10753(.A1(new_n10801_), .A2(new_n10803_), .ZN(new_n11057_));
  NOR2_X1    g10754(.A1(new_n11057_), .A2(new_n10798_), .ZN(new_n11058_));
  AOI21_X1   g10755(.A1(new_n10774_), .A2(new_n10777_), .B(new_n10775_), .ZN(new_n11059_));
  INV_X1     g10756(.I(new_n11059_), .ZN(new_n11060_));
  AOI21_X1   g10757(.A1(new_n2533_), .A2(new_n5321_), .B(new_n10782_), .ZN(new_n11061_));
  OAI21_X1   g10758(.A1(new_n796_), .A2(new_n9553_), .B(new_n10719_), .ZN(new_n11062_));
  XOR2_X1    g10759(.A1(new_n11061_), .A2(new_n11062_), .Z(new_n11063_));
  NOR2_X1    g10760(.A1(new_n11063_), .A2(new_n10715_), .ZN(new_n11064_));
  INV_X1     g10761(.I(new_n11061_), .ZN(new_n11065_));
  NOR2_X1    g10762(.A1(new_n11065_), .A2(new_n11062_), .ZN(new_n11066_));
  INV_X1     g10763(.I(new_n11066_), .ZN(new_n11067_));
  NAND2_X1   g10764(.A1(new_n11065_), .A2(new_n11062_), .ZN(new_n11068_));
  AOI21_X1   g10765(.A1(new_n11067_), .A2(new_n11068_), .B(new_n10714_), .ZN(new_n11069_));
  NOR2_X1    g10766(.A1(new_n11069_), .A2(new_n11064_), .ZN(new_n11070_));
  AOI21_X1   g10767(.A1(new_n3126_), .A2(new_n6024_), .B(new_n10762_), .ZN(new_n11071_));
  INV_X1     g10768(.I(new_n11071_), .ZN(new_n11072_));
  NAND2_X1   g10769(.A1(new_n8755_), .A2(new_n1447_), .ZN(new_n11073_));
  NOR2_X1    g10770(.A1(new_n8755_), .A2(new_n1447_), .ZN(new_n11074_));
  NOR2_X1    g10771(.A1(\a[22] ), .A2(\a[48] ), .ZN(new_n11075_));
  AOI21_X1   g10772(.A1(new_n11073_), .A2(new_n11075_), .B(new_n11074_), .ZN(new_n11076_));
  NOR2_X1    g10773(.A1(new_n268_), .A2(new_n9310_), .ZN(new_n11077_));
  OAI21_X1   g10774(.A1(new_n10765_), .A2(new_n10767_), .B(new_n11077_), .ZN(new_n11078_));
  OAI21_X1   g10775(.A1(new_n10766_), .A2(new_n10768_), .B(new_n11078_), .ZN(new_n11079_));
  XNOR2_X1   g10776(.A1(new_n11079_), .A2(new_n11076_), .ZN(new_n11080_));
  AND2_X2    g10777(.A1(new_n11079_), .A2(new_n11076_), .Z(new_n11081_));
  NOR2_X1    g10778(.A1(new_n11079_), .A2(new_n11076_), .ZN(new_n11082_));
  OAI21_X1   g10779(.A1(new_n11081_), .A2(new_n11082_), .B(new_n11072_), .ZN(new_n11083_));
  OAI21_X1   g10780(.A1(new_n11072_), .A2(new_n11080_), .B(new_n11083_), .ZN(new_n11084_));
  INV_X1     g10781(.I(new_n11084_), .ZN(new_n11085_));
  XOR2_X1    g10782(.A1(new_n11070_), .A2(new_n11085_), .Z(new_n11086_));
  NAND2_X1   g10783(.A1(new_n11086_), .A2(new_n11060_), .ZN(new_n11087_));
  NOR2_X1    g10784(.A1(new_n11070_), .A2(new_n11085_), .ZN(new_n11088_));
  NAND2_X1   g10785(.A1(new_n11070_), .A2(new_n11085_), .ZN(new_n11089_));
  INV_X1     g10786(.I(new_n11089_), .ZN(new_n11090_));
  OAI21_X1   g10787(.A1(new_n11090_), .A2(new_n11088_), .B(new_n11059_), .ZN(new_n11091_));
  NAND2_X1   g10788(.A1(new_n11087_), .A2(new_n11091_), .ZN(new_n11092_));
  AND2_X2    g10789(.A1(new_n11058_), .A2(new_n11092_), .Z(new_n11093_));
  NOR2_X1    g10790(.A1(new_n11058_), .A2(new_n11092_), .ZN(new_n11094_));
  NOR2_X1    g10791(.A1(new_n11093_), .A2(new_n11094_), .ZN(new_n11095_));
  NOR2_X1    g10792(.A1(new_n11095_), .A2(new_n11056_), .ZN(new_n11096_));
  XNOR2_X1   g10793(.A1(new_n11058_), .A2(new_n11092_), .ZN(new_n11097_));
  INV_X1     g10794(.I(new_n11097_), .ZN(new_n11098_));
  AOI21_X1   g10795(.A1(new_n11056_), .A2(new_n11098_), .B(new_n11096_), .ZN(new_n11099_));
  XNOR2_X1   g10796(.A1(new_n11099_), .A2(new_n11041_), .ZN(new_n11100_));
  NOR2_X1    g10797(.A1(new_n11100_), .A2(new_n10949_), .ZN(new_n11101_));
  NOR2_X1    g10798(.A1(new_n11099_), .A2(new_n11041_), .ZN(new_n11102_));
  INV_X1     g10799(.I(new_n11102_), .ZN(new_n11103_));
  NAND2_X1   g10800(.A1(new_n11099_), .A2(new_n11041_), .ZN(new_n11104_));
  NAND2_X1   g10801(.A1(new_n11103_), .A2(new_n11104_), .ZN(new_n11105_));
  AOI21_X1   g10802(.A1(new_n10949_), .A2(new_n11105_), .B(new_n11101_), .ZN(new_n11106_));
  NAND2_X1   g10803(.A1(new_n10810_), .A2(new_n10812_), .ZN(new_n11107_));
  NAND2_X1   g10804(.A1(new_n11107_), .A2(new_n10809_), .ZN(new_n11108_));
  INV_X1     g10805(.I(new_n10742_), .ZN(new_n11109_));
  OAI21_X1   g10806(.A1(new_n10739_), .A2(new_n10743_), .B(new_n11109_), .ZN(new_n11110_));
  NOR2_X1    g10807(.A1(new_n359_), .A2(new_n9029_), .ZN(new_n11111_));
  OAI21_X1   g10808(.A1(new_n10834_), .A2(new_n10836_), .B(new_n11111_), .ZN(new_n11112_));
  OAI21_X1   g10809(.A1(new_n10835_), .A2(new_n10837_), .B(new_n11112_), .ZN(new_n11113_));
  INV_X1     g10810(.I(new_n11113_), .ZN(new_n11114_));
  NOR2_X1    g10811(.A1(new_n10830_), .A2(new_n10819_), .ZN(new_n11115_));
  NOR2_X1    g10812(.A1(new_n11115_), .A2(new_n10829_), .ZN(new_n11116_));
  XOR2_X1    g10813(.A1(new_n11116_), .A2(new_n11114_), .Z(new_n11117_));
  AND2_X2    g10814(.A1(new_n11117_), .A2(new_n11110_), .Z(new_n11118_));
  NOR2_X1    g10815(.A1(new_n11116_), .A2(new_n11114_), .ZN(new_n11119_));
  INV_X1     g10816(.I(new_n11119_), .ZN(new_n11120_));
  NAND2_X1   g10817(.A1(new_n11116_), .A2(new_n11114_), .ZN(new_n11121_));
  AOI21_X1   g10818(.A1(new_n11120_), .A2(new_n11121_), .B(new_n11110_), .ZN(new_n11122_));
  NOR2_X1    g10819(.A1(new_n11118_), .A2(new_n11122_), .ZN(new_n11123_));
  AOI21_X1   g10820(.A1(new_n10843_), .A2(new_n10847_), .B(new_n10845_), .ZN(new_n11124_));
  AOI21_X1   g10821(.A1(new_n10730_), .A2(new_n10753_), .B(new_n10752_), .ZN(new_n11125_));
  NOR2_X1    g10822(.A1(new_n11125_), .A2(new_n11124_), .ZN(new_n11126_));
  INV_X1     g10823(.I(new_n11126_), .ZN(new_n11127_));
  NAND2_X1   g10824(.A1(new_n11125_), .A2(new_n11124_), .ZN(new_n11128_));
  AOI21_X1   g10825(.A1(new_n11127_), .A2(new_n11128_), .B(new_n11123_), .ZN(new_n11129_));
  XNOR2_X1   g10826(.A1(new_n11125_), .A2(new_n11124_), .ZN(new_n11130_));
  NOR3_X1    g10827(.A1(new_n11130_), .A2(new_n11118_), .A3(new_n11122_), .ZN(new_n11131_));
  NOR2_X1    g10828(.A1(new_n11131_), .A2(new_n11129_), .ZN(new_n11132_));
  OAI21_X1   g10829(.A1(new_n10816_), .A2(new_n10869_), .B(new_n10871_), .ZN(new_n11133_));
  XOR2_X1    g10830(.A1(new_n11132_), .A2(new_n11133_), .Z(new_n11134_));
  INV_X1     g10831(.I(new_n11132_), .ZN(new_n11135_));
  INV_X1     g10832(.I(new_n11133_), .ZN(new_n11136_));
  NOR2_X1    g10833(.A1(new_n11135_), .A2(new_n11136_), .ZN(new_n11137_));
  INV_X1     g10834(.I(new_n11137_), .ZN(new_n11138_));
  NOR2_X1    g10835(.A1(new_n11132_), .A2(new_n11133_), .ZN(new_n11139_));
  INV_X1     g10836(.I(new_n11139_), .ZN(new_n11140_));
  AOI21_X1   g10837(.A1(new_n11138_), .A2(new_n11140_), .B(new_n11108_), .ZN(new_n11141_));
  AOI21_X1   g10838(.A1(new_n11134_), .A2(new_n11108_), .B(new_n11141_), .ZN(new_n11142_));
  XNOR2_X1   g10839(.A1(new_n11106_), .A2(new_n11142_), .ZN(new_n11143_));
  NOR2_X1    g10840(.A1(new_n11143_), .A2(new_n10948_), .ZN(new_n11144_));
  NOR2_X1    g10841(.A1(new_n11106_), .A2(new_n11142_), .ZN(new_n11145_));
  INV_X1     g10842(.I(new_n11145_), .ZN(new_n11146_));
  NAND2_X1   g10843(.A1(new_n11106_), .A2(new_n11142_), .ZN(new_n11147_));
  NAND2_X1   g10844(.A1(new_n11146_), .A2(new_n11147_), .ZN(new_n11148_));
  AOI21_X1   g10845(.A1(new_n10948_), .A2(new_n11148_), .B(new_n11144_), .ZN(new_n11149_));
  NOR2_X1    g10846(.A1(new_n11149_), .A2(new_n10946_), .ZN(new_n11150_));
  INV_X1     g10847(.I(new_n11150_), .ZN(new_n11151_));
  XOR2_X1    g10848(.A1(new_n10944_), .A2(new_n11151_), .Z(new_n11152_));
  XOR2_X1    g10849(.A1(new_n11152_), .A2(new_n10937_), .Z(\asquared[72] ));
  AOI21_X1   g10850(.A1(new_n11149_), .A2(new_n10946_), .B(new_n10938_), .ZN(new_n11154_));
  INV_X1     g10851(.I(new_n11154_), .ZN(new_n11155_));
  OAI21_X1   g10852(.A1(new_n10944_), .A2(new_n11155_), .B(new_n11151_), .ZN(new_n11156_));
  OAI21_X1   g10853(.A1(new_n10949_), .A2(new_n11102_), .B(new_n11104_), .ZN(new_n11157_));
  INV_X1     g10854(.I(new_n11157_), .ZN(new_n11158_));
  AOI21_X1   g10855(.A1(new_n11108_), .A2(new_n11140_), .B(new_n11137_), .ZN(new_n11159_));
  AOI21_X1   g10856(.A1(new_n11050_), .A2(new_n11054_), .B(new_n11052_), .ZN(new_n11160_));
  NOR2_X1    g10857(.A1(new_n885_), .A2(new_n6999_), .ZN(new_n11161_));
  NOR2_X1    g10858(.A1(new_n10290_), .A2(new_n1536_), .ZN(new_n11162_));
  NAND4_X1   g10859(.A1(new_n11162_), .A2(\a[20] ), .A3(\a[52] ), .A4(new_n11161_), .ZN(new_n11163_));
  AOI21_X1   g10860(.A1(new_n11163_), .A2(new_n8005_), .B(new_n1268_), .ZN(new_n11164_));
  NOR2_X1    g10861(.A1(new_n10290_), .A2(new_n1536_), .ZN(new_n11165_));
  INV_X1     g10862(.I(new_n11165_), .ZN(new_n11166_));
  NOR2_X1    g10863(.A1(new_n2368_), .A2(new_n5745_), .ZN(new_n11167_));
  INV_X1     g10864(.I(new_n11167_), .ZN(new_n11168_));
  NOR2_X1    g10865(.A1(new_n4975_), .A2(new_n11168_), .ZN(new_n11169_));
  XOR2_X1    g10866(.A1(new_n11169_), .A2(new_n800_), .Z(new_n11170_));
  XOR2_X1    g10867(.A1(new_n11170_), .A2(\a[56] ), .Z(new_n11171_));
  NAND2_X1   g10868(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n11172_));
  XNOR2_X1   g10869(.A1(new_n1773_), .A2(new_n11172_), .ZN(new_n11173_));
  NOR2_X1    g10870(.A1(new_n11171_), .A2(new_n11173_), .ZN(new_n11174_));
  INV_X1     g10871(.I(new_n11174_), .ZN(new_n11175_));
  NAND2_X1   g10872(.A1(new_n11171_), .A2(new_n11173_), .ZN(new_n11176_));
  AOI21_X1   g10873(.A1(new_n11175_), .A2(new_n11176_), .B(new_n11166_), .ZN(new_n11177_));
  XNOR2_X1   g10874(.A1(new_n11171_), .A2(new_n11173_), .ZN(new_n11178_));
  NOR2_X1    g10875(.A1(new_n11178_), .A2(new_n11165_), .ZN(new_n11179_));
  NOR2_X1    g10876(.A1(new_n11179_), .A2(new_n11177_), .ZN(new_n11180_));
  AOI22_X1   g10877(.A1(new_n10954_), .A2(new_n1220_), .B1(new_n8676_), .B2(new_n10956_), .ZN(new_n11181_));
  AOI22_X1   g10878(.A1(new_n597_), .A2(new_n9781_), .B1(new_n9549_), .B2(new_n5183_), .ZN(new_n11182_));
  NOR4_X1    g10879(.A1(new_n9784_), .A2(new_n797_), .A3(new_n364_), .A4(new_n9310_), .ZN(new_n11183_));
  NAND2_X1   g10880(.A1(new_n11182_), .A2(new_n11183_), .ZN(new_n11184_));
  NAND2_X1   g10881(.A1(new_n6030_), .A2(new_n2277_), .ZN(new_n11185_));
  NOR2_X1    g10882(.A1(new_n566_), .A2(new_n8990_), .ZN(new_n11186_));
  XOR2_X1    g10883(.A1(new_n11185_), .A2(new_n11186_), .Z(new_n11187_));
  XNOR2_X1   g10884(.A1(new_n11187_), .A2(new_n11184_), .ZN(new_n11188_));
  NOR2_X1    g10885(.A1(new_n11188_), .A2(new_n11181_), .ZN(new_n11189_));
  NOR2_X1    g10886(.A1(new_n11187_), .A2(new_n11184_), .ZN(new_n11190_));
  INV_X1     g10887(.I(new_n11190_), .ZN(new_n11191_));
  NAND2_X1   g10888(.A1(new_n11187_), .A2(new_n11184_), .ZN(new_n11192_));
  NAND2_X1   g10889(.A1(new_n11191_), .A2(new_n11192_), .ZN(new_n11193_));
  AOI21_X1   g10890(.A1(new_n11181_), .A2(new_n11193_), .B(new_n11189_), .ZN(new_n11194_));
  XOR2_X1    g10891(.A1(new_n11180_), .A2(new_n11194_), .Z(new_n11195_));
  NOR2_X1    g10892(.A1(new_n11195_), .A2(new_n11160_), .ZN(new_n11196_));
  INV_X1     g10893(.I(new_n11180_), .ZN(new_n11197_));
  NOR2_X1    g10894(.A1(new_n11197_), .A2(new_n11194_), .ZN(new_n11198_));
  INV_X1     g10895(.I(new_n11198_), .ZN(new_n11199_));
  NAND2_X1   g10896(.A1(new_n11197_), .A2(new_n11194_), .ZN(new_n11200_));
  NAND2_X1   g10897(.A1(new_n11199_), .A2(new_n11200_), .ZN(new_n11201_));
  AOI21_X1   g10898(.A1(new_n11160_), .A2(new_n11201_), .B(new_n11196_), .ZN(new_n11202_));
  NAND2_X1   g10899(.A1(new_n11128_), .A2(new_n11123_), .ZN(new_n11203_));
  NAND2_X1   g10900(.A1(new_n11203_), .A2(new_n11127_), .ZN(new_n11204_));
  AOI21_X1   g10901(.A1(new_n11110_), .A2(new_n11121_), .B(new_n11119_), .ZN(new_n11205_));
  AOI21_X1   g10902(.A1(new_n10530_), .A2(new_n9781_), .B(new_n11019_), .ZN(new_n11206_));
  INV_X1     g10903(.I(new_n11206_), .ZN(new_n11207_));
  OAI21_X1   g10904(.A1(new_n1021_), .A2(new_n8953_), .B(new_n10960_), .ZN(new_n11208_));
  AOI21_X1   g10905(.A1(new_n2752_), .A2(new_n5488_), .B(new_n10964_), .ZN(new_n11209_));
  XOR2_X1    g10906(.A1(new_n11208_), .A2(new_n11209_), .Z(new_n11210_));
  NOR2_X1    g10907(.A1(new_n11210_), .A2(new_n11207_), .ZN(new_n11211_));
  INV_X1     g10908(.I(new_n11209_), .ZN(new_n11212_));
  NOR2_X1    g10909(.A1(new_n11212_), .A2(new_n11208_), .ZN(new_n11213_));
  INV_X1     g10910(.I(new_n11213_), .ZN(new_n11214_));
  NAND2_X1   g10911(.A1(new_n11212_), .A2(new_n11208_), .ZN(new_n11215_));
  AOI21_X1   g10912(.A1(new_n11214_), .A2(new_n11215_), .B(new_n11206_), .ZN(new_n11216_));
  NOR2_X1    g10913(.A1(new_n11211_), .A2(new_n11216_), .ZN(new_n11217_));
  AOI21_X1   g10914(.A1(new_n787_), .A2(new_n2328_), .B(new_n8678_), .ZN(new_n11218_));
  NAND4_X1   g10915(.A1(new_n11218_), .A2(new_n1018_), .A3(new_n8246_), .A4(new_n10955_), .ZN(new_n11219_));
  AOI22_X1   g10916(.A1(new_n2533_), .A2(new_n7452_), .B1(new_n5488_), .B2(new_n3037_), .ZN(new_n11220_));
  NOR4_X1    g10917(.A1(new_n5742_), .A2(new_n2797_), .A3(new_n1916_), .A4(new_n5175_), .ZN(new_n11221_));
  NAND2_X1   g10918(.A1(new_n11220_), .A2(new_n11221_), .ZN(new_n11222_));
  NAND2_X1   g10919(.A1(new_n4372_), .A2(new_n5339_), .ZN(new_n11223_));
  NOR2_X1    g10920(.A1(new_n1339_), .A2(new_n6694_), .ZN(new_n11224_));
  XOR2_X1    g10921(.A1(new_n11223_), .A2(new_n11224_), .Z(new_n11225_));
  NOR2_X1    g10922(.A1(new_n11225_), .A2(new_n11222_), .ZN(new_n11226_));
  INV_X1     g10923(.I(new_n11226_), .ZN(new_n11227_));
  NAND2_X1   g10924(.A1(new_n11225_), .A2(new_n11222_), .ZN(new_n11228_));
  AOI21_X1   g10925(.A1(new_n11227_), .A2(new_n11228_), .B(new_n11219_), .ZN(new_n11229_));
  INV_X1     g10926(.I(new_n11219_), .ZN(new_n11230_));
  XNOR2_X1   g10927(.A1(new_n11225_), .A2(new_n11222_), .ZN(new_n11231_));
  NOR2_X1    g10928(.A1(new_n11231_), .A2(new_n11230_), .ZN(new_n11232_));
  NOR2_X1    g10929(.A1(new_n11232_), .A2(new_n11229_), .ZN(new_n11233_));
  XOR2_X1    g10930(.A1(new_n11217_), .A2(new_n11233_), .Z(new_n11234_));
  NOR2_X1    g10931(.A1(new_n11234_), .A2(new_n11205_), .ZN(new_n11235_));
  INV_X1     g10932(.I(new_n11217_), .ZN(new_n11236_));
  NOR2_X1    g10933(.A1(new_n11236_), .A2(new_n11233_), .ZN(new_n11237_));
  INV_X1     g10934(.I(new_n11237_), .ZN(new_n11238_));
  NAND2_X1   g10935(.A1(new_n11236_), .A2(new_n11233_), .ZN(new_n11239_));
  NAND2_X1   g10936(.A1(new_n11238_), .A2(new_n11239_), .ZN(new_n11240_));
  AOI21_X1   g10937(.A1(new_n11205_), .A2(new_n11240_), .B(new_n11235_), .ZN(new_n11241_));
  XNOR2_X1   g10938(.A1(new_n11204_), .A2(new_n11241_), .ZN(new_n11242_));
  NOR2_X1    g10939(.A1(new_n11242_), .A2(new_n11202_), .ZN(new_n11243_));
  INV_X1     g10940(.I(new_n11202_), .ZN(new_n11244_));
  NOR2_X1    g10941(.A1(new_n11204_), .A2(new_n11241_), .ZN(new_n11245_));
  INV_X1     g10942(.I(new_n11245_), .ZN(new_n11246_));
  NAND2_X1   g10943(.A1(new_n11204_), .A2(new_n11241_), .ZN(new_n11247_));
  AOI21_X1   g10944(.A1(new_n11246_), .A2(new_n11247_), .B(new_n11244_), .ZN(new_n11248_));
  NOR2_X1    g10945(.A1(new_n11243_), .A2(new_n11248_), .ZN(new_n11249_));
  INV_X1     g10946(.I(new_n11249_), .ZN(new_n11250_));
  INV_X1     g10947(.I(new_n10953_), .ZN(new_n11251_));
  AOI21_X1   g10948(.A1(new_n11251_), .A2(new_n10995_), .B(new_n10994_), .ZN(new_n11252_));
  AOI21_X1   g10949(.A1(new_n10714_), .A2(new_n11068_), .B(new_n11066_), .ZN(new_n11253_));
  NAND2_X1   g10950(.A1(new_n10987_), .A2(new_n10989_), .ZN(new_n11254_));
  NAND2_X1   g10951(.A1(new_n11254_), .A2(new_n10986_), .ZN(new_n11255_));
  INV_X1     g10952(.I(new_n11255_), .ZN(new_n11256_));
  INV_X1     g10953(.I(new_n11005_), .ZN(new_n11257_));
  NAND2_X1   g10954(.A1(new_n11012_), .A2(new_n11257_), .ZN(new_n11258_));
  NAND2_X1   g10955(.A1(new_n11258_), .A2(new_n11011_), .ZN(new_n11259_));
  XOR2_X1    g10956(.A1(new_n11259_), .A2(new_n11256_), .Z(new_n11260_));
  NOR2_X1    g10957(.A1(new_n11260_), .A2(new_n11253_), .ZN(new_n11261_));
  INV_X1     g10958(.I(new_n11253_), .ZN(new_n11262_));
  INV_X1     g10959(.I(new_n11259_), .ZN(new_n11263_));
  NOR2_X1    g10960(.A1(new_n11263_), .A2(new_n11256_), .ZN(new_n11264_));
  NOR2_X1    g10961(.A1(new_n11259_), .A2(new_n11255_), .ZN(new_n11265_));
  NOR2_X1    g10962(.A1(new_n11264_), .A2(new_n11265_), .ZN(new_n11266_));
  NOR2_X1    g10963(.A1(new_n11266_), .A2(new_n11262_), .ZN(new_n11267_));
  NOR2_X1    g10964(.A1(new_n11267_), .A2(new_n11261_), .ZN(new_n11268_));
  INV_X1     g10965(.I(new_n10970_), .ZN(new_n11269_));
  AOI21_X1   g10966(.A1(new_n10973_), .A2(new_n11269_), .B(new_n10969_), .ZN(new_n11270_));
  INV_X1     g10967(.I(new_n11270_), .ZN(new_n11271_));
  AOI21_X1   g10968(.A1(new_n2690_), .A2(new_n5173_), .B(new_n10977_), .ZN(new_n11272_));
  AOI21_X1   g10969(.A1(new_n3981_), .A2(new_n6024_), .B(new_n10980_), .ZN(new_n11273_));
  NAND2_X1   g10970(.A1(new_n7482_), .A2(new_n1441_), .ZN(new_n11274_));
  NOR2_X1    g10971(.A1(new_n7482_), .A2(new_n1441_), .ZN(new_n11275_));
  NOR2_X1    g10972(.A1(\a[23] ), .A2(\a[48] ), .ZN(new_n11276_));
  AOI21_X1   g10973(.A1(new_n11274_), .A2(new_n11276_), .B(new_n11275_), .ZN(new_n11277_));
  XNOR2_X1   g10974(.A1(new_n11273_), .A2(new_n11277_), .ZN(new_n11278_));
  INV_X1     g10975(.I(new_n11273_), .ZN(new_n11279_));
  INV_X1     g10976(.I(new_n11277_), .ZN(new_n11280_));
  NOR2_X1    g10977(.A1(new_n11279_), .A2(new_n11280_), .ZN(new_n11281_));
  NOR2_X1    g10978(.A1(new_n11273_), .A2(new_n11277_), .ZN(new_n11282_));
  NOR2_X1    g10979(.A1(new_n11281_), .A2(new_n11282_), .ZN(new_n11283_));
  MUX2_X1    g10980(.I0(new_n11283_), .I1(new_n11278_), .S(new_n11272_), .Z(new_n11284_));
  AOI21_X1   g10981(.A1(new_n1798_), .A2(new_n6777_), .B(new_n11003_), .ZN(new_n11285_));
  NOR4_X1    g10982(.A1(new_n2868_), .A2(new_n3371_), .A3(new_n3837_), .A4(new_n3804_), .ZN(new_n11286_));
  INV_X1     g10983(.I(new_n11286_), .ZN(new_n11287_));
  NAND2_X1   g10984(.A1(new_n11007_), .A2(new_n3393_), .ZN(new_n11288_));
  NAND3_X1   g10985(.A1(new_n11288_), .A2(\a[9] ), .A3(\a[62] ), .ZN(new_n11289_));
  OAI21_X1   g10986(.A1(new_n3393_), .A2(new_n11007_), .B(new_n11289_), .ZN(new_n11290_));
  XOR2_X1    g10987(.A1(new_n11290_), .A2(new_n11287_), .Z(new_n11291_));
  INV_X1     g10988(.I(new_n11290_), .ZN(new_n11292_));
  NOR2_X1    g10989(.A1(new_n11292_), .A2(new_n11287_), .ZN(new_n11293_));
  NOR2_X1    g10990(.A1(new_n11290_), .A2(new_n11286_), .ZN(new_n11294_));
  NOR2_X1    g10991(.A1(new_n11293_), .A2(new_n11294_), .ZN(new_n11295_));
  MUX2_X1    g10992(.I0(new_n11295_), .I1(new_n11291_), .S(new_n11285_), .Z(new_n11296_));
  XOR2_X1    g10993(.A1(new_n11284_), .A2(new_n11296_), .Z(new_n11297_));
  NAND2_X1   g10994(.A1(new_n11297_), .A2(new_n11271_), .ZN(new_n11298_));
  NOR2_X1    g10995(.A1(new_n11284_), .A2(new_n11296_), .ZN(new_n11299_));
  INV_X1     g10996(.I(new_n11299_), .ZN(new_n11300_));
  NAND2_X1   g10997(.A1(new_n11284_), .A2(new_n11296_), .ZN(new_n11301_));
  NAND2_X1   g10998(.A1(new_n11300_), .A2(new_n11301_), .ZN(new_n11302_));
  NAND2_X1   g10999(.A1(new_n11302_), .A2(new_n11270_), .ZN(new_n11303_));
  NAND2_X1   g11000(.A1(new_n11303_), .A2(new_n11298_), .ZN(new_n11304_));
  XOR2_X1    g11001(.A1(new_n11268_), .A2(new_n11304_), .Z(new_n11305_));
  NOR2_X1    g11002(.A1(new_n11305_), .A2(new_n11252_), .ZN(new_n11306_));
  INV_X1     g11003(.I(new_n11304_), .ZN(new_n11307_));
  NOR2_X1    g11004(.A1(new_n11307_), .A2(new_n11268_), .ZN(new_n11308_));
  INV_X1     g11005(.I(new_n11308_), .ZN(new_n11309_));
  NAND2_X1   g11006(.A1(new_n11307_), .A2(new_n11268_), .ZN(new_n11310_));
  NAND2_X1   g11007(.A1(new_n11309_), .A2(new_n11310_), .ZN(new_n11311_));
  AOI21_X1   g11008(.A1(new_n11252_), .A2(new_n11311_), .B(new_n11306_), .ZN(new_n11312_));
  NOR2_X1    g11009(.A1(new_n11250_), .A2(new_n11312_), .ZN(new_n11313_));
  INV_X1     g11010(.I(new_n11313_), .ZN(new_n11314_));
  NAND2_X1   g11011(.A1(new_n11250_), .A2(new_n11312_), .ZN(new_n11315_));
  AOI21_X1   g11012(.A1(new_n11314_), .A2(new_n11315_), .B(new_n11159_), .ZN(new_n11316_));
  INV_X1     g11013(.I(new_n11159_), .ZN(new_n11317_));
  XOR2_X1    g11014(.A1(new_n11249_), .A2(new_n11312_), .Z(new_n11318_));
  NOR2_X1    g11015(.A1(new_n11318_), .A2(new_n11317_), .ZN(new_n11319_));
  NOR2_X1    g11016(.A1(new_n11316_), .A2(new_n11319_), .ZN(new_n11320_));
  AOI21_X1   g11017(.A1(new_n11036_), .A2(new_n11037_), .B(new_n11038_), .ZN(new_n11321_));
  INV_X1     g11018(.I(new_n11093_), .ZN(new_n11322_));
  AOI21_X1   g11019(.A1(new_n11322_), .A2(new_n11056_), .B(new_n11094_), .ZN(new_n11323_));
  OAI21_X1   g11020(.A1(new_n11059_), .A2(new_n11088_), .B(new_n11089_), .ZN(new_n11324_));
  INV_X1     g11021(.I(new_n11324_), .ZN(new_n11325_));
  INV_X1     g11022(.I(new_n11030_), .ZN(new_n11326_));
  OAI21_X1   g11023(.A1(new_n11000_), .A2(new_n11326_), .B(new_n11029_), .ZN(new_n11327_));
  INV_X1     g11024(.I(new_n11023_), .ZN(new_n11328_));
  AOI21_X1   g11025(.A1(new_n11328_), .A2(new_n11016_), .B(new_n11022_), .ZN(new_n11329_));
  NOR2_X1    g11026(.A1(new_n11072_), .A2(new_n11082_), .ZN(new_n11330_));
  NOR2_X1    g11027(.A1(new_n11330_), .A2(new_n11081_), .ZN(new_n11331_));
  OAI22_X1   g11028(.A1(new_n6578_), .A2(new_n5174_), .B1(new_n3175_), .B2(new_n3734_), .ZN(new_n11332_));
  NOR2_X1    g11029(.A1(new_n2499_), .A2(new_n4501_), .ZN(new_n11333_));
  INV_X1     g11030(.I(new_n11333_), .ZN(new_n11334_));
  NOR4_X1    g11031(.A1(new_n11332_), .A2(new_n3126_), .A3(new_n5350_), .A4(new_n11334_), .ZN(new_n11335_));
  XOR2_X1    g11032(.A1(new_n11331_), .A2(new_n11335_), .Z(new_n11336_));
  NOR2_X1    g11033(.A1(new_n11336_), .A2(new_n11329_), .ZN(new_n11337_));
  INV_X1     g11034(.I(new_n11329_), .ZN(new_n11338_));
  INV_X1     g11035(.I(new_n11335_), .ZN(new_n11339_));
  NOR2_X1    g11036(.A1(new_n11331_), .A2(new_n11339_), .ZN(new_n11340_));
  INV_X1     g11037(.I(new_n11340_), .ZN(new_n11341_));
  NAND2_X1   g11038(.A1(new_n11331_), .A2(new_n11339_), .ZN(new_n11342_));
  AOI21_X1   g11039(.A1(new_n11341_), .A2(new_n11342_), .B(new_n11338_), .ZN(new_n11343_));
  NOR2_X1    g11040(.A1(new_n11337_), .A2(new_n11343_), .ZN(new_n11344_));
  XNOR2_X1   g11041(.A1(new_n11327_), .A2(new_n11344_), .ZN(new_n11345_));
  NOR2_X1    g11042(.A1(new_n11345_), .A2(new_n11325_), .ZN(new_n11346_));
  NOR2_X1    g11043(.A1(new_n11327_), .A2(new_n11344_), .ZN(new_n11347_));
  INV_X1     g11044(.I(new_n11347_), .ZN(new_n11348_));
  NAND2_X1   g11045(.A1(new_n11327_), .A2(new_n11344_), .ZN(new_n11349_));
  AOI21_X1   g11046(.A1(new_n11348_), .A2(new_n11349_), .B(new_n11324_), .ZN(new_n11350_));
  NOR2_X1    g11047(.A1(new_n11346_), .A2(new_n11350_), .ZN(new_n11351_));
  XOR2_X1    g11048(.A1(new_n11323_), .A2(new_n11351_), .Z(new_n11352_));
  NOR2_X1    g11049(.A1(new_n11352_), .A2(new_n11321_), .ZN(new_n11353_));
  INV_X1     g11050(.I(new_n11321_), .ZN(new_n11354_));
  INV_X1     g11051(.I(new_n11323_), .ZN(new_n11355_));
  NOR2_X1    g11052(.A1(new_n11355_), .A2(new_n11351_), .ZN(new_n11356_));
  INV_X1     g11053(.I(new_n11356_), .ZN(new_n11357_));
  NAND2_X1   g11054(.A1(new_n11355_), .A2(new_n11351_), .ZN(new_n11358_));
  AOI21_X1   g11055(.A1(new_n11357_), .A2(new_n11358_), .B(new_n11354_), .ZN(new_n11359_));
  NOR2_X1    g11056(.A1(new_n11359_), .A2(new_n11353_), .ZN(new_n11360_));
  XOR2_X1    g11057(.A1(new_n11320_), .A2(new_n11360_), .Z(new_n11361_));
  NOR2_X1    g11058(.A1(new_n11361_), .A2(new_n11158_), .ZN(new_n11362_));
  INV_X1     g11059(.I(new_n11320_), .ZN(new_n11363_));
  NOR2_X1    g11060(.A1(new_n11363_), .A2(new_n11360_), .ZN(new_n11364_));
  INV_X1     g11061(.I(new_n11364_), .ZN(new_n11365_));
  NAND2_X1   g11062(.A1(new_n11363_), .A2(new_n11360_), .ZN(new_n11366_));
  AOI21_X1   g11063(.A1(new_n11365_), .A2(new_n11366_), .B(new_n11157_), .ZN(new_n11367_));
  NOR2_X1    g11064(.A1(new_n11367_), .A2(new_n11362_), .ZN(new_n11368_));
  OAI21_X1   g11065(.A1(new_n10948_), .A2(new_n11145_), .B(new_n11147_), .ZN(new_n11369_));
  NAND2_X1   g11066(.A1(new_n11368_), .A2(new_n11369_), .ZN(new_n11370_));
  OR2_X2     g11067(.A1(new_n11368_), .A2(new_n11369_), .Z(new_n11371_));
  NAND2_X1   g11068(.A1(new_n11371_), .A2(new_n11370_), .ZN(new_n11372_));
  XOR2_X1    g11069(.A1(new_n11156_), .A2(new_n11372_), .Z(\asquared[73] ));
  INV_X1     g11070(.I(new_n11156_), .ZN(new_n11374_));
  NAND2_X1   g11071(.A1(new_n11374_), .A2(new_n11370_), .ZN(new_n11375_));
  NAND2_X1   g11072(.A1(new_n11375_), .A2(new_n11371_), .ZN(new_n11376_));
  OAI21_X1   g11073(.A1(new_n11158_), .A2(new_n11364_), .B(new_n11366_), .ZN(new_n11377_));
  OAI21_X1   g11074(.A1(new_n11159_), .A2(new_n11313_), .B(new_n11315_), .ZN(new_n11378_));
  OAI21_X1   g11075(.A1(new_n11321_), .A2(new_n11356_), .B(new_n11358_), .ZN(new_n11379_));
  OAI21_X1   g11076(.A1(new_n11160_), .A2(new_n11198_), .B(new_n11200_), .ZN(new_n11380_));
  INV_X1     g11077(.I(new_n11380_), .ZN(new_n11381_));
  INV_X1     g11078(.I(new_n11181_), .ZN(new_n11382_));
  AOI21_X1   g11079(.A1(new_n11382_), .A2(new_n11192_), .B(new_n11190_), .ZN(new_n11383_));
  INV_X1     g11080(.I(new_n11294_), .ZN(new_n11384_));
  AOI21_X1   g11081(.A1(new_n11285_), .A2(new_n11384_), .B(new_n11293_), .ZN(new_n11385_));
  NAND2_X1   g11082(.A1(new_n11230_), .A2(new_n11228_), .ZN(new_n11386_));
  NAND2_X1   g11083(.A1(new_n11386_), .A2(new_n11227_), .ZN(new_n11387_));
  XOR2_X1    g11084(.A1(new_n11387_), .A2(new_n11385_), .Z(new_n11388_));
  NOR2_X1    g11085(.A1(new_n11388_), .A2(new_n11383_), .ZN(new_n11389_));
  INV_X1     g11086(.I(new_n11383_), .ZN(new_n11390_));
  INV_X1     g11087(.I(new_n11387_), .ZN(new_n11391_));
  NOR2_X1    g11088(.A1(new_n11391_), .A2(new_n11385_), .ZN(new_n11392_));
  INV_X1     g11089(.I(new_n11392_), .ZN(new_n11393_));
  NAND2_X1   g11090(.A1(new_n11391_), .A2(new_n11385_), .ZN(new_n11394_));
  AOI21_X1   g11091(.A1(new_n11393_), .A2(new_n11394_), .B(new_n11390_), .ZN(new_n11395_));
  NOR2_X1    g11092(.A1(new_n11395_), .A2(new_n11389_), .ZN(new_n11396_));
  AOI21_X1   g11093(.A1(new_n11165_), .A2(new_n11176_), .B(new_n11174_), .ZN(new_n11397_));
  NOR2_X1    g11094(.A1(new_n11164_), .A2(new_n11162_), .ZN(new_n11398_));
  AOI21_X1   g11095(.A1(new_n797_), .A2(new_n9784_), .B(new_n11182_), .ZN(new_n11399_));
  NAND2_X1   g11096(.A1(new_n6030_), .A2(new_n2277_), .ZN(new_n11400_));
  NOR2_X1    g11097(.A1(new_n6030_), .A2(new_n2277_), .ZN(new_n11401_));
  NOR2_X1    g11098(.A1(\a[12] ), .A2(\a[60] ), .ZN(new_n11402_));
  AOI21_X1   g11099(.A1(new_n11400_), .A2(new_n11402_), .B(new_n11401_), .ZN(new_n11403_));
  XOR2_X1    g11100(.A1(new_n11399_), .A2(new_n11403_), .Z(new_n11404_));
  NAND2_X1   g11101(.A1(new_n11404_), .A2(new_n11398_), .ZN(new_n11405_));
  INV_X1     g11102(.I(new_n11398_), .ZN(new_n11406_));
  AND2_X2    g11103(.A1(new_n11399_), .A2(new_n11403_), .Z(new_n11407_));
  NOR2_X1    g11104(.A1(new_n11399_), .A2(new_n11403_), .ZN(new_n11408_));
  OAI21_X1   g11105(.A1(new_n11407_), .A2(new_n11408_), .B(new_n11406_), .ZN(new_n11409_));
  NAND2_X1   g11106(.A1(new_n11409_), .A2(new_n11405_), .ZN(new_n11410_));
  NAND2_X1   g11107(.A1(new_n1339_), .A2(new_n6694_), .ZN(new_n11411_));
  AOI21_X1   g11108(.A1(new_n4372_), .A2(new_n5339_), .B(new_n11411_), .ZN(new_n11412_));
  AOI21_X1   g11109(.A1(new_n4644_), .A2(new_n5340_), .B(new_n11412_), .ZN(new_n11413_));
  OAI21_X1   g11110(.A1(new_n1773_), .A2(new_n9375_), .B(new_n8941_), .ZN(new_n11414_));
  NAND2_X1   g11111(.A1(new_n11413_), .A2(new_n11414_), .ZN(new_n11415_));
  XOR2_X1    g11112(.A1(new_n11415_), .A2(\a[13] ), .Z(new_n11416_));
  XOR2_X1    g11113(.A1(new_n11416_), .A2(\a[60] ), .Z(new_n11417_));
  XOR2_X1    g11114(.A1(new_n11417_), .A2(new_n11410_), .Z(new_n11418_));
  NOR2_X1    g11115(.A1(new_n11418_), .A2(new_n11397_), .ZN(new_n11419_));
  INV_X1     g11116(.I(new_n11410_), .ZN(new_n11420_));
  NOR2_X1    g11117(.A1(new_n11420_), .A2(new_n11417_), .ZN(new_n11421_));
  INV_X1     g11118(.I(new_n11421_), .ZN(new_n11422_));
  NAND2_X1   g11119(.A1(new_n11420_), .A2(new_n11417_), .ZN(new_n11423_));
  NAND2_X1   g11120(.A1(new_n11422_), .A2(new_n11423_), .ZN(new_n11424_));
  AOI21_X1   g11121(.A1(new_n11397_), .A2(new_n11424_), .B(new_n11419_), .ZN(new_n11425_));
  XNOR2_X1   g11122(.A1(new_n11425_), .A2(new_n11396_), .ZN(new_n11426_));
  NOR2_X1    g11123(.A1(new_n11426_), .A2(new_n11381_), .ZN(new_n11427_));
  NOR2_X1    g11124(.A1(new_n11425_), .A2(new_n11396_), .ZN(new_n11428_));
  INV_X1     g11125(.I(new_n11428_), .ZN(new_n11429_));
  NAND2_X1   g11126(.A1(new_n11425_), .A2(new_n11396_), .ZN(new_n11430_));
  AOI21_X1   g11127(.A1(new_n11429_), .A2(new_n11430_), .B(new_n11380_), .ZN(new_n11431_));
  NOR2_X1    g11128(.A1(new_n11427_), .A2(new_n11431_), .ZN(new_n11432_));
  INV_X1     g11129(.I(new_n11432_), .ZN(new_n11433_));
  NOR2_X1    g11130(.A1(new_n9297_), .A2(new_n1955_), .ZN(new_n11434_));
  NAND4_X1   g11131(.A1(new_n11434_), .A2(\a[18] ), .A3(new_n9299_), .A4(\a[24] ), .ZN(new_n11435_));
  AOI21_X1   g11132(.A1(new_n11435_), .A2(new_n8005_), .B(new_n1342_), .ZN(new_n11436_));
  NOR3_X1    g11133(.A1(new_n11436_), .A2(new_n1276_), .A3(new_n6999_), .ZN(new_n11437_));
  NOR2_X1    g11134(.A1(new_n11436_), .A2(new_n11434_), .ZN(new_n11438_));
  INV_X1     g11135(.I(new_n11438_), .ZN(new_n11439_));
  NAND2_X1   g11136(.A1(new_n9297_), .A2(new_n1955_), .ZN(new_n11440_));
  NOR2_X1    g11137(.A1(new_n11439_), .A2(new_n11440_), .ZN(new_n11441_));
  NOR2_X1    g11138(.A1(new_n11441_), .A2(new_n11437_), .ZN(new_n11442_));
  AOI22_X1   g11139(.A1(new_n4538_), .A2(new_n7000_), .B1(new_n6777_), .B2(new_n4437_), .ZN(new_n11443_));
  NOR2_X1    g11140(.A1(new_n1674_), .A2(new_n6260_), .ZN(new_n11444_));
  NAND4_X1   g11141(.A1(new_n11443_), .A2(new_n1711_), .A3(new_n8056_), .A4(new_n11444_), .ZN(new_n11445_));
  NAND2_X1   g11142(.A1(\a[23] ), .A2(\a[50] ), .ZN(new_n11446_));
  NOR2_X1    g11143(.A1(new_n11446_), .A2(new_n3837_), .ZN(new_n11447_));
  XOR2_X1    g11144(.A1(new_n11447_), .A2(new_n675_), .Z(new_n11448_));
  XOR2_X1    g11145(.A1(new_n11448_), .A2(\a[62] ), .Z(new_n11449_));
  NOR2_X1    g11146(.A1(new_n11449_), .A2(new_n11445_), .ZN(new_n11450_));
  AND2_X2    g11147(.A1(new_n11449_), .A2(new_n11445_), .Z(new_n11451_));
  OAI21_X1   g11148(.A1(new_n11451_), .A2(new_n11450_), .B(new_n11442_), .ZN(new_n11452_));
  XNOR2_X1   g11149(.A1(new_n11449_), .A2(new_n11445_), .ZN(new_n11453_));
  OAI21_X1   g11150(.A1(new_n11442_), .A2(new_n11453_), .B(new_n11452_), .ZN(new_n11454_));
  NOR2_X1    g11151(.A1(new_n11265_), .A2(new_n11253_), .ZN(new_n11455_));
  NOR2_X1    g11152(.A1(new_n11455_), .A2(new_n11264_), .ZN(new_n11456_));
  AOI22_X1   g11153(.A1(new_n1718_), .A2(new_n8676_), .B1(new_n8674_), .B2(new_n1447_), .ZN(new_n11457_));
  NOR2_X1    g11154(.A1(new_n650_), .A2(new_n8085_), .ZN(new_n11458_));
  NAND4_X1   g11155(.A1(new_n11457_), .A2(new_n1021_), .A3(new_n8246_), .A4(new_n11458_), .ZN(new_n11459_));
  NAND2_X1   g11156(.A1(new_n2533_), .A2(new_n5980_), .ZN(new_n11460_));
  NAND2_X1   g11157(.A1(\a[17] ), .A2(\a[56] ), .ZN(new_n11461_));
  XNOR2_X1   g11158(.A1(new_n11460_), .A2(new_n11461_), .ZN(new_n11462_));
  NOR2_X1    g11159(.A1(new_n800_), .A2(new_n7216_), .ZN(new_n11463_));
  OAI21_X1   g11160(.A1(new_n4974_), .A2(new_n11167_), .B(new_n11463_), .ZN(new_n11464_));
  OAI21_X1   g11161(.A1(new_n4975_), .A2(new_n11168_), .B(new_n11464_), .ZN(new_n11465_));
  INV_X1     g11162(.I(new_n11465_), .ZN(new_n11466_));
  NOR2_X1    g11163(.A1(new_n11462_), .A2(new_n11466_), .ZN(new_n11467_));
  INV_X1     g11164(.I(new_n11462_), .ZN(new_n11468_));
  NOR2_X1    g11165(.A1(new_n11468_), .A2(new_n11465_), .ZN(new_n11469_));
  NOR2_X1    g11166(.A1(new_n11469_), .A2(new_n11467_), .ZN(new_n11470_));
  NOR2_X1    g11167(.A1(new_n11470_), .A2(new_n11459_), .ZN(new_n11471_));
  INV_X1     g11168(.I(new_n11459_), .ZN(new_n11472_));
  XOR2_X1    g11169(.A1(new_n11462_), .A2(new_n11465_), .Z(new_n11473_));
  NOR2_X1    g11170(.A1(new_n11473_), .A2(new_n11472_), .ZN(new_n11474_));
  NOR2_X1    g11171(.A1(new_n11471_), .A2(new_n11474_), .ZN(new_n11475_));
  XNOR2_X1   g11172(.A1(new_n11456_), .A2(new_n11475_), .ZN(new_n11476_));
  INV_X1     g11173(.I(new_n11476_), .ZN(new_n11477_));
  NOR2_X1    g11174(.A1(new_n11456_), .A2(new_n11475_), .ZN(new_n11478_));
  INV_X1     g11175(.I(new_n11478_), .ZN(new_n11479_));
  NAND2_X1   g11176(.A1(new_n11456_), .A2(new_n11475_), .ZN(new_n11480_));
  AOI21_X1   g11177(.A1(new_n11479_), .A2(new_n11480_), .B(new_n11454_), .ZN(new_n11481_));
  AOI21_X1   g11178(.A1(new_n11477_), .A2(new_n11454_), .B(new_n11481_), .ZN(new_n11482_));
  OAI21_X1   g11179(.A1(new_n11325_), .A2(new_n11347_), .B(new_n11349_), .ZN(new_n11483_));
  AOI21_X1   g11180(.A1(new_n11338_), .A2(new_n11342_), .B(new_n11340_), .ZN(new_n11484_));
  OAI21_X1   g11181(.A1(new_n3127_), .A2(new_n5881_), .B(new_n11332_), .ZN(new_n11485_));
  AOI21_X1   g11182(.A1(new_n1447_), .A2(new_n8245_), .B(new_n11218_), .ZN(new_n11486_));
  AOI21_X1   g11183(.A1(new_n2797_), .A2(new_n5742_), .B(new_n11220_), .ZN(new_n11487_));
  INV_X1     g11184(.I(new_n11487_), .ZN(new_n11488_));
  XOR2_X1    g11185(.A1(new_n11486_), .A2(new_n11488_), .Z(new_n11489_));
  AND2_X2    g11186(.A1(new_n11486_), .A2(new_n11487_), .Z(new_n11490_));
  NOR2_X1    g11187(.A1(new_n11486_), .A2(new_n11487_), .ZN(new_n11491_));
  OAI21_X1   g11188(.A1(new_n11490_), .A2(new_n11491_), .B(new_n11485_), .ZN(new_n11492_));
  OAI21_X1   g11189(.A1(new_n11485_), .A2(new_n11489_), .B(new_n11492_), .ZN(new_n11493_));
  NAND2_X1   g11190(.A1(new_n9781_), .A2(new_n1479_), .ZN(new_n11494_));
  NAND2_X1   g11191(.A1(\a[25] ), .A2(\a[48] ), .ZN(new_n11495_));
  XNOR2_X1   g11192(.A1(new_n11494_), .A2(new_n11495_), .ZN(new_n11496_));
  INV_X1     g11193(.I(new_n11496_), .ZN(new_n11497_));
  NOR2_X1    g11194(.A1(new_n7188_), .A2(new_n10484_), .ZN(new_n11498_));
  NOR4_X1    g11195(.A1(new_n2898_), .A2(new_n5321_), .A3(new_n2178_), .A4(new_n5004_), .ZN(new_n11499_));
  NAND2_X1   g11196(.A1(new_n11498_), .A2(new_n11499_), .ZN(new_n11500_));
  AOI22_X1   g11197(.A1(new_n3487_), .A2(new_n3838_), .B1(new_n4868_), .B2(new_n5339_), .ZN(new_n11501_));
  NOR2_X1    g11198(.A1(new_n3967_), .A2(new_n4706_), .ZN(new_n11502_));
  AOI21_X1   g11199(.A1(\a[35] ), .A2(\a[38] ), .B(new_n3838_), .ZN(new_n11503_));
  NOR3_X1    g11200(.A1(new_n11502_), .A2(new_n4869_), .A3(new_n11503_), .ZN(new_n11504_));
  NAND2_X1   g11201(.A1(new_n11504_), .A2(new_n11501_), .ZN(new_n11505_));
  NOR2_X1    g11202(.A1(new_n11505_), .A2(new_n11500_), .ZN(new_n11506_));
  AOI22_X1   g11203(.A1(new_n11498_), .A2(new_n11499_), .B1(new_n11504_), .B2(new_n11501_), .ZN(new_n11507_));
  OAI21_X1   g11204(.A1(new_n11506_), .A2(new_n11507_), .B(new_n11497_), .ZN(new_n11508_));
  XOR2_X1    g11205(.A1(new_n11505_), .A2(new_n11500_), .Z(new_n11509_));
  NAND2_X1   g11206(.A1(new_n11509_), .A2(new_n11496_), .ZN(new_n11510_));
  NAND2_X1   g11207(.A1(new_n11510_), .A2(new_n11508_), .ZN(new_n11511_));
  XOR2_X1    g11208(.A1(new_n11493_), .A2(new_n11511_), .Z(new_n11512_));
  NOR2_X1    g11209(.A1(new_n11512_), .A2(new_n11484_), .ZN(new_n11513_));
  INV_X1     g11210(.I(new_n11484_), .ZN(new_n11514_));
  INV_X1     g11211(.I(new_n11511_), .ZN(new_n11515_));
  NOR2_X1    g11212(.A1(new_n11515_), .A2(new_n11493_), .ZN(new_n11516_));
  INV_X1     g11213(.I(new_n11516_), .ZN(new_n11517_));
  NAND2_X1   g11214(.A1(new_n11515_), .A2(new_n11493_), .ZN(new_n11518_));
  AOI21_X1   g11215(.A1(new_n11517_), .A2(new_n11518_), .B(new_n11514_), .ZN(new_n11519_));
  NOR2_X1    g11216(.A1(new_n11513_), .A2(new_n11519_), .ZN(new_n11520_));
  XNOR2_X1   g11217(.A1(new_n11483_), .A2(new_n11520_), .ZN(new_n11521_));
  NOR2_X1    g11218(.A1(new_n11521_), .A2(new_n11482_), .ZN(new_n11522_));
  INV_X1     g11219(.I(new_n11482_), .ZN(new_n11523_));
  NOR2_X1    g11220(.A1(new_n11483_), .A2(new_n11520_), .ZN(new_n11524_));
  INV_X1     g11221(.I(new_n11524_), .ZN(new_n11525_));
  NAND2_X1   g11222(.A1(new_n11483_), .A2(new_n11520_), .ZN(new_n11526_));
  AOI21_X1   g11223(.A1(new_n11525_), .A2(new_n11526_), .B(new_n11523_), .ZN(new_n11527_));
  NOR2_X1    g11224(.A1(new_n11522_), .A2(new_n11527_), .ZN(new_n11528_));
  NOR2_X1    g11225(.A1(new_n11528_), .A2(new_n11433_), .ZN(new_n11529_));
  NOR3_X1    g11226(.A1(new_n11522_), .A2(new_n11432_), .A3(new_n11527_), .ZN(new_n11530_));
  NOR2_X1    g11227(.A1(new_n11529_), .A2(new_n11530_), .ZN(new_n11531_));
  XOR2_X1    g11228(.A1(new_n11528_), .A2(new_n11432_), .Z(new_n11532_));
  MUX2_X1    g11229(.I0(new_n11532_), .I1(new_n11531_), .S(new_n11379_), .Z(new_n11533_));
  OAI21_X1   g11230(.A1(new_n11244_), .A2(new_n11245_), .B(new_n11247_), .ZN(new_n11534_));
  INV_X1     g11231(.I(new_n11205_), .ZN(new_n11535_));
  AOI21_X1   g11232(.A1(new_n11535_), .A2(new_n11239_), .B(new_n11237_), .ZN(new_n11536_));
  OAI21_X1   g11233(.A1(new_n11270_), .A2(new_n11299_), .B(new_n11301_), .ZN(new_n11537_));
  AOI21_X1   g11234(.A1(new_n11206_), .A2(new_n11215_), .B(new_n11213_), .ZN(new_n11538_));
  INV_X1     g11235(.I(new_n11282_), .ZN(new_n11539_));
  AOI21_X1   g11236(.A1(new_n11272_), .A2(new_n11539_), .B(new_n11281_), .ZN(new_n11540_));
  NOR2_X1    g11237(.A1(new_n2870_), .A2(new_n4184_), .ZN(new_n11541_));
  NOR2_X1    g11238(.A1(new_n11541_), .A2(new_n6390_), .ZN(new_n11542_));
  NOR2_X1    g11239(.A1(new_n2655_), .A2(new_n4769_), .ZN(new_n11543_));
  NAND4_X1   g11240(.A1(new_n11542_), .A2(new_n3852_), .A3(new_n6579_), .A4(new_n11543_), .ZN(new_n11544_));
  XNOR2_X1   g11241(.A1(new_n11540_), .A2(new_n11544_), .ZN(new_n11545_));
  NOR2_X1    g11242(.A1(new_n11545_), .A2(new_n11538_), .ZN(new_n11546_));
  INV_X1     g11243(.I(new_n11538_), .ZN(new_n11547_));
  NOR2_X1    g11244(.A1(new_n11540_), .A2(new_n11544_), .ZN(new_n11548_));
  INV_X1     g11245(.I(new_n11548_), .ZN(new_n11549_));
  NAND2_X1   g11246(.A1(new_n11540_), .A2(new_n11544_), .ZN(new_n11550_));
  AOI21_X1   g11247(.A1(new_n11549_), .A2(new_n11550_), .B(new_n11547_), .ZN(new_n11551_));
  NOR2_X1    g11248(.A1(new_n11546_), .A2(new_n11551_), .ZN(new_n11552_));
  XNOR2_X1   g11249(.A1(new_n11552_), .A2(new_n11537_), .ZN(new_n11553_));
  NOR2_X1    g11250(.A1(new_n11553_), .A2(new_n11536_), .ZN(new_n11554_));
  NOR2_X1    g11251(.A1(new_n11552_), .A2(new_n11537_), .ZN(new_n11555_));
  INV_X1     g11252(.I(new_n11555_), .ZN(new_n11556_));
  NAND2_X1   g11253(.A1(new_n11552_), .A2(new_n11537_), .ZN(new_n11557_));
  NAND2_X1   g11254(.A1(new_n11556_), .A2(new_n11557_), .ZN(new_n11558_));
  AOI21_X1   g11255(.A1(new_n11536_), .A2(new_n11558_), .B(new_n11554_), .ZN(new_n11559_));
  OAI21_X1   g11256(.A1(new_n11252_), .A2(new_n11308_), .B(new_n11310_), .ZN(new_n11560_));
  XOR2_X1    g11257(.A1(new_n11559_), .A2(new_n11560_), .Z(new_n11561_));
  NAND2_X1   g11258(.A1(new_n11534_), .A2(new_n11561_), .ZN(new_n11562_));
  NAND2_X1   g11259(.A1(new_n11559_), .A2(new_n11560_), .ZN(new_n11563_));
  OR2_X2     g11260(.A1(new_n11559_), .A2(new_n11560_), .Z(new_n11564_));
  AND2_X2    g11261(.A1(new_n11564_), .A2(new_n11563_), .Z(new_n11565_));
  OAI21_X1   g11262(.A1(new_n11534_), .A2(new_n11565_), .B(new_n11562_), .ZN(new_n11566_));
  XOR2_X1    g11263(.A1(new_n11533_), .A2(new_n11566_), .Z(new_n11567_));
  NAND2_X1   g11264(.A1(new_n11533_), .A2(new_n11566_), .ZN(new_n11568_));
  NOR2_X1    g11265(.A1(new_n11533_), .A2(new_n11566_), .ZN(new_n11569_));
  INV_X1     g11266(.I(new_n11569_), .ZN(new_n11570_));
  AOI21_X1   g11267(.A1(new_n11570_), .A2(new_n11568_), .B(new_n11378_), .ZN(new_n11571_));
  AOI21_X1   g11268(.A1(new_n11378_), .A2(new_n11567_), .B(new_n11571_), .ZN(new_n11572_));
  XNOR2_X1   g11269(.A1(new_n11377_), .A2(new_n11572_), .ZN(new_n11573_));
  NOR2_X1    g11270(.A1(new_n11377_), .A2(new_n11572_), .ZN(new_n11574_));
  NAND2_X1   g11271(.A1(new_n11377_), .A2(new_n11572_), .ZN(new_n11575_));
  INV_X1     g11272(.I(new_n11575_), .ZN(new_n11576_));
  OAI21_X1   g11273(.A1(new_n11574_), .A2(new_n11576_), .B(new_n11376_), .ZN(new_n11577_));
  OAI21_X1   g11274(.A1(new_n11376_), .A2(new_n11573_), .B(new_n11577_), .ZN(\asquared[74] ));
  INV_X1     g11275(.I(new_n11574_), .ZN(new_n11579_));
  NAND3_X1   g11276(.A1(new_n11156_), .A2(new_n11368_), .A3(new_n11369_), .ZN(new_n11580_));
  AOI21_X1   g11277(.A1(new_n11378_), .A2(new_n11568_), .B(new_n11569_), .ZN(new_n11581_));
  NAND2_X1   g11278(.A1(new_n11534_), .A2(new_n11564_), .ZN(new_n11582_));
  NAND2_X1   g11279(.A1(new_n11582_), .A2(new_n11563_), .ZN(new_n11583_));
  INV_X1     g11280(.I(new_n11583_), .ZN(new_n11584_));
  OAI21_X1   g11281(.A1(new_n11536_), .A2(new_n11555_), .B(new_n11557_), .ZN(new_n11585_));
  AOI21_X1   g11282(.A1(new_n2978_), .A2(new_n7204_), .B(new_n11443_), .ZN(new_n11586_));
  NAND2_X1   g11283(.A1(new_n9781_), .A2(new_n1479_), .ZN(new_n11587_));
  NOR2_X1    g11284(.A1(new_n9781_), .A2(new_n1479_), .ZN(new_n11588_));
  NOR2_X1    g11285(.A1(\a[25] ), .A2(\a[48] ), .ZN(new_n11589_));
  AOI21_X1   g11286(.A1(new_n11587_), .A2(new_n11589_), .B(new_n11588_), .ZN(new_n11590_));
  XNOR2_X1   g11287(.A1(new_n11586_), .A2(new_n11590_), .ZN(new_n11591_));
  NOR2_X1    g11288(.A1(new_n11439_), .A2(new_n11591_), .ZN(new_n11592_));
  INV_X1     g11289(.I(new_n11586_), .ZN(new_n11593_));
  INV_X1     g11290(.I(new_n11590_), .ZN(new_n11594_));
  NOR2_X1    g11291(.A1(new_n11593_), .A2(new_n11594_), .ZN(new_n11595_));
  NOR2_X1    g11292(.A1(new_n11586_), .A2(new_n11590_), .ZN(new_n11596_));
  NOR2_X1    g11293(.A1(new_n11595_), .A2(new_n11596_), .ZN(new_n11597_));
  NOR2_X1    g11294(.A1(new_n11597_), .A2(new_n11438_), .ZN(new_n11598_));
  NOR2_X1    g11295(.A1(new_n11592_), .A2(new_n11598_), .ZN(new_n11599_));
  AOI21_X1   g11296(.A1(new_n1719_), .A2(new_n8245_), .B(new_n11457_), .ZN(new_n11600_));
  INV_X1     g11297(.I(new_n11600_), .ZN(new_n11601_));
  NOR2_X1    g11298(.A1(new_n2533_), .A2(new_n5980_), .ZN(new_n11602_));
  NAND2_X1   g11299(.A1(new_n885_), .A2(new_n7216_), .ZN(new_n11603_));
  AOI21_X1   g11300(.A1(new_n2533_), .A2(new_n5980_), .B(new_n11603_), .ZN(new_n11604_));
  NOR2_X1    g11301(.A1(new_n11604_), .A2(new_n11602_), .ZN(new_n11605_));
  INV_X1     g11302(.I(new_n11605_), .ZN(new_n11606_));
  AOI21_X1   g11303(.A1(new_n2898_), .A2(new_n5321_), .B(new_n11498_), .ZN(new_n11607_));
  XOR2_X1    g11304(.A1(new_n11607_), .A2(new_n11606_), .Z(new_n11608_));
  NOR2_X1    g11305(.A1(new_n11608_), .A2(new_n11601_), .ZN(new_n11609_));
  INV_X1     g11306(.I(new_n11607_), .ZN(new_n11610_));
  NOR2_X1    g11307(.A1(new_n11610_), .A2(new_n11606_), .ZN(new_n11611_));
  NOR2_X1    g11308(.A1(new_n11607_), .A2(new_n11605_), .ZN(new_n11612_));
  NOR2_X1    g11309(.A1(new_n11611_), .A2(new_n11612_), .ZN(new_n11613_));
  NOR2_X1    g11310(.A1(new_n11613_), .A2(new_n11600_), .ZN(new_n11614_));
  NOR2_X1    g11311(.A1(new_n11507_), .A2(new_n11496_), .ZN(new_n11615_));
  NOR2_X1    g11312(.A1(new_n11615_), .A2(new_n11506_), .ZN(new_n11616_));
  NOR3_X1    g11313(.A1(new_n11614_), .A2(new_n11609_), .A3(new_n11616_), .ZN(new_n11617_));
  NOR2_X1    g11314(.A1(new_n11614_), .A2(new_n11609_), .ZN(new_n11618_));
  NOR3_X1    g11315(.A1(new_n11618_), .A2(new_n11506_), .A3(new_n11615_), .ZN(new_n11619_));
  NOR2_X1    g11316(.A1(new_n11619_), .A2(new_n11617_), .ZN(new_n11620_));
  NOR2_X1    g11317(.A1(new_n11620_), .A2(new_n11599_), .ZN(new_n11621_));
  XOR2_X1    g11318(.A1(new_n11618_), .A2(new_n11616_), .Z(new_n11622_));
  INV_X1     g11319(.I(new_n11622_), .ZN(new_n11623_));
  AOI21_X1   g11320(.A1(new_n11599_), .A2(new_n11623_), .B(new_n11621_), .ZN(new_n11624_));
  INV_X1     g11321(.I(new_n11624_), .ZN(new_n11625_));
  NOR2_X1    g11322(.A1(new_n11491_), .A2(new_n11485_), .ZN(new_n11626_));
  NOR2_X1    g11323(.A1(new_n11626_), .A2(new_n11490_), .ZN(new_n11627_));
  INV_X1     g11324(.I(new_n11627_), .ZN(new_n11628_));
  NAND2_X1   g11325(.A1(new_n11446_), .A2(new_n3837_), .ZN(new_n11629_));
  NAND3_X1   g11326(.A1(new_n11629_), .A2(\a[11] ), .A3(\a[62] ), .ZN(new_n11630_));
  OAI21_X1   g11327(.A1(new_n3837_), .A2(new_n11446_), .B(new_n11630_), .ZN(new_n11631_));
  NAND2_X1   g11328(.A1(\a[12] ), .A2(\a[61] ), .ZN(new_n11632_));
  NAND2_X1   g11329(.A1(\a[13] ), .A2(\a[62] ), .ZN(new_n11633_));
  XNOR2_X1   g11330(.A1(new_n11632_), .A2(new_n11633_), .ZN(new_n11634_));
  XNOR2_X1   g11331(.A1(new_n11631_), .A2(new_n11634_), .ZN(new_n11635_));
  NOR2_X1    g11332(.A1(new_n2499_), .A2(new_n5004_), .ZN(new_n11636_));
  AOI22_X1   g11333(.A1(new_n2898_), .A2(new_n5742_), .B1(new_n9347_), .B2(new_n11636_), .ZN(new_n11637_));
  NOR2_X1    g11334(.A1(new_n2461_), .A2(new_n4770_), .ZN(new_n11638_));
  AOI21_X1   g11335(.A1(new_n9348_), .A2(new_n11638_), .B(new_n11637_), .ZN(new_n11639_));
  INV_X1     g11336(.I(new_n11639_), .ZN(new_n11640_));
  XNOR2_X1   g11337(.A1(new_n9347_), .A2(new_n11638_), .ZN(new_n11641_));
  OAI21_X1   g11338(.A1(new_n2499_), .A2(new_n5004_), .B(new_n11641_), .ZN(new_n11642_));
  AND2_X2    g11339(.A1(new_n11642_), .A2(new_n11640_), .Z(new_n11643_));
  XNOR2_X1   g11340(.A1(new_n11643_), .A2(new_n11635_), .ZN(new_n11644_));
  NAND2_X1   g11341(.A1(new_n11628_), .A2(new_n11644_), .ZN(new_n11645_));
  INV_X1     g11342(.I(new_n11643_), .ZN(new_n11646_));
  NOR2_X1    g11343(.A1(new_n11646_), .A2(new_n11635_), .ZN(new_n11647_));
  NAND2_X1   g11344(.A1(new_n11646_), .A2(new_n11635_), .ZN(new_n11648_));
  INV_X1     g11345(.I(new_n11648_), .ZN(new_n11649_));
  OAI21_X1   g11346(.A1(new_n11649_), .A2(new_n11647_), .B(new_n11627_), .ZN(new_n11650_));
  NAND2_X1   g11347(.A1(new_n11645_), .A2(new_n11650_), .ZN(new_n11651_));
  INV_X1     g11348(.I(new_n11651_), .ZN(new_n11652_));
  NAND2_X1   g11349(.A1(new_n3981_), .A2(new_n5173_), .ZN(new_n11653_));
  NAND2_X1   g11350(.A1(\a[11] ), .A2(\a[63] ), .ZN(new_n11654_));
  XNOR2_X1   g11351(.A1(new_n11653_), .A2(new_n11654_), .ZN(new_n11655_));
  NAND3_X1   g11352(.A1(new_n6732_), .A2(\a[25] ), .A3(\a[56] ), .ZN(new_n11656_));
  NOR2_X1    g11353(.A1(new_n5745_), .A2(new_n7216_), .ZN(new_n11657_));
  INV_X1     g11354(.I(new_n11657_), .ZN(new_n11658_));
  AOI21_X1   g11355(.A1(new_n4519_), .A2(new_n11658_), .B(new_n11656_), .ZN(new_n11659_));
  XOR2_X1    g11356(.A1(new_n11659_), .A2(new_n5348_), .Z(new_n11660_));
  AOI22_X1   g11357(.A1(new_n2533_), .A2(new_n8198_), .B1(new_n6030_), .B2(new_n3037_), .ZN(new_n11661_));
  NOR4_X1    g11358(.A1(new_n5980_), .A2(new_n2797_), .A3(new_n1916_), .A4(new_n5750_), .ZN(new_n11662_));
  NAND2_X1   g11359(.A1(new_n11661_), .A2(new_n11662_), .ZN(new_n11663_));
  NOR2_X1    g11360(.A1(new_n11660_), .A2(new_n11663_), .ZN(new_n11664_));
  INV_X1     g11361(.I(new_n11664_), .ZN(new_n11665_));
  NAND2_X1   g11362(.A1(new_n11660_), .A2(new_n11663_), .ZN(new_n11666_));
  AOI21_X1   g11363(.A1(new_n11665_), .A2(new_n11666_), .B(new_n11655_), .ZN(new_n11667_));
  XOR2_X1    g11364(.A1(new_n11660_), .A2(new_n11663_), .Z(new_n11668_));
  AOI21_X1   g11365(.A1(new_n11655_), .A2(new_n11668_), .B(new_n11667_), .ZN(new_n11669_));
  NOR2_X1    g11366(.A1(new_n6692_), .A2(new_n6999_), .ZN(new_n11670_));
  AOI22_X1   g11367(.A1(new_n4173_), .A2(new_n7204_), .B1(new_n11670_), .B2(new_n4538_), .ZN(new_n11671_));
  NOR2_X1    g11368(.A1(new_n1674_), .A2(new_n6692_), .ZN(new_n11672_));
  NAND4_X1   g11369(.A1(new_n11671_), .A2(new_n1710_), .A3(new_n7486_), .A4(new_n11672_), .ZN(new_n11673_));
  XOR2_X1    g11370(.A1(new_n3487_), .A2(new_n4321_), .Z(new_n11674_));
  NAND2_X1   g11371(.A1(\a[50] ), .A2(\a[51] ), .ZN(new_n11675_));
  XNOR2_X1   g11372(.A1(new_n1956_), .A2(new_n11675_), .ZN(new_n11676_));
  NOR2_X1    g11373(.A1(new_n11674_), .A2(new_n11676_), .ZN(new_n11677_));
  AND2_X2    g11374(.A1(new_n11674_), .A2(new_n11676_), .Z(new_n11678_));
  NOR2_X1    g11375(.A1(new_n11678_), .A2(new_n11677_), .ZN(new_n11679_));
  NOR2_X1    g11376(.A1(new_n11679_), .A2(new_n11673_), .ZN(new_n11680_));
  INV_X1     g11377(.I(new_n11673_), .ZN(new_n11681_));
  XNOR2_X1   g11378(.A1(new_n11674_), .A2(new_n11676_), .ZN(new_n11682_));
  NOR2_X1    g11379(.A1(new_n11682_), .A2(new_n11681_), .ZN(new_n11683_));
  NOR2_X1    g11380(.A1(new_n11680_), .A2(new_n11683_), .ZN(new_n11684_));
  XNOR2_X1   g11381(.A1(new_n11669_), .A2(new_n11684_), .ZN(new_n11685_));
  NOR2_X1    g11382(.A1(new_n11685_), .A2(new_n11652_), .ZN(new_n11686_));
  NOR2_X1    g11383(.A1(new_n11669_), .A2(new_n11684_), .ZN(new_n11687_));
  INV_X1     g11384(.I(new_n11687_), .ZN(new_n11688_));
  NAND2_X1   g11385(.A1(new_n11669_), .A2(new_n11684_), .ZN(new_n11689_));
  AOI21_X1   g11386(.A1(new_n11688_), .A2(new_n11689_), .B(new_n11651_), .ZN(new_n11690_));
  NOR2_X1    g11387(.A1(new_n11686_), .A2(new_n11690_), .ZN(new_n11691_));
  NOR2_X1    g11388(.A1(new_n11625_), .A2(new_n11691_), .ZN(new_n11692_));
  NAND2_X1   g11389(.A1(new_n11625_), .A2(new_n11691_), .ZN(new_n11693_));
  INV_X1     g11390(.I(new_n11693_), .ZN(new_n11694_));
  OAI21_X1   g11391(.A1(new_n11694_), .A2(new_n11692_), .B(new_n11585_), .ZN(new_n11695_));
  XOR2_X1    g11392(.A1(new_n11691_), .A2(new_n11624_), .Z(new_n11696_));
  OAI21_X1   g11393(.A1(new_n11585_), .A2(new_n11696_), .B(new_n11695_), .ZN(new_n11697_));
  NOR3_X1    g11394(.A1(new_n11451_), .A2(new_n11437_), .A3(new_n11441_), .ZN(new_n11698_));
  NOR2_X1    g11395(.A1(new_n11698_), .A2(new_n11450_), .ZN(new_n11699_));
  NAND2_X1   g11396(.A1(new_n11547_), .A2(new_n11550_), .ZN(new_n11700_));
  NAND2_X1   g11397(.A1(new_n11700_), .A2(new_n11549_), .ZN(new_n11701_));
  AOI21_X1   g11398(.A1(new_n3851_), .A2(new_n5592_), .B(new_n11542_), .ZN(new_n11702_));
  NOR2_X1    g11399(.A1(new_n11501_), .A2(new_n11502_), .ZN(new_n11703_));
  INV_X1     g11400(.I(new_n11703_), .ZN(new_n11704_));
  NOR2_X1    g11401(.A1(new_n9556_), .A2(new_n1019_), .ZN(new_n11705_));
  NOR4_X1    g11402(.A1(new_n8676_), .A2(new_n1719_), .A3(new_n650_), .A4(new_n8990_), .ZN(new_n11706_));
  NAND2_X1   g11403(.A1(new_n11705_), .A2(new_n11706_), .ZN(new_n11707_));
  NOR2_X1    g11404(.A1(new_n11707_), .A2(new_n11704_), .ZN(new_n11708_));
  INV_X1     g11405(.I(new_n11707_), .ZN(new_n11709_));
  NOR2_X1    g11406(.A1(new_n11709_), .A2(new_n11703_), .ZN(new_n11710_));
  OAI21_X1   g11407(.A1(new_n11710_), .A2(new_n11708_), .B(new_n11702_), .ZN(new_n11711_));
  INV_X1     g11408(.I(new_n11702_), .ZN(new_n11712_));
  XOR2_X1    g11409(.A1(new_n11707_), .A2(new_n11704_), .Z(new_n11713_));
  NAND2_X1   g11410(.A1(new_n11713_), .A2(new_n11712_), .ZN(new_n11714_));
  NAND2_X1   g11411(.A1(new_n11714_), .A2(new_n11711_), .ZN(new_n11715_));
  INV_X1     g11412(.I(new_n11715_), .ZN(new_n11716_));
  XOR2_X1    g11413(.A1(new_n11701_), .A2(new_n11716_), .Z(new_n11717_));
  NOR2_X1    g11414(.A1(new_n11717_), .A2(new_n11699_), .ZN(new_n11718_));
  INV_X1     g11415(.I(new_n11699_), .ZN(new_n11719_));
  INV_X1     g11416(.I(new_n11701_), .ZN(new_n11720_));
  NOR2_X1    g11417(.A1(new_n11720_), .A2(new_n11716_), .ZN(new_n11721_));
  NOR2_X1    g11418(.A1(new_n11701_), .A2(new_n11715_), .ZN(new_n11722_));
  NOR2_X1    g11419(.A1(new_n11721_), .A2(new_n11722_), .ZN(new_n11723_));
  NOR2_X1    g11420(.A1(new_n11723_), .A2(new_n11719_), .ZN(new_n11724_));
  NOR2_X1    g11421(.A1(new_n11724_), .A2(new_n11718_), .ZN(new_n11725_));
  NAND2_X1   g11422(.A1(new_n11480_), .A2(new_n11454_), .ZN(new_n11726_));
  NAND2_X1   g11423(.A1(new_n11726_), .A2(new_n11479_), .ZN(new_n11727_));
  INV_X1     g11424(.I(new_n11727_), .ZN(new_n11728_));
  AOI21_X1   g11425(.A1(new_n11514_), .A2(new_n11518_), .B(new_n11516_), .ZN(new_n11729_));
  NOR2_X1    g11426(.A1(new_n11728_), .A2(new_n11729_), .ZN(new_n11730_));
  INV_X1     g11427(.I(new_n11730_), .ZN(new_n11731_));
  NAND2_X1   g11428(.A1(new_n11728_), .A2(new_n11729_), .ZN(new_n11732_));
  AOI21_X1   g11429(.A1(new_n11731_), .A2(new_n11732_), .B(new_n11725_), .ZN(new_n11733_));
  XOR2_X1    g11430(.A1(new_n11727_), .A2(new_n11729_), .Z(new_n11734_));
  INV_X1     g11431(.I(new_n11734_), .ZN(new_n11735_));
  AOI21_X1   g11432(.A1(new_n11725_), .A2(new_n11735_), .B(new_n11733_), .ZN(new_n11736_));
  NOR2_X1    g11433(.A1(new_n11736_), .A2(new_n11697_), .ZN(new_n11737_));
  INV_X1     g11434(.I(new_n11737_), .ZN(new_n11738_));
  NAND2_X1   g11435(.A1(new_n11736_), .A2(new_n11697_), .ZN(new_n11739_));
  AOI21_X1   g11436(.A1(new_n11738_), .A2(new_n11739_), .B(new_n11584_), .ZN(new_n11740_));
  XNOR2_X1   g11437(.A1(new_n11736_), .A2(new_n11697_), .ZN(new_n11741_));
  NOR2_X1    g11438(.A1(new_n11583_), .A2(new_n11741_), .ZN(new_n11742_));
  NOR2_X1    g11439(.A1(new_n11740_), .A2(new_n11742_), .ZN(new_n11743_));
  INV_X1     g11440(.I(new_n11530_), .ZN(new_n11744_));
  AOI21_X1   g11441(.A1(new_n11379_), .A2(new_n11744_), .B(new_n11529_), .ZN(new_n11745_));
  OAI21_X1   g11442(.A1(new_n11381_), .A2(new_n11428_), .B(new_n11430_), .ZN(new_n11746_));
  OAI21_X1   g11443(.A1(new_n11523_), .A2(new_n11524_), .B(new_n11526_), .ZN(new_n11747_));
  NOR2_X1    g11444(.A1(new_n11406_), .A2(new_n11408_), .ZN(new_n11748_));
  NOR2_X1    g11445(.A1(new_n11748_), .A2(new_n11407_), .ZN(new_n11749_));
  INV_X1     g11446(.I(new_n11749_), .ZN(new_n11750_));
  NOR2_X1    g11447(.A1(new_n599_), .A2(new_n8990_), .ZN(new_n11751_));
  OAI21_X1   g11448(.A1(new_n11413_), .A2(new_n11414_), .B(new_n11751_), .ZN(new_n11752_));
  NAND2_X1   g11449(.A1(new_n11752_), .A2(new_n11415_), .ZN(new_n11753_));
  INV_X1     g11450(.I(new_n11467_), .ZN(new_n11754_));
  OAI21_X1   g11451(.A1(new_n11459_), .A2(new_n11469_), .B(new_n11754_), .ZN(new_n11755_));
  XOR2_X1    g11452(.A1(new_n11755_), .A2(new_n11753_), .Z(new_n11756_));
  NAND2_X1   g11453(.A1(new_n11755_), .A2(new_n11753_), .ZN(new_n11757_));
  NOR2_X1    g11454(.A1(new_n11755_), .A2(new_n11753_), .ZN(new_n11758_));
  INV_X1     g11455(.I(new_n11758_), .ZN(new_n11759_));
  AOI21_X1   g11456(.A1(new_n11759_), .A2(new_n11757_), .B(new_n11750_), .ZN(new_n11760_));
  AOI21_X1   g11457(.A1(new_n11750_), .A2(new_n11756_), .B(new_n11760_), .ZN(new_n11761_));
  OAI21_X1   g11458(.A1(new_n11397_), .A2(new_n11421_), .B(new_n11423_), .ZN(new_n11762_));
  INV_X1     g11459(.I(new_n11762_), .ZN(new_n11763_));
  AOI21_X1   g11460(.A1(new_n11390_), .A2(new_n11394_), .B(new_n11392_), .ZN(new_n11764_));
  NOR2_X1    g11461(.A1(new_n11763_), .A2(new_n11764_), .ZN(new_n11765_));
  INV_X1     g11462(.I(new_n11764_), .ZN(new_n11766_));
  NOR2_X1    g11463(.A1(new_n11762_), .A2(new_n11766_), .ZN(new_n11767_));
  NOR2_X1    g11464(.A1(new_n11765_), .A2(new_n11767_), .ZN(new_n11768_));
  NOR2_X1    g11465(.A1(new_n11768_), .A2(new_n11761_), .ZN(new_n11769_));
  XOR2_X1    g11466(.A1(new_n11762_), .A2(new_n11764_), .Z(new_n11770_));
  INV_X1     g11467(.I(new_n11770_), .ZN(new_n11771_));
  AOI21_X1   g11468(.A1(new_n11761_), .A2(new_n11771_), .B(new_n11769_), .ZN(new_n11772_));
  XNOR2_X1   g11469(.A1(new_n11747_), .A2(new_n11772_), .ZN(new_n11773_));
  INV_X1     g11470(.I(new_n11773_), .ZN(new_n11774_));
  NOR2_X1    g11471(.A1(new_n11747_), .A2(new_n11772_), .ZN(new_n11775_));
  INV_X1     g11472(.I(new_n11775_), .ZN(new_n11776_));
  NAND2_X1   g11473(.A1(new_n11747_), .A2(new_n11772_), .ZN(new_n11777_));
  AOI21_X1   g11474(.A1(new_n11776_), .A2(new_n11777_), .B(new_n11746_), .ZN(new_n11778_));
  AOI21_X1   g11475(.A1(new_n11774_), .A2(new_n11746_), .B(new_n11778_), .ZN(new_n11779_));
  XOR2_X1    g11476(.A1(new_n11745_), .A2(new_n11779_), .Z(new_n11780_));
  NOR2_X1    g11477(.A1(new_n11743_), .A2(new_n11780_), .ZN(new_n11781_));
  INV_X1     g11478(.I(new_n11745_), .ZN(new_n11782_));
  NOR2_X1    g11479(.A1(new_n11782_), .A2(new_n11779_), .ZN(new_n11783_));
  INV_X1     g11480(.I(new_n11783_), .ZN(new_n11784_));
  NAND2_X1   g11481(.A1(new_n11782_), .A2(new_n11779_), .ZN(new_n11785_));
  NAND2_X1   g11482(.A1(new_n11784_), .A2(new_n11785_), .ZN(new_n11786_));
  AOI21_X1   g11483(.A1(new_n11743_), .A2(new_n11786_), .B(new_n11781_), .ZN(new_n11787_));
  NOR2_X1    g11484(.A1(new_n11787_), .A2(new_n11581_), .ZN(new_n11788_));
  XOR2_X1    g11485(.A1(new_n11580_), .A2(new_n11788_), .Z(new_n11789_));
  XOR2_X1    g11486(.A1(new_n11789_), .A2(new_n11579_), .Z(\asquared[75] ));
  INV_X1     g11487(.I(new_n11788_), .ZN(new_n11791_));
  AOI21_X1   g11488(.A1(new_n11581_), .A2(new_n11787_), .B(new_n11579_), .ZN(new_n11792_));
  INV_X1     g11489(.I(new_n11792_), .ZN(new_n11793_));
  OAI21_X1   g11490(.A1(new_n11580_), .A2(new_n11793_), .B(new_n11791_), .ZN(new_n11794_));
  INV_X1     g11491(.I(new_n11794_), .ZN(new_n11795_));
  OAI21_X1   g11492(.A1(new_n11743_), .A2(new_n11783_), .B(new_n11785_), .ZN(new_n11796_));
  NAND2_X1   g11493(.A1(new_n11776_), .A2(new_n11746_), .ZN(new_n11797_));
  NAND2_X1   g11494(.A1(new_n11797_), .A2(new_n11777_), .ZN(new_n11798_));
  INV_X1     g11495(.I(new_n11798_), .ZN(new_n11799_));
  INV_X1     g11496(.I(new_n11765_), .ZN(new_n11800_));
  OAI21_X1   g11497(.A1(new_n11762_), .A2(new_n11766_), .B(new_n11761_), .ZN(new_n11801_));
  OAI21_X1   g11498(.A1(new_n11749_), .A2(new_n11758_), .B(new_n11757_), .ZN(new_n11802_));
  INV_X1     g11499(.I(new_n11802_), .ZN(new_n11803_));
  NOR2_X1    g11500(.A1(new_n5745_), .A2(new_n7727_), .ZN(new_n11804_));
  INV_X1     g11501(.I(new_n11804_), .ZN(new_n11805_));
  NOR2_X1    g11502(.A1(new_n4703_), .A2(new_n11805_), .ZN(new_n11806_));
  NOR4_X1    g11503(.A1(new_n885_), .A2(new_n1916_), .A3(new_n5745_), .A4(new_n7647_), .ZN(new_n11807_));
  NAND2_X1   g11504(.A1(new_n11806_), .A2(new_n11807_), .ZN(new_n11808_));
  AOI21_X1   g11505(.A1(new_n11808_), .A2(new_n8246_), .B(new_n1268_), .ZN(new_n11809_));
  NOR3_X1    g11506(.A1(new_n11809_), .A2(new_n885_), .A3(new_n7647_), .ZN(new_n11810_));
  NOR3_X1    g11507(.A1(new_n11809_), .A2(new_n4702_), .A3(new_n11804_), .ZN(new_n11811_));
  NOR2_X1    g11508(.A1(new_n11810_), .A2(new_n11811_), .ZN(new_n11812_));
  AOI22_X1   g11509(.A1(new_n1718_), .A2(new_n8991_), .B1(new_n8455_), .B2(new_n1447_), .ZN(new_n11813_));
  INV_X1     g11510(.I(new_n11813_), .ZN(new_n11814_));
  NAND4_X1   g11511(.A1(new_n9553_), .A2(\a[14] ), .A3(\a[61] ), .A4(new_n1021_), .ZN(new_n11815_));
  NOR2_X1    g11512(.A1(new_n11814_), .A2(new_n11815_), .ZN(new_n11816_));
  INV_X1     g11513(.I(new_n11816_), .ZN(new_n11817_));
  NOR2_X1    g11514(.A1(new_n7693_), .A2(new_n8199_), .ZN(new_n11818_));
  NOR2_X1    g11515(.A1(new_n11818_), .A2(new_n9042_), .ZN(new_n11819_));
  NOR4_X1    g11516(.A1(new_n5980_), .A2(new_n2690_), .A3(new_n2098_), .A4(new_n5750_), .ZN(new_n11820_));
  NAND2_X1   g11517(.A1(new_n11819_), .A2(new_n11820_), .ZN(new_n11821_));
  NOR2_X1    g11518(.A1(new_n11817_), .A2(new_n11821_), .ZN(new_n11822_));
  AOI21_X1   g11519(.A1(new_n11819_), .A2(new_n11820_), .B(new_n11816_), .ZN(new_n11823_));
  NOR2_X1    g11520(.A1(new_n11822_), .A2(new_n11823_), .ZN(new_n11824_));
  XOR2_X1    g11521(.A1(new_n11821_), .A2(new_n11816_), .Z(new_n11825_));
  MUX2_X1    g11522(.I0(new_n11825_), .I1(new_n11824_), .S(new_n11812_), .Z(new_n11826_));
  NAND4_X1   g11523(.A1(\a[12] ), .A2(\a[19] ), .A3(\a[56] ), .A4(\a[63] ), .ZN(new_n11827_));
  NAND2_X1   g11524(.A1(\a[30] ), .A2(\a[45] ), .ZN(new_n11828_));
  XNOR2_X1   g11525(.A1(new_n11827_), .A2(new_n11828_), .ZN(new_n11829_));
  INV_X1     g11526(.I(new_n11829_), .ZN(new_n11830_));
  NOR2_X1    g11527(.A1(new_n2368_), .A2(new_n6692_), .ZN(new_n11831_));
  XOR2_X1    g11528(.A1(new_n3966_), .A2(new_n4321_), .Z(new_n11832_));
  NAND2_X1   g11529(.A1(\a[13] ), .A2(\a[38] ), .ZN(new_n11833_));
  NAND2_X1   g11530(.A1(\a[37] ), .A2(\a[62] ), .ZN(new_n11834_));
  XNOR2_X1   g11531(.A1(new_n11833_), .A2(new_n11834_), .ZN(new_n11835_));
  NOR2_X1    g11532(.A1(new_n11832_), .A2(new_n11835_), .ZN(new_n11836_));
  AND2_X2    g11533(.A1(new_n11832_), .A2(new_n11835_), .Z(new_n11837_));
  OAI21_X1   g11534(.A1(new_n11837_), .A2(new_n11836_), .B(new_n11830_), .ZN(new_n11838_));
  XOR2_X1    g11535(.A1(new_n11832_), .A2(new_n11835_), .Z(new_n11839_));
  NAND2_X1   g11536(.A1(new_n11839_), .A2(new_n11829_), .ZN(new_n11840_));
  NAND2_X1   g11537(.A1(new_n11840_), .A2(new_n11838_), .ZN(new_n11841_));
  XOR2_X1    g11538(.A1(new_n11826_), .A2(new_n11841_), .Z(new_n11842_));
  INV_X1     g11539(.I(new_n11841_), .ZN(new_n11843_));
  NOR2_X1    g11540(.A1(new_n11826_), .A2(new_n11843_), .ZN(new_n11844_));
  NAND2_X1   g11541(.A1(new_n11826_), .A2(new_n11843_), .ZN(new_n11845_));
  INV_X1     g11542(.I(new_n11845_), .ZN(new_n11846_));
  OAI21_X1   g11543(.A1(new_n11846_), .A2(new_n11844_), .B(new_n11803_), .ZN(new_n11847_));
  OAI21_X1   g11544(.A1(new_n11803_), .A2(new_n11842_), .B(new_n11847_), .ZN(new_n11848_));
  AOI21_X1   g11545(.A1(new_n1719_), .A2(new_n8676_), .B(new_n11705_), .ZN(new_n11849_));
  NAND2_X1   g11546(.A1(new_n9347_), .A2(new_n11638_), .ZN(new_n11850_));
  AND2_X2    g11547(.A1(new_n11637_), .A2(new_n11850_), .Z(new_n11851_));
  AOI21_X1   g11548(.A1(new_n2797_), .A2(new_n5980_), .B(new_n11661_), .ZN(new_n11852_));
  XOR2_X1    g11549(.A1(new_n11851_), .A2(new_n11852_), .Z(new_n11853_));
  NAND2_X1   g11550(.A1(new_n11853_), .A2(new_n11849_), .ZN(new_n11854_));
  INV_X1     g11551(.I(new_n11849_), .ZN(new_n11855_));
  AND2_X2    g11552(.A1(new_n11851_), .A2(new_n11852_), .Z(new_n11856_));
  NOR2_X1    g11553(.A1(new_n11851_), .A2(new_n11852_), .ZN(new_n11857_));
  OAI21_X1   g11554(.A1(new_n11857_), .A2(new_n11856_), .B(new_n11855_), .ZN(new_n11858_));
  NAND2_X1   g11555(.A1(new_n11854_), .A2(new_n11858_), .ZN(new_n11859_));
  INV_X1     g11556(.I(new_n11678_), .ZN(new_n11860_));
  AOI21_X1   g11557(.A1(new_n11860_), .A2(new_n11681_), .B(new_n11677_), .ZN(new_n11861_));
  INV_X1     g11558(.I(new_n11655_), .ZN(new_n11862_));
  NAND2_X1   g11559(.A1(new_n11666_), .A2(new_n11862_), .ZN(new_n11863_));
  AOI21_X1   g11560(.A1(new_n11665_), .A2(new_n11863_), .B(new_n11861_), .ZN(new_n11864_));
  INV_X1     g11561(.I(new_n11861_), .ZN(new_n11865_));
  NAND2_X1   g11562(.A1(new_n11863_), .A2(new_n11665_), .ZN(new_n11866_));
  NOR2_X1    g11563(.A1(new_n11866_), .A2(new_n11865_), .ZN(new_n11867_));
  OAI21_X1   g11564(.A1(new_n11864_), .A2(new_n11867_), .B(new_n11859_), .ZN(new_n11868_));
  XOR2_X1    g11565(.A1(new_n11866_), .A2(new_n11861_), .Z(new_n11869_));
  OAI21_X1   g11566(.A1(new_n11869_), .A2(new_n11859_), .B(new_n11868_), .ZN(new_n11870_));
  NAND2_X1   g11567(.A1(new_n11848_), .A2(new_n11870_), .ZN(new_n11871_));
  NOR2_X1    g11568(.A1(new_n11848_), .A2(new_n11870_), .ZN(new_n11872_));
  INV_X1     g11569(.I(new_n11872_), .ZN(new_n11873_));
  AOI22_X1   g11570(.A1(new_n11873_), .A2(new_n11871_), .B1(new_n11800_), .B2(new_n11801_), .ZN(new_n11874_));
  NAND2_X1   g11571(.A1(new_n11800_), .A2(new_n11801_), .ZN(new_n11875_));
  XNOR2_X1   g11572(.A1(new_n11848_), .A2(new_n11870_), .ZN(new_n11876_));
  NOR2_X1    g11573(.A1(new_n11876_), .A2(new_n11875_), .ZN(new_n11877_));
  NOR2_X1    g11574(.A1(new_n11877_), .A2(new_n11874_), .ZN(new_n11878_));
  INV_X1     g11575(.I(new_n11596_), .ZN(new_n11879_));
  AOI21_X1   g11576(.A1(new_n11438_), .A2(new_n11879_), .B(new_n11595_), .ZN(new_n11880_));
  INV_X1     g11577(.I(new_n11708_), .ZN(new_n11881_));
  OAI21_X1   g11578(.A1(new_n11709_), .A2(new_n11703_), .B(new_n11702_), .ZN(new_n11882_));
  NAND2_X1   g11579(.A1(new_n11882_), .A2(new_n11881_), .ZN(new_n11883_));
  NOR2_X1    g11580(.A1(new_n11612_), .A2(new_n11601_), .ZN(new_n11884_));
  NOR2_X1    g11581(.A1(new_n11884_), .A2(new_n11611_), .ZN(new_n11885_));
  XOR2_X1    g11582(.A1(new_n11885_), .A2(new_n11883_), .Z(new_n11886_));
  NOR2_X1    g11583(.A1(new_n11886_), .A2(new_n11880_), .ZN(new_n11887_));
  INV_X1     g11584(.I(new_n11880_), .ZN(new_n11888_));
  INV_X1     g11585(.I(new_n11883_), .ZN(new_n11889_));
  NOR2_X1    g11586(.A1(new_n11889_), .A2(new_n11885_), .ZN(new_n11890_));
  INV_X1     g11587(.I(new_n11890_), .ZN(new_n11891_));
  NAND2_X1   g11588(.A1(new_n11889_), .A2(new_n11885_), .ZN(new_n11892_));
  AOI21_X1   g11589(.A1(new_n11891_), .A2(new_n11892_), .B(new_n11888_), .ZN(new_n11893_));
  NOR2_X1    g11590(.A1(new_n11887_), .A2(new_n11893_), .ZN(new_n11894_));
  NAND2_X1   g11591(.A1(new_n11652_), .A2(new_n11689_), .ZN(new_n11895_));
  NAND2_X1   g11592(.A1(new_n11895_), .A2(new_n11688_), .ZN(new_n11896_));
  AOI21_X1   g11593(.A1(new_n11628_), .A2(new_n11648_), .B(new_n11647_), .ZN(new_n11897_));
  AOI21_X1   g11594(.A1(new_n1769_), .A2(new_n7485_), .B(new_n11671_), .ZN(new_n11898_));
  INV_X1     g11595(.I(new_n11898_), .ZN(new_n11899_));
  AOI21_X1   g11596(.A1(new_n3487_), .A2(new_n10498_), .B(new_n6024_), .ZN(new_n11900_));
  AOI21_X1   g11597(.A1(new_n2543_), .A2(new_n3805_), .B(new_n6779_), .ZN(new_n11901_));
  XNOR2_X1   g11598(.A1(new_n11901_), .A2(new_n11900_), .ZN(new_n11902_));
  NOR2_X1    g11599(.A1(new_n11902_), .A2(new_n11899_), .ZN(new_n11903_));
  NOR2_X1    g11600(.A1(new_n11901_), .A2(new_n11900_), .ZN(new_n11904_));
  INV_X1     g11601(.I(new_n11904_), .ZN(new_n11905_));
  NAND2_X1   g11602(.A1(new_n11901_), .A2(new_n11900_), .ZN(new_n11906_));
  AOI21_X1   g11603(.A1(new_n11905_), .A2(new_n11906_), .B(new_n11898_), .ZN(new_n11907_));
  NOR2_X1    g11604(.A1(new_n11903_), .A2(new_n11907_), .ZN(new_n11908_));
  NAND2_X1   g11605(.A1(new_n3981_), .A2(new_n5173_), .ZN(new_n11909_));
  NOR2_X1    g11606(.A1(new_n3981_), .A2(new_n5173_), .ZN(new_n11910_));
  NOR2_X1    g11607(.A1(\a[11] ), .A2(\a[63] ), .ZN(new_n11911_));
  AOI21_X1   g11608(.A1(new_n11909_), .A2(new_n11911_), .B(new_n11910_), .ZN(new_n11912_));
  NOR2_X1    g11609(.A1(\a[33] ), .A2(\a[41] ), .ZN(new_n11913_));
  AOI22_X1   g11610(.A1(new_n11656_), .A2(new_n11913_), .B1(new_n11658_), .B2(new_n4519_), .ZN(new_n11914_));
  INV_X1     g11611(.I(new_n11914_), .ZN(new_n11915_));
  NAND2_X1   g11612(.A1(new_n11631_), .A2(new_n1220_), .ZN(new_n11916_));
  OAI21_X1   g11613(.A1(new_n9785_), .A2(new_n11634_), .B(new_n11916_), .ZN(new_n11917_));
  XOR2_X1    g11614(.A1(new_n11917_), .A2(new_n11915_), .Z(new_n11918_));
  INV_X1     g11615(.I(new_n11917_), .ZN(new_n11919_));
  NOR2_X1    g11616(.A1(new_n11919_), .A2(new_n11915_), .ZN(new_n11920_));
  NOR2_X1    g11617(.A1(new_n11917_), .A2(new_n11914_), .ZN(new_n11921_));
  NOR2_X1    g11618(.A1(new_n11920_), .A2(new_n11921_), .ZN(new_n11922_));
  MUX2_X1    g11619(.I0(new_n11922_), .I1(new_n11918_), .S(new_n11912_), .Z(new_n11923_));
  XNOR2_X1   g11620(.A1(new_n11923_), .A2(new_n11908_), .ZN(new_n11924_));
  NOR2_X1    g11621(.A1(new_n11924_), .A2(new_n11897_), .ZN(new_n11925_));
  INV_X1     g11622(.I(new_n11897_), .ZN(new_n11926_));
  NOR2_X1    g11623(.A1(new_n11923_), .A2(new_n11908_), .ZN(new_n11927_));
  INV_X1     g11624(.I(new_n11927_), .ZN(new_n11928_));
  NAND2_X1   g11625(.A1(new_n11923_), .A2(new_n11908_), .ZN(new_n11929_));
  AOI21_X1   g11626(.A1(new_n11928_), .A2(new_n11929_), .B(new_n11926_), .ZN(new_n11930_));
  NOR2_X1    g11627(.A1(new_n11925_), .A2(new_n11930_), .ZN(new_n11931_));
  NOR2_X1    g11628(.A1(new_n11931_), .A2(new_n11896_), .ZN(new_n11932_));
  INV_X1     g11629(.I(new_n11896_), .ZN(new_n11933_));
  INV_X1     g11630(.I(new_n11931_), .ZN(new_n11934_));
  NOR2_X1    g11631(.A1(new_n11934_), .A2(new_n11933_), .ZN(new_n11935_));
  NOR2_X1    g11632(.A1(new_n11935_), .A2(new_n11932_), .ZN(new_n11936_));
  NOR2_X1    g11633(.A1(new_n11936_), .A2(new_n11894_), .ZN(new_n11937_));
  XOR2_X1    g11634(.A1(new_n11931_), .A2(new_n11933_), .Z(new_n11938_));
  INV_X1     g11635(.I(new_n11938_), .ZN(new_n11939_));
  AOI21_X1   g11636(.A1(new_n11894_), .A2(new_n11939_), .B(new_n11937_), .ZN(new_n11940_));
  XOR2_X1    g11637(.A1(new_n11940_), .A2(new_n11878_), .Z(new_n11941_));
  INV_X1     g11638(.I(new_n11878_), .ZN(new_n11942_));
  NOR2_X1    g11639(.A1(new_n11940_), .A2(new_n11942_), .ZN(new_n11943_));
  NAND2_X1   g11640(.A1(new_n11940_), .A2(new_n11942_), .ZN(new_n11944_));
  INV_X1     g11641(.I(new_n11944_), .ZN(new_n11945_));
  OAI21_X1   g11642(.A1(new_n11943_), .A2(new_n11945_), .B(new_n11799_), .ZN(new_n11946_));
  OAI21_X1   g11643(.A1(new_n11799_), .A2(new_n11941_), .B(new_n11946_), .ZN(new_n11947_));
  AOI21_X1   g11644(.A1(new_n11585_), .A2(new_n11693_), .B(new_n11692_), .ZN(new_n11948_));
  INV_X1     g11645(.I(new_n11948_), .ZN(new_n11949_));
  INV_X1     g11646(.I(new_n11722_), .ZN(new_n11950_));
  AOI21_X1   g11647(.A1(new_n11719_), .A2(new_n11950_), .B(new_n11721_), .ZN(new_n11951_));
  INV_X1     g11648(.I(new_n11951_), .ZN(new_n11952_));
  INV_X1     g11649(.I(new_n11619_), .ZN(new_n11953_));
  AOI21_X1   g11650(.A1(new_n11953_), .A2(new_n11599_), .B(new_n11617_), .ZN(new_n11954_));
  NOR4_X1    g11651(.A1(new_n1313_), .A2(new_n1691_), .A3(new_n6260_), .A4(new_n6945_), .ZN(new_n11955_));
  NAND3_X1   g11652(.A1(new_n11955_), .A2(new_n2383_), .A3(new_n7000_), .ZN(new_n11956_));
  AOI21_X1   g11653(.A1(new_n11956_), .A2(new_n10288_), .B(new_n1773_), .ZN(new_n11957_));
  NOR2_X1    g11654(.A1(new_n7001_), .A2(new_n2384_), .ZN(new_n11959_));
  AOI22_X1   g11655(.A1(new_n2869_), .A2(new_n5321_), .B1(new_n3981_), .B2(new_n4771_), .ZN(new_n11960_));
  NOR2_X1    g11656(.A1(new_n2655_), .A2(new_n4770_), .ZN(new_n11961_));
  NAND4_X1   g11657(.A1(new_n11960_), .A2(new_n3852_), .A3(new_n5174_), .A4(new_n11961_), .ZN(new_n11962_));
  NOR2_X1    g11658(.A1(new_n1999_), .A2(new_n6055_), .ZN(new_n11963_));
  INV_X1     g11659(.I(new_n11963_), .ZN(new_n11964_));
  NOR2_X1    g11660(.A1(new_n3371_), .A2(new_n4414_), .ZN(new_n11965_));
  INV_X1     g11661(.I(new_n11965_), .ZN(new_n11966_));
  NOR2_X1    g11662(.A1(new_n11964_), .A2(new_n11966_), .ZN(new_n11967_));
  XOR2_X1    g11663(.A1(new_n11967_), .A2(new_n1215_), .Z(new_n11968_));
  XOR2_X1    g11664(.A1(new_n11968_), .A2(\a[55] ), .Z(new_n11969_));
  NOR2_X1    g11665(.A1(new_n11969_), .A2(new_n11962_), .ZN(new_n11970_));
  AND2_X2    g11666(.A1(new_n11969_), .A2(new_n11962_), .Z(new_n11971_));
  NOR2_X1    g11667(.A1(new_n11971_), .A2(new_n11970_), .ZN(new_n11972_));
  XNOR2_X1   g11668(.A1(new_n11969_), .A2(new_n11962_), .ZN(new_n11973_));
  MUX2_X1    g11669(.I0(new_n11973_), .I1(new_n11972_), .S(new_n11959_), .Z(new_n11974_));
  NOR2_X1    g11670(.A1(new_n11954_), .A2(new_n11974_), .ZN(new_n11975_));
  NAND2_X1   g11671(.A1(new_n11954_), .A2(new_n11974_), .ZN(new_n11976_));
  INV_X1     g11672(.I(new_n11976_), .ZN(new_n11977_));
  OAI21_X1   g11673(.A1(new_n11977_), .A2(new_n11975_), .B(new_n11952_), .ZN(new_n11978_));
  XOR2_X1    g11674(.A1(new_n11954_), .A2(new_n11974_), .Z(new_n11979_));
  NAND2_X1   g11675(.A1(new_n11979_), .A2(new_n11951_), .ZN(new_n11980_));
  NAND2_X1   g11676(.A1(new_n11980_), .A2(new_n11978_), .ZN(new_n11981_));
  INV_X1     g11677(.I(new_n11981_), .ZN(new_n11982_));
  NAND2_X1   g11678(.A1(new_n11732_), .A2(new_n11725_), .ZN(new_n11983_));
  NAND2_X1   g11679(.A1(new_n11983_), .A2(new_n11731_), .ZN(new_n11984_));
  XOR2_X1    g11680(.A1(new_n11984_), .A2(new_n11982_), .Z(new_n11985_));
  INV_X1     g11681(.I(new_n11985_), .ZN(new_n11986_));
  AOI21_X1   g11682(.A1(new_n11731_), .A2(new_n11983_), .B(new_n11982_), .ZN(new_n11987_));
  NOR2_X1    g11683(.A1(new_n11984_), .A2(new_n11981_), .ZN(new_n11988_));
  NOR2_X1    g11684(.A1(new_n11987_), .A2(new_n11988_), .ZN(new_n11989_));
  NOR2_X1    g11685(.A1(new_n11989_), .A2(new_n11949_), .ZN(new_n11990_));
  AOI21_X1   g11686(.A1(new_n11949_), .A2(new_n11986_), .B(new_n11990_), .ZN(new_n11991_));
  INV_X1     g11687(.I(new_n11991_), .ZN(new_n11992_));
  OAI21_X1   g11688(.A1(new_n11584_), .A2(new_n11737_), .B(new_n11739_), .ZN(new_n11993_));
  INV_X1     g11689(.I(new_n11993_), .ZN(new_n11994_));
  NOR2_X1    g11690(.A1(new_n11994_), .A2(new_n11992_), .ZN(new_n11995_));
  NOR2_X1    g11691(.A1(new_n11993_), .A2(new_n11991_), .ZN(new_n11996_));
  OAI21_X1   g11692(.A1(new_n11995_), .A2(new_n11996_), .B(new_n11947_), .ZN(new_n11997_));
  XOR2_X1    g11693(.A1(new_n11993_), .A2(new_n11992_), .Z(new_n11998_));
  OAI21_X1   g11694(.A1(new_n11947_), .A2(new_n11998_), .B(new_n11997_), .ZN(new_n11999_));
  XOR2_X1    g11695(.A1(new_n11999_), .A2(new_n11796_), .Z(new_n12000_));
  INV_X1     g11696(.I(new_n11999_), .ZN(new_n12001_));
  NOR2_X1    g11697(.A1(new_n12001_), .A2(new_n11796_), .ZN(new_n12002_));
  INV_X1     g11698(.I(new_n12002_), .ZN(new_n12003_));
  NAND2_X1   g11699(.A1(new_n12001_), .A2(new_n11796_), .ZN(new_n12004_));
  NAND2_X1   g11700(.A1(new_n12003_), .A2(new_n12004_), .ZN(new_n12005_));
  NAND2_X1   g11701(.A1(new_n11795_), .A2(new_n12005_), .ZN(new_n12006_));
  OAI21_X1   g11702(.A1(new_n11795_), .A2(new_n12000_), .B(new_n12006_), .ZN(\asquared[76] ));
  OAI21_X1   g11703(.A1(new_n11795_), .A2(new_n12002_), .B(new_n12004_), .ZN(new_n12008_));
  NOR2_X1    g11704(.A1(new_n11988_), .A2(new_n11948_), .ZN(new_n12009_));
  NOR2_X1    g11705(.A1(new_n12009_), .A2(new_n11987_), .ZN(new_n12010_));
  NOR2_X1    g11706(.A1(new_n11977_), .A2(new_n11951_), .ZN(new_n12011_));
  NOR2_X1    g11707(.A1(new_n12011_), .A2(new_n11975_), .ZN(new_n12012_));
  INV_X1     g11708(.I(new_n11823_), .ZN(new_n12013_));
  AOI21_X1   g11709(.A1(new_n11812_), .A2(new_n12013_), .B(new_n11822_), .ZN(new_n12014_));
  AOI21_X1   g11710(.A1(new_n1719_), .A2(new_n8996_), .B(new_n11813_), .ZN(new_n12015_));
  AOI21_X1   g11711(.A1(new_n3851_), .A2(new_n5173_), .B(new_n11960_), .ZN(new_n12016_));
  XNOR2_X1   g11712(.A1(new_n12016_), .A2(new_n12015_), .ZN(new_n12017_));
  NOR3_X1    g11713(.A1(new_n12017_), .A2(new_n11806_), .A3(new_n11809_), .ZN(new_n12018_));
  NOR2_X1    g11714(.A1(new_n11809_), .A2(new_n11806_), .ZN(new_n12019_));
  INV_X1     g11715(.I(new_n12015_), .ZN(new_n12020_));
  INV_X1     g11716(.I(new_n12016_), .ZN(new_n12021_));
  NOR2_X1    g11717(.A1(new_n12021_), .A2(new_n12020_), .ZN(new_n12022_));
  NOR2_X1    g11718(.A1(new_n12016_), .A2(new_n12015_), .ZN(new_n12023_));
  NOR2_X1    g11719(.A1(new_n12022_), .A2(new_n12023_), .ZN(new_n12024_));
  NOR2_X1    g11720(.A1(new_n12024_), .A2(new_n12019_), .ZN(new_n12025_));
  NOR2_X1    g11721(.A1(new_n12025_), .A2(new_n12018_), .ZN(new_n12026_));
  NOR2_X1    g11722(.A1(new_n11837_), .A2(new_n11829_), .ZN(new_n12027_));
  NOR2_X1    g11723(.A1(new_n12027_), .A2(new_n11836_), .ZN(new_n12028_));
  XOR2_X1    g11724(.A1(new_n12026_), .A2(new_n12028_), .Z(new_n12029_));
  NOR2_X1    g11725(.A1(new_n12029_), .A2(new_n12014_), .ZN(new_n12030_));
  INV_X1     g11726(.I(new_n12014_), .ZN(new_n12031_));
  INV_X1     g11727(.I(new_n12026_), .ZN(new_n12032_));
  NOR2_X1    g11728(.A1(new_n12032_), .A2(new_n12028_), .ZN(new_n12033_));
  INV_X1     g11729(.I(new_n12033_), .ZN(new_n12034_));
  NAND2_X1   g11730(.A1(new_n12032_), .A2(new_n12028_), .ZN(new_n12035_));
  AOI21_X1   g11731(.A1(new_n12034_), .A2(new_n12035_), .B(new_n12031_), .ZN(new_n12036_));
  NOR2_X1    g11732(.A1(new_n12036_), .A2(new_n12030_), .ZN(new_n12037_));
  NAND2_X1   g11733(.A1(new_n11892_), .A2(new_n11888_), .ZN(new_n12038_));
  AOI21_X1   g11734(.A1(new_n2383_), .A2(new_n7000_), .B(new_n11957_), .ZN(new_n12039_));
  NOR2_X1    g11735(.A1(new_n8993_), .A2(new_n4049_), .ZN(new_n12040_));
  NOR4_X1    g11736(.A1(new_n8996_), .A2(new_n1275_), .A3(new_n875_), .A4(new_n8453_), .ZN(new_n12041_));
  NAND2_X1   g11737(.A1(new_n12040_), .A2(new_n12041_), .ZN(new_n12042_));
  NAND2_X1   g11738(.A1(new_n2533_), .A2(new_n6280_), .ZN(new_n12043_));
  NOR2_X1    g11739(.A1(new_n1276_), .A2(new_n7647_), .ZN(new_n12044_));
  XOR2_X1    g11740(.A1(new_n12043_), .A2(new_n12044_), .Z(new_n12045_));
  XOR2_X1    g11741(.A1(new_n12042_), .A2(new_n12045_), .Z(new_n12046_));
  NAND2_X1   g11742(.A1(new_n12046_), .A2(new_n12039_), .ZN(new_n12047_));
  NOR2_X1    g11743(.A1(new_n12042_), .A2(new_n12045_), .ZN(new_n12048_));
  NAND2_X1   g11744(.A1(new_n12042_), .A2(new_n12045_), .ZN(new_n12049_));
  INV_X1     g11745(.I(new_n12049_), .ZN(new_n12050_));
  NOR2_X1    g11746(.A1(new_n12050_), .A2(new_n12048_), .ZN(new_n12051_));
  OAI21_X1   g11747(.A1(new_n12039_), .A2(new_n12051_), .B(new_n12047_), .ZN(new_n12052_));
  AOI22_X1   g11748(.A1(new_n3354_), .A2(new_n6030_), .B1(new_n8198_), .B2(new_n2690_), .ZN(new_n12053_));
  NOR2_X1    g11749(.A1(new_n2178_), .A2(new_n5750_), .ZN(new_n12054_));
  NAND4_X1   g11750(.A1(new_n12053_), .A2(new_n3175_), .A3(new_n5793_), .A4(new_n12054_), .ZN(new_n12055_));
  NOR2_X1    g11751(.A1(new_n4240_), .A2(new_n4769_), .ZN(new_n12056_));
  AOI22_X1   g11752(.A1(new_n3487_), .A2(new_n12056_), .B1(new_n4727_), .B2(new_n5350_), .ZN(new_n12057_));
  NOR4_X1    g11753(.A1(new_n3966_), .A2(new_n5592_), .A3(new_n3371_), .A4(new_n4769_), .ZN(new_n12058_));
  NAND2_X1   g11754(.A1(new_n12057_), .A2(new_n12058_), .ZN(new_n12059_));
  NAND2_X1   g11755(.A1(\a[51] ), .A2(\a[52] ), .ZN(new_n12060_));
  XNOR2_X1   g11756(.A1(new_n2276_), .A2(new_n12060_), .ZN(new_n12061_));
  NOR2_X1    g11757(.A1(new_n12059_), .A2(new_n12061_), .ZN(new_n12062_));
  INV_X1     g11758(.I(new_n12062_), .ZN(new_n12063_));
  NAND2_X1   g11759(.A1(new_n12059_), .A2(new_n12061_), .ZN(new_n12064_));
  AOI21_X1   g11760(.A1(new_n12063_), .A2(new_n12064_), .B(new_n12055_), .ZN(new_n12065_));
  INV_X1     g11761(.I(new_n12055_), .ZN(new_n12066_));
  XNOR2_X1   g11762(.A1(new_n12059_), .A2(new_n12061_), .ZN(new_n12067_));
  NOR2_X1    g11763(.A1(new_n12067_), .A2(new_n12066_), .ZN(new_n12068_));
  NOR2_X1    g11764(.A1(new_n12068_), .A2(new_n12065_), .ZN(new_n12069_));
  XNOR2_X1   g11765(.A1(new_n12052_), .A2(new_n12069_), .ZN(new_n12070_));
  AOI21_X1   g11766(.A1(new_n11891_), .A2(new_n12038_), .B(new_n12070_), .ZN(new_n12071_));
  NAND2_X1   g11767(.A1(new_n12038_), .A2(new_n11891_), .ZN(new_n12072_));
  NOR2_X1    g11768(.A1(new_n12052_), .A2(new_n12069_), .ZN(new_n12073_));
  INV_X1     g11769(.I(new_n12073_), .ZN(new_n12074_));
  NAND2_X1   g11770(.A1(new_n12052_), .A2(new_n12069_), .ZN(new_n12075_));
  AOI21_X1   g11771(.A1(new_n12074_), .A2(new_n12075_), .B(new_n12072_), .ZN(new_n12076_));
  NOR2_X1    g11772(.A1(new_n12071_), .A2(new_n12076_), .ZN(new_n12077_));
  NOR2_X1    g11773(.A1(new_n12077_), .A2(new_n12037_), .ZN(new_n12078_));
  INV_X1     g11774(.I(new_n12037_), .ZN(new_n12079_));
  INV_X1     g11775(.I(new_n12077_), .ZN(new_n12080_));
  NOR2_X1    g11776(.A1(new_n12080_), .A2(new_n12079_), .ZN(new_n12081_));
  NOR2_X1    g11777(.A1(new_n12081_), .A2(new_n12078_), .ZN(new_n12082_));
  NOR2_X1    g11778(.A1(new_n12082_), .A2(new_n12012_), .ZN(new_n12083_));
  INV_X1     g11779(.I(new_n12012_), .ZN(new_n12084_));
  XOR2_X1    g11780(.A1(new_n12077_), .A2(new_n12079_), .Z(new_n12085_));
  NOR2_X1    g11781(.A1(new_n12084_), .A2(new_n12085_), .ZN(new_n12086_));
  NOR2_X1    g11782(.A1(new_n12086_), .A2(new_n12083_), .ZN(new_n12087_));
  AOI21_X1   g11783(.A1(new_n11802_), .A2(new_n11845_), .B(new_n11844_), .ZN(new_n12088_));
  INV_X1     g11784(.I(new_n11971_), .ZN(new_n12089_));
  AOI21_X1   g11785(.A1(new_n12089_), .A2(new_n11959_), .B(new_n11970_), .ZN(new_n12090_));
  NOR2_X1    g11786(.A1(new_n1339_), .A2(new_n9310_), .ZN(new_n12091_));
  NAND3_X1   g11787(.A1(new_n12091_), .A2(\a[12] ), .A3(\a[56] ), .ZN(new_n12092_));
  AOI22_X1   g11788(.A1(\a[12] ), .A2(\a[19] ), .B1(\a[56] ), .B2(\a[63] ), .ZN(new_n12093_));
  NOR2_X1    g11789(.A1(\a[30] ), .A2(\a[45] ), .ZN(new_n12094_));
  AOI21_X1   g11790(.A1(new_n12092_), .A2(new_n12094_), .B(new_n12093_), .ZN(new_n12095_));
  AOI21_X1   g11791(.A1(new_n2690_), .A2(new_n5980_), .B(new_n11819_), .ZN(new_n12096_));
  OAI21_X1   g11792(.A1(new_n11963_), .A2(new_n11965_), .B(new_n9499_), .ZN(new_n12097_));
  OAI21_X1   g11793(.A1(new_n11964_), .A2(new_n11966_), .B(new_n12097_), .ZN(new_n12098_));
  XOR2_X1    g11794(.A1(new_n12096_), .A2(new_n12098_), .Z(new_n12099_));
  NAND2_X1   g11795(.A1(new_n12099_), .A2(new_n12095_), .ZN(new_n12100_));
  INV_X1     g11796(.I(new_n12095_), .ZN(new_n12101_));
  AND2_X2    g11797(.A1(new_n12096_), .A2(new_n12098_), .Z(new_n12102_));
  NOR2_X1    g11798(.A1(new_n12096_), .A2(new_n12098_), .ZN(new_n12103_));
  OAI21_X1   g11799(.A1(new_n12102_), .A2(new_n12103_), .B(new_n12101_), .ZN(new_n12104_));
  NAND2_X1   g11800(.A1(new_n12100_), .A2(new_n12104_), .ZN(new_n12105_));
  INV_X1     g11801(.I(new_n11831_), .ZN(new_n12106_));
  OAI21_X1   g11802(.A1(new_n12106_), .A2(new_n3967_), .B(new_n4321_), .ZN(new_n12107_));
  NOR2_X1    g11803(.A1(new_n3804_), .A2(new_n9029_), .ZN(new_n12108_));
  AOI21_X1   g11804(.A1(\a[13] ), .A2(new_n12108_), .B(new_n5600_), .ZN(new_n12109_));
  NAND2_X1   g11805(.A1(new_n12107_), .A2(new_n12109_), .ZN(new_n12110_));
  XOR2_X1    g11806(.A1(new_n12110_), .A2(\a[14] ), .Z(new_n12111_));
  XOR2_X1    g11807(.A1(new_n12111_), .A2(\a[62] ), .Z(new_n12112_));
  NOR2_X1    g11808(.A1(new_n12105_), .A2(new_n12112_), .ZN(new_n12113_));
  INV_X1     g11809(.I(new_n12113_), .ZN(new_n12114_));
  NAND2_X1   g11810(.A1(new_n12105_), .A2(new_n12112_), .ZN(new_n12115_));
  AOI21_X1   g11811(.A1(new_n12114_), .A2(new_n12115_), .B(new_n12090_), .ZN(new_n12116_));
  INV_X1     g11812(.I(new_n12090_), .ZN(new_n12117_));
  XNOR2_X1   g11813(.A1(new_n12105_), .A2(new_n12112_), .ZN(new_n12118_));
  NOR2_X1    g11814(.A1(new_n12118_), .A2(new_n12117_), .ZN(new_n12119_));
  INV_X1     g11815(.I(new_n11921_), .ZN(new_n12120_));
  AOI21_X1   g11816(.A1(new_n11912_), .A2(new_n12120_), .B(new_n11920_), .ZN(new_n12121_));
  INV_X1     g11817(.I(new_n12121_), .ZN(new_n12122_));
  NOR2_X1    g11818(.A1(new_n11855_), .A2(new_n11857_), .ZN(new_n12123_));
  NOR2_X1    g11819(.A1(new_n12123_), .A2(new_n11856_), .ZN(new_n12124_));
  AOI21_X1   g11820(.A1(new_n11898_), .A2(new_n11906_), .B(new_n11904_), .ZN(new_n12125_));
  XOR2_X1    g11821(.A1(new_n12124_), .A2(new_n12125_), .Z(new_n12126_));
  NAND2_X1   g11822(.A1(new_n12126_), .A2(new_n12122_), .ZN(new_n12127_));
  NOR2_X1    g11823(.A1(new_n12124_), .A2(new_n12125_), .ZN(new_n12128_));
  NAND2_X1   g11824(.A1(new_n12124_), .A2(new_n12125_), .ZN(new_n12129_));
  INV_X1     g11825(.I(new_n12129_), .ZN(new_n12130_));
  OAI21_X1   g11826(.A1(new_n12130_), .A2(new_n12128_), .B(new_n12121_), .ZN(new_n12131_));
  NAND2_X1   g11827(.A1(new_n12127_), .A2(new_n12131_), .ZN(new_n12132_));
  INV_X1     g11828(.I(new_n12132_), .ZN(new_n12133_));
  NOR3_X1    g11829(.A1(new_n12119_), .A2(new_n12133_), .A3(new_n12116_), .ZN(new_n12134_));
  NOR2_X1    g11830(.A1(new_n12119_), .A2(new_n12116_), .ZN(new_n12135_));
  NOR2_X1    g11831(.A1(new_n12135_), .A2(new_n12132_), .ZN(new_n12136_));
  NOR2_X1    g11832(.A1(new_n12136_), .A2(new_n12134_), .ZN(new_n12137_));
  NOR2_X1    g11833(.A1(new_n12137_), .A2(new_n12088_), .ZN(new_n12138_));
  INV_X1     g11834(.I(new_n12088_), .ZN(new_n12139_));
  XOR2_X1    g11835(.A1(new_n12135_), .A2(new_n12133_), .Z(new_n12140_));
  NOR2_X1    g11836(.A1(new_n12140_), .A2(new_n12139_), .ZN(new_n12141_));
  NOR2_X1    g11837(.A1(new_n12141_), .A2(new_n12138_), .ZN(new_n12142_));
  XNOR2_X1   g11838(.A1(new_n12087_), .A2(new_n12142_), .ZN(new_n12143_));
  NOR2_X1    g11839(.A1(new_n12087_), .A2(new_n12142_), .ZN(new_n12144_));
  NAND2_X1   g11840(.A1(new_n12087_), .A2(new_n12142_), .ZN(new_n12145_));
  INV_X1     g11841(.I(new_n12145_), .ZN(new_n12146_));
  OAI21_X1   g11842(.A1(new_n12144_), .A2(new_n12146_), .B(new_n12010_), .ZN(new_n12147_));
  OAI21_X1   g11843(.A1(new_n12010_), .A2(new_n12143_), .B(new_n12147_), .ZN(new_n12148_));
  OAI21_X1   g11844(.A1(new_n11799_), .A2(new_n11943_), .B(new_n11944_), .ZN(new_n12149_));
  AOI21_X1   g11845(.A1(new_n11875_), .A2(new_n11871_), .B(new_n11872_), .ZN(new_n12150_));
  INV_X1     g11846(.I(new_n11932_), .ZN(new_n12151_));
  AOI21_X1   g11847(.A1(new_n11894_), .A2(new_n12151_), .B(new_n11935_), .ZN(new_n12152_));
  OAI21_X1   g11848(.A1(new_n11897_), .A2(new_n11927_), .B(new_n11929_), .ZN(new_n12153_));
  NOR2_X1    g11849(.A1(new_n11867_), .A2(new_n11859_), .ZN(new_n12154_));
  NOR2_X1    g11850(.A1(new_n12154_), .A2(new_n11864_), .ZN(new_n12155_));
  NAND2_X1   g11851(.A1(new_n3981_), .A2(new_n5742_), .ZN(new_n12156_));
  NAND2_X1   g11852(.A1(\a[13] ), .A2(\a[63] ), .ZN(new_n12157_));
  XNOR2_X1   g11853(.A1(new_n12156_), .A2(new_n12157_), .ZN(new_n12158_));
  INV_X1     g11854(.I(new_n12158_), .ZN(new_n12159_));
  NOR2_X1    g11855(.A1(new_n7422_), .A2(new_n8953_), .ZN(new_n12160_));
  NOR2_X1    g11856(.A1(new_n12160_), .A2(new_n7009_), .ZN(new_n12161_));
  INV_X1     g11857(.I(new_n12161_), .ZN(new_n12162_));
  NOR4_X1    g11858(.A1(new_n12162_), .A2(new_n4538_), .A3(new_n7483_), .A4(new_n10175_), .ZN(new_n12163_));
  INV_X1     g11859(.I(new_n12163_), .ZN(new_n12164_));
  NOR2_X1    g11860(.A1(new_n2368_), .A2(new_n6694_), .ZN(new_n12165_));
  INV_X1     g11861(.I(new_n12165_), .ZN(new_n12166_));
  NOR2_X1    g11862(.A1(new_n5563_), .A2(new_n12166_), .ZN(new_n12167_));
  XOR2_X1    g11863(.A1(new_n12167_), .A2(new_n1339_), .Z(new_n12168_));
  XOR2_X1    g11864(.A1(new_n12168_), .A2(\a[57] ), .Z(new_n12169_));
  NOR2_X1    g11865(.A1(new_n12169_), .A2(new_n12164_), .ZN(new_n12170_));
  AND2_X2    g11866(.A1(new_n12169_), .A2(new_n12164_), .Z(new_n12171_));
  OAI21_X1   g11867(.A1(new_n12171_), .A2(new_n12170_), .B(new_n12159_), .ZN(new_n12172_));
  XOR2_X1    g11868(.A1(new_n12169_), .A2(new_n12164_), .Z(new_n12173_));
  NAND2_X1   g11869(.A1(new_n12173_), .A2(new_n12158_), .ZN(new_n12174_));
  NAND2_X1   g11870(.A1(new_n12174_), .A2(new_n12172_), .ZN(new_n12175_));
  XOR2_X1    g11871(.A1(new_n12175_), .A2(new_n12155_), .Z(new_n12176_));
  INV_X1     g11872(.I(new_n12176_), .ZN(new_n12177_));
  INV_X1     g11873(.I(new_n12175_), .ZN(new_n12178_));
  NOR2_X1    g11874(.A1(new_n12178_), .A2(new_n12155_), .ZN(new_n12179_));
  INV_X1     g11875(.I(new_n12179_), .ZN(new_n12180_));
  NAND2_X1   g11876(.A1(new_n12178_), .A2(new_n12155_), .ZN(new_n12181_));
  AOI21_X1   g11877(.A1(new_n12180_), .A2(new_n12181_), .B(new_n12153_), .ZN(new_n12182_));
  AOI21_X1   g11878(.A1(new_n12153_), .A2(new_n12177_), .B(new_n12182_), .ZN(new_n12183_));
  XOR2_X1    g11879(.A1(new_n12152_), .A2(new_n12183_), .Z(new_n12184_));
  NOR2_X1    g11880(.A1(new_n12184_), .A2(new_n12150_), .ZN(new_n12185_));
  INV_X1     g11881(.I(new_n12150_), .ZN(new_n12186_));
  INV_X1     g11882(.I(new_n12152_), .ZN(new_n12187_));
  NOR2_X1    g11883(.A1(new_n12187_), .A2(new_n12183_), .ZN(new_n12188_));
  INV_X1     g11884(.I(new_n12188_), .ZN(new_n12189_));
  NAND2_X1   g11885(.A1(new_n12187_), .A2(new_n12183_), .ZN(new_n12190_));
  AOI21_X1   g11886(.A1(new_n12189_), .A2(new_n12190_), .B(new_n12186_), .ZN(new_n12191_));
  NOR2_X1    g11887(.A1(new_n12191_), .A2(new_n12185_), .ZN(new_n12192_));
  XOR2_X1    g11888(.A1(new_n12149_), .A2(new_n12192_), .Z(new_n12193_));
  NOR2_X1    g11889(.A1(new_n12149_), .A2(new_n12192_), .ZN(new_n12194_));
  INV_X1     g11890(.I(new_n12194_), .ZN(new_n12195_));
  NAND2_X1   g11891(.A1(new_n12149_), .A2(new_n12192_), .ZN(new_n12196_));
  AOI21_X1   g11892(.A1(new_n12195_), .A2(new_n12196_), .B(new_n12148_), .ZN(new_n12197_));
  AOI21_X1   g11893(.A1(new_n12148_), .A2(new_n12193_), .B(new_n12197_), .ZN(new_n12198_));
  INV_X1     g11894(.I(new_n11995_), .ZN(new_n12199_));
  OR2_X2     g11895(.A1(new_n11996_), .A2(new_n11947_), .Z(new_n12200_));
  NAND2_X1   g11896(.A1(new_n12200_), .A2(new_n12199_), .ZN(new_n12201_));
  XNOR2_X1   g11897(.A1(new_n12201_), .A2(new_n12198_), .ZN(new_n12202_));
  NAND2_X1   g11898(.A1(new_n12008_), .A2(new_n12202_), .ZN(new_n12203_));
  INV_X1     g11899(.I(new_n12201_), .ZN(new_n12204_));
  NOR2_X1    g11900(.A1(new_n12204_), .A2(new_n12198_), .ZN(new_n12205_));
  NAND2_X1   g11901(.A1(new_n12204_), .A2(new_n12198_), .ZN(new_n12206_));
  INV_X1     g11902(.I(new_n12206_), .ZN(new_n12207_));
  NOR2_X1    g11903(.A1(new_n12207_), .A2(new_n12205_), .ZN(new_n12208_));
  OAI21_X1   g11904(.A1(new_n12008_), .A2(new_n12208_), .B(new_n12203_), .ZN(\asquared[77] ));
  NOR2_X1    g11905(.A1(new_n12205_), .A2(new_n11999_), .ZN(new_n12210_));
  AOI21_X1   g11906(.A1(new_n12205_), .A2(new_n11999_), .B(new_n11796_), .ZN(new_n12211_));
  NOR2_X1    g11907(.A1(new_n12211_), .A2(new_n12210_), .ZN(new_n12212_));
  NAND2_X1   g11908(.A1(new_n11794_), .A2(new_n12212_), .ZN(new_n12213_));
  OAI21_X1   g11909(.A1(new_n12148_), .A2(new_n12194_), .B(new_n12196_), .ZN(new_n12214_));
  INV_X1     g11910(.I(new_n12214_), .ZN(new_n12215_));
  INV_X1     g11911(.I(new_n12010_), .ZN(new_n12216_));
  AOI21_X1   g11912(.A1(new_n12216_), .A2(new_n12145_), .B(new_n12144_), .ZN(new_n12217_));
  INV_X1     g11913(.I(new_n12078_), .ZN(new_n12218_));
  AOI21_X1   g11914(.A1(new_n12084_), .A2(new_n12218_), .B(new_n12081_), .ZN(new_n12219_));
  INV_X1     g11915(.I(new_n12134_), .ZN(new_n12220_));
  AOI21_X1   g11916(.A1(new_n12220_), .A2(new_n12139_), .B(new_n12136_), .ZN(new_n12221_));
  AOI21_X1   g11917(.A1(new_n12031_), .A2(new_n12035_), .B(new_n12033_), .ZN(new_n12222_));
  NAND2_X1   g11918(.A1(new_n12117_), .A2(new_n12115_), .ZN(new_n12223_));
  NAND2_X1   g11919(.A1(new_n12223_), .A2(new_n12114_), .ZN(new_n12224_));
  NOR2_X1    g11920(.A1(new_n10722_), .A2(new_n4048_), .ZN(new_n12225_));
  NOR2_X1    g11921(.A1(new_n1999_), .A2(new_n6692_), .ZN(new_n12226_));
  NAND4_X1   g11922(.A1(new_n12225_), .A2(new_n1956_), .A3(new_n10288_), .A4(new_n12226_), .ZN(new_n12227_));
  NAND2_X1   g11923(.A1(new_n3851_), .A2(new_n5742_), .ZN(new_n12228_));
  NAND2_X1   g11924(.A1(\a[16] ), .A2(\a[61] ), .ZN(new_n12229_));
  XNOR2_X1   g11925(.A1(new_n12228_), .A2(new_n12229_), .ZN(new_n12230_));
  NOR4_X1    g11926(.A1(new_n1916_), .A2(new_n3371_), .A3(new_n4501_), .A4(new_n6260_), .ZN(new_n12231_));
  XOR2_X1    g11927(.A1(new_n12231_), .A2(new_n1674_), .Z(new_n12232_));
  XOR2_X1    g11928(.A1(new_n12232_), .A2(\a[55] ), .Z(new_n12233_));
  NOR2_X1    g11929(.A1(new_n12233_), .A2(new_n12230_), .ZN(new_n12234_));
  AND2_X2    g11930(.A1(new_n12233_), .A2(new_n12230_), .Z(new_n12235_));
  NOR2_X1    g11931(.A1(new_n12235_), .A2(new_n12234_), .ZN(new_n12236_));
  NOR2_X1    g11932(.A1(new_n12236_), .A2(new_n12227_), .ZN(new_n12237_));
  INV_X1     g11933(.I(new_n12227_), .ZN(new_n12238_));
  XNOR2_X1   g11934(.A1(new_n12233_), .A2(new_n12230_), .ZN(new_n12239_));
  NOR2_X1    g11935(.A1(new_n12239_), .A2(new_n12238_), .ZN(new_n12240_));
  NOR2_X1    g11936(.A1(new_n12237_), .A2(new_n12240_), .ZN(new_n12241_));
  XOR2_X1    g11937(.A1(new_n12224_), .A2(new_n12241_), .Z(new_n12242_));
  NOR2_X1    g11938(.A1(new_n12242_), .A2(new_n12222_), .ZN(new_n12243_));
  INV_X1     g11939(.I(new_n12222_), .ZN(new_n12244_));
  INV_X1     g11940(.I(new_n12224_), .ZN(new_n12245_));
  NOR2_X1    g11941(.A1(new_n12245_), .A2(new_n12241_), .ZN(new_n12246_));
  INV_X1     g11942(.I(new_n12246_), .ZN(new_n12247_));
  NAND2_X1   g11943(.A1(new_n12245_), .A2(new_n12241_), .ZN(new_n12248_));
  AOI21_X1   g11944(.A1(new_n12247_), .A2(new_n12248_), .B(new_n12244_), .ZN(new_n12249_));
  NOR2_X1    g11945(.A1(new_n12249_), .A2(new_n12243_), .ZN(new_n12250_));
  XOR2_X1    g11946(.A1(new_n12250_), .A2(new_n12221_), .Z(new_n12251_));
  INV_X1     g11947(.I(new_n12221_), .ZN(new_n12252_));
  NOR2_X1    g11948(.A1(new_n12250_), .A2(new_n12252_), .ZN(new_n12253_));
  NAND2_X1   g11949(.A1(new_n12250_), .A2(new_n12252_), .ZN(new_n12254_));
  INV_X1     g11950(.I(new_n12254_), .ZN(new_n12255_));
  OAI21_X1   g11951(.A1(new_n12255_), .A2(new_n12253_), .B(new_n12219_), .ZN(new_n12256_));
  OAI21_X1   g11952(.A1(new_n12219_), .A2(new_n12251_), .B(new_n12256_), .ZN(new_n12257_));
  OAI21_X1   g11953(.A1(new_n12150_), .A2(new_n12188_), .B(new_n12190_), .ZN(new_n12258_));
  INV_X1     g11954(.I(new_n12258_), .ZN(new_n12259_));
  AOI21_X1   g11955(.A1(new_n12072_), .A2(new_n12075_), .B(new_n12073_), .ZN(new_n12260_));
  INV_X1     g11956(.I(new_n12023_), .ZN(new_n12261_));
  AOI21_X1   g11957(.A1(new_n12019_), .A2(new_n12261_), .B(new_n12022_), .ZN(new_n12262_));
  NOR2_X1    g11958(.A1(new_n12103_), .A2(new_n12101_), .ZN(new_n12263_));
  NOR2_X1    g11959(.A1(new_n12263_), .A2(new_n12102_), .ZN(new_n12264_));
  AOI21_X1   g11960(.A1(new_n2277_), .A2(new_n5601_), .B(new_n6777_), .ZN(new_n12265_));
  NAND2_X1   g11961(.A1(\a[17] ), .A2(\a[59] ), .ZN(new_n12266_));
  NOR2_X1    g11962(.A1(new_n1276_), .A2(new_n8990_), .ZN(new_n12267_));
  XOR2_X1    g11963(.A1(new_n12267_), .A2(new_n12266_), .Z(new_n12268_));
  XOR2_X1    g11964(.A1(new_n12268_), .A2(new_n12265_), .Z(new_n12269_));
  XNOR2_X1   g11965(.A1(new_n12264_), .A2(new_n12269_), .ZN(new_n12270_));
  NOR2_X1    g11966(.A1(new_n12264_), .A2(new_n12269_), .ZN(new_n12271_));
  NAND2_X1   g11967(.A1(new_n12264_), .A2(new_n12269_), .ZN(new_n12272_));
  INV_X1     g11968(.I(new_n12272_), .ZN(new_n12273_));
  OAI21_X1   g11969(.A1(new_n12273_), .A2(new_n12271_), .B(new_n12262_), .ZN(new_n12274_));
  OAI21_X1   g11970(.A1(new_n12270_), .A2(new_n12262_), .B(new_n12274_), .ZN(new_n12275_));
  NAND2_X1   g11971(.A1(new_n3981_), .A2(new_n5742_), .ZN(new_n12276_));
  NOR2_X1    g11972(.A1(new_n3981_), .A2(new_n5742_), .ZN(new_n12277_));
  NOR2_X1    g11973(.A1(\a[13] ), .A2(\a[63] ), .ZN(new_n12278_));
  AOI21_X1   g11974(.A1(new_n12276_), .A2(new_n12278_), .B(new_n12277_), .ZN(new_n12279_));
  INV_X1     g11975(.I(new_n12279_), .ZN(new_n12280_));
  AOI21_X1   g11976(.A1(new_n4538_), .A2(new_n7483_), .B(new_n12161_), .ZN(new_n12281_));
  AOI21_X1   g11977(.A1(new_n2898_), .A2(new_n5980_), .B(new_n12053_), .ZN(new_n12282_));
  INV_X1     g11978(.I(new_n12282_), .ZN(new_n12283_));
  XOR2_X1    g11979(.A1(new_n12281_), .A2(new_n12283_), .Z(new_n12284_));
  AND2_X2    g11980(.A1(new_n12281_), .A2(new_n12282_), .Z(new_n12285_));
  NOR2_X1    g11981(.A1(new_n12281_), .A2(new_n12282_), .ZN(new_n12286_));
  OAI21_X1   g11982(.A1(new_n12285_), .A2(new_n12286_), .B(new_n12280_), .ZN(new_n12287_));
  OAI21_X1   g11983(.A1(new_n12284_), .A2(new_n12280_), .B(new_n12287_), .ZN(new_n12288_));
  AOI21_X1   g11984(.A1(new_n1275_), .A2(new_n8996_), .B(new_n12040_), .ZN(new_n12289_));
  INV_X1     g11985(.I(new_n12289_), .ZN(new_n12290_));
  NAND2_X1   g11986(.A1(new_n2533_), .A2(new_n6280_), .ZN(new_n12291_));
  NOR2_X1    g11987(.A1(new_n2533_), .A2(new_n6280_), .ZN(new_n12292_));
  NOR2_X1    g11988(.A1(\a[18] ), .A2(\a[58] ), .ZN(new_n12293_));
  AOI21_X1   g11989(.A1(new_n12291_), .A2(new_n12293_), .B(new_n12292_), .ZN(new_n12294_));
  NOR2_X1    g11990(.A1(new_n1339_), .A2(new_n7727_), .ZN(new_n12295_));
  OAI21_X1   g11991(.A1(new_n5557_), .A2(new_n12165_), .B(new_n12295_), .ZN(new_n12296_));
  OAI21_X1   g11992(.A1(new_n5563_), .A2(new_n12166_), .B(new_n12296_), .ZN(new_n12297_));
  XNOR2_X1   g11993(.A1(new_n12297_), .A2(new_n12294_), .ZN(new_n12298_));
  AND2_X2    g11994(.A1(new_n12297_), .A2(new_n12294_), .Z(new_n12299_));
  NOR2_X1    g11995(.A1(new_n12297_), .A2(new_n12294_), .ZN(new_n12300_));
  OAI21_X1   g11996(.A1(new_n12299_), .A2(new_n12300_), .B(new_n12290_), .ZN(new_n12301_));
  OAI21_X1   g11997(.A1(new_n12290_), .A2(new_n12298_), .B(new_n12301_), .ZN(new_n12302_));
  NOR2_X1    g11998(.A1(new_n12171_), .A2(new_n12158_), .ZN(new_n12303_));
  NOR2_X1    g11999(.A1(new_n12303_), .A2(new_n12170_), .ZN(new_n12304_));
  NOR2_X1    g12000(.A1(new_n12304_), .A2(new_n12302_), .ZN(new_n12305_));
  NAND2_X1   g12001(.A1(new_n12304_), .A2(new_n12302_), .ZN(new_n12306_));
  INV_X1     g12002(.I(new_n12306_), .ZN(new_n12307_));
  OAI21_X1   g12003(.A1(new_n12307_), .A2(new_n12305_), .B(new_n12288_), .ZN(new_n12308_));
  XNOR2_X1   g12004(.A1(new_n12304_), .A2(new_n12302_), .ZN(new_n12309_));
  OAI21_X1   g12005(.A1(new_n12288_), .A2(new_n12309_), .B(new_n12308_), .ZN(new_n12310_));
  XNOR2_X1   g12006(.A1(new_n12310_), .A2(new_n12275_), .ZN(new_n12311_));
  NOR2_X1    g12007(.A1(new_n12311_), .A2(new_n12260_), .ZN(new_n12312_));
  INV_X1     g12008(.I(new_n12260_), .ZN(new_n12313_));
  NAND2_X1   g12009(.A1(new_n12310_), .A2(new_n12275_), .ZN(new_n12314_));
  NOR2_X1    g12010(.A1(new_n12310_), .A2(new_n12275_), .ZN(new_n12315_));
  INV_X1     g12011(.I(new_n12315_), .ZN(new_n12316_));
  AOI21_X1   g12012(.A1(new_n12316_), .A2(new_n12314_), .B(new_n12313_), .ZN(new_n12317_));
  NOR2_X1    g12013(.A1(new_n12312_), .A2(new_n12317_), .ZN(new_n12318_));
  AOI21_X1   g12014(.A1(new_n12153_), .A2(new_n12181_), .B(new_n12179_), .ZN(new_n12319_));
  AOI21_X1   g12015(.A1(new_n12039_), .A2(new_n12049_), .B(new_n12048_), .ZN(new_n12320_));
  NAND2_X1   g12016(.A1(new_n12066_), .A2(new_n12064_), .ZN(new_n12321_));
  NAND2_X1   g12017(.A1(new_n12321_), .A2(new_n12063_), .ZN(new_n12322_));
  NOR2_X1    g12018(.A1(new_n650_), .A2(new_n9029_), .ZN(new_n12323_));
  OAI21_X1   g12019(.A1(new_n12107_), .A2(new_n12109_), .B(new_n12323_), .ZN(new_n12324_));
  NAND2_X1   g12020(.A1(new_n12324_), .A2(new_n12110_), .ZN(new_n12325_));
  INV_X1     g12021(.I(new_n12325_), .ZN(new_n12326_));
  XOR2_X1    g12022(.A1(new_n12322_), .A2(new_n12326_), .Z(new_n12327_));
  AOI21_X1   g12023(.A1(new_n12063_), .A2(new_n12321_), .B(new_n12326_), .ZN(new_n12328_));
  NOR2_X1    g12024(.A1(new_n12322_), .A2(new_n12325_), .ZN(new_n12329_));
  OAI21_X1   g12025(.A1(new_n12329_), .A2(new_n12328_), .B(new_n12320_), .ZN(new_n12330_));
  OAI21_X1   g12026(.A1(new_n12327_), .A2(new_n12320_), .B(new_n12330_), .ZN(new_n12331_));
  NAND2_X1   g12027(.A1(\a[31] ), .A2(\a[63] ), .ZN(new_n12332_));
  NOR2_X1    g12028(.A1(new_n7139_), .A2(new_n12332_), .ZN(new_n12333_));
  NOR4_X1    g12029(.A1(new_n650_), .A2(new_n2655_), .A3(new_n5175_), .A4(new_n9310_), .ZN(new_n12337_));
  AOI22_X1   g12030(.A1(new_n3966_), .A2(new_n12056_), .B1(new_n5184_), .B2(new_n5350_), .ZN(new_n12338_));
  NOR3_X1    g12031(.A1(new_n3838_), .A2(new_n5592_), .A3(new_n5581_), .ZN(new_n12339_));
  NAND2_X1   g12032(.A1(new_n12338_), .A2(new_n12339_), .ZN(new_n12340_));
  XNOR2_X1   g12033(.A1(new_n6782_), .A2(new_n12108_), .ZN(new_n12341_));
  NOR2_X1    g12034(.A1(new_n12340_), .A2(new_n12341_), .ZN(new_n12342_));
  AND2_X2    g12035(.A1(new_n12340_), .A2(new_n12341_), .Z(new_n12343_));
  NOR2_X1    g12036(.A1(new_n12343_), .A2(new_n12342_), .ZN(new_n12344_));
  XNOR2_X1   g12037(.A1(new_n12340_), .A2(new_n12341_), .ZN(new_n12345_));
  MUX2_X1    g12038(.I0(new_n12345_), .I1(new_n12344_), .S(new_n12337_), .Z(new_n12346_));
  NOR2_X1    g12039(.A1(new_n12130_), .A2(new_n12121_), .ZN(new_n12347_));
  NOR2_X1    g12040(.A1(new_n12347_), .A2(new_n12128_), .ZN(new_n12348_));
  AOI21_X1   g12041(.A1(new_n3966_), .A2(new_n5592_), .B(new_n12057_), .ZN(new_n12349_));
  NOR2_X1    g12042(.A1(new_n8247_), .A2(new_n6638_), .ZN(new_n12350_));
  NOR4_X1    g12043(.A1(new_n8242_), .A2(new_n2978_), .A3(new_n1339_), .A4(new_n7647_), .ZN(new_n12351_));
  NAND2_X1   g12044(.A1(new_n12350_), .A2(new_n12351_), .ZN(new_n12352_));
  AOI22_X1   g12045(.A1(new_n2500_), .A2(new_n6280_), .B1(new_n6056_), .B2(new_n2797_), .ZN(new_n12353_));
  INV_X1     g12046(.I(new_n12353_), .ZN(new_n12354_));
  INV_X1     g12047(.I(new_n6028_), .ZN(new_n12355_));
  NAND4_X1   g12048(.A1(new_n12355_), .A2(\a[27] ), .A3(\a[50] ), .A4(new_n2689_), .ZN(new_n12356_));
  NOR2_X1    g12049(.A1(new_n12354_), .A2(new_n12356_), .ZN(new_n12357_));
  XNOR2_X1   g12050(.A1(new_n12352_), .A2(new_n12357_), .ZN(new_n12358_));
  NAND2_X1   g12051(.A1(new_n12358_), .A2(new_n12349_), .ZN(new_n12359_));
  INV_X1     g12052(.I(new_n12349_), .ZN(new_n12360_));
  INV_X1     g12053(.I(new_n12357_), .ZN(new_n12361_));
  NOR2_X1    g12054(.A1(new_n12361_), .A2(new_n12352_), .ZN(new_n12362_));
  NAND2_X1   g12055(.A1(new_n12361_), .A2(new_n12352_), .ZN(new_n12363_));
  INV_X1     g12056(.I(new_n12363_), .ZN(new_n12364_));
  OAI21_X1   g12057(.A1(new_n12364_), .A2(new_n12362_), .B(new_n12360_), .ZN(new_n12365_));
  NAND2_X1   g12058(.A1(new_n12359_), .A2(new_n12365_), .ZN(new_n12366_));
  INV_X1     g12059(.I(new_n12366_), .ZN(new_n12367_));
  XOR2_X1    g12060(.A1(new_n12348_), .A2(new_n12367_), .Z(new_n12368_));
  NOR3_X1    g12061(.A1(new_n12347_), .A2(new_n12128_), .A3(new_n12367_), .ZN(new_n12369_));
  NOR2_X1    g12062(.A1(new_n12348_), .A2(new_n12366_), .ZN(new_n12370_));
  OAI21_X1   g12063(.A1(new_n12370_), .A2(new_n12369_), .B(new_n12346_), .ZN(new_n12371_));
  OAI21_X1   g12064(.A1(new_n12368_), .A2(new_n12346_), .B(new_n12371_), .ZN(new_n12372_));
  NAND2_X1   g12065(.A1(new_n12372_), .A2(new_n12331_), .ZN(new_n12373_));
  NOR2_X1    g12066(.A1(new_n12372_), .A2(new_n12331_), .ZN(new_n12374_));
  INV_X1     g12067(.I(new_n12374_), .ZN(new_n12375_));
  AOI21_X1   g12068(.A1(new_n12375_), .A2(new_n12373_), .B(new_n12319_), .ZN(new_n12376_));
  INV_X1     g12069(.I(new_n12319_), .ZN(new_n12377_));
  XNOR2_X1   g12070(.A1(new_n12372_), .A2(new_n12331_), .ZN(new_n12378_));
  NOR2_X1    g12071(.A1(new_n12378_), .A2(new_n12377_), .ZN(new_n12379_));
  NOR2_X1    g12072(.A1(new_n12379_), .A2(new_n12376_), .ZN(new_n12380_));
  XOR2_X1    g12073(.A1(new_n12318_), .A2(new_n12380_), .Z(new_n12381_));
  INV_X1     g12074(.I(new_n12318_), .ZN(new_n12382_));
  NOR2_X1    g12075(.A1(new_n12382_), .A2(new_n12380_), .ZN(new_n12383_));
  NAND2_X1   g12076(.A1(new_n12382_), .A2(new_n12380_), .ZN(new_n12384_));
  INV_X1     g12077(.I(new_n12384_), .ZN(new_n12385_));
  OAI21_X1   g12078(.A1(new_n12385_), .A2(new_n12383_), .B(new_n12259_), .ZN(new_n12386_));
  OAI21_X1   g12079(.A1(new_n12259_), .A2(new_n12381_), .B(new_n12386_), .ZN(new_n12387_));
  NAND2_X1   g12080(.A1(new_n12387_), .A2(new_n12257_), .ZN(new_n12388_));
  NOR2_X1    g12081(.A1(new_n12387_), .A2(new_n12257_), .ZN(new_n12389_));
  INV_X1     g12082(.I(new_n12389_), .ZN(new_n12390_));
  AOI21_X1   g12083(.A1(new_n12390_), .A2(new_n12388_), .B(new_n12217_), .ZN(new_n12391_));
  INV_X1     g12084(.I(new_n12217_), .ZN(new_n12392_));
  XNOR2_X1   g12085(.A1(new_n12387_), .A2(new_n12257_), .ZN(new_n12393_));
  NOR2_X1    g12086(.A1(new_n12393_), .A2(new_n12392_), .ZN(new_n12394_));
  NOR2_X1    g12087(.A1(new_n12394_), .A2(new_n12391_), .ZN(new_n12395_));
  NOR2_X1    g12088(.A1(new_n12395_), .A2(new_n12215_), .ZN(new_n12396_));
  XOR2_X1    g12089(.A1(new_n12213_), .A2(new_n12396_), .Z(new_n12397_));
  XOR2_X1    g12090(.A1(new_n12397_), .A2(new_n12206_), .Z(\asquared[78] ));
  NOR2_X1    g12091(.A1(new_n12206_), .A2(new_n12215_), .ZN(new_n12399_));
  INV_X1     g12092(.I(new_n12399_), .ZN(new_n12400_));
  AOI21_X1   g12093(.A1(new_n12206_), .A2(new_n12215_), .B(new_n12395_), .ZN(new_n12401_));
  NAND3_X1   g12094(.A1(new_n11794_), .A2(new_n12212_), .A3(new_n12401_), .ZN(new_n12402_));
  NAND2_X1   g12095(.A1(new_n12402_), .A2(new_n12400_), .ZN(new_n12403_));
  INV_X1     g12096(.I(new_n12403_), .ZN(new_n12404_));
  NAND2_X1   g12097(.A1(new_n12388_), .A2(new_n12392_), .ZN(new_n12405_));
  NAND2_X1   g12098(.A1(new_n12405_), .A2(new_n12390_), .ZN(new_n12406_));
  OAI21_X1   g12099(.A1(new_n12219_), .A2(new_n12253_), .B(new_n12254_), .ZN(new_n12407_));
  INV_X1     g12100(.I(new_n12407_), .ZN(new_n12408_));
  AOI21_X1   g12101(.A1(new_n12244_), .A2(new_n12248_), .B(new_n12246_), .ZN(new_n12409_));
  NOR2_X1    g12102(.A1(new_n12273_), .A2(new_n12262_), .ZN(new_n12410_));
  NOR2_X1    g12103(.A1(new_n12410_), .A2(new_n12271_), .ZN(new_n12411_));
  NOR2_X1    g12104(.A1(new_n12286_), .A2(new_n12280_), .ZN(new_n12412_));
  NOR2_X1    g12105(.A1(new_n12412_), .A2(new_n12285_), .ZN(new_n12413_));
  INV_X1     g12106(.I(new_n12413_), .ZN(new_n12414_));
  NAND2_X1   g12107(.A1(new_n3966_), .A2(new_n5173_), .ZN(new_n12415_));
  NOR2_X1    g12108(.A1(new_n2368_), .A2(new_n6999_), .ZN(new_n12416_));
  XOR2_X1    g12109(.A1(new_n12415_), .A2(new_n12416_), .Z(new_n12417_));
  NOR2_X1    g12110(.A1(new_n1916_), .A2(new_n6692_), .ZN(new_n12418_));
  NAND4_X1   g12111(.A1(\a[37] ), .A2(\a[38] ), .A3(\a[40] ), .A4(\a[41] ), .ZN(new_n12419_));
  XOR2_X1    g12112(.A1(new_n12417_), .A2(new_n12419_), .Z(new_n12420_));
  NAND2_X1   g12113(.A1(new_n12414_), .A2(new_n12420_), .ZN(new_n12421_));
  NOR2_X1    g12114(.A1(new_n12417_), .A2(new_n12419_), .ZN(new_n12422_));
  NAND2_X1   g12115(.A1(new_n12417_), .A2(new_n12419_), .ZN(new_n12423_));
  INV_X1     g12116(.I(new_n12423_), .ZN(new_n12424_));
  OAI21_X1   g12117(.A1(new_n12422_), .A2(new_n12424_), .B(new_n12413_), .ZN(new_n12425_));
  NAND2_X1   g12118(.A1(new_n12421_), .A2(new_n12425_), .ZN(new_n12426_));
  AOI21_X1   g12119(.A1(new_n2978_), .A2(new_n8242_), .B(new_n12350_), .ZN(new_n12427_));
  OAI22_X1   g12120(.A1(new_n12268_), .A2(new_n9553_), .B1(new_n1268_), .B2(new_n12265_), .ZN(new_n12428_));
  AOI22_X1   g12121(.A1(\a[26] ), .A2(\a[51] ), .B1(\a[34] ), .B2(\a[43] ), .ZN(new_n12429_));
  NOR3_X1    g12122(.A1(new_n12429_), .A2(new_n1674_), .A3(new_n6999_), .ZN(new_n12430_));
  NOR2_X1    g12123(.A1(new_n12430_), .A2(new_n12231_), .ZN(new_n12431_));
  XOR2_X1    g12124(.A1(new_n12428_), .A2(new_n12431_), .Z(new_n12432_));
  INV_X1     g12125(.I(new_n12432_), .ZN(new_n12433_));
  INV_X1     g12126(.I(new_n12428_), .ZN(new_n12434_));
  NOR2_X1    g12127(.A1(new_n12434_), .A2(new_n12431_), .ZN(new_n12435_));
  INV_X1     g12128(.I(new_n12435_), .ZN(new_n12436_));
  NAND2_X1   g12129(.A1(new_n12434_), .A2(new_n12431_), .ZN(new_n12437_));
  AOI21_X1   g12130(.A1(new_n12436_), .A2(new_n12437_), .B(new_n12427_), .ZN(new_n12438_));
  AOI21_X1   g12131(.A1(new_n12427_), .A2(new_n12433_), .B(new_n12438_), .ZN(new_n12439_));
  XOR2_X1    g12132(.A1(new_n12426_), .A2(new_n12439_), .Z(new_n12440_));
  NOR2_X1    g12133(.A1(new_n12440_), .A2(new_n12411_), .ZN(new_n12441_));
  INV_X1     g12134(.I(new_n12411_), .ZN(new_n12442_));
  INV_X1     g12135(.I(new_n12426_), .ZN(new_n12443_));
  NOR2_X1    g12136(.A1(new_n12443_), .A2(new_n12439_), .ZN(new_n12444_));
  INV_X1     g12137(.I(new_n12444_), .ZN(new_n12445_));
  NAND2_X1   g12138(.A1(new_n12443_), .A2(new_n12439_), .ZN(new_n12446_));
  AOI21_X1   g12139(.A1(new_n12445_), .A2(new_n12446_), .B(new_n12442_), .ZN(new_n12447_));
  NOR2_X1    g12140(.A1(new_n12447_), .A2(new_n12441_), .ZN(new_n12448_));
  INV_X1     g12141(.I(new_n12448_), .ZN(new_n12449_));
  INV_X1     g12142(.I(new_n12370_), .ZN(new_n12450_));
  OR2_X2     g12143(.A1(new_n12369_), .A2(new_n12346_), .Z(new_n12451_));
  NAND2_X1   g12144(.A1(new_n12451_), .A2(new_n12450_), .ZN(new_n12452_));
  INV_X1     g12145(.I(new_n12452_), .ZN(new_n12453_));
  NOR2_X1    g12146(.A1(new_n12449_), .A2(new_n12453_), .ZN(new_n12454_));
  NOR2_X1    g12147(.A1(new_n12448_), .A2(new_n12452_), .ZN(new_n12455_));
  NOR2_X1    g12148(.A1(new_n12454_), .A2(new_n12455_), .ZN(new_n12456_));
  NOR2_X1    g12149(.A1(new_n12456_), .A2(new_n12409_), .ZN(new_n12457_));
  INV_X1     g12150(.I(new_n12409_), .ZN(new_n12458_));
  XOR2_X1    g12151(.A1(new_n12448_), .A2(new_n12453_), .Z(new_n12459_));
  NOR2_X1    g12152(.A1(new_n12458_), .A2(new_n12459_), .ZN(new_n12460_));
  NOR2_X1    g12153(.A1(new_n12457_), .A2(new_n12460_), .ZN(new_n12461_));
  INV_X1     g12154(.I(new_n12343_), .ZN(new_n12462_));
  AOI21_X1   g12155(.A1(new_n12462_), .A2(new_n12337_), .B(new_n12342_), .ZN(new_n12463_));
  AOI21_X1   g12156(.A1(new_n12349_), .A2(new_n12363_), .B(new_n12362_), .ZN(new_n12464_));
  NOR2_X1    g12157(.A1(new_n12235_), .A2(new_n12227_), .ZN(new_n12465_));
  NOR2_X1    g12158(.A1(new_n12465_), .A2(new_n12234_), .ZN(new_n12466_));
  XNOR2_X1   g12159(.A1(new_n12466_), .A2(new_n12464_), .ZN(new_n12467_));
  NOR2_X1    g12160(.A1(new_n12467_), .A2(new_n12463_), .ZN(new_n12468_));
  INV_X1     g12161(.I(new_n12463_), .ZN(new_n12469_));
  NOR2_X1    g12162(.A1(new_n12466_), .A2(new_n12464_), .ZN(new_n12470_));
  INV_X1     g12163(.I(new_n12470_), .ZN(new_n12471_));
  NAND2_X1   g12164(.A1(new_n12466_), .A2(new_n12464_), .ZN(new_n12472_));
  AOI21_X1   g12165(.A1(new_n12471_), .A2(new_n12472_), .B(new_n12469_), .ZN(new_n12473_));
  NOR2_X1    g12166(.A1(new_n12468_), .A2(new_n12473_), .ZN(new_n12474_));
  AOI21_X1   g12167(.A1(new_n3126_), .A2(new_n5980_), .B(new_n12333_), .ZN(new_n12475_));
  INV_X1     g12168(.I(new_n12475_), .ZN(new_n12476_));
  NAND2_X1   g12169(.A1(new_n3851_), .A2(new_n5742_), .ZN(new_n12477_));
  NOR2_X1    g12170(.A1(new_n3851_), .A2(new_n5742_), .ZN(new_n12478_));
  NOR2_X1    g12171(.A1(\a[16] ), .A2(\a[61] ), .ZN(new_n12479_));
  AOI21_X1   g12172(.A1(new_n12477_), .A2(new_n12479_), .B(new_n12478_), .ZN(new_n12480_));
  AOI21_X1   g12173(.A1(new_n2690_), .A2(new_n6028_), .B(new_n12353_), .ZN(new_n12481_));
  XNOR2_X1   g12174(.A1(new_n12481_), .A2(new_n12480_), .ZN(new_n12482_));
  NOR2_X1    g12175(.A1(new_n12482_), .A2(new_n12476_), .ZN(new_n12483_));
  INV_X1     g12176(.I(new_n12480_), .ZN(new_n12484_));
  INV_X1     g12177(.I(new_n12481_), .ZN(new_n12485_));
  NOR2_X1    g12178(.A1(new_n12485_), .A2(new_n12484_), .ZN(new_n12486_));
  NOR2_X1    g12179(.A1(new_n12481_), .A2(new_n12480_), .ZN(new_n12487_));
  NOR2_X1    g12180(.A1(new_n12486_), .A2(new_n12487_), .ZN(new_n12488_));
  NOR2_X1    g12181(.A1(new_n12488_), .A2(new_n12475_), .ZN(new_n12489_));
  NOR2_X1    g12182(.A1(new_n12489_), .A2(new_n12483_), .ZN(new_n12490_));
  AOI21_X1   g12183(.A1(new_n2543_), .A2(new_n7482_), .B(new_n12225_), .ZN(new_n12491_));
  INV_X1     g12184(.I(new_n12491_), .ZN(new_n12492_));
  AOI21_X1   g12185(.A1(new_n3838_), .A2(new_n5592_), .B(new_n12338_), .ZN(new_n12493_));
  AOI21_X1   g12186(.A1(\a[62] ), .A2(new_n6782_), .B(new_n5339_), .ZN(new_n12494_));
  INV_X1     g12187(.I(new_n12494_), .ZN(new_n12495_));
  XOR2_X1    g12188(.A1(new_n12493_), .A2(new_n12495_), .Z(new_n12496_));
  NOR2_X1    g12189(.A1(new_n12496_), .A2(new_n12492_), .ZN(new_n12497_));
  INV_X1     g12190(.I(new_n12493_), .ZN(new_n12498_));
  NOR2_X1    g12191(.A1(new_n12498_), .A2(new_n12495_), .ZN(new_n12499_));
  NOR2_X1    g12192(.A1(new_n12493_), .A2(new_n12494_), .ZN(new_n12500_));
  NOR2_X1    g12193(.A1(new_n12499_), .A2(new_n12500_), .ZN(new_n12501_));
  NOR2_X1    g12194(.A1(new_n12501_), .A2(new_n12491_), .ZN(new_n12502_));
  NOR2_X1    g12195(.A1(new_n12502_), .A2(new_n12497_), .ZN(new_n12503_));
  INV_X1     g12196(.I(new_n12503_), .ZN(new_n12504_));
  NOR2_X1    g12197(.A1(new_n12290_), .A2(new_n12300_), .ZN(new_n12505_));
  NOR2_X1    g12198(.A1(new_n12505_), .A2(new_n12299_), .ZN(new_n12506_));
  NOR2_X1    g12199(.A1(new_n12504_), .A2(new_n12506_), .ZN(new_n12507_));
  NOR3_X1    g12200(.A1(new_n12503_), .A2(new_n12299_), .A3(new_n12505_), .ZN(new_n12508_));
  NOR2_X1    g12201(.A1(new_n12507_), .A2(new_n12508_), .ZN(new_n12509_));
  NOR2_X1    g12202(.A1(new_n12509_), .A2(new_n12490_), .ZN(new_n12510_));
  XOR2_X1    g12203(.A1(new_n12503_), .A2(new_n12506_), .Z(new_n12511_));
  NOR3_X1    g12204(.A1(new_n12511_), .A2(new_n12483_), .A3(new_n12489_), .ZN(new_n12512_));
  NOR2_X1    g12205(.A1(new_n12510_), .A2(new_n12512_), .ZN(new_n12513_));
  INV_X1     g12206(.I(new_n12513_), .ZN(new_n12514_));
  NOR2_X1    g12207(.A1(new_n12307_), .A2(new_n12288_), .ZN(new_n12515_));
  NOR2_X1    g12208(.A1(new_n12515_), .A2(new_n12305_), .ZN(new_n12516_));
  NOR2_X1    g12209(.A1(new_n12516_), .A2(new_n12514_), .ZN(new_n12517_));
  INV_X1     g12210(.I(new_n12517_), .ZN(new_n12518_));
  NAND2_X1   g12211(.A1(new_n12516_), .A2(new_n12514_), .ZN(new_n12519_));
  AOI21_X1   g12212(.A1(new_n12518_), .A2(new_n12519_), .B(new_n12474_), .ZN(new_n12520_));
  XOR2_X1    g12213(.A1(new_n12516_), .A2(new_n12513_), .Z(new_n12521_));
  INV_X1     g12214(.I(new_n12521_), .ZN(new_n12522_));
  AOI21_X1   g12215(.A1(new_n12522_), .A2(new_n12474_), .B(new_n12520_), .ZN(new_n12523_));
  XOR2_X1    g12216(.A1(new_n12461_), .A2(new_n12523_), .Z(new_n12524_));
  NOR2_X1    g12217(.A1(new_n12524_), .A2(new_n12408_), .ZN(new_n12525_));
  INV_X1     g12218(.I(new_n12461_), .ZN(new_n12526_));
  NOR2_X1    g12219(.A1(new_n12526_), .A2(new_n12523_), .ZN(new_n12527_));
  INV_X1     g12220(.I(new_n12527_), .ZN(new_n12528_));
  NAND2_X1   g12221(.A1(new_n12526_), .A2(new_n12523_), .ZN(new_n12529_));
  AOI21_X1   g12222(.A1(new_n12528_), .A2(new_n12529_), .B(new_n12407_), .ZN(new_n12530_));
  NOR2_X1    g12223(.A1(new_n12530_), .A2(new_n12525_), .ZN(new_n12531_));
  NOR2_X1    g12224(.A1(new_n12385_), .A2(new_n12259_), .ZN(new_n12532_));
  NOR2_X1    g12225(.A1(new_n12532_), .A2(new_n12383_), .ZN(new_n12533_));
  AOI21_X1   g12226(.A1(new_n12377_), .A2(new_n12373_), .B(new_n12374_), .ZN(new_n12534_));
  NAND2_X1   g12227(.A1(new_n12314_), .A2(new_n12313_), .ZN(new_n12535_));
  NAND2_X1   g12228(.A1(new_n12535_), .A2(new_n12316_), .ZN(new_n12536_));
  NOR2_X1    g12229(.A1(new_n12329_), .A2(new_n12320_), .ZN(new_n12537_));
  NOR2_X1    g12230(.A1(new_n12537_), .A2(new_n12328_), .ZN(new_n12538_));
  NOR2_X1    g12231(.A1(new_n8675_), .A2(new_n1710_), .ZN(new_n12539_));
  NAND2_X1   g12232(.A1(\a[57] ), .A2(\a[60] ), .ZN(new_n12540_));
  NOR2_X1    g12233(.A1(new_n3889_), .A2(new_n12540_), .ZN(new_n12541_));
  NAND2_X1   g12234(.A1(new_n12539_), .A2(new_n12541_), .ZN(new_n12542_));
  AOI21_X1   g12235(.A1(new_n12542_), .A2(new_n9553_), .B(new_n1342_), .ZN(new_n12543_));
  NOR2_X1    g12236(.A1(new_n8675_), .A2(new_n1710_), .ZN(new_n12544_));
  NOR2_X1    g12237(.A1(new_n8941_), .A2(new_n10785_), .ZN(new_n12545_));
  NOR2_X1    g12238(.A1(new_n12545_), .A2(new_n9042_), .ZN(new_n12546_));
  NOR4_X1    g12239(.A1(new_n6280_), .A2(new_n2690_), .A3(new_n2098_), .A4(new_n6260_), .ZN(new_n12547_));
  NAND2_X1   g12240(.A1(new_n12546_), .A2(new_n12547_), .ZN(new_n12548_));
  AOI22_X1   g12241(.A1(new_n1719_), .A2(new_n9781_), .B1(new_n9549_), .B2(new_n1143_), .ZN(new_n12549_));
  NOR4_X1    g12242(.A1(new_n9784_), .A2(new_n1275_), .A3(new_n875_), .A4(new_n9310_), .ZN(new_n12550_));
  NAND2_X1   g12243(.A1(new_n12549_), .A2(new_n12550_), .ZN(new_n12551_));
  NOR2_X1    g12244(.A1(new_n12548_), .A2(new_n12551_), .ZN(new_n12552_));
  INV_X1     g12245(.I(new_n12548_), .ZN(new_n12553_));
  INV_X1     g12246(.I(new_n12551_), .ZN(new_n12554_));
  NOR2_X1    g12247(.A1(new_n12553_), .A2(new_n12554_), .ZN(new_n12555_));
  OAI21_X1   g12248(.A1(new_n12555_), .A2(new_n12552_), .B(new_n12544_), .ZN(new_n12556_));
  XOR2_X1    g12249(.A1(new_n12548_), .A2(new_n12554_), .Z(new_n12557_));
  OAI21_X1   g12250(.A1(new_n12544_), .A2(new_n12557_), .B(new_n12556_), .ZN(new_n12558_));
  NAND2_X1   g12251(.A1(\a[53] ), .A2(\a[54] ), .ZN(new_n12559_));
  NOR2_X1    g12252(.A1(new_n2276_), .A2(new_n12559_), .ZN(new_n12560_));
  NOR2_X1    g12253(.A1(new_n7422_), .A2(new_n2384_), .ZN(new_n12562_));
  NAND2_X1   g12254(.A1(new_n3126_), .A2(new_n6030_), .ZN(new_n12563_));
  NOR2_X1    g12255(.A1(new_n1215_), .A2(new_n7647_), .ZN(new_n12564_));
  XOR2_X1    g12256(.A1(new_n12563_), .A2(new_n12564_), .Z(new_n12565_));
  AOI22_X1   g12257(.A1(new_n3851_), .A2(new_n7452_), .B1(new_n4368_), .B2(new_n5488_), .ZN(new_n12566_));
  NAND4_X1   g12258(.A1(new_n12566_), .A2(new_n4644_), .A3(new_n5487_), .A4(new_n5743_), .ZN(new_n12567_));
  NOR2_X1    g12259(.A1(new_n12565_), .A2(new_n12567_), .ZN(new_n12568_));
  NAND2_X1   g12260(.A1(new_n12565_), .A2(new_n12567_), .ZN(new_n12569_));
  INV_X1     g12261(.I(new_n12569_), .ZN(new_n12570_));
  OAI21_X1   g12262(.A1(new_n12570_), .A2(new_n12568_), .B(new_n12562_), .ZN(new_n12571_));
  XNOR2_X1   g12263(.A1(new_n12565_), .A2(new_n12567_), .ZN(new_n12572_));
  OAI21_X1   g12264(.A1(new_n12562_), .A2(new_n12572_), .B(new_n12571_), .ZN(new_n12573_));
  XNOR2_X1   g12265(.A1(new_n12558_), .A2(new_n12573_), .ZN(new_n12574_));
  NOR2_X1    g12266(.A1(new_n12574_), .A2(new_n12538_), .ZN(new_n12575_));
  INV_X1     g12267(.I(new_n12538_), .ZN(new_n12576_));
  NAND2_X1   g12268(.A1(new_n12558_), .A2(new_n12573_), .ZN(new_n12577_));
  NOR2_X1    g12269(.A1(new_n12558_), .A2(new_n12573_), .ZN(new_n12578_));
  INV_X1     g12270(.I(new_n12578_), .ZN(new_n12579_));
  AOI21_X1   g12271(.A1(new_n12579_), .A2(new_n12577_), .B(new_n12576_), .ZN(new_n12580_));
  NOR2_X1    g12272(.A1(new_n12575_), .A2(new_n12580_), .ZN(new_n12581_));
  XNOR2_X1   g12273(.A1(new_n12536_), .A2(new_n12581_), .ZN(new_n12582_));
  NOR2_X1    g12274(.A1(new_n12536_), .A2(new_n12581_), .ZN(new_n12583_));
  NAND2_X1   g12275(.A1(new_n12536_), .A2(new_n12581_), .ZN(new_n12584_));
  INV_X1     g12276(.I(new_n12584_), .ZN(new_n12585_));
  NOR2_X1    g12277(.A1(new_n12585_), .A2(new_n12583_), .ZN(new_n12586_));
  MUX2_X1    g12278(.I0(new_n12582_), .I1(new_n12586_), .S(new_n12534_), .Z(new_n12587_));
  XOR2_X1    g12279(.A1(new_n12533_), .A2(new_n12587_), .Z(new_n12588_));
  NOR2_X1    g12280(.A1(new_n12588_), .A2(new_n12531_), .ZN(new_n12589_));
  INV_X1     g12281(.I(new_n12531_), .ZN(new_n12590_));
  INV_X1     g12282(.I(new_n12533_), .ZN(new_n12591_));
  NOR2_X1    g12283(.A1(new_n12591_), .A2(new_n12587_), .ZN(new_n12592_));
  INV_X1     g12284(.I(new_n12592_), .ZN(new_n12593_));
  NAND2_X1   g12285(.A1(new_n12591_), .A2(new_n12587_), .ZN(new_n12594_));
  AOI21_X1   g12286(.A1(new_n12593_), .A2(new_n12594_), .B(new_n12590_), .ZN(new_n12595_));
  NOR2_X1    g12287(.A1(new_n12595_), .A2(new_n12589_), .ZN(new_n12596_));
  XOR2_X1    g12288(.A1(new_n12596_), .A2(new_n12406_), .Z(new_n12597_));
  INV_X1     g12289(.I(new_n12596_), .ZN(new_n12598_));
  NAND2_X1   g12290(.A1(new_n12598_), .A2(new_n12406_), .ZN(new_n12599_));
  NAND3_X1   g12291(.A1(new_n12596_), .A2(new_n12390_), .A3(new_n12405_), .ZN(new_n12600_));
  NAND2_X1   g12292(.A1(new_n12599_), .A2(new_n12600_), .ZN(new_n12601_));
  NAND2_X1   g12293(.A1(new_n12404_), .A2(new_n12601_), .ZN(new_n12602_));
  OAI21_X1   g12294(.A1(new_n12404_), .A2(new_n12597_), .B(new_n12602_), .ZN(\asquared[79] ));
  NAND2_X1   g12295(.A1(new_n12403_), .A2(new_n12600_), .ZN(new_n12604_));
  NAND2_X1   g12296(.A1(new_n12604_), .A2(new_n12599_), .ZN(new_n12605_));
  OAI21_X1   g12297(.A1(new_n12590_), .A2(new_n12592_), .B(new_n12594_), .ZN(new_n12606_));
  OAI21_X1   g12298(.A1(new_n12408_), .A2(new_n12527_), .B(new_n12529_), .ZN(new_n12607_));
  NOR2_X1    g12299(.A1(new_n12409_), .A2(new_n12455_), .ZN(new_n12608_));
  NOR2_X1    g12300(.A1(new_n12608_), .A2(new_n12454_), .ZN(new_n12609_));
  OAI21_X1   g12301(.A1(new_n12534_), .A2(new_n12583_), .B(new_n12584_), .ZN(new_n12610_));
  OAI21_X1   g12302(.A1(new_n12538_), .A2(new_n12578_), .B(new_n12577_), .ZN(new_n12611_));
  INV_X1     g12303(.I(new_n12611_), .ZN(new_n12612_));
  NOR2_X1    g12304(.A1(new_n12543_), .A2(new_n12539_), .ZN(new_n12613_));
  INV_X1     g12305(.I(new_n12613_), .ZN(new_n12614_));
  AOI21_X1   g12306(.A1(new_n2383_), .A2(new_n7421_), .B(new_n12560_), .ZN(new_n12615_));
  INV_X1     g12307(.I(new_n12615_), .ZN(new_n12616_));
  AOI21_X1   g12308(.A1(new_n2690_), .A2(new_n6280_), .B(new_n12546_), .ZN(new_n12617_));
  XOR2_X1    g12309(.A1(new_n12617_), .A2(new_n12616_), .Z(new_n12618_));
  AND2_X2    g12310(.A1(new_n12617_), .A2(new_n12615_), .Z(new_n12619_));
  NOR2_X1    g12311(.A1(new_n12617_), .A2(new_n12615_), .ZN(new_n12620_));
  OAI21_X1   g12312(.A1(new_n12619_), .A2(new_n12620_), .B(new_n12614_), .ZN(new_n12621_));
  OAI21_X1   g12313(.A1(new_n12618_), .A2(new_n12614_), .B(new_n12621_), .ZN(new_n12622_));
  INV_X1     g12314(.I(new_n12622_), .ZN(new_n12623_));
  AOI21_X1   g12315(.A1(new_n12414_), .A2(new_n12423_), .B(new_n12422_), .ZN(new_n12624_));
  INV_X1     g12316(.I(new_n12624_), .ZN(new_n12625_));
  NAND2_X1   g12317(.A1(new_n12437_), .A2(new_n12427_), .ZN(new_n12626_));
  NAND2_X1   g12318(.A1(new_n12626_), .A2(new_n12436_), .ZN(new_n12627_));
  NAND2_X1   g12319(.A1(new_n3487_), .A2(new_n5742_), .ZN(new_n12628_));
  NOR2_X1    g12320(.A1(new_n800_), .A2(new_n9310_), .ZN(new_n12629_));
  XOR2_X1    g12321(.A1(new_n12628_), .A2(new_n12629_), .Z(new_n12630_));
  NOR2_X1    g12322(.A1(new_n2098_), .A2(new_n7216_), .ZN(new_n12631_));
  INV_X1     g12323(.I(new_n12631_), .ZN(new_n12632_));
  AOI22_X1   g12324(.A1(\a[23] ), .A2(\a[27] ), .B1(\a[52] ), .B2(\a[56] ), .ZN(new_n12633_));
  NOR3_X1    g12325(.A1(new_n12106_), .A2(new_n12632_), .A3(new_n12633_), .ZN(new_n12634_));
  XOR2_X1    g12326(.A1(new_n12634_), .A2(new_n5877_), .Z(new_n12635_));
  XOR2_X1    g12327(.A1(new_n12635_), .A2(new_n12630_), .Z(new_n12636_));
  NAND2_X1   g12328(.A1(new_n12627_), .A2(new_n12636_), .ZN(new_n12637_));
  INV_X1     g12329(.I(new_n12627_), .ZN(new_n12638_));
  NOR2_X1    g12330(.A1(new_n12635_), .A2(new_n12630_), .ZN(new_n12639_));
  NAND2_X1   g12331(.A1(new_n12635_), .A2(new_n12630_), .ZN(new_n12640_));
  INV_X1     g12332(.I(new_n12640_), .ZN(new_n12641_));
  OAI21_X1   g12333(.A1(new_n12639_), .A2(new_n12641_), .B(new_n12638_), .ZN(new_n12642_));
  AOI21_X1   g12334(.A1(new_n12637_), .A2(new_n12642_), .B(new_n12625_), .ZN(new_n12643_));
  NAND2_X1   g12335(.A1(new_n12642_), .A2(new_n12637_), .ZN(new_n12644_));
  NOR2_X1    g12336(.A1(new_n12644_), .A2(new_n12624_), .ZN(new_n12645_));
  NOR2_X1    g12337(.A1(new_n12645_), .A2(new_n12643_), .ZN(new_n12646_));
  NOR2_X1    g12338(.A1(new_n12646_), .A2(new_n12623_), .ZN(new_n12647_));
  XOR2_X1    g12339(.A1(new_n12644_), .A2(new_n12625_), .Z(new_n12648_));
  NOR2_X1    g12340(.A1(new_n12648_), .A2(new_n12622_), .ZN(new_n12649_));
  NOR2_X1    g12341(.A1(new_n12649_), .A2(new_n12647_), .ZN(new_n12650_));
  AOI21_X1   g12342(.A1(new_n12562_), .A2(new_n12569_), .B(new_n12568_), .ZN(new_n12651_));
  INV_X1     g12343(.I(new_n12651_), .ZN(new_n12652_));
  NAND2_X1   g12344(.A1(new_n2368_), .A2(new_n6999_), .ZN(new_n12653_));
  AOI21_X1   g12345(.A1(new_n3966_), .A2(new_n5173_), .B(new_n12653_), .ZN(new_n12654_));
  AOI21_X1   g12346(.A1(new_n3967_), .A2(new_n5174_), .B(new_n12654_), .ZN(new_n12655_));
  NOR4_X1    g12347(.A1(new_n3837_), .A2(new_n3804_), .A3(new_n4240_), .A4(new_n4414_), .ZN(new_n12656_));
  NAND2_X1   g12348(.A1(new_n12655_), .A2(new_n12656_), .ZN(new_n12657_));
  XOR2_X1    g12349(.A1(new_n12657_), .A2(\a[18] ), .Z(new_n12658_));
  XOR2_X1    g12350(.A1(new_n12658_), .A2(\a[61] ), .Z(new_n12659_));
  AOI21_X1   g12351(.A1(new_n1275_), .A2(new_n9784_), .B(new_n12549_), .ZN(new_n12660_));
  INV_X1     g12352(.I(new_n12660_), .ZN(new_n12661_));
  NAND2_X1   g12353(.A1(new_n3126_), .A2(new_n6030_), .ZN(new_n12662_));
  NOR2_X1    g12354(.A1(new_n3126_), .A2(new_n6030_), .ZN(new_n12663_));
  NOR2_X1    g12355(.A1(\a[20] ), .A2(\a[58] ), .ZN(new_n12664_));
  AOI21_X1   g12356(.A1(new_n12662_), .A2(new_n12664_), .B(new_n12663_), .ZN(new_n12665_));
  AOI21_X1   g12357(.A1(new_n4372_), .A2(new_n5742_), .B(new_n12566_), .ZN(new_n12666_));
  XNOR2_X1   g12358(.A1(new_n12666_), .A2(new_n12665_), .ZN(new_n12667_));
  AND2_X2    g12359(.A1(new_n12666_), .A2(new_n12665_), .Z(new_n12668_));
  NOR2_X1    g12360(.A1(new_n12666_), .A2(new_n12665_), .ZN(new_n12669_));
  OAI21_X1   g12361(.A1(new_n12668_), .A2(new_n12669_), .B(new_n12661_), .ZN(new_n12670_));
  OAI21_X1   g12362(.A1(new_n12661_), .A2(new_n12667_), .B(new_n12670_), .ZN(new_n12671_));
  INV_X1     g12363(.I(new_n12671_), .ZN(new_n12672_));
  XOR2_X1    g12364(.A1(new_n12659_), .A2(new_n12672_), .Z(new_n12673_));
  NAND2_X1   g12365(.A1(new_n12673_), .A2(new_n12652_), .ZN(new_n12674_));
  NOR2_X1    g12366(.A1(new_n12659_), .A2(new_n12672_), .ZN(new_n12675_));
  NAND2_X1   g12367(.A1(new_n12659_), .A2(new_n12672_), .ZN(new_n12676_));
  INV_X1     g12368(.I(new_n12676_), .ZN(new_n12677_));
  OAI21_X1   g12369(.A1(new_n12677_), .A2(new_n12675_), .B(new_n12651_), .ZN(new_n12678_));
  NAND2_X1   g12370(.A1(new_n12674_), .A2(new_n12678_), .ZN(new_n12679_));
  XOR2_X1    g12371(.A1(new_n12650_), .A2(new_n12679_), .Z(new_n12680_));
  INV_X1     g12372(.I(new_n12679_), .ZN(new_n12681_));
  NOR2_X1    g12373(.A1(new_n12650_), .A2(new_n12681_), .ZN(new_n12682_));
  NAND2_X1   g12374(.A1(new_n12650_), .A2(new_n12681_), .ZN(new_n12683_));
  INV_X1     g12375(.I(new_n12683_), .ZN(new_n12684_));
  OAI21_X1   g12376(.A1(new_n12684_), .A2(new_n12682_), .B(new_n12612_), .ZN(new_n12685_));
  OAI21_X1   g12377(.A1(new_n12612_), .A2(new_n12680_), .B(new_n12685_), .ZN(new_n12686_));
  XOR2_X1    g12378(.A1(new_n12610_), .A2(new_n12686_), .Z(new_n12687_));
  NOR2_X1    g12379(.A1(new_n12687_), .A2(new_n12609_), .ZN(new_n12688_));
  INV_X1     g12380(.I(new_n12686_), .ZN(new_n12689_));
  NOR2_X1    g12381(.A1(new_n12689_), .A2(new_n12610_), .ZN(new_n12690_));
  INV_X1     g12382(.I(new_n12690_), .ZN(new_n12691_));
  NAND2_X1   g12383(.A1(new_n12689_), .A2(new_n12610_), .ZN(new_n12692_));
  NAND2_X1   g12384(.A1(new_n12691_), .A2(new_n12692_), .ZN(new_n12693_));
  AOI21_X1   g12385(.A1(new_n12609_), .A2(new_n12693_), .B(new_n12688_), .ZN(new_n12694_));
  NOR2_X1    g12386(.A1(new_n3837_), .A2(new_n4769_), .ZN(new_n12695_));
  AOI22_X1   g12387(.A1(new_n6024_), .A2(new_n12695_), .B1(new_n5350_), .B2(new_n5600_), .ZN(new_n12696_));
  INV_X1     g12388(.I(new_n12696_), .ZN(new_n12697_));
  NOR2_X1    g12389(.A1(new_n5340_), .A2(new_n6579_), .ZN(new_n12698_));
  INV_X1     g12390(.I(new_n12698_), .ZN(new_n12699_));
  NOR2_X1    g12391(.A1(new_n12697_), .A2(new_n12698_), .ZN(new_n12700_));
  AOI21_X1   g12392(.A1(new_n12700_), .A2(new_n6024_), .B(\a[41] ), .ZN(new_n12701_));
  NOR2_X1    g12393(.A1(\a[37] ), .A2(\a[42] ), .ZN(new_n12702_));
  OAI21_X1   g12394(.A1(new_n12701_), .A2(new_n3804_), .B(new_n12702_), .ZN(new_n12703_));
  AND3_X2    g12395(.A1(new_n12703_), .A2(new_n12697_), .A3(new_n12699_), .Z(new_n12704_));
  OAI21_X1   g12396(.A1(new_n8005_), .A2(new_n7486_), .B(new_n7149_), .ZN(new_n12705_));
  NOR2_X1    g12397(.A1(new_n1691_), .A2(new_n6999_), .ZN(new_n12706_));
  INV_X1     g12398(.I(new_n12706_), .ZN(new_n12707_));
  NOR4_X1    g12399(.A1(new_n12705_), .A2(new_n2752_), .A3(new_n7482_), .A4(new_n12707_), .ZN(new_n12708_));
  INV_X1     g12400(.I(new_n12708_), .ZN(new_n12709_));
  NAND3_X1   g12401(.A1(\a[28] ), .A2(\a[40] ), .A3(\a[51] ), .ZN(new_n12710_));
  XOR2_X1    g12402(.A1(new_n12710_), .A2(\a[17] ), .Z(new_n12711_));
  XOR2_X1    g12403(.A1(new_n12711_), .A2(\a[62] ), .Z(new_n12712_));
  NOR2_X1    g12404(.A1(new_n12709_), .A2(new_n12712_), .ZN(new_n12713_));
  INV_X1     g12405(.I(new_n12712_), .ZN(new_n12714_));
  NOR2_X1    g12406(.A1(new_n12714_), .A2(new_n12708_), .ZN(new_n12715_));
  OAI21_X1   g12407(.A1(new_n12713_), .A2(new_n12715_), .B(new_n12704_), .ZN(new_n12716_));
  XOR2_X1    g12408(.A1(new_n12712_), .A2(new_n12708_), .Z(new_n12717_));
  OAI21_X1   g12409(.A1(new_n12704_), .A2(new_n12717_), .B(new_n12716_), .ZN(new_n12718_));
  INV_X1     g12410(.I(new_n12508_), .ZN(new_n12719_));
  AOI21_X1   g12411(.A1(new_n12719_), .A2(new_n12490_), .B(new_n12507_), .ZN(new_n12720_));
  AOI22_X1   g12412(.A1(new_n1769_), .A2(new_n8996_), .B1(new_n9554_), .B2(new_n1798_), .ZN(new_n12721_));
  NOR2_X1    g12413(.A1(new_n1339_), .A2(new_n8990_), .ZN(new_n12722_));
  NAND4_X1   g12414(.A1(new_n12721_), .A2(new_n1711_), .A3(new_n8677_), .A4(new_n12722_), .ZN(new_n12723_));
  NAND2_X1   g12415(.A1(new_n2898_), .A2(new_n6280_), .ZN(new_n12724_));
  NAND2_X1   g12416(.A1(\a[22] ), .A2(\a[57] ), .ZN(new_n12725_));
  XNOR2_X1   g12417(.A1(new_n12724_), .A2(new_n12725_), .ZN(new_n12726_));
  NOR2_X1    g12418(.A1(new_n11818_), .A2(new_n11541_), .ZN(new_n12727_));
  NOR2_X1    g12419(.A1(new_n3852_), .A2(new_n5793_), .ZN(new_n12728_));
  AOI21_X1   g12420(.A1(\a[32] ), .A2(\a[47] ), .B(new_n5909_), .ZN(new_n12729_));
  NOR4_X1    g12421(.A1(new_n12728_), .A2(new_n2655_), .A3(new_n12729_), .A4(new_n5750_), .ZN(new_n12730_));
  NAND2_X1   g12422(.A1(new_n12730_), .A2(new_n12727_), .ZN(new_n12731_));
  NOR2_X1    g12423(.A1(new_n12731_), .A2(new_n12726_), .ZN(new_n12732_));
  AND2_X2    g12424(.A1(new_n12731_), .A2(new_n12726_), .Z(new_n12733_));
  NOR2_X1    g12425(.A1(new_n12733_), .A2(new_n12732_), .ZN(new_n12734_));
  NOR2_X1    g12426(.A1(new_n12734_), .A2(new_n12723_), .ZN(new_n12735_));
  INV_X1     g12427(.I(new_n12723_), .ZN(new_n12736_));
  XNOR2_X1   g12428(.A1(new_n12731_), .A2(new_n12726_), .ZN(new_n12737_));
  NOR2_X1    g12429(.A1(new_n12737_), .A2(new_n12736_), .ZN(new_n12738_));
  NOR2_X1    g12430(.A1(new_n12735_), .A2(new_n12738_), .ZN(new_n12739_));
  XNOR2_X1   g12431(.A1(new_n12720_), .A2(new_n12739_), .ZN(new_n12740_));
  INV_X1     g12432(.I(new_n12740_), .ZN(new_n12741_));
  OR2_X2     g12433(.A1(new_n12720_), .A2(new_n12739_), .Z(new_n12742_));
  NAND2_X1   g12434(.A1(new_n12720_), .A2(new_n12739_), .ZN(new_n12743_));
  AOI21_X1   g12435(.A1(new_n12742_), .A2(new_n12743_), .B(new_n12718_), .ZN(new_n12744_));
  AOI21_X1   g12436(.A1(new_n12741_), .A2(new_n12718_), .B(new_n12744_), .ZN(new_n12745_));
  OAI21_X1   g12437(.A1(new_n12411_), .A2(new_n12444_), .B(new_n12446_), .ZN(new_n12746_));
  INV_X1     g12438(.I(new_n12487_), .ZN(new_n12747_));
  AOI21_X1   g12439(.A1(new_n12475_), .A2(new_n12747_), .B(new_n12486_), .ZN(new_n12748_));
  INV_X1     g12440(.I(new_n12748_), .ZN(new_n12749_));
  OAI21_X1   g12441(.A1(new_n12553_), .A2(new_n12554_), .B(new_n12544_), .ZN(new_n12750_));
  OAI21_X1   g12442(.A1(new_n12548_), .A2(new_n12551_), .B(new_n12750_), .ZN(new_n12751_));
  INV_X1     g12443(.I(new_n12500_), .ZN(new_n12752_));
  AOI21_X1   g12444(.A1(new_n12491_), .A2(new_n12752_), .B(new_n12499_), .ZN(new_n12753_));
  INV_X1     g12445(.I(new_n12753_), .ZN(new_n12754_));
  XOR2_X1    g12446(.A1(new_n12751_), .A2(new_n12754_), .Z(new_n12755_));
  NAND2_X1   g12447(.A1(new_n12755_), .A2(new_n12749_), .ZN(new_n12756_));
  AND2_X2    g12448(.A1(new_n12751_), .A2(new_n12754_), .Z(new_n12757_));
  NOR2_X1    g12449(.A1(new_n12751_), .A2(new_n12754_), .ZN(new_n12758_));
  OAI21_X1   g12450(.A1(new_n12757_), .A2(new_n12758_), .B(new_n12748_), .ZN(new_n12759_));
  NAND2_X1   g12451(.A1(new_n12756_), .A2(new_n12759_), .ZN(new_n12760_));
  NAND2_X1   g12452(.A1(new_n12472_), .A2(new_n12469_), .ZN(new_n12761_));
  NAND2_X1   g12453(.A1(new_n12761_), .A2(new_n12471_), .ZN(new_n12762_));
  XNOR2_X1   g12454(.A1(new_n12762_), .A2(new_n12760_), .ZN(new_n12763_));
  NAND3_X1   g12455(.A1(new_n12762_), .A2(new_n12756_), .A3(new_n12759_), .ZN(new_n12764_));
  NAND3_X1   g12456(.A1(new_n12760_), .A2(new_n12471_), .A3(new_n12761_), .ZN(new_n12765_));
  AOI21_X1   g12457(.A1(new_n12764_), .A2(new_n12765_), .B(new_n12746_), .ZN(new_n12766_));
  AOI21_X1   g12458(.A1(new_n12746_), .A2(new_n12763_), .B(new_n12766_), .ZN(new_n12767_));
  NAND2_X1   g12459(.A1(new_n12519_), .A2(new_n12474_), .ZN(new_n12768_));
  NAND2_X1   g12460(.A1(new_n12768_), .A2(new_n12518_), .ZN(new_n12769_));
  NAND2_X1   g12461(.A1(new_n12769_), .A2(new_n12767_), .ZN(new_n12770_));
  INV_X1     g12462(.I(new_n12770_), .ZN(new_n12771_));
  NOR2_X1    g12463(.A1(new_n12769_), .A2(new_n12767_), .ZN(new_n12772_));
  NOR2_X1    g12464(.A1(new_n12771_), .A2(new_n12772_), .ZN(new_n12773_));
  XOR2_X1    g12465(.A1(new_n12769_), .A2(new_n12767_), .Z(new_n12774_));
  NAND2_X1   g12466(.A1(new_n12774_), .A2(new_n12745_), .ZN(new_n12775_));
  OAI21_X1   g12467(.A1(new_n12745_), .A2(new_n12773_), .B(new_n12775_), .ZN(new_n12776_));
  XOR2_X1    g12468(.A1(new_n12694_), .A2(new_n12776_), .Z(new_n12777_));
  XNOR2_X1   g12469(.A1(new_n12694_), .A2(new_n12776_), .ZN(new_n12778_));
  MUX2_X1    g12470(.I0(new_n12778_), .I1(new_n12777_), .S(new_n12607_), .Z(new_n12779_));
  XOR2_X1    g12471(.A1(new_n12779_), .A2(new_n12606_), .Z(new_n12780_));
  NAND2_X1   g12472(.A1(new_n12605_), .A2(new_n12780_), .ZN(new_n12781_));
  NOR2_X1    g12473(.A1(new_n12779_), .A2(new_n12606_), .ZN(new_n12782_));
  NAND2_X1   g12474(.A1(new_n12779_), .A2(new_n12606_), .ZN(new_n12783_));
  INV_X1     g12475(.I(new_n12783_), .ZN(new_n12784_));
  NOR2_X1    g12476(.A1(new_n12784_), .A2(new_n12782_), .ZN(new_n12785_));
  OAI21_X1   g12477(.A1(new_n12605_), .A2(new_n12785_), .B(new_n12781_), .ZN(\asquared[80] ));
  AOI21_X1   g12478(.A1(new_n12784_), .A2(new_n12598_), .B(new_n12406_), .ZN(new_n12787_));
  AOI21_X1   g12479(.A1(new_n12596_), .A2(new_n12783_), .B(new_n12787_), .ZN(new_n12788_));
  INV_X1     g12480(.I(new_n12788_), .ZN(new_n12789_));
  AOI21_X1   g12481(.A1(new_n12402_), .A2(new_n12400_), .B(new_n12789_), .ZN(new_n12790_));
  AND2_X2    g12482(.A1(new_n12790_), .A2(new_n12782_), .Z(\asquared[81] ));
  NAND2_X1   g12483(.A1(new_n12743_), .A2(new_n12718_), .ZN(new_n12792_));
  INV_X1     g12484(.I(new_n12715_), .ZN(new_n12793_));
  AOI21_X1   g12485(.A1(new_n12704_), .A2(new_n12793_), .B(new_n12713_), .ZN(new_n12794_));
  AOI21_X1   g12486(.A1(new_n2978_), .A2(new_n8676_), .B(new_n12721_), .ZN(new_n12795_));
  NOR2_X1    g12487(.A1(new_n2898_), .A2(new_n6280_), .ZN(new_n12796_));
  NAND2_X1   g12488(.A1(new_n1674_), .A2(new_n7727_), .ZN(new_n12797_));
  AOI21_X1   g12489(.A1(new_n2898_), .A2(new_n6280_), .B(new_n12797_), .ZN(new_n12798_));
  NOR2_X1    g12490(.A1(new_n12798_), .A2(new_n12796_), .ZN(new_n12799_));
  NOR2_X1    g12491(.A1(new_n12727_), .A2(new_n12728_), .ZN(new_n12800_));
  XOR2_X1    g12492(.A1(new_n12800_), .A2(new_n12799_), .Z(new_n12801_));
  NAND2_X1   g12493(.A1(new_n12801_), .A2(new_n12795_), .ZN(new_n12802_));
  INV_X1     g12494(.I(new_n12795_), .ZN(new_n12803_));
  NOR4_X1    g12495(.A1(new_n12798_), .A2(new_n12727_), .A3(new_n12796_), .A4(new_n12728_), .ZN(new_n12804_));
  NOR2_X1    g12496(.A1(new_n12800_), .A2(new_n12799_), .ZN(new_n12805_));
  OAI21_X1   g12497(.A1(new_n12805_), .A2(new_n12804_), .B(new_n12803_), .ZN(new_n12806_));
  NAND2_X1   g12498(.A1(new_n12802_), .A2(new_n12806_), .ZN(new_n12807_));
  NOR2_X1    g12499(.A1(new_n12733_), .A2(new_n12723_), .ZN(new_n12808_));
  NOR2_X1    g12500(.A1(new_n12808_), .A2(new_n12732_), .ZN(new_n12809_));
  XNOR2_X1   g12501(.A1(new_n12807_), .A2(new_n12809_), .ZN(new_n12810_));
  NOR2_X1    g12502(.A1(new_n12807_), .A2(new_n12809_), .ZN(new_n12811_));
  NAND2_X1   g12503(.A1(new_n12807_), .A2(new_n12809_), .ZN(new_n12812_));
  INV_X1     g12504(.I(new_n12812_), .ZN(new_n12813_));
  OAI21_X1   g12505(.A1(new_n12813_), .A2(new_n12811_), .B(new_n12794_), .ZN(new_n12814_));
  OAI21_X1   g12506(.A1(new_n12794_), .A2(new_n12810_), .B(new_n12814_), .ZN(new_n12815_));
  NOR2_X1    g12507(.A1(new_n12758_), .A2(new_n12748_), .ZN(new_n12816_));
  NOR2_X1    g12508(.A1(new_n12816_), .A2(new_n12757_), .ZN(new_n12817_));
  NOR2_X1    g12509(.A1(new_n12638_), .A2(new_n12641_), .ZN(new_n12818_));
  NOR2_X1    g12510(.A1(new_n12818_), .A2(new_n12639_), .ZN(new_n12819_));
  NAND2_X1   g12511(.A1(new_n3487_), .A2(new_n5742_), .ZN(new_n12820_));
  NOR2_X1    g12512(.A1(new_n3487_), .A2(new_n5742_), .ZN(new_n12821_));
  NOR2_X1    g12513(.A1(\a[16] ), .A2(\a[63] ), .ZN(new_n12822_));
  AOI21_X1   g12514(.A1(new_n12820_), .A2(new_n12822_), .B(new_n12821_), .ZN(new_n12823_));
  INV_X1     g12515(.I(new_n12823_), .ZN(new_n12824_));
  NAND2_X1   g12516(.A1(new_n3393_), .A2(new_n4501_), .ZN(new_n12825_));
  AOI21_X1   g12517(.A1(new_n11831_), .A2(new_n12631_), .B(new_n12825_), .ZN(new_n12826_));
  NOR2_X1    g12518(.A1(new_n12826_), .A2(new_n12633_), .ZN(new_n12827_));
  OAI21_X1   g12519(.A1(new_n2753_), .A2(new_n10288_), .B(new_n12705_), .ZN(new_n12828_));
  XOR2_X1    g12520(.A1(new_n12828_), .A2(new_n12827_), .Z(new_n12829_));
  NOR2_X1    g12521(.A1(new_n12829_), .A2(new_n12824_), .ZN(new_n12830_));
  INV_X1     g12522(.I(new_n12827_), .ZN(new_n12831_));
  NOR2_X1    g12523(.A1(new_n12828_), .A2(new_n12831_), .ZN(new_n12832_));
  INV_X1     g12524(.I(new_n12832_), .ZN(new_n12833_));
  NAND2_X1   g12525(.A1(new_n12828_), .A2(new_n12831_), .ZN(new_n12834_));
  AOI21_X1   g12526(.A1(new_n12833_), .A2(new_n12834_), .B(new_n12823_), .ZN(new_n12835_));
  NOR2_X1    g12527(.A1(new_n12830_), .A2(new_n12835_), .ZN(new_n12836_));
  XOR2_X1    g12528(.A1(new_n12819_), .A2(new_n12836_), .Z(new_n12837_));
  NOR3_X1    g12529(.A1(new_n12818_), .A2(new_n12639_), .A3(new_n12836_), .ZN(new_n12838_));
  NOR3_X1    g12530(.A1(new_n12819_), .A2(new_n12830_), .A3(new_n12835_), .ZN(new_n12839_));
  OAI21_X1   g12531(.A1(new_n12839_), .A2(new_n12838_), .B(new_n12817_), .ZN(new_n12840_));
  OAI21_X1   g12532(.A1(new_n12837_), .A2(new_n12817_), .B(new_n12840_), .ZN(new_n12841_));
  XNOR2_X1   g12533(.A1(new_n12841_), .A2(new_n12815_), .ZN(new_n12842_));
  AOI21_X1   g12534(.A1(new_n12742_), .A2(new_n12792_), .B(new_n12842_), .ZN(new_n12843_));
  NAND2_X1   g12535(.A1(new_n12792_), .A2(new_n12742_), .ZN(new_n12844_));
  NAND2_X1   g12536(.A1(new_n12841_), .A2(new_n12815_), .ZN(new_n12845_));
  NOR2_X1    g12537(.A1(new_n12841_), .A2(new_n12815_), .ZN(new_n12846_));
  INV_X1     g12538(.I(new_n12846_), .ZN(new_n12847_));
  AOI21_X1   g12539(.A1(new_n12847_), .A2(new_n12845_), .B(new_n12844_), .ZN(new_n12848_));
  NOR2_X1    g12540(.A1(new_n12614_), .A2(new_n12620_), .ZN(new_n12849_));
  NOR2_X1    g12541(.A1(new_n12849_), .A2(new_n12619_), .ZN(new_n12850_));
  NOR2_X1    g12542(.A1(new_n12669_), .A2(new_n12661_), .ZN(new_n12851_));
  NOR2_X1    g12543(.A1(new_n12851_), .A2(new_n12668_), .ZN(new_n12852_));
  NOR2_X1    g12544(.A1(new_n1276_), .A2(new_n8453_), .ZN(new_n12853_));
  OAI21_X1   g12545(.A1(new_n12655_), .A2(new_n12656_), .B(new_n12853_), .ZN(new_n12854_));
  NAND2_X1   g12546(.A1(new_n12854_), .A2(new_n12657_), .ZN(new_n12855_));
  XOR2_X1    g12547(.A1(new_n12852_), .A2(new_n12855_), .Z(new_n12856_));
  NOR2_X1    g12548(.A1(new_n12856_), .A2(new_n12850_), .ZN(new_n12857_));
  INV_X1     g12549(.I(new_n12850_), .ZN(new_n12858_));
  INV_X1     g12550(.I(new_n12855_), .ZN(new_n12859_));
  NOR2_X1    g12551(.A1(new_n12852_), .A2(new_n12859_), .ZN(new_n12860_));
  INV_X1     g12552(.I(new_n12860_), .ZN(new_n12861_));
  NAND2_X1   g12553(.A1(new_n12852_), .A2(new_n12859_), .ZN(new_n12862_));
  AOI21_X1   g12554(.A1(new_n12862_), .A2(new_n12861_), .B(new_n12858_), .ZN(new_n12863_));
  NOR2_X1    g12555(.A1(new_n12863_), .A2(new_n12857_), .ZN(new_n12864_));
  INV_X1     g12556(.I(new_n12643_), .ZN(new_n12865_));
  AOI21_X1   g12557(.A1(new_n12865_), .A2(new_n12623_), .B(new_n12645_), .ZN(new_n12866_));
  OAI21_X1   g12558(.A1(new_n12651_), .A2(new_n12675_), .B(new_n12676_), .ZN(new_n12867_));
  INV_X1     g12559(.I(new_n12867_), .ZN(new_n12868_));
  NOR2_X1    g12560(.A1(new_n12866_), .A2(new_n12868_), .ZN(new_n12869_));
  AND2_X2    g12561(.A1(new_n12866_), .A2(new_n12868_), .Z(new_n12870_));
  NOR2_X1    g12562(.A1(new_n12870_), .A2(new_n12869_), .ZN(new_n12871_));
  NOR2_X1    g12563(.A1(new_n12871_), .A2(new_n12864_), .ZN(new_n12872_));
  XOR2_X1    g12564(.A1(new_n12866_), .A2(new_n12867_), .Z(new_n12873_));
  NOR3_X1    g12565(.A1(new_n12873_), .A2(new_n12857_), .A3(new_n12863_), .ZN(new_n12874_));
  NOR4_X1    g12566(.A1(new_n12843_), .A2(new_n12848_), .A3(new_n12872_), .A4(new_n12874_), .ZN(new_n12875_));
  INV_X1     g12567(.I(new_n12772_), .ZN(new_n12876_));
  AOI21_X1   g12568(.A1(new_n12745_), .A2(new_n12876_), .B(new_n12771_), .ZN(new_n12877_));
  NOR2_X1    g12569(.A1(new_n12843_), .A2(new_n12848_), .ZN(new_n12878_));
  NOR2_X1    g12570(.A1(new_n12872_), .A2(new_n12874_), .ZN(new_n12879_));
  NOR2_X1    g12571(.A1(new_n12878_), .A2(new_n12879_), .ZN(new_n12880_));
  NOR2_X1    g12572(.A1(new_n12877_), .A2(new_n12880_), .ZN(new_n12881_));
  NOR2_X1    g12573(.A1(new_n12881_), .A2(new_n12875_), .ZN(new_n12882_));
  INV_X1     g12574(.I(new_n12882_), .ZN(new_n12883_));
  AOI21_X1   g12575(.A1(new_n12844_), .A2(new_n12845_), .B(new_n12846_), .ZN(new_n12884_));
  OAI21_X1   g12576(.A1(new_n2499_), .A2(new_n6694_), .B(new_n6999_), .ZN(new_n12885_));
  AOI21_X1   g12577(.A1(new_n3037_), .A2(new_n12418_), .B(new_n12885_), .ZN(new_n12886_));
  NOR3_X1    g12578(.A1(new_n12886_), .A2(new_n2689_), .A3(new_n8056_), .ZN(new_n12887_));
  AOI21_X1   g12579(.A1(\a[29] ), .A2(\a[52] ), .B(\a[53] ), .ZN(new_n12888_));
  NOR2_X1    g12580(.A1(\a[26] ), .A2(\a[55] ), .ZN(new_n12889_));
  OAI21_X1   g12581(.A1(new_n12888_), .A2(new_n2178_), .B(new_n12889_), .ZN(new_n12890_));
  NAND2_X1   g12582(.A1(new_n12887_), .A2(new_n12890_), .ZN(new_n12891_));
  INV_X1     g12583(.I(new_n11018_), .ZN(new_n12892_));
  OAI22_X1   g12584(.A1(new_n1536_), .A2(new_n9861_), .B1(new_n12892_), .B2(new_n3889_), .ZN(new_n12893_));
  NOR4_X1    g12585(.A1(new_n8991_), .A2(new_n2978_), .A3(new_n1276_), .A4(new_n9310_), .ZN(new_n12894_));
  NAND2_X1   g12586(.A1(new_n12893_), .A2(new_n12894_), .ZN(new_n12895_));
  NOR2_X1    g12587(.A1(new_n3423_), .A2(new_n5175_), .ZN(new_n12896_));
  NOR2_X1    g12588(.A1(new_n3839_), .A2(new_n5743_), .ZN(new_n12897_));
  NAND4_X1   g12589(.A1(new_n12897_), .A2(\a[37] ), .A3(\a[44] ), .A4(new_n12896_), .ZN(new_n12898_));
  AOI21_X1   g12590(.A1(new_n12898_), .A2(new_n8424_), .B(new_n3967_), .ZN(new_n12899_));
  NOR3_X1    g12591(.A1(new_n12895_), .A2(new_n3839_), .A3(new_n5743_), .ZN(new_n12900_));
  NOR2_X1    g12592(.A1(new_n3839_), .A2(new_n5743_), .ZN(new_n12901_));
  AOI21_X1   g12593(.A1(new_n12893_), .A2(new_n12894_), .B(new_n12901_), .ZN(new_n12902_));
  NOR2_X1    g12594(.A1(new_n12900_), .A2(new_n12902_), .ZN(new_n12903_));
  XOR2_X1    g12595(.A1(new_n12895_), .A2(new_n12901_), .Z(new_n12904_));
  MUX2_X1    g12596(.I0(new_n12903_), .I1(new_n12904_), .S(new_n12891_), .Z(new_n12905_));
  INV_X1     g12597(.I(new_n12905_), .ZN(new_n12906_));
  NAND2_X1   g12598(.A1(new_n12858_), .A2(new_n12862_), .ZN(new_n12907_));
  NAND2_X1   g12599(.A1(new_n12907_), .A2(new_n12861_), .ZN(new_n12908_));
  NOR2_X1    g12600(.A1(new_n1674_), .A2(new_n8085_), .ZN(new_n12909_));
  NOR2_X1    g12601(.A1(new_n8244_), .A2(new_n1912_), .ZN(new_n12910_));
  NAND3_X1   g12602(.A1(new_n12910_), .A2(new_n5357_), .A3(new_n8460_), .ZN(new_n12911_));
  AOI21_X1   g12603(.A1(new_n12911_), .A2(new_n8677_), .B(new_n2285_), .ZN(new_n12912_));
  NOR2_X1    g12604(.A1(new_n8244_), .A2(new_n1912_), .ZN(new_n12913_));
  XNOR2_X1   g12605(.A1(new_n4372_), .A2(new_n6030_), .ZN(new_n12914_));
  NOR2_X1    g12606(.A1(new_n4240_), .A2(new_n9029_), .ZN(new_n12915_));
  XNOR2_X1   g12607(.A1(new_n8191_), .A2(new_n12915_), .ZN(new_n12916_));
  NOR2_X1    g12608(.A1(new_n12914_), .A2(new_n12916_), .ZN(new_n12917_));
  AND2_X2    g12609(.A1(new_n12914_), .A2(new_n12916_), .Z(new_n12918_));
  NOR2_X1    g12610(.A1(new_n12918_), .A2(new_n12917_), .ZN(new_n12919_));
  XNOR2_X1   g12611(.A1(new_n12914_), .A2(new_n12916_), .ZN(new_n12920_));
  MUX2_X1    g12612(.I0(new_n12920_), .I1(new_n12919_), .S(new_n12913_), .Z(new_n12921_));
  XOR2_X1    g12613(.A1(new_n12908_), .A2(new_n12921_), .Z(new_n12922_));
  INV_X1     g12614(.I(new_n12922_), .ZN(new_n12923_));
  INV_X1     g12615(.I(new_n12908_), .ZN(new_n12924_));
  NOR2_X1    g12616(.A1(new_n12924_), .A2(new_n12921_), .ZN(new_n12925_));
  INV_X1     g12617(.I(new_n12925_), .ZN(new_n12926_));
  NAND2_X1   g12618(.A1(new_n12924_), .A2(new_n12921_), .ZN(new_n12927_));
  AOI21_X1   g12619(.A1(new_n12926_), .A2(new_n12927_), .B(new_n12906_), .ZN(new_n12928_));
  AOI21_X1   g12620(.A1(new_n12906_), .A2(new_n12923_), .B(new_n12928_), .ZN(new_n12929_));
  INV_X1     g12621(.I(new_n12929_), .ZN(new_n12930_));
  INV_X1     g12622(.I(new_n12870_), .ZN(new_n12931_));
  AOI21_X1   g12623(.A1(new_n12931_), .A2(new_n12864_), .B(new_n12869_), .ZN(new_n12932_));
  NOR2_X1    g12624(.A1(new_n12932_), .A2(new_n12930_), .ZN(new_n12933_));
  INV_X1     g12625(.I(new_n12933_), .ZN(new_n12934_));
  NAND2_X1   g12626(.A1(new_n12932_), .A2(new_n12930_), .ZN(new_n12935_));
  AOI21_X1   g12627(.A1(new_n12934_), .A2(new_n12935_), .B(new_n12884_), .ZN(new_n12936_));
  INV_X1     g12628(.I(new_n12884_), .ZN(new_n12937_));
  XOR2_X1    g12629(.A1(new_n12932_), .A2(new_n12929_), .Z(new_n12938_));
  NOR2_X1    g12630(.A1(new_n12938_), .A2(new_n12937_), .ZN(new_n12939_));
  NOR2_X1    g12631(.A1(new_n12939_), .A2(new_n12936_), .ZN(new_n12940_));
  NAND2_X1   g12632(.A1(new_n12746_), .A2(new_n12765_), .ZN(new_n12941_));
  NAND2_X1   g12633(.A1(new_n12941_), .A2(new_n12764_), .ZN(new_n12942_));
  AOI22_X1   g12634(.A1(new_n2978_), .A2(new_n9554_), .B1(new_n8996_), .B2(new_n4437_), .ZN(new_n12943_));
  NOR3_X1    g12635(.A1(new_n12909_), .A2(new_n1313_), .A3(new_n7647_), .ZN(new_n12944_));
  INV_X1     g12636(.I(new_n12909_), .ZN(new_n12945_));
  AOI21_X1   g12637(.A1(\a[21] ), .A2(\a[58] ), .B(new_n12945_), .ZN(new_n12946_));
  NOR2_X1    g12638(.A1(new_n1215_), .A2(new_n8990_), .ZN(new_n12947_));
  NOR4_X1    g12639(.A1(new_n12946_), .A2(new_n12943_), .A3(new_n12944_), .A4(new_n12947_), .ZN(new_n12948_));
  AOI21_X1   g12640(.A1(\a[58] ), .A2(\a[59] ), .B(new_n12948_), .ZN(new_n12949_));
  NOR2_X1    g12641(.A1(new_n12949_), .A2(new_n1773_), .ZN(new_n12950_));
  AOI22_X1   g12642(.A1(new_n2766_), .A2(new_n6280_), .B1(new_n3126_), .B2(new_n6056_), .ZN(new_n12951_));
  NOR4_X1    g12643(.A1(new_n3981_), .A2(new_n6028_), .A3(new_n2461_), .A4(new_n6055_), .ZN(new_n12952_));
  NAND2_X1   g12644(.A1(new_n12952_), .A2(new_n12951_), .ZN(new_n12953_));
  NOR2_X1    g12645(.A1(new_n12950_), .A2(new_n12953_), .ZN(new_n12954_));
  INV_X1     g12646(.I(new_n12954_), .ZN(new_n12955_));
  NAND2_X1   g12647(.A1(new_n12950_), .A2(new_n12953_), .ZN(new_n12956_));
  NAND2_X1   g12648(.A1(new_n12955_), .A2(new_n12956_), .ZN(new_n12957_));
  XNOR2_X1   g12649(.A1(new_n12950_), .A2(new_n12953_), .ZN(new_n12958_));
  NOR2_X1    g12650(.A1(new_n12958_), .A2(new_n12700_), .ZN(new_n12959_));
  AOI21_X1   g12651(.A1(new_n12700_), .A2(new_n12957_), .B(new_n12959_), .ZN(new_n12960_));
  INV_X1     g12652(.I(new_n12960_), .ZN(new_n12961_));
  NOR2_X1    g12653(.A1(new_n7422_), .A2(new_n2679_), .ZN(new_n12962_));
  NOR2_X1    g12654(.A1(new_n6945_), .A2(new_n7727_), .ZN(new_n12964_));
  INV_X1     g12655(.I(new_n12964_), .ZN(new_n12965_));
  NOR2_X1    g12656(.A1(new_n7422_), .A2(new_n2679_), .ZN(new_n12969_));
  NAND2_X1   g12657(.A1(new_n5173_), .A2(new_n5600_), .ZN(new_n12970_));
  NAND2_X1   g12658(.A1(\a[25] ), .A2(\a[55] ), .ZN(new_n12971_));
  XNOR2_X1   g12659(.A1(new_n12970_), .A2(new_n12971_), .ZN(new_n12972_));
  NAND2_X1   g12660(.A1(\a[52] ), .A2(\a[53] ), .ZN(new_n12973_));
  XNOR2_X1   g12661(.A1(new_n2692_), .A2(new_n12973_), .ZN(new_n12974_));
  NOR2_X1    g12662(.A1(new_n12972_), .A2(new_n12974_), .ZN(new_n12975_));
  AND2_X2    g12663(.A1(new_n12972_), .A2(new_n12974_), .Z(new_n12976_));
  NOR2_X1    g12664(.A1(new_n12976_), .A2(new_n12975_), .ZN(new_n12977_));
  XNOR2_X1   g12665(.A1(new_n12972_), .A2(new_n12974_), .ZN(new_n12978_));
  MUX2_X1    g12666(.I0(new_n12978_), .I1(new_n12977_), .S(new_n12969_), .Z(new_n12979_));
  NAND4_X1   g12667(.A1(\a[17] ), .A2(\a[29] ), .A3(\a[51] ), .A4(\a[63] ), .ZN(new_n12980_));
  NAND2_X1   g12668(.A1(\a[33] ), .A2(\a[47] ), .ZN(new_n12981_));
  XNOR2_X1   g12669(.A1(new_n12980_), .A2(new_n12981_), .ZN(new_n12982_));
  AOI22_X1   g12670(.A1(new_n3487_), .A2(new_n7452_), .B1(new_n4727_), .B2(new_n5488_), .ZN(new_n12983_));
  NOR2_X1    g12671(.A1(new_n3371_), .A2(new_n5175_), .ZN(new_n12984_));
  NAND4_X1   g12672(.A1(new_n12983_), .A2(new_n3967_), .A3(new_n5743_), .A4(new_n12984_), .ZN(new_n12985_));
  AOI21_X1   g12673(.A1(\a[28] ), .A2(\a[51] ), .B(\a[40] ), .ZN(new_n12986_));
  NAND2_X1   g12674(.A1(\a[17] ), .A2(\a[62] ), .ZN(new_n12987_));
  OAI21_X1   g12675(.A1(new_n12986_), .A2(new_n12987_), .B(new_n12710_), .ZN(new_n12988_));
  NAND2_X1   g12676(.A1(\a[19] ), .A2(\a[62] ), .ZN(new_n12989_));
  XNOR2_X1   g12677(.A1(new_n12853_), .A2(new_n12989_), .ZN(new_n12990_));
  NAND2_X1   g12678(.A1(new_n12990_), .A2(new_n12988_), .ZN(new_n12991_));
  INV_X1     g12679(.I(new_n12991_), .ZN(new_n12992_));
  NOR2_X1    g12680(.A1(new_n12990_), .A2(new_n12988_), .ZN(new_n12993_));
  NOR2_X1    g12681(.A1(new_n12992_), .A2(new_n12993_), .ZN(new_n12994_));
  NOR2_X1    g12682(.A1(new_n12994_), .A2(new_n12985_), .ZN(new_n12995_));
  INV_X1     g12683(.I(new_n12985_), .ZN(new_n12996_));
  NOR3_X1    g12684(.A1(new_n12992_), .A2(new_n12996_), .A3(new_n12993_), .ZN(new_n12997_));
  NOR2_X1    g12685(.A1(new_n12995_), .A2(new_n12997_), .ZN(new_n12998_));
  NOR2_X1    g12686(.A1(new_n12998_), .A2(new_n12982_), .ZN(new_n12999_));
  INV_X1     g12687(.I(new_n12982_), .ZN(new_n13000_));
  XOR2_X1    g12688(.A1(new_n12994_), .A2(new_n12996_), .Z(new_n13001_));
  NOR2_X1    g12689(.A1(new_n13001_), .A2(new_n13000_), .ZN(new_n13002_));
  NOR2_X1    g12690(.A1(new_n13002_), .A2(new_n12999_), .ZN(new_n13003_));
  XOR2_X1    g12691(.A1(new_n13003_), .A2(new_n12979_), .Z(new_n13004_));
  NOR2_X1    g12692(.A1(new_n13003_), .A2(new_n12979_), .ZN(new_n13005_));
  INV_X1     g12693(.I(new_n13005_), .ZN(new_n13006_));
  NAND2_X1   g12694(.A1(new_n13003_), .A2(new_n12979_), .ZN(new_n13007_));
  AOI21_X1   g12695(.A1(new_n13006_), .A2(new_n13007_), .B(new_n12961_), .ZN(new_n13008_));
  AOI21_X1   g12696(.A1(new_n12961_), .A2(new_n13004_), .B(new_n13008_), .ZN(new_n13009_));
  NAND2_X1   g12697(.A1(new_n12942_), .A2(new_n13009_), .ZN(new_n13010_));
  OAI21_X1   g12698(.A1(new_n12612_), .A2(new_n12682_), .B(new_n12683_), .ZN(new_n13011_));
  INV_X1     g12699(.I(new_n13011_), .ZN(new_n13012_));
  NOR2_X1    g12700(.A1(new_n12942_), .A2(new_n13009_), .ZN(new_n13013_));
  OAI21_X1   g12701(.A1(new_n13012_), .A2(new_n13013_), .B(new_n13010_), .ZN(new_n13014_));
  NOR2_X1    g12702(.A1(new_n12813_), .A2(new_n12794_), .ZN(new_n13015_));
  NOR2_X1    g12703(.A1(new_n13015_), .A2(new_n12811_), .ZN(new_n13016_));
  NOR2_X1    g12704(.A1(new_n12838_), .A2(new_n12817_), .ZN(new_n13017_));
  NOR2_X1    g12705(.A1(new_n13017_), .A2(new_n12839_), .ZN(new_n13018_));
  NOR2_X1    g12706(.A1(new_n12805_), .A2(new_n12803_), .ZN(new_n13019_));
  NOR2_X1    g12707(.A1(new_n13019_), .A2(new_n12804_), .ZN(new_n13020_));
  NAND2_X1   g12708(.A1(new_n12834_), .A2(new_n12823_), .ZN(new_n13021_));
  NAND2_X1   g12709(.A1(new_n13021_), .A2(new_n12833_), .ZN(new_n13022_));
  NOR2_X1    g12710(.A1(new_n2098_), .A2(new_n6945_), .ZN(new_n13023_));
  XNOR2_X1   g12711(.A1(new_n5173_), .A2(new_n5339_), .ZN(new_n13024_));
  XOR2_X1    g12712(.A1(new_n13022_), .A2(new_n13024_), .Z(new_n13025_));
  NOR2_X1    g12713(.A1(new_n13025_), .A2(new_n13020_), .ZN(new_n13026_));
  INV_X1     g12714(.I(new_n13020_), .ZN(new_n13027_));
  INV_X1     g12715(.I(new_n13022_), .ZN(new_n13028_));
  NOR2_X1    g12716(.A1(new_n13028_), .A2(new_n13024_), .ZN(new_n13029_));
  INV_X1     g12717(.I(new_n13029_), .ZN(new_n13030_));
  NAND2_X1   g12718(.A1(new_n13028_), .A2(new_n13024_), .ZN(new_n13031_));
  AOI21_X1   g12719(.A1(new_n13030_), .A2(new_n13031_), .B(new_n13027_), .ZN(new_n13032_));
  NOR2_X1    g12720(.A1(new_n13032_), .A2(new_n13026_), .ZN(new_n13033_));
  XOR2_X1    g12721(.A1(new_n13018_), .A2(new_n13033_), .Z(new_n13034_));
  NOR2_X1    g12722(.A1(new_n13034_), .A2(new_n13016_), .ZN(new_n13035_));
  INV_X1     g12723(.I(new_n13016_), .ZN(new_n13036_));
  INV_X1     g12724(.I(new_n13018_), .ZN(new_n13037_));
  NOR2_X1    g12725(.A1(new_n13037_), .A2(new_n13033_), .ZN(new_n13038_));
  INV_X1     g12726(.I(new_n13038_), .ZN(new_n13039_));
  NAND2_X1   g12727(.A1(new_n13037_), .A2(new_n13033_), .ZN(new_n13040_));
  AOI21_X1   g12728(.A1(new_n13039_), .A2(new_n13040_), .B(new_n13036_), .ZN(new_n13041_));
  AOI21_X1   g12729(.A1(new_n12961_), .A2(new_n13007_), .B(new_n13005_), .ZN(new_n13042_));
  AOI21_X1   g12730(.A1(new_n2543_), .A2(new_n8242_), .B(new_n12962_), .ZN(new_n13043_));
  INV_X1     g12731(.I(new_n13043_), .ZN(new_n13044_));
  NOR2_X1    g12732(.A1(\a[25] ), .A2(\a[55] ), .ZN(new_n13045_));
  OAI21_X1   g12733(.A1(new_n5174_), .A2(new_n4706_), .B(new_n13045_), .ZN(new_n13046_));
  OAI21_X1   g12734(.A1(new_n5600_), .A2(new_n5173_), .B(new_n13046_), .ZN(new_n13047_));
  AOI21_X1   g12735(.A1(new_n2797_), .A2(new_n4415_), .B(new_n7204_), .ZN(new_n13048_));
  XNOR2_X1   g12736(.A1(new_n13047_), .A2(new_n13048_), .ZN(new_n13049_));
  NOR2_X1    g12737(.A1(new_n13049_), .A2(new_n13044_), .ZN(new_n13050_));
  NOR2_X1    g12738(.A1(new_n13047_), .A2(new_n13048_), .ZN(new_n13051_));
  INV_X1     g12739(.I(new_n13051_), .ZN(new_n13052_));
  NAND2_X1   g12740(.A1(new_n13047_), .A2(new_n13048_), .ZN(new_n13053_));
  AOI21_X1   g12741(.A1(new_n13052_), .A2(new_n13053_), .B(new_n13043_), .ZN(new_n13054_));
  NOR2_X1    g12742(.A1(new_n13050_), .A2(new_n13054_), .ZN(new_n13055_));
  INV_X1     g12743(.I(new_n12976_), .ZN(new_n13056_));
  AOI21_X1   g12744(.A1(new_n13056_), .A2(new_n12969_), .B(new_n12975_), .ZN(new_n13057_));
  NAND2_X1   g12745(.A1(new_n12956_), .A2(new_n12700_), .ZN(new_n13058_));
  NAND2_X1   g12746(.A1(new_n13058_), .A2(new_n12955_), .ZN(new_n13059_));
  INV_X1     g12747(.I(new_n13059_), .ZN(new_n13060_));
  NOR2_X1    g12748(.A1(new_n13060_), .A2(new_n13057_), .ZN(new_n13061_));
  INV_X1     g12749(.I(new_n13057_), .ZN(new_n13062_));
  NOR2_X1    g12750(.A1(new_n13059_), .A2(new_n13062_), .ZN(new_n13063_));
  NOR2_X1    g12751(.A1(new_n13061_), .A2(new_n13063_), .ZN(new_n13064_));
  NOR2_X1    g12752(.A1(new_n13064_), .A2(new_n13055_), .ZN(new_n13065_));
  XOR2_X1    g12753(.A1(new_n13059_), .A2(new_n13057_), .Z(new_n13066_));
  NOR3_X1    g12754(.A1(new_n13066_), .A2(new_n13050_), .A3(new_n13054_), .ZN(new_n13067_));
  NOR2_X1    g12755(.A1(new_n13065_), .A2(new_n13067_), .ZN(new_n13068_));
  NAND2_X1   g12756(.A1(new_n9784_), .A2(new_n2331_), .ZN(new_n13069_));
  AOI21_X1   g12757(.A1(new_n3966_), .A2(new_n5742_), .B(new_n12983_), .ZN(new_n13070_));
  NOR2_X1    g12758(.A1(new_n3849_), .A2(new_n3127_), .ZN(new_n13071_));
  NOR2_X1    g12759(.A1(new_n12545_), .A2(new_n13071_), .ZN(new_n13072_));
  NOR4_X1    g12760(.A1(new_n3981_), .A2(new_n6280_), .A3(new_n2461_), .A4(new_n6260_), .ZN(new_n13073_));
  NAND3_X1   g12761(.A1(new_n13070_), .A2(new_n13072_), .A3(new_n13073_), .ZN(new_n13074_));
  XOR2_X1    g12762(.A1(new_n13074_), .A2(new_n12993_), .Z(new_n13075_));
  XNOR2_X1   g12763(.A1(new_n13075_), .A2(new_n13069_), .ZN(new_n13076_));
  NOR2_X1    g12764(.A1(new_n2499_), .A2(new_n9310_), .ZN(new_n13077_));
  NAND2_X1   g12765(.A1(new_n7458_), .A2(new_n13077_), .ZN(new_n13078_));
  NOR2_X1    g12766(.A1(new_n6260_), .A2(new_n9310_), .ZN(new_n13079_));
  AOI21_X1   g12767(.A1(\a[17] ), .A2(\a[29] ), .B(new_n13079_), .ZN(new_n13080_));
  NOR2_X1    g12768(.A1(\a[33] ), .A2(\a[47] ), .ZN(new_n13081_));
  AOI21_X1   g12769(.A1(new_n13078_), .A2(new_n13081_), .B(new_n13080_), .ZN(new_n13082_));
  INV_X1     g12770(.I(new_n13082_), .ZN(new_n13083_));
  AOI21_X1   g12771(.A1(new_n3981_), .A2(new_n6028_), .B(new_n12951_), .ZN(new_n13084_));
  AOI21_X1   g12772(.A1(new_n4538_), .A2(new_n8676_), .B(new_n12943_), .ZN(new_n13085_));
  XNOR2_X1   g12773(.A1(new_n13084_), .A2(new_n13085_), .ZN(new_n13086_));
  NOR2_X1    g12774(.A1(new_n13086_), .A2(new_n13083_), .ZN(new_n13087_));
  INV_X1     g12775(.I(new_n13084_), .ZN(new_n13088_));
  INV_X1     g12776(.I(new_n13085_), .ZN(new_n13089_));
  NOR2_X1    g12777(.A1(new_n13088_), .A2(new_n13089_), .ZN(new_n13090_));
  NOR2_X1    g12778(.A1(new_n13084_), .A2(new_n13085_), .ZN(new_n13091_));
  NOR2_X1    g12779(.A1(new_n13090_), .A2(new_n13091_), .ZN(new_n13092_));
  NOR2_X1    g12780(.A1(new_n13092_), .A2(new_n13082_), .ZN(new_n13093_));
  NOR2_X1    g12781(.A1(new_n13093_), .A2(new_n13087_), .ZN(new_n13094_));
  INV_X1     g12782(.I(new_n13094_), .ZN(new_n13095_));
  INV_X1     g12783(.I(new_n12997_), .ZN(new_n13096_));
  AOI21_X1   g12784(.A1(new_n13096_), .A2(new_n13000_), .B(new_n12995_), .ZN(new_n13097_));
  NOR2_X1    g12785(.A1(new_n13095_), .A2(new_n13097_), .ZN(new_n13098_));
  INV_X1     g12786(.I(new_n13097_), .ZN(new_n13099_));
  NOR2_X1    g12787(.A1(new_n13099_), .A2(new_n13094_), .ZN(new_n13100_));
  NOR2_X1    g12788(.A1(new_n13098_), .A2(new_n13100_), .ZN(new_n13101_));
  NOR2_X1    g12789(.A1(new_n13101_), .A2(new_n13076_), .ZN(new_n13102_));
  INV_X1     g12790(.I(new_n13076_), .ZN(new_n13103_));
  XOR2_X1    g12791(.A1(new_n13094_), .A2(new_n13097_), .Z(new_n13104_));
  NOR2_X1    g12792(.A1(new_n13104_), .A2(new_n13103_), .ZN(new_n13105_));
  NOR2_X1    g12793(.A1(new_n13102_), .A2(new_n13105_), .ZN(new_n13106_));
  XOR2_X1    g12794(.A1(new_n13068_), .A2(new_n13106_), .Z(new_n13107_));
  INV_X1     g12795(.I(new_n13068_), .ZN(new_n13108_));
  NOR2_X1    g12796(.A1(new_n13108_), .A2(new_n13106_), .ZN(new_n13109_));
  NAND2_X1   g12797(.A1(new_n13108_), .A2(new_n13106_), .ZN(new_n13110_));
  INV_X1     g12798(.I(new_n13110_), .ZN(new_n13111_));
  OAI21_X1   g12799(.A1(new_n13111_), .A2(new_n13109_), .B(new_n13042_), .ZN(new_n13112_));
  OAI21_X1   g12800(.A1(new_n13042_), .A2(new_n13107_), .B(new_n13112_), .ZN(new_n13113_));
  OAI21_X1   g12801(.A1(new_n13035_), .A2(new_n13041_), .B(new_n13113_), .ZN(new_n13114_));
  NOR2_X1    g12802(.A1(new_n13041_), .A2(new_n13035_), .ZN(new_n13115_));
  INV_X1     g12803(.I(new_n13113_), .ZN(new_n13116_));
  NAND2_X1   g12804(.A1(new_n13116_), .A2(new_n13115_), .ZN(new_n13117_));
  NAND2_X1   g12805(.A1(new_n13117_), .A2(new_n13114_), .ZN(new_n13118_));
  XOR2_X1    g12806(.A1(new_n13113_), .A2(new_n13115_), .Z(new_n13119_));
  NOR2_X1    g12807(.A1(new_n13119_), .A2(new_n13014_), .ZN(new_n13120_));
  AOI21_X1   g12808(.A1(new_n13014_), .A2(new_n13118_), .B(new_n13120_), .ZN(new_n13121_));
  NOR2_X1    g12809(.A1(new_n13121_), .A2(new_n12940_), .ZN(new_n13122_));
  NAND2_X1   g12810(.A1(new_n13121_), .A2(new_n12940_), .ZN(new_n13123_));
  INV_X1     g12811(.I(new_n13123_), .ZN(new_n13124_));
  OAI21_X1   g12812(.A1(new_n13124_), .A2(new_n13122_), .B(new_n12883_), .ZN(new_n13125_));
  XNOR2_X1   g12813(.A1(new_n13121_), .A2(new_n12940_), .ZN(new_n13126_));
  OAI21_X1   g12814(.A1(new_n12883_), .A2(new_n13126_), .B(new_n13125_), .ZN(new_n13127_));
  XNOR2_X1   g12815(.A1(new_n12878_), .A2(new_n12879_), .ZN(new_n13128_));
  OAI21_X1   g12816(.A1(new_n12875_), .A2(new_n12880_), .B(new_n12877_), .ZN(new_n13129_));
  OAI21_X1   g12817(.A1(new_n12877_), .A2(new_n13128_), .B(new_n13129_), .ZN(new_n13130_));
  XNOR2_X1   g12818(.A1(new_n12942_), .A2(new_n13009_), .ZN(new_n13131_));
  INV_X1     g12819(.I(new_n13010_), .ZN(new_n13132_));
  OAI21_X1   g12820(.A1(new_n13132_), .A2(new_n13013_), .B(new_n13012_), .ZN(new_n13133_));
  OAI21_X1   g12821(.A1(new_n13012_), .A2(new_n13131_), .B(new_n13133_), .ZN(new_n13134_));
  OAI21_X1   g12822(.A1(new_n12609_), .A2(new_n12690_), .B(new_n12692_), .ZN(new_n13135_));
  NAND2_X1   g12823(.A1(new_n13130_), .A2(new_n13134_), .ZN(new_n13136_));
  NAND2_X1   g12824(.A1(new_n13136_), .A2(new_n13135_), .ZN(new_n13137_));
  OAI21_X1   g12825(.A1(new_n13130_), .A2(new_n13134_), .B(new_n13137_), .ZN(new_n13138_));
  XOR2_X1    g12826(.A1(new_n13127_), .A2(new_n13138_), .Z(new_n13139_));
  NAND2_X1   g12827(.A1(\asquared[81] ), .A2(new_n13139_), .ZN(new_n13140_));
  NAND2_X1   g12828(.A1(new_n13127_), .A2(new_n13138_), .ZN(new_n13141_));
  OR2_X2     g12829(.A1(new_n13127_), .A2(new_n13138_), .Z(new_n13142_));
  AND2_X2    g12830(.A1(new_n13142_), .A2(new_n13141_), .Z(new_n13143_));
  OAI21_X1   g12831(.A1(\asquared[81] ), .A2(new_n13143_), .B(new_n13140_), .ZN(\asquared[82] ));
  NAND2_X1   g12832(.A1(\asquared[81] ), .A2(new_n13142_), .ZN(new_n13145_));
  NAND2_X1   g12833(.A1(new_n13145_), .A2(new_n13141_), .ZN(new_n13146_));
  AOI21_X1   g12834(.A1(new_n12937_), .A2(new_n12935_), .B(new_n12933_), .ZN(new_n13147_));
  AOI21_X1   g12835(.A1(new_n12906_), .A2(new_n12927_), .B(new_n12925_), .ZN(new_n13148_));
  NOR2_X1    g12836(.A1(new_n12891_), .A2(new_n12902_), .ZN(new_n13149_));
  NAND2_X1   g12837(.A1(new_n7204_), .A2(new_n2690_), .ZN(new_n13150_));
  AOI21_X1   g12838(.A1(new_n3981_), .A2(new_n6280_), .B(new_n13072_), .ZN(new_n13151_));
  AOI21_X1   g12839(.A1(new_n4372_), .A2(new_n9798_), .B(new_n6030_), .ZN(new_n13152_));
  XOR2_X1    g12840(.A1(new_n13151_), .A2(new_n13152_), .Z(new_n13153_));
  INV_X1     g12841(.I(new_n13153_), .ZN(new_n13154_));
  INV_X1     g12842(.I(new_n13151_), .ZN(new_n13155_));
  NOR2_X1    g12843(.A1(new_n13155_), .A2(new_n13152_), .ZN(new_n13156_));
  INV_X1     g12844(.I(new_n13156_), .ZN(new_n13157_));
  NAND2_X1   g12845(.A1(new_n13155_), .A2(new_n13152_), .ZN(new_n13158_));
  AOI21_X1   g12846(.A1(new_n13157_), .A2(new_n13158_), .B(new_n13150_), .ZN(new_n13159_));
  AOI21_X1   g12847(.A1(new_n13150_), .A2(new_n13154_), .B(new_n13159_), .ZN(new_n13160_));
  NOR2_X1    g12848(.A1(new_n12912_), .A2(new_n12910_), .ZN(new_n13161_));
  AOI21_X1   g12849(.A1(new_n2978_), .A2(new_n8991_), .B(new_n12893_), .ZN(new_n13162_));
  INV_X1     g12850(.I(new_n13162_), .ZN(new_n13163_));
  NOR2_X1    g12851(.A1(new_n12899_), .A2(new_n12897_), .ZN(new_n13164_));
  XOR2_X1    g12852(.A1(new_n13164_), .A2(new_n13163_), .Z(new_n13165_));
  INV_X1     g12853(.I(new_n13164_), .ZN(new_n13166_));
  NOR2_X1    g12854(.A1(new_n13166_), .A2(new_n13163_), .ZN(new_n13167_));
  NOR2_X1    g12855(.A1(new_n13164_), .A2(new_n13162_), .ZN(new_n13168_));
  NOR2_X1    g12856(.A1(new_n13167_), .A2(new_n13168_), .ZN(new_n13169_));
  MUX2_X1    g12857(.I0(new_n13169_), .I1(new_n13165_), .S(new_n13161_), .Z(new_n13170_));
  XOR2_X1    g12858(.A1(new_n13170_), .A2(new_n13160_), .Z(new_n13171_));
  OAI21_X1   g12859(.A1(new_n12900_), .A2(new_n13149_), .B(new_n13171_), .ZN(new_n13172_));
  NOR2_X1    g12860(.A1(new_n13149_), .A2(new_n12900_), .ZN(new_n13173_));
  NOR2_X1    g12861(.A1(new_n13170_), .A2(new_n13160_), .ZN(new_n13174_));
  NAND2_X1   g12862(.A1(new_n13170_), .A2(new_n13160_), .ZN(new_n13175_));
  INV_X1     g12863(.I(new_n13175_), .ZN(new_n13176_));
  OAI21_X1   g12864(.A1(new_n13176_), .A2(new_n13174_), .B(new_n13173_), .ZN(new_n13177_));
  NAND2_X1   g12865(.A1(new_n13172_), .A2(new_n13177_), .ZN(new_n13178_));
  INV_X1     g12866(.I(new_n12918_), .ZN(new_n13179_));
  AOI21_X1   g12867(.A1(new_n13179_), .A2(new_n12913_), .B(new_n12917_), .ZN(new_n13180_));
  NAND2_X1   g12868(.A1(new_n12993_), .A2(new_n13070_), .ZN(new_n13181_));
  NAND2_X1   g12869(.A1(new_n13072_), .A2(new_n13073_), .ZN(new_n13182_));
  NOR2_X1    g12870(.A1(new_n13182_), .A2(new_n13069_), .ZN(new_n13183_));
  OAI21_X1   g12871(.A1(new_n12993_), .A2(new_n13070_), .B(new_n13183_), .ZN(new_n13184_));
  NAND2_X1   g12872(.A1(new_n13184_), .A2(new_n13181_), .ZN(new_n13185_));
  NOR2_X1    g12873(.A1(new_n4414_), .A2(new_n9029_), .ZN(new_n13186_));
  AOI21_X1   g12874(.A1(\a[19] ), .A2(new_n13186_), .B(new_n5592_), .ZN(new_n13187_));
  INV_X1     g12875(.I(new_n13187_), .ZN(new_n13188_));
  AOI21_X1   g12876(.A1(new_n5173_), .A2(new_n13023_), .B(new_n5339_), .ZN(new_n13189_));
  NOR2_X1    g12877(.A1(new_n13188_), .A2(new_n13189_), .ZN(new_n13190_));
  XOR2_X1    g12878(.A1(new_n13190_), .A2(new_n1339_), .Z(new_n13191_));
  XOR2_X1    g12879(.A1(new_n13191_), .A2(\a[63] ), .Z(new_n13192_));
  XNOR2_X1   g12880(.A1(new_n13192_), .A2(new_n13185_), .ZN(new_n13193_));
  NOR2_X1    g12881(.A1(new_n13193_), .A2(new_n13180_), .ZN(new_n13194_));
  NOR2_X1    g12882(.A1(new_n13192_), .A2(new_n13185_), .ZN(new_n13195_));
  INV_X1     g12883(.I(new_n13195_), .ZN(new_n13196_));
  NAND2_X1   g12884(.A1(new_n13192_), .A2(new_n13185_), .ZN(new_n13197_));
  NAND2_X1   g12885(.A1(new_n13196_), .A2(new_n13197_), .ZN(new_n13198_));
  AOI21_X1   g12886(.A1(new_n13180_), .A2(new_n13198_), .B(new_n13194_), .ZN(new_n13199_));
  XOR2_X1    g12887(.A1(new_n13178_), .A2(new_n13199_), .Z(new_n13200_));
  NOR2_X1    g12888(.A1(new_n13200_), .A2(new_n13148_), .ZN(new_n13201_));
  INV_X1     g12889(.I(new_n13178_), .ZN(new_n13202_));
  NOR2_X1    g12890(.A1(new_n13202_), .A2(new_n13199_), .ZN(new_n13203_));
  INV_X1     g12891(.I(new_n13203_), .ZN(new_n13204_));
  NAND2_X1   g12892(.A1(new_n13202_), .A2(new_n13199_), .ZN(new_n13205_));
  NAND2_X1   g12893(.A1(new_n13204_), .A2(new_n13205_), .ZN(new_n13206_));
  AOI21_X1   g12894(.A1(new_n13148_), .A2(new_n13206_), .B(new_n13201_), .ZN(new_n13207_));
  AOI21_X1   g12895(.A1(new_n13043_), .A2(new_n13053_), .B(new_n13051_), .ZN(new_n13208_));
  NOR2_X1    g12896(.A1(new_n13091_), .A2(new_n13083_), .ZN(new_n13209_));
  NOR2_X1    g12897(.A1(new_n13209_), .A2(new_n13090_), .ZN(new_n13210_));
  NOR2_X1    g12898(.A1(new_n2891_), .A2(new_n10959_), .ZN(new_n13211_));
  NAND4_X1   g12899(.A1(new_n13211_), .A2(\a[25] ), .A3(\a[57] ), .A4(new_n7219_), .ZN(new_n13212_));
  AOI21_X1   g12900(.A1(new_n13212_), .A2(new_n8005_), .B(new_n2692_), .ZN(new_n13213_));
  NOR3_X1    g12901(.A1(new_n2891_), .A2(new_n6999_), .A3(new_n7727_), .ZN(new_n13214_));
  XOR2_X1    g12902(.A1(new_n13210_), .A2(new_n13214_), .Z(new_n13215_));
  NOR2_X1    g12903(.A1(new_n13215_), .A2(new_n13208_), .ZN(new_n13216_));
  INV_X1     g12904(.I(new_n13208_), .ZN(new_n13217_));
  INV_X1     g12905(.I(new_n13214_), .ZN(new_n13218_));
  NOR2_X1    g12906(.A1(new_n13210_), .A2(new_n13218_), .ZN(new_n13219_));
  INV_X1     g12907(.I(new_n13219_), .ZN(new_n13220_));
  NAND2_X1   g12908(.A1(new_n13210_), .A2(new_n13218_), .ZN(new_n13221_));
  AOI21_X1   g12909(.A1(new_n13220_), .A2(new_n13221_), .B(new_n13217_), .ZN(new_n13222_));
  NOR2_X1    g12910(.A1(new_n13216_), .A2(new_n13222_), .ZN(new_n13223_));
  INV_X1     g12911(.I(new_n13063_), .ZN(new_n13224_));
  AOI21_X1   g12912(.A1(new_n13055_), .A2(new_n13224_), .B(new_n13061_), .ZN(new_n13225_));
  NOR2_X1    g12913(.A1(new_n13100_), .A2(new_n13076_), .ZN(new_n13226_));
  NOR2_X1    g12914(.A1(new_n13226_), .A2(new_n13098_), .ZN(new_n13227_));
  NOR2_X1    g12915(.A1(new_n13225_), .A2(new_n13227_), .ZN(new_n13228_));
  INV_X1     g12916(.I(new_n13228_), .ZN(new_n13229_));
  NAND2_X1   g12917(.A1(new_n13225_), .A2(new_n13227_), .ZN(new_n13230_));
  AOI21_X1   g12918(.A1(new_n13229_), .A2(new_n13230_), .B(new_n13223_), .ZN(new_n13231_));
  XNOR2_X1   g12919(.A1(new_n13225_), .A2(new_n13227_), .ZN(new_n13232_));
  INV_X1     g12920(.I(new_n13232_), .ZN(new_n13233_));
  AOI21_X1   g12921(.A1(new_n13233_), .A2(new_n13223_), .B(new_n13231_), .ZN(new_n13234_));
  NOR2_X1    g12922(.A1(new_n13207_), .A2(new_n13234_), .ZN(new_n13235_));
  INV_X1     g12923(.I(new_n13235_), .ZN(new_n13236_));
  NAND2_X1   g12924(.A1(new_n13207_), .A2(new_n13234_), .ZN(new_n13237_));
  AOI21_X1   g12925(.A1(new_n13236_), .A2(new_n13237_), .B(new_n13147_), .ZN(new_n13238_));
  XNOR2_X1   g12926(.A1(new_n13207_), .A2(new_n13234_), .ZN(new_n13239_));
  INV_X1     g12927(.I(new_n13239_), .ZN(new_n13240_));
  AOI21_X1   g12928(.A1(new_n13240_), .A2(new_n13147_), .B(new_n13238_), .ZN(new_n13241_));
  NAND2_X1   g12929(.A1(new_n13114_), .A2(new_n13014_), .ZN(new_n13242_));
  NAND2_X1   g12930(.A1(new_n13242_), .A2(new_n13117_), .ZN(new_n13243_));
  OAI21_X1   g12931(.A1(new_n13016_), .A2(new_n13038_), .B(new_n13040_), .ZN(new_n13244_));
  NOR2_X1    g12932(.A1(new_n13111_), .A2(new_n13042_), .ZN(new_n13245_));
  NOR2_X1    g12933(.A1(new_n13245_), .A2(new_n13109_), .ZN(new_n13246_));
  INV_X1     g12934(.I(new_n13246_), .ZN(new_n13247_));
  AOI21_X1   g12935(.A1(new_n13027_), .A2(new_n13031_), .B(new_n13029_), .ZN(new_n13248_));
  INV_X1     g12936(.I(new_n13248_), .ZN(new_n13249_));
  NOR4_X1    g12937(.A1(new_n1215_), .A2(new_n2655_), .A3(new_n6260_), .A4(new_n9029_), .ZN(new_n13250_));
  AOI21_X1   g12938(.A1(new_n2978_), .A2(new_n9784_), .B(new_n13250_), .ZN(new_n13251_));
  INV_X1     g12939(.I(new_n13251_), .ZN(new_n13252_));
  NOR2_X1    g12940(.A1(new_n2655_), .A2(new_n6260_), .ZN(new_n13253_));
  NOR2_X1    g12941(.A1(new_n1313_), .A2(new_n8453_), .ZN(new_n13254_));
  XNOR2_X1   g12942(.A1(new_n13253_), .A2(new_n13254_), .ZN(new_n13255_));
  OAI21_X1   g12943(.A1(new_n13253_), .A2(new_n13255_), .B(new_n13252_), .ZN(new_n13256_));
  OAI21_X1   g12944(.A1(new_n1215_), .A2(new_n9029_), .B(new_n13255_), .ZN(new_n13257_));
  NAND2_X1   g12945(.A1(new_n13256_), .A2(new_n13257_), .ZN(new_n13258_));
  INV_X1     g12946(.I(new_n4369_), .ZN(new_n13259_));
  INV_X1     g12947(.I(new_n6056_), .ZN(new_n13260_));
  NOR2_X1    g12948(.A1(new_n13260_), .A2(new_n7512_), .ZN(new_n13261_));
  NOR2_X1    g12949(.A1(new_n13261_), .A2(new_n13259_), .ZN(new_n13262_));
  NOR4_X1    g12950(.A1(new_n4372_), .A2(new_n6028_), .A3(new_n2765_), .A4(new_n6055_), .ZN(new_n13263_));
  NAND2_X1   g12951(.A1(new_n13262_), .A2(new_n13263_), .ZN(new_n13264_));
  AOI22_X1   g12952(.A1(new_n2383_), .A2(new_n8996_), .B1(new_n9554_), .B2(new_n2286_), .ZN(new_n13265_));
  NOR4_X1    g12953(.A1(new_n8676_), .A2(new_n2543_), .A3(new_n1674_), .A4(new_n8990_), .ZN(new_n13266_));
  NAND2_X1   g12954(.A1(new_n13265_), .A2(new_n13266_), .ZN(new_n13267_));
  NOR2_X1    g12955(.A1(new_n13264_), .A2(new_n13267_), .ZN(new_n13268_));
  INV_X1     g12956(.I(new_n13267_), .ZN(new_n13269_));
  AOI21_X1   g12957(.A1(new_n13262_), .A2(new_n13263_), .B(new_n13269_), .ZN(new_n13270_));
  NOR2_X1    g12958(.A1(new_n13268_), .A2(new_n13270_), .ZN(new_n13271_));
  NOR2_X1    g12959(.A1(new_n13271_), .A2(new_n13258_), .ZN(new_n13272_));
  INV_X1     g12960(.I(new_n13258_), .ZN(new_n13273_));
  XOR2_X1    g12961(.A1(new_n13264_), .A2(new_n13269_), .Z(new_n13274_));
  NOR2_X1    g12962(.A1(new_n13274_), .A2(new_n13273_), .ZN(new_n13275_));
  NOR2_X1    g12963(.A1(new_n13275_), .A2(new_n13272_), .ZN(new_n13276_));
  NAND2_X1   g12964(.A1(new_n5339_), .A2(new_n5321_), .ZN(new_n13277_));
  NAND2_X1   g12965(.A1(\a[26] ), .A2(\a[56] ), .ZN(new_n13278_));
  XNOR2_X1   g12966(.A1(new_n13277_), .A2(new_n13278_), .ZN(new_n13279_));
  NOR2_X1    g12967(.A1(new_n3837_), .A2(new_n5511_), .ZN(new_n13280_));
  AOI22_X1   g12968(.A1(new_n5847_), .A2(new_n13280_), .B1(new_n3966_), .B2(new_n5980_), .ZN(new_n13281_));
  INV_X1     g12969(.I(new_n13281_), .ZN(new_n13282_));
  NOR4_X1    g12970(.A1(new_n3838_), .A2(new_n5488_), .A3(new_n3423_), .A4(new_n5511_), .ZN(new_n13283_));
  NAND2_X1   g12971(.A1(new_n13282_), .A2(new_n13283_), .ZN(new_n13284_));
  NAND2_X1   g12972(.A1(\a[52] ), .A2(\a[53] ), .ZN(new_n13285_));
  XOR2_X1    g12973(.A1(new_n2898_), .A2(new_n13285_), .Z(new_n13286_));
  NOR2_X1    g12974(.A1(new_n13284_), .A2(new_n13286_), .ZN(new_n13287_));
  INV_X1     g12975(.I(new_n13287_), .ZN(new_n13288_));
  NAND2_X1   g12976(.A1(new_n13284_), .A2(new_n13286_), .ZN(new_n13289_));
  AOI21_X1   g12977(.A1(new_n13288_), .A2(new_n13289_), .B(new_n13279_), .ZN(new_n13290_));
  INV_X1     g12978(.I(new_n13279_), .ZN(new_n13291_));
  XNOR2_X1   g12979(.A1(new_n13284_), .A2(new_n13286_), .ZN(new_n13292_));
  NOR2_X1    g12980(.A1(new_n13292_), .A2(new_n13291_), .ZN(new_n13293_));
  NOR2_X1    g12981(.A1(new_n13293_), .A2(new_n13290_), .ZN(new_n13294_));
  XOR2_X1    g12982(.A1(new_n13276_), .A2(new_n13294_), .Z(new_n13295_));
  NOR2_X1    g12983(.A1(new_n13276_), .A2(new_n13294_), .ZN(new_n13296_));
  INV_X1     g12984(.I(new_n13296_), .ZN(new_n13297_));
  NAND2_X1   g12985(.A1(new_n13276_), .A2(new_n13294_), .ZN(new_n13298_));
  AOI21_X1   g12986(.A1(new_n13297_), .A2(new_n13298_), .B(new_n13249_), .ZN(new_n13299_));
  AOI21_X1   g12987(.A1(new_n13249_), .A2(new_n13295_), .B(new_n13299_), .ZN(new_n13300_));
  NOR2_X1    g12988(.A1(new_n13247_), .A2(new_n13300_), .ZN(new_n13301_));
  NAND2_X1   g12989(.A1(new_n13247_), .A2(new_n13300_), .ZN(new_n13302_));
  INV_X1     g12990(.I(new_n13302_), .ZN(new_n13303_));
  OAI21_X1   g12991(.A1(new_n13303_), .A2(new_n13301_), .B(new_n13244_), .ZN(new_n13304_));
  XOR2_X1    g12992(.A1(new_n13246_), .A2(new_n13300_), .Z(new_n13305_));
  OAI21_X1   g12993(.A1(new_n13244_), .A2(new_n13305_), .B(new_n13304_), .ZN(new_n13306_));
  NAND2_X1   g12994(.A1(new_n13306_), .A2(new_n13243_), .ZN(new_n13307_));
  NOR2_X1    g12995(.A1(new_n13306_), .A2(new_n13243_), .ZN(new_n13308_));
  INV_X1     g12996(.I(new_n13308_), .ZN(new_n13309_));
  AOI21_X1   g12997(.A1(new_n13309_), .A2(new_n13307_), .B(new_n13241_), .ZN(new_n13310_));
  XOR2_X1    g12998(.A1(new_n13306_), .A2(new_n13243_), .Z(new_n13311_));
  AOI21_X1   g12999(.A1(new_n13241_), .A2(new_n13311_), .B(new_n13310_), .ZN(new_n13312_));
  AOI21_X1   g13000(.A1(new_n12883_), .A2(new_n13123_), .B(new_n13122_), .ZN(new_n13313_));
  XOR2_X1    g13001(.A1(new_n13312_), .A2(new_n13313_), .Z(new_n13314_));
  NAND2_X1   g13002(.A1(new_n13146_), .A2(new_n13314_), .ZN(new_n13315_));
  NOR2_X1    g13003(.A1(new_n13312_), .A2(new_n13313_), .ZN(new_n13316_));
  NAND2_X1   g13004(.A1(new_n13312_), .A2(new_n13313_), .ZN(new_n13317_));
  INV_X1     g13005(.I(new_n13317_), .ZN(new_n13318_));
  NOR2_X1    g13006(.A1(new_n13318_), .A2(new_n13316_), .ZN(new_n13319_));
  OAI21_X1   g13007(.A1(new_n13146_), .A2(new_n13319_), .B(new_n13315_), .ZN(\asquared[83] ));
  INV_X1     g13008(.I(new_n13127_), .ZN(new_n13321_));
  NOR2_X1    g13009(.A1(new_n13316_), .A2(new_n13138_), .ZN(new_n13322_));
  NAND2_X1   g13010(.A1(new_n13316_), .A2(new_n13138_), .ZN(new_n13323_));
  AOI21_X1   g13011(.A1(new_n13321_), .A2(new_n13323_), .B(new_n13322_), .ZN(new_n13324_));
  NAND2_X1   g13012(.A1(\asquared[81] ), .A2(new_n13324_), .ZN(new_n13325_));
  OAI21_X1   g13013(.A1(new_n13241_), .A2(new_n13308_), .B(new_n13307_), .ZN(new_n13326_));
  INV_X1     g13014(.I(new_n13326_), .ZN(new_n13327_));
  OAI21_X1   g13015(.A1(new_n13147_), .A2(new_n13235_), .B(new_n13237_), .ZN(new_n13328_));
  INV_X1     g13016(.I(new_n13301_), .ZN(new_n13329_));
  AOI21_X1   g13017(.A1(new_n13244_), .A2(new_n13329_), .B(new_n13303_), .ZN(new_n13330_));
  OAI21_X1   g13018(.A1(new_n13173_), .A2(new_n13174_), .B(new_n13175_), .ZN(new_n13331_));
  INV_X1     g13019(.I(new_n13331_), .ZN(new_n13332_));
  AOI21_X1   g13020(.A1(new_n13249_), .A2(new_n13298_), .B(new_n13296_), .ZN(new_n13333_));
  INV_X1     g13021(.I(new_n13333_), .ZN(new_n13334_));
  AOI21_X1   g13022(.A1(new_n13253_), .A2(new_n13254_), .B(new_n13252_), .ZN(new_n13335_));
  AOI21_X1   g13023(.A1(new_n4372_), .A2(new_n6028_), .B(new_n13262_), .ZN(new_n13336_));
  XNOR2_X1   g13024(.A1(new_n13336_), .A2(new_n13335_), .ZN(new_n13337_));
  NOR3_X1    g13025(.A1(new_n13337_), .A2(new_n13211_), .A3(new_n13213_), .ZN(new_n13338_));
  NOR2_X1    g13026(.A1(new_n13213_), .A2(new_n13211_), .ZN(new_n13339_));
  INV_X1     g13027(.I(new_n13335_), .ZN(new_n13340_));
  INV_X1     g13028(.I(new_n13336_), .ZN(new_n13341_));
  NOR2_X1    g13029(.A1(new_n13341_), .A2(new_n13340_), .ZN(new_n13342_));
  NOR2_X1    g13030(.A1(new_n13336_), .A2(new_n13335_), .ZN(new_n13343_));
  NOR2_X1    g13031(.A1(new_n13342_), .A2(new_n13343_), .ZN(new_n13344_));
  NOR2_X1    g13032(.A1(new_n13344_), .A2(new_n13339_), .ZN(new_n13345_));
  NOR2_X1    g13033(.A1(new_n13338_), .A2(new_n13345_), .ZN(new_n13346_));
  AOI21_X1   g13034(.A1(new_n2543_), .A2(new_n8676_), .B(new_n13265_), .ZN(new_n13347_));
  INV_X1     g13035(.I(new_n13347_), .ZN(new_n13348_));
  NAND2_X1   g13036(.A1(new_n5339_), .A2(new_n5321_), .ZN(new_n13349_));
  NOR2_X1    g13037(.A1(new_n5339_), .A2(new_n5321_), .ZN(new_n13350_));
  NOR2_X1    g13038(.A1(\a[26] ), .A2(\a[56] ), .ZN(new_n13351_));
  AOI21_X1   g13039(.A1(new_n13349_), .A2(new_n13351_), .B(new_n13350_), .ZN(new_n13352_));
  INV_X1     g13040(.I(new_n13352_), .ZN(new_n13353_));
  AOI21_X1   g13041(.A1(new_n3838_), .A2(new_n5488_), .B(new_n13282_), .ZN(new_n13354_));
  XOR2_X1    g13042(.A1(new_n13354_), .A2(new_n13353_), .Z(new_n13355_));
  NOR2_X1    g13043(.A1(new_n13355_), .A2(new_n13348_), .ZN(new_n13356_));
  INV_X1     g13044(.I(new_n13354_), .ZN(new_n13357_));
  NOR2_X1    g13045(.A1(new_n13357_), .A2(new_n13353_), .ZN(new_n13358_));
  NOR2_X1    g13046(.A1(new_n13354_), .A2(new_n13352_), .ZN(new_n13359_));
  NOR2_X1    g13047(.A1(new_n13358_), .A2(new_n13359_), .ZN(new_n13360_));
  NOR2_X1    g13048(.A1(new_n13360_), .A2(new_n13347_), .ZN(new_n13361_));
  AOI21_X1   g13049(.A1(new_n13291_), .A2(new_n13289_), .B(new_n13287_), .ZN(new_n13362_));
  NOR3_X1    g13050(.A1(new_n13361_), .A2(new_n13356_), .A3(new_n13362_), .ZN(new_n13363_));
  INV_X1     g13051(.I(new_n13363_), .ZN(new_n13364_));
  NOR2_X1    g13052(.A1(new_n13361_), .A2(new_n13356_), .ZN(new_n13365_));
  INV_X1     g13053(.I(new_n13362_), .ZN(new_n13366_));
  NOR2_X1    g13054(.A1(new_n13365_), .A2(new_n13366_), .ZN(new_n13367_));
  INV_X1     g13055(.I(new_n13367_), .ZN(new_n13368_));
  AOI21_X1   g13056(.A1(new_n13368_), .A2(new_n13364_), .B(new_n13346_), .ZN(new_n13369_));
  XOR2_X1    g13057(.A1(new_n13365_), .A2(new_n13362_), .Z(new_n13370_));
  INV_X1     g13058(.I(new_n13370_), .ZN(new_n13371_));
  AOI21_X1   g13059(.A1(new_n13346_), .A2(new_n13371_), .B(new_n13369_), .ZN(new_n13372_));
  NOR2_X1    g13060(.A1(new_n13372_), .A2(new_n13334_), .ZN(new_n13373_));
  INV_X1     g13061(.I(new_n13373_), .ZN(new_n13374_));
  NAND2_X1   g13062(.A1(new_n13372_), .A2(new_n13334_), .ZN(new_n13375_));
  AOI21_X1   g13063(.A1(new_n13374_), .A2(new_n13375_), .B(new_n13332_), .ZN(new_n13376_));
  XOR2_X1    g13064(.A1(new_n13372_), .A2(new_n13333_), .Z(new_n13377_));
  NOR2_X1    g13065(.A1(new_n13377_), .A2(new_n13331_), .ZN(new_n13378_));
  NOR2_X1    g13066(.A1(new_n13378_), .A2(new_n13376_), .ZN(new_n13379_));
  INV_X1     g13067(.I(new_n13379_), .ZN(new_n13380_));
  AOI21_X1   g13068(.A1(new_n13150_), .A2(new_n13158_), .B(new_n13156_), .ZN(new_n13381_));
  INV_X1     g13069(.I(new_n13168_), .ZN(new_n13382_));
  AOI21_X1   g13070(.A1(new_n13161_), .A2(new_n13382_), .B(new_n13167_), .ZN(new_n13383_));
  NOR2_X1    g13071(.A1(new_n13258_), .A2(new_n13270_), .ZN(new_n13384_));
  NOR2_X1    g13072(.A1(new_n13384_), .A2(new_n13268_), .ZN(new_n13385_));
  XNOR2_X1   g13073(.A1(new_n13383_), .A2(new_n13385_), .ZN(new_n13386_));
  NOR2_X1    g13074(.A1(new_n13386_), .A2(new_n13381_), .ZN(new_n13387_));
  INV_X1     g13075(.I(new_n13381_), .ZN(new_n13388_));
  NOR2_X1    g13076(.A1(new_n13383_), .A2(new_n13385_), .ZN(new_n13389_));
  INV_X1     g13077(.I(new_n13389_), .ZN(new_n13390_));
  NAND2_X1   g13078(.A1(new_n13383_), .A2(new_n13385_), .ZN(new_n13391_));
  AOI21_X1   g13079(.A1(new_n13390_), .A2(new_n13391_), .B(new_n13388_), .ZN(new_n13392_));
  NOR2_X1    g13080(.A1(new_n13387_), .A2(new_n13392_), .ZN(new_n13393_));
  OAI21_X1   g13081(.A1(new_n13180_), .A2(new_n13195_), .B(new_n13197_), .ZN(new_n13394_));
  NAND2_X1   g13082(.A1(\a[52] ), .A2(\a[53] ), .ZN(new_n13395_));
  NOR2_X1    g13083(.A1(new_n7486_), .A2(new_n3355_), .ZN(new_n13397_));
  AOI21_X1   g13084(.A1(new_n2898_), .A2(new_n12056_), .B(new_n7204_), .ZN(new_n13398_));
  NAND2_X1   g13085(.A1(\a[23] ), .A2(\a[59] ), .ZN(new_n13399_));
  NAND2_X1   g13086(.A1(\a[24] ), .A2(\a[60] ), .ZN(new_n13400_));
  XNOR2_X1   g13087(.A1(new_n13399_), .A2(new_n13400_), .ZN(new_n13401_));
  NOR2_X1    g13088(.A1(new_n13401_), .A2(new_n13398_), .ZN(new_n13402_));
  NAND2_X1   g13089(.A1(new_n13401_), .A2(new_n13398_), .ZN(new_n13403_));
  INV_X1     g13090(.I(new_n13403_), .ZN(new_n13404_));
  NOR2_X1    g13091(.A1(new_n13404_), .A2(new_n13402_), .ZN(new_n13405_));
  NAND2_X1   g13092(.A1(new_n13188_), .A2(new_n13189_), .ZN(new_n13406_));
  AOI21_X1   g13093(.A1(new_n12091_), .A2(new_n13406_), .B(new_n13190_), .ZN(new_n13407_));
  XOR2_X1    g13094(.A1(new_n13407_), .A2(new_n13405_), .Z(new_n13408_));
  NAND2_X1   g13095(.A1(new_n13408_), .A2(new_n13397_), .ZN(new_n13409_));
  INV_X1     g13096(.I(new_n13397_), .ZN(new_n13410_));
  NOR2_X1    g13097(.A1(new_n13407_), .A2(new_n13405_), .ZN(new_n13411_));
  NAND2_X1   g13098(.A1(new_n13407_), .A2(new_n13405_), .ZN(new_n13412_));
  INV_X1     g13099(.I(new_n13412_), .ZN(new_n13413_));
  OAI21_X1   g13100(.A1(new_n13413_), .A2(new_n13411_), .B(new_n13410_), .ZN(new_n13414_));
  AOI21_X1   g13101(.A1(new_n13409_), .A2(new_n13414_), .B(new_n13394_), .ZN(new_n13415_));
  INV_X1     g13102(.I(new_n13394_), .ZN(new_n13416_));
  NAND2_X1   g13103(.A1(new_n13409_), .A2(new_n13414_), .ZN(new_n13417_));
  NOR2_X1    g13104(.A1(new_n13416_), .A2(new_n13417_), .ZN(new_n13418_));
  NOR2_X1    g13105(.A1(new_n13418_), .A2(new_n13415_), .ZN(new_n13419_));
  XOR2_X1    g13106(.A1(new_n13394_), .A2(new_n13417_), .Z(new_n13420_));
  MUX2_X1    g13107(.I0(new_n13419_), .I1(new_n13420_), .S(new_n13393_), .Z(new_n13421_));
  NOR2_X1    g13108(.A1(new_n13380_), .A2(new_n13421_), .ZN(new_n13422_));
  INV_X1     g13109(.I(new_n13422_), .ZN(new_n13423_));
  NAND2_X1   g13110(.A1(new_n13380_), .A2(new_n13421_), .ZN(new_n13424_));
  AOI21_X1   g13111(.A1(new_n13423_), .A2(new_n13424_), .B(new_n13330_), .ZN(new_n13425_));
  XNOR2_X1   g13112(.A1(new_n13379_), .A2(new_n13421_), .ZN(new_n13426_));
  AOI21_X1   g13113(.A1(new_n13330_), .A2(new_n13426_), .B(new_n13425_), .ZN(new_n13427_));
  OAI21_X1   g13114(.A1(new_n13148_), .A2(new_n13203_), .B(new_n13205_), .ZN(new_n13428_));
  INV_X1     g13115(.I(new_n13428_), .ZN(new_n13429_));
  NAND2_X1   g13116(.A1(new_n13230_), .A2(new_n13223_), .ZN(new_n13430_));
  NAND2_X1   g13117(.A1(new_n13430_), .A2(new_n13229_), .ZN(new_n13431_));
  AOI21_X1   g13118(.A1(new_n13217_), .A2(new_n13221_), .B(new_n13219_), .ZN(new_n13432_));
  NAND2_X1   g13119(.A1(new_n5321_), .A2(new_n6024_), .ZN(new_n13433_));
  NAND2_X1   g13120(.A1(\a[29] ), .A2(\a[54] ), .ZN(new_n13434_));
  XNOR2_X1   g13121(.A1(new_n13433_), .A2(new_n13434_), .ZN(new_n13435_));
  INV_X1     g13122(.I(new_n13435_), .ZN(new_n13436_));
  AOI22_X1   g13123(.A1(new_n3424_), .A2(new_n6280_), .B1(new_n4372_), .B2(new_n6056_), .ZN(new_n13437_));
  NOR4_X1    g13124(.A1(new_n3487_), .A2(new_n6028_), .A3(new_n2868_), .A4(new_n6055_), .ZN(new_n13438_));
  NAND2_X1   g13125(.A1(new_n13437_), .A2(new_n13438_), .ZN(new_n13439_));
  XOR2_X1    g13126(.A1(new_n13186_), .A2(new_n10014_), .Z(new_n13440_));
  NOR2_X1    g13127(.A1(new_n13439_), .A2(new_n13440_), .ZN(new_n13441_));
  AND2_X2    g13128(.A1(new_n13439_), .A2(new_n13440_), .Z(new_n13442_));
  OAI21_X1   g13129(.A1(new_n13441_), .A2(new_n13442_), .B(new_n13436_), .ZN(new_n13443_));
  XNOR2_X1   g13130(.A1(new_n13439_), .A2(new_n13440_), .ZN(new_n13444_));
  OAI21_X1   g13131(.A1(new_n13436_), .A2(new_n13444_), .B(new_n13443_), .ZN(new_n13445_));
  NOR2_X1    g13132(.A1(new_n1999_), .A2(new_n7647_), .ZN(new_n13446_));
  NOR4_X1    g13133(.A1(new_n1999_), .A2(new_n2765_), .A3(new_n6260_), .A4(new_n7647_), .ZN(new_n13447_));
  AOI21_X1   g13134(.A1(new_n2752_), .A2(new_n8245_), .B(new_n13447_), .ZN(new_n13448_));
  INV_X1     g13135(.I(new_n13448_), .ZN(new_n13449_));
  NOR2_X1    g13136(.A1(new_n6260_), .A2(new_n7727_), .ZN(new_n13450_));
  INV_X1     g13137(.I(new_n13450_), .ZN(new_n13451_));
  NAND4_X1   g13138(.A1(new_n13449_), .A2(new_n3500_), .A3(new_n13446_), .A4(new_n13451_), .ZN(new_n13452_));
  INV_X1     g13139(.I(new_n13452_), .ZN(new_n13453_));
  AOI22_X1   g13140(.A1(new_n3838_), .A2(new_n5512_), .B1(new_n3805_), .B2(new_n5980_), .ZN(new_n13454_));
  NOR4_X1    g13141(.A1(new_n5488_), .A2(new_n5600_), .A3(new_n3393_), .A4(new_n5511_), .ZN(new_n13455_));
  NAND2_X1   g13142(.A1(new_n13454_), .A2(new_n13455_), .ZN(new_n13456_));
  XOR2_X1    g13143(.A1(new_n9781_), .A2(new_n1949_), .Z(new_n13457_));
  NOR2_X1    g13144(.A1(new_n13456_), .A2(new_n13457_), .ZN(new_n13458_));
  INV_X1     g13145(.I(new_n13456_), .ZN(new_n13459_));
  INV_X1     g13146(.I(new_n13457_), .ZN(new_n13460_));
  NOR2_X1    g13147(.A1(new_n13459_), .A2(new_n13460_), .ZN(new_n13461_));
  OAI21_X1   g13148(.A1(new_n13458_), .A2(new_n13461_), .B(new_n13453_), .ZN(new_n13462_));
  XNOR2_X1   g13149(.A1(new_n13456_), .A2(new_n13457_), .ZN(new_n13463_));
  OAI21_X1   g13150(.A1(new_n13453_), .A2(new_n13463_), .B(new_n13462_), .ZN(new_n13464_));
  XNOR2_X1   g13151(.A1(new_n13464_), .A2(new_n13445_), .ZN(new_n13465_));
  NOR2_X1    g13152(.A1(new_n13465_), .A2(new_n13432_), .ZN(new_n13466_));
  INV_X1     g13153(.I(new_n13432_), .ZN(new_n13467_));
  NAND2_X1   g13154(.A1(new_n13464_), .A2(new_n13445_), .ZN(new_n13468_));
  NOR2_X1    g13155(.A1(new_n13464_), .A2(new_n13445_), .ZN(new_n13469_));
  INV_X1     g13156(.I(new_n13469_), .ZN(new_n13470_));
  AOI21_X1   g13157(.A1(new_n13470_), .A2(new_n13468_), .B(new_n13467_), .ZN(new_n13471_));
  NOR2_X1    g13158(.A1(new_n13466_), .A2(new_n13471_), .ZN(new_n13472_));
  XNOR2_X1   g13159(.A1(new_n13431_), .A2(new_n13472_), .ZN(new_n13473_));
  NOR2_X1    g13160(.A1(new_n13431_), .A2(new_n13472_), .ZN(new_n13474_));
  NAND2_X1   g13161(.A1(new_n13431_), .A2(new_n13472_), .ZN(new_n13475_));
  INV_X1     g13162(.I(new_n13475_), .ZN(new_n13476_));
  OAI21_X1   g13163(.A1(new_n13474_), .A2(new_n13476_), .B(new_n13429_), .ZN(new_n13477_));
  OAI21_X1   g13164(.A1(new_n13473_), .A2(new_n13429_), .B(new_n13477_), .ZN(new_n13478_));
  NAND2_X1   g13165(.A1(new_n13427_), .A2(new_n13478_), .ZN(new_n13479_));
  NOR2_X1    g13166(.A1(new_n13427_), .A2(new_n13478_), .ZN(new_n13480_));
  INV_X1     g13167(.I(new_n13480_), .ZN(new_n13481_));
  NAND2_X1   g13168(.A1(new_n13481_), .A2(new_n13479_), .ZN(new_n13482_));
  XNOR2_X1   g13169(.A1(new_n13427_), .A2(new_n13478_), .ZN(new_n13483_));
  NOR2_X1    g13170(.A1(new_n13483_), .A2(new_n13328_), .ZN(new_n13484_));
  AOI21_X1   g13171(.A1(new_n13328_), .A2(new_n13482_), .B(new_n13484_), .ZN(new_n13485_));
  NOR2_X1    g13172(.A1(new_n13485_), .A2(new_n13327_), .ZN(new_n13486_));
  XOR2_X1    g13173(.A1(new_n13325_), .A2(new_n13486_), .Z(new_n13487_));
  XOR2_X1    g13174(.A1(new_n13487_), .A2(new_n13317_), .Z(\asquared[84] ));
  NOR2_X1    g13175(.A1(new_n13317_), .A2(new_n13327_), .ZN(new_n13489_));
  INV_X1     g13176(.I(new_n13489_), .ZN(new_n13490_));
  AOI21_X1   g13177(.A1(new_n13317_), .A2(new_n13327_), .B(new_n13485_), .ZN(new_n13491_));
  NAND4_X1   g13178(.A1(new_n12790_), .A2(new_n12782_), .A3(new_n13324_), .A4(new_n13491_), .ZN(new_n13492_));
  NAND2_X1   g13179(.A1(new_n13492_), .A2(new_n13490_), .ZN(new_n13493_));
  INV_X1     g13180(.I(new_n13493_), .ZN(new_n13494_));
  NAND2_X1   g13181(.A1(new_n13479_), .A2(new_n13328_), .ZN(new_n13495_));
  NAND2_X1   g13182(.A1(new_n13495_), .A2(new_n13481_), .ZN(new_n13496_));
  OAI21_X1   g13183(.A1(new_n13330_), .A2(new_n13422_), .B(new_n13424_), .ZN(new_n13497_));
  INV_X1     g13184(.I(new_n13497_), .ZN(new_n13498_));
  OAI21_X1   g13185(.A1(new_n13429_), .A2(new_n13474_), .B(new_n13475_), .ZN(new_n13499_));
  OAI21_X1   g13186(.A1(new_n13332_), .A2(new_n13373_), .B(new_n13375_), .ZN(new_n13500_));
  OAI21_X1   g13187(.A1(new_n13432_), .A2(new_n13469_), .B(new_n13468_), .ZN(new_n13501_));
  INV_X1     g13188(.I(new_n13501_), .ZN(new_n13502_));
  NAND2_X1   g13189(.A1(new_n13368_), .A2(new_n13346_), .ZN(new_n13503_));
  NAND2_X1   g13190(.A1(new_n13503_), .A2(new_n13364_), .ZN(new_n13504_));
  OAI22_X1   g13191(.A1(new_n7486_), .A2(new_n3355_), .B1(new_n3127_), .B2(new_n13395_), .ZN(new_n13505_));
  NOR2_X1    g13192(.A1(new_n5321_), .A2(new_n6024_), .ZN(new_n13506_));
  NAND2_X1   g13193(.A1(new_n2499_), .A2(new_n6945_), .ZN(new_n13507_));
  AOI21_X1   g13194(.A1(new_n6024_), .A2(new_n5321_), .B(new_n13507_), .ZN(new_n13508_));
  NOR2_X1    g13195(.A1(new_n13508_), .A2(new_n13506_), .ZN(new_n13509_));
  AOI21_X1   g13196(.A1(new_n5881_), .A2(new_n9029_), .B(new_n1313_), .ZN(new_n13510_));
  XNOR2_X1   g13197(.A1(new_n13509_), .A2(new_n13510_), .ZN(new_n13511_));
  NOR2_X1    g13198(.A1(new_n13511_), .A2(new_n13505_), .ZN(new_n13512_));
  INV_X1     g13199(.I(new_n13505_), .ZN(new_n13513_));
  INV_X1     g13200(.I(new_n13509_), .ZN(new_n13514_));
  INV_X1     g13201(.I(new_n13510_), .ZN(new_n13515_));
  NOR2_X1    g13202(.A1(new_n13514_), .A2(new_n13515_), .ZN(new_n13516_));
  NOR2_X1    g13203(.A1(new_n13509_), .A2(new_n13510_), .ZN(new_n13517_));
  NOR2_X1    g13204(.A1(new_n13516_), .A2(new_n13517_), .ZN(new_n13518_));
  NOR2_X1    g13205(.A1(new_n13518_), .A2(new_n13513_), .ZN(new_n13519_));
  NOR2_X1    g13206(.A1(new_n13519_), .A2(new_n13512_), .ZN(new_n13520_));
  INV_X1     g13207(.I(new_n13520_), .ZN(new_n13521_));
  INV_X1     g13208(.I(new_n13458_), .ZN(new_n13522_));
  OAI21_X1   g13209(.A1(new_n13459_), .A2(new_n13460_), .B(new_n13453_), .ZN(new_n13523_));
  NAND2_X1   g13210(.A1(new_n13523_), .A2(new_n13522_), .ZN(new_n13524_));
  INV_X1     g13211(.I(new_n13524_), .ZN(new_n13525_));
  NOR2_X1    g13212(.A1(new_n13442_), .A2(new_n13435_), .ZN(new_n13526_));
  NOR2_X1    g13213(.A1(new_n13526_), .A2(new_n13441_), .ZN(new_n13527_));
  NOR2_X1    g13214(.A1(new_n13525_), .A2(new_n13527_), .ZN(new_n13528_));
  NOR3_X1    g13215(.A1(new_n13524_), .A2(new_n13441_), .A3(new_n13526_), .ZN(new_n13529_));
  OAI21_X1   g13216(.A1(new_n13528_), .A2(new_n13529_), .B(new_n13521_), .ZN(new_n13530_));
  XOR2_X1    g13217(.A1(new_n13524_), .A2(new_n13527_), .Z(new_n13531_));
  OAI21_X1   g13218(.A1(new_n13521_), .A2(new_n13531_), .B(new_n13530_), .ZN(new_n13532_));
  INV_X1     g13219(.I(new_n13532_), .ZN(new_n13533_));
  NOR2_X1    g13220(.A1(new_n13533_), .A2(new_n13504_), .ZN(new_n13534_));
  INV_X1     g13221(.I(new_n13534_), .ZN(new_n13535_));
  NAND2_X1   g13222(.A1(new_n13533_), .A2(new_n13504_), .ZN(new_n13536_));
  AOI21_X1   g13223(.A1(new_n13535_), .A2(new_n13536_), .B(new_n13502_), .ZN(new_n13537_));
  XOR2_X1    g13224(.A1(new_n13504_), .A2(new_n13532_), .Z(new_n13538_));
  NOR2_X1    g13225(.A1(new_n13538_), .A2(new_n13501_), .ZN(new_n13539_));
  NOR2_X1    g13226(.A1(new_n13539_), .A2(new_n13537_), .ZN(new_n13540_));
  XOR2_X1    g13227(.A1(new_n13540_), .A2(new_n13500_), .Z(new_n13541_));
  INV_X1     g13228(.I(new_n13541_), .ZN(new_n13542_));
  INV_X1     g13229(.I(new_n13500_), .ZN(new_n13543_));
  NOR2_X1    g13230(.A1(new_n13540_), .A2(new_n13543_), .ZN(new_n13544_));
  INV_X1     g13231(.I(new_n13544_), .ZN(new_n13545_));
  NAND2_X1   g13232(.A1(new_n13540_), .A2(new_n13543_), .ZN(new_n13546_));
  AOI21_X1   g13233(.A1(new_n13545_), .A2(new_n13546_), .B(new_n13499_), .ZN(new_n13547_));
  AOI21_X1   g13234(.A1(new_n13542_), .A2(new_n13499_), .B(new_n13547_), .ZN(new_n13548_));
  AOI21_X1   g13235(.A1(new_n13388_), .A2(new_n13391_), .B(new_n13389_), .ZN(new_n13549_));
  AOI21_X1   g13236(.A1(new_n13397_), .A2(new_n13412_), .B(new_n13411_), .ZN(new_n13550_));
  NAND2_X1   g13237(.A1(new_n8996_), .A2(new_n2543_), .ZN(new_n13551_));
  OAI21_X1   g13238(.A1(new_n1949_), .A2(new_n12632_), .B(new_n9861_), .ZN(new_n13552_));
  NOR2_X1    g13239(.A1(new_n1916_), .A2(new_n7647_), .ZN(new_n13553_));
  XNOR2_X1   g13240(.A1(new_n3981_), .A2(new_n7204_), .ZN(new_n13554_));
  INV_X1     g13241(.I(new_n13554_), .ZN(new_n13555_));
  NAND2_X1   g13242(.A1(new_n13555_), .A2(new_n13552_), .ZN(new_n13556_));
  XOR2_X1    g13243(.A1(new_n13556_), .A2(new_n13404_), .Z(new_n13557_));
  XNOR2_X1   g13244(.A1(new_n13557_), .A2(new_n13551_), .ZN(new_n13558_));
  XNOR2_X1   g13245(.A1(new_n13558_), .A2(new_n13550_), .ZN(new_n13559_));
  NOR2_X1    g13246(.A1(new_n13559_), .A2(new_n13549_), .ZN(new_n13560_));
  INV_X1     g13247(.I(new_n13549_), .ZN(new_n13561_));
  NOR2_X1    g13248(.A1(new_n13558_), .A2(new_n13550_), .ZN(new_n13562_));
  INV_X1     g13249(.I(new_n13562_), .ZN(new_n13563_));
  NAND2_X1   g13250(.A1(new_n13558_), .A2(new_n13550_), .ZN(new_n13564_));
  AOI21_X1   g13251(.A1(new_n13563_), .A2(new_n13564_), .B(new_n13561_), .ZN(new_n13565_));
  NOR2_X1    g13252(.A1(new_n13565_), .A2(new_n13560_), .ZN(new_n13566_));
  INV_X1     g13253(.I(new_n13415_), .ZN(new_n13567_));
  AOI21_X1   g13254(.A1(new_n13393_), .A2(new_n13567_), .B(new_n13418_), .ZN(new_n13568_));
  INV_X1     g13255(.I(new_n13343_), .ZN(new_n13569_));
  AOI21_X1   g13256(.A1(new_n13339_), .A2(new_n13569_), .B(new_n13342_), .ZN(new_n13570_));
  AOI21_X1   g13257(.A1(new_n3487_), .A2(new_n6028_), .B(new_n13437_), .ZN(new_n13571_));
  INV_X1     g13258(.I(new_n13571_), .ZN(new_n13572_));
  OAI21_X1   g13259(.A1(new_n3500_), .A2(new_n13451_), .B(new_n13448_), .ZN(new_n13573_));
  AOI21_X1   g13260(.A1(new_n5600_), .A2(new_n5488_), .B(new_n13454_), .ZN(new_n13574_));
  XOR2_X1    g13261(.A1(new_n13573_), .A2(new_n13574_), .Z(new_n13575_));
  NOR2_X1    g13262(.A1(new_n13575_), .A2(new_n13572_), .ZN(new_n13576_));
  INV_X1     g13263(.I(new_n13574_), .ZN(new_n13577_));
  NOR2_X1    g13264(.A1(new_n13577_), .A2(new_n13573_), .ZN(new_n13578_));
  INV_X1     g13265(.I(new_n13578_), .ZN(new_n13579_));
  NAND2_X1   g13266(.A1(new_n13577_), .A2(new_n13573_), .ZN(new_n13580_));
  AOI21_X1   g13267(.A1(new_n13579_), .A2(new_n13580_), .B(new_n13571_), .ZN(new_n13581_));
  NOR2_X1    g13268(.A1(new_n13576_), .A2(new_n13581_), .ZN(new_n13582_));
  NOR2_X1    g13269(.A1(new_n13359_), .A2(new_n13348_), .ZN(new_n13583_));
  NOR2_X1    g13270(.A1(new_n13583_), .A2(new_n13358_), .ZN(new_n13584_));
  XOR2_X1    g13271(.A1(new_n13582_), .A2(new_n13584_), .Z(new_n13585_));
  NOR2_X1    g13272(.A1(new_n13585_), .A2(new_n13570_), .ZN(new_n13586_));
  INV_X1     g13273(.I(new_n13570_), .ZN(new_n13587_));
  INV_X1     g13274(.I(new_n13582_), .ZN(new_n13588_));
  NOR2_X1    g13275(.A1(new_n13588_), .A2(new_n13584_), .ZN(new_n13589_));
  INV_X1     g13276(.I(new_n13589_), .ZN(new_n13590_));
  NAND2_X1   g13277(.A1(new_n13588_), .A2(new_n13584_), .ZN(new_n13591_));
  AOI21_X1   g13278(.A1(new_n13590_), .A2(new_n13591_), .B(new_n13587_), .ZN(new_n13592_));
  NOR2_X1    g13279(.A1(new_n13592_), .A2(new_n13586_), .ZN(new_n13593_));
  INV_X1     g13280(.I(new_n13593_), .ZN(new_n13594_));
  NOR2_X1    g13281(.A1(new_n3804_), .A2(new_n7216_), .ZN(new_n13595_));
  NAND3_X1   g13282(.A1(new_n13595_), .A2(\a[28] ), .A3(\a[46] ), .ZN(new_n13596_));
  OAI21_X1   g13283(.A1(new_n2689_), .A2(new_n8953_), .B(new_n13596_), .ZN(new_n13597_));
  NOR2_X1    g13284(.A1(new_n2499_), .A2(new_n6999_), .ZN(new_n13598_));
  NOR2_X1    g13285(.A1(new_n3804_), .A2(new_n5175_), .ZN(new_n13599_));
  XNOR2_X1   g13286(.A1(new_n13598_), .A2(new_n13599_), .ZN(new_n13600_));
  OAI21_X1   g13287(.A1(new_n2499_), .A2(new_n6999_), .B(new_n13599_), .ZN(new_n13601_));
  NAND2_X1   g13288(.A1(\a[28] ), .A2(\a[56] ), .ZN(new_n13602_));
  AOI22_X1   g13289(.A1(new_n13600_), .A2(new_n13602_), .B1(new_n13597_), .B2(new_n13601_), .ZN(new_n13603_));
  INV_X1     g13290(.I(new_n13603_), .ZN(new_n13604_));
  AOI22_X1   g13291(.A1(new_n4415_), .A2(new_n5742_), .B1(new_n7186_), .B2(new_n6024_), .ZN(new_n13605_));
  NOR2_X1    g13292(.A1(new_n5322_), .A2(new_n6579_), .ZN(new_n13606_));
  NOR2_X1    g13293(.A1(new_n5003_), .A2(new_n6772_), .ZN(new_n13607_));
  NOR4_X1    g13294(.A1(new_n13606_), .A2(new_n3783_), .A3(new_n5004_), .A4(new_n13607_), .ZN(new_n13608_));
  NAND2_X1   g13295(.A1(new_n13608_), .A2(new_n13605_), .ZN(new_n13609_));
  NAND4_X1   g13296(.A1(\a[27] ), .A2(\a[30] ), .A3(\a[54] ), .A4(\a[57] ), .ZN(new_n13610_));
  XOR2_X1    g13297(.A1(new_n13280_), .A2(new_n13610_), .Z(new_n13611_));
  NOR2_X1    g13298(.A1(new_n13609_), .A2(new_n13611_), .ZN(new_n13612_));
  INV_X1     g13299(.I(new_n13611_), .ZN(new_n13613_));
  AOI21_X1   g13300(.A1(new_n13605_), .A2(new_n13608_), .B(new_n13613_), .ZN(new_n13614_));
  NOR2_X1    g13301(.A1(new_n13612_), .A2(new_n13614_), .ZN(new_n13615_));
  NOR2_X1    g13302(.A1(new_n13615_), .A2(new_n13604_), .ZN(new_n13616_));
  XOR2_X1    g13303(.A1(new_n13609_), .A2(new_n13613_), .Z(new_n13617_));
  NOR2_X1    g13304(.A1(new_n13617_), .A2(new_n13603_), .ZN(new_n13618_));
  NOR2_X1    g13305(.A1(new_n13618_), .A2(new_n13616_), .ZN(new_n13619_));
  NOR2_X1    g13306(.A1(new_n9550_), .A2(new_n9861_), .ZN(new_n13620_));
  NOR2_X1    g13307(.A1(new_n13620_), .A2(new_n6195_), .ZN(new_n13621_));
  NOR2_X1    g13308(.A1(new_n1313_), .A2(new_n9310_), .ZN(new_n13622_));
  NAND4_X1   g13309(.A1(new_n13621_), .A2(new_n2285_), .A3(new_n9785_), .A4(new_n13622_), .ZN(new_n13623_));
  NAND2_X1   g13310(.A1(new_n8996_), .A2(new_n2277_), .ZN(new_n13624_));
  NOR2_X1    g13311(.A1(new_n2868_), .A2(new_n6260_), .ZN(new_n13625_));
  XOR2_X1    g13312(.A1(new_n13624_), .A2(new_n13625_), .Z(new_n13626_));
  AOI21_X1   g13313(.A1(new_n3487_), .A2(new_n4727_), .B(new_n13261_), .ZN(new_n13627_));
  NOR4_X1    g13314(.A1(new_n3966_), .A2(new_n6028_), .A3(new_n3371_), .A4(new_n6055_), .ZN(new_n13628_));
  NAND2_X1   g13315(.A1(new_n13627_), .A2(new_n13628_), .ZN(new_n13629_));
  NOR2_X1    g13316(.A1(new_n13629_), .A2(new_n13626_), .ZN(new_n13630_));
  INV_X1     g13317(.I(new_n13630_), .ZN(new_n13631_));
  NAND2_X1   g13318(.A1(new_n13629_), .A2(new_n13626_), .ZN(new_n13632_));
  AOI21_X1   g13319(.A1(new_n13631_), .A2(new_n13632_), .B(new_n13623_), .ZN(new_n13633_));
  INV_X1     g13320(.I(new_n13623_), .ZN(new_n13634_));
  XNOR2_X1   g13321(.A1(new_n13629_), .A2(new_n13626_), .ZN(new_n13635_));
  NOR2_X1    g13322(.A1(new_n13635_), .A2(new_n13634_), .ZN(new_n13636_));
  NOR2_X1    g13323(.A1(new_n13636_), .A2(new_n13633_), .ZN(new_n13637_));
  XOR2_X1    g13324(.A1(new_n13637_), .A2(new_n13619_), .Z(new_n13638_));
  NAND2_X1   g13325(.A1(new_n13594_), .A2(new_n13638_), .ZN(new_n13639_));
  NOR2_X1    g13326(.A1(new_n13637_), .A2(new_n13619_), .ZN(new_n13640_));
  NOR4_X1    g13327(.A1(new_n13636_), .A2(new_n13618_), .A3(new_n13616_), .A4(new_n13633_), .ZN(new_n13641_));
  OAI21_X1   g13328(.A1(new_n13640_), .A2(new_n13641_), .B(new_n13593_), .ZN(new_n13642_));
  NAND2_X1   g13329(.A1(new_n13639_), .A2(new_n13642_), .ZN(new_n13643_));
  INV_X1     g13330(.I(new_n13643_), .ZN(new_n13644_));
  NOR2_X1    g13331(.A1(new_n13644_), .A2(new_n13568_), .ZN(new_n13645_));
  INV_X1     g13332(.I(new_n13645_), .ZN(new_n13646_));
  NAND2_X1   g13333(.A1(new_n13644_), .A2(new_n13568_), .ZN(new_n13647_));
  AOI21_X1   g13334(.A1(new_n13646_), .A2(new_n13647_), .B(new_n13566_), .ZN(new_n13648_));
  XOR2_X1    g13335(.A1(new_n13643_), .A2(new_n13568_), .Z(new_n13649_));
  INV_X1     g13336(.I(new_n13649_), .ZN(new_n13650_));
  AOI21_X1   g13337(.A1(new_n13566_), .A2(new_n13650_), .B(new_n13648_), .ZN(new_n13651_));
  NOR2_X1    g13338(.A1(new_n13548_), .A2(new_n13651_), .ZN(new_n13652_));
  INV_X1     g13339(.I(new_n13652_), .ZN(new_n13653_));
  NAND2_X1   g13340(.A1(new_n13548_), .A2(new_n13651_), .ZN(new_n13654_));
  AOI21_X1   g13341(.A1(new_n13653_), .A2(new_n13654_), .B(new_n13498_), .ZN(new_n13655_));
  XNOR2_X1   g13342(.A1(new_n13548_), .A2(new_n13651_), .ZN(new_n13656_));
  NOR2_X1    g13343(.A1(new_n13656_), .A2(new_n13497_), .ZN(new_n13657_));
  NOR2_X1    g13344(.A1(new_n13657_), .A2(new_n13655_), .ZN(new_n13658_));
  XOR2_X1    g13345(.A1(new_n13496_), .A2(new_n13658_), .Z(new_n13659_));
  OAI21_X1   g13346(.A1(new_n13655_), .A2(new_n13657_), .B(new_n13496_), .ZN(new_n13660_));
  INV_X1     g13347(.I(new_n13496_), .ZN(new_n13661_));
  NAND2_X1   g13348(.A1(new_n13661_), .A2(new_n13658_), .ZN(new_n13662_));
  NAND2_X1   g13349(.A1(new_n13662_), .A2(new_n13660_), .ZN(new_n13663_));
  NAND2_X1   g13350(.A1(new_n13494_), .A2(new_n13663_), .ZN(new_n13664_));
  OAI21_X1   g13351(.A1(new_n13494_), .A2(new_n13659_), .B(new_n13664_), .ZN(\asquared[85] ));
  NAND2_X1   g13352(.A1(new_n13493_), .A2(new_n13662_), .ZN(new_n13666_));
  NAND2_X1   g13353(.A1(new_n13666_), .A2(new_n13660_), .ZN(new_n13667_));
  OAI21_X1   g13354(.A1(new_n13498_), .A2(new_n13652_), .B(new_n13654_), .ZN(new_n13668_));
  AOI21_X1   g13355(.A1(new_n13499_), .A2(new_n13546_), .B(new_n13544_), .ZN(new_n13669_));
  OAI21_X1   g13356(.A1(new_n13502_), .A2(new_n13534_), .B(new_n13536_), .ZN(new_n13670_));
  AOI21_X1   g13357(.A1(new_n13561_), .A2(new_n13564_), .B(new_n13562_), .ZN(new_n13671_));
  NOR2_X1    g13358(.A1(new_n13594_), .A2(new_n13641_), .ZN(new_n13672_));
  NOR2_X1    g13359(.A1(new_n13672_), .A2(new_n13640_), .ZN(new_n13673_));
  NOR2_X1    g13360(.A1(new_n13517_), .A2(new_n13505_), .ZN(new_n13674_));
  NOR2_X1    g13361(.A1(new_n13674_), .A2(new_n13516_), .ZN(new_n13675_));
  NAND2_X1   g13362(.A1(new_n13580_), .A2(new_n13571_), .ZN(new_n13676_));
  NAND2_X1   g13363(.A1(new_n13676_), .A2(new_n13579_), .ZN(new_n13677_));
  NAND2_X1   g13364(.A1(new_n13404_), .A2(new_n13552_), .ZN(new_n13678_));
  NOR2_X1    g13365(.A1(new_n13554_), .A2(new_n13551_), .ZN(new_n13679_));
  OAI21_X1   g13366(.A1(new_n13404_), .A2(new_n13552_), .B(new_n13679_), .ZN(new_n13680_));
  NAND2_X1   g13367(.A1(new_n13680_), .A2(new_n13678_), .ZN(new_n13681_));
  XNOR2_X1   g13368(.A1(new_n13677_), .A2(new_n13681_), .ZN(new_n13682_));
  AOI22_X1   g13369(.A1(new_n13676_), .A2(new_n13579_), .B1(new_n13678_), .B2(new_n13680_), .ZN(new_n13683_));
  NOR2_X1    g13370(.A1(new_n13677_), .A2(new_n13681_), .ZN(new_n13684_));
  OAI21_X1   g13371(.A1(new_n13684_), .A2(new_n13683_), .B(new_n13675_), .ZN(new_n13685_));
  OAI21_X1   g13372(.A1(new_n13682_), .A2(new_n13675_), .B(new_n13685_), .ZN(new_n13686_));
  XNOR2_X1   g13373(.A1(new_n13673_), .A2(new_n13686_), .ZN(new_n13687_));
  NAND2_X1   g13374(.A1(new_n13673_), .A2(new_n13686_), .ZN(new_n13688_));
  NOR2_X1    g13375(.A1(new_n13673_), .A2(new_n13686_), .ZN(new_n13689_));
  INV_X1     g13376(.I(new_n13689_), .ZN(new_n13690_));
  NAND2_X1   g13377(.A1(new_n13690_), .A2(new_n13688_), .ZN(new_n13691_));
  NAND2_X1   g13378(.A1(new_n13691_), .A2(new_n13671_), .ZN(new_n13692_));
  OAI21_X1   g13379(.A1(new_n13671_), .A2(new_n13687_), .B(new_n13692_), .ZN(new_n13693_));
  AOI21_X1   g13380(.A1(new_n13566_), .A2(new_n13647_), .B(new_n13645_), .ZN(new_n13694_));
  XOR2_X1    g13381(.A1(new_n13693_), .A2(new_n13694_), .Z(new_n13695_));
  NOR2_X1    g13382(.A1(new_n13693_), .A2(new_n13694_), .ZN(new_n13696_));
  INV_X1     g13383(.I(new_n13696_), .ZN(new_n13697_));
  NAND2_X1   g13384(.A1(new_n13693_), .A2(new_n13694_), .ZN(new_n13698_));
  AOI21_X1   g13385(.A1(new_n13697_), .A2(new_n13698_), .B(new_n13670_), .ZN(new_n13699_));
  AOI21_X1   g13386(.A1(new_n13670_), .A2(new_n13695_), .B(new_n13699_), .ZN(new_n13700_));
  INV_X1     g13387(.I(new_n13528_), .ZN(new_n13701_));
  OAI21_X1   g13388(.A1(new_n13521_), .A2(new_n13529_), .B(new_n13701_), .ZN(new_n13702_));
  NOR2_X1    g13389(.A1(new_n7001_), .A2(new_n8056_), .ZN(new_n13703_));
  NOR2_X1    g13390(.A1(new_n13703_), .A2(new_n13259_), .ZN(new_n13704_));
  NOR2_X1    g13391(.A1(new_n2765_), .A2(new_n6694_), .ZN(new_n13705_));
  NAND4_X1   g13392(.A1(new_n13704_), .A2(new_n4644_), .A3(new_n10034_), .A4(new_n13705_), .ZN(new_n13706_));
  NOR2_X1    g13393(.A1(new_n6146_), .A2(new_n4321_), .ZN(new_n13707_));
  NOR2_X1    g13394(.A1(new_n10533_), .A2(new_n13707_), .ZN(new_n13708_));
  NOR2_X1    g13395(.A1(new_n3783_), .A2(new_n5175_), .ZN(new_n13709_));
  NAND4_X1   g13396(.A1(new_n13708_), .A2(new_n6579_), .A3(new_n5743_), .A4(new_n13709_), .ZN(new_n13710_));
  NOR2_X1    g13397(.A1(new_n2178_), .A2(new_n7727_), .ZN(new_n13711_));
  NOR2_X1    g13398(.A1(new_n3423_), .A2(new_n6055_), .ZN(new_n13712_));
  NAND2_X1   g13399(.A1(new_n13711_), .A2(new_n13712_), .ZN(new_n13713_));
  XOR2_X1    g13400(.A1(new_n13713_), .A2(\a[22] ), .Z(new_n13714_));
  XOR2_X1    g13401(.A1(new_n13714_), .A2(\a[63] ), .Z(new_n13715_));
  NOR2_X1    g13402(.A1(new_n13715_), .A2(new_n13710_), .ZN(new_n13716_));
  AND2_X2    g13403(.A1(new_n13715_), .A2(new_n13710_), .Z(new_n13717_));
  NOR2_X1    g13404(.A1(new_n13717_), .A2(new_n13716_), .ZN(new_n13718_));
  NOR2_X1    g13405(.A1(new_n13718_), .A2(new_n13706_), .ZN(new_n13719_));
  INV_X1     g13406(.I(new_n13706_), .ZN(new_n13720_));
  XNOR2_X1   g13407(.A1(new_n13715_), .A2(new_n13710_), .ZN(new_n13721_));
  NOR2_X1    g13408(.A1(new_n13721_), .A2(new_n13720_), .ZN(new_n13722_));
  NOR2_X1    g13409(.A1(new_n13719_), .A2(new_n13722_), .ZN(new_n13723_));
  AOI22_X1   g13410(.A1(new_n3805_), .A2(new_n6028_), .B1(new_n3838_), .B2(new_n6027_), .ZN(new_n13724_));
  NAND4_X1   g13411(.A1(new_n13724_), .A2(new_n4706_), .A3(new_n7693_), .A4(new_n6740_), .ZN(new_n13725_));
  INV_X1     g13412(.I(new_n13725_), .ZN(new_n13726_));
  NOR2_X1    g13413(.A1(new_n12160_), .A2(new_n10761_), .ZN(new_n13727_));
  INV_X1     g13414(.I(new_n13727_), .ZN(new_n13728_));
  NAND3_X1   g13415(.A1(new_n8005_), .A2(new_n3127_), .A3(new_n7588_), .ZN(new_n13729_));
  NAND2_X1   g13416(.A1(\a[42] ), .A2(\a[62] ), .ZN(new_n13730_));
  XNOR2_X1   g13417(.A1(new_n9797_), .A2(new_n13730_), .ZN(new_n13731_));
  NOR3_X1    g13418(.A1(new_n13728_), .A2(new_n13729_), .A3(new_n13731_), .ZN(new_n13732_));
  NOR2_X1    g13419(.A1(new_n13728_), .A2(new_n13729_), .ZN(new_n13733_));
  INV_X1     g13420(.I(new_n13731_), .ZN(new_n13734_));
  NOR2_X1    g13421(.A1(new_n13733_), .A2(new_n13734_), .ZN(new_n13735_));
  OAI21_X1   g13422(.A1(new_n13735_), .A2(new_n13732_), .B(new_n13726_), .ZN(new_n13736_));
  XOR2_X1    g13423(.A1(new_n13733_), .A2(new_n13734_), .Z(new_n13737_));
  NAND2_X1   g13424(.A1(new_n13737_), .A2(new_n13725_), .ZN(new_n13738_));
  NAND2_X1   g13425(.A1(new_n13738_), .A2(new_n13736_), .ZN(new_n13739_));
  INV_X1     g13426(.I(new_n13739_), .ZN(new_n13740_));
  XOR2_X1    g13427(.A1(new_n13723_), .A2(new_n13740_), .Z(new_n13741_));
  OAI21_X1   g13428(.A1(new_n13719_), .A2(new_n13722_), .B(new_n13739_), .ZN(new_n13742_));
  NAND2_X1   g13429(.A1(new_n13723_), .A2(new_n13740_), .ZN(new_n13743_));
  AOI21_X1   g13430(.A1(new_n13743_), .A2(new_n13742_), .B(new_n13702_), .ZN(new_n13744_));
  AOI21_X1   g13431(.A1(new_n13741_), .A2(new_n13702_), .B(new_n13744_), .ZN(new_n13745_));
  NAND2_X1   g13432(.A1(new_n13591_), .A2(new_n13587_), .ZN(new_n13746_));
  AOI21_X1   g13433(.A1(new_n13598_), .A2(new_n13599_), .B(new_n13597_), .ZN(new_n13747_));
  INV_X1     g13434(.I(new_n13747_), .ZN(new_n13748_));
  NOR2_X1    g13435(.A1(new_n13606_), .A2(new_n13605_), .ZN(new_n13749_));
  INV_X1     g13436(.I(new_n13749_), .ZN(new_n13750_));
  NOR2_X1    g13437(.A1(new_n13748_), .A2(new_n13750_), .ZN(new_n13751_));
  XOR2_X1    g13438(.A1(new_n13751_), .A2(new_n1691_), .Z(new_n13752_));
  XOR2_X1    g13439(.A1(new_n13752_), .A2(\a[61] ), .Z(new_n13753_));
  INV_X1     g13440(.I(new_n13753_), .ZN(new_n13754_));
  NAND3_X1   g13441(.A1(new_n13023_), .A2(\a[30] ), .A3(\a[57] ), .ZN(new_n13755_));
  NOR2_X1    g13442(.A1(\a[37] ), .A2(\a[47] ), .ZN(new_n13756_));
  AOI22_X1   g13443(.A1(new_n13755_), .A2(new_n13756_), .B1(new_n12965_), .B2(new_n7470_), .ZN(new_n13757_));
  AOI22_X1   g13444(.A1(new_n2752_), .A2(new_n9554_), .B1(new_n2890_), .B2(new_n8996_), .ZN(new_n13758_));
  NOR4_X1    g13445(.A1(new_n2533_), .A2(new_n8676_), .A3(new_n1999_), .A4(new_n8990_), .ZN(new_n13759_));
  NAND2_X1   g13446(.A1(new_n13758_), .A2(new_n13759_), .ZN(new_n13760_));
  AOI21_X1   g13447(.A1(new_n3981_), .A2(new_n13553_), .B(new_n7204_), .ZN(new_n13761_));
  NOR2_X1    g13448(.A1(new_n13760_), .A2(new_n13761_), .ZN(new_n13762_));
  INV_X1     g13449(.I(new_n13762_), .ZN(new_n13763_));
  NAND2_X1   g13450(.A1(new_n13760_), .A2(new_n13761_), .ZN(new_n13764_));
  NAND2_X1   g13451(.A1(new_n13763_), .A2(new_n13764_), .ZN(new_n13765_));
  XNOR2_X1   g13452(.A1(new_n13760_), .A2(new_n13761_), .ZN(new_n13766_));
  NOR2_X1    g13453(.A1(new_n13766_), .A2(new_n13757_), .ZN(new_n13767_));
  AOI21_X1   g13454(.A1(new_n13757_), .A2(new_n13765_), .B(new_n13767_), .ZN(new_n13768_));
  NOR2_X1    g13455(.A1(new_n13754_), .A2(new_n13768_), .ZN(new_n13769_));
  INV_X1     g13456(.I(new_n13769_), .ZN(new_n13770_));
  NAND2_X1   g13457(.A1(new_n13754_), .A2(new_n13768_), .ZN(new_n13771_));
  AOI22_X1   g13458(.A1(new_n13770_), .A2(new_n13771_), .B1(new_n13590_), .B2(new_n13746_), .ZN(new_n13772_));
  NAND2_X1   g13459(.A1(new_n13746_), .A2(new_n13590_), .ZN(new_n13773_));
  XOR2_X1    g13460(.A1(new_n13753_), .A2(new_n13768_), .Z(new_n13774_));
  NOR2_X1    g13461(.A1(new_n13774_), .A2(new_n13773_), .ZN(new_n13775_));
  NOR2_X1    g13462(.A1(new_n13772_), .A2(new_n13775_), .ZN(new_n13776_));
  INV_X1     g13463(.I(new_n13614_), .ZN(new_n13777_));
  AOI21_X1   g13464(.A1(new_n13777_), .A2(new_n13603_), .B(new_n13612_), .ZN(new_n13778_));
  INV_X1     g13465(.I(new_n13778_), .ZN(new_n13779_));
  AOI21_X1   g13466(.A1(new_n2286_), .A2(new_n9784_), .B(new_n13621_), .ZN(new_n13780_));
  NOR2_X1    g13467(.A1(new_n8996_), .A2(new_n2277_), .ZN(new_n13781_));
  NAND2_X1   g13468(.A1(new_n2868_), .A2(new_n6260_), .ZN(new_n13782_));
  AOI21_X1   g13469(.A1(new_n2277_), .A2(new_n8996_), .B(new_n13782_), .ZN(new_n13783_));
  NOR2_X1    g13470(.A1(new_n13783_), .A2(new_n13781_), .ZN(new_n13784_));
  AOI21_X1   g13471(.A1(new_n3966_), .A2(new_n6028_), .B(new_n13627_), .ZN(new_n13785_));
  XOR2_X1    g13472(.A1(new_n13785_), .A2(new_n13784_), .Z(new_n13786_));
  NAND2_X1   g13473(.A1(new_n13786_), .A2(new_n13780_), .ZN(new_n13787_));
  INV_X1     g13474(.I(new_n13780_), .ZN(new_n13788_));
  AND2_X2    g13475(.A1(new_n13785_), .A2(new_n13784_), .Z(new_n13789_));
  NOR2_X1    g13476(.A1(new_n13785_), .A2(new_n13784_), .ZN(new_n13790_));
  OAI21_X1   g13477(.A1(new_n13789_), .A2(new_n13790_), .B(new_n13788_), .ZN(new_n13791_));
  NAND2_X1   g13478(.A1(new_n13787_), .A2(new_n13791_), .ZN(new_n13792_));
  NAND2_X1   g13479(.A1(new_n13632_), .A2(new_n13634_), .ZN(new_n13793_));
  NAND2_X1   g13480(.A1(new_n13793_), .A2(new_n13631_), .ZN(new_n13794_));
  INV_X1     g13481(.I(new_n13794_), .ZN(new_n13795_));
  XOR2_X1    g13482(.A1(new_n13792_), .A2(new_n13795_), .Z(new_n13796_));
  NAND2_X1   g13483(.A1(new_n13796_), .A2(new_n13779_), .ZN(new_n13797_));
  NOR2_X1    g13484(.A1(new_n13792_), .A2(new_n13795_), .ZN(new_n13798_));
  INV_X1     g13485(.I(new_n13798_), .ZN(new_n13799_));
  NAND2_X1   g13486(.A1(new_n13792_), .A2(new_n13795_), .ZN(new_n13800_));
  NAND2_X1   g13487(.A1(new_n13799_), .A2(new_n13800_), .ZN(new_n13801_));
  NAND2_X1   g13488(.A1(new_n13801_), .A2(new_n13778_), .ZN(new_n13802_));
  NAND2_X1   g13489(.A1(new_n13802_), .A2(new_n13797_), .ZN(new_n13803_));
  INV_X1     g13490(.I(new_n13803_), .ZN(new_n13804_));
  XOR2_X1    g13491(.A1(new_n13776_), .A2(new_n13804_), .Z(new_n13805_));
  NOR2_X1    g13492(.A1(new_n13805_), .A2(new_n13745_), .ZN(new_n13806_));
  INV_X1     g13493(.I(new_n13745_), .ZN(new_n13807_));
  NOR3_X1    g13494(.A1(new_n13804_), .A2(new_n13772_), .A3(new_n13775_), .ZN(new_n13808_));
  NOR2_X1    g13495(.A1(new_n13776_), .A2(new_n13803_), .ZN(new_n13809_));
  NOR2_X1    g13496(.A1(new_n13809_), .A2(new_n13808_), .ZN(new_n13810_));
  NOR2_X1    g13497(.A1(new_n13810_), .A2(new_n13807_), .ZN(new_n13811_));
  NOR2_X1    g13498(.A1(new_n13811_), .A2(new_n13806_), .ZN(new_n13812_));
  XNOR2_X1   g13499(.A1(new_n13700_), .A2(new_n13812_), .ZN(new_n13813_));
  XNOR2_X1   g13500(.A1(new_n13700_), .A2(new_n13812_), .ZN(new_n13814_));
  NAND2_X1   g13501(.A1(new_n13814_), .A2(new_n13669_), .ZN(new_n13815_));
  OAI21_X1   g13502(.A1(new_n13669_), .A2(new_n13813_), .B(new_n13815_), .ZN(new_n13816_));
  XOR2_X1    g13503(.A1(new_n13816_), .A2(new_n13668_), .Z(new_n13817_));
  NAND2_X1   g13504(.A1(new_n13667_), .A2(new_n13817_), .ZN(new_n13818_));
  NAND2_X1   g13505(.A1(new_n13816_), .A2(new_n13668_), .ZN(new_n13819_));
  NOR2_X1    g13506(.A1(new_n13816_), .A2(new_n13668_), .ZN(new_n13820_));
  INV_X1     g13507(.I(new_n13820_), .ZN(new_n13821_));
  AND2_X2    g13508(.A1(new_n13821_), .A2(new_n13819_), .Z(new_n13822_));
  OAI21_X1   g13509(.A1(new_n13667_), .A2(new_n13822_), .B(new_n13818_), .ZN(\asquared[86] ));
  NAND2_X1   g13510(.A1(new_n13819_), .A2(new_n13658_), .ZN(new_n13824_));
  OAI21_X1   g13511(.A1(new_n13819_), .A2(new_n13658_), .B(new_n13661_), .ZN(new_n13825_));
  NAND2_X1   g13512(.A1(new_n13825_), .A2(new_n13824_), .ZN(new_n13826_));
  NOR3_X1    g13513(.A1(new_n13494_), .A2(new_n13821_), .A3(new_n13826_), .ZN(\asquared[87] ));
  NOR2_X1    g13514(.A1(new_n13808_), .A2(new_n13807_), .ZN(new_n13828_));
  NOR2_X1    g13515(.A1(new_n13828_), .A2(new_n13809_), .ZN(new_n13829_));
  INV_X1     g13516(.I(new_n13688_), .ZN(new_n13830_));
  OAI21_X1   g13517(.A1(new_n13671_), .A2(new_n13830_), .B(new_n13690_), .ZN(new_n13831_));
  AOI21_X1   g13518(.A1(new_n13773_), .A2(new_n13771_), .B(new_n13769_), .ZN(new_n13832_));
  NAND2_X1   g13519(.A1(new_n13743_), .A2(new_n13702_), .ZN(new_n13833_));
  NAND2_X1   g13520(.A1(new_n13833_), .A2(new_n13742_), .ZN(new_n13834_));
  NOR2_X1    g13521(.A1(new_n1691_), .A2(new_n8453_), .ZN(new_n13835_));
  NAND2_X1   g13522(.A1(\a[25] ), .A2(\a[62] ), .ZN(new_n13836_));
  XNOR2_X1   g13523(.A1(new_n13835_), .A2(new_n13836_), .ZN(new_n13837_));
  NOR2_X1    g13524(.A1(new_n13790_), .A2(new_n13788_), .ZN(new_n13838_));
  NOR2_X1    g13525(.A1(new_n13838_), .A2(new_n13789_), .ZN(new_n13839_));
  INV_X1     g13526(.I(new_n13839_), .ZN(new_n13840_));
  OAI21_X1   g13527(.A1(new_n13747_), .A2(new_n13749_), .B(new_n13835_), .ZN(new_n13841_));
  OAI21_X1   g13528(.A1(new_n13748_), .A2(new_n13750_), .B(new_n13841_), .ZN(new_n13842_));
  AOI21_X1   g13529(.A1(new_n5174_), .A2(new_n9029_), .B(new_n2368_), .ZN(new_n13843_));
  XNOR2_X1   g13530(.A1(new_n13842_), .A2(new_n13843_), .ZN(new_n13844_));
  XOR2_X1    g13531(.A1(new_n13844_), .A2(new_n13840_), .Z(new_n13845_));
  XOR2_X1    g13532(.A1(new_n13845_), .A2(new_n13837_), .Z(new_n13846_));
  XNOR2_X1   g13533(.A1(new_n13846_), .A2(new_n13834_), .ZN(new_n13847_));
  NOR2_X1    g13534(.A1(new_n13847_), .A2(new_n13832_), .ZN(new_n13848_));
  NOR2_X1    g13535(.A1(new_n13846_), .A2(new_n13834_), .ZN(new_n13849_));
  INV_X1     g13536(.I(new_n13849_), .ZN(new_n13850_));
  NAND2_X1   g13537(.A1(new_n13846_), .A2(new_n13834_), .ZN(new_n13851_));
  NAND2_X1   g13538(.A1(new_n13850_), .A2(new_n13851_), .ZN(new_n13852_));
  AOI21_X1   g13539(.A1(new_n13832_), .A2(new_n13852_), .B(new_n13848_), .ZN(new_n13853_));
  XNOR2_X1   g13540(.A1(new_n13853_), .A2(new_n13831_), .ZN(new_n13854_));
  NOR2_X1    g13541(.A1(new_n13853_), .A2(new_n13831_), .ZN(new_n13855_));
  NAND2_X1   g13542(.A1(new_n13853_), .A2(new_n13831_), .ZN(new_n13856_));
  INV_X1     g13543(.I(new_n13856_), .ZN(new_n13857_));
  OAI21_X1   g13544(.A1(new_n13857_), .A2(new_n13855_), .B(new_n13829_), .ZN(new_n13858_));
  OAI21_X1   g13545(.A1(new_n13829_), .A2(new_n13854_), .B(new_n13858_), .ZN(new_n13859_));
  NOR2_X1    g13546(.A1(new_n13684_), .A2(new_n13675_), .ZN(new_n13860_));
  NOR2_X1    g13547(.A1(new_n13860_), .A2(new_n13683_), .ZN(new_n13861_));
  AOI21_X1   g13548(.A1(new_n5592_), .A2(new_n5742_), .B(new_n13708_), .ZN(new_n13862_));
  AOI21_X1   g13549(.A1(new_n5600_), .A2(new_n6030_), .B(new_n13724_), .ZN(new_n13863_));
  INV_X1     g13550(.I(new_n13863_), .ZN(new_n13864_));
  AOI21_X1   g13551(.A1(new_n3126_), .A2(new_n7483_), .B(new_n13727_), .ZN(new_n13865_));
  XOR2_X1    g13552(.A1(new_n13865_), .A2(new_n13864_), .Z(new_n13866_));
  INV_X1     g13553(.I(new_n13865_), .ZN(new_n13867_));
  NOR2_X1    g13554(.A1(new_n13867_), .A2(new_n13864_), .ZN(new_n13868_));
  NOR2_X1    g13555(.A1(new_n13865_), .A2(new_n13863_), .ZN(new_n13869_));
  NOR2_X1    g13556(.A1(new_n13868_), .A2(new_n13869_), .ZN(new_n13870_));
  MUX2_X1    g13557(.I0(new_n13870_), .I1(new_n13866_), .S(new_n13862_), .Z(new_n13871_));
  AOI21_X1   g13558(.A1(new_n4372_), .A2(new_n6777_), .B(new_n13704_), .ZN(new_n13872_));
  AOI21_X1   g13559(.A1(new_n2533_), .A2(new_n8676_), .B(new_n13758_), .ZN(new_n13873_));
  NOR2_X1    g13560(.A1(new_n1674_), .A2(new_n9310_), .ZN(new_n13874_));
  OAI21_X1   g13561(.A1(new_n13711_), .A2(new_n13712_), .B(new_n13874_), .ZN(new_n13875_));
  NAND2_X1   g13562(.A1(new_n13875_), .A2(new_n13713_), .ZN(new_n13876_));
  XOR2_X1    g13563(.A1(new_n13873_), .A2(new_n13876_), .Z(new_n13877_));
  NAND2_X1   g13564(.A1(new_n13877_), .A2(new_n13872_), .ZN(new_n13878_));
  INV_X1     g13565(.I(new_n13872_), .ZN(new_n13879_));
  AND2_X2    g13566(.A1(new_n13873_), .A2(new_n13876_), .Z(new_n13880_));
  NOR2_X1    g13567(.A1(new_n13873_), .A2(new_n13876_), .ZN(new_n13881_));
  OAI21_X1   g13568(.A1(new_n13881_), .A2(new_n13880_), .B(new_n13879_), .ZN(new_n13882_));
  NAND2_X1   g13569(.A1(new_n13882_), .A2(new_n13878_), .ZN(new_n13883_));
  XOR2_X1    g13570(.A1(new_n13871_), .A2(new_n13883_), .Z(new_n13884_));
  INV_X1     g13571(.I(new_n13883_), .ZN(new_n13885_));
  NOR2_X1    g13572(.A1(new_n13871_), .A2(new_n13885_), .ZN(new_n13886_));
  NAND2_X1   g13573(.A1(new_n13871_), .A2(new_n13885_), .ZN(new_n13887_));
  INV_X1     g13574(.I(new_n13887_), .ZN(new_n13888_));
  OAI21_X1   g13575(.A1(new_n13888_), .A2(new_n13886_), .B(new_n13861_), .ZN(new_n13889_));
  OAI21_X1   g13576(.A1(new_n13861_), .A2(new_n13884_), .B(new_n13889_), .ZN(new_n13890_));
  NAND2_X1   g13577(.A1(new_n13800_), .A2(new_n13779_), .ZN(new_n13891_));
  NAND2_X1   g13578(.A1(new_n13891_), .A2(new_n13799_), .ZN(new_n13892_));
  NAND2_X1   g13579(.A1(new_n3838_), .A2(new_n6280_), .ZN(new_n13893_));
  NAND2_X1   g13580(.A1(\a[23] ), .A2(\a[63] ), .ZN(new_n13894_));
  XNOR2_X1   g13581(.A1(new_n13893_), .A2(new_n13894_), .ZN(new_n13895_));
  INV_X1     g13582(.I(new_n13895_), .ZN(new_n13896_));
  AOI22_X1   g13583(.A1(new_n3424_), .A2(new_n7204_), .B1(new_n4372_), .B2(new_n7000_), .ZN(new_n13897_));
  NOR4_X1    g13584(.A1(new_n3487_), .A2(new_n6777_), .A3(new_n2868_), .A4(new_n6694_), .ZN(new_n13898_));
  NAND2_X1   g13585(.A1(new_n13897_), .A2(new_n13898_), .ZN(new_n13899_));
  NAND2_X1   g13586(.A1(\a[55] ), .A2(\a[57] ), .ZN(new_n13900_));
  XOR2_X1    g13587(.A1(new_n3733_), .A2(new_n13900_), .Z(new_n13901_));
  NOR2_X1    g13588(.A1(new_n13899_), .A2(new_n13901_), .ZN(new_n13902_));
  AND2_X2    g13589(.A1(new_n13899_), .A2(new_n13901_), .Z(new_n13903_));
  OAI21_X1   g13590(.A1(new_n13902_), .A2(new_n13903_), .B(new_n13896_), .ZN(new_n13904_));
  XOR2_X1    g13591(.A1(new_n13899_), .A2(new_n13901_), .Z(new_n13905_));
  NAND2_X1   g13592(.A1(new_n13905_), .A2(new_n13895_), .ZN(new_n13906_));
  NAND2_X1   g13593(.A1(new_n13906_), .A2(new_n13904_), .ZN(new_n13907_));
  AOI22_X1   g13594(.A1(new_n2533_), .A2(new_n9554_), .B1(new_n8996_), .B2(new_n3037_), .ZN(new_n13908_));
  NOR2_X1    g13595(.A1(new_n1916_), .A2(new_n8990_), .ZN(new_n13909_));
  NAND4_X1   g13596(.A1(new_n13908_), .A2(new_n2692_), .A3(new_n8677_), .A4(new_n13909_), .ZN(new_n13910_));
  NAND4_X1   g13597(.A1(\a[41] ), .A2(\a[42] ), .A3(\a[44] ), .A4(\a[45] ), .ZN(new_n13912_));
  NAND2_X1   g13598(.A1(new_n5980_), .A2(new_n6024_), .ZN(new_n13913_));
  NAND2_X1   g13599(.A1(\a[30] ), .A2(\a[56] ), .ZN(new_n13914_));
  XNOR2_X1   g13600(.A1(new_n13913_), .A2(new_n13914_), .ZN(new_n13915_));
  NOR2_X1    g13601(.A1(new_n13915_), .A2(new_n13912_), .ZN(new_n13916_));
  INV_X1     g13602(.I(new_n13912_), .ZN(new_n13917_));
  INV_X1     g13603(.I(new_n13915_), .ZN(new_n13918_));
  NOR2_X1    g13604(.A1(new_n13918_), .A2(new_n13917_), .ZN(new_n13919_));
  NOR2_X1    g13605(.A1(new_n13919_), .A2(new_n13916_), .ZN(new_n13920_));
  NOR2_X1    g13606(.A1(new_n13920_), .A2(new_n13910_), .ZN(new_n13921_));
  XOR2_X1    g13607(.A1(new_n13915_), .A2(new_n13917_), .Z(new_n13922_));
  INV_X1     g13608(.I(new_n13922_), .ZN(new_n13923_));
  AOI21_X1   g13609(.A1(new_n13910_), .A2(new_n13923_), .B(new_n13921_), .ZN(new_n13924_));
  XOR2_X1    g13610(.A1(new_n13924_), .A2(new_n13907_), .Z(new_n13925_));
  INV_X1     g13611(.I(new_n13925_), .ZN(new_n13926_));
  INV_X1     g13612(.I(new_n13907_), .ZN(new_n13927_));
  NOR2_X1    g13613(.A1(new_n13924_), .A2(new_n13927_), .ZN(new_n13928_));
  INV_X1     g13614(.I(new_n13928_), .ZN(new_n13929_));
  NAND2_X1   g13615(.A1(new_n13924_), .A2(new_n13927_), .ZN(new_n13930_));
  AOI21_X1   g13616(.A1(new_n13929_), .A2(new_n13930_), .B(new_n13892_), .ZN(new_n13931_));
  AOI21_X1   g13617(.A1(new_n13892_), .A2(new_n13926_), .B(new_n13931_), .ZN(new_n13932_));
  AOI21_X1   g13618(.A1(new_n13757_), .A2(new_n13764_), .B(new_n13762_), .ZN(new_n13933_));
  NOR2_X1    g13619(.A1(new_n13717_), .A2(new_n13706_), .ZN(new_n13934_));
  NOR2_X1    g13620(.A1(new_n13934_), .A2(new_n13716_), .ZN(new_n13935_));
  NOR2_X1    g13621(.A1(new_n13735_), .A2(new_n13725_), .ZN(new_n13936_));
  NOR2_X1    g13622(.A1(new_n13936_), .A2(new_n13732_), .ZN(new_n13937_));
  XNOR2_X1   g13623(.A1(new_n13935_), .A2(new_n13937_), .ZN(new_n13938_));
  NOR2_X1    g13624(.A1(new_n13938_), .A2(new_n13933_), .ZN(new_n13939_));
  INV_X1     g13625(.I(new_n13933_), .ZN(new_n13940_));
  NOR2_X1    g13626(.A1(new_n13935_), .A2(new_n13937_), .ZN(new_n13941_));
  INV_X1     g13627(.I(new_n13941_), .ZN(new_n13942_));
  NAND2_X1   g13628(.A1(new_n13935_), .A2(new_n13937_), .ZN(new_n13943_));
  AOI21_X1   g13629(.A1(new_n13942_), .A2(new_n13943_), .B(new_n13940_), .ZN(new_n13944_));
  NOR2_X1    g13630(.A1(new_n13939_), .A2(new_n13944_), .ZN(new_n13945_));
  NOR2_X1    g13631(.A1(new_n13932_), .A2(new_n13945_), .ZN(new_n13946_));
  NAND2_X1   g13632(.A1(new_n13932_), .A2(new_n13945_), .ZN(new_n13947_));
  INV_X1     g13633(.I(new_n13947_), .ZN(new_n13948_));
  OAI21_X1   g13634(.A1(new_n13948_), .A2(new_n13946_), .B(new_n13890_), .ZN(new_n13949_));
  XNOR2_X1   g13635(.A1(new_n13932_), .A2(new_n13945_), .ZN(new_n13950_));
  OAI21_X1   g13636(.A1(new_n13890_), .A2(new_n13950_), .B(new_n13949_), .ZN(new_n13951_));
  NOR2_X1    g13637(.A1(new_n13859_), .A2(new_n13951_), .ZN(new_n13952_));
  NAND2_X1   g13638(.A1(new_n13698_), .A2(new_n13670_), .ZN(new_n13953_));
  AOI22_X1   g13639(.A1(new_n13859_), .A2(new_n13951_), .B1(new_n13697_), .B2(new_n13953_), .ZN(new_n13954_));
  NOR2_X1    g13640(.A1(new_n13954_), .A2(new_n13952_), .ZN(new_n13955_));
  OAI21_X1   g13641(.A1(new_n13832_), .A2(new_n13849_), .B(new_n13851_), .ZN(new_n13956_));
  NAND2_X1   g13642(.A1(new_n13892_), .A2(new_n13930_), .ZN(new_n13957_));
  NAND2_X1   g13643(.A1(new_n13957_), .A2(new_n13929_), .ZN(new_n13958_));
  INV_X1     g13644(.I(new_n13869_), .ZN(new_n13959_));
  AOI21_X1   g13645(.A1(new_n13862_), .A2(new_n13959_), .B(new_n13868_), .ZN(new_n13960_));
  INV_X1     g13646(.I(new_n13902_), .ZN(new_n13961_));
  OAI21_X1   g13647(.A1(new_n13895_), .A2(new_n13903_), .B(new_n13961_), .ZN(new_n13962_));
  INV_X1     g13648(.I(new_n13916_), .ZN(new_n13963_));
  OAI21_X1   g13649(.A1(new_n13910_), .A2(new_n13919_), .B(new_n13963_), .ZN(new_n13964_));
  XNOR2_X1   g13650(.A1(new_n13964_), .A2(new_n13962_), .ZN(new_n13965_));
  NOR2_X1    g13651(.A1(new_n13965_), .A2(new_n13960_), .ZN(new_n13966_));
  INV_X1     g13652(.I(new_n13960_), .ZN(new_n13967_));
  NAND2_X1   g13653(.A1(new_n13964_), .A2(new_n13962_), .ZN(new_n13968_));
  NOR2_X1    g13654(.A1(new_n13964_), .A2(new_n13962_), .ZN(new_n13969_));
  INV_X1     g13655(.I(new_n13969_), .ZN(new_n13970_));
  AOI21_X1   g13656(.A1(new_n13970_), .A2(new_n13968_), .B(new_n13967_), .ZN(new_n13971_));
  NOR2_X1    g13657(.A1(new_n13966_), .A2(new_n13971_), .ZN(new_n13972_));
  XNOR2_X1   g13658(.A1(new_n13958_), .A2(new_n13972_), .ZN(new_n13973_));
  INV_X1     g13659(.I(new_n13973_), .ZN(new_n13974_));
  NOR2_X1    g13660(.A1(new_n13958_), .A2(new_n13972_), .ZN(new_n13975_));
  INV_X1     g13661(.I(new_n13975_), .ZN(new_n13976_));
  NAND2_X1   g13662(.A1(new_n13958_), .A2(new_n13972_), .ZN(new_n13977_));
  AOI21_X1   g13663(.A1(new_n13976_), .A2(new_n13977_), .B(new_n13956_), .ZN(new_n13978_));
  AOI21_X1   g13664(.A1(new_n13956_), .A2(new_n13974_), .B(new_n13978_), .ZN(new_n13979_));
  INV_X1     g13665(.I(new_n13979_), .ZN(new_n13980_));
  OAI21_X1   g13666(.A1(new_n13829_), .A2(new_n13855_), .B(new_n13856_), .ZN(new_n13981_));
  INV_X1     g13667(.I(new_n13981_), .ZN(new_n13982_));
  OAI21_X1   g13668(.A1(new_n13890_), .A2(new_n13946_), .B(new_n13947_), .ZN(new_n13983_));
  INV_X1     g13669(.I(new_n13983_), .ZN(new_n13984_));
  OAI21_X1   g13670(.A1(new_n13861_), .A2(new_n13886_), .B(new_n13887_), .ZN(new_n13985_));
  INV_X1     g13671(.I(new_n13842_), .ZN(new_n13986_));
  NOR2_X1    g13672(.A1(new_n13839_), .A2(new_n13986_), .ZN(new_n13987_));
  XNOR2_X1   g13673(.A1(new_n13837_), .A2(new_n13843_), .ZN(new_n13988_));
  AOI21_X1   g13674(.A1(new_n13839_), .A2(new_n13986_), .B(new_n13988_), .ZN(new_n13989_));
  NOR2_X1    g13675(.A1(new_n13989_), .A2(new_n13987_), .ZN(new_n13990_));
  NOR4_X1    g13676(.A1(new_n4414_), .A2(new_n4769_), .A3(new_n4770_), .A4(new_n5004_), .ZN(new_n13991_));
  INV_X1     g13677(.I(new_n13991_), .ZN(new_n13992_));
  NOR2_X1    g13678(.A1(\a[30] ), .A2(\a[56] ), .ZN(new_n13993_));
  OAI21_X1   g13679(.A1(new_n4321_), .A2(new_n5793_), .B(new_n13993_), .ZN(new_n13994_));
  OAI21_X1   g13680(.A1(new_n6024_), .A2(new_n5980_), .B(new_n13994_), .ZN(new_n13995_));
  AOI21_X1   g13681(.A1(new_n3733_), .A2(new_n6743_), .B(new_n10958_), .ZN(new_n13996_));
  XNOR2_X1   g13682(.A1(new_n13995_), .A2(new_n13996_), .ZN(new_n13997_));
  NOR2_X1    g13683(.A1(new_n13997_), .A2(new_n13992_), .ZN(new_n13998_));
  NOR2_X1    g13684(.A1(new_n13995_), .A2(new_n13996_), .ZN(new_n13999_));
  INV_X1     g13685(.I(new_n13999_), .ZN(new_n14000_));
  NAND2_X1   g13686(.A1(new_n13995_), .A2(new_n13996_), .ZN(new_n14001_));
  AOI21_X1   g13687(.A1(new_n14000_), .A2(new_n14001_), .B(new_n13991_), .ZN(new_n14002_));
  NOR2_X1    g13688(.A1(new_n13998_), .A2(new_n14002_), .ZN(new_n14003_));
  NAND2_X1   g13689(.A1(new_n3838_), .A2(new_n6280_), .ZN(new_n14004_));
  NOR2_X1    g13690(.A1(new_n3838_), .A2(new_n6280_), .ZN(new_n14005_));
  NOR2_X1    g13691(.A1(\a[23] ), .A2(\a[63] ), .ZN(new_n14006_));
  AOI21_X1   g13692(.A1(new_n14004_), .A2(new_n14006_), .B(new_n14005_), .ZN(new_n14007_));
  AOI21_X1   g13693(.A1(new_n3487_), .A2(new_n6777_), .B(new_n13897_), .ZN(new_n14008_));
  AOI21_X1   g13694(.A1(new_n2797_), .A2(new_n8676_), .B(new_n13908_), .ZN(new_n14009_));
  XNOR2_X1   g13695(.A1(new_n14008_), .A2(new_n14009_), .ZN(new_n14010_));
  INV_X1     g13696(.I(new_n14008_), .ZN(new_n14011_));
  INV_X1     g13697(.I(new_n14009_), .ZN(new_n14012_));
  NOR2_X1    g13698(.A1(new_n14011_), .A2(new_n14012_), .ZN(new_n14013_));
  NOR2_X1    g13699(.A1(new_n14008_), .A2(new_n14009_), .ZN(new_n14014_));
  NOR2_X1    g13700(.A1(new_n14013_), .A2(new_n14014_), .ZN(new_n14015_));
  MUX2_X1    g13701(.I0(new_n14015_), .I1(new_n14010_), .S(new_n14007_), .Z(new_n14016_));
  XNOR2_X1   g13702(.A1(new_n14016_), .A2(new_n14003_), .ZN(new_n14017_));
  NOR2_X1    g13703(.A1(new_n14017_), .A2(new_n13990_), .ZN(new_n14018_));
  INV_X1     g13704(.I(new_n13990_), .ZN(new_n14019_));
  NOR2_X1    g13705(.A1(new_n14016_), .A2(new_n14003_), .ZN(new_n14020_));
  INV_X1     g13706(.I(new_n14020_), .ZN(new_n14021_));
  NAND2_X1   g13707(.A1(new_n14016_), .A2(new_n14003_), .ZN(new_n14022_));
  AOI21_X1   g13708(.A1(new_n14021_), .A2(new_n14022_), .B(new_n14019_), .ZN(new_n14023_));
  NOR2_X1    g13709(.A1(new_n14023_), .A2(new_n14018_), .ZN(new_n14024_));
  AOI21_X1   g13710(.A1(new_n13940_), .A2(new_n13943_), .B(new_n13941_), .ZN(new_n14025_));
  INV_X1     g13711(.I(new_n14025_), .ZN(new_n14026_));
  XOR2_X1    g13712(.A1(new_n14024_), .A2(new_n14026_), .Z(new_n14027_));
  NAND2_X1   g13713(.A1(new_n14027_), .A2(new_n13985_), .ZN(new_n14028_));
  INV_X1     g13714(.I(new_n14024_), .ZN(new_n14029_));
  NOR2_X1    g13715(.A1(new_n14029_), .A2(new_n14025_), .ZN(new_n14030_));
  NOR2_X1    g13716(.A1(new_n14024_), .A2(new_n14026_), .ZN(new_n14031_));
  NOR2_X1    g13717(.A1(new_n14030_), .A2(new_n14031_), .ZN(new_n14032_));
  OAI21_X1   g13718(.A1(new_n13985_), .A2(new_n14032_), .B(new_n14028_), .ZN(new_n14033_));
  NOR2_X1    g13719(.A1(new_n6694_), .A2(new_n7727_), .ZN(new_n14034_));
  INV_X1     g13720(.I(new_n14034_), .ZN(new_n14035_));
  NOR2_X1    g13721(.A1(new_n4041_), .A2(new_n14035_), .ZN(new_n14036_));
  NOR2_X1    g13722(.A1(new_n3371_), .A2(new_n8085_), .ZN(new_n14037_));
  NAND4_X1   g13723(.A1(new_n14036_), .A2(\a[28] ), .A3(new_n14037_), .A4(\a[53] ), .ZN(new_n14038_));
  AOI21_X1   g13724(.A1(new_n14038_), .A2(new_n8675_), .B(new_n3355_), .ZN(new_n14039_));
  NAND2_X1   g13725(.A1(\a[28] ), .A2(\a[59] ), .ZN(new_n14040_));
  NOR2_X1    g13726(.A1(new_n14039_), .A2(new_n14036_), .ZN(new_n14041_));
  INV_X1     g13727(.I(new_n14041_), .ZN(new_n14042_));
  NAND2_X1   g13728(.A1(new_n4041_), .A2(new_n14035_), .ZN(new_n14043_));
  OAI22_X1   g13729(.A1(new_n14042_), .A2(new_n14043_), .B1(new_n14039_), .B2(new_n14040_), .ZN(new_n14044_));
  INV_X1     g13730(.I(new_n14044_), .ZN(new_n14045_));
  NOR2_X1    g13731(.A1(new_n2499_), .A2(new_n6692_), .ZN(new_n14046_));
  NOR2_X1    g13732(.A1(new_n3423_), .A2(new_n7647_), .ZN(new_n14047_));
  AOI22_X1   g13733(.A1(new_n3966_), .A2(new_n14047_), .B1(new_n6777_), .B2(new_n14046_), .ZN(new_n14048_));
  INV_X1     g13734(.I(new_n14048_), .ZN(new_n14049_));
  NOR2_X1    g13735(.A1(new_n2499_), .A2(new_n7647_), .ZN(new_n14050_));
  NOR2_X1    g13736(.A1(new_n3393_), .A2(new_n6260_), .ZN(new_n14051_));
  XNOR2_X1   g13737(.A1(new_n14050_), .A2(new_n14051_), .ZN(new_n14052_));
  NOR2_X1    g13738(.A1(new_n14052_), .A2(new_n14050_), .ZN(new_n14053_));
  NOR2_X1    g13739(.A1(new_n14049_), .A2(new_n14053_), .ZN(new_n14054_));
  OAI21_X1   g13740(.A1(new_n3423_), .A2(new_n6692_), .B(new_n14052_), .ZN(new_n14055_));
  INV_X1     g13741(.I(new_n14055_), .ZN(new_n14056_));
  NOR2_X1    g13742(.A1(new_n14056_), .A2(new_n14054_), .ZN(new_n14057_));
  AOI22_X1   g13743(.A1(new_n13837_), .A2(new_n2277_), .B1(new_n9784_), .B2(new_n13843_), .ZN(new_n14058_));
  XNOR2_X1   g13744(.A1(new_n14057_), .A2(new_n14058_), .ZN(new_n14059_));
  INV_X1     g13745(.I(new_n14057_), .ZN(new_n14060_));
  NOR2_X1    g13746(.A1(new_n14060_), .A2(new_n14058_), .ZN(new_n14061_));
  INV_X1     g13747(.I(new_n14061_), .ZN(new_n14062_));
  NAND2_X1   g13748(.A1(new_n14060_), .A2(new_n14058_), .ZN(new_n14063_));
  AOI21_X1   g13749(.A1(new_n14062_), .A2(new_n14063_), .B(new_n14045_), .ZN(new_n14064_));
  AOI21_X1   g13750(.A1(new_n14045_), .A2(new_n14059_), .B(new_n14064_), .ZN(new_n14065_));
  NOR2_X1    g13751(.A1(new_n13879_), .A2(new_n13881_), .ZN(new_n14066_));
  NOR2_X1    g13752(.A1(new_n14066_), .A2(new_n13880_), .ZN(new_n14067_));
  NAND2_X1   g13753(.A1(new_n2869_), .A2(new_n7421_), .ZN(new_n14068_));
  NOR2_X1    g13754(.A1(new_n4240_), .A2(new_n5511_), .ZN(new_n14069_));
  XOR2_X1    g13755(.A1(new_n14068_), .A2(new_n14069_), .Z(new_n14070_));
  NAND2_X1   g13756(.A1(\a[25] ), .A2(\a[44] ), .ZN(new_n14071_));
  NAND2_X1   g13757(.A1(\a[43] ), .A2(\a[62] ), .ZN(new_n14072_));
  XNOR2_X1   g13758(.A1(new_n14071_), .A2(new_n14072_), .ZN(new_n14073_));
  XNOR2_X1   g13759(.A1(new_n14070_), .A2(new_n14073_), .ZN(new_n14074_));
  NOR2_X1    g13760(.A1(new_n14067_), .A2(new_n14074_), .ZN(new_n14075_));
  INV_X1     g13761(.I(new_n14067_), .ZN(new_n14076_));
  NOR2_X1    g13762(.A1(new_n14070_), .A2(new_n14073_), .ZN(new_n14077_));
  INV_X1     g13763(.I(new_n14077_), .ZN(new_n14078_));
  NAND2_X1   g13764(.A1(new_n14070_), .A2(new_n14073_), .ZN(new_n14079_));
  AOI21_X1   g13765(.A1(new_n14078_), .A2(new_n14079_), .B(new_n14076_), .ZN(new_n14080_));
  NOR2_X1    g13766(.A1(new_n14080_), .A2(new_n14075_), .ZN(new_n14081_));
  NOR2_X1    g13767(.A1(new_n8992_), .A2(new_n2534_), .ZN(new_n14082_));
  NOR2_X1    g13768(.A1(new_n8992_), .A2(new_n2534_), .ZN(new_n14086_));
  INV_X1     g13769(.I(new_n14086_), .ZN(new_n14087_));
  AOI21_X1   g13770(.A1(new_n5600_), .A2(new_n5601_), .B(new_n13261_), .ZN(new_n14088_));
  NOR2_X1    g13771(.A1(new_n3837_), .A2(new_n6055_), .ZN(new_n14089_));
  AND4_X2    g13772(.A1(new_n5340_), .A2(new_n14088_), .A3(new_n12355_), .A4(new_n14089_), .Z(new_n14090_));
  NAND2_X1   g13773(.A1(new_n5350_), .A2(new_n5488_), .ZN(new_n14091_));
  NAND2_X1   g13774(.A1(\a[32] ), .A2(\a[55] ), .ZN(new_n14092_));
  XNOR2_X1   g13775(.A1(new_n14091_), .A2(new_n14092_), .ZN(new_n14093_));
  INV_X1     g13776(.I(new_n14093_), .ZN(new_n14094_));
  NAND2_X1   g13777(.A1(new_n14090_), .A2(new_n14094_), .ZN(new_n14095_));
  OR2_X2     g13778(.A1(new_n14090_), .A2(new_n14094_), .Z(new_n14096_));
  AOI21_X1   g13779(.A1(new_n14096_), .A2(new_n14095_), .B(new_n14087_), .ZN(new_n14097_));
  XOR2_X1    g13780(.A1(new_n14090_), .A2(new_n14093_), .Z(new_n14098_));
  NOR2_X1    g13781(.A1(new_n14098_), .A2(new_n14086_), .ZN(new_n14099_));
  OAI21_X1   g13782(.A1(new_n14097_), .A2(new_n14099_), .B(new_n14081_), .ZN(new_n14100_));
  NOR2_X1    g13783(.A1(new_n14099_), .A2(new_n14097_), .ZN(new_n14101_));
  OAI21_X1   g13784(.A1(new_n14075_), .A2(new_n14080_), .B(new_n14101_), .ZN(new_n14102_));
  NAND2_X1   g13785(.A1(new_n14100_), .A2(new_n14102_), .ZN(new_n14103_));
  XNOR2_X1   g13786(.A1(new_n14081_), .A2(new_n14101_), .ZN(new_n14104_));
  MUX2_X1    g13787(.I0(new_n14103_), .I1(new_n14104_), .S(new_n14065_), .Z(new_n14105_));
  NAND2_X1   g13788(.A1(new_n14033_), .A2(new_n14105_), .ZN(new_n14106_));
  NOR2_X1    g13789(.A1(new_n14033_), .A2(new_n14105_), .ZN(new_n14107_));
  INV_X1     g13790(.I(new_n14107_), .ZN(new_n14108_));
  AOI21_X1   g13791(.A1(new_n14108_), .A2(new_n14106_), .B(new_n13984_), .ZN(new_n14109_));
  XNOR2_X1   g13792(.A1(new_n14033_), .A2(new_n14105_), .ZN(new_n14110_));
  NOR2_X1    g13793(.A1(new_n14110_), .A2(new_n13983_), .ZN(new_n14111_));
  NOR2_X1    g13794(.A1(new_n14111_), .A2(new_n14109_), .ZN(new_n14112_));
  NOR2_X1    g13795(.A1(new_n14112_), .A2(new_n13982_), .ZN(new_n14113_));
  NOR3_X1    g13796(.A1(new_n14111_), .A2(new_n13981_), .A3(new_n14109_), .ZN(new_n14114_));
  OAI21_X1   g13797(.A1(new_n14113_), .A2(new_n14114_), .B(new_n13980_), .ZN(new_n14115_));
  XOR2_X1    g13798(.A1(new_n14112_), .A2(new_n13982_), .Z(new_n14116_));
  NAND2_X1   g13799(.A1(new_n14116_), .A2(new_n13979_), .ZN(new_n14117_));
  NAND2_X1   g13800(.A1(new_n14117_), .A2(new_n14115_), .ZN(new_n14118_));
  XOR2_X1    g13801(.A1(new_n14118_), .A2(new_n13955_), .Z(new_n14119_));
  NAND2_X1   g13802(.A1(\asquared[87] ), .A2(new_n14119_), .ZN(new_n14120_));
  NAND2_X1   g13803(.A1(new_n14118_), .A2(new_n13955_), .ZN(new_n14121_));
  INV_X1     g13804(.I(new_n13955_), .ZN(new_n14122_));
  INV_X1     g13805(.I(new_n14118_), .ZN(new_n14123_));
  NAND2_X1   g13806(.A1(new_n14123_), .A2(new_n14122_), .ZN(new_n14124_));
  AND2_X2    g13807(.A1(new_n14124_), .A2(new_n14121_), .Z(new_n14125_));
  OAI21_X1   g13808(.A1(\asquared[87] ), .A2(new_n14125_), .B(new_n14120_), .ZN(\asquared[88] ));
  NAND2_X1   g13809(.A1(\asquared[87] ), .A2(new_n14121_), .ZN(new_n14127_));
  NAND2_X1   g13810(.A1(new_n14127_), .A2(new_n14124_), .ZN(new_n14128_));
  NAND2_X1   g13811(.A1(new_n13956_), .A2(new_n13976_), .ZN(new_n14129_));
  NAND2_X1   g13812(.A1(new_n14129_), .A2(new_n13977_), .ZN(new_n14130_));
  OAI21_X1   g13813(.A1(new_n13990_), .A2(new_n14020_), .B(new_n14022_), .ZN(new_n14131_));
  AOI21_X1   g13814(.A1(new_n4515_), .A2(new_n9781_), .B(new_n14082_), .ZN(new_n14132_));
  INV_X1     g13815(.I(new_n14132_), .ZN(new_n14133_));
  AOI21_X1   g13816(.A1(new_n5339_), .A2(new_n6028_), .B(new_n14088_), .ZN(new_n14134_));
  XNOR2_X1   g13817(.A1(new_n14041_), .A2(new_n14134_), .ZN(new_n14135_));
  NOR2_X1    g13818(.A1(new_n14135_), .A2(new_n14133_), .ZN(new_n14136_));
  INV_X1     g13819(.I(new_n14134_), .ZN(new_n14137_));
  NOR2_X1    g13820(.A1(new_n14042_), .A2(new_n14137_), .ZN(new_n14138_));
  NOR2_X1    g13821(.A1(new_n14041_), .A2(new_n14134_), .ZN(new_n14139_));
  NOR2_X1    g13822(.A1(new_n14138_), .A2(new_n14139_), .ZN(new_n14140_));
  NOR2_X1    g13823(.A1(new_n14140_), .A2(new_n14132_), .ZN(new_n14141_));
  NOR2_X1    g13824(.A1(new_n14141_), .A2(new_n14136_), .ZN(new_n14142_));
  INV_X1     g13825(.I(new_n14142_), .ZN(new_n14143_));
  NAND2_X1   g13826(.A1(new_n14076_), .A2(new_n14079_), .ZN(new_n14144_));
  NAND2_X1   g13827(.A1(new_n14144_), .A2(new_n14078_), .ZN(new_n14145_));
  INV_X1     g13828(.I(new_n14145_), .ZN(new_n14146_));
  NAND2_X1   g13829(.A1(new_n2869_), .A2(new_n7421_), .ZN(new_n14147_));
  NOR2_X1    g13830(.A1(new_n2869_), .A2(new_n7421_), .ZN(new_n14148_));
  NOR2_X1    g13831(.A1(\a[40] ), .A2(\a[47] ), .ZN(new_n14149_));
  AOI21_X1   g13832(.A1(new_n14147_), .A2(new_n14149_), .B(new_n14148_), .ZN(new_n14150_));
  AOI21_X1   g13833(.A1(new_n14050_), .A2(new_n14051_), .B(new_n14048_), .ZN(new_n14151_));
  INV_X1     g13834(.I(new_n14151_), .ZN(new_n14152_));
  NAND2_X1   g13835(.A1(\a[54] ), .A2(\a[55] ), .ZN(new_n14153_));
  XOR2_X1    g13836(.A1(new_n4372_), .A2(new_n14153_), .Z(new_n14154_));
  NOR2_X1    g13837(.A1(new_n14152_), .A2(new_n14154_), .ZN(new_n14155_));
  INV_X1     g13838(.I(new_n14155_), .ZN(new_n14156_));
  INV_X1     g13839(.I(new_n14154_), .ZN(new_n14157_));
  NOR2_X1    g13840(.A1(new_n14157_), .A2(new_n14151_), .ZN(new_n14158_));
  INV_X1     g13841(.I(new_n14158_), .ZN(new_n14159_));
  NAND2_X1   g13842(.A1(new_n14156_), .A2(new_n14159_), .ZN(new_n14160_));
  XOR2_X1    g13843(.A1(new_n14151_), .A2(new_n14154_), .Z(new_n14161_));
  NOR2_X1    g13844(.A1(new_n14161_), .A2(new_n14150_), .ZN(new_n14162_));
  AOI21_X1   g13845(.A1(new_n14150_), .A2(new_n14160_), .B(new_n14162_), .ZN(new_n14163_));
  NOR2_X1    g13846(.A1(new_n14146_), .A2(new_n14163_), .ZN(new_n14164_));
  NAND2_X1   g13847(.A1(new_n14146_), .A2(new_n14163_), .ZN(new_n14165_));
  INV_X1     g13848(.I(new_n14165_), .ZN(new_n14166_));
  OAI21_X1   g13849(.A1(new_n14166_), .A2(new_n14164_), .B(new_n14143_), .ZN(new_n14167_));
  XOR2_X1    g13850(.A1(new_n14145_), .A2(new_n14163_), .Z(new_n14168_));
  OAI21_X1   g13851(.A1(new_n14143_), .A2(new_n14168_), .B(new_n14167_), .ZN(new_n14169_));
  OAI21_X1   g13852(.A1(new_n13960_), .A2(new_n13969_), .B(new_n13968_), .ZN(new_n14170_));
  INV_X1     g13853(.I(new_n14170_), .ZN(new_n14171_));
  XOR2_X1    g13854(.A1(new_n14169_), .A2(new_n14171_), .Z(new_n14172_));
  NOR2_X1    g13855(.A1(new_n14169_), .A2(new_n14171_), .ZN(new_n14173_));
  INV_X1     g13856(.I(new_n14173_), .ZN(new_n14174_));
  NAND2_X1   g13857(.A1(new_n14169_), .A2(new_n14171_), .ZN(new_n14175_));
  AOI21_X1   g13858(.A1(new_n14174_), .A2(new_n14175_), .B(new_n14131_), .ZN(new_n14176_));
  AOI21_X1   g13859(.A1(new_n14131_), .A2(new_n14172_), .B(new_n14176_), .ZN(new_n14177_));
  NAND2_X1   g13860(.A1(new_n14001_), .A2(new_n13991_), .ZN(new_n14178_));
  NAND2_X1   g13861(.A1(new_n14178_), .A2(new_n14000_), .ZN(new_n14179_));
  NAND2_X1   g13862(.A1(new_n5339_), .A2(new_n6280_), .ZN(new_n14180_));
  NOR2_X1    g13863(.A1(new_n2499_), .A2(new_n8085_), .ZN(new_n14181_));
  XOR2_X1    g13864(.A1(new_n14180_), .A2(new_n14181_), .Z(new_n14182_));
  NOR2_X1    g13865(.A1(new_n4240_), .A2(new_n5750_), .ZN(new_n14183_));
  NAND2_X1   g13866(.A1(\a[56] ), .A2(\a[58] ), .ZN(new_n14184_));
  XOR2_X1    g13867(.A1(new_n2766_), .A2(new_n14184_), .Z(new_n14185_));
  XOR2_X1    g13868(.A1(new_n14182_), .A2(new_n14185_), .Z(new_n14186_));
  NOR2_X1    g13869(.A1(new_n14182_), .A2(new_n14185_), .ZN(new_n14187_));
  INV_X1     g13870(.I(new_n14187_), .ZN(new_n14188_));
  NAND2_X1   g13871(.A1(new_n14182_), .A2(new_n14185_), .ZN(new_n14189_));
  AOI21_X1   g13872(.A1(new_n14188_), .A2(new_n14189_), .B(new_n14179_), .ZN(new_n14190_));
  AOI21_X1   g13873(.A1(new_n14179_), .A2(new_n14186_), .B(new_n14190_), .ZN(new_n14191_));
  NOR2_X1    g13874(.A1(new_n8574_), .A2(new_n9394_), .ZN(new_n14192_));
  NOR2_X1    g13875(.A1(new_n1916_), .A2(new_n9029_), .ZN(new_n14193_));
  NAND4_X1   g13876(.A1(new_n14192_), .A2(new_n2692_), .A3(new_n8992_), .A4(new_n14193_), .ZN(new_n14194_));
  NAND2_X1   g13877(.A1(new_n5350_), .A2(new_n5980_), .ZN(new_n14195_));
  NOR2_X1    g13878(.A1(new_n2655_), .A2(new_n7727_), .ZN(new_n14196_));
  XOR2_X1    g13879(.A1(new_n14195_), .A2(new_n14196_), .Z(new_n14197_));
  AOI21_X1   g13880(.A1(new_n3966_), .A2(new_n5184_), .B(new_n13703_), .ZN(new_n14198_));
  NOR4_X1    g13881(.A1(new_n3838_), .A2(new_n6777_), .A3(new_n3423_), .A4(new_n6694_), .ZN(new_n14199_));
  NAND2_X1   g13882(.A1(new_n14198_), .A2(new_n14199_), .ZN(new_n14200_));
  NOR2_X1    g13883(.A1(new_n14200_), .A2(new_n14197_), .ZN(new_n14201_));
  INV_X1     g13884(.I(new_n14201_), .ZN(new_n14202_));
  NAND2_X1   g13885(.A1(new_n14200_), .A2(new_n14197_), .ZN(new_n14203_));
  AOI21_X1   g13886(.A1(new_n14202_), .A2(new_n14203_), .B(new_n14194_), .ZN(new_n14204_));
  INV_X1     g13887(.I(new_n14194_), .ZN(new_n14205_));
  XNOR2_X1   g13888(.A1(new_n14200_), .A2(new_n14197_), .ZN(new_n14206_));
  NOR2_X1    g13889(.A1(new_n14206_), .A2(new_n14205_), .ZN(new_n14207_));
  NOR2_X1    g13890(.A1(new_n14207_), .A2(new_n14204_), .ZN(new_n14208_));
  NOR2_X1    g13891(.A1(new_n5350_), .A2(new_n5488_), .ZN(new_n14209_));
  NAND2_X1   g13892(.A1(new_n2765_), .A2(new_n6999_), .ZN(new_n14210_));
  AOI21_X1   g13893(.A1(new_n5350_), .A2(new_n5488_), .B(new_n14210_), .ZN(new_n14211_));
  NOR2_X1    g13894(.A1(new_n14211_), .A2(new_n14209_), .ZN(new_n14212_));
  INV_X1     g13895(.I(new_n14212_), .ZN(new_n14213_));
  NOR2_X1    g13896(.A1(new_n4770_), .A2(new_n9029_), .ZN(new_n14214_));
  AOI21_X1   g13897(.A1(\a[25] ), .A2(new_n14214_), .B(new_n5321_), .ZN(new_n14215_));
  INV_X1     g13898(.I(new_n14215_), .ZN(new_n14216_));
  NOR2_X1    g13899(.A1(new_n14213_), .A2(new_n14216_), .ZN(new_n14217_));
  XOR2_X1    g13900(.A1(new_n14217_), .A2(new_n1999_), .Z(new_n14218_));
  XOR2_X1    g13901(.A1(new_n14218_), .A2(\a[63] ), .Z(new_n14219_));
  XOR2_X1    g13902(.A1(new_n14219_), .A2(new_n14208_), .Z(new_n14220_));
  INV_X1     g13903(.I(new_n14208_), .ZN(new_n14221_));
  NOR2_X1    g13904(.A1(new_n14221_), .A2(new_n14219_), .ZN(new_n14222_));
  NAND2_X1   g13905(.A1(new_n14221_), .A2(new_n14219_), .ZN(new_n14223_));
  INV_X1     g13906(.I(new_n14223_), .ZN(new_n14224_));
  OAI21_X1   g13907(.A1(new_n14224_), .A2(new_n14222_), .B(new_n14191_), .ZN(new_n14225_));
  OAI21_X1   g13908(.A1(new_n14191_), .A2(new_n14220_), .B(new_n14225_), .ZN(new_n14226_));
  NAND2_X1   g13909(.A1(new_n14177_), .A2(new_n14226_), .ZN(new_n14227_));
  OR2_X2     g13910(.A1(new_n14177_), .A2(new_n14226_), .Z(new_n14228_));
  NAND2_X1   g13911(.A1(new_n14228_), .A2(new_n14227_), .ZN(new_n14229_));
  XNOR2_X1   g13912(.A1(new_n14177_), .A2(new_n14226_), .ZN(new_n14230_));
  NOR2_X1    g13913(.A1(new_n14230_), .A2(new_n14130_), .ZN(new_n14231_));
  AOI21_X1   g13914(.A1(new_n14130_), .A2(new_n14229_), .B(new_n14231_), .ZN(new_n14232_));
  NAND2_X1   g13915(.A1(new_n14106_), .A2(new_n13983_), .ZN(new_n14233_));
  NAND2_X1   g13916(.A1(new_n14233_), .A2(new_n14108_), .ZN(new_n14234_));
  INV_X1     g13917(.I(new_n14030_), .ZN(new_n14235_));
  OAI21_X1   g13918(.A1(new_n14024_), .A2(new_n14026_), .B(new_n13985_), .ZN(new_n14236_));
  NAND2_X1   g13919(.A1(new_n14235_), .A2(new_n14236_), .ZN(new_n14237_));
  INV_X1     g13920(.I(new_n14237_), .ZN(new_n14238_));
  AOI21_X1   g13921(.A1(new_n14045_), .A2(new_n14063_), .B(new_n14061_), .ZN(new_n14239_));
  INV_X1     g13922(.I(new_n14239_), .ZN(new_n14240_));
  NAND2_X1   g13923(.A1(new_n14096_), .A2(new_n14086_), .ZN(new_n14241_));
  NAND2_X1   g13924(.A1(new_n14241_), .A2(new_n14095_), .ZN(new_n14242_));
  INV_X1     g13925(.I(new_n14014_), .ZN(new_n14243_));
  AOI21_X1   g13926(.A1(new_n14007_), .A2(new_n14243_), .B(new_n14013_), .ZN(new_n14244_));
  XNOR2_X1   g13927(.A1(new_n14242_), .A2(new_n14244_), .ZN(new_n14245_));
  INV_X1     g13928(.I(new_n14242_), .ZN(new_n14246_));
  NOR2_X1    g13929(.A1(new_n14246_), .A2(new_n14244_), .ZN(new_n14247_));
  INV_X1     g13930(.I(new_n14247_), .ZN(new_n14248_));
  NAND2_X1   g13931(.A1(new_n14246_), .A2(new_n14244_), .ZN(new_n14249_));
  AOI21_X1   g13932(.A1(new_n14248_), .A2(new_n14249_), .B(new_n14240_), .ZN(new_n14250_));
  AOI21_X1   g13933(.A1(new_n14240_), .A2(new_n14245_), .B(new_n14250_), .ZN(new_n14251_));
  NAND2_X1   g13934(.A1(new_n14102_), .A2(new_n14065_), .ZN(new_n14252_));
  NAND2_X1   g13935(.A1(new_n14252_), .A2(new_n14100_), .ZN(new_n14253_));
  XNOR2_X1   g13936(.A1(new_n14251_), .A2(new_n14253_), .ZN(new_n14254_));
  NAND2_X1   g13937(.A1(new_n14251_), .A2(new_n14253_), .ZN(new_n14255_));
  INV_X1     g13938(.I(new_n14255_), .ZN(new_n14256_));
  NOR2_X1    g13939(.A1(new_n14251_), .A2(new_n14253_), .ZN(new_n14257_));
  OAI21_X1   g13940(.A1(new_n14256_), .A2(new_n14257_), .B(new_n14238_), .ZN(new_n14258_));
  OAI21_X1   g13941(.A1(new_n14238_), .A2(new_n14254_), .B(new_n14258_), .ZN(new_n14259_));
  INV_X1     g13942(.I(new_n14259_), .ZN(new_n14260_));
  NOR2_X1    g13943(.A1(new_n14260_), .A2(new_n14234_), .ZN(new_n14261_));
  INV_X1     g13944(.I(new_n14261_), .ZN(new_n14262_));
  NAND2_X1   g13945(.A1(new_n14260_), .A2(new_n14234_), .ZN(new_n14263_));
  AOI21_X1   g13946(.A1(new_n14262_), .A2(new_n14263_), .B(new_n14232_), .ZN(new_n14264_));
  XNOR2_X1   g13947(.A1(new_n14234_), .A2(new_n14259_), .ZN(new_n14265_));
  AOI21_X1   g13948(.A1(new_n14232_), .A2(new_n14265_), .B(new_n14264_), .ZN(new_n14266_));
  NOR2_X1    g13949(.A1(new_n14114_), .A2(new_n13980_), .ZN(new_n14267_));
  NOR2_X1    g13950(.A1(new_n14267_), .A2(new_n14113_), .ZN(new_n14268_));
  XOR2_X1    g13951(.A1(new_n14266_), .A2(new_n14268_), .Z(new_n14269_));
  NAND2_X1   g13952(.A1(new_n14128_), .A2(new_n14269_), .ZN(new_n14270_));
  NOR2_X1    g13953(.A1(new_n14266_), .A2(new_n14268_), .ZN(new_n14271_));
  INV_X1     g13954(.I(new_n14271_), .ZN(new_n14272_));
  NAND2_X1   g13955(.A1(new_n14266_), .A2(new_n14268_), .ZN(new_n14273_));
  AND2_X2    g13956(.A1(new_n14272_), .A2(new_n14273_), .Z(new_n14274_));
  OAI21_X1   g13957(.A1(new_n14128_), .A2(new_n14274_), .B(new_n14270_), .ZN(\asquared[89] ));
  AOI21_X1   g13958(.A1(new_n14271_), .A2(new_n14118_), .B(new_n14122_), .ZN(new_n14276_));
  AOI21_X1   g13959(.A1(new_n14123_), .A2(new_n14272_), .B(new_n14276_), .ZN(new_n14277_));
  NAND2_X1   g13960(.A1(\asquared[87] ), .A2(new_n14277_), .ZN(new_n14278_));
  OAI21_X1   g13961(.A1(new_n14232_), .A2(new_n14261_), .B(new_n14263_), .ZN(new_n14279_));
  INV_X1     g13962(.I(new_n14279_), .ZN(new_n14280_));
  OAI21_X1   g13963(.A1(new_n14238_), .A2(new_n14257_), .B(new_n14255_), .ZN(new_n14281_));
  AOI21_X1   g13964(.A1(new_n14240_), .A2(new_n14249_), .B(new_n14247_), .ZN(new_n14282_));
  INV_X1     g13965(.I(new_n14139_), .ZN(new_n14283_));
  AOI21_X1   g13966(.A1(new_n14132_), .A2(new_n14283_), .B(new_n14138_), .ZN(new_n14284_));
  INV_X1     g13967(.I(new_n14284_), .ZN(new_n14285_));
  NOR2_X1    g13968(.A1(new_n1999_), .A2(new_n9310_), .ZN(new_n14286_));
  OAI21_X1   g13969(.A1(new_n14212_), .A2(new_n14215_), .B(new_n14286_), .ZN(new_n14287_));
  OAI21_X1   g13970(.A1(new_n14213_), .A2(new_n14216_), .B(new_n14287_), .ZN(new_n14288_));
  NAND2_X1   g13971(.A1(new_n14159_), .A2(new_n14150_), .ZN(new_n14289_));
  NAND2_X1   g13972(.A1(new_n14289_), .A2(new_n14156_), .ZN(new_n14290_));
  XOR2_X1    g13973(.A1(new_n14290_), .A2(new_n14288_), .Z(new_n14291_));
  NAND2_X1   g13974(.A1(new_n14291_), .A2(new_n14285_), .ZN(new_n14292_));
  AND2_X2    g13975(.A1(new_n14290_), .A2(new_n14288_), .Z(new_n14293_));
  NOR2_X1    g13976(.A1(new_n14290_), .A2(new_n14288_), .ZN(new_n14294_));
  OAI21_X1   g13977(.A1(new_n14293_), .A2(new_n14294_), .B(new_n14284_), .ZN(new_n14295_));
  NAND2_X1   g13978(.A1(new_n14292_), .A2(new_n14295_), .ZN(new_n14296_));
  AOI21_X1   g13979(.A1(new_n14142_), .A2(new_n14165_), .B(new_n14164_), .ZN(new_n14297_));
  XNOR2_X1   g13980(.A1(new_n14297_), .A2(new_n14296_), .ZN(new_n14298_));
  NOR2_X1    g13981(.A1(new_n14298_), .A2(new_n14282_), .ZN(new_n14299_));
  INV_X1     g13982(.I(new_n14282_), .ZN(new_n14300_));
  NOR2_X1    g13983(.A1(new_n14297_), .A2(new_n14296_), .ZN(new_n14301_));
  INV_X1     g13984(.I(new_n14301_), .ZN(new_n14302_));
  NAND2_X1   g13985(.A1(new_n14297_), .A2(new_n14296_), .ZN(new_n14303_));
  AOI21_X1   g13986(.A1(new_n14302_), .A2(new_n14303_), .B(new_n14300_), .ZN(new_n14304_));
  NOR2_X1    g13987(.A1(new_n14299_), .A2(new_n14304_), .ZN(new_n14305_));
  INV_X1     g13988(.I(new_n14305_), .ZN(new_n14306_));
  NAND2_X1   g13989(.A1(new_n3424_), .A2(new_n7421_), .ZN(new_n14307_));
  XNOR2_X1   g13990(.A1(new_n14307_), .A2(new_n7171_), .ZN(new_n14308_));
  AOI22_X1   g13991(.A1(new_n3805_), .A2(new_n7204_), .B1(new_n3838_), .B2(new_n7000_), .ZN(new_n14309_));
  NOR4_X1    g13992(.A1(new_n6777_), .A2(new_n5600_), .A3(new_n3393_), .A4(new_n6694_), .ZN(new_n14310_));
  NAND2_X1   g13993(.A1(new_n14309_), .A2(new_n14310_), .ZN(new_n14311_));
  AOI22_X1   g13994(.A1(new_n2766_), .A2(new_n8676_), .B1(new_n3126_), .B2(new_n8674_), .ZN(new_n14312_));
  INV_X1     g13995(.I(new_n14312_), .ZN(new_n14313_));
  NAND4_X1   g13996(.A1(new_n4184_), .A2(new_n8246_), .A3(\a[30] ), .A4(\a[59] ), .ZN(new_n14314_));
  NOR3_X1    g13997(.A1(new_n14311_), .A2(new_n14313_), .A3(new_n14314_), .ZN(new_n14315_));
  INV_X1     g13998(.I(new_n14311_), .ZN(new_n14316_));
  NOR2_X1    g13999(.A1(new_n14313_), .A2(new_n14314_), .ZN(new_n14317_));
  NOR2_X1    g14000(.A1(new_n14317_), .A2(new_n14316_), .ZN(new_n14318_));
  NOR2_X1    g14001(.A1(new_n14318_), .A2(new_n14315_), .ZN(new_n14319_));
  NOR2_X1    g14002(.A1(new_n14319_), .A2(new_n14308_), .ZN(new_n14320_));
  XOR2_X1    g14003(.A1(new_n14317_), .A2(new_n14316_), .Z(new_n14321_));
  AOI21_X1   g14004(.A1(new_n14308_), .A2(new_n14321_), .B(new_n14320_), .ZN(new_n14322_));
  AOI21_X1   g14005(.A1(new_n2797_), .A2(new_n8991_), .B(new_n14192_), .ZN(new_n14323_));
  AOI21_X1   g14006(.A1(new_n3838_), .A2(new_n6777_), .B(new_n14198_), .ZN(new_n14324_));
  AOI21_X1   g14007(.A1(new_n2766_), .A2(new_n14183_), .B(new_n7648_), .ZN(new_n14325_));
  XNOR2_X1   g14008(.A1(new_n14324_), .A2(new_n14325_), .ZN(new_n14326_));
  INV_X1     g14009(.I(new_n14324_), .ZN(new_n14327_));
  NOR2_X1    g14010(.A1(new_n14327_), .A2(new_n14325_), .ZN(new_n14328_));
  INV_X1     g14011(.I(new_n14328_), .ZN(new_n14329_));
  NAND2_X1   g14012(.A1(new_n14327_), .A2(new_n14325_), .ZN(new_n14330_));
  AOI21_X1   g14013(.A1(new_n14329_), .A2(new_n14330_), .B(new_n14323_), .ZN(new_n14331_));
  AOI21_X1   g14014(.A1(new_n14323_), .A2(new_n14326_), .B(new_n14331_), .ZN(new_n14332_));
  NAND2_X1   g14015(.A1(new_n5173_), .A2(new_n5980_), .ZN(new_n14333_));
  NAND2_X1   g14016(.A1(\a[34] ), .A2(\a[55] ), .ZN(new_n14334_));
  XNOR2_X1   g14017(.A1(new_n14333_), .A2(new_n14334_), .ZN(new_n14335_));
  INV_X1     g14018(.I(new_n14335_), .ZN(new_n14336_));
  AOI21_X1   g14019(.A1(new_n4372_), .A2(new_n7186_), .B(new_n7483_), .ZN(new_n14337_));
  NAND2_X1   g14020(.A1(\a[28] ), .A2(\a[60] ), .ZN(new_n14338_));
  NAND2_X1   g14021(.A1(\a[29] ), .A2(\a[61] ), .ZN(new_n14339_));
  XNOR2_X1   g14022(.A1(new_n14338_), .A2(new_n14339_), .ZN(new_n14340_));
  XOR2_X1    g14023(.A1(new_n14340_), .A2(new_n14337_), .Z(new_n14341_));
  NAND2_X1   g14024(.A1(\a[27] ), .A2(\a[45] ), .ZN(new_n14342_));
  XOR2_X1    g14025(.A1(new_n14214_), .A2(new_n14342_), .Z(new_n14343_));
  NOR2_X1    g14026(.A1(new_n14341_), .A2(new_n14343_), .ZN(new_n14344_));
  NAND2_X1   g14027(.A1(new_n14341_), .A2(new_n14343_), .ZN(new_n14345_));
  INV_X1     g14028(.I(new_n14345_), .ZN(new_n14346_));
  OAI21_X1   g14029(.A1(new_n14346_), .A2(new_n14344_), .B(new_n14336_), .ZN(new_n14347_));
  XNOR2_X1   g14030(.A1(new_n14341_), .A2(new_n14343_), .ZN(new_n14348_));
  OAI21_X1   g14031(.A1(new_n14336_), .A2(new_n14348_), .B(new_n14347_), .ZN(new_n14349_));
  NAND2_X1   g14032(.A1(new_n14332_), .A2(new_n14349_), .ZN(new_n14350_));
  NOR2_X1    g14033(.A1(new_n14332_), .A2(new_n14349_), .ZN(new_n14351_));
  INV_X1     g14034(.I(new_n14351_), .ZN(new_n14352_));
  AOI21_X1   g14035(.A1(new_n14352_), .A2(new_n14350_), .B(new_n14322_), .ZN(new_n14353_));
  XNOR2_X1   g14036(.A1(new_n14332_), .A2(new_n14349_), .ZN(new_n14354_));
  INV_X1     g14037(.I(new_n14354_), .ZN(new_n14355_));
  AOI21_X1   g14038(.A1(new_n14355_), .A2(new_n14322_), .B(new_n14353_), .ZN(new_n14356_));
  NOR2_X1    g14039(.A1(new_n14306_), .A2(new_n14356_), .ZN(new_n14357_));
  NAND2_X1   g14040(.A1(new_n14306_), .A2(new_n14356_), .ZN(new_n14358_));
  INV_X1     g14041(.I(new_n14358_), .ZN(new_n14359_));
  OAI21_X1   g14042(.A1(new_n14359_), .A2(new_n14357_), .B(new_n14281_), .ZN(new_n14360_));
  XOR2_X1    g14043(.A1(new_n14305_), .A2(new_n14356_), .Z(new_n14361_));
  OAI21_X1   g14044(.A1(new_n14281_), .A2(new_n14361_), .B(new_n14360_), .ZN(new_n14362_));
  NAND2_X1   g14045(.A1(new_n14228_), .A2(new_n14130_), .ZN(new_n14363_));
  NAND2_X1   g14046(.A1(new_n14363_), .A2(new_n14227_), .ZN(new_n14364_));
  NAND2_X1   g14047(.A1(new_n14175_), .A2(new_n14131_), .ZN(new_n14365_));
  NAND2_X1   g14048(.A1(new_n14365_), .A2(new_n14174_), .ZN(new_n14366_));
  INV_X1     g14049(.I(new_n14191_), .ZN(new_n14367_));
  OAI21_X1   g14050(.A1(new_n14367_), .A2(new_n14222_), .B(new_n14223_), .ZN(new_n14368_));
  AOI21_X1   g14051(.A1(new_n14179_), .A2(new_n14189_), .B(new_n14187_), .ZN(new_n14369_));
  INV_X1     g14052(.I(new_n14369_), .ZN(new_n14370_));
  NAND2_X1   g14053(.A1(new_n14203_), .A2(new_n14205_), .ZN(new_n14371_));
  NAND2_X1   g14054(.A1(new_n14371_), .A2(new_n14202_), .ZN(new_n14372_));
  NAND2_X1   g14055(.A1(new_n5350_), .A2(new_n5980_), .ZN(new_n14373_));
  NOR2_X1    g14056(.A1(new_n5350_), .A2(new_n5980_), .ZN(new_n14374_));
  NOR2_X1    g14057(.A1(\a[31] ), .A2(\a[57] ), .ZN(new_n14375_));
  AOI21_X1   g14058(.A1(new_n14373_), .A2(new_n14375_), .B(new_n14374_), .ZN(new_n14376_));
  NOR2_X1    g14059(.A1(new_n5339_), .A2(new_n6280_), .ZN(new_n14377_));
  NAND2_X1   g14060(.A1(new_n2499_), .A2(new_n8085_), .ZN(new_n14378_));
  AOI21_X1   g14061(.A1(new_n5339_), .A2(new_n6280_), .B(new_n14378_), .ZN(new_n14379_));
  NOR2_X1    g14062(.A1(new_n14379_), .A2(new_n14377_), .ZN(new_n14380_));
  INV_X1     g14063(.I(new_n14380_), .ZN(new_n14381_));
  NAND2_X1   g14064(.A1(\a[26] ), .A2(\a[63] ), .ZN(new_n14382_));
  AOI21_X1   g14065(.A1(new_n6280_), .A2(new_n6024_), .B(new_n14382_), .ZN(new_n14383_));
  NAND3_X1   g14066(.A1(new_n6280_), .A2(new_n6024_), .A3(new_n14382_), .ZN(new_n14384_));
  INV_X1     g14067(.I(new_n14384_), .ZN(new_n14385_));
  NOR2_X1    g14068(.A1(new_n14385_), .A2(new_n14383_), .ZN(new_n14386_));
  NOR2_X1    g14069(.A1(new_n14381_), .A2(new_n14386_), .ZN(new_n14387_));
  NOR3_X1    g14070(.A1(new_n14380_), .A2(new_n14383_), .A3(new_n14385_), .ZN(new_n14388_));
  NOR2_X1    g14071(.A1(new_n14387_), .A2(new_n14388_), .ZN(new_n14389_));
  XOR2_X1    g14072(.A1(new_n14386_), .A2(new_n14380_), .Z(new_n14390_));
  MUX2_X1    g14073(.I0(new_n14390_), .I1(new_n14389_), .S(new_n14376_), .Z(new_n14391_));
  XNOR2_X1   g14074(.A1(new_n14391_), .A2(new_n14372_), .ZN(new_n14392_));
  NAND2_X1   g14075(.A1(new_n14392_), .A2(new_n14370_), .ZN(new_n14393_));
  INV_X1     g14076(.I(new_n14372_), .ZN(new_n14394_));
  NOR2_X1    g14077(.A1(new_n14394_), .A2(new_n14391_), .ZN(new_n14395_));
  NAND2_X1   g14078(.A1(new_n14394_), .A2(new_n14391_), .ZN(new_n14396_));
  INV_X1     g14079(.I(new_n14396_), .ZN(new_n14397_));
  OAI21_X1   g14080(.A1(new_n14397_), .A2(new_n14395_), .B(new_n14369_), .ZN(new_n14398_));
  NAND2_X1   g14081(.A1(new_n14393_), .A2(new_n14398_), .ZN(new_n14399_));
  XNOR2_X1   g14082(.A1(new_n14368_), .A2(new_n14399_), .ZN(new_n14400_));
  INV_X1     g14083(.I(new_n14399_), .ZN(new_n14401_));
  NOR2_X1    g14084(.A1(new_n14401_), .A2(new_n14368_), .ZN(new_n14402_));
  NAND2_X1   g14085(.A1(new_n14401_), .A2(new_n14368_), .ZN(new_n14403_));
  INV_X1     g14086(.I(new_n14403_), .ZN(new_n14404_));
  NOR2_X1    g14087(.A1(new_n14404_), .A2(new_n14402_), .ZN(new_n14405_));
  NOR2_X1    g14088(.A1(new_n14366_), .A2(new_n14405_), .ZN(new_n14406_));
  AOI21_X1   g14089(.A1(new_n14366_), .A2(new_n14400_), .B(new_n14406_), .ZN(new_n14407_));
  XOR2_X1    g14090(.A1(new_n14364_), .A2(new_n14407_), .Z(new_n14408_));
  NOR2_X1    g14091(.A1(new_n14364_), .A2(new_n14407_), .ZN(new_n14409_));
  INV_X1     g14092(.I(new_n14409_), .ZN(new_n14410_));
  NAND2_X1   g14093(.A1(new_n14364_), .A2(new_n14407_), .ZN(new_n14411_));
  AOI21_X1   g14094(.A1(new_n14410_), .A2(new_n14411_), .B(new_n14362_), .ZN(new_n14412_));
  AOI21_X1   g14095(.A1(new_n14362_), .A2(new_n14408_), .B(new_n14412_), .ZN(new_n14413_));
  NOR2_X1    g14096(.A1(new_n14413_), .A2(new_n14280_), .ZN(new_n14414_));
  XOR2_X1    g14097(.A1(new_n14278_), .A2(new_n14414_), .Z(new_n14415_));
  XOR2_X1    g14098(.A1(new_n14415_), .A2(new_n14273_), .Z(\asquared[90] ));
  INV_X1     g14099(.I(new_n14414_), .ZN(new_n14417_));
  AOI21_X1   g14100(.A1(new_n13492_), .A2(new_n13490_), .B(new_n13826_), .ZN(new_n14418_));
  AOI21_X1   g14101(.A1(new_n14413_), .A2(new_n14280_), .B(new_n14273_), .ZN(new_n14419_));
  NAND4_X1   g14102(.A1(new_n14418_), .A2(new_n13820_), .A3(new_n14277_), .A4(new_n14419_), .ZN(new_n14420_));
  AND2_X2    g14103(.A1(new_n14420_), .A2(new_n14417_), .Z(new_n14421_));
  NAND2_X1   g14104(.A1(new_n14410_), .A2(new_n14362_), .ZN(new_n14422_));
  AND2_X2    g14105(.A1(new_n14422_), .A2(new_n14411_), .Z(new_n14423_));
  AOI21_X1   g14106(.A1(new_n14281_), .A2(new_n14358_), .B(new_n14357_), .ZN(new_n14424_));
  AOI21_X1   g14107(.A1(new_n14365_), .A2(new_n14174_), .B(new_n14402_), .ZN(new_n14425_));
  NOR2_X1    g14108(.A1(new_n14425_), .A2(new_n14404_), .ZN(new_n14426_));
  NOR2_X1    g14109(.A1(new_n14284_), .A2(new_n14294_), .ZN(new_n14427_));
  NOR2_X1    g14110(.A1(new_n14427_), .A2(new_n14293_), .ZN(new_n14428_));
  OAI22_X1   g14111(.A1(new_n7023_), .A2(new_n5174_), .B1(new_n7693_), .B2(new_n8199_), .ZN(new_n14429_));
  OAI21_X1   g14112(.A1(new_n5322_), .A2(new_n5793_), .B(new_n14429_), .ZN(new_n14430_));
  INV_X1     g14113(.I(new_n14430_), .ZN(new_n14431_));
  AOI21_X1   g14114(.A1(new_n14431_), .A2(new_n7452_), .B(\a[47] ), .ZN(new_n14432_));
  NOR2_X1    g14115(.A1(\a[42] ), .A2(\a[48] ), .ZN(new_n14433_));
  OAI21_X1   g14116(.A1(new_n14432_), .A2(new_n4501_), .B(new_n14433_), .ZN(new_n14434_));
  AOI21_X1   g14117(.A1(new_n5321_), .A2(new_n5980_), .B(new_n14429_), .ZN(new_n14435_));
  NAND2_X1   g14118(.A1(new_n14434_), .A2(new_n14435_), .ZN(new_n14436_));
  AOI21_X1   g14119(.A1(new_n8755_), .A2(new_n10958_), .B(new_n7008_), .ZN(new_n14437_));
  NOR4_X1    g14120(.A1(new_n4372_), .A2(new_n8242_), .A3(new_n3423_), .A4(new_n6999_), .ZN(new_n14438_));
  NAND2_X1   g14121(.A1(new_n14437_), .A2(new_n14438_), .ZN(new_n14439_));
  AOI21_X1   g14122(.A1(new_n3805_), .A2(new_n3838_), .B(new_n10291_), .ZN(new_n14440_));
  INV_X1     g14123(.I(new_n14440_), .ZN(new_n14441_));
  NOR2_X1    g14124(.A1(new_n8056_), .A2(new_n4706_), .ZN(new_n14442_));
  AOI21_X1   g14125(.A1(\a[38] ), .A2(\a[52] ), .B(new_n7205_), .ZN(new_n14443_));
  OR4_X2     g14126(.A1(new_n3393_), .A2(new_n14442_), .A3(new_n6945_), .A4(new_n14443_), .Z(new_n14444_));
  NOR2_X1    g14127(.A1(new_n14441_), .A2(new_n14444_), .ZN(new_n14445_));
  INV_X1     g14128(.I(new_n14445_), .ZN(new_n14446_));
  NOR2_X1    g14129(.A1(new_n14446_), .A2(new_n14439_), .ZN(new_n14447_));
  AOI21_X1   g14130(.A1(new_n14437_), .A2(new_n14438_), .B(new_n14445_), .ZN(new_n14448_));
  NOR2_X1    g14131(.A1(new_n14447_), .A2(new_n14448_), .ZN(new_n14449_));
  NOR2_X1    g14132(.A1(new_n14436_), .A2(new_n14449_), .ZN(new_n14450_));
  INV_X1     g14133(.I(new_n14436_), .ZN(new_n14451_));
  XOR2_X1    g14134(.A1(new_n14445_), .A2(new_n14439_), .Z(new_n14452_));
  NOR2_X1    g14135(.A1(new_n14451_), .A2(new_n14452_), .ZN(new_n14453_));
  NOR2_X1    g14136(.A1(new_n14453_), .A2(new_n14450_), .ZN(new_n14454_));
  AOI21_X1   g14137(.A1(new_n5600_), .A2(new_n6777_), .B(new_n14309_), .ZN(new_n14455_));
  AOI21_X1   g14138(.A1(new_n3981_), .A2(new_n8245_), .B(new_n14312_), .ZN(new_n14456_));
  NAND2_X1   g14139(.A1(new_n6280_), .A2(new_n6024_), .ZN(new_n14457_));
  NOR2_X1    g14140(.A1(new_n6280_), .A2(new_n6024_), .ZN(new_n14458_));
  NOR2_X1    g14141(.A1(\a[26] ), .A2(\a[63] ), .ZN(new_n14459_));
  AOI21_X1   g14142(.A1(new_n14457_), .A2(new_n14459_), .B(new_n14458_), .ZN(new_n14460_));
  XNOR2_X1   g14143(.A1(new_n14456_), .A2(new_n14460_), .ZN(new_n14461_));
  INV_X1     g14144(.I(new_n14456_), .ZN(new_n14462_));
  INV_X1     g14145(.I(new_n14460_), .ZN(new_n14463_));
  NOR2_X1    g14146(.A1(new_n14462_), .A2(new_n14463_), .ZN(new_n14464_));
  NOR2_X1    g14147(.A1(new_n14456_), .A2(new_n14460_), .ZN(new_n14465_));
  NOR2_X1    g14148(.A1(new_n14464_), .A2(new_n14465_), .ZN(new_n14466_));
  MUX2_X1    g14149(.I0(new_n14466_), .I1(new_n14461_), .S(new_n14455_), .Z(new_n14467_));
  XOR2_X1    g14150(.A1(new_n14454_), .A2(new_n14467_), .Z(new_n14468_));
  NOR2_X1    g14151(.A1(new_n14468_), .A2(new_n14428_), .ZN(new_n14469_));
  INV_X1     g14152(.I(new_n14428_), .ZN(new_n14470_));
  INV_X1     g14153(.I(new_n14454_), .ZN(new_n14471_));
  NOR2_X1    g14154(.A1(new_n14471_), .A2(new_n14467_), .ZN(new_n14472_));
  INV_X1     g14155(.I(new_n14472_), .ZN(new_n14473_));
  NAND2_X1   g14156(.A1(new_n14471_), .A2(new_n14467_), .ZN(new_n14474_));
  AOI21_X1   g14157(.A1(new_n14473_), .A2(new_n14474_), .B(new_n14470_), .ZN(new_n14475_));
  NOR2_X1    g14158(.A1(new_n14475_), .A2(new_n14469_), .ZN(new_n14476_));
  AOI21_X1   g14159(.A1(new_n14370_), .A2(new_n14396_), .B(new_n14395_), .ZN(new_n14477_));
  AOI21_X1   g14160(.A1(new_n14323_), .A2(new_n14330_), .B(new_n14328_), .ZN(new_n14478_));
  INV_X1     g14161(.I(new_n14388_), .ZN(new_n14479_));
  AOI21_X1   g14162(.A1(new_n14479_), .A2(new_n14376_), .B(new_n14387_), .ZN(new_n14480_));
  NOR2_X1    g14163(.A1(new_n12545_), .A2(new_n13707_), .ZN(new_n14481_));
  INV_X1     g14164(.I(new_n14481_), .ZN(new_n14482_));
  NOR4_X1    g14165(.A1(new_n14482_), .A2(new_n5592_), .A3(new_n6280_), .A4(new_n7462_), .ZN(new_n14483_));
  XOR2_X1    g14166(.A1(new_n14480_), .A2(new_n14483_), .Z(new_n14484_));
  NOR2_X1    g14167(.A1(new_n14484_), .A2(new_n14478_), .ZN(new_n14485_));
  INV_X1     g14168(.I(new_n14483_), .ZN(new_n14486_));
  NOR2_X1    g14169(.A1(new_n14486_), .A2(new_n14480_), .ZN(new_n14487_));
  INV_X1     g14170(.I(new_n14487_), .ZN(new_n14488_));
  NAND2_X1   g14171(.A1(new_n14486_), .A2(new_n14480_), .ZN(new_n14489_));
  NAND2_X1   g14172(.A1(new_n14488_), .A2(new_n14489_), .ZN(new_n14490_));
  AOI21_X1   g14173(.A1(new_n14478_), .A2(new_n14490_), .B(new_n14485_), .ZN(new_n14491_));
  NOR2_X1    g14174(.A1(new_n13620_), .A2(new_n9042_), .ZN(new_n14492_));
  NOR2_X1    g14175(.A1(new_n2098_), .A2(new_n9310_), .ZN(new_n14493_));
  NAND4_X1   g14176(.A1(new_n14492_), .A2(new_n2689_), .A3(new_n9785_), .A4(new_n14493_), .ZN(new_n14494_));
  INV_X1     g14177(.I(new_n14337_), .ZN(new_n14495_));
  INV_X1     g14178(.I(new_n14340_), .ZN(new_n14496_));
  AOI22_X1   g14179(.A1(new_n14496_), .A2(new_n8991_), .B1(new_n2690_), .B2(new_n14495_), .ZN(new_n14497_));
  INV_X1     g14180(.I(new_n14497_), .ZN(new_n14498_));
  NOR2_X1    g14181(.A1(new_n9556_), .A2(new_n13071_), .ZN(new_n14499_));
  INV_X1     g14182(.I(new_n14499_), .ZN(new_n14500_));
  NOR2_X1    g14183(.A1(new_n2655_), .A2(new_n7647_), .ZN(new_n14501_));
  OAI22_X1   g14184(.A1(new_n8087_), .A2(new_n14501_), .B1(new_n2461_), .B2(new_n8990_), .ZN(new_n14502_));
  AOI21_X1   g14185(.A1(new_n8087_), .A2(new_n14501_), .B(new_n14502_), .ZN(new_n14503_));
  AOI21_X1   g14186(.A1(new_n14500_), .A2(new_n14503_), .B(new_n8676_), .ZN(new_n14504_));
  NOR2_X1    g14187(.A1(new_n14504_), .A2(new_n4184_), .ZN(new_n14505_));
  XOR2_X1    g14188(.A1(new_n14505_), .A2(new_n14498_), .Z(new_n14506_));
  NOR2_X1    g14189(.A1(new_n14506_), .A2(new_n14494_), .ZN(new_n14507_));
  INV_X1     g14190(.I(new_n14494_), .ZN(new_n14508_));
  NOR3_X1    g14191(.A1(new_n14504_), .A2(new_n14498_), .A3(new_n4184_), .ZN(new_n14509_));
  NOR2_X1    g14192(.A1(new_n14505_), .A2(new_n14497_), .ZN(new_n14510_));
  NOR2_X1    g14193(.A1(new_n14510_), .A2(new_n14509_), .ZN(new_n14511_));
  NOR2_X1    g14194(.A1(new_n14511_), .A2(new_n14508_), .ZN(new_n14512_));
  NOR2_X1    g14195(.A1(new_n14507_), .A2(new_n14512_), .ZN(new_n14513_));
  NOR2_X1    g14196(.A1(new_n14491_), .A2(new_n14513_), .ZN(new_n14514_));
  INV_X1     g14197(.I(new_n14514_), .ZN(new_n14515_));
  NAND2_X1   g14198(.A1(new_n14491_), .A2(new_n14513_), .ZN(new_n14516_));
  AOI21_X1   g14199(.A1(new_n14515_), .A2(new_n14516_), .B(new_n14477_), .ZN(new_n14517_));
  INV_X1     g14200(.I(new_n14477_), .ZN(new_n14518_));
  XNOR2_X1   g14201(.A1(new_n14491_), .A2(new_n14513_), .ZN(new_n14519_));
  NOR2_X1    g14202(.A1(new_n14519_), .A2(new_n14518_), .ZN(new_n14520_));
  OAI21_X1   g14203(.A1(new_n14517_), .A2(new_n14520_), .B(new_n14476_), .ZN(new_n14521_));
  NOR2_X1    g14204(.A1(new_n14520_), .A2(new_n14517_), .ZN(new_n14522_));
  OAI21_X1   g14205(.A1(new_n14469_), .A2(new_n14475_), .B(new_n14522_), .ZN(new_n14523_));
  AOI21_X1   g14206(.A1(new_n14521_), .A2(new_n14523_), .B(new_n14426_), .ZN(new_n14524_));
  XNOR2_X1   g14207(.A1(new_n14476_), .A2(new_n14522_), .ZN(new_n14525_));
  AOI21_X1   g14208(.A1(new_n14426_), .A2(new_n14525_), .B(new_n14524_), .ZN(new_n14526_));
  NAND2_X1   g14209(.A1(new_n14303_), .A2(new_n14300_), .ZN(new_n14527_));
  NAND2_X1   g14210(.A1(new_n14527_), .A2(new_n14302_), .ZN(new_n14528_));
  OAI21_X1   g14211(.A1(new_n14322_), .A2(new_n14351_), .B(new_n14350_), .ZN(new_n14529_));
  NAND2_X1   g14212(.A1(new_n3424_), .A2(new_n7421_), .ZN(new_n14530_));
  NOR2_X1    g14213(.A1(new_n3424_), .A2(new_n7421_), .ZN(new_n14531_));
  NOR2_X1    g14214(.A1(\a[41] ), .A2(\a[48] ), .ZN(new_n14532_));
  AOI21_X1   g14215(.A1(new_n14530_), .A2(new_n14532_), .B(new_n14531_), .ZN(new_n14533_));
  INV_X1     g14216(.I(new_n14533_), .ZN(new_n14534_));
  NOR2_X1    g14217(.A1(new_n5173_), .A2(new_n5980_), .ZN(new_n14535_));
  NAND2_X1   g14218(.A1(new_n3371_), .A2(new_n6999_), .ZN(new_n14536_));
  AOI21_X1   g14219(.A1(new_n5173_), .A2(new_n5980_), .B(new_n14536_), .ZN(new_n14537_));
  NOR2_X1    g14220(.A1(new_n14537_), .A2(new_n14535_), .ZN(new_n14538_));
  NOR2_X1    g14221(.A1(new_n5004_), .A2(new_n9029_), .ZN(new_n14539_));
  AOI21_X1   g14222(.A1(\a[27] ), .A2(new_n14539_), .B(new_n5742_), .ZN(new_n14540_));
  INV_X1     g14223(.I(new_n14540_), .ZN(new_n14541_));
  XOR2_X1    g14224(.A1(new_n14538_), .A2(new_n14541_), .Z(new_n14542_));
  NOR2_X1    g14225(.A1(new_n14542_), .A2(new_n14534_), .ZN(new_n14543_));
  INV_X1     g14226(.I(new_n14538_), .ZN(new_n14544_));
  NOR2_X1    g14227(.A1(new_n14544_), .A2(new_n14541_), .ZN(new_n14545_));
  NOR2_X1    g14228(.A1(new_n14538_), .A2(new_n14540_), .ZN(new_n14546_));
  NOR2_X1    g14229(.A1(new_n14545_), .A2(new_n14546_), .ZN(new_n14547_));
  NOR2_X1    g14230(.A1(new_n14547_), .A2(new_n14533_), .ZN(new_n14548_));
  NOR2_X1    g14231(.A1(new_n14548_), .A2(new_n14543_), .ZN(new_n14549_));
  AOI21_X1   g14232(.A1(new_n14336_), .A2(new_n14345_), .B(new_n14344_), .ZN(new_n14550_));
  INV_X1     g14233(.I(new_n14315_), .ZN(new_n14551_));
  OAI21_X1   g14234(.A1(new_n14308_), .A2(new_n14318_), .B(new_n14551_), .ZN(new_n14552_));
  INV_X1     g14235(.I(new_n14552_), .ZN(new_n14553_));
  NOR2_X1    g14236(.A1(new_n14553_), .A2(new_n14550_), .ZN(new_n14554_));
  INV_X1     g14237(.I(new_n14554_), .ZN(new_n14555_));
  NAND2_X1   g14238(.A1(new_n14553_), .A2(new_n14550_), .ZN(new_n14556_));
  AOI21_X1   g14239(.A1(new_n14555_), .A2(new_n14556_), .B(new_n14549_), .ZN(new_n14557_));
  XOR2_X1    g14240(.A1(new_n14550_), .A2(new_n14552_), .Z(new_n14558_));
  INV_X1     g14241(.I(new_n14558_), .ZN(new_n14559_));
  AOI21_X1   g14242(.A1(new_n14559_), .A2(new_n14549_), .B(new_n14557_), .ZN(new_n14560_));
  XOR2_X1    g14243(.A1(new_n14529_), .A2(new_n14560_), .Z(new_n14561_));
  NAND2_X1   g14244(.A1(new_n14528_), .A2(new_n14561_), .ZN(new_n14562_));
  NOR2_X1    g14245(.A1(new_n14529_), .A2(new_n14560_), .ZN(new_n14563_));
  NAND2_X1   g14246(.A1(new_n14529_), .A2(new_n14560_), .ZN(new_n14564_));
  INV_X1     g14247(.I(new_n14564_), .ZN(new_n14565_));
  NOR2_X1    g14248(.A1(new_n14565_), .A2(new_n14563_), .ZN(new_n14566_));
  OAI21_X1   g14249(.A1(new_n14528_), .A2(new_n14566_), .B(new_n14562_), .ZN(new_n14567_));
  XNOR2_X1   g14250(.A1(new_n14526_), .A2(new_n14567_), .ZN(new_n14568_));
  NOR2_X1    g14251(.A1(new_n14568_), .A2(new_n14424_), .ZN(new_n14569_));
  INV_X1     g14252(.I(new_n14424_), .ZN(new_n14570_));
  NAND2_X1   g14253(.A1(new_n14526_), .A2(new_n14567_), .ZN(new_n14571_));
  NOR2_X1    g14254(.A1(new_n14526_), .A2(new_n14567_), .ZN(new_n14572_));
  INV_X1     g14255(.I(new_n14572_), .ZN(new_n14573_));
  AOI21_X1   g14256(.A1(new_n14573_), .A2(new_n14571_), .B(new_n14570_), .ZN(new_n14574_));
  NOR2_X1    g14257(.A1(new_n14569_), .A2(new_n14574_), .ZN(new_n14575_));
  XOR2_X1    g14258(.A1(new_n14423_), .A2(new_n14575_), .Z(new_n14576_));
  INV_X1     g14259(.I(new_n14575_), .ZN(new_n14577_));
  AND2_X2    g14260(.A1(new_n14423_), .A2(new_n14577_), .Z(new_n14578_));
  NOR2_X1    g14261(.A1(new_n14423_), .A2(new_n14577_), .ZN(new_n14579_));
  OAI21_X1   g14262(.A1(new_n14578_), .A2(new_n14579_), .B(new_n14421_), .ZN(new_n14580_));
  OAI21_X1   g14263(.A1(new_n14421_), .A2(new_n14576_), .B(new_n14580_), .ZN(\asquared[91] ));
  INV_X1     g14264(.I(new_n14579_), .ZN(new_n14582_));
  AOI21_X1   g14265(.A1(new_n14421_), .A2(new_n14582_), .B(new_n14578_), .ZN(new_n14583_));
  NAND2_X1   g14266(.A1(new_n14571_), .A2(new_n14570_), .ZN(new_n14584_));
  NAND2_X1   g14267(.A1(new_n14584_), .A2(new_n14573_), .ZN(new_n14585_));
  INV_X1     g14268(.I(new_n14563_), .ZN(new_n14586_));
  AOI21_X1   g14269(.A1(new_n14528_), .A2(new_n14586_), .B(new_n14565_), .ZN(new_n14587_));
  INV_X1     g14270(.I(new_n14478_), .ZN(new_n14588_));
  AOI21_X1   g14271(.A1(new_n14588_), .A2(new_n14489_), .B(new_n14487_), .ZN(new_n14589_));
  AOI21_X1   g14272(.A1(new_n2690_), .A2(new_n9784_), .B(new_n14492_), .ZN(new_n14590_));
  AOI21_X1   g14273(.A1(new_n3981_), .A2(new_n8676_), .B(new_n14499_), .ZN(new_n14591_));
  XNOR2_X1   g14274(.A1(new_n14591_), .A2(new_n14590_), .ZN(new_n14592_));
  NOR3_X1    g14275(.A1(new_n14592_), .A2(new_n14440_), .A3(new_n14442_), .ZN(new_n14593_));
  NOR2_X1    g14276(.A1(new_n14440_), .A2(new_n14442_), .ZN(new_n14594_));
  INV_X1     g14277(.I(new_n14590_), .ZN(new_n14595_));
  INV_X1     g14278(.I(new_n14591_), .ZN(new_n14596_));
  NOR2_X1    g14279(.A1(new_n14596_), .A2(new_n14595_), .ZN(new_n14597_));
  NOR2_X1    g14280(.A1(new_n14591_), .A2(new_n14590_), .ZN(new_n14598_));
  NOR2_X1    g14281(.A1(new_n14597_), .A2(new_n14598_), .ZN(new_n14599_));
  NOR2_X1    g14282(.A1(new_n14599_), .A2(new_n14594_), .ZN(new_n14600_));
  NOR2_X1    g14283(.A1(new_n14593_), .A2(new_n14600_), .ZN(new_n14601_));
  NAND2_X1   g14284(.A1(new_n5592_), .A2(new_n6779_), .ZN(new_n14602_));
  NAND2_X1   g14285(.A1(\a[28] ), .A2(\a[63] ), .ZN(new_n14603_));
  XNOR2_X1   g14286(.A1(new_n14602_), .A2(new_n14603_), .ZN(new_n14604_));
  NAND2_X1   g14287(.A1(new_n5321_), .A2(new_n6030_), .ZN(new_n14605_));
  NAND2_X1   g14288(.A1(\a[35] ), .A2(\a[56] ), .ZN(new_n14606_));
  XNOR2_X1   g14289(.A1(new_n14605_), .A2(new_n14606_), .ZN(new_n14607_));
  NAND2_X1   g14290(.A1(\a[29] ), .A2(\a[46] ), .ZN(new_n14608_));
  XOR2_X1    g14291(.A1(new_n14539_), .A2(new_n14608_), .Z(new_n14609_));
  NOR2_X1    g14292(.A1(new_n14607_), .A2(new_n14609_), .ZN(new_n14610_));
  AND2_X2    g14293(.A1(new_n14607_), .A2(new_n14609_), .Z(new_n14611_));
  NOR2_X1    g14294(.A1(new_n14611_), .A2(new_n14610_), .ZN(new_n14612_));
  NOR2_X1    g14295(.A1(new_n14612_), .A2(new_n14604_), .ZN(new_n14613_));
  INV_X1     g14296(.I(new_n14604_), .ZN(new_n14614_));
  XNOR2_X1   g14297(.A1(new_n14607_), .A2(new_n14609_), .ZN(new_n14615_));
  NOR2_X1    g14298(.A1(new_n14615_), .A2(new_n14614_), .ZN(new_n14616_));
  NOR2_X1    g14299(.A1(new_n14613_), .A2(new_n14616_), .ZN(new_n14617_));
  XOR2_X1    g14300(.A1(new_n14601_), .A2(new_n14617_), .Z(new_n14618_));
  NOR2_X1    g14301(.A1(new_n14618_), .A2(new_n14589_), .ZN(new_n14619_));
  INV_X1     g14302(.I(new_n14589_), .ZN(new_n14620_));
  INV_X1     g14303(.I(new_n14601_), .ZN(new_n14621_));
  NOR2_X1    g14304(.A1(new_n14621_), .A2(new_n14617_), .ZN(new_n14622_));
  INV_X1     g14305(.I(new_n14622_), .ZN(new_n14623_));
  NAND2_X1   g14306(.A1(new_n14621_), .A2(new_n14617_), .ZN(new_n14624_));
  AOI21_X1   g14307(.A1(new_n14623_), .A2(new_n14624_), .B(new_n14620_), .ZN(new_n14625_));
  NOR2_X1    g14308(.A1(new_n14625_), .A2(new_n14619_), .ZN(new_n14626_));
  INV_X1     g14309(.I(new_n14546_), .ZN(new_n14627_));
  AOI21_X1   g14310(.A1(new_n14533_), .A2(new_n14627_), .B(new_n14545_), .ZN(new_n14628_));
  INV_X1     g14311(.I(new_n14465_), .ZN(new_n14629_));
  AOI21_X1   g14312(.A1(new_n14455_), .A2(new_n14629_), .B(new_n14464_), .ZN(new_n14630_));
  NAND2_X1   g14313(.A1(\a[55] ), .A2(\a[57] ), .ZN(new_n14631_));
  XOR2_X1    g14314(.A1(new_n4727_), .A2(new_n14631_), .Z(new_n14632_));
  XNOR2_X1   g14315(.A1(new_n14630_), .A2(new_n14632_), .ZN(new_n14633_));
  NOR2_X1    g14316(.A1(new_n14633_), .A2(new_n14628_), .ZN(new_n14634_));
  INV_X1     g14317(.I(new_n14628_), .ZN(new_n14635_));
  NOR2_X1    g14318(.A1(new_n14630_), .A2(new_n14632_), .ZN(new_n14636_));
  INV_X1     g14319(.I(new_n14636_), .ZN(new_n14637_));
  NAND2_X1   g14320(.A1(new_n14630_), .A2(new_n14632_), .ZN(new_n14638_));
  AOI21_X1   g14321(.A1(new_n14637_), .A2(new_n14638_), .B(new_n14635_), .ZN(new_n14639_));
  NOR2_X1    g14322(.A1(new_n14634_), .A2(new_n14639_), .ZN(new_n14640_));
  NAND2_X1   g14323(.A1(new_n14556_), .A2(new_n14549_), .ZN(new_n14641_));
  NAND2_X1   g14324(.A1(new_n14641_), .A2(new_n14555_), .ZN(new_n14642_));
  INV_X1     g14325(.I(new_n14642_), .ZN(new_n14643_));
  AOI21_X1   g14326(.A1(new_n5592_), .A2(new_n6280_), .B(new_n14481_), .ZN(new_n14644_));
  INV_X1     g14327(.I(new_n14644_), .ZN(new_n14645_));
  NOR2_X1    g14328(.A1(new_n9556_), .A2(new_n11541_), .ZN(new_n14646_));
  NOR4_X1    g14329(.A1(new_n3851_), .A2(new_n8676_), .A3(new_n2655_), .A4(new_n8990_), .ZN(new_n14647_));
  NAND2_X1   g14330(.A1(new_n14646_), .A2(new_n14647_), .ZN(new_n14648_));
  AOI22_X1   g14331(.A1(new_n5601_), .A2(new_n7482_), .B1(new_n10289_), .B2(new_n5600_), .ZN(new_n14649_));
  NOR4_X1    g14332(.A1(new_n5339_), .A2(new_n7204_), .A3(new_n3837_), .A4(new_n6945_), .ZN(new_n14650_));
  NAND2_X1   g14333(.A1(new_n14649_), .A2(new_n14650_), .ZN(new_n14651_));
  NOR2_X1    g14334(.A1(new_n14648_), .A2(new_n14651_), .ZN(new_n14652_));
  AOI22_X1   g14335(.A1(new_n14646_), .A2(new_n14647_), .B1(new_n14649_), .B2(new_n14650_), .ZN(new_n14653_));
  NOR2_X1    g14336(.A1(new_n14652_), .A2(new_n14653_), .ZN(new_n14654_));
  NOR2_X1    g14337(.A1(new_n14654_), .A2(new_n14645_), .ZN(new_n14655_));
  XOR2_X1    g14338(.A1(new_n14648_), .A2(new_n14651_), .Z(new_n14656_));
  AOI21_X1   g14339(.A1(new_n14656_), .A2(new_n14645_), .B(new_n14655_), .ZN(new_n14657_));
  NOR2_X1    g14340(.A1(new_n14643_), .A2(new_n14657_), .ZN(new_n14658_));
  INV_X1     g14341(.I(new_n14658_), .ZN(new_n14659_));
  NAND2_X1   g14342(.A1(new_n14643_), .A2(new_n14657_), .ZN(new_n14660_));
  AOI21_X1   g14343(.A1(new_n14659_), .A2(new_n14660_), .B(new_n14640_), .ZN(new_n14661_));
  XOR2_X1    g14344(.A1(new_n14642_), .A2(new_n14657_), .Z(new_n14662_));
  NOR3_X1    g14345(.A1(new_n14662_), .A2(new_n14634_), .A3(new_n14639_), .ZN(new_n14663_));
  NOR2_X1    g14346(.A1(new_n14661_), .A2(new_n14663_), .ZN(new_n14664_));
  NOR2_X1    g14347(.A1(new_n14664_), .A2(new_n14626_), .ZN(new_n14665_));
  NOR4_X1    g14348(.A1(new_n14661_), .A2(new_n14663_), .A3(new_n14619_), .A4(new_n14625_), .ZN(new_n14666_));
  NOR2_X1    g14349(.A1(new_n14665_), .A2(new_n14666_), .ZN(new_n14667_));
  NOR2_X1    g14350(.A1(new_n14587_), .A2(new_n14667_), .ZN(new_n14668_));
  XOR2_X1    g14351(.A1(new_n14664_), .A2(new_n14626_), .Z(new_n14669_));
  AOI21_X1   g14352(.A1(new_n14669_), .A2(new_n14587_), .B(new_n14668_), .ZN(new_n14670_));
  OAI21_X1   g14353(.A1(new_n14425_), .A2(new_n14404_), .B(new_n14523_), .ZN(new_n14671_));
  NAND2_X1   g14354(.A1(new_n14671_), .A2(new_n14521_), .ZN(new_n14672_));
  OAI21_X1   g14355(.A1(new_n14477_), .A2(new_n14514_), .B(new_n14516_), .ZN(new_n14673_));
  INV_X1     g14356(.I(new_n14673_), .ZN(new_n14674_));
  OAI21_X1   g14357(.A1(new_n14428_), .A2(new_n14472_), .B(new_n14474_), .ZN(new_n14675_));
  INV_X1     g14358(.I(new_n14448_), .ZN(new_n14676_));
  AOI21_X1   g14359(.A1(new_n14451_), .A2(new_n14676_), .B(new_n14447_), .ZN(new_n14677_));
  AOI21_X1   g14360(.A1(new_n4372_), .A2(new_n8242_), .B(new_n14437_), .ZN(new_n14678_));
  INV_X1     g14361(.I(new_n14678_), .ZN(new_n14679_));
  NOR2_X1    g14362(.A1(new_n14679_), .A2(new_n14430_), .ZN(new_n14680_));
  XOR2_X1    g14363(.A1(new_n14680_), .A2(new_n2461_), .Z(new_n14681_));
  XOR2_X1    g14364(.A1(new_n14681_), .A2(\a[61] ), .Z(new_n14682_));
  NOR2_X1    g14365(.A1(new_n14509_), .A2(new_n14494_), .ZN(new_n14683_));
  NOR2_X1    g14366(.A1(new_n14683_), .A2(new_n14510_), .ZN(new_n14684_));
  XOR2_X1    g14367(.A1(new_n14682_), .A2(new_n14684_), .Z(new_n14685_));
  NOR2_X1    g14368(.A1(new_n14685_), .A2(new_n14677_), .ZN(new_n14686_));
  INV_X1     g14369(.I(new_n14677_), .ZN(new_n14687_));
  INV_X1     g14370(.I(new_n14682_), .ZN(new_n14688_));
  NOR2_X1    g14371(.A1(new_n14688_), .A2(new_n14684_), .ZN(new_n14689_));
  INV_X1     g14372(.I(new_n14689_), .ZN(new_n14690_));
  NAND2_X1   g14373(.A1(new_n14688_), .A2(new_n14684_), .ZN(new_n14691_));
  AOI21_X1   g14374(.A1(new_n14690_), .A2(new_n14691_), .B(new_n14687_), .ZN(new_n14692_));
  NOR2_X1    g14375(.A1(new_n14692_), .A2(new_n14686_), .ZN(new_n14693_));
  NOR2_X1    g14376(.A1(new_n14693_), .A2(new_n14675_), .ZN(new_n14694_));
  INV_X1     g14377(.I(new_n14694_), .ZN(new_n14695_));
  NAND2_X1   g14378(.A1(new_n14693_), .A2(new_n14675_), .ZN(new_n14696_));
  AOI21_X1   g14379(.A1(new_n14695_), .A2(new_n14696_), .B(new_n14674_), .ZN(new_n14697_));
  XOR2_X1    g14380(.A1(new_n14693_), .A2(new_n14675_), .Z(new_n14698_));
  AOI21_X1   g14381(.A1(new_n14698_), .A2(new_n14674_), .B(new_n14697_), .ZN(new_n14699_));
  XNOR2_X1   g14382(.A1(new_n14699_), .A2(new_n14672_), .ZN(new_n14700_));
  NOR2_X1    g14383(.A1(new_n14700_), .A2(new_n14670_), .ZN(new_n14701_));
  XOR2_X1    g14384(.A1(new_n14699_), .A2(new_n14672_), .Z(new_n14702_));
  INV_X1     g14385(.I(new_n14702_), .ZN(new_n14703_));
  AOI21_X1   g14386(.A1(new_n14670_), .A2(new_n14703_), .B(new_n14701_), .ZN(new_n14704_));
  XNOR2_X1   g14387(.A1(new_n14704_), .A2(new_n14585_), .ZN(new_n14705_));
  NAND2_X1   g14388(.A1(new_n14583_), .A2(new_n14705_), .ZN(new_n14706_));
  INV_X1     g14389(.I(new_n14585_), .ZN(new_n14707_));
  NOR2_X1    g14390(.A1(new_n14707_), .A2(new_n14704_), .ZN(new_n14708_));
  NAND2_X1   g14391(.A1(new_n14707_), .A2(new_n14704_), .ZN(new_n14709_));
  INV_X1     g14392(.I(new_n14709_), .ZN(new_n14710_));
  NOR2_X1    g14393(.A1(new_n14710_), .A2(new_n14708_), .ZN(new_n14711_));
  OAI21_X1   g14394(.A1(new_n14583_), .A2(new_n14711_), .B(new_n14706_), .ZN(\asquared[92] ));
  NAND2_X1   g14395(.A1(new_n14578_), .A2(new_n14708_), .ZN(new_n14713_));
  NAND3_X1   g14396(.A1(new_n14420_), .A2(new_n14417_), .A3(new_n14713_), .ZN(new_n14714_));
  AND3_X2    g14397(.A1(new_n14714_), .A2(new_n14579_), .A3(new_n14710_), .Z(\asquared[93] ));
  OAI21_X1   g14398(.A1(new_n14674_), .A2(new_n14694_), .B(new_n14696_), .ZN(new_n14716_));
  INV_X1     g14399(.I(new_n14716_), .ZN(new_n14717_));
  AOI21_X1   g14400(.A1(new_n14687_), .A2(new_n14691_), .B(new_n14689_), .ZN(new_n14718_));
  INV_X1     g14401(.I(new_n6027_), .ZN(new_n14719_));
  OAI22_X1   g14402(.A1(new_n7187_), .A2(new_n12355_), .B1(new_n5322_), .B2(new_n14719_), .ZN(new_n14720_));
  NAND2_X1   g14403(.A1(new_n5742_), .A2(new_n6030_), .ZN(new_n14721_));
  NAND2_X1   g14404(.A1(new_n14720_), .A2(new_n14721_), .ZN(new_n14722_));
  INV_X1     g14405(.I(new_n14722_), .ZN(new_n14723_));
  AOI21_X1   g14406(.A1(new_n14723_), .A2(new_n5512_), .B(\a[48] ), .ZN(new_n14724_));
  NOR2_X1    g14407(.A1(\a[43] ), .A2(\a[49] ), .ZN(new_n14725_));
  OAI21_X1   g14408(.A1(new_n14724_), .A2(new_n4770_), .B(new_n14725_), .ZN(new_n14726_));
  AOI21_X1   g14409(.A1(new_n5742_), .A2(new_n6030_), .B(new_n14720_), .ZN(new_n14727_));
  NAND2_X1   g14410(.A1(new_n14726_), .A2(new_n14727_), .ZN(new_n14728_));
  NAND4_X1   g14411(.A1(\a[34] ), .A2(\a[35] ), .A3(\a[57] ), .A4(\a[58] ), .ZN(new_n14730_));
  NOR2_X1    g14412(.A1(new_n3393_), .A2(new_n7216_), .ZN(new_n14731_));
  INV_X1     g14413(.I(new_n14731_), .ZN(new_n14732_));
  NOR3_X1    g14414(.A1(new_n14732_), .A2(new_n2499_), .A3(new_n9310_), .ZN(new_n14733_));
  XOR2_X1    g14415(.A1(new_n14733_), .A2(new_n2868_), .Z(new_n14734_));
  XOR2_X1    g14416(.A1(new_n14734_), .A2(\a[59] ), .Z(new_n14735_));
  NOR2_X1    g14417(.A1(new_n14735_), .A2(new_n14730_), .ZN(new_n14736_));
  INV_X1     g14418(.I(new_n14736_), .ZN(new_n14737_));
  NAND2_X1   g14419(.A1(new_n14735_), .A2(new_n14730_), .ZN(new_n14738_));
  AOI21_X1   g14420(.A1(new_n14737_), .A2(new_n14738_), .B(new_n14728_), .ZN(new_n14739_));
  INV_X1     g14421(.I(new_n14728_), .ZN(new_n14740_));
  XNOR2_X1   g14422(.A1(new_n14735_), .A2(new_n14730_), .ZN(new_n14741_));
  NOR2_X1    g14423(.A1(new_n14741_), .A2(new_n14740_), .ZN(new_n14742_));
  NOR2_X1    g14424(.A1(new_n14742_), .A2(new_n14739_), .ZN(new_n14743_));
  NOR2_X1    g14425(.A1(new_n2461_), .A2(new_n8453_), .ZN(new_n14744_));
  NAND2_X1   g14426(.A1(\a[31] ), .A2(\a[62] ), .ZN(new_n14745_));
  XOR2_X1    g14427(.A1(new_n14744_), .A2(new_n14745_), .Z(new_n14746_));
  INV_X1     g14428(.I(new_n14746_), .ZN(new_n14747_));
  AOI22_X1   g14429(.A1(new_n4415_), .A2(new_n7204_), .B1(new_n7000_), .B2(new_n6024_), .ZN(new_n14748_));
  NOR2_X1    g14430(.A1(new_n3783_), .A2(new_n6694_), .ZN(new_n14749_));
  NAND4_X1   g14431(.A1(new_n14748_), .A2(new_n6579_), .A3(new_n10034_), .A4(new_n14749_), .ZN(new_n14750_));
  INV_X1     g14432(.I(new_n14750_), .ZN(new_n14751_));
  OAI21_X1   g14433(.A1(new_n14678_), .A2(new_n14431_), .B(new_n14744_), .ZN(new_n14752_));
  OAI21_X1   g14434(.A1(new_n14430_), .A2(new_n14679_), .B(new_n14752_), .ZN(new_n14753_));
  AOI21_X1   g14435(.A1(new_n8424_), .A2(new_n9029_), .B(new_n2499_), .ZN(new_n14754_));
  XNOR2_X1   g14436(.A1(new_n14753_), .A2(new_n14754_), .ZN(new_n14755_));
  XOR2_X1    g14437(.A1(new_n14755_), .A2(new_n14751_), .Z(new_n14756_));
  XOR2_X1    g14438(.A1(new_n14756_), .A2(new_n14747_), .Z(new_n14757_));
  XOR2_X1    g14439(.A1(new_n14757_), .A2(new_n14743_), .Z(new_n14758_));
  NOR2_X1    g14440(.A1(new_n14758_), .A2(new_n14718_), .ZN(new_n14759_));
  INV_X1     g14441(.I(new_n14718_), .ZN(new_n14760_));
  INV_X1     g14442(.I(new_n14743_), .ZN(new_n14761_));
  NOR2_X1    g14443(.A1(new_n14757_), .A2(new_n14761_), .ZN(new_n14762_));
  INV_X1     g14444(.I(new_n14762_), .ZN(new_n14763_));
  NAND2_X1   g14445(.A1(new_n14757_), .A2(new_n14761_), .ZN(new_n14764_));
  AOI21_X1   g14446(.A1(new_n14763_), .A2(new_n14764_), .B(new_n14760_), .ZN(new_n14765_));
  NOR2_X1    g14447(.A1(new_n14759_), .A2(new_n14765_), .ZN(new_n14766_));
  AOI21_X1   g14448(.A1(new_n14640_), .A2(new_n14660_), .B(new_n14658_), .ZN(new_n14767_));
  XOR2_X1    g14449(.A1(new_n14766_), .A2(new_n14767_), .Z(new_n14768_));
  NOR2_X1    g14450(.A1(new_n14768_), .A2(new_n14717_), .ZN(new_n14769_));
  INV_X1     g14451(.I(new_n14766_), .ZN(new_n14770_));
  NOR2_X1    g14452(.A1(new_n14770_), .A2(new_n14767_), .ZN(new_n14771_));
  INV_X1     g14453(.I(new_n14771_), .ZN(new_n14772_));
  NAND2_X1   g14454(.A1(new_n14770_), .A2(new_n14767_), .ZN(new_n14773_));
  AOI21_X1   g14455(.A1(new_n14772_), .A2(new_n14773_), .B(new_n14716_), .ZN(new_n14774_));
  AOI21_X1   g14456(.A1(new_n14620_), .A2(new_n14624_), .B(new_n14622_), .ZN(new_n14775_));
  AOI21_X1   g14457(.A1(new_n14635_), .A2(new_n14638_), .B(new_n14636_), .ZN(new_n14776_));
  NAND2_X1   g14458(.A1(new_n5592_), .A2(new_n6779_), .ZN(new_n14777_));
  NOR2_X1    g14459(.A1(new_n5592_), .A2(new_n6779_), .ZN(new_n14778_));
  NOR2_X1    g14460(.A1(\a[28] ), .A2(\a[63] ), .ZN(new_n14779_));
  AOI21_X1   g14461(.A1(new_n14777_), .A2(new_n14779_), .B(new_n14778_), .ZN(new_n14780_));
  AOI21_X1   g14462(.A1(new_n3851_), .A2(new_n8676_), .B(new_n14646_), .ZN(new_n14781_));
  AOI21_X1   g14463(.A1(new_n5339_), .A2(new_n7204_), .B(new_n14649_), .ZN(new_n14782_));
  XOR2_X1    g14464(.A1(new_n14781_), .A2(new_n14782_), .Z(new_n14783_));
  NAND2_X1   g14465(.A1(new_n14783_), .A2(new_n14780_), .ZN(new_n14784_));
  INV_X1     g14466(.I(new_n14780_), .ZN(new_n14785_));
  AND2_X2    g14467(.A1(new_n14781_), .A2(new_n14782_), .Z(new_n14786_));
  NOR2_X1    g14468(.A1(new_n14781_), .A2(new_n14782_), .ZN(new_n14787_));
  OAI21_X1   g14469(.A1(new_n14786_), .A2(new_n14787_), .B(new_n14785_), .ZN(new_n14788_));
  NAND2_X1   g14470(.A1(new_n14784_), .A2(new_n14788_), .ZN(new_n14789_));
  NAND2_X1   g14471(.A1(new_n5321_), .A2(new_n6030_), .ZN(new_n14790_));
  NOR2_X1    g14472(.A1(new_n5321_), .A2(new_n6030_), .ZN(new_n14791_));
  NOR2_X1    g14473(.A1(\a[35] ), .A2(\a[56] ), .ZN(new_n14792_));
  AOI21_X1   g14474(.A1(new_n14790_), .A2(new_n14792_), .B(new_n14791_), .ZN(new_n14793_));
  INV_X1     g14475(.I(new_n14793_), .ZN(new_n14794_));
  NAND2_X1   g14476(.A1(\a[32] ), .A2(\a[60] ), .ZN(new_n14795_));
  AOI21_X1   g14477(.A1(new_n7483_), .A2(new_n5600_), .B(new_n14795_), .ZN(new_n14796_));
  NAND3_X1   g14478(.A1(new_n7483_), .A2(new_n5600_), .A3(new_n14795_), .ZN(new_n14797_));
  INV_X1     g14479(.I(new_n14797_), .ZN(new_n14798_));
  NOR2_X1    g14480(.A1(new_n14798_), .A2(new_n14796_), .ZN(new_n14799_));
  AOI21_X1   g14481(.A1(new_n4727_), .A2(new_n7639_), .B(new_n10958_), .ZN(new_n14800_));
  NOR2_X1    g14482(.A1(new_n14799_), .A2(new_n14800_), .ZN(new_n14801_));
  INV_X1     g14483(.I(new_n14800_), .ZN(new_n14802_));
  NOR3_X1    g14484(.A1(new_n14802_), .A2(new_n14798_), .A3(new_n14796_), .ZN(new_n14803_));
  NOR2_X1    g14485(.A1(new_n14801_), .A2(new_n14803_), .ZN(new_n14804_));
  NOR2_X1    g14486(.A1(new_n14804_), .A2(new_n14794_), .ZN(new_n14805_));
  XOR2_X1    g14487(.A1(new_n14799_), .A2(new_n14802_), .Z(new_n14806_));
  NOR2_X1    g14488(.A1(new_n14806_), .A2(new_n14793_), .ZN(new_n14807_));
  NOR2_X1    g14489(.A1(new_n14807_), .A2(new_n14805_), .ZN(new_n14808_));
  XNOR2_X1   g14490(.A1(new_n14789_), .A2(new_n14808_), .ZN(new_n14809_));
  NOR2_X1    g14491(.A1(new_n14809_), .A2(new_n14776_), .ZN(new_n14810_));
  INV_X1     g14492(.I(new_n14776_), .ZN(new_n14811_));
  NOR2_X1    g14493(.A1(new_n14789_), .A2(new_n14808_), .ZN(new_n14812_));
  INV_X1     g14494(.I(new_n14812_), .ZN(new_n14813_));
  NAND2_X1   g14495(.A1(new_n14789_), .A2(new_n14808_), .ZN(new_n14814_));
  AOI21_X1   g14496(.A1(new_n14813_), .A2(new_n14814_), .B(new_n14811_), .ZN(new_n14815_));
  NOR2_X1    g14497(.A1(new_n14810_), .A2(new_n14815_), .ZN(new_n14816_));
  INV_X1     g14498(.I(new_n14653_), .ZN(new_n14817_));
  AOI21_X1   g14499(.A1(new_n14817_), .A2(new_n14644_), .B(new_n14652_), .ZN(new_n14818_));
  INV_X1     g14500(.I(new_n14598_), .ZN(new_n14819_));
  AOI21_X1   g14501(.A1(new_n14594_), .A2(new_n14819_), .B(new_n14597_), .ZN(new_n14820_));
  NOR2_X1    g14502(.A1(new_n14611_), .A2(new_n14604_), .ZN(new_n14821_));
  NOR2_X1    g14503(.A1(new_n14821_), .A2(new_n14610_), .ZN(new_n14822_));
  XNOR2_X1   g14504(.A1(new_n14820_), .A2(new_n14822_), .ZN(new_n14823_));
  NOR2_X1    g14505(.A1(new_n14823_), .A2(new_n14818_), .ZN(new_n14824_));
  INV_X1     g14506(.I(new_n14818_), .ZN(new_n14825_));
  NOR2_X1    g14507(.A1(new_n14820_), .A2(new_n14822_), .ZN(new_n14826_));
  INV_X1     g14508(.I(new_n14826_), .ZN(new_n14827_));
  NAND2_X1   g14509(.A1(new_n14820_), .A2(new_n14822_), .ZN(new_n14828_));
  AOI21_X1   g14510(.A1(new_n14827_), .A2(new_n14828_), .B(new_n14825_), .ZN(new_n14829_));
  NOR2_X1    g14511(.A1(new_n14824_), .A2(new_n14829_), .ZN(new_n14830_));
  XNOR2_X1   g14512(.A1(new_n14816_), .A2(new_n14830_), .ZN(new_n14831_));
  NOR2_X1    g14513(.A1(new_n14831_), .A2(new_n14775_), .ZN(new_n14832_));
  INV_X1     g14514(.I(new_n14775_), .ZN(new_n14833_));
  NOR2_X1    g14515(.A1(new_n14816_), .A2(new_n14830_), .ZN(new_n14834_));
  INV_X1     g14516(.I(new_n14834_), .ZN(new_n14835_));
  NAND2_X1   g14517(.A1(new_n14816_), .A2(new_n14830_), .ZN(new_n14836_));
  AOI21_X1   g14518(.A1(new_n14835_), .A2(new_n14836_), .B(new_n14833_), .ZN(new_n14837_));
  NOR4_X1    g14519(.A1(new_n14774_), .A2(new_n14769_), .A3(new_n14832_), .A4(new_n14837_), .ZN(new_n14838_));
  INV_X1     g14520(.I(new_n14666_), .ZN(new_n14839_));
  OAI21_X1   g14521(.A1(new_n14587_), .A2(new_n14665_), .B(new_n14839_), .ZN(new_n14840_));
  NOR2_X1    g14522(.A1(new_n14774_), .A2(new_n14769_), .ZN(new_n14841_));
  NOR2_X1    g14523(.A1(new_n14832_), .A2(new_n14837_), .ZN(new_n14842_));
  NOR2_X1    g14524(.A1(new_n14841_), .A2(new_n14842_), .ZN(new_n14843_));
  INV_X1     g14525(.I(new_n14843_), .ZN(new_n14844_));
  AOI21_X1   g14526(.A1(new_n14844_), .A2(new_n14840_), .B(new_n14838_), .ZN(new_n14845_));
  AOI21_X1   g14527(.A1(new_n14716_), .A2(new_n14773_), .B(new_n14771_), .ZN(new_n14846_));
  OAI21_X1   g14528(.A1(new_n14718_), .A2(new_n14762_), .B(new_n14764_), .ZN(new_n14847_));
  INV_X1     g14529(.I(new_n14847_), .ZN(new_n14848_));
  OAI21_X1   g14530(.A1(new_n14775_), .A2(new_n14834_), .B(new_n14836_), .ZN(new_n14849_));
  NAND2_X1   g14531(.A1(new_n6743_), .A2(new_n9507_), .ZN(new_n14850_));
  INV_X1     g14532(.I(new_n14850_), .ZN(new_n14851_));
  NOR4_X1    g14533(.A1(new_n3837_), .A2(new_n5004_), .A3(new_n5750_), .A4(new_n7216_), .ZN(new_n14852_));
  NAND2_X1   g14534(.A1(new_n14851_), .A2(new_n14852_), .ZN(new_n14853_));
  AOI21_X1   g14535(.A1(new_n14853_), .A2(new_n8953_), .B(new_n4706_), .ZN(new_n14854_));
  NOR3_X1    g14536(.A1(new_n14854_), .A2(new_n3837_), .A3(new_n7216_), .ZN(new_n14855_));
  NOR2_X1    g14537(.A1(new_n14854_), .A2(new_n14851_), .ZN(new_n14856_));
  NOR2_X1    g14538(.A1(new_n5750_), .A2(new_n6999_), .ZN(new_n14857_));
  AOI21_X1   g14539(.A1(\a[38] ), .A2(\a[45] ), .B(new_n14857_), .ZN(new_n14858_));
  AOI21_X1   g14540(.A1(new_n14856_), .A2(new_n14858_), .B(new_n14855_), .ZN(new_n14859_));
  INV_X1     g14541(.I(new_n14859_), .ZN(new_n14860_));
  AOI21_X1   g14542(.A1(new_n4771_), .A2(new_n5173_), .B(new_n12545_), .ZN(new_n14861_));
  NOR4_X1    g14543(.A1(new_n5321_), .A2(new_n6280_), .A3(new_n4769_), .A4(new_n6260_), .ZN(new_n14862_));
  NAND2_X1   g14544(.A1(new_n14861_), .A2(new_n14862_), .ZN(new_n14863_));
  NAND2_X1   g14545(.A1(\a[31] ), .A2(\a[47] ), .ZN(new_n14864_));
  NAND2_X1   g14546(.A1(\a[46] ), .A2(\a[62] ), .ZN(new_n14865_));
  XNOR2_X1   g14547(.A1(new_n14864_), .A2(new_n14865_), .ZN(new_n14866_));
  NOR2_X1    g14548(.A1(new_n14863_), .A2(new_n14866_), .ZN(new_n14867_));
  INV_X1     g14549(.I(new_n14866_), .ZN(new_n14868_));
  AOI21_X1   g14550(.A1(new_n14861_), .A2(new_n14862_), .B(new_n14868_), .ZN(new_n14869_));
  NOR2_X1    g14551(.A1(new_n14867_), .A2(new_n14869_), .ZN(new_n14870_));
  NOR2_X1    g14552(.A1(new_n14860_), .A2(new_n14870_), .ZN(new_n14871_));
  XOR2_X1    g14553(.A1(new_n14863_), .A2(new_n14868_), .Z(new_n14872_));
  INV_X1     g14554(.I(new_n14872_), .ZN(new_n14873_));
  AOI21_X1   g14555(.A1(new_n14860_), .A2(new_n14873_), .B(new_n14871_), .ZN(new_n14874_));
  NAND2_X1   g14556(.A1(new_n14828_), .A2(new_n14825_), .ZN(new_n14875_));
  NAND2_X1   g14557(.A1(new_n14875_), .A2(new_n14827_), .ZN(new_n14876_));
  NOR3_X1    g14558(.A1(new_n12965_), .A2(new_n3393_), .A3(new_n3783_), .ZN(new_n14877_));
  NAND4_X1   g14559(.A1(new_n14877_), .A2(\a[39] ), .A3(\a[54] ), .A4(new_n14047_), .ZN(new_n14878_));
  AOI21_X1   g14560(.A1(new_n14878_), .A2(new_n8246_), .B(new_n3967_), .ZN(new_n14879_));
  NOR3_X1    g14561(.A1(new_n12965_), .A2(new_n3393_), .A3(new_n3783_), .ZN(new_n14880_));
  AOI22_X1   g14562(.A1(new_n2766_), .A2(new_n11018_), .B1(new_n8973_), .B2(new_n9781_), .ZN(new_n14881_));
  NOR4_X1    g14563(.A1(new_n3851_), .A2(new_n8991_), .A3(new_n2461_), .A4(new_n9310_), .ZN(new_n14882_));
  NAND2_X1   g14564(.A1(new_n14881_), .A2(new_n14882_), .ZN(new_n14883_));
  XNOR2_X1   g14565(.A1(new_n5592_), .A2(new_n7204_), .ZN(new_n14884_));
  NOR2_X1    g14566(.A1(new_n14883_), .A2(new_n14884_), .ZN(new_n14885_));
  AND2_X2    g14567(.A1(new_n14883_), .A2(new_n14884_), .Z(new_n14886_));
  OAI21_X1   g14568(.A1(new_n14886_), .A2(new_n14885_), .B(new_n14880_), .ZN(new_n14887_));
  INV_X1     g14569(.I(new_n14880_), .ZN(new_n14888_));
  XOR2_X1    g14570(.A1(new_n14883_), .A2(new_n14884_), .Z(new_n14889_));
  NAND2_X1   g14571(.A1(new_n14889_), .A2(new_n14888_), .ZN(new_n14890_));
  NAND2_X1   g14572(.A1(new_n14890_), .A2(new_n14887_), .ZN(new_n14891_));
  INV_X1     g14573(.I(new_n14891_), .ZN(new_n14892_));
  XOR2_X1    g14574(.A1(new_n14876_), .A2(new_n14892_), .Z(new_n14893_));
  NOR2_X1    g14575(.A1(new_n14893_), .A2(new_n14874_), .ZN(new_n14894_));
  AOI21_X1   g14576(.A1(new_n14875_), .A2(new_n14827_), .B(new_n14892_), .ZN(new_n14895_));
  NOR2_X1    g14577(.A1(new_n14876_), .A2(new_n14891_), .ZN(new_n14896_));
  NOR2_X1    g14578(.A1(new_n14896_), .A2(new_n14895_), .ZN(new_n14897_));
  INV_X1     g14579(.I(new_n14897_), .ZN(new_n14898_));
  AOI21_X1   g14580(.A1(new_n14874_), .A2(new_n14898_), .B(new_n14894_), .ZN(new_n14899_));
  XNOR2_X1   g14581(.A1(new_n14849_), .A2(new_n14899_), .ZN(new_n14900_));
  NOR2_X1    g14582(.A1(new_n14849_), .A2(new_n14899_), .ZN(new_n14901_));
  NAND2_X1   g14583(.A1(new_n14849_), .A2(new_n14899_), .ZN(new_n14902_));
  INV_X1     g14584(.I(new_n14902_), .ZN(new_n14903_));
  OAI21_X1   g14585(.A1(new_n14903_), .A2(new_n14901_), .B(new_n14848_), .ZN(new_n14904_));
  OAI21_X1   g14586(.A1(new_n14848_), .A2(new_n14900_), .B(new_n14904_), .ZN(new_n14905_));
  NAND2_X1   g14587(.A1(new_n14740_), .A2(new_n14738_), .ZN(new_n14906_));
  NAND2_X1   g14588(.A1(new_n14906_), .A2(new_n14737_), .ZN(new_n14907_));
  INV_X1     g14589(.I(new_n14907_), .ZN(new_n14908_));
  NOR2_X1    g14590(.A1(new_n14803_), .A2(new_n14794_), .ZN(new_n14909_));
  NOR2_X1    g14591(.A1(new_n14909_), .A2(new_n14801_), .ZN(new_n14910_));
  NOR2_X1    g14592(.A1(new_n14787_), .A2(new_n14785_), .ZN(new_n14911_));
  NOR2_X1    g14593(.A1(new_n14911_), .A2(new_n14786_), .ZN(new_n14912_));
  XNOR2_X1   g14594(.A1(new_n14912_), .A2(new_n14910_), .ZN(new_n14913_));
  NOR2_X1    g14595(.A1(new_n14908_), .A2(new_n14913_), .ZN(new_n14914_));
  NOR2_X1    g14596(.A1(new_n14912_), .A2(new_n14910_), .ZN(new_n14915_));
  NAND2_X1   g14597(.A1(new_n14912_), .A2(new_n14910_), .ZN(new_n14916_));
  INV_X1     g14598(.I(new_n14916_), .ZN(new_n14917_));
  NOR2_X1    g14599(.A1(new_n14917_), .A2(new_n14915_), .ZN(new_n14918_));
  NOR2_X1    g14600(.A1(new_n14907_), .A2(new_n14918_), .ZN(new_n14919_));
  NOR2_X1    g14601(.A1(new_n14914_), .A2(new_n14919_), .ZN(new_n14920_));
  AOI21_X1   g14602(.A1(new_n14811_), .A2(new_n14814_), .B(new_n14812_), .ZN(new_n14921_));
  INV_X1     g14603(.I(new_n14921_), .ZN(new_n14922_));
  AND2_X2    g14604(.A1(new_n14753_), .A2(new_n14751_), .Z(new_n14923_));
  NOR2_X1    g14605(.A1(new_n14753_), .A2(new_n14751_), .ZN(new_n14924_));
  XOR2_X1    g14606(.A1(new_n14746_), .A2(new_n14754_), .Z(new_n14925_));
  NOR2_X1    g14607(.A1(new_n14924_), .A2(new_n14925_), .ZN(new_n14926_));
  NOR2_X1    g14608(.A1(new_n14926_), .A2(new_n14923_), .ZN(new_n14927_));
  AOI21_X1   g14609(.A1(new_n5592_), .A2(new_n6777_), .B(new_n14748_), .ZN(new_n14928_));
  INV_X1     g14610(.I(new_n14928_), .ZN(new_n14929_));
  NOR4_X1    g14611(.A1(new_n3371_), .A2(new_n3423_), .A3(new_n7727_), .A4(new_n7647_), .ZN(new_n14930_));
  XOR2_X1    g14612(.A1(new_n14722_), .A2(new_n14930_), .Z(new_n14931_));
  NOR2_X1    g14613(.A1(new_n14931_), .A2(new_n14929_), .ZN(new_n14932_));
  INV_X1     g14614(.I(new_n14930_), .ZN(new_n14933_));
  NOR2_X1    g14615(.A1(new_n14722_), .A2(new_n14933_), .ZN(new_n14934_));
  NOR2_X1    g14616(.A1(new_n14723_), .A2(new_n14930_), .ZN(new_n14935_));
  NOR2_X1    g14617(.A1(new_n14935_), .A2(new_n14934_), .ZN(new_n14936_));
  NOR2_X1    g14618(.A1(new_n14936_), .A2(new_n14928_), .ZN(new_n14937_));
  NOR2_X1    g14619(.A1(new_n14937_), .A2(new_n14932_), .ZN(new_n14938_));
  NAND2_X1   g14620(.A1(new_n7483_), .A2(new_n5600_), .ZN(new_n14939_));
  NOR2_X1    g14621(.A1(new_n7483_), .A2(new_n5600_), .ZN(new_n14940_));
  NOR2_X1    g14622(.A1(\a[32] ), .A2(\a[60] ), .ZN(new_n14941_));
  AOI21_X1   g14623(.A1(new_n14939_), .A2(new_n14941_), .B(new_n14940_), .ZN(new_n14942_));
  NOR2_X1    g14624(.A1(new_n13077_), .A2(new_n14731_), .ZN(new_n14943_));
  NOR3_X1    g14625(.A1(new_n14943_), .A2(new_n2868_), .A3(new_n8085_), .ZN(new_n14944_));
  NOR2_X1    g14626(.A1(new_n14944_), .A2(new_n14733_), .ZN(new_n14945_));
  AOI22_X1   g14627(.A1(new_n14747_), .A2(new_n3126_), .B1(new_n9784_), .B2(new_n14754_), .ZN(new_n14946_));
  XNOR2_X1   g14628(.A1(new_n14946_), .A2(new_n14945_), .ZN(new_n14947_));
  INV_X1     g14629(.I(new_n14947_), .ZN(new_n14948_));
  NOR2_X1    g14630(.A1(new_n14946_), .A2(new_n14945_), .ZN(new_n14949_));
  INV_X1     g14631(.I(new_n14949_), .ZN(new_n14950_));
  NAND2_X1   g14632(.A1(new_n14946_), .A2(new_n14945_), .ZN(new_n14951_));
  AOI21_X1   g14633(.A1(new_n14950_), .A2(new_n14951_), .B(new_n14942_), .ZN(new_n14952_));
  AOI21_X1   g14634(.A1(new_n14948_), .A2(new_n14942_), .B(new_n14952_), .ZN(new_n14953_));
  XNOR2_X1   g14635(.A1(new_n14953_), .A2(new_n14938_), .ZN(new_n14954_));
  NOR2_X1    g14636(.A1(new_n14954_), .A2(new_n14927_), .ZN(new_n14955_));
  INV_X1     g14637(.I(new_n14927_), .ZN(new_n14956_));
  NOR2_X1    g14638(.A1(new_n14953_), .A2(new_n14938_), .ZN(new_n14957_));
  INV_X1     g14639(.I(new_n14957_), .ZN(new_n14958_));
  NAND2_X1   g14640(.A1(new_n14953_), .A2(new_n14938_), .ZN(new_n14959_));
  AOI21_X1   g14641(.A1(new_n14959_), .A2(new_n14958_), .B(new_n14956_), .ZN(new_n14960_));
  NOR2_X1    g14642(.A1(new_n14955_), .A2(new_n14960_), .ZN(new_n14961_));
  NOR2_X1    g14643(.A1(new_n14961_), .A2(new_n14922_), .ZN(new_n14962_));
  NOR3_X1    g14644(.A1(new_n14955_), .A2(new_n14960_), .A3(new_n14921_), .ZN(new_n14963_));
  NOR2_X1    g14645(.A1(new_n14962_), .A2(new_n14963_), .ZN(new_n14964_));
  XOR2_X1    g14646(.A1(new_n14961_), .A2(new_n14922_), .Z(new_n14965_));
  NAND2_X1   g14647(.A1(new_n14965_), .A2(new_n14920_), .ZN(new_n14966_));
  OAI21_X1   g14648(.A1(new_n14920_), .A2(new_n14964_), .B(new_n14966_), .ZN(new_n14967_));
  XNOR2_X1   g14649(.A1(new_n14905_), .A2(new_n14967_), .ZN(new_n14968_));
  NOR2_X1    g14650(.A1(new_n14968_), .A2(new_n14846_), .ZN(new_n14969_));
  INV_X1     g14651(.I(new_n14846_), .ZN(new_n14970_));
  NAND2_X1   g14652(.A1(new_n14905_), .A2(new_n14967_), .ZN(new_n14971_));
  NOR2_X1    g14653(.A1(new_n14905_), .A2(new_n14967_), .ZN(new_n14972_));
  INV_X1     g14654(.I(new_n14972_), .ZN(new_n14973_));
  AOI21_X1   g14655(.A1(new_n14973_), .A2(new_n14971_), .B(new_n14970_), .ZN(new_n14974_));
  NOR2_X1    g14656(.A1(new_n14974_), .A2(new_n14969_), .ZN(new_n14975_));
  INV_X1     g14657(.I(new_n14975_), .ZN(new_n14976_));
  XOR2_X1    g14658(.A1(new_n14845_), .A2(new_n14976_), .Z(new_n14977_));
  NAND2_X1   g14659(.A1(\asquared[93] ), .A2(new_n14977_), .ZN(new_n14978_));
  NAND2_X1   g14660(.A1(new_n14845_), .A2(new_n14976_), .ZN(new_n14979_));
  OR2_X2     g14661(.A1(new_n14845_), .A2(new_n14976_), .Z(new_n14980_));
  AND2_X2    g14662(.A1(new_n14980_), .A2(new_n14979_), .Z(new_n14981_));
  OAI21_X1   g14663(.A1(\asquared[93] ), .A2(new_n14981_), .B(new_n14978_), .ZN(\asquared[94] ));
  NAND2_X1   g14664(.A1(\asquared[93] ), .A2(new_n14979_), .ZN(new_n14983_));
  NAND2_X1   g14665(.A1(new_n14983_), .A2(new_n14980_), .ZN(new_n14984_));
  OAI21_X1   g14666(.A1(new_n14848_), .A2(new_n14901_), .B(new_n14902_), .ZN(new_n14985_));
  INV_X1     g14667(.I(new_n14985_), .ZN(new_n14986_));
  INV_X1     g14668(.I(new_n14962_), .ZN(new_n14987_));
  AOI21_X1   g14669(.A1(new_n14987_), .A2(new_n14920_), .B(new_n14963_), .ZN(new_n14988_));
  NOR2_X1    g14670(.A1(new_n14908_), .A2(new_n14917_), .ZN(new_n14989_));
  NOR2_X1    g14671(.A1(new_n14989_), .A2(new_n14915_), .ZN(new_n14990_));
  NOR3_X1    g14672(.A1(new_n14334_), .A2(new_n3783_), .A3(new_n8990_), .ZN(new_n14991_));
  NOR3_X1    g14673(.A1(new_n12540_), .A2(new_n3371_), .A3(new_n3837_), .ZN(new_n14992_));
  NAND2_X1   g14674(.A1(new_n14991_), .A2(new_n14992_), .ZN(new_n14993_));
  AOI21_X1   g14675(.A1(new_n14993_), .A2(new_n10959_), .B(new_n5786_), .ZN(new_n14994_));
  NOR3_X1    g14676(.A1(new_n14994_), .A2(new_n3837_), .A3(new_n7727_), .ZN(new_n14995_));
  NOR2_X1    g14677(.A1(new_n14994_), .A2(new_n14991_), .ZN(new_n14996_));
  AOI21_X1   g14678(.A1(\a[55] ), .A2(\a[60] ), .B(new_n4868_), .ZN(new_n14997_));
  AOI21_X1   g14679(.A1(new_n14996_), .A2(new_n14997_), .B(new_n14995_), .ZN(new_n14998_));
  NOR2_X1    g14680(.A1(new_n4530_), .A2(new_n8989_), .ZN(new_n14999_));
  NAND4_X1   g14681(.A1(new_n14999_), .A2(\a[35] ), .A3(new_n8086_), .A4(\a[62] ), .ZN(new_n15000_));
  AOI21_X1   g14682(.A1(new_n15000_), .A2(new_n9785_), .B(new_n3852_), .ZN(new_n15001_));
  NOR2_X1    g14683(.A1(new_n4530_), .A2(new_n8989_), .ZN(new_n15002_));
  AOI21_X1   g14684(.A1(new_n5321_), .A2(new_n6280_), .B(new_n14861_), .ZN(new_n15003_));
  XOR2_X1    g14685(.A1(new_n15003_), .A2(new_n15002_), .Z(new_n15004_));
  AND2_X2    g14686(.A1(new_n15004_), .A2(new_n14998_), .Z(new_n15005_));
  INV_X1     g14687(.I(new_n15002_), .ZN(new_n15006_));
  INV_X1     g14688(.I(new_n15003_), .ZN(new_n15007_));
  NOR2_X1    g14689(.A1(new_n15007_), .A2(new_n15006_), .ZN(new_n15008_));
  INV_X1     g14690(.I(new_n15008_), .ZN(new_n15009_));
  NAND2_X1   g14691(.A1(new_n15007_), .A2(new_n15006_), .ZN(new_n15010_));
  AOI21_X1   g14692(.A1(new_n15009_), .A2(new_n15010_), .B(new_n14998_), .ZN(new_n15011_));
  NOR2_X1    g14693(.A1(new_n15005_), .A2(new_n15011_), .ZN(new_n15012_));
  NAND2_X1   g14694(.A1(new_n5321_), .A2(new_n6779_), .ZN(new_n15013_));
  NAND2_X1   g14695(.A1(\a[36] ), .A2(\a[58] ), .ZN(new_n15014_));
  XNOR2_X1   g14696(.A1(new_n15013_), .A2(new_n15014_), .ZN(new_n15015_));
  AOI22_X1   g14697(.A1(new_n5592_), .A2(new_n10289_), .B1(new_n12056_), .B2(new_n7482_), .ZN(new_n15016_));
  NOR3_X1    g14698(.A1(new_n8007_), .A2(new_n5350_), .A3(new_n7204_), .ZN(new_n15017_));
  NAND2_X1   g14699(.A1(new_n15017_), .A2(new_n15016_), .ZN(new_n15018_));
  NAND4_X1   g14700(.A1(\a[45] ), .A2(\a[46] ), .A3(\a[48] ), .A4(\a[49] ), .ZN(new_n15019_));
  NOR2_X1    g14701(.A1(new_n15018_), .A2(new_n15019_), .ZN(new_n15020_));
  INV_X1     g14702(.I(new_n15019_), .ZN(new_n15021_));
  AOI21_X1   g14703(.A1(new_n15017_), .A2(new_n15016_), .B(new_n15021_), .ZN(new_n15022_));
  NOR2_X1    g14704(.A1(new_n15020_), .A2(new_n15022_), .ZN(new_n15023_));
  NOR2_X1    g14705(.A1(new_n15023_), .A2(new_n15015_), .ZN(new_n15024_));
  INV_X1     g14706(.I(new_n15015_), .ZN(new_n15025_));
  XOR2_X1    g14707(.A1(new_n15018_), .A2(new_n15021_), .Z(new_n15026_));
  NOR2_X1    g14708(.A1(new_n15026_), .A2(new_n15025_), .ZN(new_n15027_));
  NOR2_X1    g14709(.A1(new_n15027_), .A2(new_n15024_), .ZN(new_n15028_));
  XOR2_X1    g14710(.A1(new_n15012_), .A2(new_n15028_), .Z(new_n15029_));
  NOR2_X1    g14711(.A1(new_n14990_), .A2(new_n15029_), .ZN(new_n15030_));
  OAI21_X1   g14712(.A1(new_n15024_), .A2(new_n15027_), .B(new_n15012_), .ZN(new_n15031_));
  OAI21_X1   g14713(.A1(new_n15005_), .A2(new_n15011_), .B(new_n15028_), .ZN(new_n15032_));
  NAND2_X1   g14714(.A1(new_n15031_), .A2(new_n15032_), .ZN(new_n15033_));
  AOI21_X1   g14715(.A1(new_n14990_), .A2(new_n15033_), .B(new_n15030_), .ZN(new_n15034_));
  NOR2_X1    g14716(.A1(new_n14860_), .A2(new_n14869_), .ZN(new_n15035_));
  INV_X1     g14717(.I(new_n14856_), .ZN(new_n15036_));
  NOR2_X1    g14718(.A1(new_n5511_), .A2(new_n9029_), .ZN(new_n15037_));
  INV_X1     g14719(.I(new_n15037_), .ZN(new_n15038_));
  OAI21_X1   g14720(.A1(new_n15038_), .A2(new_n2655_), .B(new_n5793_), .ZN(new_n15039_));
  NOR2_X1    g14721(.A1(new_n15036_), .A2(new_n15039_), .ZN(new_n15040_));
  XOR2_X1    g14722(.A1(new_n15040_), .A2(new_n2655_), .Z(new_n15041_));
  XOR2_X1    g14723(.A1(new_n15041_), .A2(\a[63] ), .Z(new_n15042_));
  NOR2_X1    g14724(.A1(new_n14879_), .A2(new_n14877_), .ZN(new_n15043_));
  AOI21_X1   g14725(.A1(new_n3851_), .A2(new_n8991_), .B(new_n14881_), .ZN(new_n15044_));
  AOI21_X1   g14726(.A1(new_n5592_), .A2(new_n14037_), .B(new_n7204_), .ZN(new_n15045_));
  XOR2_X1    g14727(.A1(new_n15044_), .A2(new_n15045_), .Z(new_n15046_));
  INV_X1     g14728(.I(new_n15046_), .ZN(new_n15047_));
  INV_X1     g14729(.I(new_n15044_), .ZN(new_n15048_));
  NOR2_X1    g14730(.A1(new_n15048_), .A2(new_n15045_), .ZN(new_n15049_));
  INV_X1     g14731(.I(new_n15049_), .ZN(new_n15050_));
  NAND2_X1   g14732(.A1(new_n15048_), .A2(new_n15045_), .ZN(new_n15051_));
  AOI21_X1   g14733(.A1(new_n15050_), .A2(new_n15051_), .B(new_n15043_), .ZN(new_n15052_));
  AOI21_X1   g14734(.A1(new_n15043_), .A2(new_n15047_), .B(new_n15052_), .ZN(new_n15053_));
  XOR2_X1    g14735(.A1(new_n15042_), .A2(new_n15053_), .Z(new_n15054_));
  OAI21_X1   g14736(.A1(new_n14867_), .A2(new_n15035_), .B(new_n15054_), .ZN(new_n15055_));
  NOR2_X1    g14737(.A1(new_n15035_), .A2(new_n14867_), .ZN(new_n15056_));
  NOR2_X1    g14738(.A1(new_n15042_), .A2(new_n15053_), .ZN(new_n15057_));
  NAND2_X1   g14739(.A1(new_n15042_), .A2(new_n15053_), .ZN(new_n15058_));
  INV_X1     g14740(.I(new_n15058_), .ZN(new_n15059_));
  OAI21_X1   g14741(.A1(new_n15059_), .A2(new_n15057_), .B(new_n15056_), .ZN(new_n15060_));
  NAND2_X1   g14742(.A1(new_n15055_), .A2(new_n15060_), .ZN(new_n15061_));
  INV_X1     g14743(.I(new_n15061_), .ZN(new_n15062_));
  NOR2_X1    g14744(.A1(new_n15062_), .A2(new_n15034_), .ZN(new_n15063_));
  INV_X1     g14745(.I(new_n15063_), .ZN(new_n15064_));
  NAND2_X1   g14746(.A1(new_n15062_), .A2(new_n15034_), .ZN(new_n15065_));
  AOI21_X1   g14747(.A1(new_n15064_), .A2(new_n15065_), .B(new_n14988_), .ZN(new_n15066_));
  XNOR2_X1   g14748(.A1(new_n15061_), .A2(new_n15034_), .ZN(new_n15067_));
  AOI21_X1   g14749(.A1(new_n14988_), .A2(new_n15067_), .B(new_n15066_), .ZN(new_n15068_));
  NOR2_X1    g14750(.A1(new_n14896_), .A2(new_n14874_), .ZN(new_n15069_));
  NOR2_X1    g14751(.A1(new_n15069_), .A2(new_n14895_), .ZN(new_n15070_));
  NOR2_X1    g14752(.A1(new_n14886_), .A2(new_n14888_), .ZN(new_n15071_));
  NOR2_X1    g14753(.A1(new_n15071_), .A2(new_n14885_), .ZN(new_n15072_));
  NAND2_X1   g14754(.A1(new_n14951_), .A2(new_n14942_), .ZN(new_n15073_));
  NAND2_X1   g14755(.A1(new_n15073_), .A2(new_n14950_), .ZN(new_n15074_));
  NOR2_X1    g14756(.A1(new_n14935_), .A2(new_n14929_), .ZN(new_n15075_));
  NOR2_X1    g14757(.A1(new_n15075_), .A2(new_n14934_), .ZN(new_n15076_));
  XOR2_X1    g14758(.A1(new_n15074_), .A2(new_n15076_), .Z(new_n15077_));
  NOR2_X1    g14759(.A1(new_n15077_), .A2(new_n15072_), .ZN(new_n15078_));
  INV_X1     g14760(.I(new_n15072_), .ZN(new_n15079_));
  INV_X1     g14761(.I(new_n15074_), .ZN(new_n15080_));
  NOR2_X1    g14762(.A1(new_n15080_), .A2(new_n15076_), .ZN(new_n15081_));
  INV_X1     g14763(.I(new_n15081_), .ZN(new_n15082_));
  NAND2_X1   g14764(.A1(new_n15080_), .A2(new_n15076_), .ZN(new_n15083_));
  AOI21_X1   g14765(.A1(new_n15082_), .A2(new_n15083_), .B(new_n15079_), .ZN(new_n15084_));
  NOR2_X1    g14766(.A1(new_n15084_), .A2(new_n15078_), .ZN(new_n15085_));
  OAI21_X1   g14767(.A1(new_n14927_), .A2(new_n14957_), .B(new_n14959_), .ZN(new_n15086_));
  XNOR2_X1   g14768(.A1(new_n15085_), .A2(new_n15086_), .ZN(new_n15087_));
  AND2_X2    g14769(.A1(new_n15085_), .A2(new_n15086_), .Z(new_n15088_));
  NOR2_X1    g14770(.A1(new_n15085_), .A2(new_n15086_), .ZN(new_n15089_));
  OAI21_X1   g14771(.A1(new_n15088_), .A2(new_n15089_), .B(new_n15070_), .ZN(new_n15090_));
  OAI21_X1   g14772(.A1(new_n15070_), .A2(new_n15087_), .B(new_n15090_), .ZN(new_n15091_));
  XNOR2_X1   g14773(.A1(new_n15068_), .A2(new_n15091_), .ZN(new_n15092_));
  NOR2_X1    g14774(.A1(new_n15092_), .A2(new_n14986_), .ZN(new_n15093_));
  NAND2_X1   g14775(.A1(new_n15068_), .A2(new_n15091_), .ZN(new_n15094_));
  NOR2_X1    g14776(.A1(new_n15068_), .A2(new_n15091_), .ZN(new_n15095_));
  INV_X1     g14777(.I(new_n15095_), .ZN(new_n15096_));
  AOI21_X1   g14778(.A1(new_n15096_), .A2(new_n15094_), .B(new_n14985_), .ZN(new_n15097_));
  NOR2_X1    g14779(.A1(new_n15093_), .A2(new_n15097_), .ZN(new_n15098_));
  AOI21_X1   g14780(.A1(new_n14970_), .A2(new_n14971_), .B(new_n14972_), .ZN(new_n15099_));
  XNOR2_X1   g14781(.A1(new_n15098_), .A2(new_n15099_), .ZN(new_n15100_));
  NAND2_X1   g14782(.A1(new_n14984_), .A2(new_n15100_), .ZN(new_n15101_));
  INV_X1     g14783(.I(new_n15098_), .ZN(new_n15102_));
  NOR2_X1    g14784(.A1(new_n15102_), .A2(new_n15099_), .ZN(new_n15103_));
  NAND2_X1   g14785(.A1(new_n15102_), .A2(new_n15099_), .ZN(new_n15104_));
  INV_X1     g14786(.I(new_n15104_), .ZN(new_n15105_));
  NOR2_X1    g14787(.A1(new_n15105_), .A2(new_n15103_), .ZN(new_n15106_));
  OAI21_X1   g14788(.A1(new_n14984_), .A2(new_n15106_), .B(new_n15101_), .ZN(\asquared[95] ));
  NOR2_X1    g14789(.A1(new_n15103_), .A2(new_n14976_), .ZN(new_n15108_));
  NAND2_X1   g14790(.A1(new_n15103_), .A2(new_n14976_), .ZN(new_n15109_));
  AOI21_X1   g14791(.A1(new_n14845_), .A2(new_n15109_), .B(new_n15108_), .ZN(new_n15110_));
  NAND4_X1   g14792(.A1(new_n14714_), .A2(new_n14579_), .A3(new_n14710_), .A4(new_n15110_), .ZN(new_n15111_));
  OAI21_X1   g14793(.A1(new_n14988_), .A2(new_n15063_), .B(new_n15065_), .ZN(new_n15112_));
  INV_X1     g14794(.I(new_n15112_), .ZN(new_n15113_));
  OAI21_X1   g14795(.A1(new_n14989_), .A2(new_n14915_), .B(new_n15032_), .ZN(new_n15114_));
  NAND2_X1   g14796(.A1(new_n15114_), .A2(new_n15031_), .ZN(new_n15115_));
  OAI21_X1   g14797(.A1(new_n15056_), .A2(new_n15057_), .B(new_n15058_), .ZN(new_n15116_));
  AOI21_X1   g14798(.A1(new_n15036_), .A2(new_n15039_), .B(new_n12332_), .ZN(new_n15117_));
  NOR2_X1    g14799(.A1(new_n15117_), .A2(new_n15040_), .ZN(new_n15118_));
  NAND2_X1   g14800(.A1(new_n15043_), .A2(new_n15051_), .ZN(new_n15119_));
  NAND2_X1   g14801(.A1(new_n15119_), .A2(new_n15050_), .ZN(new_n15120_));
  NOR4_X1    g14802(.A1(new_n5004_), .A2(new_n5175_), .A3(new_n5750_), .A4(new_n5745_), .ZN(new_n15121_));
  INV_X1     g14803(.I(new_n15121_), .ZN(new_n15122_));
  NAND2_X1   g14804(.A1(\a[35] ), .A2(\a[59] ), .ZN(new_n15123_));
  NOR2_X1    g14805(.A1(new_n3393_), .A2(new_n8990_), .ZN(new_n15124_));
  XOR2_X1    g14806(.A1(new_n15124_), .A2(new_n15123_), .Z(new_n15125_));
  XOR2_X1    g14807(.A1(new_n15125_), .A2(new_n15122_), .Z(new_n15126_));
  XOR2_X1    g14808(.A1(new_n15120_), .A2(new_n15126_), .Z(new_n15127_));
  NOR2_X1    g14809(.A1(new_n15127_), .A2(new_n15118_), .ZN(new_n15128_));
  INV_X1     g14810(.I(new_n15118_), .ZN(new_n15129_));
  INV_X1     g14811(.I(new_n15120_), .ZN(new_n15130_));
  NOR2_X1    g14812(.A1(new_n15130_), .A2(new_n15126_), .ZN(new_n15131_));
  INV_X1     g14813(.I(new_n15131_), .ZN(new_n15132_));
  NAND2_X1   g14814(.A1(new_n15130_), .A2(new_n15126_), .ZN(new_n15133_));
  AOI21_X1   g14815(.A1(new_n15132_), .A2(new_n15133_), .B(new_n15129_), .ZN(new_n15134_));
  NOR2_X1    g14816(.A1(new_n15134_), .A2(new_n15128_), .ZN(new_n15135_));
  XNOR2_X1   g14817(.A1(new_n15116_), .A2(new_n15135_), .ZN(new_n15136_));
  INV_X1     g14818(.I(new_n15136_), .ZN(new_n15137_));
  NOR2_X1    g14819(.A1(new_n15116_), .A2(new_n15135_), .ZN(new_n15138_));
  INV_X1     g14820(.I(new_n15138_), .ZN(new_n15139_));
  NAND2_X1   g14821(.A1(new_n15116_), .A2(new_n15135_), .ZN(new_n15140_));
  AOI21_X1   g14822(.A1(new_n15139_), .A2(new_n15140_), .B(new_n15115_), .ZN(new_n15141_));
  AOI21_X1   g14823(.A1(new_n15137_), .A2(new_n15115_), .B(new_n15141_), .ZN(new_n15142_));
  INV_X1     g14824(.I(new_n15142_), .ZN(new_n15143_));
  NOR2_X1    g14825(.A1(new_n15070_), .A2(new_n15089_), .ZN(new_n15144_));
  NOR2_X1    g14826(.A1(new_n15144_), .A2(new_n15088_), .ZN(new_n15145_));
  NAND2_X1   g14827(.A1(new_n15083_), .A2(new_n15079_), .ZN(new_n15146_));
  NOR2_X1    g14828(.A1(new_n3837_), .A2(new_n4240_), .ZN(new_n15147_));
  NOR2_X1    g14829(.A1(new_n6999_), .A2(new_n7647_), .ZN(new_n15148_));
  NAND4_X1   g14830(.A1(new_n4241_), .A2(new_n10958_), .A3(new_n15147_), .A4(new_n15148_), .ZN(new_n15149_));
  AOI21_X1   g14831(.A1(new_n15149_), .A2(new_n8246_), .B(new_n4706_), .ZN(new_n15150_));
  NOR2_X1    g14832(.A1(new_n8251_), .A2(new_n10959_), .ZN(new_n15152_));
  NOR2_X1    g14833(.A1(new_n5321_), .A2(new_n6779_), .ZN(new_n15153_));
  NAND2_X1   g14834(.A1(new_n3393_), .A2(new_n7647_), .ZN(new_n15154_));
  AOI21_X1   g14835(.A1(new_n5321_), .A2(new_n6779_), .B(new_n15154_), .ZN(new_n15155_));
  NOR2_X1    g14836(.A1(new_n15155_), .A2(new_n15153_), .ZN(new_n15156_));
  INV_X1     g14837(.I(new_n15156_), .ZN(new_n15157_));
  NAND2_X1   g14838(.A1(new_n4368_), .A2(new_n9781_), .ZN(new_n15158_));
  NAND2_X1   g14839(.A1(\a[41] ), .A2(\a[54] ), .ZN(new_n15159_));
  XNOR2_X1   g14840(.A1(new_n15158_), .A2(new_n15159_), .ZN(new_n15160_));
  NOR2_X1    g14841(.A1(new_n15160_), .A2(new_n15157_), .ZN(new_n15161_));
  NAND2_X1   g14842(.A1(new_n15160_), .A2(new_n15157_), .ZN(new_n15162_));
  INV_X1     g14843(.I(new_n15162_), .ZN(new_n15163_));
  OAI21_X1   g14844(.A1(new_n15163_), .A2(new_n15161_), .B(new_n15152_), .ZN(new_n15164_));
  INV_X1     g14845(.I(new_n15152_), .ZN(new_n15165_));
  XOR2_X1    g14846(.A1(new_n15160_), .A2(new_n15157_), .Z(new_n15166_));
  NAND2_X1   g14847(.A1(new_n15166_), .A2(new_n15165_), .ZN(new_n15167_));
  NAND2_X1   g14848(.A1(new_n15167_), .A2(new_n15164_), .ZN(new_n15168_));
  INV_X1     g14849(.I(new_n15168_), .ZN(new_n15169_));
  NAND2_X1   g14850(.A1(new_n5488_), .A2(new_n6280_), .ZN(new_n15170_));
  NAND2_X1   g14851(.A1(\a[39] ), .A2(\a[56] ), .ZN(new_n15171_));
  XNOR2_X1   g14852(.A1(new_n15170_), .A2(new_n15171_), .ZN(new_n15172_));
  INV_X1     g14853(.I(new_n15172_), .ZN(new_n15173_));
  AOI22_X1   g14854(.A1(new_n4771_), .A2(new_n7204_), .B1(new_n5173_), .B2(new_n7000_), .ZN(new_n15174_));
  NAND4_X1   g14855(.A1(new_n15174_), .A2(new_n5322_), .A3(new_n10034_), .A4(new_n8177_), .ZN(new_n15175_));
  NAND2_X1   g14856(.A1(\a[33] ), .A2(\a[48] ), .ZN(new_n15176_));
  XOR2_X1    g14857(.A1(new_n15037_), .A2(new_n15176_), .Z(new_n15177_));
  NOR2_X1    g14858(.A1(new_n15175_), .A2(new_n15177_), .ZN(new_n15178_));
  AND2_X2    g14859(.A1(new_n15175_), .A2(new_n15177_), .Z(new_n15179_));
  OAI21_X1   g14860(.A1(new_n15179_), .A2(new_n15178_), .B(new_n15173_), .ZN(new_n15180_));
  XOR2_X1    g14861(.A1(new_n15175_), .A2(new_n15177_), .Z(new_n15181_));
  NAND2_X1   g14862(.A1(new_n15181_), .A2(new_n15172_), .ZN(new_n15182_));
  NAND2_X1   g14863(.A1(new_n15182_), .A2(new_n15180_), .ZN(new_n15183_));
  INV_X1     g14864(.I(new_n15183_), .ZN(new_n15184_));
  NOR2_X1    g14865(.A1(new_n15169_), .A2(new_n15184_), .ZN(new_n15185_));
  INV_X1     g14866(.I(new_n15185_), .ZN(new_n15186_));
  NOR2_X1    g14867(.A1(new_n15168_), .A2(new_n15183_), .ZN(new_n15187_));
  INV_X1     g14868(.I(new_n15187_), .ZN(new_n15188_));
  AOI22_X1   g14869(.A1(new_n15186_), .A2(new_n15188_), .B1(new_n15082_), .B2(new_n15146_), .ZN(new_n15189_));
  NAND2_X1   g14870(.A1(new_n15146_), .A2(new_n15082_), .ZN(new_n15190_));
  XNOR2_X1   g14871(.A1(new_n15168_), .A2(new_n15183_), .ZN(new_n15191_));
  NOR2_X1    g14872(.A1(new_n15190_), .A2(new_n15191_), .ZN(new_n15192_));
  AOI21_X1   g14873(.A1(new_n14998_), .A2(new_n15010_), .B(new_n15008_), .ZN(new_n15193_));
  NOR2_X1    g14874(.A1(new_n15001_), .A2(new_n14999_), .ZN(new_n15194_));
  INV_X1     g14875(.I(new_n15194_), .ZN(new_n15195_));
  AOI21_X1   g14876(.A1(new_n5350_), .A2(new_n7204_), .B(new_n15016_), .ZN(new_n15196_));
  XNOR2_X1   g14877(.A1(new_n14996_), .A2(new_n15196_), .ZN(new_n15197_));
  INV_X1     g14878(.I(new_n14996_), .ZN(new_n15198_));
  INV_X1     g14879(.I(new_n15196_), .ZN(new_n15199_));
  NOR2_X1    g14880(.A1(new_n15198_), .A2(new_n15199_), .ZN(new_n15200_));
  NOR2_X1    g14881(.A1(new_n14996_), .A2(new_n15196_), .ZN(new_n15201_));
  OAI21_X1   g14882(.A1(new_n15200_), .A2(new_n15201_), .B(new_n15195_), .ZN(new_n15202_));
  OAI21_X1   g14883(.A1(new_n15195_), .A2(new_n15197_), .B(new_n15202_), .ZN(new_n15203_));
  INV_X1     g14884(.I(new_n15022_), .ZN(new_n15204_));
  AOI21_X1   g14885(.A1(new_n15025_), .A2(new_n15204_), .B(new_n15020_), .ZN(new_n15205_));
  XNOR2_X1   g14886(.A1(new_n15203_), .A2(new_n15205_), .ZN(new_n15206_));
  NOR2_X1    g14887(.A1(new_n15206_), .A2(new_n15193_), .ZN(new_n15207_));
  INV_X1     g14888(.I(new_n15193_), .ZN(new_n15208_));
  NOR2_X1    g14889(.A1(new_n15203_), .A2(new_n15205_), .ZN(new_n15209_));
  INV_X1     g14890(.I(new_n15209_), .ZN(new_n15210_));
  NAND2_X1   g14891(.A1(new_n15203_), .A2(new_n15205_), .ZN(new_n15211_));
  AOI21_X1   g14892(.A1(new_n15210_), .A2(new_n15211_), .B(new_n15208_), .ZN(new_n15212_));
  NOR2_X1    g14893(.A1(new_n15207_), .A2(new_n15212_), .ZN(new_n15213_));
  NOR3_X1    g14894(.A1(new_n15189_), .A2(new_n15192_), .A3(new_n15213_), .ZN(new_n15214_));
  NOR2_X1    g14895(.A1(new_n15192_), .A2(new_n15189_), .ZN(new_n15215_));
  INV_X1     g14896(.I(new_n15213_), .ZN(new_n15216_));
  NOR2_X1    g14897(.A1(new_n15216_), .A2(new_n15215_), .ZN(new_n15217_));
  NOR2_X1    g14898(.A1(new_n15217_), .A2(new_n15214_), .ZN(new_n15218_));
  NOR2_X1    g14899(.A1(new_n15218_), .A2(new_n15145_), .ZN(new_n15219_));
  XNOR2_X1   g14900(.A1(new_n15213_), .A2(new_n15215_), .ZN(new_n15220_));
  AOI21_X1   g14901(.A1(new_n15145_), .A2(new_n15220_), .B(new_n15219_), .ZN(new_n15221_));
  NOR2_X1    g14902(.A1(new_n15143_), .A2(new_n15221_), .ZN(new_n15222_));
  INV_X1     g14903(.I(new_n15222_), .ZN(new_n15223_));
  NAND2_X1   g14904(.A1(new_n15143_), .A2(new_n15221_), .ZN(new_n15224_));
  AOI21_X1   g14905(.A1(new_n15223_), .A2(new_n15224_), .B(new_n15113_), .ZN(new_n15225_));
  XOR2_X1    g14906(.A1(new_n15221_), .A2(new_n15142_), .Z(new_n15226_));
  NOR2_X1    g14907(.A1(new_n15226_), .A2(new_n15112_), .ZN(new_n15227_));
  NOR2_X1    g14908(.A1(new_n15225_), .A2(new_n15227_), .ZN(new_n15228_));
  AOI21_X1   g14909(.A1(new_n14985_), .A2(new_n15094_), .B(new_n15095_), .ZN(new_n15229_));
  NOR2_X1    g14910(.A1(new_n15229_), .A2(new_n15228_), .ZN(new_n15230_));
  XOR2_X1    g14911(.A1(new_n15111_), .A2(new_n15230_), .Z(new_n15231_));
  XOR2_X1    g14912(.A1(new_n15231_), .A2(new_n15104_), .Z(\asquared[96] ));
  OAI21_X1   g14913(.A1(new_n15225_), .A2(new_n15227_), .B(new_n15105_), .ZN(new_n15233_));
  AOI21_X1   g14914(.A1(new_n15104_), .A2(new_n15228_), .B(new_n15229_), .ZN(new_n15234_));
  INV_X1     g14915(.I(new_n15234_), .ZN(new_n15235_));
  OAI21_X1   g14916(.A1(new_n15111_), .A2(new_n15235_), .B(new_n15233_), .ZN(new_n15236_));
  INV_X1     g14917(.I(new_n15236_), .ZN(new_n15237_));
  INV_X1     g14918(.I(new_n15140_), .ZN(new_n15238_));
  AOI21_X1   g14919(.A1(new_n15115_), .A2(new_n15139_), .B(new_n15238_), .ZN(new_n15239_));
  INV_X1     g14920(.I(new_n15200_), .ZN(new_n15240_));
  OAI21_X1   g14921(.A1(new_n15195_), .A2(new_n15201_), .B(new_n15240_), .ZN(new_n15241_));
  NOR2_X1    g14922(.A1(new_n5174_), .A2(new_n10288_), .ZN(new_n15242_));
  NAND4_X1   g14923(.A1(new_n15242_), .A2(\a[43] ), .A3(\a[53] ), .A4(new_n8187_), .ZN(new_n15243_));
  AOI21_X1   g14924(.A1(new_n15243_), .A2(new_n8005_), .B(new_n5881_), .ZN(new_n15244_));
  NOR2_X1    g14925(.A1(new_n5174_), .A2(new_n10288_), .ZN(new_n15245_));
  AOI21_X1   g14926(.A1(new_n3424_), .A2(new_n4372_), .B(new_n13620_), .ZN(new_n15246_));
  NOR4_X1    g14927(.A1(new_n3487_), .A2(new_n9784_), .A3(new_n2868_), .A4(new_n9310_), .ZN(new_n15247_));
  NAND2_X1   g14928(.A1(new_n15246_), .A2(new_n15247_), .ZN(new_n15248_));
  XOR2_X1    g14929(.A1(new_n15248_), .A2(new_n15245_), .Z(new_n15249_));
  INV_X1     g14930(.I(new_n15249_), .ZN(new_n15250_));
  INV_X1     g14931(.I(new_n15245_), .ZN(new_n15251_));
  NOR2_X1    g14932(.A1(new_n15248_), .A2(new_n15251_), .ZN(new_n15252_));
  INV_X1     g14933(.I(new_n15252_), .ZN(new_n15253_));
  NAND2_X1   g14934(.A1(new_n15248_), .A2(new_n15251_), .ZN(new_n15254_));
  AOI21_X1   g14935(.A1(new_n15253_), .A2(new_n15254_), .B(new_n15241_), .ZN(new_n15255_));
  AOI21_X1   g14936(.A1(new_n15241_), .A2(new_n15250_), .B(new_n15255_), .ZN(new_n15256_));
  INV_X1     g14937(.I(new_n15256_), .ZN(new_n15257_));
  NAND2_X1   g14938(.A1(new_n15133_), .A2(new_n15129_), .ZN(new_n15258_));
  NAND2_X1   g14939(.A1(new_n15258_), .A2(new_n15132_), .ZN(new_n15259_));
  AOI21_X1   g14940(.A1(new_n4241_), .A2(new_n10958_), .B(new_n15150_), .ZN(new_n15260_));
  OAI22_X1   g14941(.A1(new_n15125_), .A2(new_n9553_), .B1(new_n3967_), .B2(new_n15122_), .ZN(new_n15261_));
  NAND2_X1   g14942(.A1(new_n4368_), .A2(new_n9781_), .ZN(new_n15262_));
  NOR2_X1    g14943(.A1(new_n4368_), .A2(new_n9781_), .ZN(new_n15263_));
  NOR2_X1    g14944(.A1(\a[41] ), .A2(\a[54] ), .ZN(new_n15264_));
  AOI21_X1   g14945(.A1(new_n15262_), .A2(new_n15264_), .B(new_n15263_), .ZN(new_n15265_));
  INV_X1     g14946(.I(new_n15265_), .ZN(new_n15266_));
  XOR2_X1    g14947(.A1(new_n15261_), .A2(new_n15266_), .Z(new_n15267_));
  INV_X1     g14948(.I(new_n15261_), .ZN(new_n15268_));
  NOR2_X1    g14949(.A1(new_n15268_), .A2(new_n15266_), .ZN(new_n15269_));
  NOR2_X1    g14950(.A1(new_n15261_), .A2(new_n15265_), .ZN(new_n15270_));
  NOR2_X1    g14951(.A1(new_n15269_), .A2(new_n15270_), .ZN(new_n15271_));
  MUX2_X1    g14952(.I0(new_n15271_), .I1(new_n15267_), .S(new_n15260_), .Z(new_n15272_));
  NOR2_X1    g14953(.A1(new_n15259_), .A2(new_n15272_), .ZN(new_n15273_));
  NAND2_X1   g14954(.A1(new_n15259_), .A2(new_n15272_), .ZN(new_n15274_));
  INV_X1     g14955(.I(new_n15274_), .ZN(new_n15275_));
  OAI21_X1   g14956(.A1(new_n15275_), .A2(new_n15273_), .B(new_n15257_), .ZN(new_n15276_));
  XNOR2_X1   g14957(.A1(new_n15259_), .A2(new_n15272_), .ZN(new_n15277_));
  OAI21_X1   g14958(.A1(new_n15257_), .A2(new_n15277_), .B(new_n15276_), .ZN(new_n15278_));
  AOI21_X1   g14959(.A1(new_n15152_), .A2(new_n15162_), .B(new_n15161_), .ZN(new_n15279_));
  INV_X1     g14960(.I(new_n15279_), .ZN(new_n15280_));
  NAND2_X1   g14961(.A1(new_n5488_), .A2(new_n6280_), .ZN(new_n15281_));
  NOR2_X1    g14962(.A1(new_n5488_), .A2(new_n6280_), .ZN(new_n15282_));
  NOR2_X1    g14963(.A1(\a[39] ), .A2(\a[56] ), .ZN(new_n15283_));
  AOI21_X1   g14964(.A1(new_n15281_), .A2(new_n15283_), .B(new_n15282_), .ZN(new_n15284_));
  INV_X1     g14965(.I(new_n15284_), .ZN(new_n15285_));
  AOI21_X1   g14966(.A1(new_n5321_), .A2(new_n6777_), .B(new_n15174_), .ZN(new_n15286_));
  AOI21_X1   g14967(.A1(new_n7693_), .A2(new_n9029_), .B(new_n2868_), .ZN(new_n15287_));
  INV_X1     g14968(.I(new_n15287_), .ZN(new_n15288_));
  XOR2_X1    g14969(.A1(new_n15286_), .A2(new_n15288_), .Z(new_n15289_));
  NOR2_X1    g14970(.A1(new_n15289_), .A2(new_n15285_), .ZN(new_n15290_));
  INV_X1     g14971(.I(new_n15286_), .ZN(new_n15291_));
  NOR2_X1    g14972(.A1(new_n15291_), .A2(new_n15288_), .ZN(new_n15292_));
  NOR2_X1    g14973(.A1(new_n15286_), .A2(new_n15287_), .ZN(new_n15293_));
  NOR2_X1    g14974(.A1(new_n15292_), .A2(new_n15293_), .ZN(new_n15294_));
  NOR2_X1    g14975(.A1(new_n15294_), .A2(new_n15284_), .ZN(new_n15295_));
  NOR2_X1    g14976(.A1(new_n15295_), .A2(new_n15290_), .ZN(new_n15296_));
  NOR2_X1    g14977(.A1(new_n15179_), .A2(new_n15172_), .ZN(new_n15297_));
  NOR2_X1    g14978(.A1(new_n15297_), .A2(new_n15178_), .ZN(new_n15298_));
  INV_X1     g14979(.I(new_n15298_), .ZN(new_n15299_));
  XOR2_X1    g14980(.A1(new_n15296_), .A2(new_n15299_), .Z(new_n15300_));
  NAND2_X1   g14981(.A1(new_n15300_), .A2(new_n15280_), .ZN(new_n15301_));
  NOR3_X1    g14982(.A1(new_n15295_), .A2(new_n15298_), .A3(new_n15290_), .ZN(new_n15302_));
  NOR2_X1    g14983(.A1(new_n15296_), .A2(new_n15299_), .ZN(new_n15303_));
  OAI21_X1   g14984(.A1(new_n15303_), .A2(new_n15302_), .B(new_n15279_), .ZN(new_n15304_));
  NAND2_X1   g14985(.A1(new_n15301_), .A2(new_n15304_), .ZN(new_n15305_));
  INV_X1     g14986(.I(new_n15305_), .ZN(new_n15306_));
  XOR2_X1    g14987(.A1(new_n15278_), .A2(new_n15306_), .Z(new_n15307_));
  NOR2_X1    g14988(.A1(new_n15307_), .A2(new_n15239_), .ZN(new_n15308_));
  INV_X1     g14989(.I(new_n15239_), .ZN(new_n15309_));
  AND2_X2    g14990(.A1(new_n15278_), .A2(new_n15305_), .Z(new_n15310_));
  NOR2_X1    g14991(.A1(new_n15278_), .A2(new_n15305_), .ZN(new_n15311_));
  NOR2_X1    g14992(.A1(new_n15310_), .A2(new_n15311_), .ZN(new_n15312_));
  NOR2_X1    g14993(.A1(new_n15309_), .A2(new_n15312_), .ZN(new_n15313_));
  NOR2_X1    g14994(.A1(new_n15313_), .A2(new_n15308_), .ZN(new_n15314_));
  NOR2_X1    g14995(.A1(new_n15145_), .A2(new_n15214_), .ZN(new_n15315_));
  NOR2_X1    g14996(.A1(new_n15315_), .A2(new_n15217_), .ZN(new_n15316_));
  AOI21_X1   g14997(.A1(new_n15190_), .A2(new_n15188_), .B(new_n15185_), .ZN(new_n15317_));
  NOR3_X1    g14998(.A1(new_n8424_), .A2(new_n8941_), .A3(new_n5793_), .ZN(new_n15318_));
  NOR4_X1    g14999(.A1(new_n14719_), .A2(new_n7512_), .A3(new_n5004_), .A4(new_n6260_), .ZN(new_n15319_));
  NOR2_X1    g15000(.A1(new_n15319_), .A2(new_n15318_), .ZN(new_n15320_));
  INV_X1     g15001(.I(new_n15320_), .ZN(new_n15321_));
  AOI21_X1   g15002(.A1(new_n5980_), .A2(new_n6280_), .B(new_n15321_), .ZN(new_n15322_));
  AND2_X2    g15003(.A1(new_n15322_), .A2(new_n6027_), .Z(new_n15323_));
  OAI21_X1   g15004(.A1(new_n15323_), .A2(\a[50] ), .B(\a[46] ), .ZN(new_n15324_));
  NOR2_X1    g15005(.A1(\a[45] ), .A2(\a[51] ), .ZN(new_n15325_));
  AOI21_X1   g15006(.A1(new_n15324_), .A2(new_n15325_), .B(new_n15320_), .ZN(new_n15326_));
  NOR3_X1    g15007(.A1(new_n8461_), .A2(new_n3837_), .A3(new_n4240_), .ZN(new_n15327_));
  NAND2_X1   g15008(.A1(\a[40] ), .A2(\a[60] ), .ZN(new_n15328_));
  NOR2_X1    g15009(.A1(new_n14732_), .A2(new_n15328_), .ZN(new_n15329_));
  AOI21_X1   g15010(.A1(new_n15327_), .A2(new_n15329_), .B(new_n8996_), .ZN(new_n15330_));
  OAI21_X1   g15011(.A1(new_n15330_), .A2(new_n3839_), .B(new_n15124_), .ZN(new_n15331_));
  INV_X1     g15012(.I(new_n15331_), .ZN(new_n15332_));
  AOI21_X1   g15013(.A1(new_n3838_), .A2(new_n8996_), .B(new_n15327_), .ZN(new_n15333_));
  INV_X1     g15014(.I(new_n15333_), .ZN(new_n15334_));
  NOR3_X1    g15015(.A1(new_n15334_), .A2(new_n8460_), .A3(new_n15147_), .ZN(new_n15335_));
  XNOR2_X1   g15016(.A1(new_n5339_), .A2(new_n8245_), .ZN(new_n15336_));
  NOR3_X1    g15017(.A1(new_n15335_), .A2(new_n15332_), .A3(new_n15336_), .ZN(new_n15337_));
  NOR2_X1    g15018(.A1(new_n15335_), .A2(new_n15332_), .ZN(new_n15338_));
  INV_X1     g15019(.I(new_n15336_), .ZN(new_n15339_));
  NOR2_X1    g15020(.A1(new_n15338_), .A2(new_n15339_), .ZN(new_n15340_));
  OAI21_X1   g15021(.A1(new_n15337_), .A2(new_n15340_), .B(new_n15326_), .ZN(new_n15341_));
  INV_X1     g15022(.I(new_n15326_), .ZN(new_n15342_));
  XOR2_X1    g15023(.A1(new_n15338_), .A2(new_n15339_), .Z(new_n15343_));
  NAND2_X1   g15024(.A1(new_n15342_), .A2(new_n15343_), .ZN(new_n15344_));
  NAND2_X1   g15025(.A1(new_n15211_), .A2(new_n15208_), .ZN(new_n15345_));
  AOI22_X1   g15026(.A1(new_n15344_), .A2(new_n15341_), .B1(new_n15210_), .B2(new_n15345_), .ZN(new_n15346_));
  INV_X1     g15027(.I(new_n15346_), .ZN(new_n15347_));
  NAND2_X1   g15028(.A1(new_n15344_), .A2(new_n15341_), .ZN(new_n15348_));
  NAND2_X1   g15029(.A1(new_n15345_), .A2(new_n15210_), .ZN(new_n15349_));
  NOR2_X1    g15030(.A1(new_n15348_), .A2(new_n15349_), .ZN(new_n15350_));
  INV_X1     g15031(.I(new_n15350_), .ZN(new_n15351_));
  AOI21_X1   g15032(.A1(new_n15351_), .A2(new_n15347_), .B(new_n15317_), .ZN(new_n15352_));
  XOR2_X1    g15033(.A1(new_n15348_), .A2(new_n15349_), .Z(new_n15353_));
  AOI21_X1   g15034(.A1(new_n15317_), .A2(new_n15353_), .B(new_n15352_), .ZN(new_n15354_));
  NOR2_X1    g15035(.A1(new_n15316_), .A2(new_n15354_), .ZN(new_n15355_));
  INV_X1     g15036(.I(new_n15355_), .ZN(new_n15356_));
  NAND2_X1   g15037(.A1(new_n15316_), .A2(new_n15354_), .ZN(new_n15357_));
  AOI21_X1   g15038(.A1(new_n15356_), .A2(new_n15357_), .B(new_n15314_), .ZN(new_n15358_));
  XNOR2_X1   g15039(.A1(new_n15316_), .A2(new_n15354_), .ZN(new_n15359_));
  NOR3_X1    g15040(.A1(new_n15359_), .A2(new_n15308_), .A3(new_n15313_), .ZN(new_n15360_));
  NOR2_X1    g15041(.A1(new_n15358_), .A2(new_n15360_), .ZN(new_n15361_));
  AOI21_X1   g15042(.A1(new_n15112_), .A2(new_n15224_), .B(new_n15222_), .ZN(new_n15362_));
  XOR2_X1    g15043(.A1(new_n15361_), .A2(new_n15362_), .Z(new_n15363_));
  INV_X1     g15044(.I(new_n15361_), .ZN(new_n15364_));
  NOR2_X1    g15045(.A1(new_n15364_), .A2(new_n15362_), .ZN(new_n15365_));
  INV_X1     g15046(.I(new_n15362_), .ZN(new_n15366_));
  NOR2_X1    g15047(.A1(new_n15366_), .A2(new_n15361_), .ZN(new_n15367_));
  OAI21_X1   g15048(.A1(new_n15365_), .A2(new_n15367_), .B(new_n15237_), .ZN(new_n15368_));
  OAI21_X1   g15049(.A1(new_n15237_), .A2(new_n15363_), .B(new_n15368_), .ZN(\asquared[97] ));
  NAND2_X1   g15050(.A1(new_n15364_), .A2(new_n15362_), .ZN(new_n15370_));
  OAI21_X1   g15051(.A1(new_n15236_), .A2(new_n15365_), .B(new_n15370_), .ZN(new_n15371_));
  NAND2_X1   g15052(.A1(new_n15314_), .A2(new_n15357_), .ZN(new_n15372_));
  NAND2_X1   g15053(.A1(new_n15372_), .A2(new_n15356_), .ZN(new_n15373_));
  NOR2_X1    g15054(.A1(new_n15239_), .A2(new_n15310_), .ZN(new_n15374_));
  NOR2_X1    g15055(.A1(new_n15374_), .A2(new_n15311_), .ZN(new_n15375_));
  INV_X1     g15056(.I(new_n15375_), .ZN(new_n15376_));
  OAI21_X1   g15057(.A1(new_n15317_), .A2(new_n15350_), .B(new_n15347_), .ZN(new_n15377_));
  NOR2_X1    g15058(.A1(new_n15342_), .A2(new_n15340_), .ZN(new_n15378_));
  NOR2_X1    g15059(.A1(new_n15378_), .A2(new_n15337_), .ZN(new_n15379_));
  OAI21_X1   g15060(.A1(new_n5340_), .A2(new_n8565_), .B(new_n8246_), .ZN(new_n15380_));
  NAND2_X1   g15061(.A1(new_n15322_), .A2(new_n15380_), .ZN(new_n15381_));
  XOR2_X1    g15062(.A1(new_n15381_), .A2(\a[36] ), .Z(new_n15382_));
  XOR2_X1    g15063(.A1(new_n15382_), .A2(\a[61] ), .Z(new_n15383_));
  INV_X1     g15064(.I(new_n15270_), .ZN(new_n15384_));
  AOI21_X1   g15065(.A1(new_n15260_), .A2(new_n15384_), .B(new_n15269_), .ZN(new_n15385_));
  XOR2_X1    g15066(.A1(new_n15383_), .A2(new_n15385_), .Z(new_n15386_));
  NOR2_X1    g15067(.A1(new_n15386_), .A2(new_n15379_), .ZN(new_n15387_));
  INV_X1     g15068(.I(new_n15379_), .ZN(new_n15388_));
  INV_X1     g15069(.I(new_n15383_), .ZN(new_n15389_));
  NOR2_X1    g15070(.A1(new_n15389_), .A2(new_n15385_), .ZN(new_n15390_));
  INV_X1     g15071(.I(new_n15390_), .ZN(new_n15391_));
  NAND2_X1   g15072(.A1(new_n15389_), .A2(new_n15385_), .ZN(new_n15392_));
  AOI21_X1   g15073(.A1(new_n15391_), .A2(new_n15392_), .B(new_n15388_), .ZN(new_n15393_));
  NOR2_X1    g15074(.A1(new_n15393_), .A2(new_n15387_), .ZN(new_n15394_));
  AOI21_X1   g15075(.A1(new_n15241_), .A2(new_n15254_), .B(new_n15252_), .ZN(new_n15395_));
  INV_X1     g15076(.I(new_n15293_), .ZN(new_n15396_));
  AOI21_X1   g15077(.A1(new_n15284_), .A2(new_n15396_), .B(new_n15292_), .ZN(new_n15397_));
  NAND2_X1   g15078(.A1(new_n6779_), .A2(new_n5980_), .ZN(new_n15398_));
  NOR2_X1    g15079(.A1(new_n4240_), .A2(new_n7727_), .ZN(new_n15399_));
  XOR2_X1    g15080(.A1(new_n15398_), .A2(new_n15399_), .Z(new_n15400_));
  NAND2_X1   g15081(.A1(\a[35] ), .A2(\a[49] ), .ZN(new_n15401_));
  NAND2_X1   g15082(.A1(\a[48] ), .A2(\a[62] ), .ZN(new_n15402_));
  XNOR2_X1   g15083(.A1(new_n15401_), .A2(new_n15402_), .ZN(new_n15403_));
  XNOR2_X1   g15084(.A1(new_n15400_), .A2(new_n15403_), .ZN(new_n15404_));
  NOR2_X1    g15085(.A1(new_n15397_), .A2(new_n15404_), .ZN(new_n15405_));
  NOR2_X1    g15086(.A1(new_n15400_), .A2(new_n15403_), .ZN(new_n15406_));
  INV_X1     g15087(.I(new_n15406_), .ZN(new_n15407_));
  NAND2_X1   g15088(.A1(new_n15400_), .A2(new_n15403_), .ZN(new_n15408_));
  NAND2_X1   g15089(.A1(new_n15407_), .A2(new_n15408_), .ZN(new_n15409_));
  AOI21_X1   g15090(.A1(new_n15397_), .A2(new_n15409_), .B(new_n15405_), .ZN(new_n15410_));
  NOR2_X1    g15091(.A1(new_n15244_), .A2(new_n15242_), .ZN(new_n15411_));
  AOI21_X1   g15092(.A1(new_n3487_), .A2(new_n9784_), .B(new_n15246_), .ZN(new_n15412_));
  XOR2_X1    g15093(.A1(new_n15411_), .A2(new_n15412_), .Z(new_n15413_));
  INV_X1     g15094(.I(new_n15411_), .ZN(new_n15414_));
  INV_X1     g15095(.I(new_n15412_), .ZN(new_n15415_));
  NOR2_X1    g15096(.A1(new_n15414_), .A2(new_n15415_), .ZN(new_n15416_));
  NOR2_X1    g15097(.A1(new_n15411_), .A2(new_n15412_), .ZN(new_n15417_));
  NOR2_X1    g15098(.A1(new_n15416_), .A2(new_n15417_), .ZN(new_n15418_));
  NOR2_X1    g15099(.A1(new_n15418_), .A2(new_n15333_), .ZN(new_n15419_));
  AOI21_X1   g15100(.A1(new_n15333_), .A2(new_n15413_), .B(new_n15419_), .ZN(new_n15420_));
  XNOR2_X1   g15101(.A1(new_n15420_), .A2(new_n15410_), .ZN(new_n15421_));
  NOR2_X1    g15102(.A1(new_n15420_), .A2(new_n15410_), .ZN(new_n15422_));
  NAND2_X1   g15103(.A1(new_n15420_), .A2(new_n15410_), .ZN(new_n15423_));
  INV_X1     g15104(.I(new_n15423_), .ZN(new_n15424_));
  OAI21_X1   g15105(.A1(new_n15424_), .A2(new_n15422_), .B(new_n15395_), .ZN(new_n15425_));
  OAI21_X1   g15106(.A1(new_n15395_), .A2(new_n15421_), .B(new_n15425_), .ZN(new_n15426_));
  INV_X1     g15107(.I(new_n15426_), .ZN(new_n15427_));
  XOR2_X1    g15108(.A1(new_n15394_), .A2(new_n15427_), .Z(new_n15428_));
  NOR2_X1    g15109(.A1(new_n15394_), .A2(new_n15427_), .ZN(new_n15429_));
  INV_X1     g15110(.I(new_n15429_), .ZN(new_n15430_));
  NAND2_X1   g15111(.A1(new_n15394_), .A2(new_n15427_), .ZN(new_n15431_));
  NAND2_X1   g15112(.A1(new_n15430_), .A2(new_n15431_), .ZN(new_n15432_));
  MUX2_X1    g15113(.I0(new_n15432_), .I1(new_n15428_), .S(new_n15377_), .Z(new_n15433_));
  OAI21_X1   g15114(.A1(new_n15257_), .A2(new_n15273_), .B(new_n15274_), .ZN(new_n15434_));
  INV_X1     g15115(.I(new_n15434_), .ZN(new_n15435_));
  NOR2_X1    g15116(.A1(new_n15303_), .A2(new_n15279_), .ZN(new_n15436_));
  NOR2_X1    g15117(.A1(new_n15436_), .A2(new_n15302_), .ZN(new_n15437_));
  NAND4_X1   g15118(.A1(\a[41] ), .A2(\a[42] ), .A3(\a[55] ), .A4(\a[56] ), .ZN(new_n15439_));
  AOI22_X1   g15119(.A1(new_n5601_), .A2(new_n8996_), .B1(new_n9554_), .B2(new_n5600_), .ZN(new_n15440_));
  NOR4_X1    g15120(.A1(new_n5339_), .A2(new_n8676_), .A3(new_n3837_), .A4(new_n8990_), .ZN(new_n15441_));
  NAND2_X1   g15121(.A1(new_n15440_), .A2(new_n15441_), .ZN(new_n15442_));
  INV_X1     g15122(.I(new_n15442_), .ZN(new_n15443_));
  INV_X1     g15123(.I(new_n8767_), .ZN(new_n15444_));
  NOR2_X1    g15124(.A1(new_n7187_), .A2(new_n5322_), .ZN(new_n15445_));
  NOR2_X1    g15125(.A1(new_n10291_), .A2(new_n15445_), .ZN(new_n15446_));
  INV_X1     g15126(.I(new_n15446_), .ZN(new_n15447_));
  NOR4_X1    g15127(.A1(new_n15447_), .A2(new_n5742_), .A3(new_n7204_), .A4(new_n15444_), .ZN(new_n15448_));
  AND2_X2    g15128(.A1(new_n15448_), .A2(new_n15443_), .Z(new_n15449_));
  NOR2_X1    g15129(.A1(new_n15448_), .A2(new_n15443_), .ZN(new_n15450_));
  NOR2_X1    g15130(.A1(new_n15449_), .A2(new_n15450_), .ZN(new_n15451_));
  NOR2_X1    g15131(.A1(new_n15451_), .A2(new_n15439_), .ZN(new_n15452_));
  XOR2_X1    g15132(.A1(new_n15448_), .A2(new_n15443_), .Z(new_n15453_));
  AOI21_X1   g15133(.A1(new_n15453_), .A2(new_n15439_), .B(new_n15452_), .ZN(new_n15454_));
  OR2_X2     g15134(.A1(new_n15437_), .A2(new_n15454_), .Z(new_n15455_));
  NAND2_X1   g15135(.A1(new_n15437_), .A2(new_n15454_), .ZN(new_n15456_));
  AOI21_X1   g15136(.A1(new_n15455_), .A2(new_n15456_), .B(new_n15435_), .ZN(new_n15457_));
  XOR2_X1    g15137(.A1(new_n15437_), .A2(new_n15454_), .Z(new_n15458_));
  AOI21_X1   g15138(.A1(new_n15435_), .A2(new_n15458_), .B(new_n15457_), .ZN(new_n15459_));
  XOR2_X1    g15139(.A1(new_n15433_), .A2(new_n15459_), .Z(new_n15460_));
  OR2_X2     g15140(.A1(new_n15433_), .A2(new_n15459_), .Z(new_n15461_));
  NAND2_X1   g15141(.A1(new_n15433_), .A2(new_n15459_), .ZN(new_n15462_));
  AOI21_X1   g15142(.A1(new_n15461_), .A2(new_n15462_), .B(new_n15376_), .ZN(new_n15463_));
  AOI21_X1   g15143(.A1(new_n15376_), .A2(new_n15460_), .B(new_n15463_), .ZN(new_n15464_));
  XNOR2_X1   g15144(.A1(new_n15464_), .A2(new_n15373_), .ZN(new_n15465_));
  NOR2_X1    g15145(.A1(new_n15464_), .A2(new_n15373_), .ZN(new_n15466_));
  NAND2_X1   g15146(.A1(new_n15464_), .A2(new_n15373_), .ZN(new_n15467_));
  INV_X1     g15147(.I(new_n15467_), .ZN(new_n15468_));
  OAI21_X1   g15148(.A1(new_n15466_), .A2(new_n15468_), .B(new_n15371_), .ZN(new_n15469_));
  OAI21_X1   g15149(.A1(new_n15371_), .A2(new_n15465_), .B(new_n15469_), .ZN(\asquared[98] ));
  NAND3_X1   g15150(.A1(new_n15236_), .A2(new_n15361_), .A3(new_n15366_), .ZN(new_n15471_));
  NAND2_X1   g15151(.A1(new_n15462_), .A2(new_n15376_), .ZN(new_n15472_));
  NAND2_X1   g15152(.A1(new_n15472_), .A2(new_n15461_), .ZN(new_n15473_));
  NAND2_X1   g15153(.A1(new_n15434_), .A2(new_n15456_), .ZN(new_n15474_));
  NAND2_X1   g15154(.A1(new_n15474_), .A2(new_n15455_), .ZN(new_n15475_));
  AOI22_X1   g15155(.A1(new_n6776_), .A2(new_n8198_), .B1(new_n6777_), .B2(new_n5980_), .ZN(new_n15476_));
  INV_X1     g15156(.I(new_n15476_), .ZN(new_n15477_));
  NOR2_X1    g15157(.A1(new_n7693_), .A2(new_n8941_), .ZN(new_n15478_));
  NOR2_X1    g15158(.A1(new_n15477_), .A2(new_n15478_), .ZN(new_n15479_));
  AOI21_X1   g15159(.A1(new_n15479_), .A2(new_n6056_), .B(\a[51] ), .ZN(new_n15480_));
  NOR2_X1    g15160(.A1(\a[46] ), .A2(\a[52] ), .ZN(new_n15481_));
  OAI21_X1   g15161(.A1(new_n15480_), .A2(new_n5511_), .B(new_n15481_), .ZN(new_n15482_));
  NOR2_X1    g15162(.A1(new_n15478_), .A2(new_n15476_), .ZN(new_n15483_));
  AND2_X2    g15163(.A1(new_n15482_), .A2(new_n15483_), .Z(new_n15484_));
  INV_X1     g15164(.I(new_n15484_), .ZN(new_n15485_));
  NAND2_X1   g15165(.A1(new_n8676_), .A2(new_n6024_), .ZN(new_n15486_));
  NAND2_X1   g15166(.A1(\a[45] ), .A2(\a[53] ), .ZN(new_n15487_));
  XNOR2_X1   g15167(.A1(new_n15486_), .A2(new_n15487_), .ZN(new_n15488_));
  INV_X1     g15168(.I(new_n15488_), .ZN(new_n15489_));
  AOI21_X1   g15169(.A1(new_n12355_), .A2(new_n9029_), .B(new_n3423_), .ZN(new_n15490_));
  NOR2_X1    g15170(.A1(new_n3393_), .A2(new_n8453_), .ZN(new_n15491_));
  XOR2_X1    g15171(.A1(new_n15491_), .A2(new_n11834_), .Z(new_n15492_));
  XNOR2_X1   g15172(.A1(new_n15492_), .A2(new_n15490_), .ZN(new_n15493_));
  NOR2_X1    g15173(.A1(new_n15493_), .A2(new_n15489_), .ZN(new_n15494_));
  INV_X1     g15174(.I(new_n15493_), .ZN(new_n15495_));
  NOR2_X1    g15175(.A1(new_n15495_), .A2(new_n15488_), .ZN(new_n15496_));
  NOR2_X1    g15176(.A1(new_n15496_), .A2(new_n15494_), .ZN(new_n15497_));
  NOR2_X1    g15177(.A1(new_n15485_), .A2(new_n15497_), .ZN(new_n15498_));
  XOR2_X1    g15178(.A1(new_n15493_), .A2(new_n15488_), .Z(new_n15499_));
  NOR2_X1    g15179(.A1(new_n15484_), .A2(new_n15499_), .ZN(new_n15500_));
  NOR2_X1    g15180(.A1(new_n15498_), .A2(new_n15500_), .ZN(new_n15501_));
  INV_X1     g15181(.I(new_n15408_), .ZN(new_n15502_));
  OAI21_X1   g15182(.A1(new_n15397_), .A2(new_n15502_), .B(new_n15407_), .ZN(new_n15503_));
  NOR4_X1    g15183(.A1(new_n4414_), .A2(new_n4769_), .A3(new_n6999_), .A4(new_n7216_), .ZN(new_n15504_));
  AOI21_X1   g15184(.A1(new_n5339_), .A2(new_n8676_), .B(new_n15440_), .ZN(new_n15505_));
  AOI21_X1   g15185(.A1(new_n5742_), .A2(new_n7204_), .B(new_n15446_), .ZN(new_n15506_));
  XOR2_X1    g15186(.A1(new_n15506_), .A2(new_n15505_), .Z(new_n15507_));
  INV_X1     g15187(.I(new_n15505_), .ZN(new_n15508_));
  INV_X1     g15188(.I(new_n15506_), .ZN(new_n15509_));
  NOR2_X1    g15189(.A1(new_n15509_), .A2(new_n15508_), .ZN(new_n15510_));
  NOR2_X1    g15190(.A1(new_n15506_), .A2(new_n15505_), .ZN(new_n15511_));
  NOR2_X1    g15191(.A1(new_n15510_), .A2(new_n15511_), .ZN(new_n15512_));
  NOR2_X1    g15192(.A1(new_n15512_), .A2(new_n15504_), .ZN(new_n15513_));
  AOI21_X1   g15193(.A1(new_n15504_), .A2(new_n15507_), .B(new_n15513_), .ZN(new_n15514_));
  NOR2_X1    g15194(.A1(new_n15514_), .A2(new_n15503_), .ZN(new_n15515_));
  INV_X1     g15195(.I(new_n15515_), .ZN(new_n15516_));
  NAND2_X1   g15196(.A1(new_n15514_), .A2(new_n15503_), .ZN(new_n15517_));
  AOI21_X1   g15197(.A1(new_n15516_), .A2(new_n15517_), .B(new_n15501_), .ZN(new_n15518_));
  XNOR2_X1   g15198(.A1(new_n15514_), .A2(new_n15503_), .ZN(new_n15519_));
  NOR3_X1    g15199(.A1(new_n15519_), .A2(new_n15498_), .A3(new_n15500_), .ZN(new_n15520_));
  NOR2_X1    g15200(.A1(new_n15520_), .A2(new_n15518_), .ZN(new_n15521_));
  INV_X1     g15201(.I(new_n15521_), .ZN(new_n15522_));
  INV_X1     g15202(.I(new_n15417_), .ZN(new_n15523_));
  AOI21_X1   g15203(.A1(new_n15333_), .A2(new_n15523_), .B(new_n15416_), .ZN(new_n15524_));
  OAI21_X1   g15204(.A1(new_n15322_), .A2(new_n15380_), .B(new_n15491_), .ZN(new_n15525_));
  NAND2_X1   g15205(.A1(new_n15525_), .A2(new_n15381_), .ZN(new_n15526_));
  INV_X1     g15206(.I(new_n15526_), .ZN(new_n15527_));
  INV_X1     g15207(.I(new_n15449_), .ZN(new_n15528_));
  OR2_X2     g15208(.A1(new_n15450_), .A2(new_n15439_), .Z(new_n15529_));
  NAND2_X1   g15209(.A1(new_n15529_), .A2(new_n15528_), .ZN(new_n15530_));
  XOR2_X1    g15210(.A1(new_n15530_), .A2(new_n15527_), .Z(new_n15531_));
  NOR2_X1    g15211(.A1(new_n15531_), .A2(new_n15524_), .ZN(new_n15532_));
  INV_X1     g15212(.I(new_n15524_), .ZN(new_n15533_));
  INV_X1     g15213(.I(new_n15530_), .ZN(new_n15534_));
  NOR2_X1    g15214(.A1(new_n15534_), .A2(new_n15527_), .ZN(new_n15535_));
  NOR2_X1    g15215(.A1(new_n15530_), .A2(new_n15526_), .ZN(new_n15536_));
  NOR2_X1    g15216(.A1(new_n15535_), .A2(new_n15536_), .ZN(new_n15537_));
  NOR2_X1    g15217(.A1(new_n15537_), .A2(new_n15533_), .ZN(new_n15538_));
  NOR2_X1    g15218(.A1(new_n15538_), .A2(new_n15532_), .ZN(new_n15539_));
  NOR2_X1    g15219(.A1(new_n15522_), .A2(new_n15539_), .ZN(new_n15540_));
  INV_X1     g15220(.I(new_n15539_), .ZN(new_n15541_));
  NOR2_X1    g15221(.A1(new_n15521_), .A2(new_n15541_), .ZN(new_n15542_));
  OAI21_X1   g15222(.A1(new_n15540_), .A2(new_n15542_), .B(new_n15475_), .ZN(new_n15543_));
  XOR2_X1    g15223(.A1(new_n15521_), .A2(new_n15539_), .Z(new_n15544_));
  OAI21_X1   g15224(.A1(new_n15475_), .A2(new_n15544_), .B(new_n15543_), .ZN(new_n15545_));
  INV_X1     g15225(.I(new_n15545_), .ZN(new_n15546_));
  NAND2_X1   g15226(.A1(new_n15430_), .A2(new_n15377_), .ZN(new_n15547_));
  NAND2_X1   g15227(.A1(new_n15547_), .A2(new_n15431_), .ZN(new_n15548_));
  AOI21_X1   g15228(.A1(new_n15388_), .A2(new_n15392_), .B(new_n15390_), .ZN(new_n15549_));
  INV_X1     g15229(.I(new_n15549_), .ZN(new_n15550_));
  OAI21_X1   g15230(.A1(new_n15395_), .A2(new_n15422_), .B(new_n15423_), .ZN(new_n15551_));
  NAND2_X1   g15231(.A1(new_n6779_), .A2(new_n5980_), .ZN(new_n15552_));
  NOR2_X1    g15232(.A1(new_n6779_), .A2(new_n5980_), .ZN(new_n15553_));
  NOR2_X1    g15233(.A1(\a[40] ), .A2(\a[57] ), .ZN(new_n15554_));
  AOI21_X1   g15234(.A1(new_n15552_), .A2(new_n15554_), .B(new_n15553_), .ZN(new_n15555_));
  INV_X1     g15235(.I(new_n15555_), .ZN(new_n15556_));
  XNOR2_X1   g15236(.A1(new_n8767_), .A2(new_n8955_), .ZN(new_n15557_));
  NOR2_X1    g15237(.A1(new_n3423_), .A2(new_n9310_), .ZN(new_n15558_));
  NOR2_X1    g15238(.A1(new_n15557_), .A2(new_n15558_), .ZN(new_n15559_));
  INV_X1     g15239(.I(new_n15557_), .ZN(new_n15560_));
  NOR3_X1    g15240(.A1(new_n15560_), .A2(new_n3423_), .A3(new_n9310_), .ZN(new_n15561_));
  NOR2_X1    g15241(.A1(new_n15561_), .A2(new_n15559_), .ZN(new_n15562_));
  INV_X1     g15242(.I(new_n15562_), .ZN(new_n15563_));
  NOR2_X1    g15243(.A1(new_n3804_), .A2(new_n8990_), .ZN(new_n15564_));
  XNOR2_X1   g15244(.A1(new_n5350_), .A2(new_n8242_), .ZN(new_n15565_));
  NOR2_X1    g15245(.A1(new_n15563_), .A2(new_n15565_), .ZN(new_n15566_));
  INV_X1     g15246(.I(new_n15565_), .ZN(new_n15567_));
  NOR2_X1    g15247(.A1(new_n15562_), .A2(new_n15567_), .ZN(new_n15568_));
  NOR2_X1    g15248(.A1(new_n15566_), .A2(new_n15568_), .ZN(new_n15569_));
  NOR2_X1    g15249(.A1(new_n15569_), .A2(new_n15556_), .ZN(new_n15570_));
  XOR2_X1    g15250(.A1(new_n15562_), .A2(new_n15565_), .Z(new_n15571_));
  NOR2_X1    g15251(.A1(new_n15571_), .A2(new_n15555_), .ZN(new_n15572_));
  NOR2_X1    g15252(.A1(new_n15570_), .A2(new_n15572_), .ZN(new_n15573_));
  INV_X1     g15253(.I(new_n15573_), .ZN(new_n15574_));
  XOR2_X1    g15254(.A1(new_n15551_), .A2(new_n15574_), .Z(new_n15575_));
  NAND2_X1   g15255(.A1(new_n15575_), .A2(new_n15550_), .ZN(new_n15576_));
  AND2_X2    g15256(.A1(new_n15551_), .A2(new_n15574_), .Z(new_n15577_));
  NOR2_X1    g15257(.A1(new_n15551_), .A2(new_n15574_), .ZN(new_n15578_));
  OAI21_X1   g15258(.A1(new_n15578_), .A2(new_n15577_), .B(new_n15549_), .ZN(new_n15579_));
  NAND2_X1   g15259(.A1(new_n15576_), .A2(new_n15579_), .ZN(new_n15580_));
  XOR2_X1    g15260(.A1(new_n15548_), .A2(new_n15580_), .Z(new_n15581_));
  INV_X1     g15261(.I(new_n15580_), .ZN(new_n15582_));
  NOR2_X1    g15262(.A1(new_n15548_), .A2(new_n15582_), .ZN(new_n15583_));
  NAND2_X1   g15263(.A1(new_n15548_), .A2(new_n15582_), .ZN(new_n15584_));
  INV_X1     g15264(.I(new_n15584_), .ZN(new_n15585_));
  OAI21_X1   g15265(.A1(new_n15585_), .A2(new_n15583_), .B(new_n15546_), .ZN(new_n15586_));
  OAI21_X1   g15266(.A1(new_n15546_), .A2(new_n15581_), .B(new_n15586_), .ZN(new_n15587_));
  NAND2_X1   g15267(.A1(new_n15587_), .A2(new_n15473_), .ZN(new_n15588_));
  XOR2_X1    g15268(.A1(new_n15471_), .A2(new_n15588_), .Z(new_n15589_));
  XOR2_X1    g15269(.A1(new_n15589_), .A2(new_n15466_), .Z(\asquared[99] ));
  OAI21_X1   g15270(.A1(new_n15473_), .A2(new_n15587_), .B(new_n15466_), .ZN(new_n15591_));
  OAI21_X1   g15271(.A1(new_n15471_), .A2(new_n15591_), .B(new_n15588_), .ZN(new_n15592_));
  INV_X1     g15272(.I(new_n15592_), .ZN(new_n15593_));
  NOR2_X1    g15273(.A1(new_n15549_), .A2(new_n15578_), .ZN(new_n15594_));
  NOR2_X1    g15274(.A1(new_n15594_), .A2(new_n15577_), .ZN(new_n15595_));
  INV_X1     g15275(.I(new_n15494_), .ZN(new_n15596_));
  AOI21_X1   g15276(.A1(new_n15484_), .A2(new_n15596_), .B(new_n15496_), .ZN(new_n15597_));
  NOR2_X1    g15277(.A1(new_n3393_), .A2(new_n3783_), .ZN(new_n15598_));
  AOI22_X1   g15278(.A1(new_n3805_), .A2(new_n9781_), .B1(new_n11018_), .B2(new_n15598_), .ZN(new_n15599_));
  INV_X1     g15279(.I(new_n15599_), .ZN(new_n15600_));
  NOR2_X1    g15280(.A1(new_n3393_), .A2(new_n9310_), .ZN(new_n15601_));
  NAND4_X1   g15281(.A1(new_n15600_), .A2(new_n5340_), .A3(new_n8992_), .A4(new_n15601_), .ZN(new_n15602_));
  AOI21_X1   g15282(.A1(new_n5350_), .A2(new_n15564_), .B(new_n8242_), .ZN(new_n15603_));
  NAND2_X1   g15283(.A1(new_n15490_), .A2(new_n9784_), .ZN(new_n15604_));
  OAI21_X1   g15284(.A1(new_n3839_), .A2(new_n15492_), .B(new_n15604_), .ZN(new_n15605_));
  INV_X1     g15285(.I(new_n15605_), .ZN(new_n15606_));
  NOR2_X1    g15286(.A1(new_n15606_), .A2(new_n15603_), .ZN(new_n15607_));
  INV_X1     g15287(.I(new_n15607_), .ZN(new_n15608_));
  NAND2_X1   g15288(.A1(new_n15606_), .A2(new_n15603_), .ZN(new_n15609_));
  AOI21_X1   g15289(.A1(new_n15608_), .A2(new_n15609_), .B(new_n15602_), .ZN(new_n15610_));
  INV_X1     g15290(.I(new_n15602_), .ZN(new_n15611_));
  XOR2_X1    g15291(.A1(new_n15605_), .A2(new_n15603_), .Z(new_n15612_));
  NOR2_X1    g15292(.A1(new_n15612_), .A2(new_n15611_), .ZN(new_n15613_));
  NOR2_X1    g15293(.A1(new_n15610_), .A2(new_n15613_), .ZN(new_n15614_));
  INV_X1     g15294(.I(new_n15614_), .ZN(new_n15615_));
  NAND2_X1   g15295(.A1(new_n8676_), .A2(new_n6024_), .ZN(new_n15616_));
  NOR2_X1    g15296(.A1(new_n8676_), .A2(new_n6024_), .ZN(new_n15617_));
  NOR2_X1    g15297(.A1(\a[45] ), .A2(\a[53] ), .ZN(new_n15618_));
  AOI21_X1   g15298(.A1(new_n15616_), .A2(new_n15618_), .B(new_n15617_), .ZN(new_n15619_));
  INV_X1     g15299(.I(new_n15479_), .ZN(new_n15620_));
  AOI22_X1   g15300(.A1(new_n15560_), .A2(new_n15558_), .B1(new_n5321_), .B2(new_n7483_), .ZN(new_n15621_));
  XOR2_X1    g15301(.A1(new_n15621_), .A2(new_n15620_), .Z(new_n15622_));
  INV_X1     g15302(.I(new_n15621_), .ZN(new_n15623_));
  NOR2_X1    g15303(.A1(new_n15623_), .A2(new_n15620_), .ZN(new_n15624_));
  NOR2_X1    g15304(.A1(new_n15621_), .A2(new_n15479_), .ZN(new_n15625_));
  NOR2_X1    g15305(.A1(new_n15624_), .A2(new_n15625_), .ZN(new_n15626_));
  MUX2_X1    g15306(.I0(new_n15626_), .I1(new_n15622_), .S(new_n15619_), .Z(new_n15627_));
  NOR2_X1    g15307(.A1(new_n15615_), .A2(new_n15627_), .ZN(new_n15628_));
  INV_X1     g15308(.I(new_n15628_), .ZN(new_n15629_));
  NAND2_X1   g15309(.A1(new_n15615_), .A2(new_n15627_), .ZN(new_n15630_));
  AOI21_X1   g15310(.A1(new_n15629_), .A2(new_n15630_), .B(new_n15597_), .ZN(new_n15631_));
  INV_X1     g15311(.I(new_n15597_), .ZN(new_n15632_));
  XOR2_X1    g15312(.A1(new_n15627_), .A2(new_n15614_), .Z(new_n15633_));
  NOR2_X1    g15313(.A1(new_n15633_), .A2(new_n15632_), .ZN(new_n15634_));
  NOR2_X1    g15314(.A1(new_n15634_), .A2(new_n15631_), .ZN(new_n15635_));
  INV_X1     g15315(.I(new_n15511_), .ZN(new_n15636_));
  AOI21_X1   g15316(.A1(new_n15504_), .A2(new_n15636_), .B(new_n15510_), .ZN(new_n15637_));
  NOR2_X1    g15317(.A1(new_n15568_), .A2(new_n15556_), .ZN(new_n15638_));
  NOR2_X1    g15318(.A1(new_n15638_), .A2(new_n15566_), .ZN(new_n15639_));
  NAND2_X1   g15319(.A1(\a[49] ), .A2(\a[62] ), .ZN(new_n15640_));
  XOR2_X1    g15320(.A1(new_n14089_), .A2(new_n15640_), .Z(new_n15641_));
  XNOR2_X1   g15321(.A1(new_n15639_), .A2(new_n15641_), .ZN(new_n15642_));
  NOR2_X1    g15322(.A1(new_n15642_), .A2(new_n15637_), .ZN(new_n15643_));
  INV_X1     g15323(.I(new_n15637_), .ZN(new_n15644_));
  NOR2_X1    g15324(.A1(new_n15639_), .A2(new_n15641_), .ZN(new_n15645_));
  INV_X1     g15325(.I(new_n15645_), .ZN(new_n15646_));
  NAND2_X1   g15326(.A1(new_n15639_), .A2(new_n15641_), .ZN(new_n15647_));
  AOI21_X1   g15327(.A1(new_n15646_), .A2(new_n15647_), .B(new_n15644_), .ZN(new_n15648_));
  NOR2_X1    g15328(.A1(new_n15643_), .A2(new_n15648_), .ZN(new_n15649_));
  XOR2_X1    g15329(.A1(new_n15635_), .A2(new_n15649_), .Z(new_n15650_));
  NOR2_X1    g15330(.A1(new_n15595_), .A2(new_n15650_), .ZN(new_n15651_));
  INV_X1     g15331(.I(new_n15595_), .ZN(new_n15652_));
  INV_X1     g15332(.I(new_n15635_), .ZN(new_n15653_));
  NOR2_X1    g15333(.A1(new_n15653_), .A2(new_n15649_), .ZN(new_n15654_));
  INV_X1     g15334(.I(new_n15654_), .ZN(new_n15655_));
  NAND2_X1   g15335(.A1(new_n15653_), .A2(new_n15649_), .ZN(new_n15656_));
  AOI21_X1   g15336(.A1(new_n15655_), .A2(new_n15656_), .B(new_n15652_), .ZN(new_n15657_));
  NOR2_X1    g15337(.A1(new_n15657_), .A2(new_n15651_), .ZN(new_n15658_));
  INV_X1     g15338(.I(new_n15540_), .ZN(new_n15659_));
  AOI21_X1   g15339(.A1(new_n15659_), .A2(new_n15475_), .B(new_n15542_), .ZN(new_n15660_));
  OAI21_X1   g15340(.A1(new_n15501_), .A2(new_n15515_), .B(new_n15517_), .ZN(new_n15661_));
  NOR2_X1    g15341(.A1(new_n15536_), .A2(new_n15524_), .ZN(new_n15662_));
  NOR2_X1    g15342(.A1(new_n15662_), .A2(new_n15535_), .ZN(new_n15663_));
  NOR2_X1    g15343(.A1(new_n6999_), .A2(new_n8085_), .ZN(new_n15664_));
  AOI22_X1   g15344(.A1(new_n5592_), .A2(new_n8676_), .B1(new_n6772_), .B2(new_n15664_), .ZN(new_n15665_));
  NOR2_X1    g15345(.A1(new_n4414_), .A2(new_n7647_), .ZN(new_n15666_));
  AOI21_X1   g15346(.A1(new_n8956_), .A2(new_n15666_), .B(new_n15665_), .ZN(new_n15667_));
  INV_X1     g15347(.I(new_n15667_), .ZN(new_n15668_));
  XNOR2_X1   g15348(.A1(new_n8955_), .A2(new_n15666_), .ZN(new_n15669_));
  OAI21_X1   g15349(.A1(new_n4240_), .A2(new_n8085_), .B(new_n15669_), .ZN(new_n15670_));
  AND2_X2    g15350(.A1(new_n15670_), .A2(new_n15668_), .Z(new_n15671_));
  INV_X1     g15351(.I(new_n15671_), .ZN(new_n15672_));
  NOR2_X1    g15352(.A1(new_n8026_), .A2(new_n8424_), .ZN(new_n15673_));
  NOR2_X1    g15353(.A1(new_n10291_), .A2(new_n15673_), .ZN(new_n15674_));
  NOR4_X1    g15354(.A1(new_n7204_), .A2(new_n5980_), .A3(new_n5004_), .A4(new_n6945_), .ZN(new_n15675_));
  NAND2_X1   g15355(.A1(new_n15674_), .A2(new_n15675_), .ZN(new_n15676_));
  NOR2_X1    g15356(.A1(new_n5750_), .A2(new_n6260_), .ZN(new_n15677_));
  XNOR2_X1   g15357(.A1(new_n5173_), .A2(new_n8242_), .ZN(new_n15678_));
  NOR2_X1    g15358(.A1(new_n15676_), .A2(new_n15678_), .ZN(new_n15679_));
  INV_X1     g15359(.I(new_n15678_), .ZN(new_n15680_));
  AOI21_X1   g15360(.A1(new_n15674_), .A2(new_n15675_), .B(new_n15680_), .ZN(new_n15681_));
  NOR2_X1    g15361(.A1(new_n15679_), .A2(new_n15681_), .ZN(new_n15682_));
  NOR2_X1    g15362(.A1(new_n15682_), .A2(new_n15672_), .ZN(new_n15683_));
  XOR2_X1    g15363(.A1(new_n15676_), .A2(new_n15680_), .Z(new_n15684_));
  NOR2_X1    g15364(.A1(new_n15684_), .A2(new_n15671_), .ZN(new_n15685_));
  NOR2_X1    g15365(.A1(new_n15683_), .A2(new_n15685_), .ZN(new_n15686_));
  XNOR2_X1   g15366(.A1(new_n15663_), .A2(new_n15686_), .ZN(new_n15687_));
  INV_X1     g15367(.I(new_n15687_), .ZN(new_n15688_));
  NOR2_X1    g15368(.A1(new_n15663_), .A2(new_n15686_), .ZN(new_n15689_));
  INV_X1     g15369(.I(new_n15689_), .ZN(new_n15690_));
  NAND2_X1   g15370(.A1(new_n15663_), .A2(new_n15686_), .ZN(new_n15691_));
  AOI21_X1   g15371(.A1(new_n15690_), .A2(new_n15691_), .B(new_n15661_), .ZN(new_n15692_));
  AOI21_X1   g15372(.A1(new_n15688_), .A2(new_n15661_), .B(new_n15692_), .ZN(new_n15693_));
  INV_X1     g15373(.I(new_n15693_), .ZN(new_n15694_));
  AND2_X2    g15374(.A1(new_n15660_), .A2(new_n15694_), .Z(new_n15695_));
  NOR2_X1    g15375(.A1(new_n15660_), .A2(new_n15694_), .ZN(new_n15696_));
  NOR2_X1    g15376(.A1(new_n15695_), .A2(new_n15696_), .ZN(new_n15697_));
  NOR2_X1    g15377(.A1(new_n15697_), .A2(new_n15658_), .ZN(new_n15698_));
  XOR2_X1    g15378(.A1(new_n15660_), .A2(new_n15693_), .Z(new_n15699_));
  NOR3_X1    g15379(.A1(new_n15699_), .A2(new_n15651_), .A3(new_n15657_), .ZN(new_n15700_));
  NOR2_X1    g15380(.A1(new_n15698_), .A2(new_n15700_), .ZN(new_n15701_));
  OAI21_X1   g15381(.A1(new_n15546_), .A2(new_n15583_), .B(new_n15584_), .ZN(new_n15702_));
  XNOR2_X1   g15382(.A1(new_n15701_), .A2(new_n15702_), .ZN(new_n15703_));
  NAND2_X1   g15383(.A1(new_n15701_), .A2(new_n15702_), .ZN(new_n15704_));
  NOR2_X1    g15384(.A1(new_n15701_), .A2(new_n15702_), .ZN(new_n15705_));
  INV_X1     g15385(.I(new_n15705_), .ZN(new_n15706_));
  NAND2_X1   g15386(.A1(new_n15706_), .A2(new_n15704_), .ZN(new_n15707_));
  NAND2_X1   g15387(.A1(new_n15593_), .A2(new_n15707_), .ZN(new_n15708_));
  OAI21_X1   g15388(.A1(new_n15593_), .A2(new_n15703_), .B(new_n15708_), .ZN(\asquared[100] ));
  OAI21_X1   g15389(.A1(new_n15593_), .A2(new_n15705_), .B(new_n15704_), .ZN(new_n15710_));
  INV_X1     g15390(.I(new_n15695_), .ZN(new_n15711_));
  AOI21_X1   g15391(.A1(new_n15711_), .A2(new_n15658_), .B(new_n15696_), .ZN(new_n15712_));
  INV_X1     g15392(.I(new_n15712_), .ZN(new_n15713_));
  OAI21_X1   g15393(.A1(new_n15595_), .A2(new_n15654_), .B(new_n15656_), .ZN(new_n15714_));
  AOI21_X1   g15394(.A1(new_n15661_), .A2(new_n15691_), .B(new_n15689_), .ZN(new_n15715_));
  OAI22_X1   g15395(.A1(new_n14719_), .A2(new_n7693_), .B1(new_n7001_), .B2(new_n8056_), .ZN(new_n15716_));
  OAI21_X1   g15396(.A1(new_n12355_), .A2(new_n10034_), .B(new_n15716_), .ZN(new_n15717_));
  INV_X1     g15397(.I(new_n15717_), .ZN(new_n15718_));
  AOI21_X1   g15398(.A1(new_n15718_), .A2(new_n9629_), .B(\a[52] ), .ZN(new_n15719_));
  NOR2_X1    g15399(.A1(\a[47] ), .A2(\a[53] ), .ZN(new_n15720_));
  OAI21_X1   g15400(.A1(new_n15719_), .A2(new_n5750_), .B(new_n15720_), .ZN(new_n15721_));
  AOI21_X1   g15401(.A1(new_n6028_), .A2(new_n6777_), .B(new_n15716_), .ZN(new_n15722_));
  AND2_X2    g15402(.A1(new_n15721_), .A2(new_n15722_), .Z(new_n15723_));
  INV_X1     g15403(.I(new_n15723_), .ZN(new_n15724_));
  AOI21_X1   g15404(.A1(new_n15611_), .A2(new_n15609_), .B(new_n15607_), .ZN(new_n15725_));
  INV_X1     g15405(.I(new_n15625_), .ZN(new_n15726_));
  AOI21_X1   g15406(.A1(new_n15619_), .A2(new_n15726_), .B(new_n15624_), .ZN(new_n15727_));
  XNOR2_X1   g15407(.A1(new_n15727_), .A2(new_n15725_), .ZN(new_n15728_));
  NOR2_X1    g15408(.A1(new_n15727_), .A2(new_n15725_), .ZN(new_n15729_));
  NAND2_X1   g15409(.A1(new_n15727_), .A2(new_n15725_), .ZN(new_n15730_));
  INV_X1     g15410(.I(new_n15730_), .ZN(new_n15731_));
  OAI21_X1   g15411(.A1(new_n15731_), .A2(new_n15729_), .B(new_n15724_), .ZN(new_n15732_));
  OAI21_X1   g15412(.A1(new_n15724_), .A2(new_n15728_), .B(new_n15732_), .ZN(new_n15733_));
  AOI21_X1   g15413(.A1(new_n5339_), .A2(new_n8991_), .B(new_n15600_), .ZN(new_n15734_));
  INV_X1     g15414(.I(new_n15734_), .ZN(new_n15735_));
  NAND2_X1   g15415(.A1(new_n8955_), .A2(new_n15666_), .ZN(new_n15736_));
  AND2_X2    g15416(.A1(new_n15665_), .A2(new_n15736_), .Z(new_n15737_));
  INV_X1     g15417(.I(new_n15737_), .ZN(new_n15738_));
  AOI21_X1   g15418(.A1(new_n5980_), .A2(new_n7204_), .B(new_n15674_), .ZN(new_n15739_));
  XOR2_X1    g15419(.A1(new_n15739_), .A2(new_n15738_), .Z(new_n15740_));
  NOR2_X1    g15420(.A1(new_n15740_), .A2(new_n15735_), .ZN(new_n15741_));
  INV_X1     g15421(.I(new_n15739_), .ZN(new_n15742_));
  NOR2_X1    g15422(.A1(new_n15742_), .A2(new_n15738_), .ZN(new_n15743_));
  NOR2_X1    g15423(.A1(new_n15739_), .A2(new_n15737_), .ZN(new_n15744_));
  NOR2_X1    g15424(.A1(new_n15743_), .A2(new_n15744_), .ZN(new_n15745_));
  NOR2_X1    g15425(.A1(new_n15745_), .A2(new_n15734_), .ZN(new_n15746_));
  NOR2_X1    g15426(.A1(new_n15746_), .A2(new_n15741_), .ZN(new_n15747_));
  INV_X1     g15427(.I(new_n15681_), .ZN(new_n15748_));
  AOI21_X1   g15428(.A1(new_n15671_), .A2(new_n15748_), .B(new_n15679_), .ZN(new_n15749_));
  INV_X1     g15429(.I(new_n15749_), .ZN(new_n15750_));
  AOI21_X1   g15430(.A1(new_n5173_), .A2(new_n15677_), .B(new_n8242_), .ZN(new_n15751_));
  AOI21_X1   g15431(.A1(new_n7512_), .A2(new_n9029_), .B(new_n3837_), .ZN(new_n15752_));
  INV_X1     g15432(.I(new_n15752_), .ZN(new_n15753_));
  NOR2_X1    g15433(.A1(new_n15753_), .A2(new_n15751_), .ZN(new_n15754_));
  XOR2_X1    g15434(.A1(new_n15754_), .A2(\a[37] ), .Z(new_n15755_));
  XOR2_X1    g15435(.A1(new_n15755_), .A2(new_n9310_), .Z(new_n15756_));
  NOR2_X1    g15436(.A1(new_n15756_), .A2(new_n15750_), .ZN(new_n15757_));
  INV_X1     g15437(.I(new_n15756_), .ZN(new_n15758_));
  NOR2_X1    g15438(.A1(new_n15758_), .A2(new_n15749_), .ZN(new_n15759_));
  NOR2_X1    g15439(.A1(new_n15759_), .A2(new_n15757_), .ZN(new_n15760_));
  NOR2_X1    g15440(.A1(new_n15760_), .A2(new_n15747_), .ZN(new_n15761_));
  XOR2_X1    g15441(.A1(new_n15756_), .A2(new_n15749_), .Z(new_n15762_));
  NOR3_X1    g15442(.A1(new_n15762_), .A2(new_n15741_), .A3(new_n15746_), .ZN(new_n15763_));
  NOR2_X1    g15443(.A1(new_n15761_), .A2(new_n15763_), .ZN(new_n15764_));
  XOR2_X1    g15444(.A1(new_n15764_), .A2(new_n15733_), .Z(new_n15765_));
  INV_X1     g15445(.I(new_n15733_), .ZN(new_n15766_));
  NOR2_X1    g15446(.A1(new_n15764_), .A2(new_n15766_), .ZN(new_n15767_));
  NOR3_X1    g15447(.A1(new_n15733_), .A2(new_n15761_), .A3(new_n15763_), .ZN(new_n15768_));
  OAI21_X1   g15448(.A1(new_n15767_), .A2(new_n15768_), .B(new_n15715_), .ZN(new_n15769_));
  OAI21_X1   g15449(.A1(new_n15765_), .A2(new_n15715_), .B(new_n15769_), .ZN(new_n15770_));
  OAI21_X1   g15450(.A1(new_n15597_), .A2(new_n15628_), .B(new_n15630_), .ZN(new_n15771_));
  NOR2_X1    g15451(.A1(new_n8992_), .A2(new_n4321_), .ZN(new_n15772_));
  NAND3_X1   g15452(.A1(new_n15772_), .A2(new_n12915_), .A3(new_n15564_), .ZN(new_n15773_));
  AOI21_X1   g15453(.A1(new_n15773_), .A2(new_n9785_), .B(new_n5340_), .ZN(new_n15774_));
  NOR2_X1    g15454(.A1(new_n8992_), .A2(new_n4321_), .ZN(new_n15775_));
  NOR2_X1    g15455(.A1(new_n8243_), .A2(new_n10959_), .ZN(new_n15776_));
  NOR2_X1    g15456(.A1(new_n15776_), .A2(new_n15445_), .ZN(new_n15777_));
  NOR4_X1    g15457(.A1(new_n5742_), .A2(new_n8755_), .A3(new_n4501_), .A4(new_n7727_), .ZN(new_n15778_));
  NAND2_X1   g15458(.A1(new_n15777_), .A2(new_n15778_), .ZN(new_n15779_));
  XNOR2_X1   g15459(.A1(new_n5350_), .A2(new_n8676_), .ZN(new_n15780_));
  NOR2_X1    g15460(.A1(new_n15779_), .A2(new_n15780_), .ZN(new_n15781_));
  INV_X1     g15461(.I(new_n15781_), .ZN(new_n15782_));
  NAND2_X1   g15462(.A1(new_n15779_), .A2(new_n15780_), .ZN(new_n15783_));
  NAND2_X1   g15463(.A1(new_n15782_), .A2(new_n15783_), .ZN(new_n15784_));
  XNOR2_X1   g15464(.A1(new_n15779_), .A2(new_n15780_), .ZN(new_n15785_));
  NOR2_X1    g15465(.A1(new_n15785_), .A2(new_n15775_), .ZN(new_n15786_));
  AOI21_X1   g15466(.A1(new_n15775_), .A2(new_n15784_), .B(new_n15786_), .ZN(new_n15787_));
  INV_X1     g15467(.I(new_n15787_), .ZN(new_n15788_));
  NAND2_X1   g15468(.A1(new_n15647_), .A2(new_n15644_), .ZN(new_n15789_));
  NAND2_X1   g15469(.A1(new_n15789_), .A2(new_n15646_), .ZN(new_n15790_));
  XOR2_X1    g15470(.A1(new_n15790_), .A2(new_n15788_), .Z(new_n15791_));
  NAND2_X1   g15471(.A1(new_n15791_), .A2(new_n15771_), .ZN(new_n15792_));
  AOI21_X1   g15472(.A1(new_n15789_), .A2(new_n15646_), .B(new_n15787_), .ZN(new_n15793_));
  NOR2_X1    g15473(.A1(new_n15790_), .A2(new_n15788_), .ZN(new_n15794_));
  NOR2_X1    g15474(.A1(new_n15794_), .A2(new_n15793_), .ZN(new_n15795_));
  OAI21_X1   g15475(.A1(new_n15771_), .A2(new_n15795_), .B(new_n15792_), .ZN(new_n15796_));
  XNOR2_X1   g15476(.A1(new_n15770_), .A2(new_n15796_), .ZN(new_n15797_));
  INV_X1     g15477(.I(new_n15797_), .ZN(new_n15798_));
  NAND2_X1   g15478(.A1(new_n15770_), .A2(new_n15796_), .ZN(new_n15799_));
  NOR2_X1    g15479(.A1(new_n15770_), .A2(new_n15796_), .ZN(new_n15800_));
  INV_X1     g15480(.I(new_n15800_), .ZN(new_n15801_));
  AOI21_X1   g15481(.A1(new_n15801_), .A2(new_n15799_), .B(new_n15714_), .ZN(new_n15802_));
  AOI21_X1   g15482(.A1(new_n15798_), .A2(new_n15714_), .B(new_n15802_), .ZN(new_n15803_));
  NOR2_X1    g15483(.A1(new_n15713_), .A2(new_n15803_), .ZN(new_n15804_));
  INV_X1     g15484(.I(new_n15804_), .ZN(new_n15805_));
  NAND2_X1   g15485(.A1(new_n15713_), .A2(new_n15803_), .ZN(new_n15806_));
  NAND2_X1   g15486(.A1(new_n15805_), .A2(new_n15806_), .ZN(new_n15807_));
  XOR2_X1    g15487(.A1(new_n15710_), .A2(new_n15807_), .Z(\asquared[101] ));
  NOR2_X1    g15488(.A1(new_n15806_), .A2(new_n15701_), .ZN(new_n15809_));
  NOR2_X1    g15489(.A1(new_n15809_), .A2(new_n15702_), .ZN(new_n15810_));
  AOI21_X1   g15490(.A1(new_n15701_), .A2(new_n15806_), .B(new_n15810_), .ZN(new_n15811_));
  NAND2_X1   g15491(.A1(new_n15592_), .A2(new_n15811_), .ZN(new_n15812_));
  AOI21_X1   g15492(.A1(new_n15714_), .A2(new_n15799_), .B(new_n15800_), .ZN(new_n15813_));
  NOR2_X1    g15493(.A1(new_n15767_), .A2(new_n15715_), .ZN(new_n15814_));
  NOR2_X1    g15494(.A1(new_n15814_), .A2(new_n15768_), .ZN(new_n15815_));
  INV_X1     g15495(.I(new_n15794_), .ZN(new_n15816_));
  AOI21_X1   g15496(.A1(new_n15816_), .A2(new_n15771_), .B(new_n15793_), .ZN(new_n15817_));
  INV_X1     g15497(.I(new_n15757_), .ZN(new_n15818_));
  AOI21_X1   g15498(.A1(new_n15818_), .A2(new_n15747_), .B(new_n15759_), .ZN(new_n15819_));
  INV_X1     g15499(.I(new_n15819_), .ZN(new_n15820_));
  AOI21_X1   g15500(.A1(new_n5742_), .A2(new_n8755_), .B(new_n15777_), .ZN(new_n15821_));
  AOI21_X1   g15501(.A1(new_n5350_), .A2(new_n8933_), .B(new_n8676_), .ZN(new_n15822_));
  XOR2_X1    g15502(.A1(new_n15821_), .A2(new_n15822_), .Z(new_n15823_));
  NOR3_X1    g15503(.A1(new_n15823_), .A2(new_n15772_), .A3(new_n15774_), .ZN(new_n15824_));
  NOR2_X1    g15504(.A1(new_n15774_), .A2(new_n15772_), .ZN(new_n15825_));
  INV_X1     g15505(.I(new_n15821_), .ZN(new_n15826_));
  NOR2_X1    g15506(.A1(new_n15826_), .A2(new_n15822_), .ZN(new_n15827_));
  INV_X1     g15507(.I(new_n15827_), .ZN(new_n15828_));
  NAND2_X1   g15508(.A1(new_n15826_), .A2(new_n15822_), .ZN(new_n15829_));
  AOI21_X1   g15509(.A1(new_n15828_), .A2(new_n15829_), .B(new_n15825_), .ZN(new_n15830_));
  NOR2_X1    g15510(.A1(new_n15830_), .A2(new_n15824_), .ZN(new_n15831_));
  NAND2_X1   g15511(.A1(new_n15783_), .A2(new_n15775_), .ZN(new_n15832_));
  NAND2_X1   g15512(.A1(new_n15832_), .A2(new_n15782_), .ZN(new_n15833_));
  INV_X1     g15513(.I(new_n15833_), .ZN(new_n15834_));
  NOR2_X1    g15514(.A1(new_n15744_), .A2(new_n15735_), .ZN(new_n15835_));
  NOR2_X1    g15515(.A1(new_n15835_), .A2(new_n15743_), .ZN(new_n15836_));
  NOR2_X1    g15516(.A1(new_n15834_), .A2(new_n15836_), .ZN(new_n15837_));
  INV_X1     g15517(.I(new_n15837_), .ZN(new_n15838_));
  NAND2_X1   g15518(.A1(new_n15834_), .A2(new_n15836_), .ZN(new_n15839_));
  AOI21_X1   g15519(.A1(new_n15838_), .A2(new_n15839_), .B(new_n15831_), .ZN(new_n15840_));
  XOR2_X1    g15520(.A1(new_n15836_), .A2(new_n15833_), .Z(new_n15841_));
  NOR3_X1    g15521(.A1(new_n15841_), .A2(new_n15824_), .A3(new_n15830_), .ZN(new_n15842_));
  NOR2_X1    g15522(.A1(new_n15842_), .A2(new_n15840_), .ZN(new_n15843_));
  NOR2_X1    g15523(.A1(new_n15820_), .A2(new_n15843_), .ZN(new_n15844_));
  NOR3_X1    g15524(.A1(new_n15819_), .A2(new_n15840_), .A3(new_n15842_), .ZN(new_n15845_));
  NOR2_X1    g15525(.A1(new_n15844_), .A2(new_n15845_), .ZN(new_n15846_));
  NOR2_X1    g15526(.A1(new_n15846_), .A2(new_n15817_), .ZN(new_n15847_));
  XNOR2_X1   g15527(.A1(new_n15843_), .A2(new_n15819_), .ZN(new_n15848_));
  AOI21_X1   g15528(.A1(new_n15817_), .A2(new_n15848_), .B(new_n15847_), .ZN(new_n15849_));
  AOI21_X1   g15529(.A1(new_n15723_), .A2(new_n15730_), .B(new_n15729_), .ZN(new_n15850_));
  NOR2_X1    g15530(.A1(new_n7187_), .A2(new_n8244_), .ZN(new_n15851_));
  NOR2_X1    g15531(.A1(new_n4769_), .A2(new_n5004_), .ZN(new_n15852_));
  INV_X1     g15532(.I(new_n15852_), .ZN(new_n15853_));
  NOR2_X1    g15533(.A1(new_n7187_), .A2(new_n8244_), .ZN(new_n15857_));
  NOR2_X1    g15534(.A1(new_n8565_), .A2(new_n11805_), .ZN(new_n15859_));
  NOR4_X1    g15535(.A1(new_n4770_), .A2(new_n5745_), .A3(new_n6692_), .A4(new_n7727_), .ZN(new_n15863_));
  INV_X1     g15536(.I(new_n15863_), .ZN(new_n15864_));
  NAND2_X1   g15537(.A1(new_n7483_), .A2(new_n5980_), .ZN(new_n15865_));
  NAND2_X1   g15538(.A1(\a[38] ), .A2(\a[63] ), .ZN(new_n15866_));
  XNOR2_X1   g15539(.A1(new_n15865_), .A2(new_n15866_), .ZN(new_n15867_));
  NOR2_X1    g15540(.A1(new_n15867_), .A2(new_n15864_), .ZN(new_n15868_));
  INV_X1     g15541(.I(new_n15868_), .ZN(new_n15869_));
  NAND2_X1   g15542(.A1(new_n15867_), .A2(new_n15864_), .ZN(new_n15870_));
  NAND2_X1   g15543(.A1(new_n15869_), .A2(new_n15870_), .ZN(new_n15871_));
  XOR2_X1    g15544(.A1(new_n15867_), .A2(new_n15863_), .Z(new_n15872_));
  NOR2_X1    g15545(.A1(new_n15872_), .A2(new_n15857_), .ZN(new_n15873_));
  AOI21_X1   g15546(.A1(new_n15857_), .A2(new_n15871_), .B(new_n15873_), .ZN(new_n15874_));
  NAND2_X1   g15547(.A1(\a[41] ), .A2(\a[61] ), .ZN(new_n15875_));
  XNOR2_X1   g15548(.A1(new_n15328_), .A2(new_n15875_), .ZN(new_n15876_));
  INV_X1     g15549(.I(new_n15876_), .ZN(new_n15877_));
  NAND2_X1   g15550(.A1(new_n15718_), .A2(new_n15877_), .ZN(new_n15878_));
  NOR2_X1    g15551(.A1(new_n15718_), .A2(new_n15877_), .ZN(new_n15879_));
  INV_X1     g15552(.I(new_n15879_), .ZN(new_n15880_));
  AND2_X2    g15553(.A1(new_n15880_), .A2(new_n15878_), .Z(new_n15881_));
  NAND2_X1   g15554(.A1(new_n15753_), .A2(new_n15751_), .ZN(new_n15882_));
  NOR2_X1    g15555(.A1(new_n3837_), .A2(new_n9310_), .ZN(new_n15883_));
  AOI21_X1   g15556(.A1(new_n15882_), .A2(new_n15883_), .B(new_n15754_), .ZN(new_n15884_));
  NAND2_X1   g15557(.A1(\a[50] ), .A2(\a[62] ), .ZN(new_n15885_));
  XOR2_X1    g15558(.A1(new_n7461_), .A2(new_n15885_), .Z(new_n15886_));
  NOR2_X1    g15559(.A1(new_n15884_), .A2(new_n15886_), .ZN(new_n15887_));
  INV_X1     g15560(.I(new_n15887_), .ZN(new_n15888_));
  NAND2_X1   g15561(.A1(new_n15884_), .A2(new_n15886_), .ZN(new_n15889_));
  AOI21_X1   g15562(.A1(new_n15888_), .A2(new_n15889_), .B(new_n15881_), .ZN(new_n15890_));
  INV_X1     g15563(.I(new_n15881_), .ZN(new_n15891_));
  XNOR2_X1   g15564(.A1(new_n15884_), .A2(new_n15886_), .ZN(new_n15892_));
  NOR2_X1    g15565(.A1(new_n15891_), .A2(new_n15892_), .ZN(new_n15893_));
  NOR2_X1    g15566(.A1(new_n15893_), .A2(new_n15890_), .ZN(new_n15894_));
  XNOR2_X1   g15567(.A1(new_n15894_), .A2(new_n15874_), .ZN(new_n15895_));
  NOR2_X1    g15568(.A1(new_n15894_), .A2(new_n15874_), .ZN(new_n15896_));
  INV_X1     g15569(.I(new_n15896_), .ZN(new_n15897_));
  NAND2_X1   g15570(.A1(new_n15894_), .A2(new_n15874_), .ZN(new_n15898_));
  NAND2_X1   g15571(.A1(new_n15897_), .A2(new_n15898_), .ZN(new_n15899_));
  NAND2_X1   g15572(.A1(new_n15899_), .A2(new_n15850_), .ZN(new_n15900_));
  OAI21_X1   g15573(.A1(new_n15850_), .A2(new_n15895_), .B(new_n15900_), .ZN(new_n15901_));
  NAND2_X1   g15574(.A1(new_n15849_), .A2(new_n15901_), .ZN(new_n15902_));
  NOR2_X1    g15575(.A1(new_n15849_), .A2(new_n15901_), .ZN(new_n15903_));
  INV_X1     g15576(.I(new_n15903_), .ZN(new_n15904_));
  AOI21_X1   g15577(.A1(new_n15904_), .A2(new_n15902_), .B(new_n15815_), .ZN(new_n15905_));
  XOR2_X1    g15578(.A1(new_n15849_), .A2(new_n15901_), .Z(new_n15906_));
  AOI21_X1   g15579(.A1(new_n15815_), .A2(new_n15906_), .B(new_n15905_), .ZN(new_n15907_));
  NOR2_X1    g15580(.A1(new_n15907_), .A2(new_n15813_), .ZN(new_n15908_));
  XOR2_X1    g15581(.A1(new_n15812_), .A2(new_n15908_), .Z(new_n15909_));
  XOR2_X1    g15582(.A1(new_n15909_), .A2(new_n15805_), .Z(\asquared[102] ));
  NOR2_X1    g15583(.A1(new_n15805_), .A2(new_n15813_), .ZN(new_n15911_));
  INV_X1     g15584(.I(new_n15911_), .ZN(new_n15912_));
  AOI21_X1   g15585(.A1(new_n15805_), .A2(new_n15813_), .B(new_n15907_), .ZN(new_n15913_));
  NAND3_X1   g15586(.A1(new_n15592_), .A2(new_n15811_), .A3(new_n15913_), .ZN(new_n15914_));
  AND2_X2    g15587(.A1(new_n15914_), .A2(new_n15912_), .Z(new_n15915_));
  OAI21_X1   g15588(.A1(new_n15768_), .A2(new_n15814_), .B(new_n15902_), .ZN(new_n15916_));
  NAND2_X1   g15589(.A1(new_n15916_), .A2(new_n15904_), .ZN(new_n15917_));
  INV_X1     g15590(.I(new_n15845_), .ZN(new_n15918_));
  OAI21_X1   g15591(.A1(new_n15817_), .A2(new_n15844_), .B(new_n15918_), .ZN(new_n15919_));
  INV_X1     g15592(.I(new_n15898_), .ZN(new_n15920_));
  OAI21_X1   g15593(.A1(new_n15850_), .A2(new_n15920_), .B(new_n15897_), .ZN(new_n15921_));
  INV_X1     g15594(.I(new_n15921_), .ZN(new_n15922_));
  AOI21_X1   g15595(.A1(new_n6028_), .A2(new_n7204_), .B(new_n15859_), .ZN(new_n15923_));
  NOR2_X1    g15596(.A1(new_n7483_), .A2(new_n5980_), .ZN(new_n15924_));
  NAND2_X1   g15597(.A1(new_n3804_), .A2(new_n9310_), .ZN(new_n15925_));
  AOI21_X1   g15598(.A1(new_n5980_), .A2(new_n7483_), .B(new_n15925_), .ZN(new_n15926_));
  NOR2_X1    g15599(.A1(new_n15926_), .A2(new_n15924_), .ZN(new_n15927_));
  AOI21_X1   g15600(.A1(\a[62] ), .A2(new_n7461_), .B(new_n6779_), .ZN(new_n15928_));
  XOR2_X1    g15601(.A1(new_n15927_), .A2(new_n15928_), .Z(new_n15929_));
  NAND2_X1   g15602(.A1(new_n15929_), .A2(new_n15923_), .ZN(new_n15930_));
  INV_X1     g15603(.I(new_n15923_), .ZN(new_n15931_));
  AND2_X2    g15604(.A1(new_n15927_), .A2(new_n15928_), .Z(new_n15932_));
  NOR2_X1    g15605(.A1(new_n15927_), .A2(new_n15928_), .ZN(new_n15933_));
  OAI21_X1   g15606(.A1(new_n15932_), .A2(new_n15933_), .B(new_n15931_), .ZN(new_n15934_));
  NAND2_X1   g15607(.A1(new_n15930_), .A2(new_n15934_), .ZN(new_n15935_));
  INV_X1     g15608(.I(new_n15935_), .ZN(new_n15936_));
  NAND2_X1   g15609(.A1(new_n15829_), .A2(new_n15825_), .ZN(new_n15937_));
  NAND2_X1   g15610(.A1(new_n15937_), .A2(new_n15828_), .ZN(new_n15938_));
  INV_X1     g15611(.I(new_n15938_), .ZN(new_n15939_));
  NAND2_X1   g15612(.A1(new_n15870_), .A2(new_n15857_), .ZN(new_n15940_));
  NAND2_X1   g15613(.A1(new_n15940_), .A2(new_n15869_), .ZN(new_n15941_));
  INV_X1     g15614(.I(new_n15941_), .ZN(new_n15942_));
  NOR2_X1    g15615(.A1(new_n15939_), .A2(new_n15942_), .ZN(new_n15943_));
  NOR2_X1    g15616(.A1(new_n15938_), .A2(new_n15941_), .ZN(new_n15944_));
  NOR2_X1    g15617(.A1(new_n15943_), .A2(new_n15944_), .ZN(new_n15945_));
  NOR2_X1    g15618(.A1(new_n15945_), .A2(new_n15936_), .ZN(new_n15946_));
  XOR2_X1    g15619(.A1(new_n15938_), .A2(new_n15942_), .Z(new_n15947_));
  NOR2_X1    g15620(.A1(new_n15947_), .A2(new_n15935_), .ZN(new_n15948_));
  NOR2_X1    g15621(.A1(new_n15946_), .A2(new_n15948_), .ZN(new_n15949_));
  AOI21_X1   g15622(.A1(new_n15831_), .A2(new_n15839_), .B(new_n15837_), .ZN(new_n15950_));
  XOR2_X1    g15623(.A1(new_n15949_), .A2(new_n15950_), .Z(new_n15951_));
  NOR2_X1    g15624(.A1(new_n15951_), .A2(new_n15922_), .ZN(new_n15952_));
  INV_X1     g15625(.I(new_n15949_), .ZN(new_n15953_));
  NOR2_X1    g15626(.A1(new_n15953_), .A2(new_n15950_), .ZN(new_n15954_));
  INV_X1     g15627(.I(new_n15954_), .ZN(new_n15955_));
  NAND2_X1   g15628(.A1(new_n15953_), .A2(new_n15950_), .ZN(new_n15956_));
  AOI21_X1   g15629(.A1(new_n15955_), .A2(new_n15956_), .B(new_n15921_), .ZN(new_n15957_));
  NOR2_X1    g15630(.A1(new_n15957_), .A2(new_n15952_), .ZN(new_n15958_));
  OAI22_X1   g15631(.A1(new_n13260_), .A2(new_n12355_), .B1(new_n10288_), .B2(new_n10290_), .ZN(new_n15959_));
  OAI21_X1   g15632(.A1(new_n7512_), .A2(new_n8056_), .B(new_n15959_), .ZN(new_n15960_));
  INV_X1     g15633(.I(new_n15960_), .ZN(new_n15961_));
  AOI21_X1   g15634(.A1(new_n15961_), .A2(new_n6776_), .B(\a[53] ), .ZN(new_n15962_));
  NOR2_X1    g15635(.A1(\a[48] ), .A2(\a[54] ), .ZN(new_n15963_));
  OAI21_X1   g15636(.A1(new_n15962_), .A2(new_n5745_), .B(new_n15963_), .ZN(new_n15964_));
  AOI21_X1   g15637(.A1(new_n6280_), .A2(new_n7204_), .B(new_n15959_), .ZN(new_n15965_));
  NAND2_X1   g15638(.A1(new_n15964_), .A2(new_n15965_), .ZN(new_n15966_));
  NOR2_X1    g15639(.A1(new_n15776_), .A2(new_n15673_), .ZN(new_n15967_));
  NOR4_X1    g15640(.A1(new_n8755_), .A2(new_n5980_), .A3(new_n5004_), .A4(new_n7727_), .ZN(new_n15968_));
  NAND2_X1   g15641(.A1(new_n15967_), .A2(new_n15968_), .ZN(new_n15969_));
  XNOR2_X1   g15642(.A1(new_n5321_), .A2(new_n8676_), .ZN(new_n15970_));
  NOR2_X1    g15643(.A1(new_n15969_), .A2(new_n15970_), .ZN(new_n15971_));
  INV_X1     g15644(.I(new_n15969_), .ZN(new_n15972_));
  INV_X1     g15645(.I(new_n15970_), .ZN(new_n15973_));
  NOR2_X1    g15646(.A1(new_n15972_), .A2(new_n15973_), .ZN(new_n15974_));
  NOR2_X1    g15647(.A1(new_n15974_), .A2(new_n15971_), .ZN(new_n15975_));
  NOR2_X1    g15648(.A1(new_n15966_), .A2(new_n15975_), .ZN(new_n15976_));
  XOR2_X1    g15649(.A1(new_n15969_), .A2(new_n15970_), .Z(new_n15977_));
  AOI21_X1   g15650(.A1(new_n15966_), .A2(new_n15977_), .B(new_n15976_), .ZN(new_n15978_));
  INV_X1     g15651(.I(new_n15978_), .ZN(new_n15979_));
  NOR2_X1    g15652(.A1(new_n6579_), .A2(new_n8992_), .ZN(new_n15980_));
  AOI21_X1   g15653(.A1(new_n5173_), .A2(new_n8676_), .B(new_n15851_), .ZN(new_n15981_));
  NOR2_X1    g15654(.A1(new_n5881_), .A2(new_n8992_), .ZN(new_n15982_));
  NOR2_X1    g15655(.A1(new_n5881_), .A2(new_n8992_), .ZN(new_n15986_));
  NAND2_X1   g15656(.A1(new_n15981_), .A2(new_n15986_), .ZN(new_n15987_));
  XOR2_X1    g15657(.A1(new_n15879_), .A2(new_n15987_), .Z(new_n15988_));
  XOR2_X1    g15658(.A1(new_n15988_), .A2(new_n15980_), .Z(new_n15989_));
  AOI21_X1   g15659(.A1(new_n15891_), .A2(new_n15889_), .B(new_n15887_), .ZN(new_n15990_));
  XNOR2_X1   g15660(.A1(new_n15989_), .A2(new_n15990_), .ZN(new_n15991_));
  INV_X1     g15661(.I(new_n15991_), .ZN(new_n15992_));
  NOR2_X1    g15662(.A1(new_n15989_), .A2(new_n15990_), .ZN(new_n15993_));
  NAND2_X1   g15663(.A1(new_n15989_), .A2(new_n15990_), .ZN(new_n15994_));
  INV_X1     g15664(.I(new_n15994_), .ZN(new_n15995_));
  NOR2_X1    g15665(.A1(new_n15995_), .A2(new_n15993_), .ZN(new_n15996_));
  NOR2_X1    g15666(.A1(new_n15996_), .A2(new_n15979_), .ZN(new_n15997_));
  AOI21_X1   g15667(.A1(new_n15979_), .A2(new_n15992_), .B(new_n15997_), .ZN(new_n15998_));
  NOR2_X1    g15668(.A1(new_n15958_), .A2(new_n15998_), .ZN(new_n15999_));
  INV_X1     g15669(.I(new_n15958_), .ZN(new_n16000_));
  INV_X1     g15670(.I(new_n15998_), .ZN(new_n16001_));
  NOR2_X1    g15671(.A1(new_n16000_), .A2(new_n16001_), .ZN(new_n16002_));
  NOR2_X1    g15672(.A1(new_n16002_), .A2(new_n15999_), .ZN(new_n16003_));
  XOR2_X1    g15673(.A1(new_n15958_), .A2(new_n16001_), .Z(new_n16004_));
  MUX2_X1    g15674(.I0(new_n16004_), .I1(new_n16003_), .S(new_n15919_), .Z(new_n16005_));
  INV_X1     g15675(.I(new_n16005_), .ZN(new_n16006_));
  NAND2_X1   g15676(.A1(new_n16006_), .A2(new_n15917_), .ZN(new_n16007_));
  INV_X1     g15677(.I(new_n16007_), .ZN(new_n16008_));
  NOR2_X1    g15678(.A1(new_n16006_), .A2(new_n15917_), .ZN(new_n16009_));
  NOR2_X1    g15679(.A1(new_n16008_), .A2(new_n16009_), .ZN(new_n16010_));
  XOR2_X1    g15680(.A1(new_n15915_), .A2(new_n16010_), .Z(\asquared[103] ));
  AOI21_X1   g15681(.A1(new_n15915_), .A2(new_n16007_), .B(new_n16009_), .ZN(new_n16012_));
  INV_X1     g15682(.I(new_n15999_), .ZN(new_n16013_));
  AOI21_X1   g15683(.A1(new_n15919_), .A2(new_n16013_), .B(new_n16002_), .ZN(new_n16014_));
  AOI21_X1   g15684(.A1(new_n15921_), .A2(new_n15956_), .B(new_n15954_), .ZN(new_n16015_));
  INV_X1     g15685(.I(new_n15971_), .ZN(new_n16016_));
  OAI21_X1   g15686(.A1(new_n15966_), .A2(new_n15974_), .B(new_n16016_), .ZN(new_n16017_));
  INV_X1     g15687(.I(new_n16017_), .ZN(new_n16018_));
  NOR2_X1    g15688(.A1(new_n15879_), .A2(new_n15981_), .ZN(new_n16019_));
  NOR3_X1    g15689(.A1(new_n16019_), .A2(new_n6579_), .A3(new_n8992_), .ZN(new_n16020_));
  AOI22_X1   g15690(.A1(new_n16020_), .A2(new_n15986_), .B1(new_n15879_), .B2(new_n15981_), .ZN(new_n16021_));
  NOR2_X1    g15691(.A1(new_n15931_), .A2(new_n15933_), .ZN(new_n16022_));
  NOR2_X1    g15692(.A1(new_n16022_), .A2(new_n15932_), .ZN(new_n16023_));
  XNOR2_X1   g15693(.A1(new_n16021_), .A2(new_n16023_), .ZN(new_n16024_));
  NOR2_X1    g15694(.A1(new_n16021_), .A2(new_n16023_), .ZN(new_n16025_));
  NAND2_X1   g15695(.A1(new_n16021_), .A2(new_n16023_), .ZN(new_n16026_));
  INV_X1     g15696(.I(new_n16026_), .ZN(new_n16027_));
  OAI21_X1   g15697(.A1(new_n16027_), .A2(new_n16025_), .B(new_n16018_), .ZN(new_n16028_));
  OAI21_X1   g15698(.A1(new_n16018_), .A2(new_n16024_), .B(new_n16028_), .ZN(new_n16029_));
  INV_X1     g15699(.I(new_n16029_), .ZN(new_n16030_));
  AOI21_X1   g15700(.A1(new_n15979_), .A2(new_n15994_), .B(new_n15993_), .ZN(new_n16031_));
  NOR2_X1    g15701(.A1(new_n15944_), .A2(new_n15935_), .ZN(new_n16032_));
  NOR2_X1    g15702(.A1(new_n16032_), .A2(new_n15943_), .ZN(new_n16033_));
  NOR2_X1    g15703(.A1(new_n16031_), .A2(new_n16033_), .ZN(new_n16034_));
  INV_X1     g15704(.I(new_n16034_), .ZN(new_n16035_));
  NAND2_X1   g15705(.A1(new_n16031_), .A2(new_n16033_), .ZN(new_n16036_));
  AOI21_X1   g15706(.A1(new_n16035_), .A2(new_n16036_), .B(new_n16030_), .ZN(new_n16037_));
  XNOR2_X1   g15707(.A1(new_n16031_), .A2(new_n16033_), .ZN(new_n16038_));
  NOR2_X1    g15708(.A1(new_n16038_), .A2(new_n16029_), .ZN(new_n16039_));
  NOR2_X1    g15709(.A1(new_n16039_), .A2(new_n16037_), .ZN(new_n16040_));
  INV_X1     g15710(.I(new_n16040_), .ZN(new_n16041_));
  NOR4_X1    g15711(.A1(new_n15853_), .A2(new_n7647_), .A3(new_n8085_), .A4(new_n8453_), .ZN(new_n16042_));
  NOR3_X1    g15712(.A1(new_n7023_), .A2(new_n5743_), .A3(new_n8989_), .ZN(new_n16043_));
  NOR2_X1    g15713(.A1(new_n16043_), .A2(new_n16042_), .ZN(new_n16044_));
  INV_X1     g15714(.I(new_n16044_), .ZN(new_n16045_));
  NOR3_X1    g15715(.A1(new_n16045_), .A2(new_n4769_), .A3(new_n8453_), .ZN(new_n16046_));
  NOR3_X1    g15716(.A1(new_n16045_), .A2(new_n5742_), .A3(new_n8676_), .ZN(new_n16047_));
  NOR2_X1    g15717(.A1(new_n16047_), .A2(new_n16046_), .ZN(new_n16048_));
  AOI21_X1   g15718(.A1(new_n4415_), .A2(new_n9781_), .B(new_n15982_), .ZN(new_n16049_));
  AOI21_X1   g15719(.A1(new_n5321_), .A2(new_n12915_), .B(new_n8676_), .ZN(new_n16050_));
  INV_X1     g15720(.I(new_n16050_), .ZN(new_n16051_));
  AND2_X2    g15721(.A1(new_n16049_), .A2(new_n16051_), .Z(new_n16052_));
  NOR2_X1    g15722(.A1(new_n16049_), .A2(new_n16051_), .ZN(new_n16053_));
  OAI21_X1   g15723(.A1(new_n16052_), .A2(new_n16053_), .B(new_n16048_), .ZN(new_n16054_));
  XOR2_X1    g15724(.A1(new_n16049_), .A2(new_n16050_), .Z(new_n16055_));
  OAI21_X1   g15725(.A1(new_n16048_), .A2(new_n16055_), .B(new_n16054_), .ZN(new_n16056_));
  NAND2_X1   g15726(.A1(new_n8242_), .A2(new_n5980_), .ZN(new_n16057_));
  NAND2_X1   g15727(.A1(\a[43] ), .A2(\a[60] ), .ZN(new_n16058_));
  XNOR2_X1   g15728(.A1(new_n16057_), .A2(new_n16058_), .ZN(new_n16059_));
  AOI22_X1   g15729(.A1(new_n6056_), .A2(new_n7483_), .B1(new_n6028_), .B2(new_n7485_), .ZN(new_n16060_));
  NAND4_X1   g15730(.A1(new_n16060_), .A2(new_n7512_), .A3(new_n10288_), .A4(new_n14857_), .ZN(new_n16061_));
  NOR2_X1    g15731(.A1(new_n6692_), .A2(\a[51] ), .ZN(new_n16062_));
  XOR2_X1    g15732(.A1(new_n13186_), .A2(new_n16062_), .Z(new_n16063_));
  NOR2_X1    g15733(.A1(new_n16061_), .A2(new_n16063_), .ZN(new_n16064_));
  INV_X1     g15734(.I(new_n16064_), .ZN(new_n16065_));
  NAND2_X1   g15735(.A1(new_n16061_), .A2(new_n16063_), .ZN(new_n16066_));
  AOI21_X1   g15736(.A1(new_n16065_), .A2(new_n16066_), .B(new_n16059_), .ZN(new_n16067_));
  INV_X1     g15737(.I(new_n16059_), .ZN(new_n16068_));
  XNOR2_X1   g15738(.A1(new_n16061_), .A2(new_n16063_), .ZN(new_n16069_));
  NOR2_X1    g15739(.A1(new_n16069_), .A2(new_n16068_), .ZN(new_n16070_));
  NOR2_X1    g15740(.A1(new_n16070_), .A2(new_n16067_), .ZN(new_n16071_));
  AOI21_X1   g15741(.A1(new_n5980_), .A2(new_n8755_), .B(new_n15967_), .ZN(new_n16072_));
  INV_X1     g15742(.I(new_n16072_), .ZN(new_n16073_));
  NOR2_X1    g15743(.A1(new_n16073_), .A2(new_n15960_), .ZN(new_n16074_));
  XOR2_X1    g15744(.A1(new_n16074_), .A2(new_n4240_), .Z(new_n16075_));
  XOR2_X1    g15745(.A1(new_n16075_), .A2(\a[63] ), .Z(new_n16076_));
  INV_X1     g15746(.I(new_n16076_), .ZN(new_n16077_));
  NAND2_X1   g15747(.A1(new_n16077_), .A2(new_n16071_), .ZN(new_n16078_));
  NOR2_X1    g15748(.A1(new_n16077_), .A2(new_n16071_), .ZN(new_n16079_));
  INV_X1     g15749(.I(new_n16079_), .ZN(new_n16080_));
  NAND2_X1   g15750(.A1(new_n16080_), .A2(new_n16078_), .ZN(new_n16081_));
  XOR2_X1    g15751(.A1(new_n16076_), .A2(new_n16071_), .Z(new_n16082_));
  NOR2_X1    g15752(.A1(new_n16082_), .A2(new_n16056_), .ZN(new_n16083_));
  AOI21_X1   g15753(.A1(new_n16056_), .A2(new_n16081_), .B(new_n16083_), .ZN(new_n16084_));
  NOR2_X1    g15754(.A1(new_n16041_), .A2(new_n16084_), .ZN(new_n16085_));
  INV_X1     g15755(.I(new_n16084_), .ZN(new_n16086_));
  NOR2_X1    g15756(.A1(new_n16040_), .A2(new_n16086_), .ZN(new_n16087_));
  NOR2_X1    g15757(.A1(new_n16085_), .A2(new_n16087_), .ZN(new_n16088_));
  NOR2_X1    g15758(.A1(new_n16088_), .A2(new_n16015_), .ZN(new_n16089_));
  INV_X1     g15759(.I(new_n16015_), .ZN(new_n16090_));
  XOR2_X1    g15760(.A1(new_n16040_), .A2(new_n16084_), .Z(new_n16091_));
  NOR2_X1    g15761(.A1(new_n16091_), .A2(new_n16090_), .ZN(new_n16092_));
  NOR2_X1    g15762(.A1(new_n16089_), .A2(new_n16092_), .ZN(new_n16093_));
  XOR2_X1    g15763(.A1(new_n16093_), .A2(new_n16014_), .Z(new_n16094_));
  NAND2_X1   g15764(.A1(new_n16012_), .A2(new_n16094_), .ZN(new_n16095_));
  NOR2_X1    g15765(.A1(new_n16093_), .A2(new_n16014_), .ZN(new_n16096_));
  NAND2_X1   g15766(.A1(new_n16093_), .A2(new_n16014_), .ZN(new_n16097_));
  INV_X1     g15767(.I(new_n16097_), .ZN(new_n16098_));
  NOR2_X1    g15768(.A1(new_n16098_), .A2(new_n16096_), .ZN(new_n16099_));
  OAI21_X1   g15769(.A1(new_n16012_), .A2(new_n16099_), .B(new_n16095_), .ZN(\asquared[104] ));
  NAND2_X1   g15770(.A1(new_n16009_), .A2(new_n16096_), .ZN(new_n16101_));
  NAND3_X1   g15771(.A1(new_n15914_), .A2(new_n15912_), .A3(new_n16101_), .ZN(new_n16102_));
  NAND2_X1   g15772(.A1(new_n16102_), .A2(new_n16008_), .ZN(new_n16103_));
  INV_X1     g15773(.I(new_n16087_), .ZN(new_n16104_));
  AOI21_X1   g15774(.A1(new_n16090_), .A2(new_n16104_), .B(new_n16085_), .ZN(new_n16105_));
  AOI21_X1   g15775(.A1(new_n16030_), .A2(new_n16036_), .B(new_n16034_), .ZN(new_n16106_));
  INV_X1     g15776(.I(new_n16106_), .ZN(new_n16107_));
  AOI21_X1   g15777(.A1(new_n16056_), .A2(new_n16078_), .B(new_n16079_), .ZN(new_n16108_));
  AOI21_X1   g15778(.A1(new_n16017_), .A2(new_n16026_), .B(new_n16025_), .ZN(new_n16109_));
  NOR2_X1    g15779(.A1(new_n4769_), .A2(new_n9310_), .ZN(new_n16110_));
  XNOR2_X1   g15780(.A1(new_n13186_), .A2(new_n16110_), .ZN(new_n16111_));
  NAND2_X1   g15781(.A1(\a[40] ), .A2(\a[63] ), .ZN(new_n16112_));
  AOI21_X1   g15782(.A1(new_n16073_), .A2(new_n15960_), .B(new_n16112_), .ZN(new_n16113_));
  NOR2_X1    g15783(.A1(new_n16113_), .A2(new_n16074_), .ZN(new_n16114_));
  INV_X1     g15784(.I(new_n16053_), .ZN(new_n16115_));
  AOI21_X1   g15785(.A1(new_n16048_), .A2(new_n16115_), .B(new_n16052_), .ZN(new_n16116_));
  OAI21_X1   g15786(.A1(new_n13186_), .A2(\a[51] ), .B(\a[52] ), .ZN(new_n16117_));
  XOR2_X1    g15787(.A1(new_n16116_), .A2(new_n16117_), .Z(new_n16118_));
  XNOR2_X1   g15788(.A1(new_n16118_), .A2(new_n16114_), .ZN(new_n16119_));
  XNOR2_X1   g15789(.A1(new_n16119_), .A2(new_n16111_), .ZN(new_n16120_));
  XOR2_X1    g15790(.A1(new_n16120_), .A2(new_n16109_), .Z(new_n16121_));
  INV_X1     g15791(.I(new_n16109_), .ZN(new_n16122_));
  NOR2_X1    g15792(.A1(new_n16120_), .A2(new_n16122_), .ZN(new_n16123_));
  NAND2_X1   g15793(.A1(new_n16120_), .A2(new_n16122_), .ZN(new_n16124_));
  INV_X1     g15794(.I(new_n16124_), .ZN(new_n16125_));
  OAI21_X1   g15795(.A1(new_n16125_), .A2(new_n16123_), .B(new_n16108_), .ZN(new_n16126_));
  OAI21_X1   g15796(.A1(new_n16108_), .A2(new_n16121_), .B(new_n16126_), .ZN(new_n16127_));
  AOI21_X1   g15797(.A1(new_n5742_), .A2(new_n8676_), .B(new_n16045_), .ZN(new_n16128_));
  NAND2_X1   g15798(.A1(new_n8242_), .A2(new_n5980_), .ZN(new_n16129_));
  NOR2_X1    g15799(.A1(new_n8242_), .A2(new_n5980_), .ZN(new_n16130_));
  NOR2_X1    g15800(.A1(\a[43] ), .A2(\a[60] ), .ZN(new_n16131_));
  AOI21_X1   g15801(.A1(new_n16129_), .A2(new_n16131_), .B(new_n16130_), .ZN(new_n16132_));
  AOI21_X1   g15802(.A1(new_n6280_), .A2(new_n7482_), .B(new_n16060_), .ZN(new_n16133_));
  XNOR2_X1   g15803(.A1(new_n16133_), .A2(new_n16132_), .ZN(new_n16134_));
  INV_X1     g15804(.I(new_n16134_), .ZN(new_n16135_));
  AND2_X2    g15805(.A1(new_n16133_), .A2(new_n16132_), .Z(new_n16136_));
  INV_X1     g15806(.I(new_n16136_), .ZN(new_n16137_));
  NOR2_X1    g15807(.A1(new_n16133_), .A2(new_n16132_), .ZN(new_n16138_));
  INV_X1     g15808(.I(new_n16138_), .ZN(new_n16139_));
  AOI21_X1   g15809(.A1(new_n16137_), .A2(new_n16139_), .B(new_n16128_), .ZN(new_n16140_));
  AOI21_X1   g15810(.A1(new_n16135_), .A2(new_n16128_), .B(new_n16140_), .ZN(new_n16141_));
  AOI21_X1   g15811(.A1(new_n16068_), .A2(new_n16066_), .B(new_n16064_), .ZN(new_n16142_));
  AOI22_X1   g15812(.A1(new_n5321_), .A2(new_n5742_), .B1(new_n8991_), .B2(new_n8996_), .ZN(new_n16143_));
  NOR2_X1    g15813(.A1(new_n4770_), .A2(new_n8990_), .ZN(new_n16144_));
  NAND4_X1   g15814(.A1(new_n16143_), .A2(new_n7187_), .A3(new_n8989_), .A4(new_n16144_), .ZN(new_n16145_));
  AOI22_X1   g15815(.A1(new_n7648_), .A2(new_n8198_), .B1(new_n8245_), .B2(new_n5980_), .ZN(new_n16146_));
  INV_X1     g15816(.I(new_n16146_), .ZN(new_n16147_));
  NOR4_X1    g15817(.A1(new_n6030_), .A2(new_n8242_), .A3(new_n5175_), .A4(new_n7647_), .ZN(new_n16148_));
  NAND2_X1   g15818(.A1(new_n16147_), .A2(new_n16148_), .ZN(new_n16149_));
  AOI22_X1   g15819(.A1(new_n6280_), .A2(new_n9299_), .B1(new_n7000_), .B2(new_n7483_), .ZN(new_n16150_));
  NOR2_X1    g15820(.A1(new_n8941_), .A2(new_n10288_), .ZN(new_n16151_));
  AOI21_X1   g15821(.A1(\a[50] ), .A2(\a[54] ), .B(new_n7000_), .ZN(new_n16152_));
  NOR4_X1    g15822(.A1(new_n16151_), .A2(new_n5745_), .A3(new_n6999_), .A4(new_n16152_), .ZN(new_n16153_));
  NAND2_X1   g15823(.A1(new_n16153_), .A2(new_n16150_), .ZN(new_n16154_));
  NOR2_X1    g15824(.A1(new_n16154_), .A2(new_n16149_), .ZN(new_n16155_));
  INV_X1     g15825(.I(new_n16155_), .ZN(new_n16156_));
  NAND2_X1   g15826(.A1(new_n16154_), .A2(new_n16149_), .ZN(new_n16157_));
  AOI21_X1   g15827(.A1(new_n16156_), .A2(new_n16157_), .B(new_n16145_), .ZN(new_n16158_));
  XOR2_X1    g15828(.A1(new_n16154_), .A2(new_n16149_), .Z(new_n16159_));
  AOI21_X1   g15829(.A1(new_n16145_), .A2(new_n16159_), .B(new_n16158_), .ZN(new_n16160_));
  NOR2_X1    g15830(.A1(new_n16160_), .A2(new_n16142_), .ZN(new_n16161_));
  NAND2_X1   g15831(.A1(new_n16160_), .A2(new_n16142_), .ZN(new_n16162_));
  INV_X1     g15832(.I(new_n16162_), .ZN(new_n16163_));
  NOR2_X1    g15833(.A1(new_n16163_), .A2(new_n16161_), .ZN(new_n16164_));
  XOR2_X1    g15834(.A1(new_n16160_), .A2(new_n16142_), .Z(new_n16165_));
  NAND2_X1   g15835(.A1(new_n16165_), .A2(new_n16141_), .ZN(new_n16166_));
  OAI21_X1   g15836(.A1(new_n16141_), .A2(new_n16164_), .B(new_n16166_), .ZN(new_n16167_));
  NAND2_X1   g15837(.A1(new_n16127_), .A2(new_n16167_), .ZN(new_n16168_));
  INV_X1     g15838(.I(new_n16168_), .ZN(new_n16169_));
  NOR2_X1    g15839(.A1(new_n16127_), .A2(new_n16167_), .ZN(new_n16170_));
  OAI21_X1   g15840(.A1(new_n16169_), .A2(new_n16170_), .B(new_n16107_), .ZN(new_n16171_));
  XOR2_X1    g15841(.A1(new_n16127_), .A2(new_n16167_), .Z(new_n16172_));
  NAND2_X1   g15842(.A1(new_n16172_), .A2(new_n16106_), .ZN(new_n16173_));
  AOI21_X1   g15843(.A1(new_n16173_), .A2(new_n16171_), .B(new_n16105_), .ZN(new_n16174_));
  XOR2_X1    g15844(.A1(new_n16103_), .A2(new_n16174_), .Z(new_n16175_));
  XOR2_X1    g15845(.A1(new_n16175_), .A2(new_n16097_), .Z(\asquared[105] ));
  OR2_X2     g15846(.A1(new_n16097_), .A2(new_n16105_), .Z(new_n16177_));
  AOI22_X1   g15847(.A1(new_n16097_), .A2(new_n16105_), .B1(new_n16173_), .B2(new_n16171_), .ZN(new_n16178_));
  NAND3_X1   g15848(.A1(new_n16102_), .A2(new_n16008_), .A3(new_n16178_), .ZN(new_n16179_));
  NAND2_X1   g15849(.A1(new_n16179_), .A2(new_n16177_), .ZN(new_n16180_));
  NOR2_X1    g15850(.A1(new_n16116_), .A2(new_n16114_), .ZN(new_n16181_));
  XOR2_X1    g15851(.A1(new_n16111_), .A2(new_n16117_), .Z(new_n16182_));
  AOI21_X1   g15852(.A1(new_n16116_), .A2(new_n16114_), .B(new_n16182_), .ZN(new_n16183_));
  NOR2_X1    g15853(.A1(new_n16183_), .A2(new_n16181_), .ZN(new_n16184_));
  AOI21_X1   g15854(.A1(new_n7186_), .A2(new_n8455_), .B(new_n16143_), .ZN(new_n16185_));
  INV_X1     g15855(.I(new_n16185_), .ZN(new_n16186_));
  AOI21_X1   g15856(.A1(new_n6030_), .A2(new_n8242_), .B(new_n16147_), .ZN(new_n16187_));
  NOR2_X1    g15857(.A1(new_n16151_), .A2(new_n16150_), .ZN(new_n16188_));
  INV_X1     g15858(.I(new_n16188_), .ZN(new_n16189_));
  XOR2_X1    g15859(.A1(new_n16187_), .A2(new_n16189_), .Z(new_n16190_));
  NOR2_X1    g15860(.A1(new_n16190_), .A2(new_n16186_), .ZN(new_n16191_));
  INV_X1     g15861(.I(new_n16187_), .ZN(new_n16192_));
  NOR2_X1    g15862(.A1(new_n16192_), .A2(new_n16189_), .ZN(new_n16193_));
  NOR2_X1    g15863(.A1(new_n16187_), .A2(new_n16188_), .ZN(new_n16194_));
  NOR2_X1    g15864(.A1(new_n16193_), .A2(new_n16194_), .ZN(new_n16195_));
  NOR2_X1    g15865(.A1(new_n16195_), .A2(new_n16185_), .ZN(new_n16196_));
  NOR2_X1    g15866(.A1(new_n16196_), .A2(new_n16191_), .ZN(new_n16197_));
  INV_X1     g15867(.I(new_n16145_), .ZN(new_n16198_));
  AOI21_X1   g15868(.A1(new_n16198_), .A2(new_n16157_), .B(new_n16155_), .ZN(new_n16199_));
  XOR2_X1    g15869(.A1(new_n16197_), .A2(new_n16199_), .Z(new_n16200_));
  NOR2_X1    g15870(.A1(new_n16200_), .A2(new_n16184_), .ZN(new_n16201_));
  INV_X1     g15871(.I(new_n16197_), .ZN(new_n16202_));
  NOR2_X1    g15872(.A1(new_n16202_), .A2(new_n16199_), .ZN(new_n16203_));
  NAND2_X1   g15873(.A1(new_n16202_), .A2(new_n16199_), .ZN(new_n16204_));
  INV_X1     g15874(.I(new_n16204_), .ZN(new_n16205_));
  NOR2_X1    g15875(.A1(new_n16205_), .A2(new_n16203_), .ZN(new_n16206_));
  INV_X1     g15876(.I(new_n16206_), .ZN(new_n16207_));
  AOI21_X1   g15877(.A1(new_n16207_), .A2(new_n16184_), .B(new_n16201_), .ZN(new_n16208_));
  OAI21_X1   g15878(.A1(new_n16108_), .A2(new_n16123_), .B(new_n16124_), .ZN(new_n16209_));
  AND2_X2    g15879(.A1(new_n16162_), .A2(new_n16141_), .Z(new_n16210_));
  NOR2_X1    g15880(.A1(new_n16210_), .A2(new_n16161_), .ZN(new_n16211_));
  NAND2_X1   g15881(.A1(new_n16128_), .A2(new_n16139_), .ZN(new_n16212_));
  NOR2_X1    g15882(.A1(new_n10786_), .A2(new_n12160_), .ZN(new_n16213_));
  INV_X1     g15883(.I(new_n16213_), .ZN(new_n16214_));
  NOR4_X1    g15884(.A1(new_n16214_), .A2(new_n6779_), .A3(new_n7483_), .A4(new_n11658_), .ZN(new_n16215_));
  NAND2_X1   g15885(.A1(\a[43] ), .A2(\a[53] ), .ZN(new_n16216_));
  NAND2_X1   g15886(.A1(\a[52] ), .A2(\a[62] ), .ZN(new_n16217_));
  XNOR2_X1   g15887(.A1(new_n16216_), .A2(new_n16217_), .ZN(new_n16218_));
  XOR2_X1    g15888(.A1(new_n16215_), .A2(new_n16218_), .Z(new_n16219_));
  AOI21_X1   g15889(.A1(new_n16137_), .A2(new_n16212_), .B(new_n16219_), .ZN(new_n16220_));
  NAND2_X1   g15890(.A1(new_n16212_), .A2(new_n16137_), .ZN(new_n16221_));
  INV_X1     g15891(.I(new_n16215_), .ZN(new_n16222_));
  NOR2_X1    g15892(.A1(new_n16222_), .A2(new_n16218_), .ZN(new_n16223_));
  INV_X1     g15893(.I(new_n16223_), .ZN(new_n16224_));
  NAND2_X1   g15894(.A1(new_n16222_), .A2(new_n16218_), .ZN(new_n16225_));
  AOI21_X1   g15895(.A1(new_n16224_), .A2(new_n16225_), .B(new_n16221_), .ZN(new_n16226_));
  NOR2_X1    g15896(.A1(new_n16220_), .A2(new_n16226_), .ZN(new_n16227_));
  AOI22_X1   g15897(.A1(new_n4771_), .A2(new_n9781_), .B1(new_n11018_), .B2(new_n15852_), .ZN(new_n16228_));
  INV_X1     g15898(.I(new_n16228_), .ZN(new_n16229_));
  NAND4_X1   g15899(.A1(new_n16229_), .A2(new_n5743_), .A3(new_n8992_), .A4(new_n16110_), .ZN(new_n16230_));
  NAND2_X1   g15900(.A1(new_n16117_), .A2(new_n5350_), .ZN(new_n16231_));
  OAI21_X1   g15901(.A1(new_n16111_), .A2(new_n9550_), .B(new_n16231_), .ZN(new_n16232_));
  OAI22_X1   g15902(.A1(new_n8675_), .A2(new_n8677_), .B1(new_n8199_), .B2(new_n5793_), .ZN(new_n16233_));
  NAND4_X1   g15903(.A1(new_n7693_), .A2(new_n8246_), .A3(\a[46] ), .A4(\a[59] ), .ZN(new_n16234_));
  NOR2_X1    g15904(.A1(new_n16233_), .A2(new_n16234_), .ZN(new_n16235_));
  XNOR2_X1   g15905(.A1(new_n16232_), .A2(new_n16235_), .ZN(new_n16236_));
  NOR2_X1    g15906(.A1(new_n16236_), .A2(new_n16230_), .ZN(new_n16237_));
  INV_X1     g15907(.I(new_n16230_), .ZN(new_n16238_));
  INV_X1     g15908(.I(new_n16232_), .ZN(new_n16239_));
  INV_X1     g15909(.I(new_n16235_), .ZN(new_n16240_));
  NOR2_X1    g15910(.A1(new_n16239_), .A2(new_n16240_), .ZN(new_n16241_));
  NOR2_X1    g15911(.A1(new_n16232_), .A2(new_n16235_), .ZN(new_n16242_));
  NOR2_X1    g15912(.A1(new_n16241_), .A2(new_n16242_), .ZN(new_n16243_));
  NOR2_X1    g15913(.A1(new_n16243_), .A2(new_n16238_), .ZN(new_n16244_));
  NOR2_X1    g15914(.A1(new_n16244_), .A2(new_n16237_), .ZN(new_n16245_));
  XNOR2_X1   g15915(.A1(new_n16227_), .A2(new_n16245_), .ZN(new_n16246_));
  NOR2_X1    g15916(.A1(new_n16246_), .A2(new_n16211_), .ZN(new_n16247_));
  OAI22_X1   g15917(.A1(new_n16220_), .A2(new_n16226_), .B1(new_n16237_), .B2(new_n16244_), .ZN(new_n16248_));
  NAND2_X1   g15918(.A1(new_n16227_), .A2(new_n16245_), .ZN(new_n16249_));
  NAND2_X1   g15919(.A1(new_n16249_), .A2(new_n16248_), .ZN(new_n16250_));
  AOI21_X1   g15920(.A1(new_n16211_), .A2(new_n16250_), .B(new_n16247_), .ZN(new_n16251_));
  NOR2_X1    g15921(.A1(new_n16209_), .A2(new_n16251_), .ZN(new_n16252_));
  INV_X1     g15922(.I(new_n16252_), .ZN(new_n16253_));
  NAND2_X1   g15923(.A1(new_n16209_), .A2(new_n16251_), .ZN(new_n16254_));
  AOI21_X1   g15924(.A1(new_n16253_), .A2(new_n16254_), .B(new_n16208_), .ZN(new_n16255_));
  XOR2_X1    g15925(.A1(new_n16209_), .A2(new_n16251_), .Z(new_n16256_));
  AOI21_X1   g15926(.A1(new_n16208_), .A2(new_n16256_), .B(new_n16255_), .ZN(new_n16257_));
  AOI21_X1   g15927(.A1(new_n16107_), .A2(new_n16168_), .B(new_n16170_), .ZN(new_n16258_));
  XNOR2_X1   g15928(.A1(new_n16257_), .A2(new_n16258_), .ZN(new_n16259_));
  NAND2_X1   g15929(.A1(new_n16180_), .A2(new_n16259_), .ZN(new_n16260_));
  XNOR2_X1   g15930(.A1(new_n16257_), .A2(new_n16258_), .ZN(new_n16261_));
  OAI21_X1   g15931(.A1(new_n16180_), .A2(new_n16261_), .B(new_n16260_), .ZN(\asquared[106] ));
  INV_X1     g15932(.I(new_n16258_), .ZN(new_n16263_));
  NAND2_X1   g15933(.A1(new_n16263_), .A2(new_n16257_), .ZN(new_n16264_));
  OAI21_X1   g15934(.A1(new_n16257_), .A2(new_n16263_), .B(new_n16180_), .ZN(new_n16265_));
  NAND2_X1   g15935(.A1(new_n16265_), .A2(new_n16264_), .ZN(new_n16266_));
  NOR2_X1    g15936(.A1(new_n16205_), .A2(new_n16184_), .ZN(new_n16267_));
  NOR2_X1    g15937(.A1(new_n16267_), .A2(new_n16203_), .ZN(new_n16268_));
  OAI22_X1   g15938(.A1(new_n8941_), .A2(new_n11001_), .B1(new_n7422_), .B2(new_n8953_), .ZN(new_n16269_));
  OAI21_X1   g15939(.A1(new_n10034_), .A2(new_n8005_), .B(new_n16269_), .ZN(new_n16270_));
  NOR2_X1    g15940(.A1(new_n16270_), .A2(new_n10290_), .ZN(new_n16271_));
  OAI21_X1   g15941(.A1(new_n16271_), .A2(\a[55] ), .B(\a[51] ), .ZN(new_n16272_));
  NAND3_X1   g15942(.A1(new_n16272_), .A2(new_n6055_), .A3(new_n7216_), .ZN(new_n16273_));
  AOI21_X1   g15943(.A1(new_n6777_), .A2(new_n7483_), .B(new_n16269_), .ZN(new_n16274_));
  NAND2_X1   g15944(.A1(new_n16273_), .A2(new_n16274_), .ZN(new_n16275_));
  INV_X1     g15945(.I(new_n16194_), .ZN(new_n16276_));
  AOI21_X1   g15946(.A1(new_n16185_), .A2(new_n16276_), .B(new_n16193_), .ZN(new_n16277_));
  AOI21_X1   g15947(.A1(new_n6027_), .A2(new_n6030_), .B(new_n8678_), .ZN(new_n16278_));
  NOR2_X1    g15948(.A1(new_n5511_), .A2(new_n8085_), .ZN(new_n16279_));
  NAND4_X1   g15949(.A1(new_n16278_), .A2(new_n12355_), .A3(new_n8246_), .A4(new_n16279_), .ZN(new_n16280_));
  INV_X1     g15950(.I(new_n16280_), .ZN(new_n16281_));
  NAND2_X1   g15951(.A1(new_n16277_), .A2(new_n16281_), .ZN(new_n16282_));
  INV_X1     g15952(.I(new_n16277_), .ZN(new_n16283_));
  NAND2_X1   g15953(.A1(new_n16283_), .A2(new_n16280_), .ZN(new_n16284_));
  AOI21_X1   g15954(.A1(new_n16284_), .A2(new_n16282_), .B(new_n16275_), .ZN(new_n16285_));
  INV_X1     g15955(.I(new_n16275_), .ZN(new_n16286_));
  NOR2_X1    g15956(.A1(new_n16277_), .A2(new_n16280_), .ZN(new_n16287_));
  NOR2_X1    g15957(.A1(new_n16283_), .A2(new_n16281_), .ZN(new_n16288_));
  NOR2_X1    g15958(.A1(new_n16288_), .A2(new_n16287_), .ZN(new_n16289_));
  NOR2_X1    g15959(.A1(new_n16289_), .A2(new_n16286_), .ZN(new_n16290_));
  NOR2_X1    g15960(.A1(new_n16290_), .A2(new_n16285_), .ZN(new_n16291_));
  INV_X1     g15961(.I(new_n16291_), .ZN(new_n16292_));
  AOI21_X1   g15962(.A1(new_n5742_), .A2(new_n8991_), .B(new_n16229_), .ZN(new_n16293_));
  INV_X1     g15963(.I(new_n16293_), .ZN(new_n16294_));
  NOR2_X1    g15964(.A1(new_n8424_), .A2(new_n8992_), .ZN(new_n16295_));
  NAND4_X1   g15965(.A1(new_n16295_), .A2(\a[46] ), .A3(new_n14214_), .A4(\a[60] ), .ZN(new_n16296_));
  AOI21_X1   g15966(.A1(new_n16296_), .A2(new_n9785_), .B(new_n5743_), .ZN(new_n16297_));
  NOR2_X1    g15967(.A1(new_n8424_), .A2(new_n8992_), .ZN(new_n16298_));
  INV_X1     g15968(.I(new_n16298_), .ZN(new_n16299_));
  OAI21_X1   g15969(.A1(new_n7693_), .A2(new_n8246_), .B(new_n16233_), .ZN(new_n16300_));
  NOR2_X1    g15970(.A1(new_n16300_), .A2(new_n16299_), .ZN(new_n16301_));
  INV_X1     g15971(.I(new_n16301_), .ZN(new_n16302_));
  NAND2_X1   g15972(.A1(new_n16300_), .A2(new_n16299_), .ZN(new_n16303_));
  AOI21_X1   g15973(.A1(new_n16302_), .A2(new_n16303_), .B(new_n16294_), .ZN(new_n16304_));
  XOR2_X1    g15974(.A1(new_n16300_), .A2(new_n16298_), .Z(new_n16305_));
  NOR2_X1    g15975(.A1(new_n16305_), .A2(new_n16293_), .ZN(new_n16306_));
  NOR2_X1    g15976(.A1(new_n16306_), .A2(new_n16304_), .ZN(new_n16307_));
  NOR2_X1    g15977(.A1(new_n16292_), .A2(new_n16307_), .ZN(new_n16308_));
  NOR3_X1    g15978(.A1(new_n16291_), .A2(new_n16304_), .A3(new_n16306_), .ZN(new_n16309_));
  NOR2_X1    g15979(.A1(new_n16308_), .A2(new_n16309_), .ZN(new_n16310_));
  NOR2_X1    g15980(.A1(new_n16310_), .A2(new_n16268_), .ZN(new_n16311_));
  INV_X1     g15981(.I(new_n16268_), .ZN(new_n16312_));
  XOR2_X1    g15982(.A1(new_n16291_), .A2(new_n16307_), .Z(new_n16313_));
  NOR2_X1    g15983(.A1(new_n16313_), .A2(new_n16312_), .ZN(new_n16314_));
  NOR2_X1    g15984(.A1(new_n16311_), .A2(new_n16314_), .ZN(new_n16315_));
  AOI21_X1   g15985(.A1(new_n16221_), .A2(new_n16225_), .B(new_n16223_), .ZN(new_n16316_));
  INV_X1     g15986(.I(new_n16316_), .ZN(new_n16317_));
  NOR2_X1    g15987(.A1(new_n16242_), .A2(new_n16230_), .ZN(new_n16318_));
  NOR2_X1    g15988(.A1(new_n16318_), .A2(new_n16241_), .ZN(new_n16319_));
  INV_X1     g15989(.I(new_n16319_), .ZN(new_n16320_));
  AOI21_X1   g15990(.A1(new_n6779_), .A2(new_n7483_), .B(new_n16213_), .ZN(new_n16321_));
  INV_X1     g15991(.I(new_n16321_), .ZN(new_n16322_));
  NOR2_X1    g15992(.A1(new_n7204_), .A2(\a[62] ), .ZN(new_n16323_));
  OAI21_X1   g15993(.A1(new_n16322_), .A2(new_n16323_), .B(\a[43] ), .ZN(new_n16324_));
  XOR2_X1    g15994(.A1(new_n16324_), .A2(\a[63] ), .Z(new_n16325_));
  XOR2_X1    g15995(.A1(new_n16325_), .A2(new_n16320_), .Z(new_n16326_));
  NAND2_X1   g15996(.A1(new_n16326_), .A2(new_n16317_), .ZN(new_n16327_));
  NOR2_X1    g15997(.A1(new_n16325_), .A2(new_n16320_), .ZN(new_n16328_));
  NAND2_X1   g15998(.A1(new_n16325_), .A2(new_n16320_), .ZN(new_n16329_));
  INV_X1     g15999(.I(new_n16329_), .ZN(new_n16330_));
  OAI21_X1   g16000(.A1(new_n16330_), .A2(new_n16328_), .B(new_n16316_), .ZN(new_n16331_));
  NAND2_X1   g16001(.A1(new_n16327_), .A2(new_n16331_), .ZN(new_n16332_));
  INV_X1     g16002(.I(new_n16332_), .ZN(new_n16333_));
  OAI21_X1   g16003(.A1(new_n16210_), .A2(new_n16161_), .B(new_n16248_), .ZN(new_n16334_));
  NAND2_X1   g16004(.A1(new_n16334_), .A2(new_n16249_), .ZN(new_n16335_));
  NAND2_X1   g16005(.A1(new_n16333_), .A2(new_n16335_), .ZN(new_n16336_));
  INV_X1     g16006(.I(new_n16336_), .ZN(new_n16337_));
  NOR2_X1    g16007(.A1(new_n16333_), .A2(new_n16335_), .ZN(new_n16338_));
  NOR2_X1    g16008(.A1(new_n16337_), .A2(new_n16338_), .ZN(new_n16339_));
  XNOR2_X1   g16009(.A1(new_n16335_), .A2(new_n16332_), .ZN(new_n16340_));
  NAND2_X1   g16010(.A1(new_n16315_), .A2(new_n16340_), .ZN(new_n16341_));
  OAI21_X1   g16011(.A1(new_n16315_), .A2(new_n16339_), .B(new_n16341_), .ZN(new_n16342_));
  NAND2_X1   g16012(.A1(new_n16253_), .A2(new_n16208_), .ZN(new_n16343_));
  NAND2_X1   g16013(.A1(new_n16343_), .A2(new_n16254_), .ZN(new_n16344_));
  NOR2_X1    g16014(.A1(new_n16344_), .A2(new_n16342_), .ZN(new_n16345_));
  INV_X1     g16015(.I(new_n16345_), .ZN(new_n16346_));
  NAND2_X1   g16016(.A1(new_n16344_), .A2(new_n16342_), .ZN(new_n16347_));
  NAND2_X1   g16017(.A1(new_n16346_), .A2(new_n16347_), .ZN(new_n16348_));
  XOR2_X1    g16018(.A1(new_n16266_), .A2(new_n16348_), .Z(\asquared[107] ));
  NAND2_X1   g16019(.A1(new_n16347_), .A2(new_n16257_), .ZN(new_n16350_));
  OAI21_X1   g16020(.A1(new_n16347_), .A2(new_n16257_), .B(new_n16258_), .ZN(new_n16351_));
  NAND2_X1   g16021(.A1(new_n16351_), .A2(new_n16350_), .ZN(new_n16352_));
  AOI21_X1   g16022(.A1(new_n16179_), .A2(new_n16177_), .B(new_n16352_), .ZN(new_n16353_));
  OAI21_X1   g16023(.A1(new_n16315_), .A2(new_n16338_), .B(new_n16336_), .ZN(new_n16354_));
  INV_X1     g16024(.I(new_n16354_), .ZN(new_n16355_));
  INV_X1     g16025(.I(new_n16309_), .ZN(new_n16356_));
  AOI21_X1   g16026(.A1(new_n16312_), .A2(new_n16356_), .B(new_n16308_), .ZN(new_n16357_));
  OAI21_X1   g16027(.A1(new_n16316_), .A2(new_n16328_), .B(new_n16329_), .ZN(new_n16358_));
  INV_X1     g16028(.I(new_n16358_), .ZN(new_n16359_));
  NOR2_X1    g16029(.A1(new_n16297_), .A2(new_n16295_), .ZN(new_n16360_));
  AOI21_X1   g16030(.A1(new_n6028_), .A2(new_n8245_), .B(new_n16278_), .ZN(new_n16361_));
  NOR4_X1    g16031(.A1(new_n4770_), .A2(new_n5750_), .A3(new_n8085_), .A4(new_n9310_), .ZN(new_n16362_));
  AOI21_X1   g16032(.A1(new_n6028_), .A2(new_n8676_), .B(new_n16362_), .ZN(new_n16363_));
  INV_X1     g16033(.I(new_n16363_), .ZN(new_n16364_));
  NOR2_X1    g16034(.A1(new_n7647_), .A2(new_n9310_), .ZN(new_n16365_));
  NOR4_X1    g16035(.A1(new_n8072_), .A2(new_n16365_), .A3(new_n5750_), .A4(new_n8085_), .ZN(new_n16366_));
  NAND2_X1   g16036(.A1(new_n16364_), .A2(new_n16366_), .ZN(new_n16367_));
  INV_X1     g16037(.I(new_n16367_), .ZN(new_n16368_));
  AND2_X2    g16038(.A1(new_n16361_), .A2(new_n16368_), .Z(new_n16369_));
  NOR2_X1    g16039(.A1(new_n16361_), .A2(new_n16368_), .ZN(new_n16370_));
  OAI21_X1   g16040(.A1(new_n16369_), .A2(new_n16370_), .B(new_n16360_), .ZN(new_n16371_));
  INV_X1     g16041(.I(new_n16360_), .ZN(new_n16372_));
  XOR2_X1    g16042(.A1(new_n16361_), .A2(new_n16368_), .Z(new_n16373_));
  NAND2_X1   g16043(.A1(new_n16373_), .A2(new_n16372_), .ZN(new_n16374_));
  NAND2_X1   g16044(.A1(new_n16374_), .A2(new_n16371_), .ZN(new_n16375_));
  NAND2_X1   g16045(.A1(\a[46] ), .A2(\a[60] ), .ZN(new_n16376_));
  NAND2_X1   g16046(.A1(\a[47] ), .A2(\a[61] ), .ZN(new_n16377_));
  XNOR2_X1   g16047(.A1(new_n16376_), .A2(new_n16377_), .ZN(new_n16378_));
  XOR2_X1    g16048(.A1(new_n16270_), .A2(new_n16378_), .Z(new_n16379_));
  AOI22_X1   g16049(.A1(new_n6779_), .A2(new_n10958_), .B1(new_n6776_), .B2(new_n8242_), .ZN(new_n16380_));
  NOR2_X1    g16050(.A1(new_n10034_), .A2(new_n8953_), .ZN(new_n16381_));
  AOI21_X1   g16051(.A1(\a[51] ), .A2(\a[56] ), .B(new_n11670_), .ZN(new_n16382_));
  NOR4_X1    g16052(.A1(new_n16381_), .A2(new_n6055_), .A3(new_n7727_), .A4(new_n16382_), .ZN(new_n16383_));
  NAND2_X1   g16053(.A1(new_n16383_), .A2(new_n16380_), .ZN(new_n16384_));
  NOR2_X1    g16054(.A1(new_n6945_), .A2(\a[53] ), .ZN(new_n16385_));
  XOR2_X1    g16055(.A1(new_n14539_), .A2(new_n16385_), .Z(new_n16386_));
  NOR2_X1    g16056(.A1(new_n16384_), .A2(new_n16386_), .ZN(new_n16387_));
  INV_X1     g16057(.I(new_n16387_), .ZN(new_n16388_));
  NAND2_X1   g16058(.A1(new_n16384_), .A2(new_n16386_), .ZN(new_n16389_));
  AOI21_X1   g16059(.A1(new_n16388_), .A2(new_n16389_), .B(new_n16379_), .ZN(new_n16390_));
  INV_X1     g16060(.I(new_n16379_), .ZN(new_n16391_));
  XNOR2_X1   g16061(.A1(new_n16384_), .A2(new_n16386_), .ZN(new_n16392_));
  NOR2_X1    g16062(.A1(new_n16391_), .A2(new_n16392_), .ZN(new_n16393_));
  NOR2_X1    g16063(.A1(new_n16393_), .A2(new_n16390_), .ZN(new_n16394_));
  XOR2_X1    g16064(.A1(new_n16375_), .A2(new_n16394_), .Z(new_n16395_));
  INV_X1     g16065(.I(new_n16375_), .ZN(new_n16396_));
  NOR2_X1    g16066(.A1(new_n16396_), .A2(new_n16394_), .ZN(new_n16397_));
  NAND2_X1   g16067(.A1(new_n16396_), .A2(new_n16394_), .ZN(new_n16398_));
  INV_X1     g16068(.I(new_n16398_), .ZN(new_n16399_));
  OAI21_X1   g16069(.A1(new_n16397_), .A2(new_n16399_), .B(new_n16359_), .ZN(new_n16400_));
  OAI21_X1   g16070(.A1(new_n16359_), .A2(new_n16395_), .B(new_n16400_), .ZN(new_n16401_));
  NOR2_X1    g16071(.A1(new_n16288_), .A2(new_n16275_), .ZN(new_n16402_));
  NOR2_X1    g16072(.A1(new_n16402_), .A2(new_n16287_), .ZN(new_n16403_));
  NAND2_X1   g16073(.A1(new_n16303_), .A2(new_n16293_), .ZN(new_n16404_));
  NAND2_X1   g16074(.A1(new_n16404_), .A2(new_n16302_), .ZN(new_n16405_));
  AOI21_X1   g16075(.A1(new_n8056_), .A2(new_n9029_), .B(new_n4501_), .ZN(new_n16406_));
  INV_X1     g16076(.I(new_n16406_), .ZN(new_n16407_));
  NOR2_X1    g16077(.A1(new_n4501_), .A2(new_n9310_), .ZN(new_n16408_));
  OAI21_X1   g16078(.A1(new_n16321_), .A2(new_n16406_), .B(new_n16408_), .ZN(new_n16409_));
  OAI21_X1   g16079(.A1(new_n16322_), .A2(new_n16407_), .B(new_n16409_), .ZN(new_n16410_));
  XNOR2_X1   g16080(.A1(new_n16410_), .A2(new_n16405_), .ZN(new_n16411_));
  AND2_X2    g16081(.A1(new_n16410_), .A2(new_n16405_), .Z(new_n16412_));
  NOR2_X1    g16082(.A1(new_n16410_), .A2(new_n16405_), .ZN(new_n16413_));
  OAI21_X1   g16083(.A1(new_n16412_), .A2(new_n16413_), .B(new_n16403_), .ZN(new_n16414_));
  OAI21_X1   g16084(.A1(new_n16403_), .A2(new_n16411_), .B(new_n16414_), .ZN(new_n16415_));
  XNOR2_X1   g16085(.A1(new_n16401_), .A2(new_n16415_), .ZN(new_n16416_));
  NOR2_X1    g16086(.A1(new_n16416_), .A2(new_n16357_), .ZN(new_n16417_));
  INV_X1     g16087(.I(new_n16357_), .ZN(new_n16418_));
  NAND2_X1   g16088(.A1(new_n16401_), .A2(new_n16415_), .ZN(new_n16419_));
  NOR2_X1    g16089(.A1(new_n16401_), .A2(new_n16415_), .ZN(new_n16420_));
  INV_X1     g16090(.I(new_n16420_), .ZN(new_n16421_));
  AOI21_X1   g16091(.A1(new_n16421_), .A2(new_n16419_), .B(new_n16418_), .ZN(new_n16422_));
  NOR2_X1    g16092(.A1(new_n16417_), .A2(new_n16422_), .ZN(new_n16423_));
  NOR2_X1    g16093(.A1(new_n16423_), .A2(new_n16355_), .ZN(new_n16424_));
  XOR2_X1    g16094(.A1(new_n16353_), .A2(new_n16424_), .Z(new_n16425_));
  XOR2_X1    g16095(.A1(new_n16425_), .A2(new_n16345_), .Z(\asquared[108] ));
  AOI21_X1   g16096(.A1(new_n16355_), .A2(new_n16423_), .B(new_n16346_), .ZN(new_n16427_));
  AOI21_X1   g16097(.A1(new_n16353_), .A2(new_n16427_), .B(new_n16424_), .ZN(new_n16428_));
  AOI21_X1   g16098(.A1(new_n16418_), .A2(new_n16419_), .B(new_n16420_), .ZN(new_n16429_));
  AOI21_X1   g16099(.A1(new_n16358_), .A2(new_n16398_), .B(new_n16397_), .ZN(new_n16430_));
  INV_X1     g16100(.I(new_n16412_), .ZN(new_n16431_));
  OAI21_X1   g16101(.A1(new_n16403_), .A2(new_n16413_), .B(new_n16431_), .ZN(new_n16432_));
  INV_X1     g16102(.I(new_n16432_), .ZN(new_n16433_));
  OAI22_X1   g16103(.A1(new_n16270_), .A2(new_n5793_), .B1(new_n8992_), .B2(new_n16378_), .ZN(new_n16434_));
  NOR2_X1    g16104(.A1(new_n13620_), .A2(new_n15673_), .ZN(new_n16435_));
  NOR4_X1    g16105(.A1(new_n9784_), .A2(new_n5980_), .A3(new_n5004_), .A4(new_n9310_), .ZN(new_n16436_));
  NAND2_X1   g16106(.A1(new_n16435_), .A2(new_n16436_), .ZN(new_n16437_));
  NOR2_X1    g16107(.A1(new_n13260_), .A2(new_n12355_), .ZN(new_n16438_));
  NOR2_X1    g16108(.A1(new_n9556_), .A2(new_n16438_), .ZN(new_n16439_));
  NOR4_X1    g16109(.A1(new_n6280_), .A2(new_n8676_), .A3(new_n5750_), .A4(new_n8990_), .ZN(new_n16440_));
  NAND2_X1   g16110(.A1(new_n16439_), .A2(new_n16440_), .ZN(new_n16441_));
  XNOR2_X1   g16111(.A1(new_n16437_), .A2(new_n16441_), .ZN(new_n16442_));
  INV_X1     g16112(.I(new_n16442_), .ZN(new_n16443_));
  NOR2_X1    g16113(.A1(new_n16437_), .A2(new_n16441_), .ZN(new_n16444_));
  INV_X1     g16114(.I(new_n16444_), .ZN(new_n16445_));
  NAND2_X1   g16115(.A1(new_n16437_), .A2(new_n16441_), .ZN(new_n16446_));
  AOI21_X1   g16116(.A1(new_n16445_), .A2(new_n16446_), .B(new_n16434_), .ZN(new_n16447_));
  AOI21_X1   g16117(.A1(new_n16434_), .A2(new_n16443_), .B(new_n16447_), .ZN(new_n16448_));
  AOI21_X1   g16118(.A1(new_n8072_), .A2(new_n16365_), .B(new_n16364_), .ZN(new_n16449_));
  INV_X1     g16119(.I(new_n16449_), .ZN(new_n16450_));
  NOR2_X1    g16120(.A1(new_n16381_), .A2(new_n16380_), .ZN(new_n16451_));
  OAI21_X1   g16121(.A1(new_n14539_), .A2(\a[53] ), .B(\a[54] ), .ZN(new_n16452_));
  INV_X1     g16122(.I(new_n16452_), .ZN(new_n16453_));
  XOR2_X1    g16123(.A1(new_n16451_), .A2(new_n16453_), .Z(new_n16454_));
  NOR2_X1    g16124(.A1(new_n16454_), .A2(new_n16450_), .ZN(new_n16455_));
  INV_X1     g16125(.I(new_n16451_), .ZN(new_n16456_));
  NOR2_X1    g16126(.A1(new_n16456_), .A2(new_n16453_), .ZN(new_n16457_));
  NOR2_X1    g16127(.A1(new_n16451_), .A2(new_n16452_), .ZN(new_n16458_));
  NOR2_X1    g16128(.A1(new_n16457_), .A2(new_n16458_), .ZN(new_n16459_));
  NOR2_X1    g16129(.A1(new_n16459_), .A2(new_n16449_), .ZN(new_n16460_));
  NOR2_X1    g16130(.A1(new_n16460_), .A2(new_n16455_), .ZN(new_n16461_));
  XNOR2_X1   g16131(.A1(new_n16448_), .A2(new_n16461_), .ZN(new_n16462_));
  NOR2_X1    g16132(.A1(new_n16433_), .A2(new_n16462_), .ZN(new_n16463_));
  NOR2_X1    g16133(.A1(new_n16448_), .A2(new_n16461_), .ZN(new_n16464_));
  INV_X1     g16134(.I(new_n16464_), .ZN(new_n16465_));
  NAND2_X1   g16135(.A1(new_n16448_), .A2(new_n16461_), .ZN(new_n16466_));
  AOI21_X1   g16136(.A1(new_n16465_), .A2(new_n16466_), .B(new_n16432_), .ZN(new_n16467_));
  NOR2_X1    g16137(.A1(new_n16463_), .A2(new_n16467_), .ZN(new_n16468_));
  NOR2_X1    g16138(.A1(new_n16372_), .A2(new_n16370_), .ZN(new_n16469_));
  NOR2_X1    g16139(.A1(new_n16469_), .A2(new_n16369_), .ZN(new_n16470_));
  AOI22_X1   g16140(.A1(new_n6777_), .A2(new_n10958_), .B1(new_n7000_), .B2(new_n8242_), .ZN(new_n16471_));
  INV_X1     g16141(.I(new_n16471_), .ZN(new_n16472_));
  NAND2_X1   g16142(.A1(new_n7204_), .A2(new_n8755_), .ZN(new_n16473_));
  NAND2_X1   g16143(.A1(new_n16472_), .A2(new_n16473_), .ZN(new_n16474_));
  OAI21_X1   g16144(.A1(new_n16474_), .A2(new_n7486_), .B(new_n7216_), .ZN(new_n16475_));
  NAND2_X1   g16145(.A1(new_n6260_), .A2(new_n7727_), .ZN(new_n16476_));
  AOI21_X1   g16146(.A1(new_n16475_), .A2(\a[52] ), .B(new_n16476_), .ZN(new_n16477_));
  NAND2_X1   g16147(.A1(new_n16471_), .A2(new_n16473_), .ZN(new_n16478_));
  NOR2_X1    g16148(.A1(new_n16477_), .A2(new_n16478_), .ZN(new_n16479_));
  INV_X1     g16149(.I(new_n16479_), .ZN(new_n16480_));
  NAND2_X1   g16150(.A1(new_n16391_), .A2(new_n16389_), .ZN(new_n16481_));
  NAND2_X1   g16151(.A1(new_n16481_), .A2(new_n16388_), .ZN(new_n16482_));
  INV_X1     g16152(.I(new_n16482_), .ZN(new_n16483_));
  NOR2_X1    g16153(.A1(new_n16483_), .A2(new_n16480_), .ZN(new_n16484_));
  NOR2_X1    g16154(.A1(new_n16482_), .A2(new_n16479_), .ZN(new_n16485_));
  NOR2_X1    g16155(.A1(new_n16484_), .A2(new_n16485_), .ZN(new_n16486_));
  NOR2_X1    g16156(.A1(new_n16486_), .A2(new_n16470_), .ZN(new_n16487_));
  INV_X1     g16157(.I(new_n16470_), .ZN(new_n16488_));
  XOR2_X1    g16158(.A1(new_n16482_), .A2(new_n16480_), .Z(new_n16489_));
  NOR2_X1    g16159(.A1(new_n16489_), .A2(new_n16488_), .ZN(new_n16490_));
  NOR2_X1    g16160(.A1(new_n16487_), .A2(new_n16490_), .ZN(new_n16491_));
  INV_X1     g16161(.I(new_n16491_), .ZN(new_n16492_));
  NAND2_X1   g16162(.A1(new_n16468_), .A2(new_n16492_), .ZN(new_n16493_));
  NOR2_X1    g16163(.A1(new_n16468_), .A2(new_n16492_), .ZN(new_n16494_));
  INV_X1     g16164(.I(new_n16494_), .ZN(new_n16495_));
  AOI21_X1   g16165(.A1(new_n16495_), .A2(new_n16493_), .B(new_n16430_), .ZN(new_n16496_));
  XOR2_X1    g16166(.A1(new_n16468_), .A2(new_n16492_), .Z(new_n16497_));
  AOI21_X1   g16167(.A1(new_n16430_), .A2(new_n16497_), .B(new_n16496_), .ZN(new_n16498_));
  NOR2_X1    g16168(.A1(new_n16498_), .A2(new_n16429_), .ZN(new_n16499_));
  NAND2_X1   g16169(.A1(new_n16498_), .A2(new_n16429_), .ZN(new_n16500_));
  INV_X1     g16170(.I(new_n16500_), .ZN(new_n16501_));
  NOR2_X1    g16171(.A1(new_n16501_), .A2(new_n16499_), .ZN(new_n16502_));
  XOR2_X1    g16172(.A1(new_n16428_), .A2(new_n16502_), .Z(\asquared[109] ));
  INV_X1     g16173(.I(new_n16499_), .ZN(new_n16504_));
  NAND2_X1   g16174(.A1(new_n16428_), .A2(new_n16504_), .ZN(new_n16505_));
  NAND2_X1   g16175(.A1(new_n16505_), .A2(new_n16500_), .ZN(new_n16506_));
  OAI21_X1   g16176(.A1(new_n16433_), .A2(new_n16464_), .B(new_n16466_), .ZN(new_n16507_));
  INV_X1     g16177(.I(new_n16485_), .ZN(new_n16508_));
  AOI21_X1   g16178(.A1(new_n16488_), .A2(new_n16508_), .B(new_n16484_), .ZN(new_n16509_));
  OAI22_X1   g16179(.A1(new_n9556_), .A2(new_n16438_), .B1(new_n7512_), .B2(new_n8677_), .ZN(new_n16510_));
  NOR2_X1    g16180(.A1(new_n16474_), .A2(new_n16510_), .ZN(new_n16511_));
  XOR2_X1    g16181(.A1(new_n16511_), .A2(new_n5175_), .Z(new_n16512_));
  XOR2_X1    g16182(.A1(new_n16512_), .A2(\a[63] ), .Z(new_n16513_));
  AOI21_X1   g16183(.A1(new_n5980_), .A2(new_n9784_), .B(new_n16435_), .ZN(new_n16514_));
  AOI22_X1   g16184(.A1(new_n6056_), .A2(new_n8991_), .B1(new_n6028_), .B2(new_n8455_), .ZN(new_n16515_));
  NOR4_X1    g16185(.A1(new_n6280_), .A2(new_n8996_), .A3(new_n5750_), .A4(new_n8453_), .ZN(new_n16516_));
  NAND2_X1   g16186(.A1(new_n16515_), .A2(new_n16516_), .ZN(new_n16517_));
  AOI21_X1   g16187(.A1(new_n6777_), .A2(new_n7000_), .B(new_n8247_), .ZN(new_n16518_));
  NOR4_X1    g16188(.A1(new_n7204_), .A2(new_n8242_), .A3(new_n6260_), .A4(new_n7647_), .ZN(new_n16519_));
  NAND2_X1   g16189(.A1(new_n16518_), .A2(new_n16519_), .ZN(new_n16520_));
  XOR2_X1    g16190(.A1(new_n16520_), .A2(new_n16517_), .Z(new_n16521_));
  NAND2_X1   g16191(.A1(new_n16521_), .A2(new_n16514_), .ZN(new_n16522_));
  INV_X1     g16192(.I(new_n16514_), .ZN(new_n16523_));
  NOR2_X1    g16193(.A1(new_n16520_), .A2(new_n16517_), .ZN(new_n16524_));
  NAND2_X1   g16194(.A1(new_n16520_), .A2(new_n16517_), .ZN(new_n16525_));
  INV_X1     g16195(.I(new_n16525_), .ZN(new_n16526_));
  OAI21_X1   g16196(.A1(new_n16526_), .A2(new_n16524_), .B(new_n16523_), .ZN(new_n16527_));
  NAND2_X1   g16197(.A1(new_n16522_), .A2(new_n16527_), .ZN(new_n16528_));
  XOR2_X1    g16198(.A1(new_n16513_), .A2(new_n16528_), .Z(new_n16529_));
  NOR2_X1    g16199(.A1(new_n16509_), .A2(new_n16529_), .ZN(new_n16530_));
  INV_X1     g16200(.I(new_n16528_), .ZN(new_n16531_));
  NOR2_X1    g16201(.A1(new_n16513_), .A2(new_n16531_), .ZN(new_n16532_));
  INV_X1     g16202(.I(new_n16532_), .ZN(new_n16533_));
  NAND2_X1   g16203(.A1(new_n16513_), .A2(new_n16531_), .ZN(new_n16534_));
  NAND2_X1   g16204(.A1(new_n16533_), .A2(new_n16534_), .ZN(new_n16535_));
  AOI21_X1   g16205(.A1(new_n16509_), .A2(new_n16535_), .B(new_n16530_), .ZN(new_n16536_));
  AOI21_X1   g16206(.A1(new_n16434_), .A2(new_n16446_), .B(new_n16444_), .ZN(new_n16537_));
  NOR2_X1    g16207(.A1(new_n16450_), .A2(new_n16458_), .ZN(new_n16538_));
  NOR2_X1    g16208(.A1(new_n16538_), .A2(new_n16457_), .ZN(new_n16539_));
  NOR2_X1    g16209(.A1(new_n6999_), .A2(\a[54] ), .ZN(new_n16540_));
  XOR2_X1    g16210(.A1(new_n15037_), .A2(new_n16540_), .Z(new_n16541_));
  XNOR2_X1   g16211(.A1(new_n16539_), .A2(new_n16541_), .ZN(new_n16542_));
  NOR2_X1    g16212(.A1(new_n16539_), .A2(new_n16541_), .ZN(new_n16543_));
  INV_X1     g16213(.I(new_n16543_), .ZN(new_n16544_));
  NAND2_X1   g16214(.A1(new_n16539_), .A2(new_n16541_), .ZN(new_n16545_));
  NAND2_X1   g16215(.A1(new_n16544_), .A2(new_n16545_), .ZN(new_n16546_));
  NAND2_X1   g16216(.A1(new_n16546_), .A2(new_n16537_), .ZN(new_n16547_));
  OAI21_X1   g16217(.A1(new_n16537_), .A2(new_n16542_), .B(new_n16547_), .ZN(new_n16548_));
  XOR2_X1    g16218(.A1(new_n16536_), .A2(new_n16548_), .Z(new_n16549_));
  NAND2_X1   g16219(.A1(new_n16549_), .A2(new_n16507_), .ZN(new_n16550_));
  XOR2_X1    g16220(.A1(new_n16536_), .A2(new_n16548_), .Z(new_n16551_));
  OAI21_X1   g16221(.A1(new_n16507_), .A2(new_n16551_), .B(new_n16550_), .ZN(new_n16552_));
  OAI21_X1   g16222(.A1(new_n16430_), .A2(new_n16494_), .B(new_n16493_), .ZN(new_n16553_));
  XNOR2_X1   g16223(.A1(new_n16552_), .A2(new_n16553_), .ZN(new_n16554_));
  XNOR2_X1   g16224(.A1(new_n16552_), .A2(new_n16553_), .ZN(new_n16555_));
  NAND2_X1   g16225(.A1(new_n16506_), .A2(new_n16555_), .ZN(new_n16556_));
  OAI21_X1   g16226(.A1(new_n16506_), .A2(new_n16554_), .B(new_n16556_), .ZN(\asquared[110] ));
  NOR2_X1    g16227(.A1(new_n16552_), .A2(new_n16553_), .ZN(new_n16558_));
  NAND3_X1   g16228(.A1(new_n16501_), .A2(new_n16552_), .A3(new_n16553_), .ZN(new_n16559_));
  AOI21_X1   g16229(.A1(new_n16428_), .A2(new_n16559_), .B(new_n16504_), .ZN(new_n16560_));
  AND2_X2    g16230(.A1(new_n16560_), .A2(new_n16558_), .Z(\asquared[111] ));
  OAI21_X1   g16231(.A1(new_n16509_), .A2(new_n16532_), .B(new_n16534_), .ZN(new_n16562_));
  NOR2_X1    g16232(.A1(new_n5750_), .A2(new_n9310_), .ZN(new_n16563_));
  XNOR2_X1   g16233(.A1(new_n15037_), .A2(new_n16563_), .ZN(new_n16564_));
  INV_X1     g16234(.I(new_n16564_), .ZN(new_n16565_));
  NAND2_X1   g16235(.A1(\a[46] ), .A2(\a[63] ), .ZN(new_n16566_));
  AOI21_X1   g16236(.A1(new_n16474_), .A2(new_n16510_), .B(new_n16566_), .ZN(new_n16567_));
  NOR2_X1    g16237(.A1(new_n16567_), .A2(new_n16511_), .ZN(new_n16568_));
  NAND3_X1   g16238(.A1(new_n7653_), .A2(\a[52] ), .A3(\a[56] ), .ZN(new_n16569_));
  OAI21_X1   g16239(.A1(new_n8056_), .A2(new_n8246_), .B(new_n16569_), .ZN(new_n16570_));
  NOR2_X1    g16240(.A1(new_n10288_), .A2(new_n8243_), .ZN(new_n16571_));
  INV_X1     g16241(.I(new_n16571_), .ZN(new_n16572_));
  NOR2_X1    g16242(.A1(new_n16570_), .A2(new_n16571_), .ZN(new_n16573_));
  AOI21_X1   g16243(.A1(new_n16573_), .A2(new_n7421_), .B(\a[57] ), .ZN(new_n16574_));
  NOR2_X1    g16244(.A1(\a[52] ), .A2(\a[58] ), .ZN(new_n16575_));
  OAI21_X1   g16245(.A1(new_n16574_), .A2(new_n6694_), .B(new_n16575_), .ZN(new_n16576_));
  NAND3_X1   g16246(.A1(new_n16576_), .A2(new_n16570_), .A3(new_n16572_), .ZN(new_n16577_));
  AOI21_X1   g16247(.A1(new_n15038_), .A2(new_n6945_), .B(new_n6999_), .ZN(new_n16578_));
  XOR2_X1    g16248(.A1(new_n16577_), .A2(new_n16578_), .Z(new_n16579_));
  XOR2_X1    g16249(.A1(new_n16579_), .A2(new_n16568_), .Z(new_n16580_));
  XOR2_X1    g16250(.A1(new_n16580_), .A2(new_n16565_), .Z(new_n16581_));
  AND2_X2    g16251(.A1(new_n16581_), .A2(new_n16562_), .Z(new_n16582_));
  INV_X1     g16252(.I(new_n16545_), .ZN(new_n16583_));
  OAI21_X1   g16253(.A1(new_n16537_), .A2(new_n16583_), .B(new_n16544_), .ZN(new_n16584_));
  AOI21_X1   g16254(.A1(new_n6280_), .A2(new_n8996_), .B(new_n16515_), .ZN(new_n16585_));
  AOI21_X1   g16255(.A1(new_n7204_), .A2(new_n8242_), .B(new_n16518_), .ZN(new_n16586_));
  INV_X1     g16256(.I(new_n16586_), .ZN(new_n16587_));
  NOR2_X1    g16257(.A1(new_n8993_), .A2(new_n10786_), .ZN(new_n16588_));
  NOR4_X1    g16258(.A1(new_n6779_), .A2(new_n8996_), .A3(new_n5745_), .A4(new_n8453_), .ZN(new_n16589_));
  NAND2_X1   g16259(.A1(new_n16588_), .A2(new_n16589_), .ZN(new_n16590_));
  NOR2_X1    g16260(.A1(new_n16587_), .A2(new_n16590_), .ZN(new_n16591_));
  AOI21_X1   g16261(.A1(new_n16588_), .A2(new_n16589_), .B(new_n16586_), .ZN(new_n16592_));
  NOR2_X1    g16262(.A1(new_n16591_), .A2(new_n16592_), .ZN(new_n16593_));
  XOR2_X1    g16263(.A1(new_n16586_), .A2(new_n16590_), .Z(new_n16594_));
  MUX2_X1    g16264(.I0(new_n16594_), .I1(new_n16593_), .S(new_n16585_), .Z(new_n16595_));
  AOI21_X1   g16265(.A1(new_n16514_), .A2(new_n16525_), .B(new_n16524_), .ZN(new_n16596_));
  XOR2_X1    g16266(.A1(new_n16595_), .A2(new_n16596_), .Z(new_n16597_));
  AND2_X2    g16267(.A1(new_n16597_), .A2(new_n16584_), .Z(new_n16598_));
  OR2_X2     g16268(.A1(new_n16595_), .A2(new_n16596_), .Z(new_n16599_));
  NAND2_X1   g16269(.A1(new_n16595_), .A2(new_n16596_), .ZN(new_n16600_));
  AOI21_X1   g16270(.A1(new_n16599_), .A2(new_n16600_), .B(new_n16584_), .ZN(new_n16601_));
  NOR2_X1    g16271(.A1(new_n16581_), .A2(new_n16562_), .ZN(new_n16602_));
  NOR3_X1    g16272(.A1(new_n16602_), .A2(new_n16598_), .A3(new_n16601_), .ZN(new_n16603_));
  NOR2_X1    g16273(.A1(new_n16603_), .A2(new_n16582_), .ZN(new_n16604_));
  NOR2_X1    g16274(.A1(new_n16577_), .A2(new_n16568_), .ZN(new_n16605_));
  XNOR2_X1   g16275(.A1(new_n16564_), .A2(new_n16578_), .ZN(new_n16606_));
  AOI21_X1   g16276(.A1(new_n16577_), .A2(new_n16568_), .B(new_n16606_), .ZN(new_n16607_));
  AOI21_X1   g16277(.A1(new_n6779_), .A2(new_n8996_), .B(new_n16588_), .ZN(new_n16608_));
  INV_X1     g16278(.I(new_n16608_), .ZN(new_n16609_));
  OAI22_X1   g16279(.A1(new_n16564_), .A2(new_n9550_), .B1(new_n7693_), .B2(new_n16578_), .ZN(new_n16610_));
  XNOR2_X1   g16280(.A1(new_n16610_), .A2(new_n16573_), .ZN(new_n16611_));
  NOR2_X1    g16281(.A1(new_n16611_), .A2(new_n16609_), .ZN(new_n16612_));
  AND2_X2    g16282(.A1(new_n16610_), .A2(new_n16573_), .Z(new_n16613_));
  INV_X1     g16283(.I(new_n16613_), .ZN(new_n16614_));
  NOR2_X1    g16284(.A1(new_n16610_), .A2(new_n16573_), .ZN(new_n16615_));
  INV_X1     g16285(.I(new_n16615_), .ZN(new_n16616_));
  AOI21_X1   g16286(.A1(new_n16614_), .A2(new_n16616_), .B(new_n16608_), .ZN(new_n16617_));
  NOR2_X1    g16287(.A1(new_n16617_), .A2(new_n16612_), .ZN(new_n16618_));
  INV_X1     g16288(.I(new_n16592_), .ZN(new_n16619_));
  AOI21_X1   g16289(.A1(new_n16619_), .A2(new_n16585_), .B(new_n16591_), .ZN(new_n16620_));
  XNOR2_X1   g16290(.A1(new_n16618_), .A2(new_n16620_), .ZN(new_n16621_));
  OAI21_X1   g16291(.A1(new_n16605_), .A2(new_n16607_), .B(new_n16621_), .ZN(new_n16622_));
  NOR2_X1    g16292(.A1(new_n16607_), .A2(new_n16605_), .ZN(new_n16623_));
  NOR3_X1    g16293(.A1(new_n16620_), .A2(new_n16617_), .A3(new_n16612_), .ZN(new_n16624_));
  INV_X1     g16294(.I(new_n16620_), .ZN(new_n16625_));
  NOR2_X1    g16295(.A1(new_n16625_), .A2(new_n16618_), .ZN(new_n16626_));
  OAI21_X1   g16296(.A1(new_n16626_), .A2(new_n16624_), .B(new_n16623_), .ZN(new_n16627_));
  NAND2_X1   g16297(.A1(new_n16622_), .A2(new_n16627_), .ZN(new_n16628_));
  NAND2_X1   g16298(.A1(new_n16600_), .A2(new_n16584_), .ZN(new_n16629_));
  AOI22_X1   g16299(.A1(new_n6056_), .A2(new_n15677_), .B1(new_n9781_), .B2(new_n11018_), .ZN(new_n16630_));
  NAND4_X1   g16300(.A1(new_n16630_), .A2(new_n8941_), .A3(new_n8992_), .A4(new_n16563_), .ZN(new_n16631_));
  NOR2_X1    g16301(.A1(new_n8678_), .A2(new_n10722_), .ZN(new_n16632_));
  NOR2_X1    g16302(.A1(new_n10288_), .A2(new_n8246_), .ZN(new_n16633_));
  NOR2_X1    g16303(.A1(new_n6694_), .A2(new_n7647_), .ZN(new_n16634_));
  NOR2_X1    g16304(.A1(new_n12964_), .A2(new_n16634_), .ZN(new_n16635_));
  NOR4_X1    g16305(.A1(new_n16633_), .A2(new_n6692_), .A3(new_n8085_), .A4(new_n16635_), .ZN(new_n16636_));
  NAND2_X1   g16306(.A1(new_n16636_), .A2(new_n16632_), .ZN(new_n16637_));
  NAND2_X1   g16307(.A1(\a[55] ), .A2(\a[62] ), .ZN(new_n16638_));
  XOR2_X1    g16308(.A1(new_n11657_), .A2(new_n16638_), .Z(new_n16639_));
  NOR2_X1    g16309(.A1(new_n16637_), .A2(new_n16639_), .ZN(new_n16640_));
  INV_X1     g16310(.I(new_n16640_), .ZN(new_n16641_));
  NAND2_X1   g16311(.A1(new_n16637_), .A2(new_n16639_), .ZN(new_n16642_));
  AOI21_X1   g16312(.A1(new_n16641_), .A2(new_n16642_), .B(new_n16631_), .ZN(new_n16643_));
  INV_X1     g16313(.I(new_n16631_), .ZN(new_n16644_));
  XNOR2_X1   g16314(.A1(new_n16637_), .A2(new_n16639_), .ZN(new_n16645_));
  NOR2_X1    g16315(.A1(new_n16645_), .A2(new_n16644_), .ZN(new_n16646_));
  NOR2_X1    g16316(.A1(new_n16646_), .A2(new_n16643_), .ZN(new_n16647_));
  AOI21_X1   g16317(.A1(new_n16629_), .A2(new_n16599_), .B(new_n16647_), .ZN(new_n16648_));
  NAND2_X1   g16318(.A1(new_n16629_), .A2(new_n16599_), .ZN(new_n16649_));
  INV_X1     g16319(.I(new_n16647_), .ZN(new_n16650_));
  NOR2_X1    g16320(.A1(new_n16649_), .A2(new_n16650_), .ZN(new_n16651_));
  OAI21_X1   g16321(.A1(new_n16648_), .A2(new_n16651_), .B(new_n16628_), .ZN(new_n16652_));
  XOR2_X1    g16322(.A1(new_n16649_), .A2(new_n16650_), .Z(new_n16653_));
  NAND3_X1   g16323(.A1(new_n16653_), .A2(new_n16622_), .A3(new_n16627_), .ZN(new_n16654_));
  NAND2_X1   g16324(.A1(new_n16654_), .A2(new_n16652_), .ZN(new_n16655_));
  XOR2_X1    g16325(.A1(new_n16604_), .A2(new_n16655_), .Z(new_n16656_));
  NAND2_X1   g16326(.A1(\asquared[111] ), .A2(new_n16656_), .ZN(new_n16657_));
  NAND2_X1   g16327(.A1(new_n16604_), .A2(new_n16655_), .ZN(new_n16658_));
  INV_X1     g16328(.I(new_n16604_), .ZN(new_n16659_));
  INV_X1     g16329(.I(new_n16655_), .ZN(new_n16660_));
  NAND2_X1   g16330(.A1(new_n16659_), .A2(new_n16660_), .ZN(new_n16661_));
  AND2_X2    g16331(.A1(new_n16661_), .A2(new_n16658_), .Z(new_n16662_));
  OAI21_X1   g16332(.A1(\asquared[111] ), .A2(new_n16662_), .B(new_n16657_), .ZN(\asquared[112] ));
  NAND2_X1   g16333(.A1(\asquared[111] ), .A2(new_n16658_), .ZN(new_n16664_));
  NAND2_X1   g16334(.A1(new_n16664_), .A2(new_n16661_), .ZN(new_n16665_));
  NOR2_X1    g16335(.A1(new_n16626_), .A2(new_n16623_), .ZN(new_n16666_));
  NOR2_X1    g16336(.A1(new_n16666_), .A2(new_n16624_), .ZN(new_n16667_));
  NOR2_X1    g16337(.A1(new_n9861_), .A2(new_n6692_), .ZN(new_n16668_));
  NOR2_X1    g16338(.A1(new_n12892_), .A2(new_n6260_), .ZN(new_n16669_));
  NOR3_X1    g16339(.A1(new_n16668_), .A2(new_n16669_), .A3(\a[49] ), .ZN(new_n16670_));
  NOR3_X1    g16340(.A1(new_n16670_), .A2(new_n10034_), .A3(new_n8992_), .ZN(new_n16671_));
  INV_X1     g16341(.I(new_n16671_), .ZN(new_n16672_));
  NOR2_X1    g16342(.A1(new_n5745_), .A2(new_n9310_), .ZN(new_n16673_));
  NOR2_X1    g16343(.A1(new_n6777_), .A2(new_n8991_), .ZN(new_n16674_));
  AOI21_X1   g16344(.A1(new_n16672_), .A2(new_n16673_), .B(new_n16674_), .ZN(new_n16675_));
  AOI22_X1   g16345(.A1(new_n7482_), .A2(new_n8676_), .B1(new_n14034_), .B2(new_n15664_), .ZN(new_n16676_));
  INV_X1     g16346(.I(new_n16676_), .ZN(new_n16677_));
  NOR2_X1    g16347(.A1(new_n8005_), .A2(new_n8246_), .ZN(new_n16678_));
  NOR2_X1    g16348(.A1(new_n16677_), .A2(new_n16678_), .ZN(new_n16679_));
  NAND2_X1   g16349(.A1(new_n16679_), .A2(new_n10958_), .ZN(new_n16680_));
  AOI21_X1   g16350(.A1(new_n16680_), .A2(new_n7647_), .B(new_n6945_), .ZN(new_n16681_));
  NOR3_X1    g16351(.A1(new_n16681_), .A2(\a[53] ), .A3(\a[59] ), .ZN(new_n16682_));
  NOR2_X1    g16352(.A1(new_n16678_), .A2(new_n16676_), .ZN(new_n16683_));
  INV_X1     g16353(.I(new_n16683_), .ZN(new_n16684_));
  NOR2_X1    g16354(.A1(new_n16682_), .A2(new_n16684_), .ZN(new_n16685_));
  AOI21_X1   g16355(.A1(new_n6779_), .A2(new_n8991_), .B(new_n16630_), .ZN(new_n16686_));
  INV_X1     g16356(.I(new_n16686_), .ZN(new_n16687_));
  XOR2_X1    g16357(.A1(new_n16685_), .A2(new_n16687_), .Z(new_n16688_));
  INV_X1     g16358(.I(new_n16685_), .ZN(new_n16689_));
  NOR2_X1    g16359(.A1(new_n16689_), .A2(new_n16687_), .ZN(new_n16690_));
  NOR2_X1    g16360(.A1(new_n16685_), .A2(new_n16686_), .ZN(new_n16691_));
  NOR2_X1    g16361(.A1(new_n16690_), .A2(new_n16691_), .ZN(new_n16692_));
  MUX2_X1    g16362(.I0(new_n16692_), .I1(new_n16688_), .S(new_n16675_), .Z(new_n16693_));
  OAI22_X1   g16363(.A1(new_n8678_), .A2(new_n10722_), .B1(new_n10288_), .B2(new_n8246_), .ZN(new_n16694_));
  NOR2_X1    g16364(.A1(new_n7216_), .A2(new_n9029_), .ZN(new_n16695_));
  INV_X1     g16365(.I(new_n16695_), .ZN(new_n16696_));
  OAI21_X1   g16366(.A1(new_n5745_), .A2(new_n16696_), .B(new_n8953_), .ZN(new_n16697_));
  NOR2_X1    g16367(.A1(new_n16694_), .A2(new_n16697_), .ZN(new_n16698_));
  XOR2_X1    g16368(.A1(new_n16698_), .A2(new_n6055_), .Z(new_n16699_));
  XOR2_X1    g16369(.A1(new_n16699_), .A2(\a[62] ), .Z(new_n16700_));
  NAND2_X1   g16370(.A1(new_n16616_), .A2(new_n16608_), .ZN(new_n16701_));
  NAND2_X1   g16371(.A1(new_n16701_), .A2(new_n16614_), .ZN(new_n16702_));
  INV_X1     g16372(.I(new_n16702_), .ZN(new_n16703_));
  NAND2_X1   g16373(.A1(new_n16642_), .A2(new_n16644_), .ZN(new_n16704_));
  NAND2_X1   g16374(.A1(new_n16704_), .A2(new_n16641_), .ZN(new_n16705_));
  INV_X1     g16375(.I(new_n16705_), .ZN(new_n16706_));
  NOR2_X1    g16376(.A1(new_n16703_), .A2(new_n16706_), .ZN(new_n16707_));
  NOR2_X1    g16377(.A1(new_n16702_), .A2(new_n16705_), .ZN(new_n16708_));
  NOR2_X1    g16378(.A1(new_n16707_), .A2(new_n16708_), .ZN(new_n16709_));
  NOR2_X1    g16379(.A1(new_n16709_), .A2(new_n16700_), .ZN(new_n16710_));
  INV_X1     g16380(.I(new_n16700_), .ZN(new_n16711_));
  XNOR2_X1   g16381(.A1(new_n16702_), .A2(new_n16705_), .ZN(new_n16712_));
  NOR2_X1    g16382(.A1(new_n16712_), .A2(new_n16711_), .ZN(new_n16713_));
  NOR2_X1    g16383(.A1(new_n16710_), .A2(new_n16713_), .ZN(new_n16714_));
  XNOR2_X1   g16384(.A1(new_n16714_), .A2(new_n16693_), .ZN(new_n16715_));
  NOR2_X1    g16385(.A1(new_n16715_), .A2(new_n16667_), .ZN(new_n16716_));
  NOR2_X1    g16386(.A1(new_n16714_), .A2(new_n16693_), .ZN(new_n16717_));
  INV_X1     g16387(.I(new_n16717_), .ZN(new_n16718_));
  NAND2_X1   g16388(.A1(new_n16714_), .A2(new_n16693_), .ZN(new_n16719_));
  NAND2_X1   g16389(.A1(new_n16718_), .A2(new_n16719_), .ZN(new_n16720_));
  AOI21_X1   g16390(.A1(new_n16667_), .A2(new_n16720_), .B(new_n16716_), .ZN(new_n16721_));
  INV_X1     g16391(.I(new_n16721_), .ZN(new_n16722_));
  NOR2_X1    g16392(.A1(new_n16628_), .A2(new_n16651_), .ZN(new_n16723_));
  NOR2_X1    g16393(.A1(new_n16723_), .A2(new_n16648_), .ZN(new_n16724_));
  NOR2_X1    g16394(.A1(new_n16722_), .A2(new_n16724_), .ZN(new_n16725_));
  INV_X1     g16395(.I(new_n16725_), .ZN(new_n16726_));
  NAND2_X1   g16396(.A1(new_n16722_), .A2(new_n16724_), .ZN(new_n16727_));
  NAND2_X1   g16397(.A1(new_n16726_), .A2(new_n16727_), .ZN(new_n16728_));
  XOR2_X1    g16398(.A1(new_n16665_), .A2(new_n16728_), .Z(\asquared[113] ));
  INV_X1     g16399(.I(new_n16424_), .ZN(new_n16730_));
  INV_X1     g16400(.I(new_n16352_), .ZN(new_n16731_));
  NAND3_X1   g16401(.A1(new_n16180_), .A2(new_n16731_), .A3(new_n16427_), .ZN(new_n16732_));
  NAND3_X1   g16402(.A1(new_n16732_), .A2(new_n16730_), .A3(new_n16559_), .ZN(new_n16733_));
  AOI21_X1   g16403(.A1(new_n16725_), .A2(new_n16655_), .B(new_n16659_), .ZN(new_n16734_));
  AOI21_X1   g16404(.A1(new_n16660_), .A2(new_n16726_), .B(new_n16734_), .ZN(new_n16735_));
  NAND4_X1   g16405(.A1(new_n16733_), .A2(new_n16499_), .A3(new_n16558_), .A4(new_n16735_), .ZN(new_n16736_));
  OAI21_X1   g16406(.A1(new_n16667_), .A2(new_n16717_), .B(new_n16719_), .ZN(new_n16737_));
  INV_X1     g16407(.I(new_n16737_), .ZN(new_n16738_));
  INV_X1     g16408(.I(new_n16691_), .ZN(new_n16739_));
  AOI21_X1   g16409(.A1(new_n16675_), .A2(new_n16739_), .B(new_n16690_), .ZN(new_n16740_));
  INV_X1     g16410(.I(new_n16740_), .ZN(new_n16741_));
  NAND2_X1   g16411(.A1(\a[52] ), .A2(\a[60] ), .ZN(new_n16742_));
  NAND2_X1   g16412(.A1(\a[53] ), .A2(\a[61] ), .ZN(new_n16743_));
  XOR2_X1    g16413(.A1(new_n16742_), .A2(new_n16743_), .Z(new_n16744_));
  XOR2_X1    g16414(.A1(new_n16679_), .A2(new_n16744_), .Z(new_n16745_));
  AOI21_X1   g16415(.A1(new_n16694_), .A2(new_n16697_), .B(new_n15885_), .ZN(new_n16746_));
  NOR2_X1    g16416(.A1(new_n16746_), .A2(new_n16698_), .ZN(new_n16747_));
  XOR2_X1    g16417(.A1(new_n16745_), .A2(new_n16747_), .Z(new_n16748_));
  NAND2_X1   g16418(.A1(new_n16741_), .A2(new_n16748_), .ZN(new_n16749_));
  OR2_X2     g16419(.A1(new_n16745_), .A2(new_n16747_), .Z(new_n16750_));
  NAND2_X1   g16420(.A1(new_n16745_), .A2(new_n16747_), .ZN(new_n16751_));
  NAND2_X1   g16421(.A1(new_n16750_), .A2(new_n16751_), .ZN(new_n16752_));
  NAND2_X1   g16422(.A1(new_n16740_), .A2(new_n16752_), .ZN(new_n16753_));
  NAND2_X1   g16423(.A1(new_n16749_), .A2(new_n16753_), .ZN(new_n16754_));
  INV_X1     g16424(.I(new_n16754_), .ZN(new_n16755_));
  INV_X1     g16425(.I(new_n16708_), .ZN(new_n16756_));
  AOI21_X1   g16426(.A1(new_n16700_), .A2(new_n16756_), .B(new_n16707_), .ZN(new_n16757_));
  NAND2_X1   g16427(.A1(new_n6777_), .A2(new_n8991_), .ZN(new_n16758_));
  INV_X1     g16428(.I(new_n16758_), .ZN(new_n16759_));
  NAND2_X1   g16429(.A1(new_n7483_), .A2(new_n8676_), .ZN(new_n16760_));
  NOR2_X1    g16430(.A1(new_n6055_), .A2(new_n9310_), .ZN(new_n16761_));
  XOR2_X1    g16431(.A1(new_n16760_), .A2(new_n16761_), .Z(new_n16762_));
  XNOR2_X1   g16432(.A1(new_n13450_), .A2(new_n16695_), .ZN(new_n16763_));
  XNOR2_X1   g16433(.A1(new_n16762_), .A2(new_n16763_), .ZN(new_n16764_));
  NOR2_X1    g16434(.A1(new_n16764_), .A2(new_n16759_), .ZN(new_n16765_));
  NOR2_X1    g16435(.A1(new_n16762_), .A2(new_n16763_), .ZN(new_n16766_));
  INV_X1     g16436(.I(new_n16766_), .ZN(new_n16767_));
  NAND2_X1   g16437(.A1(new_n16762_), .A2(new_n16763_), .ZN(new_n16768_));
  AOI21_X1   g16438(.A1(new_n16767_), .A2(new_n16768_), .B(new_n16758_), .ZN(new_n16769_));
  NOR2_X1    g16439(.A1(new_n16765_), .A2(new_n16769_), .ZN(new_n16770_));
  INV_X1     g16440(.I(new_n16770_), .ZN(new_n16771_));
  AND2_X2    g16441(.A1(new_n16757_), .A2(new_n16771_), .Z(new_n16772_));
  NOR2_X1    g16442(.A1(new_n16757_), .A2(new_n16771_), .ZN(new_n16773_));
  NOR2_X1    g16443(.A1(new_n16772_), .A2(new_n16773_), .ZN(new_n16774_));
  NOR2_X1    g16444(.A1(new_n16755_), .A2(new_n16774_), .ZN(new_n16775_));
  XOR2_X1    g16445(.A1(new_n16757_), .A2(new_n16770_), .Z(new_n16776_));
  NOR2_X1    g16446(.A1(new_n16754_), .A2(new_n16776_), .ZN(new_n16777_));
  NOR2_X1    g16447(.A1(new_n16775_), .A2(new_n16777_), .ZN(new_n16778_));
  NOR2_X1    g16448(.A1(new_n16778_), .A2(new_n16738_), .ZN(new_n16779_));
  XOR2_X1    g16449(.A1(new_n16736_), .A2(new_n16779_), .Z(new_n16780_));
  XOR2_X1    g16450(.A1(new_n16780_), .A2(new_n16727_), .Z(\asquared[114] ));
  INV_X1     g16451(.I(new_n16779_), .ZN(new_n16782_));
  AOI21_X1   g16452(.A1(new_n16738_), .A2(new_n16778_), .B(new_n16727_), .ZN(new_n16783_));
  INV_X1     g16453(.I(new_n16783_), .ZN(new_n16784_));
  OAI21_X1   g16454(.A1(new_n16736_), .A2(new_n16784_), .B(new_n16782_), .ZN(new_n16785_));
  INV_X1     g16455(.I(new_n16772_), .ZN(new_n16786_));
  AOI21_X1   g16456(.A1(new_n16755_), .A2(new_n16786_), .B(new_n16773_), .ZN(new_n16787_));
  NAND2_X1   g16457(.A1(new_n16741_), .A2(new_n16751_), .ZN(new_n16788_));
  OAI22_X1   g16458(.A1(new_n7422_), .A2(new_n8005_), .B1(new_n9553_), .B2(new_n9555_), .ZN(new_n16789_));
  OAI21_X1   g16459(.A1(new_n8677_), .A2(new_n8953_), .B(new_n16789_), .ZN(new_n16790_));
  OAI21_X1   g16460(.A1(new_n16790_), .A2(new_n8244_), .B(new_n8085_), .ZN(new_n16791_));
  NAND2_X1   g16461(.A1(new_n16791_), .A2(\a[55] ), .ZN(new_n16792_));
  NAND3_X1   g16462(.A1(new_n16792_), .A2(new_n6945_), .A3(new_n8990_), .ZN(new_n16793_));
  AOI21_X1   g16463(.A1(new_n8676_), .A2(new_n8755_), .B(new_n16789_), .ZN(new_n16794_));
  NAND2_X1   g16464(.A1(new_n16793_), .A2(new_n16794_), .ZN(new_n16795_));
  NAND2_X1   g16465(.A1(new_n16768_), .A2(new_n16758_), .ZN(new_n16796_));
  NAND2_X1   g16466(.A1(new_n16796_), .A2(new_n16767_), .ZN(new_n16797_));
  AOI22_X1   g16467(.A1(new_n6777_), .A2(new_n9781_), .B1(new_n7000_), .B2(new_n9549_), .ZN(new_n16798_));
  NAND4_X1   g16468(.A1(new_n16798_), .A2(new_n8056_), .A3(new_n9785_), .A4(new_n13079_), .ZN(new_n16799_));
  XOR2_X1    g16469(.A1(new_n16797_), .A2(new_n16799_), .Z(new_n16800_));
  AOI21_X1   g16470(.A1(new_n16796_), .A2(new_n16767_), .B(new_n16799_), .ZN(new_n16801_));
  INV_X1     g16471(.I(new_n16799_), .ZN(new_n16802_));
  NOR2_X1    g16472(.A1(new_n16797_), .A2(new_n16802_), .ZN(new_n16803_));
  OAI21_X1   g16473(.A1(new_n16801_), .A2(new_n16803_), .B(new_n16795_), .ZN(new_n16804_));
  OAI21_X1   g16474(.A1(new_n16795_), .A2(new_n16800_), .B(new_n16804_), .ZN(new_n16805_));
  AOI22_X1   g16475(.A1(new_n16679_), .A2(new_n7204_), .B1(new_n16744_), .B2(new_n8991_), .ZN(new_n16806_));
  INV_X1     g16476(.I(new_n16806_), .ZN(new_n16807_));
  NOR2_X1    g16477(.A1(new_n7483_), .A2(new_n8676_), .ZN(new_n16808_));
  NAND2_X1   g16478(.A1(new_n6055_), .A2(new_n9310_), .ZN(new_n16809_));
  AOI21_X1   g16479(.A1(new_n7483_), .A2(new_n8676_), .B(new_n16809_), .ZN(new_n16810_));
  NOR2_X1    g16480(.A1(new_n16810_), .A2(new_n16808_), .ZN(new_n16811_));
  AOI21_X1   g16481(.A1(new_n8243_), .A2(new_n9029_), .B(new_n6260_), .ZN(new_n16812_));
  XNOR2_X1   g16482(.A1(new_n16811_), .A2(new_n16812_), .ZN(new_n16813_));
  INV_X1     g16483(.I(new_n16813_), .ZN(new_n16814_));
  INV_X1     g16484(.I(new_n16811_), .ZN(new_n16815_));
  INV_X1     g16485(.I(new_n16812_), .ZN(new_n16816_));
  NOR2_X1    g16486(.A1(new_n16815_), .A2(new_n16816_), .ZN(new_n16817_));
  NOR2_X1    g16487(.A1(new_n16811_), .A2(new_n16812_), .ZN(new_n16818_));
  NOR2_X1    g16488(.A1(new_n16817_), .A2(new_n16818_), .ZN(new_n16819_));
  NOR2_X1    g16489(.A1(new_n16807_), .A2(new_n16819_), .ZN(new_n16820_));
  AOI21_X1   g16490(.A1(new_n16807_), .A2(new_n16814_), .B(new_n16820_), .ZN(new_n16821_));
  XOR2_X1    g16491(.A1(new_n16805_), .A2(new_n16821_), .Z(new_n16822_));
  AOI21_X1   g16492(.A1(new_n16788_), .A2(new_n16750_), .B(new_n16822_), .ZN(new_n16823_));
  NAND2_X1   g16493(.A1(new_n16788_), .A2(new_n16750_), .ZN(new_n16824_));
  INV_X1     g16494(.I(new_n16821_), .ZN(new_n16825_));
  NAND2_X1   g16495(.A1(new_n16805_), .A2(new_n16825_), .ZN(new_n16826_));
  NOR2_X1    g16496(.A1(new_n16805_), .A2(new_n16825_), .ZN(new_n16827_));
  INV_X1     g16497(.I(new_n16827_), .ZN(new_n16828_));
  AOI21_X1   g16498(.A1(new_n16828_), .A2(new_n16826_), .B(new_n16824_), .ZN(new_n16829_));
  NOR2_X1    g16499(.A1(new_n16829_), .A2(new_n16823_), .ZN(new_n16830_));
  XNOR2_X1   g16500(.A1(new_n16830_), .A2(new_n16787_), .ZN(new_n16831_));
  INV_X1     g16501(.I(new_n16830_), .ZN(new_n16832_));
  NAND2_X1   g16502(.A1(new_n16832_), .A2(new_n16787_), .ZN(new_n16833_));
  INV_X1     g16503(.I(new_n16787_), .ZN(new_n16834_));
  NAND2_X1   g16504(.A1(new_n16834_), .A2(new_n16830_), .ZN(new_n16835_));
  NAND2_X1   g16505(.A1(new_n16833_), .A2(new_n16835_), .ZN(new_n16836_));
  MUX2_X1    g16506(.I0(new_n16836_), .I1(new_n16831_), .S(new_n16785_), .Z(\asquared[115] ));
  NAND2_X1   g16507(.A1(new_n16785_), .A2(new_n16833_), .ZN(new_n16838_));
  NAND2_X1   g16508(.A1(new_n16838_), .A2(new_n16835_), .ZN(new_n16839_));
  AOI21_X1   g16509(.A1(new_n16824_), .A2(new_n16826_), .B(new_n16827_), .ZN(new_n16840_));
  INV_X1     g16510(.I(new_n16817_), .ZN(new_n16841_));
  OAI21_X1   g16511(.A1(new_n16806_), .A2(new_n16818_), .B(new_n16841_), .ZN(new_n16842_));
  AOI22_X1   g16512(.A1(new_n7421_), .A2(new_n8991_), .B1(new_n7483_), .B2(new_n8455_), .ZN(new_n16843_));
  NOR4_X1    g16513(.A1(new_n8755_), .A2(new_n8996_), .A3(new_n6945_), .A4(new_n8453_), .ZN(new_n16844_));
  NAND2_X1   g16514(.A1(new_n16843_), .A2(new_n16844_), .ZN(new_n16845_));
  NAND2_X1   g16515(.A1(\a[57] ), .A2(\a[62] ), .ZN(new_n16846_));
  XOR2_X1    g16516(.A1(new_n16634_), .A2(new_n16846_), .Z(new_n16847_));
  XNOR2_X1   g16517(.A1(new_n16845_), .A2(new_n16847_), .ZN(new_n16848_));
  INV_X1     g16518(.I(new_n16848_), .ZN(new_n16849_));
  NOR2_X1    g16519(.A1(new_n16845_), .A2(new_n16847_), .ZN(new_n16850_));
  NAND2_X1   g16520(.A1(new_n16845_), .A2(new_n16847_), .ZN(new_n16851_));
  INV_X1     g16521(.I(new_n16851_), .ZN(new_n16852_));
  NOR2_X1    g16522(.A1(new_n16852_), .A2(new_n16850_), .ZN(new_n16853_));
  NOR2_X1    g16523(.A1(new_n16842_), .A2(new_n16853_), .ZN(new_n16854_));
  AOI21_X1   g16524(.A1(new_n16842_), .A2(new_n16849_), .B(new_n16854_), .ZN(new_n16855_));
  NOR2_X1    g16525(.A1(new_n16795_), .A2(new_n16803_), .ZN(new_n16856_));
  NOR2_X1    g16526(.A1(new_n16856_), .A2(new_n16801_), .ZN(new_n16857_));
  INV_X1     g16527(.I(new_n16798_), .ZN(new_n16858_));
  OAI21_X1   g16528(.A1(new_n8056_), .A2(new_n9785_), .B(new_n16858_), .ZN(new_n16859_));
  NOR2_X1    g16529(.A1(new_n16859_), .A2(new_n16790_), .ZN(new_n16860_));
  XOR2_X1    g16530(.A1(new_n16860_), .A2(new_n6692_), .Z(new_n16861_));
  XOR2_X1    g16531(.A1(new_n16861_), .A2(\a[63] ), .Z(new_n16862_));
  XNOR2_X1   g16532(.A1(new_n16857_), .A2(new_n16862_), .ZN(new_n16863_));
  NOR2_X1    g16533(.A1(new_n16863_), .A2(new_n16855_), .ZN(new_n16864_));
  INV_X1     g16534(.I(new_n16855_), .ZN(new_n16865_));
  XOR2_X1    g16535(.A1(new_n16857_), .A2(new_n16862_), .Z(new_n16866_));
  NOR2_X1    g16536(.A1(new_n16866_), .A2(new_n16865_), .ZN(new_n16867_));
  NOR2_X1    g16537(.A1(new_n16864_), .A2(new_n16867_), .ZN(new_n16868_));
  XNOR2_X1   g16538(.A1(new_n16840_), .A2(new_n16868_), .ZN(new_n16869_));
  NAND2_X1   g16539(.A1(new_n16839_), .A2(new_n16869_), .ZN(new_n16870_));
  INV_X1     g16540(.I(new_n16840_), .ZN(new_n16871_));
  NOR2_X1    g16541(.A1(new_n16871_), .A2(new_n16868_), .ZN(new_n16872_));
  NOR3_X1    g16542(.A1(new_n16840_), .A2(new_n16864_), .A3(new_n16867_), .ZN(new_n16873_));
  NOR2_X1    g16543(.A1(new_n16872_), .A2(new_n16873_), .ZN(new_n16874_));
  OAI21_X1   g16544(.A1(new_n16839_), .A2(new_n16874_), .B(new_n16870_), .ZN(\asquared[116] ));
  NAND4_X1   g16545(.A1(new_n16560_), .A2(new_n16558_), .A3(new_n16735_), .A4(new_n16783_), .ZN(new_n16876_));
  NOR2_X1    g16546(.A1(new_n16832_), .A2(new_n16873_), .ZN(new_n16877_));
  AOI21_X1   g16547(.A1(new_n16832_), .A2(new_n16873_), .B(new_n16834_), .ZN(new_n16878_));
  NOR2_X1    g16548(.A1(new_n16878_), .A2(new_n16877_), .ZN(new_n16879_));
  INV_X1     g16549(.I(new_n16879_), .ZN(new_n16880_));
  AOI21_X1   g16550(.A1(new_n16876_), .A2(new_n16782_), .B(new_n16880_), .ZN(new_n16881_));
  AND2_X2    g16551(.A1(new_n16881_), .A2(new_n16872_), .Z(\asquared[117] ));
  NAND2_X1   g16552(.A1(\a[53] ), .A2(\a[62] ), .ZN(new_n16883_));
  NOR2_X1    g16553(.A1(new_n6945_), .A2(new_n9310_), .ZN(new_n16884_));
  XOR2_X1    g16554(.A1(new_n16884_), .A2(new_n16883_), .Z(new_n16885_));
  AOI21_X1   g16555(.A1(new_n8755_), .A2(new_n8996_), .B(new_n16843_), .ZN(new_n16886_));
  AOI22_X1   g16556(.A1(new_n8455_), .A2(new_n8755_), .B1(new_n8991_), .B2(new_n10958_), .ZN(new_n16887_));
  NAND2_X1   g16557(.A1(new_n8242_), .A2(new_n8996_), .ZN(new_n16888_));
  AOI21_X1   g16558(.A1(new_n8242_), .A2(new_n8996_), .B(new_n16887_), .ZN(new_n16889_));
  AOI21_X1   g16559(.A1(new_n16889_), .A2(new_n8674_), .B(\a[60] ), .ZN(new_n16890_));
  NOR2_X1    g16560(.A1(\a[55] ), .A2(\a[61] ), .ZN(new_n16891_));
  OAI21_X1   g16561(.A1(new_n16890_), .A2(new_n7216_), .B(new_n16891_), .ZN(new_n16892_));
  NAND3_X1   g16562(.A1(new_n16892_), .A2(new_n16887_), .A3(new_n16888_), .ZN(new_n16893_));
  AOI21_X1   g16563(.A1(new_n8246_), .A2(new_n9029_), .B(new_n6694_), .ZN(new_n16894_));
  XOR2_X1    g16564(.A1(new_n16893_), .A2(new_n16894_), .Z(new_n16895_));
  XOR2_X1    g16565(.A1(new_n16895_), .A2(new_n16886_), .Z(new_n16896_));
  XOR2_X1    g16566(.A1(new_n16896_), .A2(new_n16885_), .Z(new_n16897_));
  NAND2_X1   g16567(.A1(\a[52] ), .A2(\a[63] ), .ZN(new_n16898_));
  AOI21_X1   g16568(.A1(new_n16859_), .A2(new_n16790_), .B(new_n16898_), .ZN(new_n16899_));
  NOR2_X1    g16569(.A1(new_n16899_), .A2(new_n16860_), .ZN(new_n16900_));
  NOR2_X1    g16570(.A1(new_n16897_), .A2(new_n16900_), .ZN(new_n16901_));
  AOI21_X1   g16571(.A1(new_n16842_), .A2(new_n16851_), .B(new_n16850_), .ZN(new_n16902_));
  AOI21_X1   g16572(.A1(new_n16897_), .A2(new_n16900_), .B(new_n16902_), .ZN(new_n16903_));
  NOR2_X1    g16573(.A1(new_n16903_), .A2(new_n16901_), .ZN(new_n16904_));
  INV_X1     g16574(.I(new_n16886_), .ZN(new_n16905_));
  NOR2_X1    g16575(.A1(new_n16893_), .A2(new_n16905_), .ZN(new_n16906_));
  XOR2_X1    g16576(.A1(new_n16885_), .A2(new_n16894_), .Z(new_n16907_));
  AOI21_X1   g16577(.A1(new_n16893_), .A2(new_n16905_), .B(new_n16907_), .ZN(new_n16908_));
  NOR2_X1    g16578(.A1(new_n16908_), .A2(new_n16906_), .ZN(new_n16909_));
  INV_X1     g16579(.I(new_n16909_), .ZN(new_n16910_));
  INV_X1     g16580(.I(new_n16885_), .ZN(new_n16911_));
  NOR2_X1    g16581(.A1(new_n16911_), .A2(new_n16894_), .ZN(new_n16912_));
  NOR2_X1    g16582(.A1(new_n10288_), .A2(new_n9550_), .ZN(new_n16913_));
  INV_X1     g16583(.I(new_n16913_), .ZN(new_n16914_));
  INV_X1     g16584(.I(new_n16889_), .ZN(new_n16915_));
  AOI22_X1   g16585(.A1(new_n7421_), .A2(new_n12964_), .B1(new_n9781_), .B2(new_n11018_), .ZN(new_n16916_));
  NAND4_X1   g16586(.A1(new_n16916_), .A2(new_n8243_), .A3(new_n8992_), .A4(new_n16884_), .ZN(new_n16917_));
  NOR2_X1    g16587(.A1(new_n16915_), .A2(new_n16917_), .ZN(new_n16918_));
  XOR2_X1    g16588(.A1(new_n16918_), .A2(new_n16914_), .Z(new_n16919_));
  XOR2_X1    g16589(.A1(new_n16919_), .A2(new_n16912_), .Z(new_n16920_));
  NAND2_X1   g16590(.A1(\a[58] ), .A2(\a[62] ), .ZN(new_n16921_));
  XOR2_X1    g16591(.A1(new_n15664_), .A2(new_n16921_), .Z(new_n16922_));
  NOR2_X1    g16592(.A1(new_n16920_), .A2(new_n16922_), .ZN(new_n16923_));
  NAND2_X1   g16593(.A1(new_n16920_), .A2(new_n16922_), .ZN(new_n16924_));
  INV_X1     g16594(.I(new_n16924_), .ZN(new_n16925_));
  OAI21_X1   g16595(.A1(new_n16925_), .A2(new_n16923_), .B(new_n16910_), .ZN(new_n16926_));
  XNOR2_X1   g16596(.A1(new_n16920_), .A2(new_n16922_), .ZN(new_n16927_));
  OAI21_X1   g16597(.A1(new_n16927_), .A2(new_n16910_), .B(new_n16926_), .ZN(new_n16928_));
  INV_X1     g16598(.I(new_n16928_), .ZN(new_n16929_));
  XOR2_X1    g16599(.A1(new_n16904_), .A2(new_n16929_), .Z(new_n16930_));
  NAND2_X1   g16600(.A1(\asquared[117] ), .A2(new_n16930_), .ZN(new_n16931_));
  XOR2_X1    g16601(.A1(new_n16904_), .A2(new_n16929_), .Z(new_n16932_));
  OAI21_X1   g16602(.A1(\asquared[117] ), .A2(new_n16932_), .B(new_n16931_), .ZN(\asquared[118] ));
  NOR2_X1    g16603(.A1(new_n16904_), .A2(new_n16929_), .ZN(new_n16934_));
  NAND2_X1   g16604(.A1(new_n16904_), .A2(new_n16929_), .ZN(new_n16935_));
  AOI21_X1   g16605(.A1(\asquared[117] ), .A2(new_n16935_), .B(new_n16934_), .ZN(new_n16936_));
  NOR2_X1    g16606(.A1(new_n16925_), .A2(new_n16909_), .ZN(new_n16937_));
  NOR2_X1    g16607(.A1(new_n16937_), .A2(new_n16923_), .ZN(new_n16938_));
  AOI21_X1   g16608(.A1(new_n8242_), .A2(new_n8991_), .B(new_n16916_), .ZN(new_n16939_));
  INV_X1     g16609(.I(new_n16939_), .ZN(new_n16940_));
  NOR2_X1    g16610(.A1(new_n8676_), .A2(\a[62] ), .ZN(new_n16941_));
  OAI21_X1   g16611(.A1(new_n16940_), .A2(new_n16941_), .B(\a[55] ), .ZN(new_n16942_));
  XOR2_X1    g16612(.A1(new_n16942_), .A2(\a[63] ), .Z(new_n16943_));
  NOR2_X1    g16613(.A1(new_n16915_), .A2(new_n16914_), .ZN(new_n16944_));
  NOR2_X1    g16614(.A1(new_n16889_), .A2(new_n16913_), .ZN(new_n16945_));
  NOR4_X1    g16615(.A1(new_n16945_), .A2(new_n16911_), .A3(new_n16894_), .A4(new_n16917_), .ZN(new_n16946_));
  NOR2_X1    g16616(.A1(new_n16946_), .A2(new_n16944_), .ZN(new_n16947_));
  AOI22_X1   g16617(.A1(new_n8242_), .A2(new_n16695_), .B1(new_n9784_), .B2(new_n9554_), .ZN(new_n16948_));
  INV_X1     g16618(.I(new_n16948_), .ZN(new_n16949_));
  NOR2_X1    g16619(.A1(new_n8246_), .A2(new_n8992_), .ZN(new_n16950_));
  AOI21_X1   g16620(.A1(\a[57] ), .A2(\a[61] ), .B(new_n9554_), .ZN(new_n16951_));
  NOR4_X1    g16621(.A1(new_n16949_), .A2(new_n16696_), .A3(new_n16950_), .A4(new_n16951_), .ZN(new_n16952_));
  INV_X1     g16622(.I(new_n16952_), .ZN(new_n16953_));
  NOR2_X1    g16623(.A1(new_n16947_), .A2(new_n16953_), .ZN(new_n16954_));
  NOR3_X1    g16624(.A1(new_n16946_), .A2(new_n16944_), .A3(new_n16952_), .ZN(new_n16955_));
  NOR2_X1    g16625(.A1(new_n16954_), .A2(new_n16955_), .ZN(new_n16956_));
  NOR2_X1    g16626(.A1(new_n16956_), .A2(new_n16943_), .ZN(new_n16957_));
  INV_X1     g16627(.I(new_n16943_), .ZN(new_n16958_));
  XOR2_X1    g16628(.A1(new_n16947_), .A2(new_n16952_), .Z(new_n16959_));
  NOR2_X1    g16629(.A1(new_n16959_), .A2(new_n16958_), .ZN(new_n16960_));
  NOR2_X1    g16630(.A1(new_n16960_), .A2(new_n16957_), .ZN(new_n16961_));
  XOR2_X1    g16631(.A1(new_n16938_), .A2(new_n16961_), .Z(new_n16962_));
  NOR3_X1    g16632(.A1(new_n16937_), .A2(new_n16923_), .A3(new_n16961_), .ZN(new_n16963_));
  NOR3_X1    g16633(.A1(new_n16938_), .A2(new_n16957_), .A3(new_n16960_), .ZN(new_n16964_));
  OAI21_X1   g16634(.A1(new_n16963_), .A2(new_n16964_), .B(new_n16936_), .ZN(new_n16965_));
  OAI21_X1   g16635(.A1(new_n16936_), .A2(new_n16962_), .B(new_n16965_), .ZN(\asquared[119] ));
  NOR2_X1    g16636(.A1(new_n16964_), .A2(new_n16928_), .ZN(new_n16967_));
  NAND2_X1   g16637(.A1(new_n16964_), .A2(new_n16928_), .ZN(new_n16968_));
  AOI21_X1   g16638(.A1(new_n16904_), .A2(new_n16968_), .B(new_n16967_), .ZN(new_n16969_));
  NAND4_X1   g16639(.A1(new_n16785_), .A2(new_n16872_), .A3(new_n16879_), .A4(new_n16969_), .ZN(new_n16970_));
  NOR2_X1    g16640(.A1(new_n16950_), .A2(new_n16948_), .ZN(new_n16971_));
  XNOR2_X1   g16641(.A1(new_n8454_), .A2(new_n16365_), .ZN(new_n16972_));
  XNOR2_X1   g16642(.A1(new_n16971_), .A2(new_n16972_), .ZN(new_n16973_));
  AOI21_X1   g16643(.A1(new_n8677_), .A2(new_n9029_), .B(new_n6999_), .ZN(new_n16974_));
  INV_X1     g16644(.I(new_n16974_), .ZN(new_n16975_));
  NOR2_X1    g16645(.A1(new_n6999_), .A2(new_n9310_), .ZN(new_n16976_));
  OAI21_X1   g16646(.A1(new_n16939_), .A2(new_n16974_), .B(new_n16976_), .ZN(new_n16977_));
  OAI21_X1   g16647(.A1(new_n16940_), .A2(new_n16975_), .B(new_n16977_), .ZN(new_n16978_));
  NAND2_X1   g16648(.A1(\a[59] ), .A2(\a[62] ), .ZN(new_n16979_));
  XNOR2_X1   g16649(.A1(new_n12540_), .A2(new_n16979_), .ZN(new_n16980_));
  XOR2_X1    g16650(.A1(new_n16978_), .A2(new_n16980_), .Z(new_n16981_));
  NOR2_X1    g16651(.A1(new_n16981_), .A2(new_n16973_), .ZN(new_n16982_));
  INV_X1     g16652(.I(new_n16973_), .ZN(new_n16983_));
  INV_X1     g16653(.I(new_n16978_), .ZN(new_n16984_));
  NOR2_X1    g16654(.A1(new_n16984_), .A2(new_n16980_), .ZN(new_n16985_));
  INV_X1     g16655(.I(new_n16985_), .ZN(new_n16986_));
  NAND2_X1   g16656(.A1(new_n16984_), .A2(new_n16980_), .ZN(new_n16987_));
  AOI21_X1   g16657(.A1(new_n16986_), .A2(new_n16987_), .B(new_n16983_), .ZN(new_n16988_));
  NOR2_X1    g16658(.A1(new_n16988_), .A2(new_n16982_), .ZN(new_n16989_));
  INV_X1     g16659(.I(new_n16989_), .ZN(new_n16990_));
  NOR2_X1    g16660(.A1(new_n16958_), .A2(new_n16955_), .ZN(new_n16991_));
  NOR2_X1    g16661(.A1(new_n16991_), .A2(new_n16954_), .ZN(new_n16992_));
  INV_X1     g16662(.I(new_n16992_), .ZN(new_n16993_));
  NAND2_X1   g16663(.A1(new_n16990_), .A2(new_n16993_), .ZN(new_n16994_));
  XOR2_X1    g16664(.A1(new_n16970_), .A2(new_n16994_), .Z(new_n16995_));
  XOR2_X1    g16665(.A1(new_n16995_), .A2(new_n16963_), .Z(\asquared[120] ));
  NAND2_X1   g16666(.A1(new_n16963_), .A2(new_n16990_), .ZN(new_n16997_));
  OAI21_X1   g16667(.A1(new_n16963_), .A2(new_n16990_), .B(new_n16993_), .ZN(new_n16998_));
  OAI21_X1   g16668(.A1(new_n16970_), .A2(new_n16998_), .B(new_n16997_), .ZN(new_n16999_));
  AOI22_X1   g16669(.A1(new_n8245_), .A2(new_n9781_), .B1(new_n8674_), .B2(new_n9549_), .ZN(new_n17000_));
  NAND2_X1   g16670(.A1(new_n8676_), .A2(new_n9784_), .ZN(new_n17001_));
  AOI21_X1   g16671(.A1(new_n8676_), .A2(new_n9784_), .B(new_n17000_), .ZN(new_n17002_));
  AOI21_X1   g16672(.A1(new_n17002_), .A2(new_n8455_), .B(\a[62] ), .ZN(new_n17003_));
  NOR2_X1    g16673(.A1(\a[57] ), .A2(\a[63] ), .ZN(new_n17004_));
  OAI21_X1   g16674(.A1(new_n17003_), .A2(new_n7647_), .B(new_n17004_), .ZN(new_n17005_));
  INV_X1     g16675(.I(new_n16971_), .ZN(new_n17006_));
  OAI22_X1   g16676(.A1(new_n17006_), .A2(new_n8244_), .B1(new_n9861_), .B2(new_n16972_), .ZN(new_n17007_));
  AOI21_X1   g16677(.A1(\a[57] ), .A2(new_n9153_), .B(new_n8996_), .ZN(new_n17008_));
  XOR2_X1    g16678(.A1(new_n17007_), .A2(new_n17008_), .Z(new_n17009_));
  NAND4_X1   g16679(.A1(new_n17009_), .A2(new_n17000_), .A3(new_n17001_), .A4(new_n17005_), .ZN(new_n17010_));
  NAND3_X1   g16680(.A1(new_n17005_), .A2(new_n17000_), .A3(new_n17001_), .ZN(new_n17011_));
  NAND2_X1   g16681(.A1(new_n17007_), .A2(new_n17008_), .ZN(new_n17012_));
  INV_X1     g16682(.I(new_n17012_), .ZN(new_n17013_));
  NOR2_X1    g16683(.A1(new_n17007_), .A2(new_n17008_), .ZN(new_n17014_));
  OAI21_X1   g16684(.A1(new_n17013_), .A2(new_n17014_), .B(new_n17011_), .ZN(new_n17015_));
  NAND2_X1   g16685(.A1(new_n17010_), .A2(new_n17015_), .ZN(new_n17016_));
  AOI21_X1   g16686(.A1(new_n16983_), .A2(new_n16987_), .B(new_n16985_), .ZN(new_n17017_));
  XOR2_X1    g16687(.A1(new_n17016_), .A2(new_n17017_), .Z(new_n17018_));
  INV_X1     g16688(.I(new_n17016_), .ZN(new_n17019_));
  INV_X1     g16689(.I(new_n17017_), .ZN(new_n17020_));
  NAND2_X1   g16690(.A1(new_n17019_), .A2(new_n17020_), .ZN(new_n17021_));
  NAND2_X1   g16691(.A1(new_n17016_), .A2(new_n17017_), .ZN(new_n17022_));
  NAND2_X1   g16692(.A1(new_n17021_), .A2(new_n17022_), .ZN(new_n17023_));
  MUX2_X1    g16693(.I0(new_n17023_), .I1(new_n17018_), .S(new_n16999_), .Z(\asquared[121] ));
  NAND2_X1   g16694(.A1(new_n16999_), .A2(new_n17022_), .ZN(new_n17025_));
  NAND2_X1   g16695(.A1(new_n17025_), .A2(new_n17021_), .ZN(new_n17026_));
  OAI21_X1   g16696(.A1(new_n17011_), .A2(new_n17014_), .B(new_n17012_), .ZN(new_n17027_));
  INV_X1     g16697(.I(new_n17002_), .ZN(new_n17028_));
  XNOR2_X1   g16698(.A1(new_n8455_), .A2(new_n9153_), .ZN(new_n17029_));
  NOR2_X1    g16699(.A1(new_n17028_), .A2(new_n17029_), .ZN(new_n17030_));
  XOR2_X1    g16700(.A1(new_n17030_), .A2(new_n7647_), .Z(new_n17031_));
  XOR2_X1    g16701(.A1(new_n17031_), .A2(\a[63] ), .Z(new_n17032_));
  XOR2_X1    g16702(.A1(new_n17032_), .A2(new_n17027_), .Z(new_n17033_));
  NAND2_X1   g16703(.A1(new_n17026_), .A2(new_n17033_), .ZN(new_n17034_));
  NOR2_X1    g16704(.A1(new_n17032_), .A2(new_n17027_), .ZN(new_n17035_));
  NAND2_X1   g16705(.A1(new_n17032_), .A2(new_n17027_), .ZN(new_n17036_));
  INV_X1     g16706(.I(new_n17036_), .ZN(new_n17037_));
  NOR2_X1    g16707(.A1(new_n17037_), .A2(new_n17035_), .ZN(new_n17038_));
  OAI21_X1   g16708(.A1(new_n17026_), .A2(new_n17038_), .B(new_n17034_), .ZN(\asquared[122] ));
  INV_X1     g16709(.I(new_n16998_), .ZN(new_n17040_));
  NAND4_X1   g16710(.A1(new_n16881_), .A2(new_n16872_), .A3(new_n16969_), .A4(new_n17040_), .ZN(new_n17041_));
  AOI21_X1   g16711(.A1(new_n17037_), .A2(new_n17016_), .B(new_n17020_), .ZN(new_n17042_));
  AOI21_X1   g16712(.A1(new_n17019_), .A2(new_n17036_), .B(new_n17042_), .ZN(new_n17043_));
  INV_X1     g16713(.I(new_n17043_), .ZN(new_n17044_));
  AOI21_X1   g16714(.A1(new_n17041_), .A2(new_n16997_), .B(new_n17044_), .ZN(new_n17045_));
  INV_X1     g16715(.I(new_n16365_), .ZN(new_n17046_));
  AOI21_X1   g16716(.A1(new_n17028_), .A2(new_n17029_), .B(new_n17046_), .ZN(new_n17047_));
  NOR2_X1    g16717(.A1(new_n17047_), .A2(new_n17030_), .ZN(new_n17048_));
  AOI21_X1   g16718(.A1(\a[59] ), .A2(\a[63] ), .B(new_n9153_), .ZN(new_n17049_));
  AOI21_X1   g16719(.A1(new_n8992_), .A2(new_n9029_), .B(new_n8085_), .ZN(new_n17050_));
  OAI21_X1   g16720(.A1(new_n17050_), .A2(new_n17049_), .B(new_n9549_), .ZN(new_n17051_));
  XOR2_X1    g16721(.A1(new_n17051_), .A2(new_n8996_), .Z(new_n17052_));
  NOR2_X1    g16722(.A1(new_n17048_), .A2(new_n17052_), .ZN(new_n17053_));
  XOR2_X1    g16723(.A1(new_n17045_), .A2(new_n17053_), .Z(new_n17054_));
  XOR2_X1    g16724(.A1(new_n17054_), .A2(new_n17035_), .Z(\asquared[123] ));
  INV_X1     g16725(.I(new_n17048_), .ZN(new_n17056_));
  NOR2_X1    g16726(.A1(new_n17035_), .A2(new_n17056_), .ZN(new_n17057_));
  NOR2_X1    g16727(.A1(new_n17057_), .A2(new_n17052_), .ZN(new_n17058_));
  AOI22_X1   g16728(.A1(new_n17045_), .A2(new_n17058_), .B1(new_n17035_), .B2(new_n17056_), .ZN(new_n17059_));
  AOI22_X1   g16729(.A1(new_n17050_), .A2(new_n9549_), .B1(new_n8996_), .B2(new_n17049_), .ZN(new_n17060_));
  AOI21_X1   g16730(.A1(new_n8453_), .A2(\a[62] ), .B(new_n12892_), .ZN(new_n17061_));
  NOR3_X1    g16731(.A1(new_n11018_), .A2(\a[61] ), .A3(new_n9029_), .ZN(new_n17062_));
  NOR2_X1    g16732(.A1(new_n17061_), .A2(new_n17062_), .ZN(new_n17063_));
  XOR2_X1    g16733(.A1(new_n17060_), .A2(new_n17063_), .Z(new_n17064_));
  INV_X1     g16734(.I(new_n17060_), .ZN(new_n17065_));
  NOR2_X1    g16735(.A1(new_n17065_), .A2(new_n17063_), .ZN(new_n17066_));
  INV_X1     g16736(.I(new_n17063_), .ZN(new_n17067_));
  NOR2_X1    g16737(.A1(new_n17067_), .A2(new_n17060_), .ZN(new_n17068_));
  OAI21_X1   g16738(.A1(new_n17066_), .A2(new_n17068_), .B(new_n17059_), .ZN(new_n17069_));
  OAI21_X1   g16739(.A1(new_n17059_), .A2(new_n17064_), .B(new_n17069_), .ZN(\asquared[124] ));
  NAND2_X1   g16740(.A1(new_n9549_), .A2(new_n8990_), .ZN(new_n17071_));
  NAND2_X1   g16741(.A1(new_n9550_), .A2(\a[60] ), .ZN(new_n17072_));
  AOI21_X1   g16742(.A1(new_n17072_), .A2(new_n17071_), .B(new_n8453_), .ZN(new_n17073_));
  NOR2_X1    g16743(.A1(new_n17073_), .A2(new_n9153_), .ZN(new_n17074_));
  INV_X1     g16744(.I(new_n17074_), .ZN(new_n17075_));
  NOR2_X1    g16745(.A1(new_n17068_), .A2(new_n17075_), .ZN(new_n17076_));
  OAI21_X1   g16746(.A1(new_n17059_), .A2(new_n17066_), .B(new_n17076_), .ZN(new_n17077_));
  NAND3_X1   g16747(.A1(new_n17077_), .A2(\a[62] ), .A3(new_n9861_), .ZN(new_n17078_));
  NAND2_X1   g16748(.A1(new_n17077_), .A2(\a[62] ), .ZN(new_n17079_));
  NAND2_X1   g16749(.A1(new_n17079_), .A2(new_n9781_), .ZN(new_n17080_));
  NAND2_X1   g16750(.A1(new_n17080_), .A2(new_n17078_), .ZN(\asquared[125] ));
  NAND2_X1   g16751(.A1(new_n17035_), .A2(new_n17056_), .ZN(new_n17082_));
  NAND3_X1   g16752(.A1(new_n16999_), .A2(new_n17043_), .A3(new_n17058_), .ZN(new_n17083_));
  NAND2_X1   g16753(.A1(new_n17083_), .A2(new_n17082_), .ZN(new_n17084_));
  AOI21_X1   g16754(.A1(new_n17075_), .A2(new_n17067_), .B(new_n17065_), .ZN(new_n17085_));
  AOI21_X1   g16755(.A1(new_n17063_), .A2(new_n17074_), .B(new_n17085_), .ZN(new_n17086_));
  NAND3_X1   g16756(.A1(new_n17084_), .A2(new_n8453_), .A3(new_n17086_), .ZN(new_n17087_));
  NAND2_X1   g16757(.A1(new_n17087_), .A2(new_n9310_), .ZN(new_n17088_));
  NAND3_X1   g16758(.A1(new_n17088_), .A2(new_n8453_), .A3(\a[62] ), .ZN(new_n17089_));
  OAI21_X1   g16759(.A1(new_n9029_), .A2(new_n9310_), .B(\a[61] ), .ZN(new_n17090_));
  NAND2_X1   g16760(.A1(new_n17089_), .A2(new_n17090_), .ZN(\asquared[126] ));
  NAND2_X1   g16761(.A1(new_n17084_), .A2(new_n17086_), .ZN(new_n17092_));
  AOI21_X1   g16762(.A1(new_n17092_), .A2(new_n8453_), .B(new_n9029_), .ZN(\asquared[127] ));
  assign     \asquared[1]  = 1'b1;
  BUF_X16    g16763(.I(\a[0] ), .Z(\asquared[0] ));
endmodule


