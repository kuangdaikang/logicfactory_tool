// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:57 2022

module in1  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    \v16.0 , \v16.1 , \v16.2 , \v16.3 , \v16.4 , \v16.5 , \v16.6 , \v16.7 ,
    \v16.8 , \v16.9 , \v16.10 , \v16.11 , \v16.12 , \v16.13 , \v16.14 ,
    \v16.15 , \v16.16   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15;
  output \v16.0 , \v16.1 , \v16.2 , \v16.3 , \v16.4 , \v16.5 , \v16.6 ,
    \v16.7 , \v16.8 , \v16.9 , \v16.10 , \v16.11 , \v16.12 , \v16.13 ,
    \v16.14 , \v16.15 , \v16.16 ;
  wire new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_,
    new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_,
    new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_;
  assign new_n34_ = ~v1 & v15;
  assign new_n35_ = ~v14 & ~v15;
  assign new_n36_ = ~new_n34_ & ~new_n35_;
  assign new_n37_ = v0 & ~new_n36_;
  assign new_n38_ = ~v14 & v15;
  assign new_n39_ = ~v0 & new_n38_;
  assign new_n40_ = ~v14 & ~new_n39_;
  assign new_n41_ = ~new_n37_ & new_n40_;
  assign new_n42_ = v12 & ~new_n41_;
  assign new_n43_ = v0 & v15;
  assign new_n44_ = ~v8 & v9;
  assign new_n45_ = ~v8 & ~new_n44_;
  assign new_n46_ = ~new_n43_ & ~new_n45_;
  assign new_n47_ = ~v14 & new_n46_;
  assign new_n48_ = v7 & new_n47_;
  assign new_n49_ = ~v6 & new_n48_;
  assign new_n50_ = ~v5 & new_n49_;
  assign new_n51_ = v4 & new_n50_;
  assign new_n52_ = ~v0 & v14;
  assign new_n53_ = ~new_n51_ & ~new_n52_;
  assign new_n54_ = ~v12 & ~new_n53_;
  assign new_n55_ = ~new_n42_ & ~new_n54_;
  assign new_n56_ = ~v11 & ~new_n55_;
  assign new_n57_ = v8 & ~v14;
  assign new_n58_ = v15 & ~new_n57_;
  assign new_n59_ = v6 & v7;
  assign new_n60_ = v0 & ~new_n59_;
  assign new_n61_ = ~new_n58_ & ~new_n60_;
  assign new_n62_ = ~v8 & v14;
  assign new_n63_ = ~v6 & ~new_n62_;
  assign new_n64_ = ~v0 & new_n63_;
  assign new_n65_ = ~new_n61_ & ~new_n64_;
  assign new_n66_ = v5 & ~new_n65_;
  assign new_n67_ = ~v8 & ~v9;
  assign new_n68_ = ~v7 & ~new_n67_;
  assign new_n69_ = ~v8 & ~v14;
  assign new_n70_ = v7 & new_n69_;
  assign new_n71_ = ~new_n68_ & ~new_n70_;
  assign new_n72_ = ~v15 & ~new_n71_;
  assign new_n73_ = ~v6 & new_n72_;
  assign new_n74_ = ~v0 & new_n73_;
  assign new_n75_ = ~new_n66_ & ~new_n74_;
  assign new_n76_ = ~v12 & ~new_n75_;
  assign new_n77_ = v7 & ~v9;
  assign new_n78_ = ~v9 & ~new_n77_;
  assign new_n79_ = ~v14 & ~new_n78_;
  assign new_n80_ = v12 & new_n79_;
  assign new_n81_ = ~v8 & new_n80_;
  assign new_n82_ = ~v6 & new_n81_;
  assign new_n83_ = ~v5 & new_n82_;
  assign new_n84_ = v4 & new_n83_;
  assign new_n85_ = ~v0 & new_n84_;
  assign new_n86_ = ~new_n76_ & ~new_n85_;
  assign new_n87_ = v11 & ~new_n86_;
  assign new_n88_ = ~new_n56_ & ~new_n87_;
  assign new_n89_ = v10 & ~new_n88_;
  assign new_n90_ = ~v7 & v12;
  assign new_n91_ = ~v1 & new_n90_;
  assign new_n92_ = ~v7 & ~new_n91_;
  assign new_n93_ = ~v1 & new_n92_;
  assign new_n94_ = v15 & ~new_n93_;
  assign new_n95_ = v6 & new_n94_;
  assign new_n96_ = ~v7 & v8;
  assign new_n97_ = v6 & ~new_n96_;
  assign new_n98_ = ~v15 & ~new_n97_;
  assign new_n99_ = ~v12 & new_n98_;
  assign new_n100_ = ~new_n95_ & ~new_n99_;
  assign new_n101_ = ~v14 & ~new_n100_;
  assign new_n102_ = v14 & v15;
  assign new_n103_ = v8 & ~v15;
  assign new_n104_ = v1 & new_n103_;
  assign new_n105_ = ~new_n102_ & ~new_n104_;
  assign new_n106_ = ~v6 & ~new_n105_;
  assign new_n107_ = new_n96_ & new_n102_;
  assign new_n108_ = ~new_n106_ & ~new_n107_;
  assign new_n109_ = ~v12 & ~new_n108_;
  assign new_n110_ = ~new_n101_ & ~new_n109_;
  assign new_n111_ = ~v0 & ~new_n110_;
  assign new_n112_ = ~new_n35_ & ~new_n102_;
  assign new_n113_ = ~v12 & ~new_n112_;
  assign new_n114_ = v8 & new_n113_;
  assign new_n115_ = v7 & new_n114_;
  assign new_n116_ = v6 & new_n115_;
  assign new_n117_ = ~new_n111_ & ~new_n116_;
  assign new_n118_ = v5 & ~new_n117_;
  assign new_n119_ = ~v5 & ~v6;
  assign new_n120_ = new_n96_ & new_n119_;
  assign new_n121_ = v9 & v12;
  assign new_n122_ = new_n35_ & new_n121_;
  assign new_n123_ = new_n120_ & new_n122_;
  assign new_n124_ = ~new_n118_ & ~new_n123_;
  assign new_n125_ = v11 & ~new_n124_;
  assign new_n126_ = ~v6 & v15;
  assign new_n127_ = v15 & ~new_n126_;
  assign new_n128_ = ~v14 & ~new_n127_;
  assign new_n129_ = ~v14 & ~new_n128_;
  assign new_n130_ = v12 & ~new_n129_;
  assign new_n131_ = ~v11 & new_n130_;
  assign new_n132_ = ~new_n125_ & ~new_n131_;
  assign new_n133_ = v4 & ~new_n132_;
  assign new_n134_ = ~v5 & ~v14;
  assign new_n135_ = ~v12 & ~new_n134_;
  assign new_n136_ = ~v11 & ~new_n135_;
  assign new_n137_ = ~v4 & new_n136_;
  assign new_n138_ = ~new_n133_ & ~new_n137_;
  assign new_n139_ = ~v10 & ~new_n138_;
  assign new_n140_ = ~new_n89_ & ~new_n139_;
  assign new_n141_ = ~v13 & ~new_n140_;
  assign new_n142_ = ~v1 & ~v7;
  assign new_n143_ = v11 & ~new_n142_;
  assign new_n144_ = ~v10 & new_n143_;
  assign new_n145_ = v6 & new_n144_;
  assign new_n146_ = v5 & new_n145_;
  assign new_n147_ = v4 & new_n146_;
  assign new_n148_ = ~v2 & new_n147_;
  assign new_n149_ = ~v0 & new_n148_;
  assign new_n150_ = v7 & v8;
  assign new_n151_ = ~v4 & new_n150_;
  assign new_n152_ = ~v11 & v15;
  assign new_n153_ = v10 & new_n152_;
  assign new_n154_ = new_n151_ & new_n153_;
  assign new_n155_ = ~new_n149_ & ~new_n154_;
  assign new_n156_ = ~v10 & v11;
  assign new_n157_ = ~v5 & new_n156_;
  assign new_n158_ = ~v6 & new_n44_;
  assign new_n159_ = v8 & ~v9;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_ = ~v7 & ~new_n160_;
  assign new_n162_ = v7 & ~v8;
  assign new_n163_ = ~new_n161_ & ~new_n162_;
  assign new_n164_ = ~v4 & ~new_n163_;
  assign new_n165_ = ~v4 & ~new_n164_;
  assign new_n166_ = v15 & ~new_n165_;
  assign new_n167_ = ~v11 & new_n166_;
  assign new_n168_ = v10 & new_n167_;
  assign new_n169_ = ~new_n157_ & ~new_n168_;
  assign new_n170_ = new_n155_ & new_n169_;
  assign new_n171_ = ~v14 & ~new_n170_;
  assign new_n172_ = v8 & new_n156_;
  assign new_n173_ = ~v6 & new_n172_;
  assign new_n174_ = v5 & new_n173_;
  assign new_n175_ = v4 & new_n174_;
  assign new_n176_ = v1 & new_n175_;
  assign new_n177_ = ~v0 & new_n176_;
  assign new_n178_ = v10 & ~v11;
  assign new_n179_ = ~new_n177_ & ~new_n178_;
  assign new_n180_ = ~v15 & ~new_n179_;
  assign new_n181_ = v14 & new_n180_;
  assign new_n182_ = ~new_n171_ & ~new_n181_;
  assign new_n183_ = v12 & ~new_n182_;
  assign new_n184_ = v4 & ~v5;
  assign new_n185_ = ~v6 & ~v7;
  assign new_n186_ = new_n184_ & new_n185_;
  assign new_n187_ = ~v9 & ~v10;
  assign new_n188_ = v11 & new_n38_;
  assign new_n189_ = new_n187_ & new_n188_;
  assign new_n190_ = new_n186_ & new_n189_;
  assign new_n191_ = v14 & ~v15;
  assign new_n192_ = new_n178_ & new_n191_;
  assign new_n193_ = ~new_n190_ & ~new_n192_;
  assign new_n194_ = v8 & ~new_n193_;
  assign new_n195_ = v9 & v11;
  assign new_n196_ = ~v8 & new_n195_;
  assign new_n197_ = ~v7 & new_n196_;
  assign new_n198_ = ~v6 & new_n197_;
  assign new_n199_ = ~v5 & new_n198_;
  assign new_n200_ = ~v10 & ~v11;
  assign new_n201_ = ~new_n199_ & ~new_n200_;
  assign new_n202_ = v15 & ~new_n201_;
  assign new_n203_ = ~v11 & ~v15;
  assign new_n204_ = ~v10 & new_n203_;
  assign new_n205_ = ~new_n202_ & ~new_n204_;
  assign new_n206_ = v14 & ~new_n205_;
  assign new_n207_ = ~v11 & ~v14;
  assign new_n208_ = ~v10 & new_n207_;
  assign new_n209_ = ~new_n206_ & ~new_n208_;
  assign new_n210_ = v4 & ~new_n209_;
  assign new_n211_ = v9 & v14;
  assign new_n212_ = new_n162_ & new_n211_;
  assign new_n213_ = v14 & ~new_n212_;
  assign new_n214_ = ~v11 & ~new_n213_;
  assign new_n215_ = v10 & new_n214_;
  assign new_n216_ = ~new_n210_ & ~new_n215_;
  assign new_n217_ = ~new_n194_ & new_n216_;
  assign new_n218_ = ~v12 & ~new_n217_;
  assign new_n219_ = new_n35_ & new_n178_;
  assign new_n220_ = ~new_n218_ & ~new_n219_;
  assign new_n221_ = ~new_n183_ & new_n220_;
  assign new_n222_ = v13 & ~new_n221_;
  assign new_n223_ = ~v4 & ~v10;
  assign new_n224_ = ~v12 & ~v15;
  assign new_n225_ = ~v11 & new_n224_;
  assign new_n226_ = new_n223_ & new_n225_;
  assign new_n227_ = ~new_n222_ & ~new_n226_;
  assign \v16.0  = new_n141_ | ~new_n227_;
  assign new_n229_ = v4 & v9;
  assign new_n230_ = v4 & ~new_n229_;
  assign new_n231_ = v15 & ~new_n142_;
  assign new_n232_ = ~v10 & new_n231_;
  assign new_n233_ = v6 & new_n232_;
  assign new_n234_ = v5 & new_n233_;
  assign new_n235_ = ~v6 & v7;
  assign new_n236_ = ~v5 & new_n235_;
  assign new_n237_ = v10 & v12;
  assign new_n238_ = ~v8 & new_n237_;
  assign new_n239_ = new_n236_ & new_n238_;
  assign new_n240_ = ~new_n234_ & ~new_n239_;
  assign new_n241_ = v11 & ~new_n240_;
  assign new_n242_ = v8 & v10;
  assign new_n243_ = ~v11 & ~v12;
  assign new_n244_ = new_n242_ & new_n243_;
  assign new_n245_ = new_n236_ & new_n244_;
  assign new_n246_ = ~new_n241_ & ~new_n245_;
  assign new_n247_ = ~v0 & ~new_n246_;
  assign new_n248_ = new_n119_ & new_n150_;
  assign new_n249_ = new_n178_ & new_n224_;
  assign new_n250_ = new_n248_ & new_n249_;
  assign new_n251_ = ~new_n247_ & ~new_n250_;
  assign new_n252_ = ~new_n230_ & ~new_n251_;
  assign new_n253_ = ~v1 & v4;
  assign new_n254_ = ~v7 & v9;
  assign new_n255_ = new_n253_ & new_n254_;
  assign new_n256_ = v4 & ~new_n255_;
  assign new_n257_ = v11 & ~new_n256_;
  assign new_n258_ = v5 & new_n257_;
  assign new_n259_ = ~v0 & new_n258_;
  assign new_n260_ = v1 & ~v4;
  assign new_n261_ = ~v11 & ~new_n260_;
  assign new_n262_ = ~new_n259_ & ~new_n261_;
  assign new_n263_ = v6 & ~new_n262_;
  assign new_n264_ = ~v6 & ~v11;
  assign new_n265_ = v4 & new_n264_;
  assign new_n266_ = ~new_n263_ & ~new_n265_;
  assign new_n267_ = v15 & ~new_n266_;
  assign new_n268_ = ~v5 & new_n185_;
  assign new_n269_ = v8 & new_n195_;
  assign new_n270_ = new_n268_ & new_n269_;
  assign new_n271_ = v11 & ~new_n270_;
  assign new_n272_ = v4 & ~new_n271_;
  assign new_n273_ = ~v4 & new_n119_;
  assign new_n274_ = new_n96_ & new_n195_;
  assign new_n275_ = new_n273_ & new_n274_;
  assign new_n276_ = ~new_n272_ & ~new_n275_;
  assign new_n277_ = ~v15 & ~new_n276_;
  assign new_n278_ = ~new_n267_ & ~new_n277_;
  assign new_n279_ = ~v10 & ~new_n278_;
  assign new_n280_ = ~new_n77_ & ~new_n254_;
  assign new_n281_ = v4 & ~new_n280_;
  assign new_n282_ = ~v4 & v9;
  assign new_n283_ = ~new_n281_ & ~new_n282_;
  assign new_n284_ = v11 & ~new_n283_;
  assign new_n285_ = ~v8 & new_n284_;
  assign new_n286_ = ~v6 & new_n285_;
  assign new_n287_ = ~v5 & new_n286_;
  assign new_n288_ = ~new_n152_ & ~new_n287_;
  assign new_n289_ = ~v0 & ~new_n288_;
  assign new_n290_ = v0 & new_n203_;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = v10 & ~new_n291_;
  assign new_n293_ = ~new_n279_ & ~new_n292_;
  assign new_n294_ = v12 & ~new_n293_;
  assign new_n295_ = ~v10 & ~v15;
  assign new_n296_ = ~v4 & new_n295_;
  assign new_n297_ = ~v10 & ~new_n296_;
  assign new_n298_ = v6 & ~v8;
  assign new_n299_ = ~v0 & ~new_n298_;
  assign new_n300_ = v6 & new_n150_;
  assign new_n301_ = ~new_n299_ & ~new_n300_;
  assign new_n302_ = ~new_n297_ & ~new_n301_;
  assign new_n303_ = v5 & new_n302_;
  assign new_n304_ = ~v0 & new_n235_;
  assign new_n305_ = v10 & ~v15;
  assign new_n306_ = ~v8 & new_n305_;
  assign new_n307_ = new_n304_ & new_n306_;
  assign new_n308_ = ~new_n303_ & ~new_n307_;
  assign new_n309_ = v11 & ~new_n308_;
  assign new_n310_ = ~new_n44_ & ~new_n159_;
  assign new_n311_ = v4 & ~new_n310_;
  assign new_n312_ = ~new_n282_ & ~new_n311_;
  assign new_n313_ = ~new_n43_ & ~new_n312_;
  assign new_n314_ = ~v11 & new_n313_;
  assign new_n315_ = v10 & new_n314_;
  assign new_n316_ = v7 & new_n315_;
  assign new_n317_ = ~v6 & new_n316_;
  assign new_n318_ = ~v5 & new_n317_;
  assign new_n319_ = ~new_n309_ & ~new_n318_;
  assign new_n320_ = ~v12 & ~new_n319_;
  assign new_n321_ = ~v4 & ~v5;
  assign new_n322_ = new_n200_ & new_n321_;
  assign new_n323_ = ~new_n320_ & ~new_n322_;
  assign new_n324_ = ~new_n294_ & new_n323_;
  assign new_n325_ = ~new_n252_ & new_n324_;
  assign new_n326_ = ~v14 & ~new_n325_;
  assign new_n327_ = ~v12 & v14;
  assign new_n328_ = ~v10 & new_n327_;
  assign new_n329_ = v12 & v15;
  assign new_n330_ = v10 & new_n329_;
  assign new_n331_ = ~new_n328_ & ~new_n330_;
  assign new_n332_ = v0 & ~new_n331_;
  assign new_n333_ = ~v10 & ~v12;
  assign new_n334_ = new_n102_ & new_n333_;
  assign new_n335_ = ~new_n332_ & ~new_n334_;
  assign new_n336_ = ~v1 & ~new_n335_;
  assign new_n337_ = v4 & ~v10;
  assign new_n338_ = v10 & v14;
  assign new_n339_ = ~v0 & new_n338_;
  assign new_n340_ = ~new_n337_ & ~new_n339_;
  assign new_n341_ = ~v12 & ~new_n340_;
  assign new_n342_ = v4 & v14;
  assign new_n343_ = v4 & ~new_n342_;
  assign new_n344_ = v12 & ~new_n343_;
  assign new_n345_ = ~v10 & new_n344_;
  assign new_n346_ = ~new_n341_ & ~new_n345_;
  assign new_n347_ = ~new_n336_ & new_n346_;
  assign new_n348_ = ~v11 & ~new_n347_;
  assign new_n349_ = ~v4 & v8;
  assign new_n350_ = ~v10 & new_n102_;
  assign new_n351_ = new_n349_ & new_n350_;
  assign new_n352_ = ~new_n305_ & ~new_n351_;
  assign new_n353_ = ~new_n60_ & ~new_n352_;
  assign new_n354_ = new_n102_ & new_n223_;
  assign new_n355_ = ~new_n242_ & ~new_n354_;
  assign new_n356_ = ~v6 & ~new_n355_;
  assign new_n357_ = ~v0 & new_n356_;
  assign new_n358_ = ~new_n353_ & ~new_n357_;
  assign new_n359_ = v5 & ~new_n358_;
  assign new_n360_ = v10 & ~new_n67_;
  assign new_n361_ = ~v7 & new_n360_;
  assign new_n362_ = ~v6 & new_n361_;
  assign new_n363_ = ~v0 & new_n362_;
  assign new_n364_ = v1 & v4;
  assign new_n365_ = ~v6 & v8;
  assign new_n366_ = v5 & new_n365_;
  assign new_n367_ = new_n364_ & new_n366_;
  assign new_n368_ = v14 & ~new_n367_;
  assign new_n369_ = ~v10 & new_n368_;
  assign new_n370_ = ~new_n363_ & ~new_n369_;
  assign new_n371_ = ~v15 & ~new_n370_;
  assign new_n372_ = ~new_n359_ & ~new_n371_;
  assign new_n373_ = ~v12 & ~new_n372_;
  assign new_n374_ = v11 & new_n373_;
  assign new_n375_ = ~new_n348_ & ~new_n374_;
  assign new_n376_ = ~new_n326_ & new_n375_;
  assign new_n377_ = ~v13 & ~new_n376_;
  assign new_n378_ = ~new_n142_ & ~new_n230_;
  assign new_n379_ = v6 & new_n378_;
  assign new_n380_ = v5 & new_n379_;
  assign new_n381_ = ~v2 & new_n380_;
  assign new_n382_ = ~v0 & new_n381_;
  assign new_n383_ = v5 & ~new_n382_;
  assign new_n384_ = v11 & ~new_n383_;
  assign new_n385_ = ~v10 & new_n384_;
  assign new_n386_ = ~v7 & ~new_n161_;
  assign new_n387_ = ~v4 & ~new_n386_;
  assign new_n388_ = ~v4 & ~new_n387_;
  assign new_n389_ = v15 & ~new_n388_;
  assign new_n390_ = ~v11 & new_n389_;
  assign new_n391_ = v10 & new_n390_;
  assign new_n392_ = ~new_n385_ & ~new_n391_;
  assign new_n393_ = v12 & ~new_n392_;
  assign new_n394_ = ~v9 & v11;
  assign new_n395_ = v8 & new_n394_;
  assign new_n396_ = new_n268_ & new_n395_;
  assign new_n397_ = v11 & ~new_n396_;
  assign new_n398_ = v4 & ~new_n397_;
  assign new_n399_ = new_n96_ & new_n394_;
  assign new_n400_ = new_n273_ & new_n399_;
  assign new_n401_ = ~new_n398_ & ~new_n400_;
  assign new_n402_ = v15 & ~new_n401_;
  assign new_n403_ = v4 & new_n203_;
  assign new_n404_ = ~new_n402_ & ~new_n403_;
  assign new_n405_ = ~v10 & ~new_n404_;
  assign new_n406_ = ~new_n178_ & ~new_n405_;
  assign new_n407_ = ~v12 & ~new_n406_;
  assign new_n408_ = v10 & new_n203_;
  assign new_n409_ = ~new_n407_ & ~new_n408_;
  assign new_n410_ = ~new_n393_ & new_n409_;
  assign new_n411_ = ~v14 & ~new_n410_;
  assign new_n412_ = ~v12 & v15;
  assign new_n413_ = v9 & new_n412_;
  assign new_n414_ = ~v8 & new_n413_;
  assign new_n415_ = ~v7 & new_n414_;
  assign new_n416_ = ~v5 & new_n415_;
  assign new_n417_ = ~v0 & v1;
  assign new_n418_ = ~v4 & v5;
  assign new_n419_ = new_n417_ & new_n418_;
  assign new_n420_ = v8 & ~v10;
  assign new_n421_ = v12 & ~v15;
  assign new_n422_ = new_n420_ & new_n421_;
  assign new_n423_ = new_n419_ & new_n422_;
  assign new_n424_ = ~new_n416_ & ~new_n423_;
  assign new_n425_ = v11 & ~new_n424_;
  assign new_n426_ = ~v6 & new_n425_;
  assign new_n427_ = v4 & new_n333_;
  assign new_n428_ = ~new_n237_ & ~new_n427_;
  assign new_n429_ = v7 & new_n44_;
  assign new_n430_ = ~new_n103_ & ~new_n429_;
  assign new_n431_ = ~v12 & ~new_n430_;
  assign new_n432_ = v10 & new_n431_;
  assign new_n433_ = new_n428_ & ~new_n432_;
  assign new_n434_ = ~v11 & ~new_n433_;
  assign new_n435_ = ~new_n426_ & ~new_n434_;
  assign new_n436_ = v14 & ~new_n435_;
  assign new_n437_ = v5 & ~v10;
  assign new_n438_ = ~v11 & new_n412_;
  assign new_n439_ = new_n437_ & new_n438_;
  assign new_n440_ = ~new_n436_ & ~new_n439_;
  assign new_n441_ = ~new_n411_ & new_n440_;
  assign new_n442_ = v13 & ~new_n441_;
  assign new_n443_ = v5 & new_n38_;
  assign new_n444_ = ~v4 & ~v15;
  assign new_n445_ = ~new_n443_ & ~new_n444_;
  assign new_n446_ = ~v12 & ~new_n445_;
  assign new_n447_ = ~v11 & new_n446_;
  assign new_n448_ = ~v10 & new_n447_;
  assign new_n449_ = ~new_n442_ & ~new_n448_;
  assign \v16.1  = new_n377_ | ~new_n449_;
  assign new_n451_ = ~v1 & ~v10;
  assign new_n452_ = new_n327_ & new_n451_;
  assign new_n453_ = new_n35_ & new_n237_;
  assign new_n454_ = ~new_n452_ & ~new_n453_;
  assign new_n455_ = v0 & ~new_n454_;
  assign new_n456_ = v12 & ~v14;
  assign new_n457_ = v6 & new_n456_;
  assign new_n458_ = ~new_n327_ & ~new_n457_;
  assign new_n459_ = ~v1 & ~new_n458_;
  assign new_n460_ = v4 & v12;
  assign new_n461_ = ~new_n459_ & ~new_n460_;
  assign new_n462_ = v15 & ~new_n461_;
  assign new_n463_ = ~v4 & ~new_n135_;
  assign new_n464_ = v12 & ~new_n421_;
  assign new_n465_ = v4 & ~new_n464_;
  assign new_n466_ = ~new_n463_ & ~new_n465_;
  assign new_n467_ = ~new_n462_ & new_n466_;
  assign new_n468_ = ~v10 & ~new_n467_;
  assign new_n469_ = ~v4 & ~new_n67_;
  assign new_n470_ = v4 & ~new_n45_;
  assign new_n471_ = ~new_n469_ & ~new_n470_;
  assign new_n472_ = ~new_n43_ & ~new_n471_;
  assign new_n473_ = ~v14 & new_n472_;
  assign new_n474_ = v7 & new_n473_;
  assign new_n475_ = ~v6 & new_n474_;
  assign new_n476_ = ~v5 & new_n475_;
  assign new_n477_ = ~new_n52_ & ~new_n476_;
  assign new_n478_ = ~v12 & ~new_n477_;
  assign new_n479_ = v12 & ~new_n40_;
  assign new_n480_ = ~new_n478_ & ~new_n479_;
  assign new_n481_ = v10 & ~new_n480_;
  assign new_n482_ = ~new_n468_ & ~new_n481_;
  assign new_n483_ = ~new_n455_ & new_n482_;
  assign new_n484_ = ~v11 & ~new_n483_;
  assign new_n485_ = v4 & ~new_n93_;
  assign new_n486_ = ~v7 & ~v12;
  assign new_n487_ = ~v1 & new_n486_;
  assign new_n488_ = ~v4 & ~new_n487_;
  assign new_n489_ = ~new_n485_ & ~new_n488_;
  assign new_n490_ = v15 & ~new_n489_;
  assign new_n491_ = v6 & new_n490_;
  assign new_n492_ = ~v15 & ~new_n298_;
  assign new_n493_ = ~v12 & new_n492_;
  assign new_n494_ = ~v4 & new_n493_;
  assign new_n495_ = ~new_n491_ & ~new_n494_;
  assign new_n496_ = ~v10 & ~new_n495_;
  assign new_n497_ = ~v12 & ~new_n298_;
  assign new_n498_ = v10 & new_n497_;
  assign new_n499_ = ~new_n496_ & ~new_n498_;
  assign new_n500_ = v5 & ~new_n499_;
  assign new_n501_ = ~v7 & ~v9;
  assign new_n502_ = ~v4 & ~new_n501_;
  assign new_n503_ = v4 & v7;
  assign new_n504_ = ~new_n502_ & ~new_n503_;
  assign new_n505_ = v12 & ~new_n504_;
  assign new_n506_ = ~v5 & new_n505_;
  assign new_n507_ = v7 & new_n224_;
  assign new_n508_ = ~new_n506_ & ~new_n507_;
  assign new_n509_ = v10 & ~new_n508_;
  assign new_n510_ = ~v8 & new_n509_;
  assign new_n511_ = ~v6 & new_n510_;
  assign new_n512_ = ~new_n500_ & ~new_n511_;
  assign new_n513_ = ~v14 & ~new_n512_;
  assign new_n514_ = v15 & ~new_n298_;
  assign new_n515_ = v14 & new_n514_;
  assign new_n516_ = ~v4 & new_n515_;
  assign new_n517_ = ~v6 & new_n103_;
  assign new_n518_ = new_n364_ & new_n517_;
  assign new_n519_ = ~new_n516_ & ~new_n518_;
  assign new_n520_ = ~v10 & ~new_n519_;
  assign new_n521_ = v15 & ~new_n365_;
  assign new_n522_ = v10 & ~new_n521_;
  assign new_n523_ = ~new_n520_ & ~new_n522_;
  assign new_n524_ = v5 & ~new_n523_;
  assign new_n525_ = ~v15 & ~new_n67_;
  assign new_n526_ = v10 & new_n525_;
  assign new_n527_ = ~v7 & new_n526_;
  assign new_n528_ = ~v6 & new_n527_;
  assign new_n529_ = ~new_n524_ & ~new_n528_;
  assign new_n530_ = ~v12 & ~new_n529_;
  assign new_n531_ = ~new_n513_ & ~new_n530_;
  assign new_n532_ = ~v0 & ~new_n531_;
  assign new_n533_ = v8 & ~new_n112_;
  assign new_n534_ = v7 & new_n533_;
  assign new_n535_ = v6 & new_n534_;
  assign new_n536_ = v5 & new_n535_;
  assign new_n537_ = ~new_n191_ & ~new_n536_;
  assign new_n538_ = ~v4 & ~new_n537_;
  assign new_n539_ = v1 & v5;
  assign new_n540_ = new_n365_ & new_n539_;
  assign new_n541_ = ~v15 & ~new_n540_;
  assign new_n542_ = v14 & new_n541_;
  assign new_n543_ = ~new_n538_ & ~new_n542_;
  assign new_n544_ = ~v12 & ~new_n543_;
  assign new_n545_ = v12 & new_n35_;
  assign new_n546_ = v9 & new_n545_;
  assign new_n547_ = v8 & new_n546_;
  assign new_n548_ = ~v7 & new_n547_;
  assign new_n549_ = ~v6 & new_n548_;
  assign new_n550_ = ~v5 & new_n549_;
  assign new_n551_ = ~new_n544_ & ~new_n550_;
  assign new_n552_ = ~v10 & ~new_n551_;
  assign new_n553_ = ~v12 & ~new_n58_;
  assign new_n554_ = v10 & new_n553_;
  assign new_n555_ = v7 & new_n554_;
  assign new_n556_ = v6 & new_n555_;
  assign new_n557_ = v5 & new_n556_;
  assign new_n558_ = ~new_n552_ & ~new_n557_;
  assign new_n559_ = ~new_n532_ & new_n558_;
  assign new_n560_ = v11 & ~new_n559_;
  assign new_n561_ = ~new_n484_ & ~new_n560_;
  assign new_n562_ = ~v13 & ~new_n561_;
  assign new_n563_ = ~v14 & ~new_n388_;
  assign new_n564_ = ~v14 & ~new_n563_;
  assign new_n565_ = v12 & ~new_n564_;
  assign new_n566_ = v10 & new_n565_;
  assign new_n567_ = ~v12 & ~new_n321_;
  assign new_n568_ = ~v10 & new_n567_;
  assign new_n569_ = ~new_n566_ & ~new_n568_;
  assign new_n570_ = ~v11 & ~new_n569_;
  assign new_n571_ = ~v8 & new_n211_;
  assign new_n572_ = ~v10 & ~v14;
  assign new_n573_ = new_n159_ & new_n572_;
  assign new_n574_ = ~new_n571_ & ~new_n573_;
  assign new_n575_ = ~v4 & ~new_n574_;
  assign new_n576_ = v4 & v8;
  assign new_n577_ = ~v9 & new_n572_;
  assign new_n578_ = new_n576_ & new_n577_;
  assign new_n579_ = ~new_n575_ & ~new_n578_;
  assign new_n580_ = ~v12 & ~new_n579_;
  assign new_n581_ = ~v7 & new_n580_;
  assign new_n582_ = ~v6 & new_n581_;
  assign new_n583_ = ~v10 & new_n456_;
  assign new_n584_ = ~new_n582_ & ~new_n583_;
  assign new_n585_ = v11 & ~new_n584_;
  assign new_n586_ = ~v5 & new_n585_;
  assign new_n587_ = ~new_n570_ & ~new_n586_;
  assign new_n588_ = v15 & ~new_n587_;
  assign new_n589_ = v6 & ~v14;
  assign new_n590_ = ~v2 & new_n589_;
  assign new_n591_ = new_n191_ & new_n365_;
  assign new_n592_ = ~new_n590_ & ~new_n591_;
  assign new_n593_ = v1 & ~new_n592_;
  assign new_n594_ = ~v2 & v6;
  assign new_n595_ = v7 & ~v14;
  assign new_n596_ = new_n594_ & new_n595_;
  assign new_n597_ = ~new_n593_ & ~new_n596_;
  assign new_n598_ = v12 & ~new_n597_;
  assign new_n599_ = v11 & new_n598_;
  assign new_n600_ = v5 & new_n599_;
  assign new_n601_ = ~v0 & new_n600_;
  assign new_n602_ = ~new_n225_ & ~new_n601_;
  assign new_n603_ = v4 & ~new_n602_;
  assign new_n604_ = v5 & ~new_n597_;
  assign new_n605_ = ~v4 & new_n604_;
  assign new_n606_ = ~v0 & new_n605_;
  assign new_n607_ = ~v5 & new_n35_;
  assign new_n608_ = ~new_n606_ & ~new_n607_;
  assign new_n609_ = v12 & ~new_n608_;
  assign new_n610_ = v11 & new_n609_;
  assign new_n611_ = ~new_n603_ & ~new_n610_;
  assign new_n612_ = ~v10 & ~new_n611_;
  assign new_n613_ = ~new_n421_ & ~new_n431_;
  assign new_n614_ = v14 & ~new_n613_;
  assign new_n615_ = ~new_n35_ & ~new_n614_;
  assign new_n616_ = ~v11 & ~new_n615_;
  assign new_n617_ = v10 & new_n616_;
  assign new_n618_ = ~new_n612_ & ~new_n617_;
  assign new_n619_ = ~new_n588_ & new_n618_;
  assign new_n620_ = v13 & ~new_n619_;
  assign new_n621_ = ~new_n448_ & ~new_n620_;
  assign \v16.2  = new_n562_ | ~new_n621_;
  assign new_n623_ = ~v1 & v6;
  assign new_n624_ = ~v4 & ~new_n623_;
  assign new_n625_ = v15 & ~new_n624_;
  assign new_n626_ = v4 & ~v15;
  assign new_n627_ = ~new_n625_ & ~new_n626_;
  assign new_n628_ = ~v10 & ~new_n627_;
  assign new_n629_ = ~v0 & v15;
  assign new_n630_ = v0 & ~v15;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign new_n632_ = v10 & ~new_n631_;
  assign new_n633_ = ~new_n628_ & ~new_n632_;
  assign new_n634_ = v12 & ~new_n633_;
  assign new_n635_ = ~v12 & new_n472_;
  assign new_n636_ = v10 & new_n635_;
  assign new_n637_ = v7 & new_n636_;
  assign new_n638_ = ~v6 & new_n637_;
  assign new_n639_ = ~v5 & new_n638_;
  assign new_n640_ = ~new_n634_ & ~new_n639_;
  assign new_n641_ = ~v14 & ~new_n640_;
  assign new_n642_ = ~v0 & new_n444_;
  assign new_n643_ = ~v15 & ~new_n642_;
  assign new_n644_ = v14 & ~new_n643_;
  assign new_n645_ = ~v12 & new_n644_;
  assign new_n646_ = ~v10 & new_n645_;
  assign new_n647_ = ~new_n332_ & ~new_n646_;
  assign new_n648_ = ~v1 & ~new_n647_;
  assign new_n649_ = ~v10 & ~new_n337_;
  assign new_n650_ = v12 & ~new_n649_;
  assign new_n651_ = v10 & ~v12;
  assign new_n652_ = ~v0 & new_n651_;
  assign new_n653_ = ~new_n650_ & ~new_n652_;
  assign new_n654_ = v14 & ~new_n653_;
  assign new_n655_ = ~new_n427_ & ~new_n654_;
  assign new_n656_ = ~new_n648_ & new_n655_;
  assign new_n657_ = ~new_n641_ & new_n656_;
  assign new_n658_ = ~v11 & ~new_n657_;
  assign new_n659_ = v4 & ~new_n97_;
  assign new_n660_ = ~v4 & ~new_n298_;
  assign new_n661_ = ~new_n659_ & ~new_n660_;
  assign new_n662_ = ~v15 & ~new_n661_;
  assign new_n663_ = ~v12 & new_n662_;
  assign new_n664_ = ~v4 & v12;
  assign new_n665_ = new_n142_ & ~new_n664_;
  assign new_n666_ = v15 & ~new_n665_;
  assign new_n667_ = v6 & new_n666_;
  assign new_n668_ = ~new_n663_ & ~new_n667_;
  assign new_n669_ = ~v14 & ~new_n668_;
  assign new_n670_ = ~v12 & ~new_n519_;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = ~v10 & ~new_n671_;
  assign new_n673_ = new_n58_ & ~new_n63_;
  assign new_n674_ = ~v12 & ~new_n673_;
  assign new_n675_ = v10 & new_n674_;
  assign new_n676_ = ~new_n672_ & ~new_n675_;
  assign new_n677_ = v5 & ~new_n676_;
  assign new_n678_ = ~v14 & ~new_n508_;
  assign new_n679_ = ~v8 & new_n678_;
  assign new_n680_ = ~v12 & new_n525_;
  assign new_n681_ = ~v7 & new_n680_;
  assign new_n682_ = ~new_n679_ & ~new_n681_;
  assign new_n683_ = v10 & ~new_n682_;
  assign new_n684_ = ~v6 & new_n683_;
  assign new_n685_ = ~new_n677_ & ~new_n684_;
  assign new_n686_ = ~v0 & ~new_n685_;
  assign new_n687_ = ~v7 & new_n121_;
  assign new_n688_ = new_n119_ & new_n687_;
  assign new_n689_ = v5 & v6;
  assign new_n690_ = v7 & ~v12;
  assign new_n691_ = new_n689_ & new_n690_;
  assign new_n692_ = ~new_n688_ & ~new_n691_;
  assign new_n693_ = ~v14 & ~new_n692_;
  assign new_n694_ = v8 & new_n693_;
  assign new_n695_ = ~v12 & new_n368_;
  assign new_n696_ = ~new_n694_ & ~new_n695_;
  assign new_n697_ = ~v15 & ~new_n696_;
  assign new_n698_ = new_n59_ & new_n418_;
  assign new_n699_ = v8 & ~v12;
  assign new_n700_ = new_n102_ & new_n699_;
  assign new_n701_ = new_n698_ & new_n700_;
  assign new_n702_ = ~new_n697_ & ~new_n701_;
  assign new_n703_ = ~v10 & ~new_n702_;
  assign new_n704_ = ~new_n557_ & ~new_n703_;
  assign new_n705_ = ~new_n686_ & new_n704_;
  assign new_n706_ = v11 & ~new_n705_;
  assign new_n707_ = ~new_n658_ & ~new_n706_;
  assign new_n708_ = ~v13 & ~new_n707_;
  assign new_n709_ = v14 & ~new_n430_;
  assign new_n710_ = v14 & ~new_n709_;
  assign new_n711_ = ~v12 & ~new_n710_;
  assign new_n712_ = ~new_n35_ & ~new_n711_;
  assign new_n713_ = ~v11 & ~new_n712_;
  assign new_n714_ = v10 & new_n713_;
  assign new_n715_ = ~new_n612_ & ~new_n714_;
  assign new_n716_ = ~new_n588_ & new_n715_;
  assign new_n717_ = v13 & ~new_n716_;
  assign new_n718_ = v5 & new_n200_;
  assign new_n719_ = ~v12 & new_n38_;
  assign new_n720_ = new_n718_ & new_n719_;
  assign new_n721_ = ~new_n717_ & ~new_n720_;
  assign \v16.3  = new_n708_ | ~new_n721_;
  assign new_n723_ = ~new_n223_ & ~new_n638_;
  assign new_n724_ = ~v5 & ~new_n723_;
  assign new_n725_ = ~new_n634_ & ~new_n724_;
  assign new_n726_ = ~v14 & ~new_n725_;
  assign new_n727_ = new_n347_ & ~new_n726_;
  assign new_n728_ = ~v11 & ~new_n727_;
  assign new_n729_ = ~new_n112_ & ~new_n298_;
  assign new_n730_ = ~v12 & new_n729_;
  assign new_n731_ = v15 & ~new_n487_;
  assign new_n732_ = ~v14 & new_n731_;
  assign new_n733_ = v6 & new_n732_;
  assign new_n734_ = ~new_n730_ & ~new_n733_;
  assign new_n735_ = ~v4 & ~new_n734_;
  assign new_n736_ = ~v14 & new_n231_;
  assign new_n737_ = v6 & new_n736_;
  assign new_n738_ = v4 & new_n737_;
  assign new_n739_ = ~new_n735_ & ~new_n738_;
  assign new_n740_ = ~v10 & ~new_n739_;
  assign new_n741_ = ~new_n675_ & ~new_n740_;
  assign new_n742_ = v5 & ~new_n741_;
  assign new_n743_ = v4 & ~new_n78_;
  assign new_n744_ = ~new_n502_ & ~new_n743_;
  assign new_n745_ = v12 & ~new_n744_;
  assign new_n746_ = ~v5 & new_n745_;
  assign new_n747_ = ~new_n507_ & ~new_n746_;
  assign new_n748_ = ~v14 & ~new_n747_;
  assign new_n749_ = ~v8 & new_n748_;
  assign new_n750_ = ~new_n681_ & ~new_n749_;
  assign new_n751_ = v10 & ~new_n750_;
  assign new_n752_ = ~v6 & new_n751_;
  assign new_n753_ = ~new_n742_ & ~new_n752_;
  assign new_n754_ = ~v0 & ~new_n753_;
  assign new_n755_ = v7 & new_n113_;
  assign new_n756_ = v6 & new_n755_;
  assign new_n757_ = v5 & new_n756_;
  assign new_n758_ = new_n122_ & new_n268_;
  assign new_n759_ = ~new_n757_ & ~new_n758_;
  assign new_n760_ = v8 & ~new_n759_;
  assign new_n761_ = ~v15 & ~new_n367_;
  assign new_n762_ = v14 & new_n761_;
  assign new_n763_ = ~v12 & new_n762_;
  assign new_n764_ = ~new_n760_ & ~new_n763_;
  assign new_n765_ = ~v10 & ~new_n764_;
  assign new_n766_ = ~new_n557_ & ~new_n765_;
  assign new_n767_ = ~new_n754_ & new_n766_;
  assign new_n768_ = v11 & ~new_n767_;
  assign new_n769_ = ~new_n728_ & ~new_n768_;
  assign new_n770_ = ~v13 & ~new_n769_;
  assign new_n771_ = v6 & ~new_n142_;
  assign new_n772_ = v5 & new_n771_;
  assign new_n773_ = ~v2 & new_n772_;
  assign new_n774_ = ~v0 & new_n773_;
  assign new_n775_ = v5 & ~new_n774_;
  assign new_n776_ = v11 & ~new_n775_;
  assign new_n777_ = ~v10 & new_n776_;
  assign new_n778_ = ~new_n391_ & ~new_n777_;
  assign new_n779_ = v12 & ~new_n778_;
  assign new_n780_ = ~new_n407_ & ~new_n779_;
  assign new_n781_ = ~v14 & ~new_n780_;
  assign new_n782_ = new_n440_ & ~new_n781_;
  assign new_n783_ = v13 & ~new_n782_;
  assign new_n784_ = ~new_n448_ & ~new_n783_;
  assign \v16.4  = new_n770_ | ~new_n784_;
  assign new_n786_ = v13 & ~v14;
  assign new_n787_ = v10 & new_n786_;
  assign new_n788_ = ~new_n296_ & ~new_n787_;
  assign new_n789_ = ~v12 & ~new_n788_;
  assign new_n790_ = ~v10 & ~new_n135_;
  assign new_n791_ = ~v4 & new_n790_;
  assign new_n792_ = v0 & new_n34_;
  assign new_n793_ = ~v14 & ~new_n792_;
  assign new_n794_ = v12 & ~new_n793_;
  assign new_n795_ = v10 & new_n794_;
  assign new_n796_ = ~new_n791_ & ~new_n795_;
  assign new_n797_ = ~v13 & ~new_n796_;
  assign new_n798_ = v12 & v14;
  assign new_n799_ = ~new_n35_ & ~new_n798_;
  assign new_n800_ = v13 & ~new_n799_;
  assign new_n801_ = v10 & new_n800_;
  assign new_n802_ = ~new_n797_ & ~new_n801_;
  assign new_n803_ = ~new_n789_ & new_n802_;
  assign \v16.5  = ~v11 & ~new_n803_;
  assign new_n805_ = ~v11 & new_n42_;
  assign new_n806_ = v11 & new_n76_;
  assign new_n807_ = ~new_n805_ & ~new_n806_;
  assign new_n808_ = ~v13 & ~new_n807_;
  assign new_n809_ = ~v12 & ~new_n431_;
  assign new_n810_ = v14 & ~new_n809_;
  assign new_n811_ = ~v14 & ~new_n329_;
  assign new_n812_ = ~new_n810_ & ~new_n811_;
  assign new_n813_ = v13 & ~new_n812_;
  assign new_n814_ = ~v11 & new_n813_;
  assign new_n815_ = ~new_n808_ & ~new_n814_;
  assign new_n816_ = v10 & ~new_n815_;
  assign new_n817_ = v4 & v13;
  assign new_n818_ = new_n102_ & new_n817_;
  assign new_n819_ = ~new_n444_ & ~new_n818_;
  assign new_n820_ = ~v12 & ~new_n819_;
  assign new_n821_ = v4 & new_n130_;
  assign new_n822_ = ~new_n463_ & ~new_n821_;
  assign new_n823_ = ~v13 & ~new_n822_;
  assign new_n824_ = ~new_n820_ & ~new_n823_;
  assign new_n825_ = ~v11 & ~new_n824_;
  assign new_n826_ = ~v10 & new_n825_;
  assign \v16.6  = new_n816_ | new_n826_;
  assign new_n828_ = v15 & ~new_n458_;
  assign new_n829_ = ~v10 & new_n828_;
  assign new_n830_ = ~new_n332_ & ~new_n829_;
  assign new_n831_ = ~v1 & ~new_n830_;
  assign new_n832_ = ~new_n478_ & ~new_n798_;
  assign new_n833_ = v10 & ~new_n832_;
  assign new_n834_ = v6 & v12;
  assign new_n835_ = new_n38_ & new_n834_;
  assign new_n836_ = v12 & ~new_n835_;
  assign new_n837_ = v4 & ~new_n836_;
  assign new_n838_ = ~new_n463_ & ~new_n837_;
  assign new_n839_ = ~v10 & ~new_n838_;
  assign new_n840_ = ~new_n833_ & ~new_n839_;
  assign new_n841_ = ~new_n831_ & new_n840_;
  assign new_n842_ = ~v11 & ~new_n841_;
  assign new_n843_ = ~new_n491_ & ~new_n663_;
  assign new_n844_ = ~v14 & ~new_n843_;
  assign new_n845_ = v15 & ~new_n661_;
  assign new_n846_ = v14 & new_n845_;
  assign new_n847_ = ~new_n518_ & ~new_n846_;
  assign new_n848_ = ~v12 & ~new_n847_;
  assign new_n849_ = ~new_n844_ & ~new_n848_;
  assign new_n850_ = ~v0 & ~new_n849_;
  assign new_n851_ = ~new_n116_ & ~new_n850_;
  assign new_n852_ = v5 & ~new_n851_;
  assign new_n853_ = v8 & v9;
  assign new_n854_ = new_n456_ & new_n853_;
  assign new_n855_ = new_n268_ & new_n854_;
  assign new_n856_ = ~new_n327_ & ~new_n855_;
  assign new_n857_ = ~v4 & ~new_n856_;
  assign new_n858_ = v4 & new_n185_;
  assign new_n859_ = new_n854_ & new_n858_;
  assign new_n860_ = ~new_n327_ & ~new_n859_;
  assign new_n861_ = ~v5 & ~new_n860_;
  assign new_n862_ = v1 & new_n365_;
  assign new_n863_ = v14 & ~new_n862_;
  assign new_n864_ = ~v12 & new_n863_;
  assign new_n865_ = ~new_n861_ & ~new_n864_;
  assign new_n866_ = ~new_n857_ & new_n865_;
  assign new_n867_ = ~v15 & ~new_n866_;
  assign new_n868_ = ~new_n852_ & ~new_n867_;
  assign new_n869_ = ~v10 & ~new_n868_;
  assign new_n870_ = ~v14 & ~new_n744_;
  assign new_n871_ = v12 & new_n870_;
  assign new_n872_ = v10 & new_n871_;
  assign new_n873_ = ~v8 & new_n872_;
  assign new_n874_ = ~v6 & new_n873_;
  assign new_n875_ = ~v5 & new_n874_;
  assign new_n876_ = ~v0 & new_n875_;
  assign new_n877_ = ~new_n869_ & ~new_n876_;
  assign new_n878_ = v11 & ~new_n877_;
  assign new_n879_ = ~new_n842_ & ~new_n878_;
  assign new_n880_ = ~v13 & ~new_n879_;
  assign new_n881_ = ~v14 & ~new_n775_;
  assign new_n882_ = v8 & new_n191_;
  assign new_n883_ = ~v6 & new_n882_;
  assign new_n884_ = v5 & new_n883_;
  assign new_n885_ = v1 & new_n884_;
  assign new_n886_ = ~v0 & new_n885_;
  assign new_n887_ = ~new_n881_ & ~new_n886_;
  assign new_n888_ = v12 & ~new_n887_;
  assign new_n889_ = ~v9 & ~v14;
  assign new_n890_ = v8 & new_n889_;
  assign new_n891_ = ~new_n571_ & ~new_n890_;
  assign new_n892_ = v4 & ~new_n891_;
  assign new_n893_ = new_n349_ & new_n889_;
  assign new_n894_ = ~new_n892_ & ~new_n893_;
  assign new_n895_ = v15 & ~new_n894_;
  assign new_n896_ = ~v12 & new_n895_;
  assign new_n897_ = ~v7 & new_n896_;
  assign new_n898_ = ~v6 & new_n897_;
  assign new_n899_ = ~v5 & new_n898_;
  assign new_n900_ = ~new_n888_ & ~new_n899_;
  assign new_n901_ = ~v10 & ~new_n900_;
  assign new_n902_ = v4 & v10;
  assign new_n903_ = v4 & ~new_n902_;
  assign new_n904_ = v15 & ~new_n903_;
  assign new_n905_ = v14 & new_n904_;
  assign new_n906_ = ~v12 & new_n905_;
  assign new_n907_ = v9 & new_n906_;
  assign new_n908_ = ~v8 & new_n907_;
  assign new_n909_ = ~v7 & new_n908_;
  assign new_n910_ = ~v6 & new_n909_;
  assign new_n911_ = ~v5 & new_n910_;
  assign new_n912_ = ~new_n901_ & ~new_n911_;
  assign new_n913_ = v11 & ~new_n912_;
  assign new_n914_ = v15 & ~new_n564_;
  assign new_n915_ = ~new_n191_ & ~new_n914_;
  assign new_n916_ = v12 & ~new_n915_;
  assign new_n917_ = ~new_n811_ & ~new_n916_;
  assign new_n918_ = v10 & ~new_n917_;
  assign new_n919_ = v14 & ~new_n191_;
  assign new_n920_ = v4 & ~new_n919_;
  assign new_n921_ = v5 & v15;
  assign new_n922_ = ~new_n920_ & ~new_n921_;
  assign new_n923_ = ~v12 & ~new_n922_;
  assign new_n924_ = ~v10 & new_n923_;
  assign new_n925_ = ~new_n918_ & ~new_n924_;
  assign new_n926_ = ~v11 & ~new_n925_;
  assign new_n927_ = ~new_n913_ & ~new_n926_;
  assign new_n928_ = v13 & ~new_n927_;
  assign new_n929_ = ~new_n448_ & ~new_n928_;
  assign \v16.7  = new_n880_ | ~new_n929_;
  assign new_n931_ = ~v14 & ~new_n37_;
  assign new_n932_ = ~v11 & ~new_n931_;
  assign new_n933_ = v11 & new_n79_;
  assign new_n934_ = ~v8 & new_n933_;
  assign new_n935_ = ~v6 & new_n934_;
  assign new_n936_ = ~v5 & new_n935_;
  assign new_n937_ = v4 & new_n936_;
  assign new_n938_ = ~v0 & new_n937_;
  assign new_n939_ = ~new_n932_ & ~new_n938_;
  assign new_n940_ = v10 & ~new_n939_;
  assign new_n941_ = v6 & v15;
  assign new_n942_ = v5 & new_n941_;
  assign new_n943_ = ~v1 & new_n942_;
  assign new_n944_ = ~v0 & new_n943_;
  assign new_n945_ = v9 & ~v15;
  assign new_n946_ = v8 & new_n945_;
  assign new_n947_ = new_n119_ & new_n946_;
  assign new_n948_ = ~new_n944_ & ~new_n947_;
  assign new_n949_ = ~v14 & ~new_n948_;
  assign new_n950_ = v11 & new_n949_;
  assign new_n951_ = ~v7 & new_n950_;
  assign new_n952_ = v4 & new_n951_;
  assign new_n953_ = ~v4 & ~v11;
  assign new_n954_ = ~new_n952_ & ~new_n953_;
  assign new_n955_ = ~v10 & ~new_n954_;
  assign new_n956_ = ~new_n940_ & ~new_n955_;
  assign new_n957_ = v12 & ~new_n956_;
  assign new_n958_ = ~v5 & new_n162_;
  assign new_n959_ = v9 & new_n178_;
  assign new_n960_ = new_n958_ & new_n959_;
  assign new_n961_ = v11 & ~v15;
  assign new_n962_ = new_n437_ & new_n961_;
  assign new_n963_ = ~new_n960_ & ~new_n962_;
  assign new_n964_ = ~v0 & ~new_n963_;
  assign new_n965_ = v9 & v10;
  assign new_n966_ = new_n203_ & new_n965_;
  assign new_n967_ = new_n958_ & new_n966_;
  assign new_n968_ = ~new_n964_ & ~new_n967_;
  assign new_n969_ = ~v14 & ~new_n968_;
  assign new_n970_ = v11 & ~new_n105_;
  assign new_n971_ = ~v10 & new_n970_;
  assign new_n972_ = v5 & new_n971_;
  assign new_n973_ = ~v0 & new_n972_;
  assign new_n974_ = ~new_n969_ & ~new_n973_;
  assign new_n975_ = ~v6 & ~new_n974_;
  assign new_n976_ = ~v0 & ~v7;
  assign new_n977_ = ~new_n59_ & ~new_n976_;
  assign new_n978_ = ~new_n112_ & ~new_n977_;
  assign new_n979_ = v11 & new_n978_;
  assign new_n980_ = ~v10 & new_n979_;
  assign new_n981_ = v8 & new_n980_;
  assign new_n982_ = v5 & new_n981_;
  assign new_n983_ = ~new_n975_ & ~new_n982_;
  assign new_n984_ = ~v12 & ~new_n983_;
  assign new_n985_ = v11 & new_n736_;
  assign new_n986_ = ~v10 & new_n985_;
  assign new_n987_ = v6 & new_n986_;
  assign new_n988_ = v5 & new_n987_;
  assign new_n989_ = ~v0 & new_n988_;
  assign new_n990_ = ~new_n984_ & ~new_n989_;
  assign new_n991_ = v4 & ~new_n990_;
  assign new_n992_ = new_n208_ & new_n321_;
  assign new_n993_ = ~new_n991_ & ~new_n992_;
  assign new_n994_ = ~new_n957_ & new_n993_;
  assign new_n995_ = ~v13 & ~new_n994_;
  assign new_n996_ = v12 & new_n191_;
  assign new_n997_ = v5 & new_n996_;
  assign new_n998_ = v1 & new_n997_;
  assign new_n999_ = ~v0 & new_n998_;
  assign new_n1000_ = ~v5 & new_n501_;
  assign new_n1001_ = new_n719_ & new_n1000_;
  assign new_n1002_ = ~new_n999_ & ~new_n1001_;
  assign new_n1003_ = v8 & ~new_n1002_;
  assign new_n1004_ = ~v7 & ~v8;
  assign new_n1005_ = ~v5 & new_n1004_;
  assign new_n1006_ = v9 & ~v12;
  assign new_n1007_ = new_n102_ & new_n1006_;
  assign new_n1008_ = new_n1005_ & new_n1007_;
  assign new_n1009_ = ~new_n1003_ & ~new_n1008_;
  assign new_n1010_ = ~v6 & ~new_n1009_;
  assign new_n1011_ = ~v14 & ~new_n142_;
  assign new_n1012_ = v12 & new_n1011_;
  assign new_n1013_ = v6 & new_n1012_;
  assign new_n1014_ = v5 & new_n1013_;
  assign new_n1015_ = ~v2 & new_n1014_;
  assign new_n1016_ = ~v0 & new_n1015_;
  assign new_n1017_ = ~new_n1010_ & ~new_n1016_;
  assign new_n1018_ = v11 & ~new_n1017_;
  assign new_n1019_ = ~v12 & ~new_n919_;
  assign new_n1020_ = ~v11 & new_n1019_;
  assign new_n1021_ = ~new_n1018_ & ~new_n1020_;
  assign new_n1022_ = v4 & ~new_n1021_;
  assign new_n1023_ = v11 & new_n456_;
  assign new_n1024_ = ~v5 & new_n1023_;
  assign new_n1025_ = ~new_n1022_ & ~new_n1024_;
  assign new_n1026_ = ~v10 & ~new_n1025_;
  assign new_n1027_ = v7 & ~v11;
  assign new_n1028_ = v4 & new_n119_;
  assign new_n1029_ = v11 & v15;
  assign new_n1030_ = ~v7 & new_n1029_;
  assign new_n1031_ = new_n1028_ & new_n1030_;
  assign new_n1032_ = ~new_n1027_ & ~new_n1031_;
  assign new_n1033_ = v9 & ~new_n1032_;
  assign new_n1034_ = ~v8 & new_n1033_;
  assign new_n1035_ = v8 & new_n203_;
  assign new_n1036_ = ~new_n1034_ & ~new_n1035_;
  assign new_n1037_ = ~v12 & ~new_n1036_;
  assign new_n1038_ = ~v11 & v12;
  assign new_n1039_ = ~new_n1037_ & ~new_n1038_;
  assign new_n1040_ = v14 & ~new_n1039_;
  assign new_n1041_ = ~v11 & new_n811_;
  assign new_n1042_ = ~new_n1040_ & ~new_n1041_;
  assign new_n1043_ = v10 & ~new_n1042_;
  assign new_n1044_ = ~new_n1026_ & ~new_n1043_;
  assign new_n1045_ = v13 & ~new_n1044_;
  assign new_n1046_ = ~new_n226_ & ~new_n1045_;
  assign \v16.8  = new_n995_ | ~new_n1046_;
  assign new_n1048_ = v11 & v12;
  assign new_n1049_ = new_n1004_ & new_n1048_;
  assign new_n1050_ = new_n150_ & new_n243_;
  assign new_n1051_ = ~new_n1049_ & ~new_n1050_;
  assign new_n1052_ = ~v0 & ~new_n1051_;
  assign new_n1053_ = new_n150_ & new_n225_;
  assign new_n1054_ = ~new_n1052_ & ~new_n1053_;
  assign new_n1055_ = ~v14 & ~new_n1054_;
  assign new_n1056_ = ~v13 & new_n1055_;
  assign new_n1057_ = ~v8 & v11;
  assign new_n1058_ = ~v7 & new_n1057_;
  assign new_n1059_ = ~v12 & v13;
  assign new_n1060_ = new_n102_ & new_n1059_;
  assign new_n1061_ = new_n1058_ & new_n1060_;
  assign new_n1062_ = ~new_n1056_ & ~new_n1061_;
  assign new_n1063_ = v9 & ~new_n1062_;
  assign new_n1064_ = ~v14 & ~new_n43_;
  assign new_n1065_ = ~v13 & new_n1064_;
  assign new_n1066_ = ~v12 & new_n1065_;
  assign new_n1067_ = ~v11 & new_n1066_;
  assign new_n1068_ = ~v9 & new_n1067_;
  assign new_n1069_ = v8 & new_n1068_;
  assign new_n1070_ = v7 & new_n1069_;
  assign new_n1071_ = ~new_n1063_ & ~new_n1070_;
  assign new_n1072_ = ~v6 & ~new_n1071_;
  assign new_n1073_ = ~v5 & new_n1072_;
  assign new_n1074_ = v4 & new_n1073_;
  assign new_n1075_ = ~v13 & v15;
  assign new_n1076_ = v0 & ~v1;
  assign new_n1077_ = new_n1075_ & new_n1076_;
  assign new_n1078_ = ~v14 & ~new_n1077_;
  assign new_n1079_ = v12 & ~new_n1078_;
  assign new_n1080_ = v13 & new_n811_;
  assign new_n1081_ = ~new_n1079_ & ~new_n1080_;
  assign new_n1082_ = ~v11 & ~new_n1081_;
  assign new_n1083_ = ~new_n1074_ & ~new_n1082_;
  assign new_n1084_ = v10 & ~new_n1083_;
  assign new_n1085_ = ~v6 & new_n38_;
  assign new_n1086_ = ~v14 & ~new_n1085_;
  assign new_n1087_ = v12 & ~new_n1086_;
  assign new_n1088_ = v4 & new_n1087_;
  assign new_n1089_ = ~new_n463_ & ~new_n1088_;
  assign new_n1090_ = ~v11 & ~new_n1089_;
  assign new_n1091_ = ~v6 & new_n96_;
  assign new_n1092_ = new_n184_ & new_n1091_;
  assign new_n1093_ = new_n195_ & new_n545_;
  assign new_n1094_ = new_n1092_ & new_n1093_;
  assign new_n1095_ = ~new_n1090_ & ~new_n1094_;
  assign new_n1096_ = ~v13 & ~new_n1095_;
  assign new_n1097_ = new_n224_ & new_n953_;
  assign new_n1098_ = ~new_n1096_ & ~new_n1097_;
  assign new_n1099_ = ~v10 & ~new_n1098_;
  assign \v16.9  = new_n1084_ | new_n1099_;
  assign new_n1101_ = ~v0 & ~v15;
  assign new_n1102_ = ~v13 & ~new_n1101_;
  assign new_n1103_ = ~v1 & new_n1102_;
  assign new_n1104_ = ~new_n817_ & ~new_n1103_;
  assign new_n1105_ = v14 & ~new_n1104_;
  assign new_n1106_ = ~v13 & v14;
  assign new_n1107_ = v5 & ~new_n1106_;
  assign new_n1108_ = v4 & new_n786_;
  assign new_n1109_ = ~new_n1107_ & ~new_n1108_;
  assign new_n1110_ = v15 & ~new_n1109_;
  assign new_n1111_ = v13 & new_n35_;
  assign new_n1112_ = v13 & ~new_n1111_;
  assign new_n1113_ = v4 & ~new_n1112_;
  assign new_n1114_ = ~new_n444_ & ~new_n1113_;
  assign new_n1115_ = ~new_n1110_ & new_n1114_;
  assign new_n1116_ = ~new_n1105_ & new_n1115_;
  assign new_n1117_ = ~v12 & ~new_n1116_;
  assign new_n1118_ = ~v13 & ~new_n135_;
  assign new_n1119_ = ~v4 & new_n1118_;
  assign new_n1120_ = ~new_n1117_ & ~new_n1119_;
  assign new_n1121_ = ~v10 & ~new_n1120_;
  assign new_n1122_ = ~v13 & ~new_n931_;
  assign new_n1123_ = ~v4 & new_n162_;
  assign new_n1124_ = ~v4 & ~new_n1123_;
  assign new_n1125_ = v15 & ~new_n1124_;
  assign new_n1126_ = ~v14 & new_n1125_;
  assign new_n1127_ = ~v14 & ~new_n1126_;
  assign new_n1128_ = v13 & ~new_n1127_;
  assign new_n1129_ = ~new_n1122_ & ~new_n1128_;
  assign new_n1130_ = v12 & ~new_n1129_;
  assign new_n1131_ = ~v0 & new_n1106_;
  assign new_n1132_ = ~new_n786_ & ~new_n1131_;
  assign new_n1133_ = ~v12 & ~new_n1132_;
  assign new_n1134_ = ~new_n1111_ & ~new_n1133_;
  assign new_n1135_ = ~new_n1130_ & new_n1134_;
  assign new_n1136_ = v10 & ~new_n1135_;
  assign new_n1137_ = ~new_n1121_ & ~new_n1136_;
  assign new_n1138_ = ~v11 & ~new_n1137_;
  assign new_n1139_ = v6 & new_n231_;
  assign new_n1140_ = ~new_n99_ & ~new_n1139_;
  assign new_n1141_ = ~v10 & ~new_n1140_;
  assign new_n1142_ = v5 & new_n1141_;
  assign new_n1143_ = ~v9 & new_n237_;
  assign new_n1144_ = ~v8 & new_n1143_;
  assign new_n1145_ = v7 & new_n1144_;
  assign new_n1146_ = ~v6 & new_n1145_;
  assign new_n1147_ = ~v5 & new_n1146_;
  assign new_n1148_ = ~new_n1142_ & ~new_n1147_;
  assign new_n1149_ = ~v13 & ~new_n1148_;
  assign new_n1150_ = v13 & ~new_n142_;
  assign new_n1151_ = v12 & new_n1150_;
  assign new_n1152_ = ~v10 & new_n1151_;
  assign new_n1153_ = v6 & new_n1152_;
  assign new_n1154_ = v5 & new_n1153_;
  assign new_n1155_ = ~v2 & new_n1154_;
  assign new_n1156_ = ~new_n1149_ & ~new_n1155_;
  assign new_n1157_ = ~v14 & ~new_n1156_;
  assign new_n1158_ = v13 & v14;
  assign new_n1159_ = v12 & new_n1158_;
  assign new_n1160_ = ~v12 & ~v13;
  assign new_n1161_ = ~new_n1159_ & ~new_n1160_;
  assign new_n1162_ = ~v15 & ~new_n1161_;
  assign new_n1163_ = v8 & new_n1162_;
  assign new_n1164_ = v1 & new_n1163_;
  assign new_n1165_ = new_n102_ & new_n1160_;
  assign new_n1166_ = ~new_n1164_ & ~new_n1165_;
  assign new_n1167_ = ~v6 & ~new_n1166_;
  assign new_n1168_ = ~v7 & new_n699_;
  assign new_n1169_ = ~v13 & new_n102_;
  assign new_n1170_ = new_n1168_ & new_n1169_;
  assign new_n1171_ = ~new_n1167_ & ~new_n1170_;
  assign new_n1172_ = ~v10 & ~new_n1171_;
  assign new_n1173_ = v5 & new_n1172_;
  assign new_n1174_ = ~new_n1157_ & ~new_n1173_;
  assign new_n1175_ = ~v0 & ~new_n1174_;
  assign new_n1176_ = ~v13 & ~new_n112_;
  assign new_n1177_ = v7 & new_n1176_;
  assign new_n1178_ = v6 & new_n1177_;
  assign new_n1179_ = v5 & new_n1178_;
  assign new_n1180_ = ~v9 & v13;
  assign new_n1181_ = new_n38_ & new_n1180_;
  assign new_n1182_ = new_n268_ & new_n1181_;
  assign new_n1183_ = ~new_n1179_ & ~new_n1182_;
  assign new_n1184_ = v8 & ~new_n1183_;
  assign new_n1185_ = new_n119_ & new_n1004_;
  assign new_n1186_ = v9 & v13;
  assign new_n1187_ = new_n102_ & new_n1186_;
  assign new_n1188_ = new_n1185_ & new_n1187_;
  assign new_n1189_ = ~new_n1184_ & ~new_n1188_;
  assign new_n1190_ = ~v12 & ~new_n1189_;
  assign new_n1191_ = ~v10 & new_n1190_;
  assign new_n1192_ = ~new_n1175_ & ~new_n1191_;
  assign new_n1193_ = v11 & ~new_n1192_;
  assign new_n1194_ = v4 & new_n1193_;
  assign \v16.10  = new_n1138_ | new_n1194_;
  assign new_n1196_ = v12 & ~new_n931_;
  assign new_n1197_ = ~new_n54_ & ~new_n1196_;
  assign new_n1198_ = ~v13 & ~new_n1197_;
  assign new_n1199_ = new_n44_ & new_n185_;
  assign new_n1200_ = ~v7 & ~new_n501_;
  assign new_n1201_ = v8 & ~new_n1200_;
  assign new_n1202_ = ~new_n1199_ & ~new_n1201_;
  assign new_n1203_ = ~v14 & ~new_n1202_;
  assign new_n1204_ = ~v4 & new_n1203_;
  assign new_n1205_ = ~v14 & ~new_n1204_;
  assign new_n1206_ = v15 & ~new_n1205_;
  assign new_n1207_ = ~new_n191_ & ~new_n1206_;
  assign new_n1208_ = v12 & ~new_n1207_;
  assign new_n1209_ = new_n712_ & ~new_n1208_;
  assign new_n1210_ = v13 & ~new_n1209_;
  assign new_n1211_ = ~new_n1198_ & ~new_n1210_;
  assign new_n1212_ = v10 & ~new_n1211_;
  assign new_n1213_ = v15 & ~new_n260_;
  assign new_n1214_ = v12 & new_n1213_;
  assign new_n1215_ = v6 & new_n1214_;
  assign new_n1216_ = ~new_n321_ & ~new_n1215_;
  assign new_n1217_ = ~v13 & ~new_n1216_;
  assign new_n1218_ = v4 & new_n1059_;
  assign new_n1219_ = ~new_n1217_ & ~new_n1218_;
  assign new_n1220_ = ~v14 & ~new_n1219_;
  assign new_n1221_ = v12 & ~v13;
  assign new_n1222_ = ~new_n224_ & ~new_n1221_;
  assign new_n1223_ = ~v4 & ~new_n1222_;
  assign new_n1224_ = v4 & ~v12;
  assign new_n1225_ = v13 & new_n191_;
  assign new_n1226_ = new_n1224_ & new_n1225_;
  assign new_n1227_ = ~new_n1223_ & ~new_n1226_;
  assign new_n1228_ = ~new_n1220_ & new_n1227_;
  assign new_n1229_ = ~v10 & ~new_n1228_;
  assign new_n1230_ = ~new_n1212_ & ~new_n1229_;
  assign new_n1231_ = ~v11 & ~new_n1230_;
  assign new_n1232_ = ~v0 & new_n539_;
  assign new_n1233_ = v12 & v13;
  assign new_n1234_ = new_n365_ & new_n1233_;
  assign new_n1235_ = new_n1232_ & new_n1234_;
  assign new_n1236_ = ~new_n1160_ & ~new_n1235_;
  assign new_n1237_ = ~v4 & ~new_n1236_;
  assign new_n1238_ = ~v13 & ~new_n540_;
  assign new_n1239_ = ~v12 & new_n1238_;
  assign new_n1240_ = ~new_n1237_ & ~new_n1239_;
  assign new_n1241_ = v14 & ~new_n1240_;
  assign new_n1242_ = ~v5 & v12;
  assign new_n1243_ = new_n786_ & new_n1242_;
  assign new_n1244_ = ~new_n1241_ & ~new_n1243_;
  assign new_n1245_ = ~v15 & ~new_n1244_;
  assign new_n1246_ = v13 & new_n38_;
  assign new_n1247_ = new_n1242_ & new_n1246_;
  assign new_n1248_ = ~new_n1245_ & ~new_n1247_;
  assign new_n1249_ = ~v10 & ~new_n1248_;
  assign new_n1250_ = ~v13 & ~v14;
  assign new_n1251_ = v12 & new_n1250_;
  assign new_n1252_ = ~v0 & new_n1251_;
  assign new_n1253_ = v13 & new_n102_;
  assign new_n1254_ = new_n486_ & new_n1253_;
  assign new_n1255_ = ~new_n1252_ & ~new_n1254_;
  assign new_n1256_ = v10 & ~new_n1255_;
  assign new_n1257_ = v9 & new_n1256_;
  assign new_n1258_ = ~v8 & new_n1257_;
  assign new_n1259_ = ~v6 & new_n1258_;
  assign new_n1260_ = ~v5 & new_n1259_;
  assign new_n1261_ = v4 & new_n1260_;
  assign new_n1262_ = ~new_n1249_ & ~new_n1261_;
  assign new_n1263_ = v11 & ~new_n1262_;
  assign \v16.11  = new_n1231_ | new_n1263_;
  assign new_n1265_ = ~v2 & new_n1233_;
  assign new_n1266_ = ~new_n1075_ & ~new_n1265_;
  assign new_n1267_ = ~new_n142_ & ~new_n1266_;
  assign new_n1268_ = v12 & new_n1075_;
  assign new_n1269_ = ~new_n1267_ & ~new_n1268_;
  assign new_n1270_ = v6 & ~new_n1269_;
  assign new_n1271_ = ~v13 & new_n492_;
  assign new_n1272_ = ~v12 & new_n1271_;
  assign new_n1273_ = ~new_n1270_ & ~new_n1272_;
  assign new_n1274_ = ~v4 & ~new_n1273_;
  assign new_n1275_ = v6 & new_n329_;
  assign new_n1276_ = ~v1 & new_n1275_;
  assign new_n1277_ = v8 & new_n224_;
  assign new_n1278_ = ~new_n1276_ & ~new_n1277_;
  assign new_n1279_ = ~v7 & ~new_n1278_;
  assign new_n1280_ = ~v6 & new_n224_;
  assign new_n1281_ = ~new_n1279_ & ~new_n1280_;
  assign new_n1282_ = ~v13 & ~new_n1281_;
  assign new_n1283_ = v4 & new_n1282_;
  assign new_n1284_ = ~new_n1274_ & ~new_n1283_;
  assign new_n1285_ = ~v10 & ~new_n1284_;
  assign new_n1286_ = ~v13 & ~new_n298_;
  assign new_n1287_ = ~v12 & new_n1286_;
  assign new_n1288_ = v10 & new_n1287_;
  assign new_n1289_ = ~new_n1285_ & ~new_n1288_;
  assign new_n1290_ = v5 & ~new_n1289_;
  assign new_n1291_ = v7 & v9;
  assign new_n1292_ = v4 & new_n1291_;
  assign new_n1293_ = ~new_n502_ & ~new_n1292_;
  assign new_n1294_ = v12 & ~new_n1293_;
  assign new_n1295_ = ~v5 & new_n1294_;
  assign new_n1296_ = ~new_n507_ & ~new_n1295_;
  assign new_n1297_ = ~v13 & ~new_n1296_;
  assign new_n1298_ = v10 & new_n1297_;
  assign new_n1299_ = ~v8 & new_n1298_;
  assign new_n1300_ = ~v6 & new_n1299_;
  assign new_n1301_ = ~new_n1290_ & ~new_n1300_;
  assign new_n1302_ = ~v0 & ~new_n1301_;
  assign new_n1303_ = v13 & v15;
  assign new_n1304_ = ~v9 & new_n1303_;
  assign new_n1305_ = new_n268_ & new_n1304_;
  assign new_n1306_ = ~v13 & ~v15;
  assign new_n1307_ = v7 & new_n1306_;
  assign new_n1308_ = new_n689_ & new_n1307_;
  assign new_n1309_ = ~new_n1305_ & ~new_n1308_;
  assign new_n1310_ = ~v12 & ~new_n1309_;
  assign new_n1311_ = new_n185_ & new_n321_;
  assign new_n1312_ = new_n121_ & new_n1306_;
  assign new_n1313_ = new_n1311_ & new_n1312_;
  assign new_n1314_ = ~new_n1310_ & ~new_n1313_;
  assign new_n1315_ = ~v10 & ~new_n1314_;
  assign new_n1316_ = v5 & new_n59_;
  assign new_n1317_ = v10 & new_n1160_;
  assign new_n1318_ = new_n1316_ & new_n1317_;
  assign new_n1319_ = ~new_n1315_ & ~new_n1318_;
  assign new_n1320_ = v8 & ~new_n1319_;
  assign new_n1321_ = ~v5 & ~v10;
  assign new_n1322_ = v13 & ~v15;
  assign new_n1323_ = v12 & new_n1322_;
  assign new_n1324_ = new_n1321_ & new_n1323_;
  assign new_n1325_ = ~new_n1320_ & ~new_n1324_;
  assign new_n1326_ = ~new_n1302_ & new_n1325_;
  assign new_n1327_ = v11 & ~new_n1326_;
  assign new_n1328_ = v12 & ~new_n627_;
  assign new_n1329_ = ~new_n321_ & ~new_n1328_;
  assign new_n1330_ = ~v10 & ~new_n1329_;
  assign new_n1331_ = v7 & new_n635_;
  assign new_n1332_ = ~v6 & new_n1331_;
  assign new_n1333_ = ~v5 & new_n1332_;
  assign new_n1334_ = ~v0 & new_n329_;
  assign new_n1335_ = ~new_n1333_ & ~new_n1334_;
  assign new_n1336_ = v10 & ~new_n1335_;
  assign new_n1337_ = ~new_n1330_ & ~new_n1336_;
  assign new_n1338_ = ~v13 & ~new_n1337_;
  assign new_n1339_ = v7 & new_n159_;
  assign new_n1340_ = ~new_n161_ & ~new_n1339_;
  assign new_n1341_ = v15 & ~new_n1340_;
  assign new_n1342_ = v12 & new_n1341_;
  assign new_n1343_ = ~v4 & new_n1342_;
  assign new_n1344_ = new_n329_ & ~new_n1343_;
  assign new_n1345_ = v10 & ~new_n1344_;
  assign new_n1346_ = new_n337_ & new_n412_;
  assign new_n1347_ = ~new_n1345_ & ~new_n1346_;
  assign new_n1348_ = v13 & ~new_n1347_;
  assign new_n1349_ = ~new_n1338_ & ~new_n1348_;
  assign new_n1350_ = ~v11 & ~new_n1349_;
  assign new_n1351_ = ~new_n1327_ & ~new_n1350_;
  assign new_n1352_ = ~v14 & ~new_n1351_;
  assign new_n1353_ = v4 & new_n1160_;
  assign new_n1354_ = new_n664_ & new_n1158_;
  assign new_n1355_ = ~new_n1353_ & ~new_n1354_;
  assign new_n1356_ = ~v15 & ~new_n1355_;
  assign new_n1357_ = v8 & new_n1356_;
  assign new_n1358_ = v1 & new_n1357_;
  assign new_n1359_ = ~v12 & new_n1169_;
  assign new_n1360_ = ~new_n1358_ & ~new_n1359_;
  assign new_n1361_ = ~v6 & ~new_n1360_;
  assign new_n1362_ = v4 & ~v7;
  assign new_n1363_ = v4 & ~new_n1362_;
  assign new_n1364_ = v15 & ~new_n1363_;
  assign new_n1365_ = v14 & new_n1364_;
  assign new_n1366_ = ~v13 & new_n1365_;
  assign new_n1367_ = ~v12 & new_n1366_;
  assign new_n1368_ = v8 & new_n1367_;
  assign new_n1369_ = ~new_n1361_ & ~new_n1368_;
  assign new_n1370_ = ~v0 & ~new_n1369_;
  assign new_n1371_ = v8 & new_n1359_;
  assign new_n1372_ = v7 & new_n1371_;
  assign new_n1373_ = v6 & new_n1372_;
  assign new_n1374_ = ~new_n1370_ & ~new_n1373_;
  assign new_n1375_ = v5 & ~new_n1374_;
  assign new_n1376_ = new_n44_ & new_n1303_;
  assign new_n1377_ = new_n858_ & new_n1376_;
  assign new_n1378_ = ~new_n1306_ & ~new_n1377_;
  assign new_n1379_ = ~v5 & ~new_n1378_;
  assign new_n1380_ = new_n364_ & new_n365_;
  assign new_n1381_ = ~v15 & ~new_n1380_;
  assign new_n1382_ = ~v13 & new_n1381_;
  assign new_n1383_ = ~new_n1379_ & ~new_n1382_;
  assign new_n1384_ = v14 & ~new_n1383_;
  assign new_n1385_ = ~v12 & new_n1384_;
  assign new_n1386_ = ~new_n1375_ & ~new_n1385_;
  assign new_n1387_ = ~v10 & ~new_n1386_;
  assign new_n1388_ = v5 & ~new_n521_;
  assign new_n1389_ = ~v7 & new_n525_;
  assign new_n1390_ = ~v6 & new_n1389_;
  assign new_n1391_ = ~new_n1388_ & ~new_n1390_;
  assign new_n1392_ = ~v0 & ~new_n1391_;
  assign new_n1393_ = v7 & ~v15;
  assign new_n1394_ = new_n689_ & new_n1393_;
  assign new_n1395_ = ~new_n1392_ & ~new_n1394_;
  assign new_n1396_ = ~v13 & ~new_n1395_;
  assign new_n1397_ = v10 & new_n1396_;
  assign new_n1398_ = new_n44_ & new_n1253_;
  assign new_n1399_ = new_n1311_ & new_n1398_;
  assign new_n1400_ = ~new_n1397_ & ~new_n1399_;
  assign new_n1401_ = ~v12 & ~new_n1400_;
  assign new_n1402_ = ~new_n1387_ & ~new_n1401_;
  assign new_n1403_ = v11 & ~new_n1402_;
  assign new_n1404_ = new_n1224_ & new_n1253_;
  assign new_n1405_ = ~new_n1223_ & ~new_n1404_;
  assign new_n1406_ = ~v10 & ~new_n1405_;
  assign new_n1407_ = v10 & new_n1079_;
  assign new_n1408_ = ~new_n1406_ & ~new_n1407_;
  assign new_n1409_ = ~v11 & ~new_n1408_;
  assign new_n1410_ = ~new_n1403_ & ~new_n1409_;
  assign \v16.12  = new_n1352_ | ~new_n1410_;
  assign new_n1412_ = v4 & new_n44_;
  assign new_n1413_ = ~new_n469_ & ~new_n1412_;
  assign new_n1414_ = ~new_n43_ & ~new_n1413_;
  assign new_n1415_ = ~v14 & new_n1414_;
  assign new_n1416_ = ~v12 & new_n1415_;
  assign new_n1417_ = v7 & new_n1416_;
  assign new_n1418_ = ~v6 & new_n1417_;
  assign new_n1419_ = ~v5 & new_n1418_;
  assign new_n1420_ = ~new_n1196_ & ~new_n1419_;
  assign new_n1421_ = v10 & ~new_n1420_;
  assign new_n1422_ = ~new_n191_ & ~new_n1085_;
  assign new_n1423_ = v4 & ~new_n1422_;
  assign new_n1424_ = v4 & ~new_n1423_;
  assign new_n1425_ = v12 & ~new_n1424_;
  assign new_n1426_ = ~v4 & new_n134_;
  assign new_n1427_ = ~new_n1425_ & ~new_n1426_;
  assign new_n1428_ = ~v10 & ~new_n1427_;
  assign new_n1429_ = ~new_n1421_ & ~new_n1428_;
  assign new_n1430_ = ~v11 & ~new_n1429_;
  assign new_n1431_ = v4 & ~v9;
  assign new_n1432_ = v4 & ~new_n1431_;
  assign new_n1433_ = ~new_n142_ & ~new_n1432_;
  assign new_n1434_ = ~new_n664_ & ~new_n1433_;
  assign new_n1435_ = v15 & ~new_n1434_;
  assign new_n1436_ = v6 & new_n1435_;
  assign new_n1437_ = ~new_n494_ & ~new_n1436_;
  assign new_n1438_ = ~v14 & ~new_n1437_;
  assign new_n1439_ = ~v12 & new_n515_;
  assign new_n1440_ = ~v4 & new_n1439_;
  assign new_n1441_ = ~new_n1438_ & ~new_n1440_;
  assign new_n1442_ = ~v0 & ~new_n1441_;
  assign new_n1443_ = ~v4 & new_n116_;
  assign new_n1444_ = ~new_n1442_ & ~new_n1443_;
  assign new_n1445_ = v5 & ~new_n1444_;
  assign new_n1446_ = ~new_n550_ & ~new_n1445_;
  assign new_n1447_ = ~v10 & ~new_n1446_;
  assign new_n1448_ = ~v14 & ~new_n1293_;
  assign new_n1449_ = v12 & new_n1448_;
  assign new_n1450_ = v10 & new_n1449_;
  assign new_n1451_ = ~v8 & new_n1450_;
  assign new_n1452_ = ~v6 & new_n1451_;
  assign new_n1453_ = ~v5 & new_n1452_;
  assign new_n1454_ = ~v0 & new_n1453_;
  assign new_n1455_ = ~new_n1447_ & ~new_n1454_;
  assign new_n1456_ = v11 & ~new_n1455_;
  assign new_n1457_ = ~new_n1430_ & ~new_n1456_;
  assign new_n1458_ = ~v13 & ~new_n1457_;
  assign new_n1459_ = v6 & new_n1433_;
  assign new_n1460_ = v5 & new_n1459_;
  assign new_n1461_ = ~v2 & new_n1460_;
  assign new_n1462_ = ~v0 & new_n1461_;
  assign new_n1463_ = ~v5 & v15;
  assign new_n1464_ = ~new_n1462_ & ~new_n1463_;
  assign new_n1465_ = v12 & ~new_n1464_;
  assign new_n1466_ = new_n159_ & new_n412_;
  assign new_n1467_ = new_n1311_ & new_n1466_;
  assign new_n1468_ = ~new_n1465_ & ~new_n1467_;
  assign new_n1469_ = ~v14 & ~new_n1468_;
  assign new_n1470_ = v5 & ~v6;
  assign new_n1471_ = v4 & new_n1470_;
  assign new_n1472_ = new_n417_ & new_n1471_;
  assign new_n1473_ = new_n159_ & new_n996_;
  assign new_n1474_ = new_n1472_ & new_n1473_;
  assign new_n1475_ = ~new_n1469_ & ~new_n1474_;
  assign new_n1476_ = ~v10 & ~new_n1475_;
  assign new_n1477_ = ~v12 & new_n102_;
  assign new_n1478_ = new_n44_ & new_n1477_;
  assign new_n1479_ = new_n1311_ & new_n1478_;
  assign new_n1480_ = ~new_n1476_ & ~new_n1479_;
  assign new_n1481_ = v11 & ~new_n1480_;
  assign new_n1482_ = v14 & ~new_n798_;
  assign new_n1483_ = v10 & ~new_n1482_;
  assign new_n1484_ = ~new_n427_ & ~new_n1483_;
  assign new_n1485_ = ~v15 & ~new_n1484_;
  assign new_n1486_ = ~v4 & v7;
  assign new_n1487_ = new_n890_ & new_n1486_;
  assign new_n1488_ = ~v14 & ~new_n1487_;
  assign new_n1489_ = v15 & ~new_n1488_;
  assign new_n1490_ = v12 & new_n1489_;
  assign new_n1491_ = ~v12 & ~v14;
  assign new_n1492_ = ~new_n1490_ & ~new_n1491_;
  assign new_n1493_ = v10 & ~new_n1492_;
  assign new_n1494_ = ~new_n1485_ & ~new_n1493_;
  assign new_n1495_ = ~v11 & ~new_n1494_;
  assign new_n1496_ = ~new_n1481_ & ~new_n1495_;
  assign new_n1497_ = v13 & ~new_n1496_;
  assign new_n1498_ = ~new_n226_ & ~new_n1497_;
  assign \v16.13  = new_n1458_ | ~new_n1498_;
  assign new_n1500_ = ~v0 & v4;
  assign new_n1501_ = new_n689_ & new_n1500_;
  assign new_n1502_ = v12 & new_n38_;
  assign new_n1503_ = new_n501_ & new_n1502_;
  assign new_n1504_ = new_n1501_ & new_n1503_;
  assign new_n1505_ = ~v12 & new_n191_;
  assign new_n1506_ = ~new_n1504_ & ~new_n1505_;
  assign new_n1507_ = ~v1 & ~new_n1506_;
  assign new_n1508_ = ~v0 & ~v6;
  assign new_n1509_ = ~new_n300_ & ~new_n1508_;
  assign new_n1510_ = v8 & ~new_n1363_;
  assign new_n1511_ = ~v0 & new_n1510_;
  assign new_n1512_ = new_n1509_ & ~new_n1511_;
  assign new_n1513_ = ~new_n112_ & ~new_n1512_;
  assign new_n1514_ = ~v0 & new_n364_;
  assign new_n1515_ = new_n517_ & new_n1514_;
  assign new_n1516_ = ~new_n1513_ & ~new_n1515_;
  assign new_n1517_ = ~v12 & ~new_n1516_;
  assign new_n1518_ = ~new_n378_ & ~new_n664_;
  assign new_n1519_ = v15 & ~new_n1518_;
  assign new_n1520_ = ~v14 & new_n1519_;
  assign new_n1521_ = v6 & new_n1520_;
  assign new_n1522_ = ~v0 & new_n1521_;
  assign new_n1523_ = ~new_n1517_ & ~new_n1522_;
  assign new_n1524_ = v5 & ~new_n1523_;
  assign new_n1525_ = v14 & ~new_n365_;
  assign new_n1526_ = ~v12 & new_n1525_;
  assign new_n1527_ = ~new_n861_ & ~new_n1526_;
  assign new_n1528_ = ~new_n857_ & new_n1527_;
  assign new_n1529_ = ~v15 & ~new_n1528_;
  assign new_n1530_ = ~new_n1524_ & ~new_n1529_;
  assign new_n1531_ = ~new_n1507_ & new_n1530_;
  assign new_n1532_ = ~v13 & ~new_n1531_;
  assign new_n1533_ = ~new_n230_ & ~new_n597_;
  assign new_n1534_ = v5 & new_n1533_;
  assign new_n1535_ = ~v0 & new_n1534_;
  assign new_n1536_ = ~v5 & new_n38_;
  assign new_n1537_ = ~new_n1535_ & ~new_n1536_;
  assign new_n1538_ = v12 & ~new_n1537_;
  assign new_n1539_ = ~new_n899_ & ~new_n1538_;
  assign new_n1540_ = v13 & ~new_n1539_;
  assign new_n1541_ = ~new_n1532_ & ~new_n1540_;
  assign new_n1542_ = v11 & ~new_n1541_;
  assign new_n1543_ = ~v14 & ~new_n624_;
  assign new_n1544_ = ~new_n342_ & ~new_n1543_;
  assign new_n1545_ = v15 & ~new_n1544_;
  assign new_n1546_ = v4 & new_n191_;
  assign new_n1547_ = ~new_n1545_ & ~new_n1546_;
  assign new_n1548_ = v12 & ~new_n1547_;
  assign new_n1549_ = ~new_n463_ & ~new_n1548_;
  assign new_n1550_ = ~v13 & ~new_n1549_;
  assign new_n1551_ = v14 & ~new_n102_;
  assign new_n1552_ = v13 & ~new_n1551_;
  assign new_n1553_ = v4 & new_n1552_;
  assign new_n1554_ = ~new_n444_ & ~new_n1553_;
  assign new_n1555_ = ~v12 & ~new_n1554_;
  assign new_n1556_ = ~new_n1550_ & ~new_n1555_;
  assign new_n1557_ = ~v11 & ~new_n1556_;
  assign new_n1558_ = ~new_n1542_ & ~new_n1557_;
  assign new_n1559_ = ~v10 & ~new_n1558_;
  assign new_n1560_ = new_n44_ & new_n327_;
  assign new_n1561_ = ~v4 & new_n159_;
  assign new_n1562_ = new_n1502_ & new_n1561_;
  assign new_n1563_ = ~new_n1560_ & ~new_n1562_;
  assign new_n1564_ = v7 & ~new_n1563_;
  assign new_n1565_ = ~v4 & new_n161_;
  assign new_n1566_ = ~v4 & ~new_n1565_;
  assign new_n1567_ = ~v14 & ~new_n1566_;
  assign new_n1568_ = ~v14 & ~new_n1567_;
  assign new_n1569_ = v15 & ~new_n1568_;
  assign new_n1570_ = ~new_n191_ & ~new_n1569_;
  assign new_n1571_ = v12 & ~new_n1570_;
  assign new_n1572_ = v14 & ~new_n882_;
  assign new_n1573_ = ~v12 & ~new_n1572_;
  assign new_n1574_ = ~new_n35_ & ~new_n1573_;
  assign new_n1575_ = ~new_n1571_ & new_n1574_;
  assign new_n1576_ = ~new_n1564_ & new_n1575_;
  assign new_n1577_ = v13 & ~new_n1576_;
  assign new_n1578_ = v9 & new_n1064_;
  assign new_n1579_ = v7 & new_n1578_;
  assign new_n1580_ = ~v6 & new_n1579_;
  assign new_n1581_ = ~v5 & new_n1580_;
  assign new_n1582_ = v4 & new_n1581_;
  assign new_n1583_ = ~new_n52_ & ~new_n1582_;
  assign new_n1584_ = ~v12 & ~new_n1583_;
  assign new_n1585_ = ~new_n794_ & ~new_n1584_;
  assign new_n1586_ = ~v13 & ~new_n1585_;
  assign new_n1587_ = ~new_n1577_ & ~new_n1586_;
  assign new_n1588_ = ~v11 & ~new_n1587_;
  assign new_n1589_ = ~v9 & ~v15;
  assign new_n1590_ = ~v9 & ~new_n1589_;
  assign new_n1591_ = v7 & ~new_n1590_;
  assign new_n1592_ = ~new_n254_ & ~new_n1591_;
  assign new_n1593_ = v4 & ~new_n1592_;
  assign new_n1594_ = ~new_n502_ & ~new_n1593_;
  assign new_n1595_ = ~v14 & ~new_n1594_;
  assign new_n1596_ = ~v13 & new_n1595_;
  assign new_n1597_ = v12 & new_n1596_;
  assign new_n1598_ = v11 & new_n1597_;
  assign new_n1599_ = ~v8 & new_n1598_;
  assign new_n1600_ = ~v6 & new_n1599_;
  assign new_n1601_ = ~v5 & new_n1600_;
  assign new_n1602_ = ~v0 & new_n1601_;
  assign new_n1603_ = ~new_n1588_ & ~new_n1602_;
  assign new_n1604_ = v10 & ~new_n1603_;
  assign new_n1605_ = ~v6 & new_n1004_;
  assign new_n1606_ = new_n321_ & new_n1605_;
  assign new_n1607_ = v11 & ~v12;
  assign new_n1608_ = v9 & new_n1607_;
  assign new_n1609_ = new_n1253_ & new_n1608_;
  assign new_n1610_ = new_n1606_ & new_n1609_;
  assign new_n1611_ = ~new_n1604_ & ~new_n1610_;
  assign \v16.14  = new_n1559_ | ~new_n1611_;
  assign new_n1613_ = v12 & ~new_n1422_;
  assign new_n1614_ = v12 & ~new_n1613_;
  assign new_n1615_ = v4 & ~new_n1614_;
  assign new_n1616_ = ~new_n463_ & ~new_n1615_;
  assign new_n1617_ = ~v10 & ~new_n1616_;
  assign new_n1618_ = ~new_n43_ & ~new_n310_;
  assign new_n1619_ = ~v14 & new_n1618_;
  assign new_n1620_ = v7 & new_n1619_;
  assign new_n1621_ = ~v6 & new_n1620_;
  assign new_n1622_ = ~v5 & new_n1621_;
  assign new_n1623_ = v4 & new_n1622_;
  assign new_n1624_ = ~new_n52_ & ~new_n1623_;
  assign new_n1625_ = ~v12 & ~new_n1624_;
  assign new_n1626_ = ~new_n798_ & ~new_n1625_;
  assign new_n1627_ = v10 & ~new_n1626_;
  assign new_n1628_ = ~new_n1617_ & ~new_n1627_;
  assign new_n1629_ = ~new_n336_ & new_n1628_;
  assign new_n1630_ = ~v11 & ~new_n1629_;
  assign new_n1631_ = v6 & v9;
  assign new_n1632_ = new_n38_ & new_n1631_;
  assign new_n1633_ = new_n224_ & new_n365_;
  assign new_n1634_ = ~new_n1632_ & ~new_n1633_;
  assign new_n1635_ = v1 & ~new_n1634_;
  assign new_n1636_ = v15 & ~new_n92_;
  assign new_n1637_ = v9 & new_n1636_;
  assign new_n1638_ = v6 & new_n1637_;
  assign new_n1639_ = ~new_n99_ & ~new_n1638_;
  assign new_n1640_ = ~v14 & ~new_n1639_;
  assign new_n1641_ = v15 & ~new_n97_;
  assign new_n1642_ = v14 & new_n1641_;
  assign new_n1643_ = ~v12 & new_n1642_;
  assign new_n1644_ = ~new_n1640_ & ~new_n1643_;
  assign new_n1645_ = ~new_n1635_ & new_n1644_;
  assign new_n1646_ = ~v10 & ~new_n1645_;
  assign new_n1647_ = v4 & new_n1646_;
  assign new_n1648_ = ~new_n675_ & ~new_n1647_;
  assign new_n1649_ = v5 & ~new_n1648_;
  assign new_n1650_ = v4 & ~new_n503_;
  assign new_n1651_ = v12 & ~new_n1650_;
  assign new_n1652_ = v9 & new_n1651_;
  assign new_n1653_ = ~v5 & new_n1652_;
  assign new_n1654_ = ~new_n507_ & ~new_n1653_;
  assign new_n1655_ = ~v14 & ~new_n1654_;
  assign new_n1656_ = ~v8 & new_n1655_;
  assign new_n1657_ = ~new_n681_ & ~new_n1656_;
  assign new_n1658_ = v10 & ~new_n1657_;
  assign new_n1659_ = ~v6 & new_n1658_;
  assign new_n1660_ = ~new_n1649_ & ~new_n1659_;
  assign new_n1661_ = ~v0 & ~new_n1660_;
  assign new_n1662_ = ~v10 & ~new_n112_;
  assign new_n1663_ = v4 & new_n1662_;
  assign new_n1664_ = v10 & ~v14;
  assign new_n1665_ = ~new_n1663_ & ~new_n1664_;
  assign new_n1666_ = v8 & ~new_n1665_;
  assign new_n1667_ = ~new_n305_ & ~new_n1666_;
  assign new_n1668_ = ~v12 & ~new_n1667_;
  assign new_n1669_ = v7 & new_n1668_;
  assign new_n1670_ = v6 & new_n1669_;
  assign new_n1671_ = v5 & new_n1670_;
  assign new_n1672_ = ~new_n1661_ & ~new_n1671_;
  assign new_n1673_ = v11 & ~new_n1672_;
  assign new_n1674_ = ~new_n1630_ & ~new_n1673_;
  assign new_n1675_ = ~v13 & ~new_n1674_;
  assign new_n1676_ = v11 & ~new_n597_;
  assign new_n1677_ = ~v10 & new_n1676_;
  assign new_n1678_ = v9 & new_n1677_;
  assign new_n1679_ = v5 & new_n1678_;
  assign new_n1680_ = ~v0 & new_n1679_;
  assign new_n1681_ = new_n38_ & new_n178_;
  assign new_n1682_ = ~new_n1680_ & ~new_n1681_;
  assign new_n1683_ = v4 & ~new_n1682_;
  assign new_n1684_ = v8 & ~new_n853_;
  assign new_n1685_ = v7 & ~new_n1684_;
  assign new_n1686_ = ~v7 & new_n159_;
  assign new_n1687_ = ~new_n1685_ & ~new_n1686_;
  assign new_n1688_ = ~v14 & ~new_n1687_;
  assign new_n1689_ = ~v4 & new_n1688_;
  assign new_n1690_ = ~v14 & ~new_n1689_;
  assign new_n1691_ = v15 & ~new_n1690_;
  assign new_n1692_ = ~new_n191_ & ~new_n1691_;
  assign new_n1693_ = ~v11 & ~new_n1692_;
  assign new_n1694_ = v10 & new_n1693_;
  assign new_n1695_ = new_n188_ & new_n1321_;
  assign new_n1696_ = ~new_n1694_ & ~new_n1695_;
  assign new_n1697_ = ~new_n1683_ & new_n1696_;
  assign new_n1698_ = v12 & ~new_n1697_;
  assign new_n1699_ = new_n196_ & new_n268_;
  assign new_n1700_ = v11 & ~new_n1699_;
  assign new_n1701_ = v14 & ~new_n1700_;
  assign new_n1702_ = v4 & new_n1701_;
  assign new_n1703_ = v5 & ~v11;
  assign new_n1704_ = ~new_n1702_ & ~new_n1703_;
  assign new_n1705_ = v15 & ~new_n1704_;
  assign new_n1706_ = ~v10 & new_n1705_;
  assign new_n1707_ = v10 & new_n207_;
  assign new_n1708_ = ~new_n1706_ & ~new_n1707_;
  assign new_n1709_ = ~v12 & ~new_n1708_;
  assign new_n1710_ = ~new_n219_ & ~new_n1709_;
  assign new_n1711_ = ~new_n1698_ & new_n1710_;
  assign new_n1712_ = v13 & ~new_n1711_;
  assign new_n1713_ = ~new_n448_ & ~new_n1712_;
  assign \v16.15  = new_n1675_ | ~new_n1713_;
  assign new_n1715_ = v4 & new_n159_;
  assign new_n1716_ = ~new_n469_ & ~new_n1715_;
  assign new_n1717_ = ~new_n43_ & ~new_n1716_;
  assign new_n1718_ = ~v14 & new_n1717_;
  assign new_n1719_ = v7 & new_n1718_;
  assign new_n1720_ = ~v6 & new_n1719_;
  assign new_n1721_ = ~v5 & new_n1720_;
  assign new_n1722_ = ~new_n52_ & ~new_n1721_;
  assign new_n1723_ = ~v12 & ~new_n1722_;
  assign new_n1724_ = ~new_n42_ & ~new_n1723_;
  assign new_n1725_ = ~v11 & ~new_n1724_;
  assign new_n1726_ = ~v9 & v15;
  assign new_n1727_ = v7 & new_n1726_;
  assign new_n1728_ = ~new_n254_ & ~new_n1727_;
  assign new_n1729_ = v4 & ~new_n1728_;
  assign new_n1730_ = ~new_n502_ & ~new_n1729_;
  assign new_n1731_ = v12 & ~new_n1730_;
  assign new_n1732_ = ~v5 & new_n1731_;
  assign new_n1733_ = ~new_n507_ & ~new_n1732_;
  assign new_n1734_ = ~v8 & ~new_n1733_;
  assign new_n1735_ = v5 & ~v12;
  assign new_n1736_ = ~new_n1734_ & ~new_n1735_;
  assign new_n1737_ = ~v14 & ~new_n1736_;
  assign new_n1738_ = v5 & v8;
  assign new_n1739_ = ~new_n1389_ & ~new_n1738_;
  assign new_n1740_ = ~v12 & ~new_n1739_;
  assign new_n1741_ = ~new_n1737_ & ~new_n1740_;
  assign new_n1742_ = ~v6 & ~new_n1741_;
  assign new_n1743_ = v5 & new_n553_;
  assign new_n1744_ = ~new_n1742_ & ~new_n1743_;
  assign new_n1745_ = ~v0 & ~new_n1744_;
  assign new_n1746_ = v7 & new_n553_;
  assign new_n1747_ = v6 & new_n1746_;
  assign new_n1748_ = v5 & new_n1747_;
  assign new_n1749_ = ~new_n1745_ & ~new_n1748_;
  assign new_n1750_ = v11 & ~new_n1749_;
  assign new_n1751_ = ~new_n1725_ & ~new_n1750_;
  assign new_n1752_ = v10 & ~new_n1751_;
  assign new_n1753_ = v6 & ~v11;
  assign new_n1754_ = new_n1502_ & new_n1753_;
  assign new_n1755_ = new_n191_ & new_n1607_;
  assign new_n1756_ = ~new_n1754_ & ~new_n1755_;
  assign new_n1757_ = ~v1 & ~new_n1756_;
  assign new_n1758_ = ~v14 & ~new_n301_;
  assign new_n1759_ = v5 & new_n1758_;
  assign new_n1760_ = ~v14 & ~new_n1759_;
  assign new_n1761_ = ~v4 & ~new_n1760_;
  assign new_n1762_ = v14 & ~new_n366_;
  assign new_n1763_ = ~new_n1761_ & ~new_n1762_;
  assign new_n1764_ = ~v12 & ~new_n1763_;
  assign new_n1765_ = v9 & new_n456_;
  assign new_n1766_ = v8 & new_n1765_;
  assign new_n1767_ = ~v7 & new_n1766_;
  assign new_n1768_ = ~v6 & new_n1767_;
  assign new_n1769_ = ~v5 & new_n1768_;
  assign new_n1770_ = ~new_n1764_ & ~new_n1769_;
  assign new_n1771_ = ~v15 & ~new_n1770_;
  assign new_n1772_ = v8 & new_n327_;
  assign new_n1773_ = ~v0 & ~v14;
  assign new_n1774_ = ~new_n1772_ & ~new_n1773_;
  assign new_n1775_ = v7 & ~new_n1774_;
  assign new_n1776_ = ~v1 & ~v12;
  assign new_n1777_ = ~v14 & ~new_n1776_;
  assign new_n1778_ = ~v0 & new_n1777_;
  assign new_n1779_ = ~new_n1775_ & ~new_n1778_;
  assign new_n1780_ = v6 & ~new_n1779_;
  assign new_n1781_ = v14 & ~new_n298_;
  assign new_n1782_ = ~v12 & new_n1781_;
  assign new_n1783_ = ~v0 & new_n1782_;
  assign new_n1784_ = ~new_n1780_ & ~new_n1783_;
  assign new_n1785_ = v15 & ~new_n1784_;
  assign new_n1786_ = v5 & new_n1785_;
  assign new_n1787_ = ~v4 & new_n1786_;
  assign new_n1788_ = ~new_n1771_ & ~new_n1787_;
  assign new_n1789_ = v11 & ~new_n1788_;
  assign new_n1790_ = v15 & ~new_n941_;
  assign new_n1791_ = ~v14 & ~new_n1790_;
  assign new_n1792_ = ~new_n102_ & ~new_n1791_;
  assign new_n1793_ = v12 & ~new_n1792_;
  assign new_n1794_ = v4 & new_n1793_;
  assign new_n1795_ = ~new_n463_ & ~new_n1794_;
  assign new_n1796_ = ~v11 & ~new_n1795_;
  assign new_n1797_ = ~new_n1789_ & ~new_n1796_;
  assign new_n1798_ = ~new_n1757_ & new_n1797_;
  assign new_n1799_ = ~v10 & ~new_n1798_;
  assign new_n1800_ = ~new_n1752_ & ~new_n1799_;
  assign new_n1801_ = ~v13 & ~new_n1800_;
  assign new_n1802_ = v5 & new_n598_;
  assign new_n1803_ = ~v0 & new_n1802_;
  assign new_n1804_ = ~v9 & ~v12;
  assign new_n1805_ = new_n38_ & new_n1804_;
  assign new_n1806_ = new_n120_ & new_n1805_;
  assign new_n1807_ = ~new_n1803_ & ~new_n1806_;
  assign new_n1808_ = ~v4 & ~new_n1807_;
  assign new_n1809_ = new_n858_ & new_n1466_;
  assign new_n1810_ = ~new_n421_ & ~new_n1809_;
  assign new_n1811_ = ~v14 & ~new_n1810_;
  assign new_n1812_ = ~v5 & new_n1811_;
  assign new_n1813_ = ~new_n1808_ & ~new_n1812_;
  assign new_n1814_ = v11 & ~new_n1813_;
  assign new_n1815_ = ~v14 & ~new_n38_;
  assign new_n1816_ = ~v12 & ~new_n1815_;
  assign new_n1817_ = ~v11 & new_n1816_;
  assign new_n1818_ = v4 & new_n1817_;
  assign new_n1819_ = ~new_n1814_ & ~new_n1818_;
  assign new_n1820_ = ~v10 & ~new_n1819_;
  assign new_n1821_ = v11 & new_n904_;
  assign new_n1822_ = ~v7 & new_n1821_;
  assign new_n1823_ = ~v6 & new_n1822_;
  assign new_n1824_ = ~v5 & new_n1823_;
  assign new_n1825_ = v7 & new_n178_;
  assign new_n1826_ = ~new_n1824_ & ~new_n1825_;
  assign new_n1827_ = v9 & ~new_n1826_;
  assign new_n1828_ = ~v8 & new_n1827_;
  assign new_n1829_ = new_n203_ & new_n242_;
  assign new_n1830_ = ~new_n1828_ & ~new_n1829_;
  assign new_n1831_ = ~v12 & ~new_n1830_;
  assign new_n1832_ = v10 & new_n1038_;
  assign new_n1833_ = ~new_n1831_ & ~new_n1832_;
  assign new_n1834_ = v14 & ~new_n1833_;
  assign new_n1835_ = v15 & ~new_n160_;
  assign new_n1836_ = v12 & new_n1835_;
  assign new_n1837_ = ~v7 & new_n1836_;
  assign new_n1838_ = ~v4 & new_n1837_;
  assign new_n1839_ = new_n329_ & ~new_n1838_;
  assign new_n1840_ = ~v14 & ~new_n1839_;
  assign new_n1841_ = ~v11 & new_n1840_;
  assign new_n1842_ = v10 & new_n1841_;
  assign new_n1843_ = ~new_n1834_ & ~new_n1842_;
  assign new_n1844_ = ~new_n1820_ & new_n1843_;
  assign new_n1845_ = v13 & ~new_n1844_;
  assign new_n1846_ = ~new_n226_ & ~new_n1845_;
  assign \v16.16  = new_n1801_ | ~new_n1846_;
endmodule


