// Benchmark "c2670.blif" written by ABC on Fri Feb 25 15:12:55 2022

module c2670  ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
    G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
    G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
    G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
    G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
    G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
    G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136,
    G137, G138, G139, G140, G141, G142, \IN-G169 , \IN-G174 , \IN-G177 ,
    \IN-G178 , \IN-G179 , \IN-G180 , \IN-G181 , \IN-G182 , \IN-G183 ,
    \IN-G184 , \IN-G185 , \IN-G186 , \IN-G189 , \IN-G190 , \IN-G191 ,
    \IN-G192 , \IN-G193 , \IN-G194 , \IN-G195 , \IN-G196 , \IN-G197 ,
    \IN-G198 , \IN-G199 , \IN-G200 , \IN-G201 , \IN-G202 , \IN-G203 ,
    \IN-G204 , \IN-G205 , \IN-G206 , \IN-G207 , \IN-G208 , \IN-G209 ,
    \IN-G210 , \IN-G211 , \IN-G212 , \IN-G213 , \IN-G214 , \IN-G215 ,
    \IN-G239 , \IN-G240 , \IN-G241 , \IN-G242 , \IN-G243 , \IN-G244 ,
    \IN-G245 , \IN-G246 , \IN-G247 , \IN-G248 , \IN-G249 , \IN-G250 ,
    \IN-G251 , \IN-G252 , \IN-G253 , \IN-G254 , \IN-G255 , \IN-G256 ,
    \IN-G257 , \IN-G262 , \IN-G263 , \IN-G264 , \IN-G265 , \IN-G266 ,
    \IN-G267 , \IN-G268 , \IN-G269 , \IN-G270 , \IN-G271 , \IN-G272 ,
    \IN-G273 , \IN-G274 , \IN-G275 , \IN-G276 , \IN-G277 , \IN-G278 ,
    \IN-G279 , G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083,
    G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986,
    G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100,
    G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451,
    G2454, G2474, G2678,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G350, G335, G409, G369, G367, G411, G337, G384,
    G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173,
    G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171,
    G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
    G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145,
    G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20,
    G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36,
    G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74,
    G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90,
    G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105,
    G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
    G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135,
    G136, G137, G138, G139, G140, G141, G142, \IN-G169 , \IN-G174 ,
    \IN-G177 , \IN-G178 , \IN-G179 , \IN-G180 , \IN-G181 , \IN-G182 ,
    \IN-G183 , \IN-G184 , \IN-G185 , \IN-G186 , \IN-G189 , \IN-G190 ,
    \IN-G191 , \IN-G192 , \IN-G193 , \IN-G194 , \IN-G195 , \IN-G196 ,
    \IN-G197 , \IN-G198 , \IN-G199 , \IN-G200 , \IN-G201 , \IN-G202 ,
    \IN-G203 , \IN-G204 , \IN-G205 , \IN-G206 , \IN-G207 , \IN-G208 ,
    \IN-G209 , \IN-G210 , \IN-G211 , \IN-G212 , \IN-G213 , \IN-G214 ,
    \IN-G215 , \IN-G239 , \IN-G240 , \IN-G241 , \IN-G242 , \IN-G243 ,
    \IN-G244 , \IN-G245 , \IN-G246 , \IN-G247 , \IN-G248 , \IN-G249 ,
    \IN-G250 , \IN-G251 , \IN-G252 , \IN-G253 , \IN-G254 , \IN-G255 ,
    \IN-G256 , \IN-G257 , \IN-G262 , \IN-G263 , \IN-G264 , \IN-G265 ,
    \IN-G266 , \IN-G267 , \IN-G268 , \IN-G269 , \IN-G270 , \IN-G271 ,
    \IN-G272 , \IN-G273 , \IN-G274 , \IN-G275 , \IN-G276 , \IN-G277 ,
    \IN-G278 , \IN-G279 , G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185,
    G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199,
    G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211,
    G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
    G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262,
    G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274,
    G275, G276, G277, G278, G279, G350, G335, G409, G369, G367, G411, G337,
    G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391,
    G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168,
    G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284,
    G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
    G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire new_n375_, new_n376_, new_n378_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n391_, new_n392_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n473_,
    new_n474_, new_n476_, new_n477_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n536_, new_n537_, new_n539_, new_n540_, new_n541_,
    new_n543_, new_n544_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_;
  assign new_n375_ = G2084 & G2090;
  assign new_n376_ = G2078 & new_n375_;
  assign G158 = ~G2072 | ~new_n376_;
  assign new_n378_ = G2 & G15;
  assign G259 = ~G661 | ~new_n378_;
  assign G173 = G94 & G452;
  assign G223 = ~G7 | ~G661;
  assign G234 = ~G567 | G223;
  assign G217 = ~G2106 | G223;
  assign new_n384_ = G57 & G120;
  assign new_n385_ = G108 & new_n384_;
  assign new_n386_ = G69 & new_n385_;
  assign new_n387_ = G82 & G132;
  assign new_n388_ = G96 & new_n387_;
  assign new_n389_ = G44 & new_n388_;
  assign G325 = new_n386_ & new_n389_;
  assign new_n391_ = G2106 & ~new_n389_;
  assign new_n392_ = G567 & ~new_n386_;
  assign G319 = ~new_n391_ & ~new_n392_;
  assign new_n394_ = G137 & ~G2104;
  assign new_n395_ = ~G2105 & new_n394_;
  assign new_n396_ = G101 & G2104;
  assign new_n397_ = ~G2105 & new_n396_;
  assign new_n398_ = G125 & ~G2104;
  assign new_n399_ = G2105 & new_n398_;
  assign new_n400_ = G113 & G2104;
  assign new_n401_ = G2105 & new_n400_;
  assign new_n402_ = ~new_n395_ & ~new_n397_;
  assign new_n403_ = ~new_n399_ & ~new_n401_;
  assign G160 = new_n402_ & new_n403_;
  assign new_n405_ = G136 & ~G2104;
  assign new_n406_ = ~G2105 & new_n405_;
  assign new_n407_ = G100 & G2104;
  assign new_n408_ = ~G2105 & new_n407_;
  assign new_n409_ = G124 & ~G2104;
  assign new_n410_ = G2105 & new_n409_;
  assign new_n411_ = G112 & G2104;
  assign new_n412_ = G2105 & new_n411_;
  assign new_n413_ = ~new_n406_ & ~new_n408_;
  assign new_n414_ = ~new_n410_ & ~new_n412_;
  assign G162 = new_n413_ & new_n414_;
  assign new_n416_ = G138 & ~G2104;
  assign new_n417_ = ~G2105 & new_n416_;
  assign new_n418_ = G102 & G2104;
  assign new_n419_ = ~G2105 & new_n418_;
  assign new_n420_ = G126 & ~G2104;
  assign new_n421_ = G2105 & new_n420_;
  assign new_n422_ = G114 & G2104;
  assign new_n423_ = G2105 & new_n422_;
  assign new_n424_ = ~new_n417_ & ~new_n419_;
  assign new_n425_ = ~new_n421_ & ~new_n423_;
  assign G164 = new_n424_ & new_n425_;
  assign new_n427_ = G88 & ~G543;
  assign new_n428_ = ~G651 & new_n427_;
  assign new_n429_ = G50 & G543;
  assign new_n430_ = ~G651 & new_n429_;
  assign new_n431_ = G62 & ~G543;
  assign new_n432_ = G651 & new_n431_;
  assign new_n433_ = G75 & G543;
  assign new_n434_ = G651 & new_n433_;
  assign new_n435_ = ~new_n428_ & ~new_n430_;
  assign new_n436_ = ~new_n432_ & ~new_n434_;
  assign G166 = new_n435_ & new_n436_;
  assign new_n438_ = G89 & ~G543;
  assign new_n439_ = ~G651 & new_n438_;
  assign new_n440_ = G51 & G543;
  assign new_n441_ = ~G651 & new_n440_;
  assign new_n442_ = G63 & ~G543;
  assign new_n443_ = G651 & new_n442_;
  assign new_n444_ = G76 & G543;
  assign new_n445_ = G651 & new_n444_;
  assign new_n446_ = ~new_n439_ & ~new_n441_;
  assign new_n447_ = ~new_n443_ & ~new_n445_;
  assign G168 = new_n446_ & new_n447_;
  assign new_n449_ = G90 & ~G543;
  assign new_n450_ = ~G651 & new_n449_;
  assign new_n451_ = G52 & G543;
  assign new_n452_ = ~G651 & new_n451_;
  assign new_n453_ = G64 & ~G543;
  assign new_n454_ = G651 & new_n453_;
  assign new_n455_ = G77 & G543;
  assign new_n456_ = G651 & new_n455_;
  assign new_n457_ = ~new_n450_ & ~new_n452_;
  assign new_n458_ = ~new_n454_ & ~new_n456_;
  assign G171 = new_n457_ & new_n458_;
  assign new_n460_ = G81 & ~G543;
  assign new_n461_ = ~G651 & new_n460_;
  assign new_n462_ = G43 & G543;
  assign new_n463_ = ~G651 & new_n462_;
  assign new_n464_ = G56 & ~G543;
  assign new_n465_ = G651 & new_n464_;
  assign new_n466_ = G68 & G543;
  assign new_n467_ = G651 & new_n466_;
  assign new_n468_ = ~new_n461_ & ~new_n463_;
  assign new_n469_ = ~new_n465_ & ~new_n467_;
  assign new_n470_ = new_n468_ & new_n469_;
  assign new_n471_ = G860 & ~new_n470_;
  assign G153 = ~G860 | new_n471_;
  assign new_n473_ = G483 & G661;
  assign new_n474_ = G36 & new_n473_;
  assign G176 = ~G319 | ~new_n474_;
  assign new_n476_ = G1 & G3;
  assign new_n477_ = G319 & new_n473_;
  assign G188 = new_n476_ | ~new_n477_;
  assign new_n479_ = G91 & ~G543;
  assign new_n480_ = ~G651 & new_n479_;
  assign new_n481_ = G53 & G543;
  assign new_n482_ = ~G651 & new_n481_;
  assign new_n483_ = G65 & ~G543;
  assign new_n484_ = G651 & new_n483_;
  assign new_n485_ = G78 & G543;
  assign new_n486_ = G651 & new_n485_;
  assign new_n487_ = ~new_n480_ & ~new_n482_;
  assign new_n488_ = ~new_n484_ & ~new_n486_;
  assign G299 = ~new_n487_ | ~new_n488_;
  assign new_n490_ = G87 & ~G543;
  assign new_n491_ = ~G651 & new_n490_;
  assign new_n492_ = G49 & G543;
  assign new_n493_ = ~G651 & new_n492_;
  assign new_n494_ = ~G543 & G651;
  assign new_n495_ = G74 & G543;
  assign new_n496_ = G651 & new_n495_;
  assign new_n497_ = ~new_n491_ & ~new_n493_;
  assign new_n498_ = ~new_n494_ & ~new_n496_;
  assign G288 = ~new_n497_ | ~new_n498_;
  assign new_n500_ = G86 & ~G543;
  assign new_n501_ = ~G651 & new_n500_;
  assign new_n502_ = G48 & G543;
  assign new_n503_ = ~G651 & new_n502_;
  assign new_n504_ = G61 & ~G543;
  assign new_n505_ = G651 & new_n504_;
  assign new_n506_ = G73 & G543;
  assign new_n507_ = G651 & new_n506_;
  assign new_n508_ = ~new_n501_ & ~new_n503_;
  assign new_n509_ = ~new_n505_ & ~new_n507_;
  assign G305 = ~new_n508_ | ~new_n509_;
  assign new_n511_ = G85 & ~G543;
  assign new_n512_ = ~G651 & new_n511_;
  assign new_n513_ = G47 & G543;
  assign new_n514_ = ~G651 & new_n513_;
  assign new_n515_ = G60 & ~G543;
  assign new_n516_ = G651 & new_n515_;
  assign new_n517_ = G72 & G543;
  assign new_n518_ = G651 & new_n517_;
  assign new_n519_ = ~new_n512_ & ~new_n514_;
  assign new_n520_ = ~new_n516_ & ~new_n518_;
  assign G290 = ~new_n519_ | ~new_n520_;
  assign new_n522_ = G92 & ~G543;
  assign new_n523_ = ~G651 & new_n522_;
  assign new_n524_ = G54 & G543;
  assign new_n525_ = ~G651 & new_n524_;
  assign new_n526_ = G66 & ~G543;
  assign new_n527_ = G651 & new_n526_;
  assign new_n528_ = G79 & G543;
  assign new_n529_ = G651 & new_n528_;
  assign new_n530_ = ~new_n523_ & ~new_n525_;
  assign new_n531_ = ~new_n527_ & ~new_n529_;
  assign new_n532_ = new_n530_ & new_n531_;
  assign new_n533_ = ~G868 & ~new_n532_;
  assign new_n534_ = G868 & ~G171;
  assign G284 = new_n533_ | new_n534_;
  assign new_n536_ = ~G868 & G299;
  assign new_n537_ = G868 & ~G168;
  assign G297 = new_n536_ | new_n537_;
  assign new_n539_ = ~G559 & new_n532_;
  assign new_n540_ = ~G860 & ~new_n539_;
  assign new_n541_ = G860 & ~new_n532_;
  assign G148 = new_n540_ | new_n541_;
  assign new_n543_ = ~G868 & ~new_n470_;
  assign new_n544_ = G868 & ~new_n539_;
  assign G282 = new_n543_ | new_n544_;
  assign new_n546_ = ~G2104 & ~G2105;
  assign new_n547_ = G2104 & ~G2105;
  assign new_n548_ = ~G2104 & G2105;
  assign new_n549_ = G2104 & G2105;
  assign new_n550_ = ~new_n546_ & ~new_n547_;
  assign new_n551_ = ~new_n548_ & ~new_n549_;
  assign new_n552_ = new_n550_ & new_n551_;
  assign new_n553_ = ~G2100 & ~new_n552_;
  assign new_n554_ = ~G2100 & ~new_n553_;
  assign new_n555_ = ~new_n552_ & ~new_n553_;
  assign new_n556_ = ~new_n554_ & ~new_n555_;
  assign new_n557_ = G135 & ~G2104;
  assign new_n558_ = ~G2105 & new_n557_;
  assign new_n559_ = G99 & G2104;
  assign new_n560_ = ~G2105 & new_n559_;
  assign new_n561_ = G123 & ~G2104;
  assign new_n562_ = G2105 & new_n561_;
  assign new_n563_ = G111 & G2104;
  assign new_n564_ = G2105 & new_n563_;
  assign new_n565_ = ~new_n558_ & ~new_n560_;
  assign new_n566_ = ~new_n562_ & ~new_n564_;
  assign new_n567_ = new_n565_ & new_n566_;
  assign new_n568_ = ~G2096 & ~new_n567_;
  assign new_n569_ = ~G2096 & ~new_n568_;
  assign new_n570_ = ~new_n567_ & ~new_n568_;
  assign new_n571_ = ~new_n569_ & ~new_n570_;
  assign G156 = ~new_n556_ | ~new_n571_;
  assign new_n573_ = ~G2451 & G2454;
  assign new_n574_ = G2451 & ~G2454;
  assign new_n575_ = ~new_n573_ & ~new_n574_;
  assign new_n576_ = G1341 & ~G1348;
  assign new_n577_ = ~G1341 & G1348;
  assign new_n578_ = ~new_n576_ & ~new_n577_;
  assign new_n579_ = ~new_n575_ & new_n578_;
  assign new_n580_ = new_n575_ & ~new_n578_;
  assign new_n581_ = ~new_n579_ & ~new_n580_;
  assign new_n582_ = ~G2427 & G2430;
  assign new_n583_ = G2427 & ~G2430;
  assign new_n584_ = ~new_n582_ & ~new_n583_;
  assign new_n585_ = ~G2435 & G2438;
  assign new_n586_ = G2435 & ~G2438;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = ~G2443 & G2446;
  assign new_n589_ = G2443 & ~G2446;
  assign new_n590_ = ~new_n588_ & ~new_n589_;
  assign new_n591_ = ~new_n584_ & new_n587_;
  assign new_n592_ = new_n590_ & new_n591_;
  assign new_n593_ = new_n584_ & new_n587_;
  assign new_n594_ = ~new_n590_ & new_n593_;
  assign new_n595_ = ~new_n592_ & ~new_n594_;
  assign new_n596_ = new_n584_ & ~new_n587_;
  assign new_n597_ = new_n590_ & new_n596_;
  assign new_n598_ = ~new_n584_ & ~new_n587_;
  assign new_n599_ = ~new_n590_ & new_n598_;
  assign new_n600_ = ~new_n597_ & ~new_n599_;
  assign new_n601_ = new_n595_ & new_n600_;
  assign new_n602_ = ~new_n581_ & new_n601_;
  assign new_n603_ = new_n581_ & ~new_n601_;
  assign new_n604_ = ~new_n602_ & ~new_n603_;
  assign G401 = G14 & new_n604_;
  assign new_n606_ = G2096 & ~G2100;
  assign new_n607_ = ~G2096 & G2100;
  assign new_n608_ = ~new_n606_ & ~new_n607_;
  assign new_n609_ = ~G2067 & G2678;
  assign new_n610_ = G2067 & ~G2678;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign new_n612_ = G2072 & ~G2078;
  assign new_n613_ = ~G2072 & G2078;
  assign new_n614_ = ~new_n612_ & ~new_n613_;
  assign new_n615_ = G2084 & ~G2090;
  assign new_n616_ = ~G2084 & G2090;
  assign new_n617_ = ~new_n615_ & ~new_n616_;
  assign new_n618_ = ~new_n611_ & new_n614_;
  assign new_n619_ = new_n617_ & new_n618_;
  assign new_n620_ = new_n611_ & new_n614_;
  assign new_n621_ = ~new_n617_ & new_n620_;
  assign new_n622_ = ~new_n619_ & ~new_n621_;
  assign new_n623_ = new_n611_ & ~new_n614_;
  assign new_n624_ = new_n617_ & new_n623_;
  assign new_n625_ = ~new_n611_ & ~new_n614_;
  assign new_n626_ = ~new_n617_ & new_n625_;
  assign new_n627_ = ~new_n624_ & ~new_n626_;
  assign new_n628_ = new_n622_ & new_n627_;
  assign new_n629_ = ~new_n608_ & new_n628_;
  assign new_n630_ = new_n608_ & ~new_n628_;
  assign G227 = ~new_n629_ & ~new_n630_;
  assign new_n632_ = G1981 & ~G1986;
  assign new_n633_ = ~G1981 & G1986;
  assign new_n634_ = ~new_n632_ & ~new_n633_;
  assign new_n635_ = G1991 & ~G1996;
  assign new_n636_ = ~G1991 & G1996;
  assign new_n637_ = ~new_n635_ & ~new_n636_;
  assign new_n638_ = ~new_n634_ & new_n637_;
  assign new_n639_ = new_n634_ & ~new_n637_;
  assign new_n640_ = ~new_n638_ & ~new_n639_;
  assign new_n641_ = ~G1956 & G2474;
  assign new_n642_ = G1956 & ~G2474;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign new_n644_ = G1961 & ~G1966;
  assign new_n645_ = ~G1961 & G1966;
  assign new_n646_ = ~new_n644_ & ~new_n645_;
  assign new_n647_ = G1971 & ~G1976;
  assign new_n648_ = ~G1971 & G1976;
  assign new_n649_ = ~new_n647_ & ~new_n648_;
  assign new_n650_ = ~new_n643_ & new_n646_;
  assign new_n651_ = new_n649_ & new_n650_;
  assign new_n652_ = new_n643_ & new_n646_;
  assign new_n653_ = ~new_n649_ & new_n652_;
  assign new_n654_ = ~new_n651_ & ~new_n653_;
  assign new_n655_ = new_n643_ & ~new_n646_;
  assign new_n656_ = new_n649_ & new_n655_;
  assign new_n657_ = ~new_n643_ & ~new_n646_;
  assign new_n658_ = ~new_n649_ & new_n657_;
  assign new_n659_ = ~new_n656_ & ~new_n658_;
  assign new_n660_ = new_n654_ & new_n659_;
  assign new_n661_ = ~new_n640_ & new_n660_;
  assign new_n662_ = new_n640_ & ~new_n660_;
  assign G229 = ~new_n661_ & ~new_n662_;
  assign new_n664_ = G25 & ~G29;
  assign new_n665_ = G131 & ~G2104;
  assign new_n666_ = ~G2105 & new_n665_;
  assign new_n667_ = G95 & G2104;
  assign new_n668_ = ~G2105 & new_n667_;
  assign new_n669_ = G119 & ~G2104;
  assign new_n670_ = G2105 & new_n669_;
  assign new_n671_ = G107 & G2104;
  assign new_n672_ = G2105 & new_n671_;
  assign new_n673_ = ~new_n666_ & ~new_n668_;
  assign new_n674_ = ~new_n670_ & ~new_n672_;
  assign new_n675_ = new_n673_ & new_n674_;
  assign new_n676_ = G29 & ~new_n675_;
  assign new_n677_ = ~new_n664_ & ~new_n676_;
  assign new_n678_ = G1991 & ~new_n677_;
  assign new_n679_ = ~G1991 & new_n677_;
  assign new_n680_ = ~new_n678_ & ~new_n679_;
  assign new_n681_ = ~G16 & G24;
  assign new_n682_ = G16 & G290;
  assign new_n683_ = ~new_n681_ & ~new_n682_;
  assign new_n684_ = G1986 & ~new_n683_;
  assign new_n685_ = ~G1986 & new_n683_;
  assign new_n686_ = ~new_n684_ & ~new_n685_;
  assign new_n687_ = G6 & ~G16;
  assign new_n688_ = G16 & G305;
  assign new_n689_ = ~new_n687_ & ~new_n688_;
  assign new_n690_ = G1981 & ~new_n689_;
  assign new_n691_ = ~G1981 & new_n689_;
  assign new_n692_ = ~new_n690_ & ~new_n691_;
  assign new_n693_ = ~G16 & G23;
  assign new_n694_ = G16 & G288;
  assign new_n695_ = ~new_n693_ & ~new_n694_;
  assign new_n696_ = G1976 & ~new_n695_;
  assign new_n697_ = ~G1976 & new_n695_;
  assign new_n698_ = ~new_n696_ & ~new_n697_;
  assign new_n699_ = ~G16 & G22;
  assign new_n700_ = G16 & ~G166;
  assign new_n701_ = ~new_n699_ & ~new_n700_;
  assign new_n702_ = G1971 & ~new_n701_;
  assign new_n703_ = ~G1971 & new_n701_;
  assign new_n704_ = ~new_n702_ & ~new_n703_;
  assign new_n705_ = new_n680_ & new_n686_;
  assign new_n706_ = new_n692_ & new_n705_;
  assign new_n707_ = new_n698_ & new_n706_;
  assign new_n708_ = new_n704_ & new_n707_;
  assign new_n709_ = ~G16 & G21;
  assign new_n710_ = G16 & ~G168;
  assign new_n711_ = ~new_n709_ & ~new_n710_;
  assign new_n712_ = G1966 & ~new_n711_;
  assign new_n713_ = ~G1966 & new_n711_;
  assign new_n714_ = ~new_n712_ & ~new_n713_;
  assign new_n715_ = G5 & ~G16;
  assign new_n716_ = G16 & ~G171;
  assign new_n717_ = ~new_n715_ & ~new_n716_;
  assign new_n718_ = G1961 & ~new_n717_;
  assign new_n719_ = ~G1961 & new_n717_;
  assign new_n720_ = ~new_n718_ & ~new_n719_;
  assign new_n721_ = ~G16 & G20;
  assign new_n722_ = G16 & G299;
  assign new_n723_ = ~new_n721_ & ~new_n722_;
  assign new_n724_ = G1956 & ~new_n723_;
  assign new_n725_ = ~G1956 & new_n723_;
  assign new_n726_ = ~new_n724_ & ~new_n725_;
  assign new_n727_ = G4 & ~G16;
  assign new_n728_ = G16 & ~new_n532_;
  assign new_n729_ = ~new_n727_ & ~new_n728_;
  assign new_n730_ = G1348 & ~new_n729_;
  assign new_n731_ = ~G1348 & new_n729_;
  assign new_n732_ = ~new_n730_ & ~new_n731_;
  assign new_n733_ = ~G16 & G19;
  assign new_n734_ = G16 & ~new_n470_;
  assign new_n735_ = ~new_n733_ & ~new_n734_;
  assign new_n736_ = G1341 & ~new_n735_;
  assign new_n737_ = ~G1341 & new_n735_;
  assign new_n738_ = ~new_n736_ & ~new_n737_;
  assign new_n739_ = new_n714_ & new_n720_;
  assign new_n740_ = new_n726_ & new_n739_;
  assign new_n741_ = new_n732_ & new_n740_;
  assign new_n742_ = new_n738_ & new_n741_;
  assign new_n743_ = new_n708_ & new_n742_;
  assign new_n744_ = G28 & ~G29;
  assign new_n745_ = G29 & ~new_n567_;
  assign new_n746_ = ~new_n744_ & ~new_n745_;
  assign new_n747_ = ~G29 & G35;
  assign new_n748_ = G29 & ~G162;
  assign new_n749_ = ~new_n747_ & ~new_n748_;
  assign new_n750_ = G2090 & ~new_n749_;
  assign new_n751_ = ~G2090 & new_n749_;
  assign new_n752_ = ~new_n750_ & ~new_n751_;
  assign new_n753_ = ~new_n746_ & new_n752_;
  assign new_n754_ = ~G29 & G34;
  assign new_n755_ = G29 & ~G160;
  assign new_n756_ = ~new_n754_ & ~new_n755_;
  assign new_n757_ = G2084 & ~new_n756_;
  assign new_n758_ = ~G2084 & new_n756_;
  assign new_n759_ = ~new_n757_ & ~new_n758_;
  assign new_n760_ = G27 & ~G29;
  assign new_n761_ = G29 & ~G164;
  assign new_n762_ = ~new_n760_ & ~new_n761_;
  assign new_n763_ = G2078 & ~new_n762_;
  assign new_n764_ = ~G2078 & new_n762_;
  assign new_n765_ = ~new_n763_ & ~new_n764_;
  assign new_n766_ = ~G29 & G33;
  assign new_n767_ = G139 & ~G2104;
  assign new_n768_ = ~G2105 & new_n767_;
  assign new_n769_ = G103 & G2104;
  assign new_n770_ = ~G2105 & new_n769_;
  assign new_n771_ = G127 & ~G2104;
  assign new_n772_ = G2105 & new_n771_;
  assign new_n773_ = G115 & G2104;
  assign new_n774_ = G2105 & new_n773_;
  assign new_n775_ = ~new_n768_ & ~new_n770_;
  assign new_n776_ = ~new_n772_ & ~new_n774_;
  assign new_n777_ = new_n775_ & new_n776_;
  assign new_n778_ = G29 & ~new_n777_;
  assign new_n779_ = ~new_n766_ & ~new_n778_;
  assign new_n780_ = G2072 & ~new_n779_;
  assign new_n781_ = ~G2072 & new_n779_;
  assign new_n782_ = ~new_n780_ & ~new_n781_;
  assign new_n783_ = G26 & ~G29;
  assign new_n784_ = G140 & ~G2104;
  assign new_n785_ = ~G2105 & new_n784_;
  assign new_n786_ = G104 & G2104;
  assign new_n787_ = ~G2105 & new_n786_;
  assign new_n788_ = G128 & ~G2104;
  assign new_n789_ = G2105 & new_n788_;
  assign new_n790_ = G116 & G2104;
  assign new_n791_ = G2105 & new_n790_;
  assign new_n792_ = ~new_n785_ & ~new_n787_;
  assign new_n793_ = ~new_n789_ & ~new_n791_;
  assign new_n794_ = new_n792_ & new_n793_;
  assign new_n795_ = G29 & ~new_n794_;
  assign new_n796_ = ~new_n783_ & ~new_n795_;
  assign new_n797_ = G2067 & ~new_n796_;
  assign new_n798_ = ~G2067 & new_n796_;
  assign new_n799_ = ~new_n797_ & ~new_n798_;
  assign new_n800_ = ~G29 & G32;
  assign new_n801_ = G141 & ~G2104;
  assign new_n802_ = ~G2105 & new_n801_;
  assign new_n803_ = G105 & G2104;
  assign new_n804_ = ~G2105 & new_n803_;
  assign new_n805_ = G129 & ~G2104;
  assign new_n806_ = G2105 & new_n805_;
  assign new_n807_ = G117 & G2104;
  assign new_n808_ = G2105 & new_n807_;
  assign new_n809_ = ~new_n802_ & ~new_n804_;
  assign new_n810_ = ~new_n806_ & ~new_n808_;
  assign new_n811_ = new_n809_ & new_n810_;
  assign new_n812_ = G29 & ~new_n811_;
  assign new_n813_ = ~new_n800_ & ~new_n812_;
  assign new_n814_ = G1996 & ~new_n813_;
  assign new_n815_ = ~G1996 & new_n813_;
  assign new_n816_ = ~new_n814_ & ~new_n815_;
  assign new_n817_ = new_n759_ & new_n765_;
  assign new_n818_ = new_n782_ & new_n817_;
  assign new_n819_ = new_n799_ & new_n818_;
  assign new_n820_ = new_n816_ & new_n819_;
  assign new_n821_ = new_n753_ & new_n820_;
  assign new_n822_ = G11 & ~G868;
  assign new_n823_ = G11 & G868;
  assign new_n824_ = ~new_n822_ & ~new_n823_;
  assign new_n825_ = new_n743_ & new_n821_;
  assign G311 = ~new_n824_ & new_n825_;
  assign new_n827_ = ~new_n470_ & new_n532_;
  assign new_n828_ = new_n470_ & ~new_n532_;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign new_n830_ = ~new_n539_ & ~new_n829_;
  assign new_n831_ = new_n539_ & new_n829_;
  assign new_n832_ = ~new_n830_ & ~new_n831_;
  assign new_n833_ = G93 & ~G543;
  assign new_n834_ = ~G651 & new_n833_;
  assign new_n835_ = G55 & G543;
  assign new_n836_ = ~G651 & new_n835_;
  assign new_n837_ = G67 & ~G543;
  assign new_n838_ = G651 & new_n837_;
  assign new_n839_ = G80 & G543;
  assign new_n840_ = G651 & new_n839_;
  assign new_n841_ = ~new_n834_ & ~new_n836_;
  assign new_n842_ = ~new_n838_ & ~new_n840_;
  assign new_n843_ = new_n841_ & new_n842_;
  assign new_n844_ = ~new_n832_ & new_n843_;
  assign new_n845_ = new_n832_ & ~new_n843_;
  assign new_n846_ = ~new_n844_ & ~new_n845_;
  assign new_n847_ = ~G860 & ~new_n846_;
  assign new_n848_ = G860 & ~new_n843_;
  assign G145 = new_n847_ | new_n848_;
  assign new_n850_ = ~G160 & G162;
  assign new_n851_ = G160 & ~G162;
  assign new_n852_ = ~new_n850_ & ~new_n851_;
  assign new_n853_ = new_n552_ & ~new_n567_;
  assign new_n854_ = ~new_n552_ & new_n567_;
  assign new_n855_ = ~new_n853_ & ~new_n854_;
  assign new_n856_ = ~new_n852_ & new_n855_;
  assign new_n857_ = new_n852_ & ~new_n855_;
  assign new_n858_ = ~new_n856_ & ~new_n857_;
  assign new_n859_ = G142 & ~G2104;
  assign new_n860_ = ~G2105 & new_n859_;
  assign new_n861_ = G106 & G2104;
  assign new_n862_ = ~G2105 & new_n861_;
  assign new_n863_ = G130 & ~G2104;
  assign new_n864_ = G2105 & new_n863_;
  assign new_n865_ = G118 & G2104;
  assign new_n866_ = G2105 & new_n865_;
  assign new_n867_ = ~new_n860_ & ~new_n862_;
  assign new_n868_ = ~new_n864_ & ~new_n866_;
  assign new_n869_ = new_n867_ & new_n868_;
  assign new_n870_ = new_n675_ & ~new_n869_;
  assign new_n871_ = ~new_n675_ & new_n869_;
  assign new_n872_ = ~new_n870_ & ~new_n871_;
  assign new_n873_ = new_n794_ & ~new_n811_;
  assign new_n874_ = ~new_n794_ & new_n811_;
  assign new_n875_ = ~new_n873_ & ~new_n874_;
  assign new_n876_ = G164 & ~new_n777_;
  assign new_n877_ = ~G164 & new_n777_;
  assign new_n878_ = ~new_n876_ & ~new_n877_;
  assign new_n879_ = ~new_n872_ & new_n875_;
  assign new_n880_ = new_n878_ & new_n879_;
  assign new_n881_ = new_n872_ & new_n875_;
  assign new_n882_ = ~new_n878_ & new_n881_;
  assign new_n883_ = ~new_n880_ & ~new_n882_;
  assign new_n884_ = new_n872_ & ~new_n875_;
  assign new_n885_ = new_n878_ & new_n884_;
  assign new_n886_ = ~new_n872_ & ~new_n875_;
  assign new_n887_ = ~new_n878_ & new_n886_;
  assign new_n888_ = ~new_n885_ & ~new_n887_;
  assign new_n889_ = new_n883_ & new_n888_;
  assign new_n890_ = ~new_n858_ & new_n889_;
  assign new_n891_ = new_n858_ & ~new_n889_;
  assign new_n892_ = ~new_n890_ & ~new_n891_;
  assign G395 = ~G37 & new_n892_;
  assign new_n894_ = ~G868 & ~new_n843_;
  assign new_n895_ = G166 & G288;
  assign new_n896_ = ~G166 & ~G288;
  assign new_n897_ = ~new_n895_ & ~new_n896_;
  assign new_n898_ = ~G305 & G290;
  assign new_n899_ = G305 & ~G290;
  assign new_n900_ = ~new_n898_ & ~new_n899_;
  assign new_n901_ = ~new_n897_ & new_n900_;
  assign new_n902_ = new_n897_ & ~new_n900_;
  assign new_n903_ = ~new_n901_ & ~new_n902_;
  assign new_n904_ = ~new_n470_ & new_n843_;
  assign new_n905_ = new_n470_ & ~new_n843_;
  assign new_n906_ = ~new_n904_ & ~new_n905_;
  assign new_n907_ = G299 & new_n532_;
  assign new_n908_ = ~G299 & ~new_n532_;
  assign new_n909_ = ~new_n907_ & ~new_n908_;
  assign new_n910_ = ~new_n539_ & new_n906_;
  assign new_n911_ = new_n909_ & new_n910_;
  assign new_n912_ = new_n539_ & new_n906_;
  assign new_n913_ = ~new_n909_ & new_n912_;
  assign new_n914_ = ~new_n911_ & ~new_n913_;
  assign new_n915_ = new_n539_ & ~new_n906_;
  assign new_n916_ = new_n909_ & new_n915_;
  assign new_n917_ = ~new_n539_ & ~new_n906_;
  assign new_n918_ = ~new_n909_ & new_n917_;
  assign new_n919_ = ~new_n916_ & ~new_n918_;
  assign new_n920_ = new_n914_ & new_n919_;
  assign new_n921_ = ~new_n903_ & new_n920_;
  assign new_n922_ = new_n903_ & ~new_n920_;
  assign new_n923_ = ~new_n921_ & ~new_n922_;
  assign new_n924_ = G868 & ~new_n923_;
  assign G295 = new_n894_ | new_n924_;
  assign new_n926_ = ~G168 & G171;
  assign new_n927_ = G168 & ~G171;
  assign new_n928_ = ~new_n926_ & ~new_n927_;
  assign new_n929_ = ~new_n906_ & new_n909_;
  assign new_n930_ = new_n928_ & new_n929_;
  assign new_n931_ = new_n906_ & new_n909_;
  assign new_n932_ = ~new_n928_ & new_n931_;
  assign new_n933_ = ~new_n930_ & ~new_n932_;
  assign new_n934_ = new_n906_ & ~new_n909_;
  assign new_n935_ = new_n928_ & new_n934_;
  assign new_n936_ = ~new_n906_ & ~new_n909_;
  assign new_n937_ = ~new_n928_ & new_n936_;
  assign new_n938_ = ~new_n935_ & ~new_n937_;
  assign new_n939_ = new_n933_ & new_n938_;
  assign new_n940_ = ~new_n903_ & new_n939_;
  assign new_n941_ = new_n903_ & ~new_n939_;
  assign new_n942_ = ~new_n940_ & ~new_n941_;
  assign G397 = ~G37 & new_n942_;
  assign new_n944_ = ~G1384 & ~G164;
  assign new_n945_ = G160 & new_n944_;
  assign new_n946_ = G40 & new_n945_;
  assign new_n947_ = ~G2067 & ~new_n946_;
  assign new_n948_ = G40 & G160;
  assign new_n949_ = ~new_n944_ & new_n948_;
  assign new_n950_ = new_n947_ & new_n949_;
  assign new_n951_ = ~new_n794_ & ~new_n946_;
  assign new_n952_ = new_n949_ & new_n951_;
  assign new_n953_ = new_n950_ & ~new_n952_;
  assign new_n954_ = ~new_n950_ & ~new_n952_;
  assign new_n955_ = new_n950_ & new_n952_;
  assign new_n956_ = ~new_n954_ & ~new_n955_;
  assign new_n957_ = ~G1996 & ~new_n946_;
  assign new_n958_ = new_n949_ & new_n957_;
  assign new_n959_ = ~new_n811_ & ~new_n946_;
  assign new_n960_ = new_n949_ & new_n959_;
  assign new_n961_ = new_n958_ & ~new_n960_;
  assign new_n962_ = ~new_n956_ & new_n961_;
  assign new_n963_ = ~new_n958_ & ~new_n960_;
  assign new_n964_ = new_n958_ & new_n960_;
  assign new_n965_ = ~new_n963_ & ~new_n964_;
  assign new_n966_ = ~G1991 & ~new_n946_;
  assign new_n967_ = new_n949_ & new_n966_;
  assign new_n968_ = ~new_n675_ & ~new_n946_;
  assign new_n969_ = new_n949_ & new_n968_;
  assign new_n970_ = new_n967_ & ~new_n969_;
  assign new_n971_ = ~new_n956_ & ~new_n965_;
  assign new_n972_ = new_n970_ & new_n971_;
  assign new_n973_ = ~new_n967_ & ~new_n969_;
  assign new_n974_ = new_n967_ & new_n969_;
  assign new_n975_ = ~new_n973_ & ~new_n974_;
  assign new_n976_ = G290 & ~new_n946_;
  assign new_n977_ = new_n949_ & new_n976_;
  assign new_n978_ = ~G1986 & ~new_n946_;
  assign new_n979_ = new_n949_ & new_n978_;
  assign new_n980_ = ~new_n977_ & new_n979_;
  assign new_n981_ = ~new_n956_ & ~new_n975_;
  assign new_n982_ = new_n980_ & new_n981_;
  assign new_n983_ = ~new_n965_ & new_n982_;
  assign new_n984_ = ~new_n953_ & ~new_n962_;
  assign new_n985_ = ~new_n972_ & ~new_n983_;
  assign new_n986_ = new_n984_ & new_n985_;
  assign new_n987_ = ~G1981 & ~new_n946_;
  assign new_n988_ = G8 & new_n987_;
  assign new_n989_ = G305 & ~new_n946_;
  assign new_n990_ = G8 & new_n989_;
  assign new_n991_ = new_n988_ & ~new_n990_;
  assign new_n992_ = ~new_n988_ & ~new_n990_;
  assign new_n993_ = new_n988_ & new_n990_;
  assign new_n994_ = ~new_n992_ & ~new_n993_;
  assign new_n995_ = ~G1976 & ~new_n946_;
  assign new_n996_ = G8 & new_n995_;
  assign new_n997_ = G288 & ~new_n946_;
  assign new_n998_ = G8 & new_n997_;
  assign new_n999_ = new_n996_ & ~new_n998_;
  assign new_n1000_ = ~new_n994_ & new_n999_;
  assign new_n1001_ = ~new_n996_ & ~new_n998_;
  assign new_n1002_ = new_n996_ & new_n998_;
  assign new_n1003_ = ~new_n1001_ & ~new_n1002_;
  assign new_n1004_ = ~G2090 & new_n946_;
  assign new_n1005_ = ~G1971 & ~new_n946_;
  assign new_n1006_ = ~new_n1004_ & ~new_n1005_;
  assign new_n1007_ = G8 & ~new_n1006_;
  assign new_n1008_ = ~G166 & ~new_n946_;
  assign new_n1009_ = ~G166 & new_n946_;
  assign new_n1010_ = ~new_n1008_ & ~new_n1009_;
  assign new_n1011_ = G8 & ~new_n1010_;
  assign new_n1012_ = new_n1007_ & ~new_n1011_;
  assign new_n1013_ = ~new_n994_ & ~new_n1003_;
  assign new_n1014_ = new_n1012_ & new_n1013_;
  assign new_n1015_ = ~new_n1007_ & ~new_n1011_;
  assign new_n1016_ = new_n1007_ & new_n1011_;
  assign new_n1017_ = ~new_n1015_ & ~new_n1016_;
  assign new_n1018_ = ~G2084 & new_n946_;
  assign new_n1019_ = ~G1966 & ~new_n946_;
  assign new_n1020_ = ~new_n1018_ & ~new_n1019_;
  assign new_n1021_ = G8 & ~new_n1020_;
  assign new_n1022_ = ~G168 & ~new_n946_;
  assign new_n1023_ = ~G168 & new_n946_;
  assign new_n1024_ = ~new_n1022_ & ~new_n1023_;
  assign new_n1025_ = G8 & ~new_n1024_;
  assign new_n1026_ = new_n1021_ & ~new_n1025_;
  assign new_n1027_ = ~new_n994_ & ~new_n1017_;
  assign new_n1028_ = new_n1026_ & new_n1027_;
  assign new_n1029_ = ~new_n1003_ & new_n1028_;
  assign new_n1030_ = ~new_n1021_ & ~new_n1025_;
  assign new_n1031_ = new_n1021_ & new_n1025_;
  assign new_n1032_ = ~new_n1030_ & ~new_n1031_;
  assign new_n1033_ = ~G2078 & new_n946_;
  assign new_n1034_ = ~G1961 & ~new_n946_;
  assign new_n1035_ = ~new_n1033_ & ~new_n1034_;
  assign new_n1036_ = G171 & ~new_n1035_;
  assign new_n1037_ = ~new_n1017_ & ~new_n1032_;
  assign new_n1038_ = ~new_n994_ & new_n1037_;
  assign new_n1039_ = new_n1036_ & new_n1038_;
  assign new_n1040_ = ~new_n1003_ & new_n1039_;
  assign new_n1041_ = ~new_n991_ & ~new_n1000_;
  assign new_n1042_ = ~new_n1014_ & new_n1041_;
  assign new_n1043_ = ~new_n1029_ & ~new_n1040_;
  assign new_n1044_ = new_n1042_ & new_n1043_;
  assign new_n1045_ = G171 & new_n1035_;
  assign new_n1046_ = ~G171 & ~new_n1035_;
  assign new_n1047_ = ~new_n1045_ & ~new_n1046_;
  assign new_n1048_ = ~new_n1003_ & ~new_n1047_;
  assign new_n1049_ = ~new_n1017_ & new_n1048_;
  assign new_n1050_ = ~new_n994_ & new_n1049_;
  assign new_n1051_ = ~new_n1032_ & new_n1050_;
  assign new_n1052_ = ~G2072 & new_n946_;
  assign new_n1053_ = ~G1956 & ~new_n946_;
  assign new_n1054_ = ~new_n1052_ & ~new_n1053_;
  assign new_n1055_ = ~G299 & ~new_n1054_;
  assign new_n1056_ = ~G299 & new_n1054_;
  assign new_n1057_ = G299 & ~new_n1054_;
  assign new_n1058_ = ~new_n1056_ & ~new_n1057_;
  assign new_n1059_ = ~G2067 & new_n946_;
  assign new_n1060_ = ~G1348 & ~new_n946_;
  assign new_n1061_ = ~new_n1059_ & ~new_n1060_;
  assign new_n1062_ = new_n532_ & ~new_n1061_;
  assign new_n1063_ = ~new_n1058_ & new_n1062_;
  assign new_n1064_ = new_n532_ & new_n1061_;
  assign new_n1065_ = ~new_n532_ & ~new_n1061_;
  assign new_n1066_ = ~new_n1064_ & ~new_n1065_;
  assign new_n1067_ = ~G1996 & new_n946_;
  assign new_n1068_ = ~G1341 & ~new_n946_;
  assign new_n1069_ = ~new_n1067_ & ~new_n1068_;
  assign new_n1070_ = new_n470_ & ~new_n1069_;
  assign new_n1071_ = ~new_n1058_ & ~new_n1066_;
  assign new_n1072_ = new_n1070_ & new_n1071_;
  assign new_n1073_ = ~new_n1055_ & ~new_n1063_;
  assign new_n1074_ = ~new_n1072_ & new_n1073_;
  assign new_n1075_ = new_n1051_ & ~new_n1074_;
  assign new_n1076_ = new_n1044_ & ~new_n1075_;
  assign new_n1077_ = ~new_n986_ & new_n1076_;
  assign new_n1078_ = ~new_n977_ & ~new_n979_;
  assign new_n1079_ = new_n977_ & new_n979_;
  assign new_n1080_ = ~new_n1078_ & ~new_n1079_;
  assign new_n1081_ = ~new_n965_ & ~new_n1080_;
  assign new_n1082_ = ~new_n975_ & new_n1081_;
  assign new_n1083_ = ~new_n956_ & new_n1082_;
  assign new_n1084_ = new_n986_ & ~new_n1083_;
  assign new_n1085_ = ~new_n1076_ & ~new_n1084_;
  assign G329 = new_n1077_ | new_n1085_;
  assign new_n1087_ = ~G395 & ~G397;
  assign new_n1088_ = ~G227 & new_n1087_;
  assign new_n1089_ = ~G401 & ~G229;
  assign new_n1090_ = new_n1088_ & new_n1089_;
  assign G308 = G319 & new_n1090_;
  assign G231 = 1'b0;
  assign G218 = ~G44;
  assign G219 = ~G132;
  assign G220 = ~G82;
  assign G221 = ~G96;
  assign G235 = ~G69;
  assign G236 = ~G120;
  assign G237 = ~G57;
  assign G238 = ~G108;
  assign G261 = ~G325;
  assign G301 = ~G171;
  assign G286 = ~G168;
  assign G303 = ~G166;
  assign G150 = ~G311;
  assign G225 = ~G308;
  assign G169 = \IN-G169 ;
  assign G174 = \IN-G174 ;
  assign G177 = \IN-G177 ;
  assign G178 = \IN-G178 ;
  assign G179 = \IN-G179 ;
  assign G180 = \IN-G180 ;
  assign G181 = \IN-G181 ;
  assign G182 = \IN-G182 ;
  assign G183 = \IN-G183 ;
  assign G184 = \IN-G184 ;
  assign G185 = \IN-G185 ;
  assign G186 = \IN-G186 ;
  assign G189 = \IN-G189 ;
  assign G190 = \IN-G190 ;
  assign G191 = \IN-G191 ;
  assign G192 = \IN-G192 ;
  assign G193 = \IN-G193 ;
  assign G194 = \IN-G194 ;
  assign G195 = \IN-G195 ;
  assign G196 = \IN-G196 ;
  assign G197 = \IN-G197 ;
  assign G198 = \IN-G198 ;
  assign G199 = \IN-G199 ;
  assign G200 = \IN-G200 ;
  assign G201 = \IN-G201 ;
  assign G202 = \IN-G202 ;
  assign G203 = \IN-G203 ;
  assign G204 = \IN-G204 ;
  assign G205 = \IN-G205 ;
  assign G206 = \IN-G206 ;
  assign G207 = \IN-G207 ;
  assign G208 = \IN-G208 ;
  assign G209 = \IN-G209 ;
  assign G210 = \IN-G210 ;
  assign G211 = \IN-G211 ;
  assign G212 = \IN-G212 ;
  assign G213 = \IN-G213 ;
  assign G214 = \IN-G214 ;
  assign G215 = \IN-G215 ;
  assign G239 = \IN-G239 ;
  assign G240 = \IN-G240 ;
  assign G241 = \IN-G241 ;
  assign G242 = \IN-G242 ;
  assign G243 = \IN-G243 ;
  assign G244 = \IN-G244 ;
  assign G245 = \IN-G245 ;
  assign G246 = \IN-G246 ;
  assign G247 = \IN-G247 ;
  assign G248 = \IN-G248 ;
  assign G249 = \IN-G249 ;
  assign G250 = \IN-G250 ;
  assign G251 = \IN-G251 ;
  assign G252 = \IN-G252 ;
  assign G253 = \IN-G253 ;
  assign G254 = \IN-G254 ;
  assign G255 = \IN-G255 ;
  assign G256 = \IN-G256 ;
  assign G257 = \IN-G257 ;
  assign G262 = \IN-G262 ;
  assign G263 = \IN-G263 ;
  assign G264 = \IN-G264 ;
  assign G265 = \IN-G265 ;
  assign G266 = \IN-G266 ;
  assign G267 = \IN-G267 ;
  assign G268 = \IN-G268 ;
  assign G269 = \IN-G269 ;
  assign G270 = \IN-G270 ;
  assign G271 = \IN-G271 ;
  assign G272 = \IN-G272 ;
  assign G273 = \IN-G273 ;
  assign G274 = \IN-G274 ;
  assign G275 = \IN-G275 ;
  assign G276 = \IN-G276 ;
  assign G277 = \IN-G277 ;
  assign G278 = \IN-G278 ;
  assign G279 = \IN-G279 ;
  assign G350 = G452;
  assign G335 = G452;
  assign G409 = G452;
  assign G369 = G1083;
  assign G367 = G1083;
  assign G411 = G2066;
  assign G337 = G2066;
  assign G384 = G2066;
  assign G391 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;
endmodule


