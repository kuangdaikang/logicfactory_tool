// Benchmark "sin" written by ABC on Fri Sep 15 11:23:57 2023

module sin ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ;
  output \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24] ;
  wire new_n50_, new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_,
    new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_,
    new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_,
    new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_,
    new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_,
    new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_,
    new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_,
    new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_,
    new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_,
    new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_,
    new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_,
    new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_,
    new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_,
    new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_,
    new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_,
    new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_,
    new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_,
    new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_,
    new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_,
    new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_,
    new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_,
    new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_,
    new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_,
    new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_,
    new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_,
    new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_,
    new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_,
    new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_,
    new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_,
    new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_,
    new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_,
    new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_,
    new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_,
    new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_,
    new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_,
    new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_,
    new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_,
    new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_,
    new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_,
    new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_,
    new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_,
    new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_,
    new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_,
    new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_,
    new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_,
    new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_,
    new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_,
    new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_,
    new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_,
    new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_,
    new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_,
    new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_,
    new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_,
    new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_,
    new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_,
    new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_,
    new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_,
    new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_,
    new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_,
    new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_,
    new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_,
    new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_,
    new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_,
    new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_,
    new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_,
    new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_,
    new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_,
    new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_,
    new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_,
    new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_,
    new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_,
    new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_,
    new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_,
    new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_,
    new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_,
    new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_,
    new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_,
    new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_,
    new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_,
    new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_,
    new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_,
    new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_,
    new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_,
    new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_,
    new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_,
    new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_,
    new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_,
    new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_,
    new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_,
    new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_,
    new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_,
    new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_,
    new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_,
    new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_,
    new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_,
    new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_,
    new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_,
    new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_,
    new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_,
    new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_,
    new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_,
    new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_,
    new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_,
    new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_,
    new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_,
    new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_,
    new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_,
    new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_,
    new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_,
    new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_,
    new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_,
    new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_,
    new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_,
    new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_,
    new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_,
    new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_,
    new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_,
    new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_,
    new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_,
    new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_,
    new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_,
    new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_,
    new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_,
    new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_,
    new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_,
    new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_,
    new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_,
    new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_,
    new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_,
    new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_,
    new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_,
    new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_,
    new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_,
    new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_,
    new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_,
    new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_,
    new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_,
    new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_,
    new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_,
    new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_,
    new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_,
    new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_,
    new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_,
    new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_,
    new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_,
    new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_,
    new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_,
    new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_,
    new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_,
    new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_,
    new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_,
    new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_,
    new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_,
    new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_,
    new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_,
    new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_,
    new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_,
    new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_,
    new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_,
    new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_,
    new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_,
    new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_,
    new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_,
    new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_,
    new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_,
    new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_,
    new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_,
    new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_,
    new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_,
    new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_,
    new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_,
    new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_,
    new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_,
    new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_,
    new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_,
    new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_,
    new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_,
    new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_,
    new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_,
    new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_,
    new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_,
    new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_,
    new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_,
    new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_,
    new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_,
    new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_,
    new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_,
    new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_,
    new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_,
    new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_,
    new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_,
    new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_,
    new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_,
    new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_,
    new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_,
    new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_,
    new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_,
    new_n4071_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_,
    new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_,
    new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_,
    new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_,
    new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_,
    new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_,
    new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_,
    new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_,
    new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_,
    new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_,
    new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_,
    new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_,
    new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_,
    new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_,
    new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_,
    new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_,
    new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_,
    new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_,
    new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_,
    new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_,
    new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_,
    new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_,
    new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_,
    new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_,
    new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_,
    new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_,
    new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_,
    new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_,
    new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4385_, new_n4386_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4515_, new_n4516_, new_n4517_, new_n4518_,
    new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_,
    new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_,
    new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_,
    new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_,
    new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_,
    new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_,
    new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_,
    new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_,
    new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_,
    new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_,
    new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_,
    new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_,
    new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_,
    new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_,
    new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_,
    new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_,
    new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_,
    new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_,
    new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_,
    new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_,
    new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_,
    new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_,
    new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_,
    new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_,
    new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_,
    new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_,
    new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_,
    new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_,
    new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_,
    new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_,
    new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_,
    new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_,
    new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_,
    new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_,
    new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_,
    new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_,
    new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_,
    new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_,
    new_n4833_, new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_,
    new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_,
    new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_,
    new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_,
    new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_,
    new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_,
    new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_,
    new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_,
    new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_,
    new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_,
    new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_,
    new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_,
    new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_,
    new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_,
    new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4924_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_,
    new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_,
    new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_,
    new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_,
    new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_,
    new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_,
    new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_,
    new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_,
    new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_,
    new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_,
    new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_,
    new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_,
    new_n5009_, new_n5010_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5069_, new_n5070_,
    new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_,
    new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_,
    new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_,
    new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_,
    new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_,
    new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_,
    new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_,
    new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_,
    new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5168_,
    new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_,
    new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_,
    new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_,
    new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_,
    new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_,
    new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_,
    new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_,
    new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_,
    new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_,
    new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_,
    new_n5229_, new_n5230_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_,
    new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_,
    new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_,
    new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_,
    new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_,
    new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_,
    new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_,
    new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_,
    new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_,
    new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_,
    new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_,
    new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_,
    new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_,
    new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_,
    new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_,
    new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_,
    new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_,
    new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_,
    new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_,
    new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_,
    new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_,
    new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_,
    new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_,
    new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_,
    new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_,
    new_n5455_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5480_,
    new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_,
    new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_,
    new_n5493_, new_n5494_, new_n5495_, new_n5497_, new_n5498_, new_n5499_,
    new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_,
    new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5512_,
    new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_,
    new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_,
    new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_,
    new_n5531_, new_n5532_, new_n5534_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5553_, new_n5554_, new_n5555_, new_n5556_,
    new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_,
    new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5582_,
    new_n5583_, new_n5584_, new_n5585_;
  NOR2_X1    g0000(.A1(\a[0] ), .A2(\a[1] ), .ZN(new_n50_));
  NOR2_X1    g0001(.A1(new_n50_), .A2(\a[22] ), .ZN(new_n51_));
  XOR2_X1    g0002(.A1(new_n51_), .A2(\a[2] ), .Z(new_n52_));
  INV_X1     g0003(.I(\a[2] ), .ZN(new_n53_));
  INV_X1     g0004(.I(new_n50_), .ZN(new_n54_));
  NOR2_X1    g0005(.A1(new_n54_), .A2(new_n53_), .ZN(new_n55_));
  INV_X1     g0006(.I(new_n55_), .ZN(new_n56_));
  INV_X1     g0007(.I(\a[22] ), .ZN(new_n57_));
  OR3_X2     g0008(.A1(\a[4] ), .A2(\a[5] ), .A3(\a[6] ), .Z(new_n58_));
  OR4_X2     g0009(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[2] ), .A4(\a[3] ), .Z(new_n59_));
  NOR2_X1    g0010(.A1(new_n59_), .A2(new_n58_), .ZN(new_n60_));
  NOR3_X1    g0011(.A1(\a[7] ), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n61_));
  NOR3_X1    g0012(.A1(\a[10] ), .A2(\a[11] ), .A3(\a[12] ), .ZN(new_n62_));
  NOR2_X1    g0013(.A1(\a[13] ), .A2(\a[14] ), .ZN(new_n63_));
  NAND4_X1   g0014(.A1(new_n60_), .A2(new_n61_), .A3(new_n62_), .A4(new_n63_), .ZN(new_n64_));
  AOI21_X1   g0015(.A1(new_n64_), .A2(new_n57_), .B(\a[15] ), .ZN(new_n65_));
  INV_X1     g0016(.I(\a[15] ), .ZN(new_n66_));
  NOR3_X1    g0017(.A1(\a[4] ), .A2(\a[5] ), .A3(\a[6] ), .ZN(new_n67_));
  NOR4_X1    g0018(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[2] ), .A4(\a[3] ), .ZN(new_n68_));
  NAND4_X1   g0019(.A1(new_n68_), .A2(new_n67_), .A3(new_n61_), .A4(new_n62_), .ZN(new_n69_));
  INV_X1     g0020(.I(new_n63_), .ZN(new_n70_));
  NOR2_X1    g0021(.A1(new_n69_), .A2(new_n70_), .ZN(new_n71_));
  NOR3_X1    g0022(.A1(new_n71_), .A2(new_n66_), .A3(\a[22] ), .ZN(new_n72_));
  NOR2_X1    g0023(.A1(new_n65_), .A2(new_n72_), .ZN(new_n73_));
  INV_X1     g0024(.I(\a[20] ), .ZN(new_n74_));
  INV_X1     g0025(.I(\a[21] ), .ZN(new_n75_));
  NOR3_X1    g0026(.A1(new_n74_), .A2(new_n75_), .A3(new_n57_), .ZN(new_n76_));
  NOR3_X1    g0027(.A1(\a[15] ), .A2(\a[16] ), .A3(\a[17] ), .ZN(new_n77_));
  INV_X1     g0028(.I(new_n77_), .ZN(new_n78_));
  NOR2_X1    g0029(.A1(\a[18] ), .A2(\a[19] ), .ZN(new_n79_));
  INV_X1     g0030(.I(new_n79_), .ZN(new_n80_));
  NOR4_X1    g0031(.A1(new_n69_), .A2(new_n70_), .A3(new_n78_), .A4(new_n80_), .ZN(new_n81_));
  NAND2_X1   g0032(.A1(new_n81_), .A2(\a[20] ), .ZN(new_n82_));
  OR3_X2     g0033(.A1(\a[7] ), .A2(\a[8] ), .A3(\a[9] ), .Z(new_n83_));
  OR3_X2     g0034(.A1(\a[10] ), .A2(\a[11] ), .A3(\a[12] ), .Z(new_n84_));
  NOR4_X1    g0035(.A1(new_n59_), .A2(new_n58_), .A3(new_n83_), .A4(new_n84_), .ZN(new_n85_));
  NAND4_X1   g0036(.A1(new_n85_), .A2(new_n63_), .A3(new_n77_), .A4(new_n79_), .ZN(new_n86_));
  NAND2_X1   g0037(.A1(new_n86_), .A2(new_n74_), .ZN(new_n87_));
  NOR2_X1    g0038(.A1(\a[21] ), .A2(\a[22] ), .ZN(new_n88_));
  INV_X1     g0039(.I(new_n88_), .ZN(new_n89_));
  AOI21_X1   g0040(.A1(new_n87_), .A2(new_n82_), .B(new_n89_), .ZN(new_n90_));
  OAI21_X1   g0041(.A1(new_n90_), .A2(new_n76_), .B(new_n73_), .ZN(new_n91_));
  INV_X1     g0042(.I(\a[19] ), .ZN(new_n92_));
  NAND3_X1   g0043(.A1(new_n85_), .A2(new_n63_), .A3(new_n77_), .ZN(new_n93_));
  NAND2_X1   g0044(.A1(new_n93_), .A2(new_n57_), .ZN(new_n94_));
  INV_X1     g0045(.I(\a[18] ), .ZN(new_n95_));
  NOR3_X1    g0046(.A1(new_n69_), .A2(new_n70_), .A3(new_n78_), .ZN(new_n96_));
  OAI21_X1   g0047(.A1(new_n96_), .A2(\a[22] ), .B(new_n95_), .ZN(new_n97_));
  NAND2_X1   g0048(.A1(new_n92_), .A2(\a[18] ), .ZN(new_n98_));
  OAI22_X1   g0049(.A1(new_n94_), .A2(new_n98_), .B1(new_n97_), .B2(new_n92_), .ZN(new_n99_));
  INV_X1     g0050(.I(\a[16] ), .ZN(new_n100_));
  NOR4_X1    g0051(.A1(new_n69_), .A2(\a[15] ), .A3(new_n100_), .A4(new_n70_), .ZN(new_n101_));
  NOR3_X1    g0052(.A1(new_n69_), .A2(\a[15] ), .A3(new_n70_), .ZN(new_n102_));
  NOR2_X1    g0053(.A1(new_n102_), .A2(\a[16] ), .ZN(new_n103_));
  OAI21_X1   g0054(.A1(new_n103_), .A2(new_n101_), .B(new_n57_), .ZN(new_n104_));
  INV_X1     g0055(.I(\a[17] ), .ZN(new_n105_));
  NOR2_X1    g0056(.A1(new_n100_), .A2(new_n105_), .ZN(new_n106_));
  INV_X1     g0057(.I(new_n106_), .ZN(new_n107_));
  OAI22_X1   g0058(.A1(new_n104_), .A2(\a[17] ), .B1(new_n57_), .B2(new_n107_), .ZN(new_n108_));
  NAND2_X1   g0059(.A1(new_n108_), .A2(new_n99_), .ZN(new_n109_));
  NOR2_X1    g0060(.A1(new_n109_), .A2(new_n91_), .ZN(new_n110_));
  NOR3_X1    g0061(.A1(new_n59_), .A2(new_n58_), .A3(new_n83_), .ZN(new_n111_));
  NAND4_X1   g0062(.A1(new_n111_), .A2(new_n66_), .A3(new_n62_), .A4(new_n63_), .ZN(new_n112_));
  NAND2_X1   g0063(.A1(new_n112_), .A2(new_n57_), .ZN(new_n113_));
  OAI21_X1   g0064(.A1(new_n102_), .A2(\a[22] ), .B(new_n100_), .ZN(new_n114_));
  OAI22_X1   g0065(.A1(new_n113_), .A2(new_n107_), .B1(new_n114_), .B2(\a[17] ), .ZN(new_n115_));
  NOR2_X1    g0066(.A1(new_n98_), .A2(new_n57_), .ZN(new_n116_));
  INV_X1     g0067(.I(new_n116_), .ZN(new_n117_));
  NOR4_X1    g0068(.A1(new_n69_), .A2(new_n95_), .A3(new_n70_), .A4(new_n78_), .ZN(new_n118_));
  NOR2_X1    g0069(.A1(new_n96_), .A2(\a[18] ), .ZN(new_n119_));
  OAI21_X1   g0070(.A1(new_n119_), .A2(new_n118_), .B(new_n57_), .ZN(new_n120_));
  OAI21_X1   g0071(.A1(new_n120_), .A2(new_n92_), .B(new_n117_), .ZN(new_n121_));
  NAND2_X1   g0072(.A1(new_n121_), .A2(new_n115_), .ZN(new_n122_));
  OAI21_X1   g0073(.A1(new_n71_), .A2(\a[22] ), .B(new_n66_), .ZN(new_n123_));
  NAND3_X1   g0074(.A1(new_n64_), .A2(\a[15] ), .A3(new_n57_), .ZN(new_n124_));
  NAND2_X1   g0075(.A1(new_n124_), .A2(new_n123_), .ZN(new_n125_));
  OAI21_X1   g0076(.A1(new_n90_), .A2(new_n76_), .B(new_n125_), .ZN(new_n126_));
  NOR2_X1    g0077(.A1(new_n122_), .A2(new_n126_), .ZN(new_n127_));
  NAND2_X1   g0078(.A1(new_n81_), .A2(new_n74_), .ZN(new_n128_));
  AOI21_X1   g0079(.A1(new_n128_), .A2(new_n57_), .B(\a[21] ), .ZN(new_n129_));
  NOR4_X1    g0080(.A1(new_n64_), .A2(\a[20] ), .A3(new_n78_), .A4(new_n80_), .ZN(new_n130_));
  NOR3_X1    g0081(.A1(new_n130_), .A2(new_n75_), .A3(\a[22] ), .ZN(new_n131_));
  OAI21_X1   g0082(.A1(new_n81_), .A2(\a[22] ), .B(new_n74_), .ZN(new_n132_));
  NAND3_X1   g0083(.A1(new_n86_), .A2(\a[20] ), .A3(new_n57_), .ZN(new_n133_));
  NAND2_X1   g0084(.A1(new_n133_), .A2(new_n132_), .ZN(new_n134_));
  OAI21_X1   g0085(.A1(new_n129_), .A2(new_n131_), .B(new_n134_), .ZN(new_n135_));
  NAND2_X1   g0086(.A1(new_n105_), .A2(\a[16] ), .ZN(new_n136_));
  OAI22_X1   g0087(.A1(new_n113_), .A2(new_n136_), .B1(new_n114_), .B2(new_n105_), .ZN(new_n137_));
  NAND2_X1   g0088(.A1(new_n99_), .A2(new_n137_), .ZN(new_n138_));
  NOR3_X1    g0089(.A1(new_n135_), .A2(new_n138_), .A3(new_n73_), .ZN(new_n139_));
  NOR3_X1    g0090(.A1(new_n110_), .A2(new_n139_), .A3(new_n127_), .ZN(new_n140_));
  INV_X1     g0091(.I(new_n140_), .ZN(new_n141_));
  NAND2_X1   g0092(.A1(\a[18] ), .A2(\a[19] ), .ZN(new_n142_));
  NOR2_X1    g0093(.A1(new_n142_), .A2(new_n57_), .ZN(new_n143_));
  INV_X1     g0094(.I(new_n143_), .ZN(new_n144_));
  OAI21_X1   g0095(.A1(new_n120_), .A2(\a[19] ), .B(new_n144_), .ZN(new_n145_));
  AOI21_X1   g0096(.A1(new_n86_), .A2(new_n57_), .B(\a[20] ), .ZN(new_n146_));
  NOR3_X1    g0097(.A1(new_n81_), .A2(new_n74_), .A3(\a[22] ), .ZN(new_n147_));
  NAND2_X1   g0098(.A1(\a[21] ), .A2(\a[22] ), .ZN(new_n148_));
  NAND2_X1   g0099(.A1(new_n89_), .A2(new_n148_), .ZN(new_n149_));
  NOR3_X1    g0100(.A1(new_n146_), .A2(new_n147_), .A3(new_n149_), .ZN(new_n150_));
  NAND4_X1   g0101(.A1(new_n108_), .A2(new_n145_), .A3(new_n73_), .A4(new_n150_), .ZN(new_n151_));
  NOR2_X1    g0102(.A1(new_n136_), .A2(new_n57_), .ZN(new_n152_));
  INV_X1     g0103(.I(new_n152_), .ZN(new_n153_));
  OAI21_X1   g0104(.A1(new_n104_), .A2(new_n105_), .B(new_n153_), .ZN(new_n154_));
  NAND2_X1   g0105(.A1(new_n154_), .A2(new_n99_), .ZN(new_n155_));
  NOR2_X1    g0106(.A1(new_n155_), .A2(new_n91_), .ZN(new_n156_));
  INV_X1     g0107(.I(new_n156_), .ZN(new_n157_));
  NAND2_X1   g0108(.A1(new_n145_), .A2(new_n115_), .ZN(new_n158_));
  NOR2_X1    g0109(.A1(new_n158_), .A2(new_n126_), .ZN(new_n159_));
  INV_X1     g0110(.I(new_n159_), .ZN(new_n160_));
  NAND3_X1   g0111(.A1(new_n160_), .A2(new_n157_), .A3(new_n151_), .ZN(new_n161_));
  OAI22_X1   g0112(.A1(new_n94_), .A2(new_n142_), .B1(new_n97_), .B2(\a[19] ), .ZN(new_n162_));
  NAND2_X1   g0113(.A1(new_n108_), .A2(new_n162_), .ZN(new_n163_));
  NOR2_X1    g0114(.A1(new_n163_), .A2(new_n126_), .ZN(new_n164_));
  OAI21_X1   g0115(.A1(new_n130_), .A2(\a[22] ), .B(new_n75_), .ZN(new_n165_));
  NAND3_X1   g0116(.A1(new_n128_), .A2(\a[21] ), .A3(new_n57_), .ZN(new_n166_));
  NAND4_X1   g0117(.A1(new_n134_), .A2(new_n165_), .A3(new_n125_), .A4(new_n166_), .ZN(new_n167_));
  NOR2_X1    g0118(.A1(new_n109_), .A2(new_n167_), .ZN(new_n168_));
  NOR4_X1    g0119(.A1(new_n141_), .A2(new_n161_), .A3(new_n164_), .A4(new_n168_), .ZN(new_n169_));
  INV_X1     g0120(.I(new_n169_), .ZN(new_n170_));
  INV_X1     g0121(.I(new_n149_), .ZN(new_n171_));
  NAND3_X1   g0122(.A1(new_n133_), .A2(new_n132_), .A3(new_n171_), .ZN(new_n172_));
  NAND3_X1   g0123(.A1(new_n121_), .A2(new_n73_), .A3(new_n137_), .ZN(new_n173_));
  NAND3_X1   g0124(.A1(new_n145_), .A2(new_n125_), .A3(new_n115_), .ZN(new_n174_));
  AOI21_X1   g0125(.A1(new_n173_), .A2(new_n174_), .B(new_n172_), .ZN(new_n175_));
  INV_X1     g0126(.I(new_n175_), .ZN(new_n176_));
  NOR2_X1    g0127(.A1(new_n155_), .A2(new_n126_), .ZN(new_n177_));
  NAND2_X1   g0128(.A1(new_n108_), .A2(new_n121_), .ZN(new_n178_));
  NOR2_X1    g0129(.A1(new_n178_), .A2(new_n167_), .ZN(new_n179_));
  NOR2_X1    g0130(.A1(new_n179_), .A2(new_n177_), .ZN(new_n180_));
  NAND2_X1   g0131(.A1(new_n165_), .A2(new_n166_), .ZN(new_n181_));
  NOR2_X1    g0132(.A1(new_n146_), .A2(new_n147_), .ZN(new_n182_));
  NOR2_X1    g0133(.A1(new_n182_), .A2(new_n125_), .ZN(new_n183_));
  NAND2_X1   g0134(.A1(new_n183_), .A2(new_n181_), .ZN(new_n184_));
  NOR2_X1    g0135(.A1(new_n184_), .A2(new_n122_), .ZN(new_n185_));
  NAND2_X1   g0136(.A1(new_n121_), .A2(new_n154_), .ZN(new_n186_));
  NOR2_X1    g0137(.A1(new_n184_), .A2(new_n186_), .ZN(new_n187_));
  NOR2_X1    g0138(.A1(new_n122_), .A2(new_n167_), .ZN(new_n188_));
  NOR3_X1    g0139(.A1(new_n185_), .A2(new_n187_), .A3(new_n188_), .ZN(new_n189_));
  NAND4_X1   g0140(.A1(new_n154_), .A2(new_n73_), .A3(new_n150_), .A4(new_n99_), .ZN(new_n190_));
  INV_X1     g0141(.I(new_n190_), .ZN(new_n191_));
  NAND3_X1   g0142(.A1(new_n181_), .A2(new_n125_), .A3(new_n134_), .ZN(new_n192_));
  NOR2_X1    g0143(.A1(new_n192_), .A2(new_n186_), .ZN(new_n193_));
  NAND2_X1   g0144(.A1(new_n99_), .A2(new_n115_), .ZN(new_n194_));
  NAND4_X1   g0145(.A1(new_n125_), .A2(new_n132_), .A3(new_n133_), .A4(new_n171_), .ZN(new_n195_));
  NOR2_X1    g0146(.A1(new_n194_), .A2(new_n195_), .ZN(new_n196_));
  NOR2_X1    g0147(.A1(new_n184_), .A2(new_n138_), .ZN(new_n197_));
  NOR4_X1    g0148(.A1(new_n197_), .A2(new_n193_), .A3(new_n191_), .A4(new_n196_), .ZN(new_n198_));
  NAND4_X1   g0149(.A1(new_n198_), .A2(new_n189_), .A3(new_n176_), .A4(new_n180_), .ZN(new_n199_));
  NOR2_X1    g0150(.A1(new_n163_), .A2(new_n167_), .ZN(new_n200_));
  NOR2_X1    g0151(.A1(new_n158_), .A2(new_n167_), .ZN(new_n201_));
  NOR2_X1    g0152(.A1(new_n186_), .A2(new_n167_), .ZN(new_n202_));
  NAND4_X1   g0153(.A1(new_n73_), .A2(new_n132_), .A3(new_n133_), .A4(new_n171_), .ZN(new_n203_));
  NAND2_X1   g0154(.A1(new_n145_), .A2(new_n154_), .ZN(new_n204_));
  NOR2_X1    g0155(.A1(new_n204_), .A2(new_n203_), .ZN(new_n205_));
  NOR4_X1    g0156(.A1(new_n200_), .A2(new_n202_), .A3(new_n205_), .A4(new_n201_), .ZN(new_n206_));
  NOR2_X1    g0157(.A1(new_n126_), .A2(new_n194_), .ZN(new_n207_));
  NOR2_X1    g0158(.A1(new_n204_), .A2(new_n167_), .ZN(new_n208_));
  NAND2_X1   g0159(.A1(new_n108_), .A2(new_n145_), .ZN(new_n209_));
  NOR2_X1    g0160(.A1(new_n192_), .A2(new_n209_), .ZN(new_n210_));
  NOR3_X1    g0161(.A1(new_n210_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n211_));
  INV_X1     g0162(.I(new_n76_), .ZN(new_n212_));
  NOR4_X1    g0163(.A1(new_n64_), .A2(new_n74_), .A3(new_n78_), .A4(new_n80_), .ZN(new_n213_));
  NOR2_X1    g0164(.A1(new_n81_), .A2(\a[20] ), .ZN(new_n214_));
  OAI21_X1   g0165(.A1(new_n213_), .A2(new_n214_), .B(new_n88_), .ZN(new_n215_));
  NAND2_X1   g0166(.A1(new_n215_), .A2(new_n212_), .ZN(new_n216_));
  AOI21_X1   g0167(.A1(new_n112_), .A2(new_n57_), .B(\a[16] ), .ZN(new_n217_));
  NOR3_X1    g0168(.A1(new_n102_), .A2(\a[22] ), .A3(new_n107_), .ZN(new_n218_));
  AOI21_X1   g0169(.A1(new_n217_), .A2(new_n105_), .B(new_n218_), .ZN(new_n219_));
  AOI21_X1   g0170(.A1(new_n93_), .A2(new_n57_), .B(\a[18] ), .ZN(new_n220_));
  NOR3_X1    g0171(.A1(new_n96_), .A2(\a[22] ), .A3(new_n142_), .ZN(new_n221_));
  AOI21_X1   g0172(.A1(new_n220_), .A2(new_n92_), .B(new_n221_), .ZN(new_n222_));
  NOR2_X1    g0173(.A1(new_n222_), .A2(new_n219_), .ZN(new_n223_));
  NAND3_X1   g0174(.A1(new_n223_), .A2(new_n216_), .A3(new_n73_), .ZN(new_n224_));
  NAND3_X1   g0175(.A1(new_n108_), .A2(new_n73_), .A3(new_n162_), .ZN(new_n225_));
  OAI21_X1   g0176(.A1(new_n172_), .A2(new_n225_), .B(new_n224_), .ZN(new_n226_));
  NOR4_X1    g0177(.A1(new_n182_), .A2(new_n131_), .A3(new_n73_), .A4(new_n129_), .ZN(new_n227_));
  NAND2_X1   g0178(.A1(new_n227_), .A2(new_n223_), .ZN(new_n228_));
  AOI22_X1   g0179(.A1(new_n165_), .A2(new_n166_), .B1(new_n132_), .B2(new_n133_), .ZN(new_n229_));
  NAND4_X1   g0180(.A1(new_n229_), .A2(new_n125_), .A3(new_n145_), .A4(new_n154_), .ZN(new_n230_));
  NAND2_X1   g0181(.A1(new_n230_), .A2(new_n228_), .ZN(new_n231_));
  NAND2_X1   g0182(.A1(new_n145_), .A2(new_n137_), .ZN(new_n232_));
  NAND2_X1   g0183(.A1(new_n154_), .A2(new_n162_), .ZN(new_n233_));
  AOI21_X1   g0184(.A1(new_n232_), .A2(new_n233_), .B(new_n91_), .ZN(new_n234_));
  NOR4_X1    g0185(.A1(new_n182_), .A2(new_n131_), .A3(new_n125_), .A4(new_n129_), .ZN(new_n235_));
  NAND3_X1   g0186(.A1(new_n235_), .A2(new_n137_), .A3(new_n145_), .ZN(new_n236_));
  NOR3_X1    g0187(.A1(new_n96_), .A2(\a[22] ), .A3(new_n98_), .ZN(new_n237_));
  AOI21_X1   g0188(.A1(new_n220_), .A2(\a[19] ), .B(new_n237_), .ZN(new_n238_));
  NOR2_X1    g0189(.A1(new_n238_), .A2(new_n219_), .ZN(new_n239_));
  NAND2_X1   g0190(.A1(new_n227_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1   g0191(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  NOR4_X1    g0192(.A1(new_n226_), .A2(new_n231_), .A3(new_n241_), .A4(new_n234_), .ZN(new_n242_));
  NOR2_X1    g0193(.A1(new_n90_), .A2(new_n76_), .ZN(new_n243_));
  NOR2_X1    g0194(.A1(new_n173_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1    g0195(.A1(new_n167_), .A2(new_n138_), .ZN(new_n245_));
  NOR2_X1    g0196(.A1(new_n163_), .A2(new_n195_), .ZN(new_n246_));
  NOR3_X1    g0197(.A1(new_n246_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n247_));
  NAND4_X1   g0198(.A1(new_n242_), .A2(new_n206_), .A3(new_n211_), .A4(new_n247_), .ZN(new_n248_));
  NAND2_X1   g0199(.A1(new_n121_), .A2(new_n137_), .ZN(new_n249_));
  NOR3_X1    g0200(.A1(new_n249_), .A2(new_n135_), .A3(new_n73_), .ZN(new_n250_));
  NOR2_X1    g0201(.A1(new_n131_), .A2(new_n129_), .ZN(new_n251_));
  NAND2_X1   g0202(.A1(new_n134_), .A2(new_n73_), .ZN(new_n252_));
  NOR3_X1    g0203(.A1(new_n155_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  NOR2_X1    g0204(.A1(new_n155_), .A2(new_n167_), .ZN(new_n254_));
  NAND4_X1   g0205(.A1(new_n229_), .A2(new_n125_), .A3(new_n108_), .A4(new_n121_), .ZN(new_n255_));
  INV_X1     g0206(.I(new_n255_), .ZN(new_n256_));
  NOR4_X1    g0207(.A1(new_n256_), .A2(new_n250_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n257_));
  INV_X1     g0208(.I(new_n257_), .ZN(new_n258_));
  NOR2_X1    g0209(.A1(new_n184_), .A2(new_n249_), .ZN(new_n259_));
  NAND4_X1   g0210(.A1(new_n183_), .A2(new_n181_), .A3(new_n108_), .A4(new_n145_), .ZN(new_n260_));
  INV_X1     g0211(.I(new_n260_), .ZN(new_n261_));
  NOR2_X1    g0212(.A1(new_n186_), .A2(new_n91_), .ZN(new_n262_));
  NOR2_X1    g0213(.A1(new_n204_), .A2(new_n126_), .ZN(new_n263_));
  NOR4_X1    g0214(.A1(new_n261_), .A2(new_n259_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n264_));
  NOR2_X1    g0215(.A1(new_n233_), .A2(new_n167_), .ZN(new_n265_));
  NAND4_X1   g0216(.A1(new_n134_), .A2(new_n165_), .A3(new_n73_), .A4(new_n166_), .ZN(new_n266_));
  NOR2_X1    g0217(.A1(new_n209_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1    g0218(.A1(new_n267_), .A2(new_n265_), .ZN(new_n268_));
  NOR2_X1    g0219(.A1(new_n91_), .A2(new_n138_), .ZN(new_n269_));
  NAND2_X1   g0220(.A1(new_n162_), .A2(new_n137_), .ZN(new_n270_));
  NOR2_X1    g0221(.A1(new_n167_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1    g0222(.A1(new_n126_), .A2(new_n270_), .ZN(new_n272_));
  NOR3_X1    g0223(.A1(new_n269_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND3_X1   g0224(.A1(new_n264_), .A2(new_n273_), .A3(new_n268_), .ZN(new_n274_));
  NAND4_X1   g0225(.A1(new_n183_), .A2(new_n181_), .A3(new_n115_), .A4(new_n145_), .ZN(new_n275_));
  INV_X1     g0226(.I(new_n275_), .ZN(new_n276_));
  NOR3_X1    g0227(.A1(new_n204_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n277_));
  NOR2_X1    g0228(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NOR3_X1    g0229(.A1(new_n102_), .A2(\a[22] ), .A3(new_n136_), .ZN(new_n279_));
  AOI21_X1   g0230(.A1(new_n217_), .A2(\a[17] ), .B(new_n279_), .ZN(new_n280_));
  INV_X1     g0231(.I(new_n118_), .ZN(new_n281_));
  NAND2_X1   g0232(.A1(new_n93_), .A2(new_n95_), .ZN(new_n282_));
  AOI21_X1   g0233(.A1(new_n282_), .A2(new_n281_), .B(\a[22] ), .ZN(new_n283_));
  AOI21_X1   g0234(.A1(new_n283_), .A2(new_n92_), .B(new_n143_), .ZN(new_n284_));
  NOR3_X1    g0235(.A1(new_n284_), .A2(new_n203_), .A3(new_n280_), .ZN(new_n285_));
  AOI21_X1   g0236(.A1(new_n283_), .A2(\a[19] ), .B(new_n116_), .ZN(new_n286_));
  INV_X1     g0237(.I(new_n101_), .ZN(new_n287_));
  NAND2_X1   g0238(.A1(new_n112_), .A2(new_n100_), .ZN(new_n288_));
  AOI21_X1   g0239(.A1(new_n288_), .A2(new_n287_), .B(\a[22] ), .ZN(new_n289_));
  AOI21_X1   g0240(.A1(new_n289_), .A2(\a[17] ), .B(new_n152_), .ZN(new_n290_));
  NOR3_X1    g0241(.A1(new_n286_), .A2(new_n290_), .A3(new_n195_), .ZN(new_n291_));
  NOR2_X1    g0242(.A1(new_n291_), .A2(new_n285_), .ZN(new_n292_));
  NAND4_X1   g0243(.A1(new_n216_), .A2(new_n108_), .A3(new_n145_), .A4(new_n73_), .ZN(new_n293_));
  INV_X1     g0244(.I(new_n293_), .ZN(new_n294_));
  AOI22_X1   g0245(.A1(new_n289_), .A2(new_n105_), .B1(\a[22] ), .B2(new_n106_), .ZN(new_n295_));
  NOR3_X1    g0246(.A1(new_n295_), .A2(new_n238_), .A3(new_n195_), .ZN(new_n296_));
  NOR2_X1    g0247(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1   g0248(.A1(new_n278_), .A2(new_n297_), .A3(new_n292_), .ZN(new_n298_));
  NOR3_X1    g0249(.A1(new_n290_), .A2(new_n195_), .A3(new_n222_), .ZN(new_n299_));
  INV_X1     g0250(.I(new_n299_), .ZN(new_n300_));
  NAND4_X1   g0251(.A1(new_n154_), .A2(new_n73_), .A3(new_n150_), .A4(new_n162_), .ZN(new_n301_));
  NOR3_X1    g0252(.A1(new_n182_), .A2(new_n131_), .A3(new_n129_), .ZN(new_n302_));
  NAND4_X1   g0253(.A1(new_n302_), .A2(new_n125_), .A3(new_n121_), .A4(new_n137_), .ZN(new_n303_));
  NAND3_X1   g0254(.A1(new_n300_), .A2(new_n303_), .A3(new_n301_), .ZN(new_n304_));
  NOR4_X1    g0255(.A1(new_n274_), .A2(new_n258_), .A3(new_n298_), .A4(new_n304_), .ZN(new_n305_));
  INV_X1     g0256(.I(new_n305_), .ZN(new_n306_));
  NOR4_X1    g0257(.A1(new_n306_), .A2(new_n170_), .A3(new_n199_), .A4(new_n248_), .ZN(new_n307_));
  INV_X1     g0258(.I(new_n307_), .ZN(new_n308_));
  AOI21_X1   g0259(.A1(new_n209_), .A2(new_n270_), .B(new_n243_), .ZN(new_n309_));
  NOR2_X1    g0260(.A1(new_n178_), .A2(new_n266_), .ZN(new_n310_));
  NOR2_X1    g0261(.A1(new_n310_), .A2(new_n262_), .ZN(new_n311_));
  NOR2_X1    g0262(.A1(new_n186_), .A2(new_n126_), .ZN(new_n312_));
  NOR2_X1    g0263(.A1(new_n109_), .A2(new_n266_), .ZN(new_n313_));
  NOR2_X1    g0264(.A1(new_n313_), .A2(new_n312_), .ZN(new_n314_));
  AOI21_X1   g0265(.A1(new_n215_), .A2(new_n212_), .B(new_n125_), .ZN(new_n315_));
  NAND2_X1   g0266(.A1(new_n239_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1   g0267(.A1(new_n155_), .A2(new_n249_), .B(new_n126_), .ZN(new_n317_));
  NOR2_X1    g0268(.A1(new_n168_), .A2(new_n207_), .ZN(new_n318_));
  INV_X1     g0269(.I(new_n318_), .ZN(new_n319_));
  NAND3_X1   g0270(.A1(new_n134_), .A2(new_n165_), .A3(new_n166_), .ZN(new_n320_));
  NOR2_X1    g0271(.A1(new_n173_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1    g0272(.A1(new_n179_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1     g0273(.I(new_n322_), .ZN(new_n323_));
  NOR2_X1    g0274(.A1(new_n320_), .A2(new_n138_), .ZN(new_n324_));
  NOR4_X1    g0275(.A1(new_n323_), .A2(new_n319_), .A3(new_n317_), .A4(new_n324_), .ZN(new_n325_));
  NAND4_X1   g0276(.A1(new_n325_), .A2(new_n311_), .A3(new_n314_), .A4(new_n316_), .ZN(new_n326_));
  NOR2_X1    g0277(.A1(new_n232_), .A2(new_n167_), .ZN(new_n327_));
  NOR2_X1    g0278(.A1(new_n110_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1   g0279(.A1(new_n227_), .A2(new_n108_), .A3(new_n145_), .ZN(new_n329_));
  NOR2_X1    g0280(.A1(new_n232_), .A2(new_n266_), .ZN(new_n330_));
  NAND3_X1   g0281(.A1(new_n145_), .A2(new_n73_), .A3(new_n115_), .ZN(new_n331_));
  NOR2_X1    g0282(.A1(new_n331_), .A2(new_n243_), .ZN(new_n332_));
  NOR2_X1    g0283(.A1(new_n332_), .A2(new_n330_), .ZN(new_n333_));
  NAND4_X1   g0284(.A1(new_n328_), .A2(new_n333_), .A3(new_n160_), .A4(new_n329_), .ZN(new_n334_));
  NOR4_X1    g0285(.A1(new_n326_), .A2(new_n234_), .A3(new_n309_), .A4(new_n334_), .ZN(new_n335_));
  NAND3_X1   g0286(.A1(new_n162_), .A2(new_n115_), .A3(new_n73_), .ZN(new_n336_));
  NOR2_X1    g0287(.A1(new_n336_), .A2(new_n243_), .ZN(new_n337_));
  NOR2_X1    g0288(.A1(new_n233_), .A2(new_n126_), .ZN(new_n338_));
  NOR3_X1    g0289(.A1(new_n91_), .A2(new_n284_), .A3(new_n290_), .ZN(new_n339_));
  NOR4_X1    g0290(.A1(new_n263_), .A2(new_n338_), .A3(new_n339_), .A4(new_n337_), .ZN(new_n340_));
  NOR2_X1    g0291(.A1(new_n158_), .A2(new_n266_), .ZN(new_n341_));
  NOR2_X1    g0292(.A1(new_n164_), .A2(new_n341_), .ZN(new_n342_));
  AOI21_X1   g0293(.A1(new_n109_), .A2(new_n138_), .B(new_n126_), .ZN(new_n343_));
  INV_X1     g0294(.I(new_n343_), .ZN(new_n344_));
  NOR4_X1    g0295(.A1(new_n295_), .A2(new_n243_), .A3(new_n125_), .A4(new_n222_), .ZN(new_n345_));
  NOR2_X1    g0296(.A1(new_n204_), .A2(new_n266_), .ZN(new_n346_));
  NOR3_X1    g0297(.A1(new_n346_), .A2(new_n345_), .A3(new_n269_), .ZN(new_n347_));
  NAND3_X1   g0298(.A1(new_n347_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n348_));
  NOR3_X1    g0299(.A1(new_n348_), .A2(new_n201_), .A3(new_n208_), .ZN(new_n349_));
  NAND3_X1   g0300(.A1(new_n315_), .A2(new_n108_), .A3(new_n121_), .ZN(new_n350_));
  NAND2_X1   g0301(.A1(new_n235_), .A2(new_n239_), .ZN(new_n351_));
  NAND3_X1   g0302(.A1(new_n240_), .A2(new_n351_), .A3(new_n350_), .ZN(new_n352_));
  NOR2_X1    g0303(.A1(new_n178_), .A2(new_n126_), .ZN(new_n353_));
  NOR4_X1    g0304(.A1(new_n244_), .A2(new_n353_), .A3(new_n254_), .A4(new_n127_), .ZN(new_n354_));
  INV_X1     g0305(.I(new_n354_), .ZN(new_n355_));
  NOR2_X1    g0306(.A1(new_n155_), .A2(new_n266_), .ZN(new_n356_));
  NOR2_X1    g0307(.A1(new_n122_), .A2(new_n91_), .ZN(new_n357_));
  NOR4_X1    g0308(.A1(new_n355_), .A2(new_n352_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n358_));
  NAND2_X1   g0309(.A1(new_n162_), .A2(new_n115_), .ZN(new_n359_));
  NOR2_X1    g0310(.A1(new_n126_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1    g0311(.A1(new_n232_), .A2(new_n126_), .ZN(new_n361_));
  NOR4_X1    g0312(.A1(new_n267_), .A2(new_n156_), .A3(new_n361_), .A4(new_n360_), .ZN(new_n362_));
  NAND4_X1   g0313(.A1(new_n358_), .A2(new_n349_), .A3(new_n340_), .A4(new_n362_), .ZN(new_n363_));
  INV_X1     g0314(.I(new_n363_), .ZN(new_n364_));
  NAND2_X1   g0315(.A1(new_n335_), .A2(new_n364_), .ZN(new_n365_));
  NOR2_X1    g0316(.A1(new_n238_), .A2(new_n280_), .ZN(new_n366_));
  NAND3_X1   g0317(.A1(new_n229_), .A2(new_n366_), .A3(new_n125_), .ZN(new_n367_));
  NAND4_X1   g0318(.A1(new_n183_), .A2(new_n181_), .A3(new_n99_), .A4(new_n154_), .ZN(new_n368_));
  NAND3_X1   g0319(.A1(new_n239_), .A2(new_n183_), .A3(new_n181_), .ZN(new_n369_));
  NAND4_X1   g0320(.A1(new_n229_), .A2(new_n125_), .A3(new_n99_), .A4(new_n154_), .ZN(new_n370_));
  NAND4_X1   g0321(.A1(new_n370_), .A2(new_n367_), .A3(new_n368_), .A4(new_n369_), .ZN(new_n371_));
  NAND4_X1   g0322(.A1(new_n229_), .A2(new_n125_), .A3(new_n108_), .A4(new_n145_), .ZN(new_n372_));
  NOR2_X1    g0323(.A1(new_n192_), .A2(new_n232_), .ZN(new_n373_));
  INV_X1     g0324(.I(new_n373_), .ZN(new_n374_));
  NAND4_X1   g0325(.A1(new_n374_), .A2(new_n372_), .A3(new_n230_), .A4(new_n260_), .ZN(new_n375_));
  NOR2_X1    g0326(.A1(new_n359_), .A2(new_n203_), .ZN(new_n376_));
  NOR2_X1    g0327(.A1(new_n186_), .A2(new_n266_), .ZN(new_n377_));
  NOR2_X1    g0328(.A1(new_n122_), .A2(new_n266_), .ZN(new_n378_));
  NOR3_X1    g0329(.A1(new_n377_), .A2(new_n378_), .A3(new_n376_), .ZN(new_n379_));
  NOR2_X1    g0330(.A1(new_n202_), .A2(new_n188_), .ZN(new_n380_));
  NOR2_X1    g0331(.A1(new_n359_), .A2(new_n195_), .ZN(new_n381_));
  NOR3_X1    g0332(.A1(new_n232_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n382_));
  NOR2_X1    g0333(.A1(new_n382_), .A2(new_n381_), .ZN(new_n383_));
  NAND4_X1   g0334(.A1(new_n278_), .A2(new_n379_), .A3(new_n380_), .A4(new_n383_), .ZN(new_n384_));
  NOR2_X1    g0335(.A1(new_n384_), .A2(new_n375_), .ZN(new_n385_));
  NAND4_X1   g0336(.A1(new_n229_), .A2(new_n125_), .A3(new_n99_), .A4(new_n108_), .ZN(new_n386_));
  INV_X1     g0337(.I(new_n386_), .ZN(new_n387_));
  NOR2_X1    g0338(.A1(new_n192_), .A2(new_n158_), .ZN(new_n388_));
  NOR2_X1    g0339(.A1(new_n184_), .A2(new_n109_), .ZN(new_n389_));
  NOR4_X1    g0340(.A1(new_n387_), .A2(new_n197_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n390_));
  AND2_X2    g0341(.A1(new_n385_), .A2(new_n390_), .Z(new_n391_));
  NOR2_X1    g0342(.A1(new_n172_), .A2(new_n125_), .ZN(new_n392_));
  NAND3_X1   g0343(.A1(new_n392_), .A2(new_n137_), .A3(new_n145_), .ZN(new_n393_));
  NOR2_X1    g0344(.A1(new_n172_), .A2(new_n73_), .ZN(new_n394_));
  NAND3_X1   g0345(.A1(new_n394_), .A2(new_n99_), .A3(new_n108_), .ZN(new_n395_));
  AOI21_X1   g0346(.A1(new_n204_), .A2(new_n331_), .B(new_n172_), .ZN(new_n396_));
  INV_X1     g0347(.I(new_n396_), .ZN(new_n397_));
  NAND3_X1   g0348(.A1(new_n392_), .A2(new_n99_), .A3(new_n108_), .ZN(new_n398_));
  NAND4_X1   g0349(.A1(new_n397_), .A2(new_n393_), .A3(new_n395_), .A4(new_n398_), .ZN(new_n399_));
  NOR2_X1    g0350(.A1(new_n167_), .A2(new_n359_), .ZN(new_n400_));
  NOR2_X1    g0351(.A1(new_n158_), .A2(new_n195_), .ZN(new_n401_));
  NOR2_X1    g0352(.A1(new_n336_), .A2(new_n320_), .ZN(new_n402_));
  NOR3_X1    g0353(.A1(new_n401_), .A2(new_n402_), .A3(new_n400_), .ZN(new_n403_));
  NAND3_X1   g0354(.A1(new_n162_), .A2(new_n137_), .A3(new_n73_), .ZN(new_n404_));
  OAI22_X1   g0355(.A1(new_n233_), .A2(new_n266_), .B1(new_n404_), .B2(new_n320_), .ZN(new_n405_));
  INV_X1     g0356(.I(new_n405_), .ZN(new_n406_));
  NOR2_X1    g0357(.A1(new_n222_), .A2(new_n280_), .ZN(new_n407_));
  NAND2_X1   g0358(.A1(new_n227_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1    g0359(.A1(new_n295_), .A2(new_n222_), .ZN(new_n409_));
  NAND2_X1   g0360(.A1(new_n409_), .A2(new_n235_), .ZN(new_n410_));
  NAND2_X1   g0361(.A1(new_n410_), .A2(new_n408_), .ZN(new_n411_));
  NAND3_X1   g0362(.A1(new_n394_), .A2(new_n108_), .A3(new_n145_), .ZN(new_n412_));
  NAND2_X1   g0363(.A1(new_n303_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1    g0364(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1    g0365(.A1(new_n138_), .A2(new_n203_), .ZN(new_n415_));
  NAND3_X1   g0366(.A1(new_n394_), .A2(new_n137_), .A3(new_n145_), .ZN(new_n416_));
  NAND2_X1   g0367(.A1(new_n416_), .A2(new_n151_), .ZN(new_n417_));
  NOR4_X1    g0368(.A1(new_n417_), .A2(new_n200_), .A3(new_n265_), .A4(new_n415_), .ZN(new_n418_));
  NAND4_X1   g0369(.A1(new_n414_), .A2(new_n403_), .A3(new_n418_), .A4(new_n406_), .ZN(new_n419_));
  NOR2_X1    g0370(.A1(new_n419_), .A2(new_n399_), .ZN(new_n420_));
  NAND2_X1   g0371(.A1(new_n391_), .A2(new_n420_), .ZN(new_n421_));
  NOR2_X1    g0372(.A1(new_n421_), .A2(new_n371_), .ZN(new_n422_));
  INV_X1     g0373(.I(new_n422_), .ZN(new_n423_));
  NOR2_X1    g0374(.A1(new_n377_), .A2(new_n378_), .ZN(new_n424_));
  NOR2_X1    g0375(.A1(new_n138_), .A2(new_n195_), .ZN(new_n425_));
  NOR2_X1    g0376(.A1(new_n178_), .A2(new_n203_), .ZN(new_n426_));
  NOR2_X1    g0377(.A1(new_n426_), .A2(new_n425_), .ZN(new_n427_));
  INV_X1     g0378(.I(new_n427_), .ZN(new_n428_));
  NAND2_X1   g0379(.A1(new_n394_), .A2(new_n239_), .ZN(new_n429_));
  NAND2_X1   g0380(.A1(new_n429_), .A2(new_n190_), .ZN(new_n430_));
  NAND3_X1   g0381(.A1(new_n392_), .A2(new_n121_), .A3(new_n137_), .ZN(new_n431_));
  NAND2_X1   g0382(.A1(new_n392_), .A2(new_n239_), .ZN(new_n432_));
  NAND3_X1   g0383(.A1(new_n394_), .A2(new_n99_), .A3(new_n154_), .ZN(new_n433_));
  NAND3_X1   g0384(.A1(new_n431_), .A2(new_n433_), .A3(new_n432_), .ZN(new_n434_));
  NOR2_X1    g0385(.A1(new_n186_), .A2(new_n203_), .ZN(new_n435_));
  INV_X1     g0386(.I(new_n435_), .ZN(new_n436_));
  NOR2_X1    g0387(.A1(new_n178_), .A2(new_n195_), .ZN(new_n437_));
  INV_X1     g0388(.I(new_n437_), .ZN(new_n438_));
  NAND3_X1   g0389(.A1(new_n394_), .A2(new_n121_), .A3(new_n137_), .ZN(new_n439_));
  NAND3_X1   g0390(.A1(new_n438_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  NOR4_X1    g0391(.A1(new_n440_), .A2(new_n428_), .A3(new_n430_), .A4(new_n434_), .ZN(new_n441_));
  AND4_X2    g0392(.A1(new_n424_), .A2(new_n420_), .A3(new_n380_), .A4(new_n441_), .Z(new_n442_));
  NOR4_X1    g0393(.A1(new_n290_), .A2(new_n125_), .A3(new_n172_), .A4(new_n222_), .ZN(new_n443_));
  NOR2_X1    g0394(.A1(new_n122_), .A2(new_n203_), .ZN(new_n444_));
  NOR2_X1    g0395(.A1(new_n444_), .A2(new_n299_), .ZN(new_n445_));
  INV_X1     g0396(.I(new_n445_), .ZN(new_n446_));
  NAND2_X1   g0397(.A1(new_n394_), .A2(new_n407_), .ZN(new_n447_));
  INV_X1     g0398(.I(new_n447_), .ZN(new_n448_));
  NOR4_X1    g0399(.A1(new_n446_), .A2(new_n246_), .A3(new_n443_), .A4(new_n448_), .ZN(new_n449_));
  NOR4_X1    g0400(.A1(new_n172_), .A2(new_n222_), .A3(new_n280_), .A4(new_n125_), .ZN(new_n450_));
  INV_X1     g0401(.I(new_n450_), .ZN(new_n451_));
  NOR2_X1    g0402(.A1(new_n225_), .A2(new_n172_), .ZN(new_n452_));
  NAND3_X1   g0403(.A1(new_n394_), .A2(new_n115_), .A3(new_n121_), .ZN(new_n453_));
  INV_X1     g0404(.I(new_n453_), .ZN(new_n454_));
  NOR2_X1    g0405(.A1(new_n454_), .A2(new_n452_), .ZN(new_n455_));
  NAND3_X1   g0406(.A1(new_n449_), .A2(new_n451_), .A3(new_n455_), .ZN(new_n456_));
  NOR2_X1    g0407(.A1(new_n456_), .A2(new_n291_), .ZN(new_n457_));
  NAND2_X1   g0408(.A1(new_n442_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1   g0409(.A1(new_n423_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1     g0410(.I(\a[13] ), .ZN(new_n460_));
  NAND2_X1   g0411(.A1(new_n69_), .A2(new_n57_), .ZN(new_n461_));
  XOR2_X1    g0412(.A1(new_n461_), .A2(new_n460_), .Z(new_n462_));
  INV_X1     g0413(.I(\a[14] ), .ZN(new_n463_));
  OAI21_X1   g0414(.A1(new_n69_), .A2(\a[13] ), .B(new_n57_), .ZN(new_n464_));
  XOR2_X1    g0415(.A1(new_n464_), .A2(new_n463_), .Z(new_n465_));
  XOR2_X1    g0416(.A1(new_n465_), .A2(new_n462_), .Z(new_n466_));
  XOR2_X1    g0417(.A1(new_n459_), .A2(new_n466_), .Z(new_n467_));
  NAND2_X1   g0418(.A1(new_n467_), .A2(new_n365_), .ZN(new_n468_));
  INV_X1     g0419(.I(new_n365_), .ZN(new_n469_));
  INV_X1     g0420(.I(new_n111_), .ZN(new_n470_));
  NOR2_X1    g0421(.A1(new_n470_), .A2(\a[10] ), .ZN(new_n471_));
  NOR2_X1    g0422(.A1(new_n471_), .A2(\a[22] ), .ZN(new_n472_));
  XOR2_X1    g0423(.A1(new_n472_), .A2(\a[11] ), .Z(new_n473_));
  INV_X1     g0424(.I(new_n473_), .ZN(new_n474_));
  INV_X1     g0425(.I(\a[11] ), .ZN(new_n475_));
  AOI21_X1   g0426(.A1(new_n471_), .A2(new_n475_), .B(\a[22] ), .ZN(new_n476_));
  XOR2_X1    g0427(.A1(new_n476_), .A2(\a[12] ), .Z(new_n477_));
  INV_X1     g0428(.I(new_n477_), .ZN(new_n478_));
  NOR2_X1    g0429(.A1(new_n478_), .A2(new_n474_), .ZN(new_n479_));
  INV_X1     g0430(.I(new_n479_), .ZN(new_n480_));
  NAND4_X1   g0431(.A1(new_n183_), .A2(new_n181_), .A3(new_n145_), .A4(new_n154_), .ZN(new_n481_));
  AOI21_X1   g0432(.A1(new_n215_), .A2(new_n212_), .B(new_n73_), .ZN(new_n482_));
  NAND3_X1   g0433(.A1(new_n482_), .A2(new_n108_), .A3(new_n121_), .ZN(new_n483_));
  NAND3_X1   g0434(.A1(new_n481_), .A2(new_n316_), .A3(new_n483_), .ZN(new_n484_));
  NOR2_X1    g0435(.A1(new_n192_), .A2(new_n204_), .ZN(new_n485_));
  NOR2_X1    g0436(.A1(new_n485_), .A2(new_n400_), .ZN(new_n486_));
  OAI22_X1   g0437(.A1(new_n163_), .A2(new_n266_), .B1(new_n186_), .B2(new_n203_), .ZN(new_n487_));
  INV_X1     g0438(.I(new_n487_), .ZN(new_n488_));
  NAND2_X1   g0439(.A1(new_n488_), .A2(new_n486_), .ZN(new_n489_));
  NOR3_X1    g0440(.A1(new_n222_), .A2(new_n280_), .A3(new_n125_), .ZN(new_n490_));
  NAND2_X1   g0441(.A1(new_n302_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1    g0442(.A1(new_n209_), .A2(new_n167_), .ZN(new_n492_));
  NOR2_X1    g0443(.A1(new_n492_), .A2(new_n360_), .ZN(new_n493_));
  NOR2_X1    g0444(.A1(new_n249_), .A2(new_n203_), .ZN(new_n494_));
  NOR3_X1    g0445(.A1(new_n126_), .A2(new_n295_), .A3(new_n284_), .ZN(new_n495_));
  NOR3_X1    g0446(.A1(new_n332_), .A2(new_n495_), .A3(new_n494_), .ZN(new_n496_));
  NOR2_X1    g0447(.A1(new_n155_), .A2(new_n195_), .ZN(new_n497_));
  NOR2_X1    g0448(.A1(new_n497_), .A2(new_n339_), .ZN(new_n498_));
  NAND4_X1   g0449(.A1(new_n496_), .A2(new_n493_), .A3(new_n498_), .A4(new_n491_), .ZN(new_n499_));
  NOR2_X1    g0450(.A1(new_n188_), .A2(new_n159_), .ZN(new_n500_));
  NAND3_X1   g0451(.A1(new_n500_), .A2(new_n372_), .A3(new_n255_), .ZN(new_n501_));
  NOR4_X1    g0452(.A1(new_n499_), .A2(new_n489_), .A3(new_n484_), .A4(new_n501_), .ZN(new_n502_));
  NOR2_X1    g0453(.A1(new_n178_), .A2(new_n91_), .ZN(new_n503_));
  NOR2_X1    g0454(.A1(new_n312_), .A2(new_n337_), .ZN(new_n504_));
  INV_X1     g0455(.I(new_n504_), .ZN(new_n505_));
  NOR3_X1    g0456(.A1(new_n505_), .A2(new_n191_), .A3(new_n503_), .ZN(new_n506_));
  NOR3_X1    g0457(.A1(new_n338_), .A2(new_n207_), .A3(new_n196_), .ZN(new_n507_));
  NOR2_X1    g0458(.A1(new_n276_), .A2(new_n200_), .ZN(new_n508_));
  NOR3_X1    g0459(.A1(new_n122_), .A2(new_n135_), .A3(new_n73_), .ZN(new_n509_));
  NOR4_X1    g0460(.A1(new_n187_), .A2(new_n378_), .A3(new_n509_), .A4(new_n402_), .ZN(new_n510_));
  NAND4_X1   g0461(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1     g0462(.I(new_n202_), .ZN(new_n512_));
  NOR2_X1    g0463(.A1(new_n286_), .A2(new_n219_), .ZN(new_n513_));
  OAI21_X1   g0464(.A1(new_n513_), .A2(new_n407_), .B(new_n315_), .ZN(new_n514_));
  NOR2_X1    g0465(.A1(new_n249_), .A2(new_n167_), .ZN(new_n515_));
  NOR2_X1    g0466(.A1(new_n184_), .A2(new_n178_), .ZN(new_n516_));
  NOR3_X1    g0467(.A1(new_n516_), .A2(new_n110_), .A3(new_n515_), .ZN(new_n517_));
  NAND4_X1   g0468(.A1(new_n517_), .A2(new_n512_), .A3(new_n383_), .A4(new_n514_), .ZN(new_n518_));
  INV_X1     g0469(.I(new_n234_), .ZN(new_n519_));
  NOR4_X1    g0470(.A1(new_n193_), .A2(new_n377_), .A3(new_n437_), .A4(new_n127_), .ZN(new_n520_));
  NOR3_X1    g0471(.A1(new_n343_), .A2(new_n164_), .A3(new_n361_), .ZN(new_n521_));
  NAND4_X1   g0472(.A1(new_n520_), .A2(new_n519_), .A3(new_n521_), .A4(new_n427_), .ZN(new_n522_));
  NOR2_X1    g0473(.A1(new_n522_), .A2(new_n518_), .ZN(new_n523_));
  NOR3_X1    g0474(.A1(new_n135_), .A2(new_n194_), .A3(new_n73_), .ZN(new_n524_));
  NOR2_X1    g0475(.A1(new_n294_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1    g0476(.A1(new_n185_), .A2(new_n373_), .ZN(new_n526_));
  INV_X1     g0477(.I(new_n526_), .ZN(new_n527_));
  NAND2_X1   g0478(.A1(new_n392_), .A2(new_n223_), .ZN(new_n528_));
  NAND2_X1   g0479(.A1(new_n157_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1   g0480(.A1(new_n216_), .A2(new_n73_), .A3(new_n121_), .A4(new_n137_), .ZN(new_n530_));
  INV_X1     g0481(.I(new_n250_), .ZN(new_n531_));
  NAND4_X1   g0482(.A1(new_n531_), .A2(new_n530_), .A3(new_n432_), .A4(new_n439_), .ZN(new_n532_));
  NOR4_X1    g0483(.A1(new_n527_), .A2(new_n532_), .A3(new_n317_), .A4(new_n529_), .ZN(new_n533_));
  NAND3_X1   g0484(.A1(new_n523_), .A2(new_n525_), .A3(new_n533_), .ZN(new_n534_));
  NOR2_X1    g0485(.A1(new_n534_), .A2(new_n511_), .ZN(new_n535_));
  NOR2_X1    g0486(.A1(new_n233_), .A2(new_n266_), .ZN(new_n536_));
  NOR3_X1    g0487(.A1(new_n274_), .A2(new_n345_), .A3(new_n536_), .ZN(new_n537_));
  NAND3_X1   g0488(.A1(new_n535_), .A2(new_n502_), .A3(new_n537_), .ZN(new_n538_));
  NOR2_X1    g0489(.A1(new_n252_), .A2(new_n251_), .ZN(new_n539_));
  NAND2_X1   g0490(.A1(new_n539_), .A2(new_n366_), .ZN(new_n540_));
  NOR2_X1    g0491(.A1(new_n495_), .A2(new_n444_), .ZN(new_n541_));
  NAND4_X1   g0492(.A1(new_n541_), .A2(new_n429_), .A3(new_n540_), .A4(new_n433_), .ZN(new_n542_));
  NOR3_X1    g0493(.A1(new_n244_), .A2(new_n313_), .A3(new_n378_), .ZN(new_n543_));
  NOR4_X1    g0494(.A1(new_n295_), .A2(new_n284_), .A3(new_n125_), .A4(new_n172_), .ZN(new_n544_));
  NOR2_X1    g0495(.A1(new_n163_), .A2(new_n266_), .ZN(new_n545_));
  NOR4_X1    g0496(.A1(new_n388_), .A2(new_n544_), .A3(new_n545_), .A4(new_n207_), .ZN(new_n546_));
  NAND2_X1   g0497(.A1(new_n546_), .A2(new_n543_), .ZN(new_n547_));
  NOR3_X1    g0498(.A1(new_n295_), .A2(new_n284_), .A3(new_n195_), .ZN(new_n548_));
  INV_X1     g0499(.I(new_n432_), .ZN(new_n549_));
  NOR3_X1    g0500(.A1(new_n549_), .A2(new_n381_), .A3(new_n548_), .ZN(new_n550_));
  NAND4_X1   g0501(.A1(new_n229_), .A2(new_n125_), .A3(new_n108_), .A4(new_n162_), .ZN(new_n551_));
  INV_X1     g0502(.I(new_n551_), .ZN(new_n552_));
  NOR2_X1    g0503(.A1(new_n552_), .A2(new_n341_), .ZN(new_n553_));
  NAND4_X1   g0504(.A1(new_n553_), .A2(new_n206_), .A3(new_n550_), .A4(new_n255_), .ZN(new_n554_));
  INV_X1     g0505(.I(new_n377_), .ZN(new_n555_));
  NAND2_X1   g0506(.A1(new_n394_), .A2(new_n366_), .ZN(new_n556_));
  NOR2_X1    g0507(.A1(new_n266_), .A2(new_n138_), .ZN(new_n557_));
  NOR3_X1    g0508(.A1(new_n524_), .A2(new_n327_), .A3(new_n557_), .ZN(new_n558_));
  NAND3_X1   g0509(.A1(new_n558_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n559_));
  NOR4_X1    g0510(.A1(new_n554_), .A2(new_n542_), .A3(new_n547_), .A4(new_n559_), .ZN(new_n560_));
  NOR2_X1    g0511(.A1(new_n91_), .A2(new_n194_), .ZN(new_n561_));
  NOR3_X1    g0512(.A1(new_n503_), .A2(new_n353_), .A3(new_n156_), .ZN(new_n562_));
  NAND3_X1   g0513(.A1(new_n394_), .A2(new_n121_), .A3(new_n154_), .ZN(new_n563_));
  NAND2_X1   g0514(.A1(new_n393_), .A2(new_n563_), .ZN(new_n564_));
  NAND4_X1   g0515(.A1(new_n183_), .A2(new_n181_), .A3(new_n108_), .A4(new_n121_), .ZN(new_n565_));
  NAND3_X1   g0516(.A1(new_n315_), .A2(new_n137_), .A3(new_n145_), .ZN(new_n566_));
  NAND2_X1   g0517(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR3_X1    g0518(.A1(new_n564_), .A2(new_n567_), .A3(new_n343_), .ZN(new_n568_));
  OAI22_X1   g0519(.A1(new_n204_), .A2(new_n126_), .B1(new_n232_), .B2(new_n195_), .ZN(new_n569_));
  NOR4_X1    g0520(.A1(new_n569_), .A2(new_n259_), .A3(new_n317_), .A4(new_n330_), .ZN(new_n570_));
  NAND3_X1   g0521(.A1(new_n568_), .A2(new_n570_), .A3(new_n562_), .ZN(new_n571_));
  NOR3_X1    g0522(.A1(new_n571_), .A2(new_n561_), .A3(new_n454_), .ZN(new_n572_));
  NOR3_X1    g0523(.A1(new_n270_), .A2(new_n252_), .A3(new_n251_), .ZN(new_n573_));
  NOR2_X1    g0524(.A1(new_n250_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1    g0525(.A1(new_n286_), .A2(new_n290_), .ZN(new_n575_));
  OAI21_X1   g0526(.A1(new_n315_), .A2(new_n482_), .B(new_n575_), .ZN(new_n576_));
  NAND3_X1   g0527(.A1(new_n574_), .A2(new_n576_), .A3(new_n372_), .ZN(new_n577_));
  NAND3_X1   g0528(.A1(new_n482_), .A2(new_n137_), .A3(new_n145_), .ZN(new_n578_));
  NOR3_X1    g0529(.A1(new_n389_), .A2(new_n208_), .A3(new_n346_), .ZN(new_n579_));
  NOR3_X1    g0530(.A1(new_n135_), .A2(new_n270_), .A3(new_n73_), .ZN(new_n580_));
  INV_X1     g0531(.I(new_n580_), .ZN(new_n581_));
  NAND4_X1   g0532(.A1(new_n579_), .A2(new_n303_), .A3(new_n578_), .A4(new_n581_), .ZN(new_n582_));
  NAND4_X1   g0533(.A1(new_n216_), .A2(new_n73_), .A3(new_n145_), .A4(new_n115_), .ZN(new_n583_));
  NOR3_X1    g0534(.A1(new_n168_), .A2(new_n339_), .A3(new_n376_), .ZN(new_n584_));
  NOR2_X1    g0535(.A1(new_n387_), .A2(new_n191_), .ZN(new_n585_));
  NAND4_X1   g0536(.A1(new_n585_), .A2(new_n584_), .A3(new_n500_), .A4(new_n583_), .ZN(new_n586_));
  NOR2_X1    g0537(.A1(new_n184_), .A2(new_n163_), .ZN(new_n587_));
  NOR3_X1    g0538(.A1(new_n261_), .A2(new_n587_), .A3(new_n452_), .ZN(new_n588_));
  NOR3_X1    g0539(.A1(new_n294_), .A2(new_n110_), .A3(new_n269_), .ZN(new_n589_));
  NAND2_X1   g0540(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NOR4_X1    g0541(.A1(new_n586_), .A2(new_n582_), .A3(new_n577_), .A4(new_n590_), .ZN(new_n591_));
  NAND3_X1   g0542(.A1(new_n560_), .A2(new_n591_), .A3(new_n572_), .ZN(new_n592_));
  NAND2_X1   g0543(.A1(new_n538_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1   g0544(.A1(new_n593_), .A2(new_n423_), .ZN(new_n594_));
  OAI21_X1   g0545(.A1(new_n473_), .A2(new_n477_), .B(new_n594_), .ZN(new_n595_));
  AOI21_X1   g0546(.A1(new_n595_), .A2(new_n480_), .B(new_n469_), .ZN(new_n596_));
  INV_X1     g0547(.I(new_n596_), .ZN(new_n597_));
  INV_X1     g0548(.I(new_n465_), .ZN(new_n598_));
  INV_X1     g0549(.I(new_n458_), .ZN(new_n599_));
  NAND2_X1   g0550(.A1(new_n599_), .A2(new_n365_), .ZN(new_n600_));
  NAND2_X1   g0551(.A1(new_n469_), .A2(new_n458_), .ZN(new_n601_));
  OAI21_X1   g0552(.A1(new_n598_), .A2(new_n601_), .B(new_n600_), .ZN(new_n602_));
  NOR2_X1    g0553(.A1(new_n599_), .A2(new_n423_), .ZN(new_n603_));
  NOR2_X1    g0554(.A1(new_n458_), .A2(new_n465_), .ZN(new_n604_));
  OR2_X2     g0555(.A1(new_n603_), .A2(new_n604_), .Z(new_n605_));
  AOI22_X1   g0556(.A1(new_n602_), .A2(new_n423_), .B1(new_n605_), .B2(new_n365_), .ZN(new_n606_));
  AND2_X2    g0557(.A1(new_n606_), .A2(new_n597_), .Z(new_n607_));
  NAND2_X1   g0558(.A1(new_n365_), .A2(new_n462_), .ZN(new_n608_));
  NOR2_X1    g0559(.A1(new_n606_), .A2(new_n597_), .ZN(new_n609_));
  NOR2_X1    g0560(.A1(new_n609_), .A2(new_n608_), .ZN(new_n610_));
  NOR2_X1    g0561(.A1(new_n610_), .A2(new_n607_), .ZN(new_n611_));
  XOR2_X1    g0562(.A1(new_n611_), .A2(new_n468_), .Z(new_n612_));
  NAND2_X1   g0563(.A1(new_n599_), .A2(new_n422_), .ZN(new_n613_));
  NAND2_X1   g0564(.A1(new_n613_), .A2(new_n459_), .ZN(new_n614_));
  NOR2_X1    g0565(.A1(new_n423_), .A2(new_n458_), .ZN(new_n615_));
  NOR2_X1    g0566(.A1(new_n615_), .A2(new_n365_), .ZN(new_n616_));
  INV_X1     g0567(.I(new_n616_), .ZN(new_n617_));
  NAND2_X1   g0568(.A1(new_n617_), .A2(new_n614_), .ZN(new_n618_));
  NAND2_X1   g0569(.A1(new_n618_), .A2(new_n462_), .ZN(new_n619_));
  INV_X1     g0570(.I(new_n462_), .ZN(new_n620_));
  NAND2_X1   g0571(.A1(new_n614_), .A2(new_n600_), .ZN(new_n621_));
  NAND2_X1   g0572(.A1(new_n621_), .A2(new_n620_), .ZN(new_n622_));
  INV_X1     g0573(.I(new_n459_), .ZN(new_n623_));
  NOR2_X1    g0574(.A1(new_n623_), .A2(new_n615_), .ZN(new_n624_));
  NAND2_X1   g0575(.A1(new_n617_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1   g0576(.A1(new_n625_), .A2(new_n465_), .ZN(new_n626_));
  XNOR2_X1   g0577(.A1(new_n458_), .A2(new_n422_), .ZN(new_n627_));
  NAND2_X1   g0578(.A1(new_n627_), .A2(new_n469_), .ZN(new_n628_));
  NAND2_X1   g0579(.A1(new_n628_), .A2(new_n598_), .ZN(new_n629_));
  AOI22_X1   g0580(.A1(new_n619_), .A2(new_n622_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1   g0581(.A1(new_n477_), .A2(new_n473_), .ZN(new_n631_));
  NOR2_X1    g0582(.A1(new_n469_), .A2(new_n631_), .ZN(new_n632_));
  XOR2_X1    g0583(.A1(new_n594_), .A2(new_n632_), .Z(new_n633_));
  NOR2_X1    g0584(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1    g0585(.A1(new_n422_), .A2(new_n592_), .ZN(new_n635_));
  INV_X1     g0586(.I(new_n592_), .ZN(new_n636_));
  NOR3_X1    g0587(.A1(new_n423_), .A2(new_n598_), .A3(new_n636_), .ZN(new_n637_));
  OAI21_X1   g0588(.A1(new_n637_), .A2(new_n635_), .B(new_n538_), .ZN(new_n638_));
  INV_X1     g0589(.I(new_n638_), .ZN(new_n639_));
  AOI21_X1   g0590(.A1(new_n465_), .A2(new_n636_), .B(new_n594_), .ZN(new_n640_));
  NOR2_X1    g0591(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1    g0592(.A1(new_n469_), .A2(new_n474_), .ZN(new_n642_));
  NAND2_X1   g0593(.A1(new_n618_), .A2(new_n477_), .ZN(new_n643_));
  NAND2_X1   g0594(.A1(new_n621_), .A2(new_n478_), .ZN(new_n644_));
  NAND2_X1   g0595(.A1(new_n625_), .A2(new_n462_), .ZN(new_n645_));
  NAND2_X1   g0596(.A1(new_n628_), .A2(new_n620_), .ZN(new_n646_));
  AOI22_X1   g0597(.A1(new_n643_), .A2(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NOR2_X1    g0598(.A1(new_n641_), .A2(new_n642_), .ZN(new_n648_));
  NOR2_X1    g0599(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1   g0600(.A1(new_n641_), .A2(new_n642_), .B(new_n649_), .ZN(new_n650_));
  AOI21_X1   g0601(.A1(new_n630_), .A2(new_n633_), .B(new_n650_), .ZN(new_n651_));
  NOR2_X1    g0602(.A1(new_n651_), .A2(new_n634_), .ZN(new_n652_));
  NOR2_X1    g0603(.A1(new_n607_), .A2(new_n609_), .ZN(new_n653_));
  XOR2_X1    g0604(.A1(new_n653_), .A2(new_n608_), .Z(new_n654_));
  NOR2_X1    g0605(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1   g0606(.A1(new_n652_), .A2(new_n654_), .ZN(new_n656_));
  INV_X1     g0607(.I(new_n656_), .ZN(new_n657_));
  XNOR2_X1   g0608(.A1(new_n641_), .A2(new_n642_), .ZN(new_n658_));
  XOR2_X1    g0609(.A1(new_n658_), .A2(new_n647_), .Z(new_n659_));
  INV_X1     g0610(.I(new_n60_), .ZN(new_n660_));
  OR2_X2     g0611(.A1(\a[7] ), .A2(\a[8] ), .Z(new_n661_));
  OAI21_X1   g0612(.A1(new_n660_), .A2(new_n661_), .B(new_n57_), .ZN(new_n662_));
  XNOR2_X1   g0613(.A1(new_n662_), .A2(\a[9] ), .ZN(new_n663_));
  INV_X1     g0614(.I(new_n663_), .ZN(new_n664_));
  INV_X1     g0615(.I(\a[10] ), .ZN(new_n665_));
  NAND2_X1   g0616(.A1(new_n470_), .A2(new_n57_), .ZN(new_n666_));
  NAND2_X1   g0617(.A1(new_n666_), .A2(new_n665_), .ZN(new_n667_));
  INV_X1     g0618(.I(new_n667_), .ZN(new_n668_));
  NOR2_X1    g0619(.A1(new_n666_), .A2(new_n665_), .ZN(new_n669_));
  NOR2_X1    g0620(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1     g0621(.I(new_n670_), .ZN(new_n671_));
  NOR2_X1    g0622(.A1(new_n671_), .A2(new_n664_), .ZN(new_n672_));
  INV_X1     g0623(.I(new_n672_), .ZN(new_n673_));
  NAND3_X1   g0624(.A1(new_n227_), .A2(new_n145_), .A3(new_n154_), .ZN(new_n674_));
  INV_X1     g0625(.I(new_n245_), .ZN(new_n675_));
  NAND3_X1   g0626(.A1(new_n394_), .A2(new_n108_), .A3(new_n162_), .ZN(new_n676_));
  NAND4_X1   g0627(.A1(new_n216_), .A2(new_n108_), .A3(new_n73_), .A4(new_n162_), .ZN(new_n677_));
  NAND4_X1   g0628(.A1(new_n675_), .A2(new_n674_), .A3(new_n676_), .A4(new_n677_), .ZN(new_n678_));
  NOR4_X1    g0629(.A1(new_n191_), .A2(new_n253_), .A3(new_n341_), .A4(new_n548_), .ZN(new_n679_));
  NOR3_X1    g0630(.A1(new_n388_), .A2(new_n339_), .A3(new_n401_), .ZN(new_n680_));
  NAND3_X1   g0631(.A1(new_n680_), .A2(new_n679_), .A3(new_n273_), .ZN(new_n681_));
  NAND2_X1   g0632(.A1(new_n374_), .A2(new_n236_), .ZN(new_n682_));
  NOR4_X1    g0633(.A1(new_n681_), .A2(new_n161_), .A3(new_n678_), .A4(new_n682_), .ZN(new_n683_));
  NAND4_X1   g0634(.A1(new_n183_), .A2(new_n181_), .A3(new_n108_), .A4(new_n99_), .ZN(new_n684_));
  NAND4_X1   g0635(.A1(new_n183_), .A2(new_n181_), .A3(new_n154_), .A4(new_n162_), .ZN(new_n685_));
  NAND4_X1   g0636(.A1(new_n528_), .A2(new_n684_), .A3(new_n685_), .A4(new_n447_), .ZN(new_n686_));
  NOR3_X1    g0637(.A1(new_n284_), .A2(new_n290_), .A3(new_n195_), .ZN(new_n687_));
  NOR4_X1    g0638(.A1(new_n587_), .A2(new_n277_), .A3(new_n327_), .A4(new_n687_), .ZN(new_n688_));
  INV_X1     g0639(.I(new_n688_), .ZN(new_n689_));
  NOR2_X1    g0640(.A1(new_n552_), .A2(new_n536_), .ZN(new_n690_));
  NOR2_X1    g0641(.A1(new_n192_), .A2(new_n233_), .ZN(new_n691_));
  NOR3_X1    g0642(.A1(new_n564_), .A2(new_n139_), .A3(new_n691_), .ZN(new_n692_));
  NOR2_X1    g0643(.A1(new_n404_), .A2(new_n320_), .ZN(new_n693_));
  NOR2_X1    g0644(.A1(new_n187_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1    g0645(.A1(new_n158_), .A2(new_n203_), .ZN(new_n695_));
  NOR2_X1    g0646(.A1(new_n695_), .A2(new_n450_), .ZN(new_n696_));
  NAND4_X1   g0647(.A1(new_n692_), .A2(new_n690_), .A3(new_n694_), .A4(new_n696_), .ZN(new_n697_));
  NOR2_X1    g0648(.A1(new_n266_), .A2(new_n194_), .ZN(new_n698_));
  NOR2_X1    g0649(.A1(new_n263_), .A2(new_n698_), .ZN(new_n699_));
  OAI22_X1   g0650(.A1(new_n331_), .A2(new_n243_), .B1(new_n155_), .B2(new_n266_), .ZN(new_n700_));
  INV_X1     g0651(.I(new_n700_), .ZN(new_n701_));
  NOR2_X1    g0652(.A1(new_n346_), .A2(new_n254_), .ZN(new_n702_));
  NAND4_X1   g0653(.A1(new_n701_), .A2(new_n699_), .A3(new_n702_), .A4(new_n541_), .ZN(new_n703_));
  NOR4_X1    g0654(.A1(new_n697_), .A2(new_n686_), .A3(new_n689_), .A4(new_n703_), .ZN(new_n704_));
  NAND4_X1   g0655(.A1(new_n704_), .A2(new_n523_), .A3(new_n525_), .A4(new_n683_), .ZN(new_n705_));
  NAND3_X1   g0656(.A1(new_n676_), .A2(new_n260_), .A3(new_n398_), .ZN(new_n706_));
  NOR4_X1    g0657(.A1(new_n706_), .A2(new_n310_), .A3(new_n387_), .A4(new_n503_), .ZN(new_n707_));
  NOR4_X1    g0658(.A1(new_n587_), .A2(new_n127_), .A3(new_n330_), .A4(new_n327_), .ZN(new_n708_));
  NOR2_X1    g0659(.A1(new_n346_), .A2(new_n265_), .ZN(new_n709_));
  NAND3_X1   g0660(.A1(new_n315_), .A2(new_n115_), .A3(new_n121_), .ZN(new_n710_));
  NAND2_X1   g0661(.A1(new_n431_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1    g0662(.A1(new_n711_), .A2(new_n337_), .ZN(new_n712_));
  NAND4_X1   g0663(.A1(new_n708_), .A2(new_n712_), .A3(new_n491_), .A4(new_n709_), .ZN(new_n713_));
  NAND2_X1   g0664(.A1(new_n223_), .A2(new_n482_), .ZN(new_n714_));
  NAND2_X1   g0665(.A1(new_n453_), .A2(new_n714_), .ZN(new_n715_));
  NOR3_X1    g0666(.A1(new_n715_), .A2(new_n139_), .A3(new_n388_), .ZN(new_n716_));
  NAND3_X1   g0667(.A1(new_n223_), .A2(new_n183_), .A3(new_n181_), .ZN(new_n717_));
  INV_X1     g0668(.I(new_n717_), .ZN(new_n718_));
  NOR4_X1    g0669(.A1(new_n718_), .A2(new_n338_), .A3(new_n345_), .A4(new_n687_), .ZN(new_n719_));
  NAND2_X1   g0670(.A1(new_n716_), .A2(new_n719_), .ZN(new_n720_));
  NOR2_X1    g0671(.A1(new_n713_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1    g0672(.A1(new_n167_), .A2(new_n194_), .ZN(new_n722_));
  NOR3_X1    g0673(.A1(new_n155_), .A2(new_n135_), .A3(new_n73_), .ZN(new_n723_));
  NOR3_X1    g0674(.A1(new_n256_), .A2(new_n723_), .A3(new_n722_), .ZN(new_n724_));
  NAND2_X1   g0675(.A1(new_n724_), .A2(new_n189_), .ZN(new_n725_));
  NAND2_X1   g0676(.A1(new_n316_), .A2(new_n483_), .ZN(new_n726_));
  NAND2_X1   g0677(.A1(new_n303_), .A2(new_n563_), .ZN(new_n727_));
  NOR4_X1    g0678(.A1(new_n727_), .A2(new_n726_), .A3(new_n201_), .A4(new_n245_), .ZN(new_n728_));
  NOR2_X1    g0679(.A1(new_n232_), .A2(new_n195_), .ZN(new_n729_));
  NAND2_X1   g0680(.A1(new_n230_), .A2(new_n151_), .ZN(new_n730_));
  OAI21_X1   g0681(.A1(new_n249_), .A2(new_n184_), .B(new_n432_), .ZN(new_n731_));
  NOR4_X1    g0682(.A1(new_n731_), .A2(new_n730_), .A3(new_n164_), .A4(new_n729_), .ZN(new_n732_));
  NAND2_X1   g0683(.A1(new_n732_), .A2(new_n728_), .ZN(new_n733_));
  NOR2_X1    g0684(.A1(new_n733_), .A2(new_n725_), .ZN(new_n734_));
  INV_X1     g0685(.I(new_n379_), .ZN(new_n735_));
  NOR3_X1    g0686(.A1(new_n233_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n736_));
  NOR4_X1    g0687(.A1(new_n313_), .A2(new_n736_), .A3(new_n356_), .A4(new_n425_), .ZN(new_n737_));
  INV_X1     g0688(.I(new_n737_), .ZN(new_n738_));
  NAND4_X1   g0689(.A1(new_n108_), .A2(new_n121_), .A3(new_n73_), .A4(new_n150_), .ZN(new_n739_));
  NAND3_X1   g0690(.A1(new_n407_), .A2(new_n183_), .A3(new_n181_), .ZN(new_n740_));
  NOR2_X1    g0691(.A1(new_n373_), .A2(new_n177_), .ZN(new_n741_));
  NAND4_X1   g0692(.A1(new_n741_), .A2(new_n739_), .A3(new_n740_), .A4(new_n696_), .ZN(new_n742_));
  INV_X1     g0693(.I(new_n207_), .ZN(new_n743_));
  NAND4_X1   g0694(.A1(new_n183_), .A2(new_n181_), .A3(new_n137_), .A4(new_n145_), .ZN(new_n744_));
  NOR2_X1    g0695(.A1(new_n249_), .A2(new_n195_), .ZN(new_n745_));
  NOR4_X1    g0696(.A1(new_n524_), .A2(new_n497_), .A3(new_n745_), .A4(new_n443_), .ZN(new_n746_));
  NAND3_X1   g0697(.A1(new_n746_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n747_));
  NOR4_X1    g0698(.A1(new_n742_), .A2(new_n747_), .A3(new_n735_), .A4(new_n738_), .ZN(new_n748_));
  NAND4_X1   g0699(.A1(new_n734_), .A2(new_n721_), .A3(new_n748_), .A4(new_n707_), .ZN(new_n749_));
  NAND2_X1   g0700(.A1(new_n705_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1   g0701(.A1(new_n750_), .A2(new_n592_), .ZN(new_n751_));
  INV_X1     g0702(.I(new_n751_), .ZN(new_n752_));
  NOR2_X1    g0703(.A1(new_n670_), .A2(new_n663_), .ZN(new_n753_));
  OAI21_X1   g0704(.A1(new_n752_), .A2(new_n753_), .B(new_n673_), .ZN(new_n754_));
  NAND2_X1   g0705(.A1(new_n754_), .A2(new_n365_), .ZN(new_n755_));
  AND2_X2    g0706(.A1(new_n659_), .A2(new_n755_), .Z(new_n756_));
  INV_X1     g0707(.I(new_n594_), .ZN(new_n757_));
  NOR2_X1    g0708(.A1(new_n538_), .A2(new_n592_), .ZN(new_n758_));
  INV_X1     g0709(.I(new_n758_), .ZN(new_n759_));
  NAND2_X1   g0710(.A1(new_n759_), .A2(new_n593_), .ZN(new_n760_));
  INV_X1     g0711(.I(new_n760_), .ZN(new_n761_));
  NOR2_X1    g0712(.A1(new_n761_), .A2(new_n757_), .ZN(new_n762_));
  INV_X1     g0713(.I(new_n762_), .ZN(new_n763_));
  NAND2_X1   g0714(.A1(new_n763_), .A2(new_n620_), .ZN(new_n764_));
  NOR2_X1    g0715(.A1(new_n758_), .A2(new_n423_), .ZN(new_n765_));
  NOR2_X1    g0716(.A1(new_n761_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1     g0717(.I(new_n766_), .ZN(new_n767_));
  NAND2_X1   g0718(.A1(new_n767_), .A2(new_n462_), .ZN(new_n768_));
  NAND3_X1   g0719(.A1(new_n759_), .A2(new_n423_), .A3(new_n593_), .ZN(new_n769_));
  NAND2_X1   g0720(.A1(new_n769_), .A2(new_n465_), .ZN(new_n770_));
  NAND3_X1   g0721(.A1(new_n759_), .A2(new_n422_), .A3(new_n593_), .ZN(new_n771_));
  NAND2_X1   g0722(.A1(new_n771_), .A2(new_n598_), .ZN(new_n772_));
  AOI22_X1   g0723(.A1(new_n768_), .A2(new_n764_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1     g0724(.I(new_n773_), .ZN(new_n774_));
  NOR2_X1    g0725(.A1(new_n624_), .A2(new_n616_), .ZN(new_n775_));
  NOR2_X1    g0726(.A1(new_n775_), .A2(new_n474_), .ZN(new_n776_));
  AOI21_X1   g0727(.A1(new_n614_), .A2(new_n600_), .B(new_n473_), .ZN(new_n777_));
  NOR2_X1    g0728(.A1(new_n614_), .A2(new_n616_), .ZN(new_n778_));
  NOR2_X1    g0729(.A1(new_n778_), .A2(new_n478_), .ZN(new_n779_));
  AOI21_X1   g0730(.A1(new_n627_), .A2(new_n469_), .B(new_n477_), .ZN(new_n780_));
  OAI22_X1   g0731(.A1(new_n776_), .A2(new_n777_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1   g0732(.A1(new_n774_), .A2(new_n781_), .ZN(new_n782_));
  NOR2_X1    g0733(.A1(new_n469_), .A2(new_n664_), .ZN(new_n783_));
  INV_X1     g0734(.I(new_n783_), .ZN(new_n784_));
  INV_X1     g0735(.I(new_n705_), .ZN(new_n785_));
  NOR2_X1    g0736(.A1(new_n290_), .A2(new_n222_), .ZN(new_n786_));
  NAND2_X1   g0737(.A1(new_n786_), .A2(new_n227_), .ZN(new_n787_));
  NAND3_X1   g0738(.A1(new_n235_), .A2(new_n145_), .A3(new_n154_), .ZN(new_n788_));
  NAND3_X1   g0739(.A1(new_n787_), .A2(new_n788_), .A3(new_n491_), .ZN(new_n789_));
  NOR3_X1    g0740(.A1(new_n789_), .A2(new_n337_), .A3(new_n711_), .ZN(new_n790_));
  NAND2_X1   g0741(.A1(new_n786_), .A2(new_n482_), .ZN(new_n791_));
  NAND3_X1   g0742(.A1(new_n394_), .A2(new_n145_), .A3(new_n154_), .ZN(new_n792_));
  NAND4_X1   g0743(.A1(new_n791_), .A2(new_n677_), .A3(new_n792_), .A4(new_n717_), .ZN(new_n793_));
  NOR4_X1    g0744(.A1(new_n793_), .A2(new_n139_), .A3(new_n388_), .A4(new_n715_), .ZN(new_n794_));
  NAND4_X1   g0745(.A1(new_n794_), .A2(new_n707_), .A3(new_n790_), .A4(new_n708_), .ZN(new_n795_));
  NAND4_X1   g0746(.A1(new_n732_), .A2(new_n728_), .A3(new_n189_), .A4(new_n724_), .ZN(new_n796_));
  NAND3_X1   g0747(.A1(new_n392_), .A2(new_n115_), .A3(new_n145_), .ZN(new_n797_));
  NAND4_X1   g0748(.A1(new_n451_), .A2(new_n740_), .A3(new_n797_), .A4(new_n739_), .ZN(new_n798_));
  NOR3_X1    g0749(.A1(new_n798_), .A2(new_n177_), .A3(new_n373_), .ZN(new_n799_));
  NAND3_X1   g0750(.A1(new_n229_), .A2(new_n239_), .A3(new_n125_), .ZN(new_n800_));
  NAND4_X1   g0751(.A1(new_n800_), .A2(new_n433_), .A3(new_n439_), .A4(new_n301_), .ZN(new_n801_));
  NOR3_X1    g0752(.A1(new_n801_), .A2(new_n207_), .A3(new_n382_), .ZN(new_n802_));
  NAND4_X1   g0753(.A1(new_n802_), .A2(new_n799_), .A3(new_n379_), .A4(new_n737_), .ZN(new_n803_));
  NOR3_X1    g0754(.A1(new_n795_), .A2(new_n796_), .A3(new_n803_), .ZN(new_n804_));
  NOR3_X1    g0755(.A1(new_n592_), .A2(new_n598_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1   g0756(.A1(new_n592_), .A2(new_n804_), .B(new_n805_), .ZN(new_n806_));
  NOR2_X1    g0757(.A1(new_n749_), .A2(new_n598_), .ZN(new_n807_));
  OAI22_X1   g0758(.A1(new_n806_), .A2(new_n785_), .B1(new_n751_), .B2(new_n807_), .ZN(new_n808_));
  NOR2_X1    g0759(.A1(new_n808_), .A2(new_n784_), .ZN(new_n809_));
  NOR2_X1    g0760(.A1(new_n762_), .A2(new_n477_), .ZN(new_n810_));
  NOR2_X1    g0761(.A1(new_n766_), .A2(new_n478_), .ZN(new_n811_));
  INV_X1     g0762(.I(new_n769_), .ZN(new_n812_));
  NOR2_X1    g0763(.A1(new_n812_), .A2(new_n620_), .ZN(new_n813_));
  INV_X1     g0764(.I(new_n771_), .ZN(new_n814_));
  NOR2_X1    g0765(.A1(new_n814_), .A2(new_n462_), .ZN(new_n815_));
  OAI22_X1   g0766(.A1(new_n810_), .A2(new_n811_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1   g0767(.A1(new_n808_), .A2(new_n784_), .ZN(new_n817_));
  AOI21_X1   g0768(.A1(new_n816_), .A2(new_n817_), .B(new_n809_), .ZN(new_n818_));
  NOR2_X1    g0769(.A1(new_n774_), .A2(new_n781_), .ZN(new_n819_));
  OAI21_X1   g0770(.A1(new_n818_), .A2(new_n819_), .B(new_n782_), .ZN(new_n820_));
  INV_X1     g0771(.I(new_n820_), .ZN(new_n821_));
  NOR2_X1    g0772(.A1(new_n659_), .A2(new_n755_), .ZN(new_n822_));
  NOR2_X1    g0773(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NOR2_X1    g0774(.A1(new_n823_), .A2(new_n756_), .ZN(new_n824_));
  XNOR2_X1   g0775(.A1(new_n630_), .A2(new_n633_), .ZN(new_n825_));
  XOR2_X1    g0776(.A1(new_n825_), .A2(new_n650_), .Z(new_n826_));
  XOR2_X1    g0777(.A1(new_n824_), .A2(new_n826_), .Z(new_n827_));
  INV_X1     g0778(.I(new_n782_), .ZN(new_n828_));
  NOR2_X1    g0779(.A1(new_n828_), .A2(new_n819_), .ZN(new_n829_));
  XOR2_X1    g0780(.A1(new_n829_), .A2(new_n818_), .Z(new_n830_));
  XNOR2_X1   g0781(.A1(new_n670_), .A2(new_n663_), .ZN(new_n831_));
  NOR2_X1    g0782(.A1(new_n469_), .A2(new_n831_), .ZN(new_n832_));
  XOR2_X1    g0783(.A1(new_n832_), .A2(new_n751_), .Z(new_n833_));
  NOR2_X1    g0784(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1   g0785(.A1(new_n618_), .A2(new_n670_), .ZN(new_n835_));
  NAND2_X1   g0786(.A1(new_n621_), .A2(new_n671_), .ZN(new_n836_));
  NAND2_X1   g0787(.A1(new_n625_), .A2(new_n473_), .ZN(new_n837_));
  NAND2_X1   g0788(.A1(new_n628_), .A2(new_n474_), .ZN(new_n838_));
  AOI22_X1   g0789(.A1(new_n835_), .A2(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1     g0790(.I(\a[7] ), .ZN(new_n840_));
  NAND2_X1   g0791(.A1(new_n660_), .A2(new_n57_), .ZN(new_n841_));
  XOR2_X1    g0792(.A1(new_n841_), .A2(new_n840_), .Z(new_n842_));
  INV_X1     g0793(.I(new_n842_), .ZN(new_n843_));
  AOI21_X1   g0794(.A1(new_n60_), .A2(new_n840_), .B(\a[22] ), .ZN(new_n844_));
  XOR2_X1    g0795(.A1(new_n844_), .A2(\a[8] ), .Z(new_n845_));
  INV_X1     g0796(.I(new_n845_), .ZN(new_n846_));
  NOR2_X1    g0797(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1     g0798(.I(new_n847_), .ZN(new_n848_));
  INV_X1     g0799(.I(new_n179_), .ZN(new_n849_));
  NOR3_X1    g0800(.A1(new_n139_), .A2(new_n330_), .A3(new_n722_), .ZN(new_n850_));
  NOR2_X1    g0801(.A1(new_n261_), .A2(new_n197_), .ZN(new_n851_));
  NOR3_X1    g0802(.A1(new_n246_), .A2(new_n263_), .A3(new_n402_), .ZN(new_n852_));
  NAND4_X1   g0803(.A1(new_n851_), .A2(new_n852_), .A3(new_n850_), .A4(new_n849_), .ZN(new_n853_));
  INV_X1     g0804(.I(new_n398_), .ZN(new_n854_));
  NOR3_X1    g0805(.A1(new_n854_), .A2(new_n545_), .A3(new_n191_), .ZN(new_n855_));
  NOR2_X1    g0806(.A1(new_n232_), .A2(new_n91_), .ZN(new_n856_));
  NOR2_X1    g0807(.A1(new_n201_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1    g0808(.A1(new_n437_), .A2(new_n245_), .ZN(new_n858_));
  NAND4_X1   g0809(.A1(new_n855_), .A2(new_n455_), .A3(new_n858_), .A4(new_n857_), .ZN(new_n859_));
  NAND4_X1   g0810(.A1(new_n743_), .A2(new_n255_), .A3(new_n583_), .A4(new_n800_), .ZN(new_n860_));
  INV_X1     g0811(.I(new_n860_), .ZN(new_n861_));
  NOR4_X1    g0812(.A1(new_n159_), .A2(new_n205_), .A3(new_n495_), .A4(new_n361_), .ZN(new_n862_));
  NAND4_X1   g0813(.A1(new_n370_), .A2(new_n408_), .A3(new_n369_), .A4(new_n412_), .ZN(new_n863_));
  NAND2_X1   g0814(.A1(new_n407_), .A2(new_n482_), .ZN(new_n864_));
  NAND3_X1   g0815(.A1(new_n368_), .A2(new_n864_), .A3(new_n530_), .ZN(new_n865_));
  NOR2_X1    g0816(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1   g0817(.A1(new_n674_), .A2(new_n293_), .A3(new_n316_), .ZN(new_n867_));
  AOI21_X1   g0818(.A1(new_n122_), .A2(new_n233_), .B(new_n126_), .ZN(new_n868_));
  OAI21_X1   g0819(.A1(new_n167_), .A2(new_n232_), .B(new_n792_), .ZN(new_n869_));
  NAND3_X1   g0820(.A1(new_n235_), .A2(new_n108_), .A3(new_n145_), .ZN(new_n870_));
  NAND3_X1   g0821(.A1(new_n315_), .A2(new_n145_), .A3(new_n154_), .ZN(new_n871_));
  NAND4_X1   g0822(.A1(new_n787_), .A2(new_n870_), .A3(new_n871_), .A4(new_n528_), .ZN(new_n872_));
  NOR4_X1    g0823(.A1(new_n872_), .A2(new_n867_), .A3(new_n868_), .A4(new_n869_), .ZN(new_n873_));
  NAND4_X1   g0824(.A1(new_n873_), .A2(new_n861_), .A3(new_n862_), .A4(new_n866_), .ZN(new_n874_));
  NAND2_X1   g0825(.A1(new_n394_), .A2(new_n223_), .ZN(new_n875_));
  NAND2_X1   g0826(.A1(new_n744_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1   g0827(.A1(new_n315_), .A2(new_n99_), .A3(new_n108_), .ZN(new_n877_));
  NAND2_X1   g0828(.A1(new_n565_), .A2(new_n877_), .ZN(new_n878_));
  NOR4_X1    g0829(.A1(new_n876_), .A2(new_n878_), .A3(new_n202_), .A4(new_n515_), .ZN(new_n879_));
  NOR4_X1    g0830(.A1(new_n210_), .A2(new_n317_), .A3(new_n254_), .A4(new_n497_), .ZN(new_n880_));
  NAND2_X1   g0831(.A1(new_n395_), .A2(new_n431_), .ZN(new_n881_));
  NOR4_X1    g0832(.A1(new_n387_), .A2(new_n881_), .A3(new_n168_), .A4(new_n378_), .ZN(new_n882_));
  NAND4_X1   g0833(.A1(new_n882_), .A2(new_n879_), .A3(new_n514_), .A4(new_n880_), .ZN(new_n883_));
  NOR4_X1    g0834(.A1(new_n874_), .A2(new_n853_), .A3(new_n859_), .A4(new_n883_), .ZN(new_n884_));
  NOR3_X1    g0835(.A1(new_n251_), .A2(new_n73_), .A3(new_n182_), .ZN(new_n885_));
  NOR2_X1    g0836(.A1(new_n290_), .A2(new_n238_), .ZN(new_n886_));
  AOI22_X1   g0837(.A1(new_n885_), .A2(new_n223_), .B1(new_n886_), .B2(new_n235_), .ZN(new_n887_));
  NOR4_X1    g0838(.A1(new_n691_), .A2(new_n267_), .A3(new_n693_), .A4(new_n580_), .ZN(new_n888_));
  NAND3_X1   g0839(.A1(new_n227_), .A2(new_n115_), .A3(new_n121_), .ZN(new_n889_));
  NAND2_X1   g0840(.A1(new_n235_), .A2(new_n366_), .ZN(new_n890_));
  NAND4_X1   g0841(.A1(new_n889_), .A2(new_n236_), .A3(new_n890_), .A4(new_n224_), .ZN(new_n891_));
  NAND3_X1   g0842(.A1(new_n227_), .A2(new_n115_), .A3(new_n145_), .ZN(new_n892_));
  NAND3_X1   g0843(.A1(new_n892_), .A2(new_n275_), .A3(new_n685_), .ZN(new_n893_));
  NOR2_X1    g0844(.A1(new_n891_), .A2(new_n893_), .ZN(new_n894_));
  NAND4_X1   g0845(.A1(new_n894_), .A2(new_n445_), .A3(new_n887_), .A4(new_n888_), .ZN(new_n895_));
  NOR3_X1    g0846(.A1(new_n524_), .A2(new_n357_), .A3(new_n856_), .ZN(new_n896_));
  NOR3_X1    g0847(.A1(new_n294_), .A2(new_n382_), .A3(new_n296_), .ZN(new_n897_));
  NAND3_X1   g0848(.A1(new_n897_), .A2(new_n543_), .A3(new_n896_), .ZN(new_n898_));
  NAND3_X1   g0849(.A1(new_n235_), .A2(new_n115_), .A3(new_n145_), .ZN(new_n899_));
  NAND3_X1   g0850(.A1(new_n482_), .A2(new_n108_), .A3(new_n145_), .ZN(new_n900_));
  NAND4_X1   g0851(.A1(new_n899_), .A2(new_n301_), .A3(new_n900_), .A4(new_n739_), .ZN(new_n901_));
  NAND3_X1   g0852(.A1(new_n482_), .A2(new_n99_), .A3(new_n108_), .ZN(new_n902_));
  NAND2_X1   g0853(.A1(new_n565_), .A2(new_n902_), .ZN(new_n903_));
  NOR3_X1    g0854(.A1(new_n901_), .A2(new_n175_), .A3(new_n903_), .ZN(new_n904_));
  NAND2_X1   g0855(.A1(new_n684_), .A2(new_n740_), .ZN(new_n905_));
  OAI22_X1   g0856(.A1(new_n204_), .A2(new_n195_), .B1(new_n336_), .B2(new_n320_), .ZN(new_n906_));
  NOR4_X1    g0857(.A1(new_n905_), .A2(new_n256_), .A3(new_n569_), .A4(new_n906_), .ZN(new_n907_));
  NAND3_X1   g0858(.A1(new_n315_), .A2(new_n121_), .A3(new_n154_), .ZN(new_n908_));
  NAND3_X1   g0859(.A1(new_n235_), .A2(new_n108_), .A3(new_n121_), .ZN(new_n909_));
  NAND4_X1   g0860(.A1(new_n909_), .A2(new_n329_), .A3(new_n151_), .A4(new_n908_), .ZN(new_n910_));
  NAND4_X1   g0861(.A1(new_n302_), .A2(new_n73_), .A3(new_n121_), .A4(new_n137_), .ZN(new_n911_));
  NAND2_X1   g0862(.A1(new_n490_), .A2(new_n216_), .ZN(new_n912_));
  NAND3_X1   g0863(.A1(new_n911_), .A2(new_n912_), .A3(new_n578_), .ZN(new_n913_));
  NAND2_X1   g0864(.A1(new_n676_), .A2(new_n429_), .ZN(new_n914_));
  NOR3_X1    g0865(.A1(new_n910_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  OAI22_X1   g0866(.A1(new_n192_), .A2(new_n158_), .B1(new_n109_), .B2(new_n167_), .ZN(new_n916_));
  NOR4_X1    g0867(.A1(new_n916_), .A2(new_n245_), .A3(new_n718_), .A4(new_n338_), .ZN(new_n917_));
  NAND4_X1   g0868(.A1(new_n915_), .A2(new_n904_), .A3(new_n907_), .A4(new_n917_), .ZN(new_n918_));
  NOR3_X1    g0869(.A1(new_n194_), .A2(new_n252_), .A3(new_n251_), .ZN(new_n919_));
  NOR4_X1    g0870(.A1(new_n723_), .A2(new_n271_), .A3(new_n919_), .A4(new_n548_), .ZN(new_n920_));
  NAND2_X1   g0871(.A1(new_n366_), .A2(new_n315_), .ZN(new_n921_));
  NAND4_X1   g0872(.A1(new_n372_), .A2(new_n551_), .A3(new_n921_), .A4(new_n556_), .ZN(new_n922_));
  NOR2_X1    g0873(.A1(new_n922_), .A2(new_n352_), .ZN(new_n923_));
  OAI22_X1   g0874(.A1(new_n178_), .A2(new_n167_), .B1(new_n155_), .B2(new_n126_), .ZN(new_n924_));
  OAI22_X1   g0875(.A1(new_n204_), .A2(new_n91_), .B1(new_n155_), .B2(new_n195_), .ZN(new_n925_));
  NAND2_X1   g0876(.A1(new_n563_), .A2(new_n677_), .ZN(new_n926_));
  NOR4_X1    g0877(.A1(new_n926_), .A2(new_n924_), .A3(new_n925_), .A4(new_n254_), .ZN(new_n927_));
  NAND4_X1   g0878(.A1(new_n923_), .A2(new_n588_), .A3(new_n927_), .A4(new_n920_), .ZN(new_n928_));
  NOR4_X1    g0879(.A1(new_n918_), .A2(new_n928_), .A3(new_n895_), .A4(new_n898_), .ZN(new_n929_));
  OAI21_X1   g0880(.A1(new_n884_), .A2(new_n929_), .B(new_n749_), .ZN(new_n930_));
  OAI21_X1   g0881(.A1(new_n842_), .A2(new_n845_), .B(new_n930_), .ZN(new_n931_));
  AOI21_X1   g0882(.A1(new_n931_), .A2(new_n848_), .B(new_n469_), .ZN(new_n932_));
  NOR2_X1    g0883(.A1(new_n839_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1   g0884(.A1(new_n618_), .A2(new_n663_), .ZN(new_n934_));
  NAND2_X1   g0885(.A1(new_n621_), .A2(new_n664_), .ZN(new_n935_));
  NAND2_X1   g0886(.A1(new_n625_), .A2(new_n670_), .ZN(new_n936_));
  NAND2_X1   g0887(.A1(new_n628_), .A2(new_n671_), .ZN(new_n937_));
  AOI22_X1   g0888(.A1(new_n934_), .A2(new_n935_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  INV_X1     g0889(.I(new_n750_), .ZN(new_n939_));
  NOR2_X1    g0890(.A1(new_n705_), .A2(new_n749_), .ZN(new_n940_));
  AOI21_X1   g0891(.A1(new_n636_), .A2(new_n940_), .B(new_n939_), .ZN(new_n941_));
  NAND2_X1   g0892(.A1(new_n941_), .A2(new_n620_), .ZN(new_n942_));
  INV_X1     g0893(.I(new_n940_), .ZN(new_n943_));
  OAI21_X1   g0894(.A1(new_n636_), .A2(new_n750_), .B(new_n943_), .ZN(new_n944_));
  INV_X1     g0895(.I(new_n944_), .ZN(new_n945_));
  NAND2_X1   g0896(.A1(new_n945_), .A2(new_n462_), .ZN(new_n946_));
  NAND3_X1   g0897(.A1(new_n943_), .A2(new_n592_), .A3(new_n750_), .ZN(new_n947_));
  NAND2_X1   g0898(.A1(new_n947_), .A2(new_n465_), .ZN(new_n948_));
  NAND3_X1   g0899(.A1(new_n943_), .A2(new_n636_), .A3(new_n750_), .ZN(new_n949_));
  NAND2_X1   g0900(.A1(new_n949_), .A2(new_n598_), .ZN(new_n950_));
  AOI22_X1   g0901(.A1(new_n942_), .A2(new_n946_), .B1(new_n948_), .B2(new_n950_), .ZN(new_n951_));
  NOR2_X1    g0902(.A1(new_n938_), .A2(new_n951_), .ZN(new_n952_));
  NAND2_X1   g0903(.A1(new_n763_), .A2(new_n474_), .ZN(new_n953_));
  NAND2_X1   g0904(.A1(new_n767_), .A2(new_n473_), .ZN(new_n954_));
  NOR2_X1    g0905(.A1(new_n812_), .A2(new_n478_), .ZN(new_n955_));
  AOI21_X1   g0906(.A1(new_n478_), .A2(new_n771_), .B(new_n955_), .ZN(new_n956_));
  AOI21_X1   g0907(.A1(new_n953_), .A2(new_n954_), .B(new_n956_), .ZN(new_n957_));
  AOI21_X1   g0908(.A1(new_n938_), .A2(new_n951_), .B(new_n957_), .ZN(new_n958_));
  NOR2_X1    g0909(.A1(new_n958_), .A2(new_n952_), .ZN(new_n959_));
  INV_X1     g0910(.I(new_n959_), .ZN(new_n960_));
  NAND2_X1   g0911(.A1(new_n839_), .A2(new_n932_), .ZN(new_n961_));
  AOI21_X1   g0912(.A1(new_n960_), .A2(new_n961_), .B(new_n933_), .ZN(new_n962_));
  AOI21_X1   g0913(.A1(new_n830_), .A2(new_n833_), .B(new_n962_), .ZN(new_n963_));
  NOR2_X1    g0914(.A1(new_n963_), .A2(new_n834_), .ZN(new_n964_));
  INV_X1     g0915(.I(new_n964_), .ZN(new_n965_));
  NOR2_X1    g0916(.A1(new_n756_), .A2(new_n822_), .ZN(new_n966_));
  XOR2_X1    g0917(.A1(new_n966_), .A2(new_n821_), .Z(new_n967_));
  INV_X1     g0918(.I(new_n967_), .ZN(new_n968_));
  NOR2_X1    g0919(.A1(new_n965_), .A2(new_n968_), .ZN(new_n969_));
  INV_X1     g0920(.I(new_n969_), .ZN(new_n970_));
  NOR2_X1    g0921(.A1(new_n469_), .A2(new_n843_), .ZN(new_n971_));
  INV_X1     g0922(.I(new_n853_), .ZN(new_n972_));
  INV_X1     g0923(.I(new_n859_), .ZN(new_n973_));
  INV_X1     g0924(.I(new_n862_), .ZN(new_n974_));
  NOR3_X1    g0925(.A1(new_n253_), .A2(new_n244_), .A3(new_n272_), .ZN(new_n975_));
  NAND2_X1   g0926(.A1(new_n920_), .A2(new_n975_), .ZN(new_n976_));
  OAI22_X1   g0927(.A1(new_n204_), .A2(new_n167_), .B1(new_n91_), .B2(new_n194_), .ZN(new_n977_));
  NOR3_X1    g0928(.A1(new_n977_), .A2(new_n294_), .A3(new_n868_), .ZN(new_n978_));
  NOR2_X1    g0929(.A1(new_n327_), .A2(new_n687_), .ZN(new_n979_));
  NOR4_X1    g0930(.A1(new_n267_), .A2(new_n265_), .A3(new_n339_), .A4(new_n376_), .ZN(new_n980_));
  NAND3_X1   g0931(.A1(new_n978_), .A2(new_n980_), .A3(new_n979_), .ZN(new_n981_));
  NOR4_X1    g0932(.A1(new_n981_), .A2(new_n860_), .A3(new_n976_), .A4(new_n974_), .ZN(new_n982_));
  AOI21_X1   g0933(.A1(new_n115_), .A2(new_n121_), .B(new_n407_), .ZN(new_n983_));
  NOR2_X1    g0934(.A1(new_n983_), .A2(new_n91_), .ZN(new_n984_));
  NOR2_X1    g0935(.A1(new_n295_), .A2(new_n238_), .ZN(new_n985_));
  INV_X1     g0936(.I(new_n178_), .ZN(new_n986_));
  AOI22_X1   g0937(.A1(new_n986_), .A2(new_n539_), .B1(new_n985_), .B2(new_n315_), .ZN(new_n987_));
  NAND4_X1   g0938(.A1(new_n987_), .A2(new_n383_), .A3(new_n512_), .A4(new_n303_), .ZN(new_n988_));
  NAND3_X1   g0939(.A1(new_n227_), .A2(new_n99_), .A3(new_n154_), .ZN(new_n989_));
  NOR2_X1    g0940(.A1(new_n286_), .A2(new_n280_), .ZN(new_n990_));
  OAI21_X1   g0941(.A1(new_n990_), .A2(new_n886_), .B(new_n482_), .ZN(new_n991_));
  NAND4_X1   g0942(.A1(new_n991_), .A2(new_n372_), .A3(new_n989_), .A4(new_n433_), .ZN(new_n992_));
  INV_X1     g0943(.I(new_n168_), .ZN(new_n993_));
  NAND2_X1   g0944(.A1(new_n513_), .A2(new_n235_), .ZN(new_n994_));
  NOR2_X1    g0945(.A1(new_n494_), .A2(new_n296_), .ZN(new_n995_));
  NAND4_X1   g0946(.A1(new_n995_), .A2(new_n993_), .A3(new_n994_), .A4(new_n386_), .ZN(new_n996_));
  NOR4_X1    g0947(.A1(new_n988_), .A2(new_n984_), .A3(new_n996_), .A4(new_n992_), .ZN(new_n997_));
  NAND4_X1   g0948(.A1(new_n982_), .A2(new_n972_), .A3(new_n997_), .A4(new_n973_), .ZN(new_n998_));
  OAI22_X1   g0949(.A1(new_n192_), .A2(new_n359_), .B1(new_n155_), .B2(new_n266_), .ZN(new_n999_));
  NAND2_X1   g0950(.A1(new_n885_), .A2(new_n786_), .ZN(new_n1000_));
  NAND4_X1   g0951(.A1(new_n581_), .A2(new_n1000_), .A3(new_n870_), .A4(new_n491_), .ZN(new_n1001_));
  NOR4_X1    g0952(.A1(new_n188_), .A2(new_n330_), .A3(new_n557_), .A4(new_n337_), .ZN(new_n1002_));
  NOR3_X1    g0953(.A1(new_n276_), .A2(new_n201_), .A3(new_n736_), .ZN(new_n1003_));
  NAND2_X1   g0954(.A1(new_n1003_), .A2(new_n1002_), .ZN(new_n1004_));
  NOR4_X1    g0955(.A1(new_n1004_), .A2(new_n446_), .A3(new_n999_), .A4(new_n1001_), .ZN(new_n1005_));
  INV_X1     g0956(.I(new_n898_), .ZN(new_n1006_));
  NOR4_X1    g0957(.A1(new_n426_), .A2(new_n341_), .A3(new_n495_), .A4(new_n443_), .ZN(new_n1007_));
  AOI22_X1   g0958(.A1(new_n986_), .A2(new_n539_), .B1(new_n985_), .B2(new_n482_), .ZN(new_n1008_));
  NAND3_X1   g0959(.A1(new_n1007_), .A2(new_n1008_), .A3(new_n176_), .ZN(new_n1009_));
  NOR2_X1    g0960(.A1(new_n263_), .A2(new_n729_), .ZN(new_n1010_));
  OAI21_X1   g0961(.A1(new_n985_), .A2(new_n407_), .B(new_n539_), .ZN(new_n1011_));
  NOR2_X1    g0962(.A1(new_n402_), .A2(new_n687_), .ZN(new_n1012_));
  NAND4_X1   g0963(.A1(new_n1010_), .A2(new_n1011_), .A3(new_n1012_), .A4(new_n255_), .ZN(new_n1013_));
  NOR3_X1    g0964(.A1(new_n262_), .A2(new_n492_), .A3(new_n544_), .ZN(new_n1014_));
  NOR2_X1    g0965(.A1(new_n404_), .A2(new_n243_), .ZN(new_n1015_));
  NOR3_X1    g0966(.A1(new_n321_), .A2(new_n361_), .A3(new_n1015_), .ZN(new_n1016_));
  NOR2_X1    g0967(.A1(new_n246_), .A2(new_n196_), .ZN(new_n1017_));
  NAND4_X1   g0968(.A1(new_n1014_), .A2(new_n1016_), .A3(new_n1017_), .A4(new_n909_), .ZN(new_n1018_));
  INV_X1     g0969(.I(new_n158_), .ZN(new_n1019_));
  AOI22_X1   g0970(.A1(new_n1019_), .A2(new_n885_), .B1(new_n985_), .B2(new_n227_), .ZN(new_n1020_));
  NAND4_X1   g0971(.A1(new_n1020_), .A2(new_n675_), .A3(new_n791_), .A4(new_n717_), .ZN(new_n1021_));
  NOR4_X1    g0972(.A1(new_n1018_), .A2(new_n1009_), .A3(new_n1021_), .A4(new_n1013_), .ZN(new_n1022_));
  INV_X1     g0973(.I(new_n452_), .ZN(new_n1023_));
  NAND2_X1   g0974(.A1(new_n409_), .A2(new_n539_), .ZN(new_n1024_));
  NAND3_X1   g0975(.A1(new_n1023_), .A2(new_n1024_), .A3(new_n260_), .ZN(new_n1025_));
  NOR3_X1    g0976(.A1(new_n503_), .A2(new_n722_), .A3(new_n698_), .ZN(new_n1026_));
  NOR2_X1    g0977(.A1(new_n269_), .A2(new_n425_), .ZN(new_n1027_));
  NAND4_X1   g0978(.A1(new_n1026_), .A2(new_n372_), .A3(new_n551_), .A4(new_n1027_), .ZN(new_n1028_));
  NOR3_X1    g0979(.A1(new_n254_), .A2(new_n345_), .A3(new_n291_), .ZN(new_n1029_));
  NAND3_X1   g0980(.A1(new_n1029_), .A2(new_n180_), .A3(new_n498_), .ZN(new_n1030_));
  NOR4_X1    g0981(.A1(new_n1028_), .A2(new_n1030_), .A3(new_n1025_), .A4(new_n863_), .ZN(new_n1031_));
  NAND4_X1   g0982(.A1(new_n1022_), .A2(new_n1005_), .A3(new_n1031_), .A4(new_n1006_), .ZN(new_n1032_));
  NOR2_X1    g0983(.A1(new_n1032_), .A2(new_n804_), .ZN(new_n1033_));
  NAND2_X1   g0984(.A1(new_n1032_), .A2(new_n804_), .ZN(new_n1034_));
  NOR2_X1    g0985(.A1(new_n1034_), .A2(new_n598_), .ZN(new_n1035_));
  OAI21_X1   g0986(.A1(new_n1035_), .A2(new_n1033_), .B(new_n998_), .ZN(new_n1036_));
  INV_X1     g0987(.I(new_n1036_), .ZN(new_n1037_));
  AOI21_X1   g0988(.A1(new_n465_), .A2(new_n929_), .B(new_n930_), .ZN(new_n1038_));
  NOR2_X1    g0989(.A1(new_n1037_), .A2(new_n1038_), .ZN(new_n1039_));
  INV_X1     g0990(.I(new_n971_), .ZN(new_n1040_));
  INV_X1     g0991(.I(new_n1039_), .ZN(new_n1041_));
  NOR2_X1    g0992(.A1(new_n944_), .A2(new_n478_), .ZN(new_n1042_));
  AOI21_X1   g0993(.A1(new_n478_), .A2(new_n941_), .B(new_n1042_), .ZN(new_n1043_));
  NOR3_X1    g0994(.A1(new_n939_), .A2(new_n592_), .A3(new_n940_), .ZN(new_n1044_));
  NOR2_X1    g0995(.A1(new_n1044_), .A2(new_n462_), .ZN(new_n1045_));
  AOI21_X1   g0996(.A1(new_n462_), .A2(new_n947_), .B(new_n1045_), .ZN(new_n1046_));
  NOR2_X1    g0997(.A1(new_n1043_), .A2(new_n1046_), .ZN(new_n1047_));
  AOI21_X1   g0998(.A1(new_n1040_), .A2(new_n1041_), .B(new_n1047_), .ZN(new_n1048_));
  AOI21_X1   g0999(.A1(new_n971_), .A2(new_n1039_), .B(new_n1048_), .ZN(new_n1049_));
  AOI21_X1   g1000(.A1(new_n998_), .A2(new_n1032_), .B(new_n804_), .ZN(new_n1050_));
  NOR2_X1    g1001(.A1(new_n843_), .A2(new_n845_), .ZN(new_n1051_));
  NOR2_X1    g1002(.A1(new_n846_), .A2(new_n842_), .ZN(new_n1052_));
  NOR2_X1    g1003(.A1(new_n1051_), .A2(new_n1052_), .ZN(new_n1053_));
  NOR2_X1    g1004(.A1(new_n1050_), .A2(new_n1053_), .ZN(new_n1054_));
  NOR2_X1    g1005(.A1(new_n842_), .A2(new_n845_), .ZN(new_n1055_));
  NOR2_X1    g1006(.A1(new_n847_), .A2(new_n1055_), .ZN(new_n1056_));
  NAND2_X1   g1007(.A1(new_n365_), .A2(new_n1056_), .ZN(new_n1057_));
  AOI22_X1   g1008(.A1(new_n1057_), .A2(new_n1050_), .B1(new_n1054_), .B2(new_n365_), .ZN(new_n1058_));
  NOR2_X1    g1009(.A1(new_n1049_), .A2(new_n1058_), .ZN(new_n1059_));
  NOR2_X1    g1010(.A1(new_n775_), .A2(new_n846_), .ZN(new_n1060_));
  AOI21_X1   g1011(.A1(new_n621_), .A2(new_n846_), .B(new_n1060_), .ZN(new_n1061_));
  NOR2_X1    g1012(.A1(new_n778_), .A2(new_n664_), .ZN(new_n1062_));
  AOI21_X1   g1013(.A1(new_n628_), .A2(new_n664_), .B(new_n1062_), .ZN(new_n1063_));
  NOR2_X1    g1014(.A1(new_n1061_), .A2(new_n1063_), .ZN(new_n1064_));
  NAND3_X1   g1015(.A1(new_n892_), .A2(new_n717_), .A3(new_n871_), .ZN(new_n1065_));
  NAND3_X1   g1016(.A1(new_n369_), .A2(new_n447_), .A3(new_n739_), .ZN(new_n1066_));
  NOR4_X1    g1017(.A1(new_n411_), .A2(new_n337_), .A3(new_n1065_), .A4(new_n1066_), .ZN(new_n1067_));
  NAND2_X1   g1018(.A1(new_n539_), .A2(new_n575_), .ZN(new_n1068_));
  NAND2_X1   g1019(.A1(new_n1068_), .A2(new_n491_), .ZN(new_n1069_));
  NAND4_X1   g1020(.A1(new_n989_), .A2(new_n684_), .A3(new_n797_), .A4(new_n432_), .ZN(new_n1070_));
  NAND4_X1   g1021(.A1(new_n160_), .A2(new_n994_), .A3(new_n889_), .A4(new_n350_), .ZN(new_n1071_));
  NOR4_X1    g1022(.A1(new_n1071_), .A2(new_n1069_), .A3(new_n175_), .A4(new_n1070_), .ZN(new_n1072_));
  OAI21_X1   g1023(.A1(new_n513_), .A2(new_n786_), .B(new_n482_), .ZN(new_n1073_));
  NAND4_X1   g1024(.A1(new_n1073_), .A2(new_n674_), .A3(new_n293_), .A4(new_n316_), .ZN(new_n1074_));
  NOR2_X1    g1025(.A1(new_n544_), .A2(new_n495_), .ZN(new_n1075_));
  NAND4_X1   g1026(.A1(new_n1075_), .A2(new_n849_), .A3(new_n292_), .A4(new_n540_), .ZN(new_n1076_));
  NOR3_X1    g1027(.A1(new_n580_), .A2(new_n327_), .A3(new_n402_), .ZN(new_n1077_));
  INV_X1     g1028(.I(new_n1077_), .ZN(new_n1078_));
  NAND3_X1   g1029(.A1(new_n227_), .A2(new_n108_), .A3(new_n162_), .ZN(new_n1079_));
  NOR3_X1    g1030(.A1(new_n515_), .A2(new_n443_), .A3(new_n299_), .ZN(new_n1080_));
  NOR2_X1    g1031(.A1(new_n332_), .A2(new_n497_), .ZN(new_n1081_));
  NAND4_X1   g1032(.A1(new_n1080_), .A2(new_n1081_), .A3(new_n1079_), .A4(new_n230_), .ZN(new_n1082_));
  NOR4_X1    g1033(.A1(new_n1082_), .A2(new_n1076_), .A3(new_n1074_), .A4(new_n1078_), .ZN(new_n1083_));
  NAND2_X1   g1034(.A1(new_n302_), .A2(new_n366_), .ZN(new_n1084_));
  NAND3_X1   g1035(.A1(new_n392_), .A2(new_n115_), .A3(new_n121_), .ZN(new_n1085_));
  NOR3_X1    g1036(.A1(new_n238_), .A2(new_n280_), .A3(new_n125_), .ZN(new_n1086_));
  OAI21_X1   g1037(.A1(new_n985_), .A2(new_n1086_), .B(new_n150_), .ZN(new_n1087_));
  NAND4_X1   g1038(.A1(new_n1087_), .A2(new_n1084_), .A3(new_n744_), .A4(new_n1085_), .ZN(new_n1088_));
  AOI21_X1   g1039(.A1(new_n409_), .A2(new_n482_), .B(new_n450_), .ZN(new_n1089_));
  NOR2_X1    g1040(.A1(new_n330_), .A2(new_n687_), .ZN(new_n1090_));
  NAND4_X1   g1041(.A1(new_n887_), .A2(new_n1090_), .A3(new_n1089_), .A4(new_n255_), .ZN(new_n1091_));
  NAND4_X1   g1042(.A1(new_n229_), .A2(new_n125_), .A3(new_n115_), .A4(new_n121_), .ZN(new_n1092_));
  AOI22_X1   g1043(.A1(new_n990_), .A2(new_n482_), .B1(new_n239_), .B2(new_n235_), .ZN(new_n1093_));
  NAND4_X1   g1044(.A1(new_n1093_), .A2(new_n514_), .A3(new_n368_), .A4(new_n1092_), .ZN(new_n1094_));
  NOR4_X1    g1045(.A1(new_n1091_), .A2(new_n577_), .A3(new_n1094_), .A4(new_n1088_), .ZN(new_n1095_));
  NAND4_X1   g1046(.A1(new_n1083_), .A2(new_n1095_), .A3(new_n1067_), .A4(new_n1072_), .ZN(new_n1096_));
  NAND2_X1   g1047(.A1(new_n122_), .A2(new_n270_), .ZN(new_n1097_));
  NAND2_X1   g1048(.A1(new_n178_), .A2(new_n359_), .ZN(new_n1098_));
  OAI21_X1   g1049(.A1(new_n1098_), .A2(new_n1097_), .B(new_n394_), .ZN(new_n1099_));
  NAND2_X1   g1050(.A1(new_n488_), .A2(new_n1099_), .ZN(new_n1100_));
  NOR4_X1    g1051(.A1(new_n1100_), .A2(new_n317_), .A3(new_n428_), .A4(new_n730_), .ZN(new_n1101_));
  NOR4_X1    g1052(.A1(new_n127_), .A2(new_n312_), .A3(new_n401_), .A4(new_n729_), .ZN(new_n1102_));
  INV_X1     g1053(.I(new_n1102_), .ZN(new_n1103_));
  NAND3_X1   g1054(.A1(new_n300_), .A2(new_n902_), .A3(new_n677_), .ZN(new_n1104_));
  NOR3_X1    g1055(.A1(new_n1103_), .A2(new_n396_), .A3(new_n1104_), .ZN(new_n1105_));
  INV_X1     g1056(.I(new_n424_), .ZN(new_n1106_));
  OAI22_X1   g1057(.A1(new_n135_), .A2(new_n359_), .B1(new_n266_), .B2(new_n194_), .ZN(new_n1107_));
  INV_X1     g1058(.I(new_n1107_), .ZN(new_n1108_));
  NAND3_X1   g1059(.A1(new_n579_), .A2(new_n850_), .A3(new_n1108_), .ZN(new_n1109_));
  INV_X1     g1060(.I(new_n185_), .ZN(new_n1110_));
  INV_X1     g1061(.I(new_n313_), .ZN(new_n1111_));
  NAND4_X1   g1062(.A1(new_n1110_), .A2(new_n1111_), .A3(new_n1000_), .A4(new_n565_), .ZN(new_n1112_));
  NOR3_X1    g1063(.A1(new_n254_), .A2(new_n736_), .A3(new_n515_), .ZN(new_n1113_));
  NAND3_X1   g1064(.A1(new_n154_), .A2(new_n73_), .A3(new_n162_), .ZN(new_n1114_));
  AOI21_X1   g1065(.A1(new_n1114_), .A2(new_n336_), .B(new_n243_), .ZN(new_n1115_));
  NOR3_X1    g1066(.A1(new_n1115_), .A2(new_n492_), .A3(new_n360_), .ZN(new_n1116_));
  NAND4_X1   g1067(.A1(new_n1116_), .A2(new_n1113_), .A3(new_n1020_), .A4(new_n255_), .ZN(new_n1117_));
  NOR4_X1    g1068(.A1(new_n1117_), .A2(new_n1109_), .A3(new_n1112_), .A4(new_n1106_), .ZN(new_n1118_));
  NOR3_X1    g1069(.A1(new_n382_), .A2(new_n444_), .A3(new_n324_), .ZN(new_n1119_));
  NOR2_X1    g1070(.A1(new_n126_), .A2(new_n138_), .ZN(new_n1120_));
  NOR4_X1    g1071(.A1(new_n191_), .A2(new_n495_), .A3(new_n361_), .A4(new_n1120_), .ZN(new_n1121_));
  NAND4_X1   g1072(.A1(new_n1121_), .A2(new_n311_), .A3(new_n1119_), .A4(new_n1087_), .ZN(new_n1122_));
  NOR2_X1    g1073(.A1(new_n509_), .A2(new_n253_), .ZN(new_n1123_));
  NAND3_X1   g1074(.A1(new_n108_), .A2(new_n145_), .A3(new_n73_), .ZN(new_n1124_));
  AOI21_X1   g1075(.A1(new_n1124_), .A2(new_n173_), .B(new_n243_), .ZN(new_n1125_));
  NOR2_X1    g1076(.A1(new_n1125_), .A2(new_n405_), .ZN(new_n1126_));
  NAND3_X1   g1077(.A1(new_n1126_), .A2(new_n701_), .A3(new_n1123_), .ZN(new_n1127_));
  NOR3_X1    g1078(.A1(new_n277_), .A2(new_n353_), .A3(new_n561_), .ZN(new_n1128_));
  NOR3_X1    g1079(.A1(new_n193_), .A2(new_n400_), .A3(new_n246_), .ZN(new_n1129_));
  NAND3_X1   g1080(.A1(new_n1129_), .A2(new_n1128_), .A3(new_n896_), .ZN(new_n1130_));
  NOR3_X1    g1081(.A1(new_n1122_), .A2(new_n1130_), .A3(new_n1127_), .ZN(new_n1131_));
  NAND4_X1   g1082(.A1(new_n1118_), .A2(new_n1131_), .A3(new_n1101_), .A4(new_n1105_), .ZN(new_n1132_));
  NAND2_X1   g1083(.A1(new_n1132_), .A2(new_n1096_), .ZN(new_n1133_));
  NAND2_X1   g1084(.A1(new_n1133_), .A2(new_n1032_), .ZN(new_n1134_));
  INV_X1     g1085(.I(new_n1067_), .ZN(new_n1135_));
  INV_X1     g1086(.I(new_n1070_), .ZN(new_n1136_));
  NOR4_X1    g1087(.A1(new_n188_), .A2(new_n503_), .A3(new_n378_), .A4(new_n159_), .ZN(new_n1137_));
  NAND4_X1   g1088(.A1(new_n1136_), .A2(new_n1137_), .A3(new_n694_), .A4(new_n176_), .ZN(new_n1138_));
  NAND2_X1   g1089(.A1(new_n900_), .A2(new_n151_), .ZN(new_n1139_));
  NOR4_X1    g1090(.A1(new_n564_), .A2(new_n1139_), .A3(new_n179_), .A4(new_n197_), .ZN(new_n1140_));
  NAND4_X1   g1091(.A1(new_n230_), .A2(new_n1079_), .A3(new_n583_), .A4(new_n433_), .ZN(new_n1141_));
  NOR2_X1    g1092(.A1(new_n1141_), .A2(new_n304_), .ZN(new_n1142_));
  NAND4_X1   g1093(.A1(new_n1142_), .A2(new_n978_), .A3(new_n1140_), .A4(new_n1077_), .ZN(new_n1143_));
  AOI21_X1   g1094(.A1(new_n91_), .A2(new_n126_), .B(new_n186_), .ZN(new_n1144_));
  NOR4_X1    g1095(.A1(new_n1144_), .A2(new_n210_), .A3(new_n250_), .A4(new_n573_), .ZN(new_n1145_));
  INV_X1     g1096(.I(new_n1086_), .ZN(new_n1146_));
  AOI21_X1   g1097(.A1(new_n1146_), .A2(new_n109_), .B(new_n172_), .ZN(new_n1147_));
  NAND3_X1   g1098(.A1(new_n744_), .A2(new_n1085_), .A3(new_n1084_), .ZN(new_n1148_));
  NOR2_X1    g1099(.A1(new_n1148_), .A2(new_n1147_), .ZN(new_n1149_));
  OAI21_X1   g1100(.A1(new_n126_), .A2(new_n163_), .B(new_n451_), .ZN(new_n1150_));
  OAI22_X1   g1101(.A1(new_n204_), .A2(new_n195_), .B1(new_n232_), .B2(new_n266_), .ZN(new_n1151_));
  NOR4_X1    g1102(.A1(new_n1150_), .A2(new_n999_), .A3(new_n256_), .A4(new_n1151_), .ZN(new_n1152_));
  NAND2_X1   g1103(.A1(new_n1092_), .A2(new_n368_), .ZN(new_n1153_));
  OAI22_X1   g1104(.A1(new_n126_), .A2(new_n249_), .B1(new_n266_), .B2(new_n194_), .ZN(new_n1154_));
  NOR3_X1    g1105(.A1(new_n1153_), .A2(new_n984_), .A3(new_n1154_), .ZN(new_n1155_));
  NAND4_X1   g1106(.A1(new_n1152_), .A2(new_n1155_), .A3(new_n1149_), .A4(new_n1145_), .ZN(new_n1156_));
  NOR4_X1    g1107(.A1(new_n1143_), .A2(new_n1156_), .A3(new_n1135_), .A4(new_n1138_), .ZN(new_n1157_));
  NOR2_X1    g1108(.A1(new_n59_), .A2(\a[4] ), .ZN(new_n1158_));
  INV_X1     g1109(.I(new_n1158_), .ZN(new_n1159_));
  OAI21_X1   g1110(.A1(new_n1159_), .A2(\a[5] ), .B(new_n57_), .ZN(new_n1160_));
  XNOR2_X1   g1111(.A1(new_n1160_), .A2(\a[6] ), .ZN(new_n1161_));
  INV_X1     g1112(.I(new_n1161_), .ZN(new_n1162_));
  NOR2_X1    g1113(.A1(new_n469_), .A2(new_n1162_), .ZN(new_n1163_));
  NOR2_X1    g1114(.A1(new_n1163_), .A2(new_n1157_), .ZN(new_n1164_));
  INV_X1     g1115(.I(new_n1164_), .ZN(new_n1165_));
  NAND2_X1   g1116(.A1(new_n1163_), .A2(new_n1157_), .ZN(new_n1166_));
  INV_X1     g1117(.I(new_n1166_), .ZN(new_n1167_));
  AOI21_X1   g1118(.A1(new_n1134_), .A2(new_n1165_), .B(new_n1167_), .ZN(new_n1168_));
  INV_X1     g1119(.I(new_n1168_), .ZN(new_n1169_));
  NOR2_X1    g1120(.A1(new_n1064_), .A2(new_n1169_), .ZN(new_n1170_));
  NAND2_X1   g1121(.A1(new_n763_), .A2(new_n671_), .ZN(new_n1171_));
  NAND2_X1   g1122(.A1(new_n767_), .A2(new_n670_), .ZN(new_n1172_));
  NOR2_X1    g1123(.A1(new_n812_), .A2(new_n474_), .ZN(new_n1173_));
  AOI21_X1   g1124(.A1(new_n474_), .A2(new_n771_), .B(new_n1173_), .ZN(new_n1174_));
  AOI21_X1   g1125(.A1(new_n1171_), .A2(new_n1172_), .B(new_n1174_), .ZN(new_n1175_));
  NOR3_X1    g1126(.A1(new_n1061_), .A2(new_n1063_), .A3(new_n1168_), .ZN(new_n1176_));
  NOR2_X1    g1127(.A1(new_n1176_), .A2(new_n1175_), .ZN(new_n1177_));
  NOR2_X1    g1128(.A1(new_n1177_), .A2(new_n1170_), .ZN(new_n1178_));
  AOI21_X1   g1129(.A1(new_n1049_), .A2(new_n1058_), .B(new_n1178_), .ZN(new_n1179_));
  NOR2_X1    g1130(.A1(new_n1179_), .A2(new_n1059_), .ZN(new_n1180_));
  XNOR2_X1   g1131(.A1(new_n839_), .A2(new_n932_), .ZN(new_n1181_));
  XNOR2_X1   g1132(.A1(new_n959_), .A2(new_n1181_), .ZN(new_n1182_));
  NOR2_X1    g1133(.A1(new_n1182_), .A2(new_n1180_), .ZN(new_n1183_));
  NAND2_X1   g1134(.A1(new_n1182_), .A2(new_n1180_), .ZN(new_n1184_));
  XOR2_X1    g1135(.A1(new_n808_), .A2(new_n783_), .Z(new_n1185_));
  XNOR2_X1   g1136(.A1(new_n816_), .A2(new_n1185_), .ZN(new_n1186_));
  AOI21_X1   g1137(.A1(new_n1184_), .A2(new_n1186_), .B(new_n1183_), .ZN(new_n1187_));
  INV_X1     g1138(.I(new_n1187_), .ZN(new_n1188_));
  XNOR2_X1   g1139(.A1(new_n830_), .A2(new_n833_), .ZN(new_n1189_));
  XOR2_X1    g1140(.A1(new_n1189_), .A2(new_n962_), .Z(new_n1190_));
  INV_X1     g1141(.I(new_n1190_), .ZN(new_n1191_));
  INV_X1     g1142(.I(new_n1183_), .ZN(new_n1192_));
  NAND2_X1   g1143(.A1(new_n1192_), .A2(new_n1184_), .ZN(new_n1193_));
  XOR2_X1    g1144(.A1(new_n1193_), .A2(new_n1186_), .Z(new_n1194_));
  INV_X1     g1145(.I(new_n1194_), .ZN(new_n1195_));
  XNOR2_X1   g1146(.A1(new_n1049_), .A2(new_n1058_), .ZN(new_n1196_));
  XNOR2_X1   g1147(.A1(new_n1196_), .A2(new_n1178_), .ZN(new_n1197_));
  XNOR2_X1   g1148(.A1(new_n938_), .A2(new_n951_), .ZN(new_n1198_));
  XNOR2_X1   g1149(.A1(new_n1198_), .A2(new_n957_), .ZN(new_n1199_));
  OR2_X2     g1150(.A1(new_n1197_), .A2(new_n1199_), .Z(new_n1200_));
  XOR2_X1    g1151(.A1(new_n1039_), .A2(new_n1040_), .Z(new_n1201_));
  XOR2_X1    g1152(.A1(new_n1201_), .A2(new_n1047_), .Z(new_n1202_));
  INV_X1     g1153(.I(new_n1202_), .ZN(new_n1203_));
  NOR2_X1    g1154(.A1(new_n1170_), .A2(new_n1176_), .ZN(new_n1204_));
  XOR2_X1    g1155(.A1(new_n1204_), .A2(new_n1175_), .Z(new_n1205_));
  NOR2_X1    g1156(.A1(new_n1205_), .A2(new_n1203_), .ZN(new_n1206_));
  NAND2_X1   g1157(.A1(new_n618_), .A2(new_n842_), .ZN(new_n1207_));
  NAND2_X1   g1158(.A1(new_n621_), .A2(new_n843_), .ZN(new_n1208_));
  NAND2_X1   g1159(.A1(new_n625_), .A2(new_n845_), .ZN(new_n1209_));
  NAND2_X1   g1160(.A1(new_n628_), .A2(new_n846_), .ZN(new_n1210_));
  AOI22_X1   g1161(.A1(new_n1209_), .A2(new_n1210_), .B1(new_n1207_), .B2(new_n1208_), .ZN(new_n1211_));
  NOR2_X1    g1162(.A1(new_n884_), .A2(new_n1032_), .ZN(new_n1212_));
  NOR2_X1    g1163(.A1(new_n998_), .A2(new_n929_), .ZN(new_n1213_));
  OAI21_X1   g1164(.A1(new_n1212_), .A2(new_n1213_), .B(new_n804_), .ZN(new_n1214_));
  NAND2_X1   g1165(.A1(new_n1214_), .A2(new_n598_), .ZN(new_n1215_));
  OAI21_X1   g1166(.A1(new_n1212_), .A2(new_n1213_), .B(new_n749_), .ZN(new_n1216_));
  NAND2_X1   g1167(.A1(new_n1216_), .A2(new_n465_), .ZN(new_n1217_));
  NOR2_X1    g1168(.A1(new_n884_), .A2(new_n929_), .ZN(new_n1218_));
  NOR2_X1    g1169(.A1(new_n998_), .A2(new_n1032_), .ZN(new_n1219_));
  AOI21_X1   g1170(.A1(new_n804_), .A2(new_n1219_), .B(new_n1218_), .ZN(new_n1220_));
  NAND2_X1   g1171(.A1(new_n1220_), .A2(new_n620_), .ZN(new_n1221_));
  OAI21_X1   g1172(.A1(new_n1219_), .A2(new_n1218_), .B(new_n1034_), .ZN(new_n1222_));
  NAND2_X1   g1173(.A1(new_n1222_), .A2(new_n462_), .ZN(new_n1223_));
  AOI22_X1   g1174(.A1(new_n1221_), .A2(new_n1223_), .B1(new_n1215_), .B2(new_n1217_), .ZN(new_n1224_));
  NOR2_X1    g1175(.A1(new_n1211_), .A2(new_n1224_), .ZN(new_n1225_));
  NOR2_X1    g1176(.A1(new_n762_), .A2(new_n663_), .ZN(new_n1226_));
  NOR2_X1    g1177(.A1(new_n766_), .A2(new_n664_), .ZN(new_n1227_));
  NOR2_X1    g1178(.A1(new_n812_), .A2(new_n671_), .ZN(new_n1228_));
  NOR2_X1    g1179(.A1(new_n814_), .A2(new_n670_), .ZN(new_n1229_));
  OAI22_X1   g1180(.A1(new_n1226_), .A2(new_n1227_), .B1(new_n1228_), .B2(new_n1229_), .ZN(new_n1230_));
  NAND2_X1   g1181(.A1(new_n1211_), .A2(new_n1224_), .ZN(new_n1231_));
  AOI21_X1   g1182(.A1(new_n1230_), .A2(new_n1231_), .B(new_n1225_), .ZN(new_n1232_));
  XNOR2_X1   g1183(.A1(new_n1204_), .A2(new_n1175_), .ZN(new_n1233_));
  NOR2_X1    g1184(.A1(new_n1233_), .A2(new_n1202_), .ZN(new_n1234_));
  NOR2_X1    g1185(.A1(new_n1234_), .A2(new_n1232_), .ZN(new_n1235_));
  NOR2_X1    g1186(.A1(new_n1235_), .A2(new_n1206_), .ZN(new_n1236_));
  NAND2_X1   g1187(.A1(new_n1197_), .A2(new_n1199_), .ZN(new_n1237_));
  INV_X1     g1188(.I(new_n1237_), .ZN(new_n1238_));
  OAI21_X1   g1189(.A1(new_n1236_), .A2(new_n1238_), .B(new_n1200_), .ZN(new_n1239_));
  NOR2_X1    g1190(.A1(new_n1195_), .A2(new_n1239_), .ZN(new_n1240_));
  INV_X1     g1191(.I(new_n1240_), .ZN(new_n1241_));
  NAND2_X1   g1192(.A1(new_n1195_), .A2(new_n1239_), .ZN(new_n1242_));
  NAND2_X1   g1193(.A1(new_n1241_), .A2(new_n1242_), .ZN(new_n1243_));
  INV_X1     g1194(.I(new_n1134_), .ZN(new_n1244_));
  NOR2_X1    g1195(.A1(new_n1167_), .A2(new_n1164_), .ZN(new_n1245_));
  XOR2_X1    g1196(.A1(new_n1245_), .A2(new_n1244_), .Z(new_n1246_));
  INV_X1     g1197(.I(new_n1246_), .ZN(new_n1247_));
  NOR2_X1    g1198(.A1(new_n1132_), .A2(new_n929_), .ZN(new_n1248_));
  INV_X1     g1199(.I(new_n730_), .ZN(new_n1249_));
  AOI21_X1   g1200(.A1(new_n108_), .A2(new_n121_), .B(new_n223_), .ZN(new_n1250_));
  AOI21_X1   g1201(.A1(new_n983_), .A2(new_n1250_), .B(new_n195_), .ZN(new_n1251_));
  NOR3_X1    g1202(.A1(new_n1251_), .A2(new_n317_), .A3(new_n487_), .ZN(new_n1252_));
  NAND3_X1   g1203(.A1(new_n1252_), .A2(new_n427_), .A3(new_n1249_), .ZN(new_n1253_));
  NOR2_X1    g1204(.A1(new_n1104_), .A2(new_n396_), .ZN(new_n1254_));
  NAND2_X1   g1205(.A1(new_n1254_), .A2(new_n1102_), .ZN(new_n1255_));
  NAND3_X1   g1206(.A1(new_n674_), .A2(new_n788_), .A3(new_n684_), .ZN(new_n1256_));
  NAND3_X1   g1207(.A1(new_n236_), .A2(new_n367_), .A3(new_n240_), .ZN(new_n1257_));
  NOR3_X1    g1208(.A1(new_n1256_), .A2(new_n1257_), .A3(new_n1107_), .ZN(new_n1258_));
  NOR4_X1    g1209(.A1(new_n185_), .A2(new_n516_), .A3(new_n691_), .A4(new_n313_), .ZN(new_n1259_));
  NAND4_X1   g1210(.A1(new_n989_), .A2(new_n255_), .A3(new_n303_), .A4(new_n685_), .ZN(new_n1260_));
  NAND4_X1   g1211(.A1(new_n216_), .A2(new_n73_), .A3(new_n154_), .A4(new_n162_), .ZN(new_n1261_));
  NAND4_X1   g1212(.A1(new_n329_), .A2(new_n224_), .A3(new_n714_), .A4(new_n1261_), .ZN(new_n1262_));
  NOR3_X1    g1213(.A1(new_n1260_), .A2(new_n1262_), .A3(new_n916_), .ZN(new_n1263_));
  NAND4_X1   g1214(.A1(new_n1263_), .A2(new_n1258_), .A3(new_n424_), .A4(new_n1259_), .ZN(new_n1264_));
  NAND2_X1   g1215(.A1(new_n909_), .A2(new_n908_), .ZN(new_n1265_));
  NAND2_X1   g1216(.A1(new_n366_), .A2(new_n482_), .ZN(new_n1266_));
  NAND4_X1   g1217(.A1(new_n1266_), .A2(new_n578_), .A3(new_n900_), .A4(new_n190_), .ZN(new_n1267_));
  NOR4_X1    g1218(.A1(new_n1267_), .A2(new_n1148_), .A3(new_n1265_), .A4(new_n1147_), .ZN(new_n1268_));
  NOR4_X1    g1219(.A1(new_n1153_), .A2(new_n405_), .A3(new_n700_), .A4(new_n1125_), .ZN(new_n1269_));
  NAND2_X1   g1220(.A1(new_n710_), .A2(new_n566_), .ZN(new_n1270_));
  NAND4_X1   g1221(.A1(new_n229_), .A2(new_n125_), .A3(new_n121_), .A4(new_n154_), .ZN(new_n1271_));
  NAND3_X1   g1222(.A1(new_n1271_), .A2(new_n228_), .A3(new_n676_), .ZN(new_n1272_));
  NOR4_X1    g1223(.A1(new_n1272_), .A2(new_n484_), .A3(new_n524_), .A4(new_n1270_), .ZN(new_n1273_));
  NAND3_X1   g1224(.A1(new_n1268_), .A2(new_n1273_), .A3(new_n1269_), .ZN(new_n1274_));
  NOR4_X1    g1225(.A1(new_n1264_), .A2(new_n1274_), .A3(new_n1253_), .A4(new_n1255_), .ZN(new_n1275_));
  NOR3_X1    g1226(.A1(new_n1032_), .A2(new_n1275_), .A3(new_n598_), .ZN(new_n1276_));
  OAI21_X1   g1227(.A1(new_n1276_), .A2(new_n1248_), .B(new_n1096_), .ZN(new_n1277_));
  INV_X1     g1228(.I(new_n1277_), .ZN(new_n1278_));
  AOI21_X1   g1229(.A1(new_n465_), .A2(new_n1275_), .B(new_n1134_), .ZN(new_n1279_));
  NOR2_X1    g1230(.A1(new_n1279_), .A2(new_n1278_), .ZN(new_n1280_));
  NOR2_X1    g1231(.A1(new_n1280_), .A2(new_n1157_), .ZN(new_n1281_));
  INV_X1     g1232(.I(new_n1281_), .ZN(new_n1282_));
  NOR2_X1    g1233(.A1(new_n1158_), .A2(\a[22] ), .ZN(new_n1283_));
  NOR2_X1    g1234(.A1(new_n1283_), .A2(\a[5] ), .ZN(new_n1284_));
  NAND2_X1   g1235(.A1(new_n1283_), .A2(\a[5] ), .ZN(new_n1285_));
  INV_X1     g1236(.I(new_n1285_), .ZN(new_n1286_));
  NOR2_X1    g1237(.A1(new_n1286_), .A2(new_n1284_), .ZN(new_n1287_));
  INV_X1     g1238(.I(new_n1287_), .ZN(new_n1288_));
  NOR2_X1    g1239(.A1(new_n469_), .A2(new_n1288_), .ZN(new_n1289_));
  NAND2_X1   g1240(.A1(new_n1280_), .A2(new_n1157_), .ZN(new_n1290_));
  NAND2_X1   g1241(.A1(new_n1290_), .A2(new_n1289_), .ZN(new_n1291_));
  NAND2_X1   g1242(.A1(new_n1291_), .A2(new_n1282_), .ZN(new_n1292_));
  NOR2_X1    g1243(.A1(new_n1247_), .A2(new_n1292_), .ZN(new_n1293_));
  NAND2_X1   g1244(.A1(new_n941_), .A2(new_n474_), .ZN(new_n1294_));
  NAND2_X1   g1245(.A1(new_n945_), .A2(new_n473_), .ZN(new_n1295_));
  NAND2_X1   g1246(.A1(new_n947_), .A2(new_n477_), .ZN(new_n1296_));
  NAND2_X1   g1247(.A1(new_n949_), .A2(new_n478_), .ZN(new_n1297_));
  AOI22_X1   g1248(.A1(new_n1295_), .A2(new_n1294_), .B1(new_n1296_), .B2(new_n1297_), .ZN(new_n1298_));
  AOI21_X1   g1249(.A1(new_n1247_), .A2(new_n1292_), .B(new_n1298_), .ZN(new_n1299_));
  NOR2_X1    g1250(.A1(new_n1299_), .A2(new_n1293_), .ZN(new_n1300_));
  NOR2_X1    g1251(.A1(new_n1234_), .A2(new_n1206_), .ZN(new_n1301_));
  XOR2_X1    g1252(.A1(new_n1301_), .A2(new_n1232_), .Z(new_n1302_));
  NOR2_X1    g1253(.A1(new_n1302_), .A2(new_n1300_), .ZN(new_n1303_));
  NOR2_X1    g1254(.A1(new_n944_), .A2(new_n671_), .ZN(new_n1304_));
  AOI21_X1   g1255(.A1(new_n671_), .A2(new_n941_), .B(new_n1304_), .ZN(new_n1305_));
  NOR2_X1    g1256(.A1(new_n1044_), .A2(new_n473_), .ZN(new_n1306_));
  AOI21_X1   g1257(.A1(new_n473_), .A2(new_n947_), .B(new_n1306_), .ZN(new_n1307_));
  NOR2_X1    g1258(.A1(new_n1305_), .A2(new_n1307_), .ZN(new_n1308_));
  NAND2_X1   g1259(.A1(new_n998_), .A2(new_n929_), .ZN(new_n1309_));
  NAND2_X1   g1260(.A1(new_n884_), .A2(new_n1032_), .ZN(new_n1310_));
  AOI21_X1   g1261(.A1(new_n1310_), .A2(new_n1309_), .B(new_n749_), .ZN(new_n1311_));
  NOR2_X1    g1262(.A1(new_n1311_), .A2(new_n462_), .ZN(new_n1312_));
  AOI21_X1   g1263(.A1(new_n462_), .A2(new_n1216_), .B(new_n1312_), .ZN(new_n1313_));
  NAND2_X1   g1264(.A1(new_n998_), .A2(new_n1032_), .ZN(new_n1314_));
  NAND2_X1   g1265(.A1(new_n884_), .A2(new_n929_), .ZN(new_n1315_));
  OAI21_X1   g1266(.A1(new_n749_), .A2(new_n1315_), .B(new_n1314_), .ZN(new_n1316_));
  NOR2_X1    g1267(.A1(new_n1316_), .A2(new_n477_), .ZN(new_n1317_));
  AOI21_X1   g1268(.A1(new_n477_), .A2(new_n1222_), .B(new_n1317_), .ZN(new_n1318_));
  NOR2_X1    g1269(.A1(new_n1318_), .A2(new_n1313_), .ZN(new_n1319_));
  NOR2_X1    g1270(.A1(new_n1308_), .A2(new_n1319_), .ZN(new_n1320_));
  NOR2_X1    g1271(.A1(new_n762_), .A2(new_n845_), .ZN(new_n1321_));
  NOR2_X1    g1272(.A1(new_n766_), .A2(new_n846_), .ZN(new_n1322_));
  NOR2_X1    g1273(.A1(new_n812_), .A2(new_n664_), .ZN(new_n1323_));
  NOR2_X1    g1274(.A1(new_n814_), .A2(new_n663_), .ZN(new_n1324_));
  OAI22_X1   g1275(.A1(new_n1321_), .A2(new_n1322_), .B1(new_n1323_), .B2(new_n1324_), .ZN(new_n1325_));
  NAND2_X1   g1276(.A1(new_n1308_), .A2(new_n1319_), .ZN(new_n1326_));
  AOI21_X1   g1277(.A1(new_n1325_), .A2(new_n1326_), .B(new_n1320_), .ZN(new_n1327_));
  INV_X1     g1278(.I(new_n1327_), .ZN(new_n1328_));
  XOR2_X1    g1279(.A1(new_n1211_), .A2(new_n1224_), .Z(new_n1329_));
  XOR2_X1    g1280(.A1(new_n1329_), .A2(new_n1230_), .Z(new_n1330_));
  NAND2_X1   g1281(.A1(new_n1330_), .A2(new_n1328_), .ZN(new_n1331_));
  INV_X1     g1282(.I(new_n1331_), .ZN(new_n1332_));
  NOR2_X1    g1283(.A1(new_n775_), .A2(new_n1162_), .ZN(new_n1333_));
  INV_X1     g1284(.I(new_n1333_), .ZN(new_n1334_));
  NAND2_X1   g1285(.A1(new_n621_), .A2(new_n1162_), .ZN(new_n1335_));
  NOR2_X1    g1286(.A1(new_n778_), .A2(new_n843_), .ZN(new_n1336_));
  INV_X1     g1287(.I(new_n1336_), .ZN(new_n1337_));
  NAND2_X1   g1288(.A1(new_n628_), .A2(new_n843_), .ZN(new_n1338_));
  AOI22_X1   g1289(.A1(new_n1334_), .A2(new_n1335_), .B1(new_n1337_), .B2(new_n1338_), .ZN(new_n1339_));
  NOR2_X1    g1290(.A1(new_n1132_), .A2(new_n1157_), .ZN(new_n1340_));
  NOR2_X1    g1291(.A1(new_n1275_), .A2(new_n1096_), .ZN(new_n1341_));
  OAI21_X1   g1292(.A1(new_n1340_), .A2(new_n1341_), .B(new_n929_), .ZN(new_n1342_));
  NAND2_X1   g1293(.A1(new_n1275_), .A2(new_n1096_), .ZN(new_n1343_));
  NAND2_X1   g1294(.A1(new_n1132_), .A2(new_n1157_), .ZN(new_n1344_));
  AOI21_X1   g1295(.A1(new_n1344_), .A2(new_n1343_), .B(new_n929_), .ZN(new_n1345_));
  NOR2_X1    g1296(.A1(new_n1345_), .A2(new_n598_), .ZN(new_n1346_));
  AOI21_X1   g1297(.A1(new_n598_), .A2(new_n1342_), .B(new_n1346_), .ZN(new_n1347_));
  NAND2_X1   g1298(.A1(new_n1275_), .A2(new_n1157_), .ZN(new_n1348_));
  NAND3_X1   g1299(.A1(new_n1132_), .A2(new_n1032_), .A3(new_n1096_), .ZN(new_n1349_));
  NAND2_X1   g1300(.A1(new_n1349_), .A2(new_n1348_), .ZN(new_n1350_));
  NOR2_X1    g1301(.A1(new_n1350_), .A2(new_n620_), .ZN(new_n1351_));
  INV_X1     g1302(.I(new_n1248_), .ZN(new_n1352_));
  NOR2_X1    g1303(.A1(new_n1340_), .A2(new_n1341_), .ZN(new_n1353_));
  NAND2_X1   g1304(.A1(new_n1353_), .A2(new_n1352_), .ZN(new_n1354_));
  AOI21_X1   g1305(.A1(new_n620_), .A2(new_n1354_), .B(new_n1351_), .ZN(new_n1355_));
  NOR2_X1    g1306(.A1(new_n1355_), .A2(new_n1347_), .ZN(new_n1356_));
  INV_X1     g1307(.I(new_n1356_), .ZN(new_n1357_));
  NOR2_X1    g1308(.A1(new_n68_), .A2(\a[22] ), .ZN(new_n1358_));
  XOR2_X1    g1309(.A1(new_n1358_), .A2(\a[4] ), .Z(new_n1359_));
  INV_X1     g1310(.I(new_n1359_), .ZN(new_n1360_));
  NOR2_X1    g1311(.A1(new_n469_), .A2(new_n1360_), .ZN(new_n1361_));
  NOR2_X1    g1312(.A1(new_n1361_), .A2(new_n1096_), .ZN(new_n1362_));
  NAND2_X1   g1313(.A1(new_n1361_), .A2(new_n1096_), .ZN(new_n1363_));
  OAI21_X1   g1314(.A1(new_n1357_), .A2(new_n1362_), .B(new_n1363_), .ZN(new_n1364_));
  OR2_X2     g1315(.A1(new_n1339_), .A2(new_n1364_), .Z(new_n1365_));
  NAND2_X1   g1316(.A1(new_n941_), .A2(new_n664_), .ZN(new_n1366_));
  NAND2_X1   g1317(.A1(new_n945_), .A2(new_n663_), .ZN(new_n1367_));
  NAND2_X1   g1318(.A1(new_n947_), .A2(new_n670_), .ZN(new_n1368_));
  NAND2_X1   g1319(.A1(new_n949_), .A2(new_n671_), .ZN(new_n1369_));
  AOI22_X1   g1320(.A1(new_n1366_), .A2(new_n1367_), .B1(new_n1368_), .B2(new_n1369_), .ZN(new_n1370_));
  NAND2_X1   g1321(.A1(new_n1214_), .A2(new_n478_), .ZN(new_n1371_));
  NAND2_X1   g1322(.A1(new_n1216_), .A2(new_n477_), .ZN(new_n1372_));
  NAND2_X1   g1323(.A1(new_n1220_), .A2(new_n474_), .ZN(new_n1373_));
  NAND2_X1   g1324(.A1(new_n1222_), .A2(new_n473_), .ZN(new_n1374_));
  AOI22_X1   g1325(.A1(new_n1373_), .A2(new_n1374_), .B1(new_n1371_), .B2(new_n1372_), .ZN(new_n1375_));
  NOR2_X1    g1326(.A1(new_n1370_), .A2(new_n1375_), .ZN(new_n1376_));
  NOR2_X1    g1327(.A1(new_n762_), .A2(new_n842_), .ZN(new_n1377_));
  NOR2_X1    g1328(.A1(new_n766_), .A2(new_n843_), .ZN(new_n1378_));
  NOR2_X1    g1329(.A1(new_n812_), .A2(new_n846_), .ZN(new_n1379_));
  NOR2_X1    g1330(.A1(new_n814_), .A2(new_n845_), .ZN(new_n1380_));
  OAI22_X1   g1331(.A1(new_n1377_), .A2(new_n1378_), .B1(new_n1379_), .B2(new_n1380_), .ZN(new_n1381_));
  NAND2_X1   g1332(.A1(new_n1370_), .A2(new_n1375_), .ZN(new_n1382_));
  AOI21_X1   g1333(.A1(new_n1381_), .A2(new_n1382_), .B(new_n1376_), .ZN(new_n1383_));
  NAND2_X1   g1334(.A1(new_n1339_), .A2(new_n1364_), .ZN(new_n1384_));
  INV_X1     g1335(.I(new_n1384_), .ZN(new_n1385_));
  OAI21_X1   g1336(.A1(new_n1385_), .A2(new_n1383_), .B(new_n1365_), .ZN(new_n1386_));
  XNOR2_X1   g1337(.A1(new_n1329_), .A2(new_n1230_), .ZN(new_n1387_));
  NAND2_X1   g1338(.A1(new_n1387_), .A2(new_n1327_), .ZN(new_n1388_));
  AOI21_X1   g1339(.A1(new_n1386_), .A2(new_n1388_), .B(new_n1332_), .ZN(new_n1389_));
  INV_X1     g1340(.I(new_n1389_), .ZN(new_n1390_));
  NAND2_X1   g1341(.A1(new_n1302_), .A2(new_n1300_), .ZN(new_n1391_));
  AOI21_X1   g1342(.A1(new_n1390_), .A2(new_n1391_), .B(new_n1303_), .ZN(new_n1392_));
  INV_X1     g1343(.I(new_n1392_), .ZN(new_n1393_));
  NAND2_X1   g1344(.A1(new_n1200_), .A2(new_n1237_), .ZN(new_n1394_));
  XOR2_X1    g1345(.A1(new_n1394_), .A2(new_n1236_), .Z(new_n1395_));
  NOR2_X1    g1346(.A1(new_n1393_), .A2(new_n1395_), .ZN(new_n1396_));
  INV_X1     g1347(.I(new_n1396_), .ZN(new_n1397_));
  NAND2_X1   g1348(.A1(new_n1393_), .A2(new_n1395_), .ZN(new_n1398_));
  INV_X1     g1349(.I(new_n1300_), .ZN(new_n1399_));
  XNOR2_X1   g1350(.A1(new_n1301_), .A2(new_n1232_), .ZN(new_n1400_));
  NAND2_X1   g1351(.A1(new_n1400_), .A2(new_n1399_), .ZN(new_n1401_));
  NAND2_X1   g1352(.A1(new_n1401_), .A2(new_n1391_), .ZN(new_n1402_));
  NOR2_X1    g1353(.A1(new_n1402_), .A2(new_n1390_), .ZN(new_n1403_));
  NOR2_X1    g1354(.A1(new_n1400_), .A2(new_n1399_), .ZN(new_n1404_));
  NOR2_X1    g1355(.A1(new_n1404_), .A2(new_n1303_), .ZN(new_n1405_));
  NOR2_X1    g1356(.A1(new_n1405_), .A2(new_n1389_), .ZN(new_n1406_));
  XOR2_X1    g1357(.A1(new_n1246_), .A2(new_n1292_), .Z(new_n1407_));
  XOR2_X1    g1358(.A1(new_n1407_), .A2(new_n1298_), .Z(new_n1408_));
  INV_X1     g1359(.I(new_n1408_), .ZN(new_n1409_));
  INV_X1     g1360(.I(new_n1326_), .ZN(new_n1410_));
  OR2_X2     g1361(.A1(new_n1410_), .A2(new_n1320_), .Z(new_n1411_));
  XOR2_X1    g1362(.A1(new_n1411_), .A2(new_n1325_), .Z(new_n1412_));
  AOI21_X1   g1363(.A1(new_n1290_), .A2(new_n1277_), .B(new_n1289_), .ZN(new_n1413_));
  NAND3_X1   g1364(.A1(new_n1282_), .A2(new_n1289_), .A3(new_n1290_), .ZN(new_n1414_));
  INV_X1     g1365(.I(new_n1414_), .ZN(new_n1415_));
  NOR2_X1    g1366(.A1(new_n1415_), .A2(new_n1413_), .ZN(new_n1416_));
  NOR2_X1    g1367(.A1(new_n1412_), .A2(new_n1416_), .ZN(new_n1417_));
  XNOR2_X1   g1368(.A1(new_n1411_), .A2(new_n1325_), .ZN(new_n1418_));
  INV_X1     g1369(.I(new_n1416_), .ZN(new_n1419_));
  NOR2_X1    g1370(.A1(new_n1418_), .A2(new_n1419_), .ZN(new_n1420_));
  NAND2_X1   g1371(.A1(new_n618_), .A2(new_n1287_), .ZN(new_n1421_));
  NAND2_X1   g1372(.A1(new_n621_), .A2(new_n1288_), .ZN(new_n1422_));
  NAND2_X1   g1373(.A1(new_n625_), .A2(new_n1161_), .ZN(new_n1423_));
  NAND2_X1   g1374(.A1(new_n628_), .A2(new_n1162_), .ZN(new_n1424_));
  AOI22_X1   g1375(.A1(new_n1423_), .A2(new_n1424_), .B1(new_n1421_), .B2(new_n1422_), .ZN(new_n1425_));
  NOR2_X1    g1376(.A1(new_n1345_), .A2(new_n620_), .ZN(new_n1426_));
  AOI21_X1   g1377(.A1(new_n620_), .A2(new_n1342_), .B(new_n1426_), .ZN(new_n1427_));
  NOR2_X1    g1378(.A1(new_n1350_), .A2(new_n478_), .ZN(new_n1428_));
  AOI21_X1   g1379(.A1(new_n478_), .A2(new_n1354_), .B(new_n1428_), .ZN(new_n1429_));
  NOR2_X1    g1380(.A1(new_n1429_), .A2(new_n1427_), .ZN(new_n1430_));
  NAND2_X1   g1381(.A1(new_n885_), .A2(new_n223_), .ZN(new_n1431_));
  NAND4_X1   g1382(.A1(new_n1431_), .A2(new_n275_), .A3(new_n875_), .A4(new_n556_), .ZN(new_n1432_));
  INV_X1     g1383(.I(new_n402_), .ZN(new_n1433_));
  NAND3_X1   g1384(.A1(new_n1433_), .A2(new_n410_), .A3(new_n433_), .ZN(new_n1434_));
  NAND2_X1   g1385(.A1(new_n565_), .A2(new_n528_), .ZN(new_n1435_));
  OR3_X2     g1386(.A1(new_n1432_), .A2(new_n1434_), .A3(new_n1435_), .Z(new_n1436_));
  NOR4_X1    g1387(.A1(new_n544_), .A2(new_n168_), .A3(new_n262_), .A4(new_n356_), .ZN(new_n1437_));
  NOR4_X1    g1388(.A1(new_n256_), .A2(new_n693_), .A3(new_n548_), .A4(new_n580_), .ZN(new_n1438_));
  NAND3_X1   g1389(.A1(new_n1438_), .A2(new_n1437_), .A3(new_n690_), .ZN(new_n1439_));
  OAI22_X1   g1390(.A1(new_n163_), .A2(new_n126_), .B1(new_n158_), .B2(new_n266_), .ZN(new_n1440_));
  NAND2_X1   g1391(.A1(new_n788_), .A2(new_n677_), .ZN(new_n1441_));
  NOR4_X1    g1392(.A1(new_n1441_), .A2(new_n269_), .A3(new_n1440_), .A4(new_n343_), .ZN(new_n1442_));
  NOR4_X1    g1393(.A1(new_n187_), .A2(new_n159_), .A3(new_n312_), .A4(new_n444_), .ZN(new_n1443_));
  NOR3_X1    g1394(.A1(new_n691_), .A2(new_n509_), .A3(new_n435_), .ZN(new_n1444_));
  NAND4_X1   g1395(.A1(new_n1442_), .A2(new_n526_), .A3(new_n1443_), .A4(new_n1444_), .ZN(new_n1445_));
  NOR4_X1    g1396(.A1(new_n248_), .A2(new_n1436_), .A3(new_n1445_), .A4(new_n1439_), .ZN(new_n1446_));
  AOI21_X1   g1397(.A1(new_n465_), .A2(new_n1446_), .B(new_n1157_), .ZN(new_n1447_));
  NOR2_X1    g1398(.A1(new_n1430_), .A2(new_n1447_), .ZN(new_n1448_));
  INV_X1     g1399(.I(\a[1] ), .ZN(new_n1449_));
  NOR2_X1    g1400(.A1(\a[0] ), .A2(\a[2] ), .ZN(new_n1450_));
  AOI21_X1   g1401(.A1(new_n1450_), .A2(new_n1449_), .B(\a[22] ), .ZN(new_n1451_));
  XOR2_X1    g1402(.A1(new_n1451_), .A2(\a[3] ), .Z(new_n1452_));
  INV_X1     g1403(.I(new_n1452_), .ZN(new_n1453_));
  NOR2_X1    g1404(.A1(new_n469_), .A2(new_n1453_), .ZN(new_n1454_));
  AND2_X2    g1405(.A1(new_n1430_), .A2(new_n1447_), .Z(new_n1455_));
  NOR2_X1    g1406(.A1(new_n1455_), .A2(new_n1454_), .ZN(new_n1456_));
  NOR2_X1    g1407(.A1(new_n1456_), .A2(new_n1448_), .ZN(new_n1457_));
  NOR2_X1    g1408(.A1(new_n1457_), .A2(new_n1425_), .ZN(new_n1458_));
  NAND2_X1   g1409(.A1(new_n769_), .A2(new_n842_), .ZN(new_n1459_));
  OAI21_X1   g1410(.A1(new_n814_), .A2(new_n842_), .B(new_n1459_), .ZN(new_n1460_));
  INV_X1     g1411(.I(new_n538_), .ZN(new_n1461_));
  NAND2_X1   g1412(.A1(new_n1461_), .A2(new_n592_), .ZN(new_n1462_));
  AOI21_X1   g1413(.A1(new_n423_), .A2(new_n1162_), .B(new_n538_), .ZN(new_n1463_));
  AOI21_X1   g1414(.A1(new_n422_), .A2(new_n1161_), .B(new_n636_), .ZN(new_n1464_));
  OAI21_X1   g1415(.A1(new_n1463_), .A2(new_n1464_), .B(new_n1462_), .ZN(new_n1465_));
  NAND2_X1   g1416(.A1(new_n1460_), .A2(new_n1465_), .ZN(new_n1466_));
  NOR2_X1    g1417(.A1(new_n1311_), .A2(new_n473_), .ZN(new_n1467_));
  AOI21_X1   g1418(.A1(new_n473_), .A2(new_n1216_), .B(new_n1467_), .ZN(new_n1468_));
  NOR2_X1    g1419(.A1(new_n1316_), .A2(new_n670_), .ZN(new_n1469_));
  AOI21_X1   g1420(.A1(new_n670_), .A2(new_n1222_), .B(new_n1469_), .ZN(new_n1470_));
  NOR2_X1    g1421(.A1(new_n1470_), .A2(new_n1468_), .ZN(new_n1471_));
  INV_X1     g1422(.I(new_n1471_), .ZN(new_n1472_));
  NAND2_X1   g1423(.A1(new_n1466_), .A2(new_n1472_), .ZN(new_n1473_));
  NAND2_X1   g1424(.A1(new_n941_), .A2(new_n846_), .ZN(new_n1474_));
  INV_X1     g1425(.I(new_n1474_), .ZN(new_n1475_));
  NOR2_X1    g1426(.A1(new_n944_), .A2(new_n846_), .ZN(new_n1476_));
  INV_X1     g1427(.I(new_n947_), .ZN(new_n1477_));
  NOR2_X1    g1428(.A1(new_n1477_), .A2(new_n664_), .ZN(new_n1478_));
  NOR2_X1    g1429(.A1(new_n1044_), .A2(new_n663_), .ZN(new_n1479_));
  OAI22_X1   g1430(.A1(new_n1475_), .A2(new_n1476_), .B1(new_n1478_), .B2(new_n1479_), .ZN(new_n1480_));
  NAND3_X1   g1431(.A1(new_n1460_), .A2(new_n1465_), .A3(new_n1471_), .ZN(new_n1481_));
  NAND2_X1   g1432(.A1(new_n1481_), .A2(new_n1480_), .ZN(new_n1482_));
  NAND2_X1   g1433(.A1(new_n1482_), .A2(new_n1473_), .ZN(new_n1483_));
  NAND2_X1   g1434(.A1(new_n1457_), .A2(new_n1425_), .ZN(new_n1484_));
  AOI21_X1   g1435(.A1(new_n1483_), .A2(new_n1484_), .B(new_n1458_), .ZN(new_n1485_));
  NOR2_X1    g1436(.A1(new_n1420_), .A2(new_n1485_), .ZN(new_n1486_));
  NOR2_X1    g1437(.A1(new_n1486_), .A2(new_n1417_), .ZN(new_n1487_));
  NOR2_X1    g1438(.A1(new_n1487_), .A2(new_n1409_), .ZN(new_n1488_));
  AND2_X2    g1439(.A1(new_n1388_), .A2(new_n1331_), .Z(new_n1489_));
  XOR2_X1    g1440(.A1(new_n1489_), .A2(new_n1386_), .Z(new_n1490_));
  NAND2_X1   g1441(.A1(new_n1487_), .A2(new_n1409_), .ZN(new_n1491_));
  AOI21_X1   g1442(.A1(new_n1490_), .A2(new_n1491_), .B(new_n1488_), .ZN(new_n1492_));
  INV_X1     g1443(.I(new_n1492_), .ZN(new_n1493_));
  OAI21_X1   g1444(.A1(new_n1406_), .A2(new_n1403_), .B(new_n1493_), .ZN(new_n1494_));
  NAND2_X1   g1445(.A1(new_n1405_), .A2(new_n1389_), .ZN(new_n1495_));
  NAND2_X1   g1446(.A1(new_n1402_), .A2(new_n1390_), .ZN(new_n1496_));
  NAND3_X1   g1447(.A1(new_n1495_), .A2(new_n1496_), .A3(new_n1492_), .ZN(new_n1497_));
  XNOR2_X1   g1448(.A1(new_n1489_), .A2(new_n1386_), .ZN(new_n1498_));
  INV_X1     g1449(.I(new_n1382_), .ZN(new_n1499_));
  NOR2_X1    g1450(.A1(new_n1499_), .A2(new_n1376_), .ZN(new_n1500_));
  XNOR2_X1   g1451(.A1(new_n1500_), .A2(new_n1381_), .ZN(new_n1501_));
  INV_X1     g1452(.I(new_n1501_), .ZN(new_n1502_));
  NAND2_X1   g1453(.A1(new_n613_), .A2(new_n1452_), .ZN(new_n1503_));
  NAND3_X1   g1454(.A1(new_n1503_), .A2(new_n365_), .A3(new_n459_), .ZN(new_n1504_));
  NAND2_X1   g1455(.A1(new_n206_), .A2(new_n211_), .ZN(new_n1505_));
  NOR2_X1    g1456(.A1(new_n452_), .A2(new_n337_), .ZN(new_n1506_));
  NOR3_X1    g1457(.A1(new_n234_), .A2(new_n330_), .A3(new_n722_), .ZN(new_n1507_));
  NAND4_X1   g1458(.A1(new_n486_), .A2(new_n1507_), .A3(new_n247_), .A4(new_n1506_), .ZN(new_n1508_));
  NOR2_X1    g1459(.A1(new_n1508_), .A2(new_n1505_), .ZN(new_n1509_));
  NOR3_X1    g1460(.A1(new_n1432_), .A2(new_n1434_), .A3(new_n1435_), .ZN(new_n1510_));
  OAI21_X1   g1461(.A1(new_n233_), .A2(new_n266_), .B(new_n551_), .ZN(new_n1511_));
  NAND3_X1   g1462(.A1(new_n993_), .A2(new_n151_), .A3(new_n908_), .ZN(new_n1512_));
  NAND4_X1   g1463(.A1(new_n581_), .A2(new_n255_), .A3(new_n491_), .A4(new_n412_), .ZN(new_n1513_));
  NOR4_X1    g1464(.A1(new_n1513_), .A2(new_n1512_), .A3(new_n356_), .A4(new_n1511_), .ZN(new_n1514_));
  INV_X1     g1465(.I(new_n312_), .ZN(new_n1515_));
  NAND4_X1   g1466(.A1(new_n1515_), .A2(new_n160_), .A3(new_n1068_), .A4(new_n1085_), .ZN(new_n1516_));
  NAND3_X1   g1467(.A1(new_n436_), .A2(new_n1092_), .A3(new_n1000_), .ZN(new_n1517_));
  NOR4_X1    g1468(.A1(new_n348_), .A2(new_n527_), .A3(new_n1516_), .A4(new_n1517_), .ZN(new_n1518_));
  NAND4_X1   g1469(.A1(new_n1509_), .A2(new_n1518_), .A3(new_n1510_), .A4(new_n1514_), .ZN(new_n1519_));
  NOR2_X1    g1470(.A1(new_n1519_), .A2(new_n462_), .ZN(new_n1520_));
  NOR2_X1    g1471(.A1(new_n1446_), .A2(new_n465_), .ZN(new_n1521_));
  OAI21_X1   g1472(.A1(new_n1520_), .A2(new_n1521_), .B(new_n1096_), .ZN(new_n1522_));
  NOR2_X1    g1473(.A1(new_n1446_), .A2(new_n1096_), .ZN(new_n1523_));
  NAND2_X1   g1474(.A1(new_n1523_), .A2(new_n465_), .ZN(new_n1524_));
  NAND2_X1   g1475(.A1(new_n1522_), .A2(new_n1524_), .ZN(new_n1525_));
  INV_X1     g1476(.I(new_n1525_), .ZN(new_n1526_));
  NOR2_X1    g1477(.A1(new_n1504_), .A2(new_n1526_), .ZN(new_n1527_));
  NOR2_X1    g1478(.A1(new_n778_), .A2(new_n1288_), .ZN(new_n1528_));
  AOI21_X1   g1479(.A1(new_n628_), .A2(new_n1288_), .B(new_n1528_), .ZN(new_n1529_));
  NOR2_X1    g1480(.A1(new_n775_), .A2(new_n1360_), .ZN(new_n1530_));
  AOI21_X1   g1481(.A1(new_n621_), .A2(new_n1360_), .B(new_n1530_), .ZN(new_n1531_));
  NOR3_X1    g1482(.A1(new_n1531_), .A2(new_n1529_), .A3(new_n1527_), .ZN(new_n1532_));
  INV_X1     g1483(.I(new_n1527_), .ZN(new_n1533_));
  NAND2_X1   g1484(.A1(new_n628_), .A2(new_n1288_), .ZN(new_n1534_));
  OAI21_X1   g1485(.A1(new_n778_), .A2(new_n1288_), .B(new_n1534_), .ZN(new_n1535_));
  NAND2_X1   g1486(.A1(new_n621_), .A2(new_n1360_), .ZN(new_n1536_));
  OAI21_X1   g1487(.A1(new_n775_), .A2(new_n1360_), .B(new_n1536_), .ZN(new_n1537_));
  AOI21_X1   g1488(.A1(new_n1537_), .A2(new_n1535_), .B(new_n1533_), .ZN(new_n1538_));
  NOR2_X1    g1489(.A1(new_n1532_), .A2(new_n1538_), .ZN(new_n1539_));
  NAND2_X1   g1490(.A1(new_n769_), .A2(new_n1161_), .ZN(new_n1540_));
  NAND2_X1   g1491(.A1(new_n771_), .A2(new_n1162_), .ZN(new_n1541_));
  NOR2_X1    g1492(.A1(new_n422_), .A2(new_n1287_), .ZN(new_n1542_));
  NOR2_X1    g1493(.A1(new_n423_), .A2(new_n1288_), .ZN(new_n1543_));
  OAI22_X1   g1494(.A1(new_n1543_), .A2(new_n636_), .B1(new_n538_), .B2(new_n1542_), .ZN(new_n1544_));
  AOI22_X1   g1495(.A1(new_n1540_), .A2(new_n1541_), .B1(new_n1462_), .B2(new_n1544_), .ZN(new_n1545_));
  INV_X1     g1496(.I(new_n1545_), .ZN(new_n1546_));
  AOI21_X1   g1497(.A1(new_n1310_), .A2(new_n1309_), .B(new_n804_), .ZN(new_n1547_));
  NOR2_X1    g1498(.A1(new_n1547_), .A2(new_n671_), .ZN(new_n1548_));
  AOI21_X1   g1499(.A1(new_n671_), .A2(new_n1214_), .B(new_n1548_), .ZN(new_n1549_));
  NOR2_X1    g1500(.A1(new_n1316_), .A2(new_n663_), .ZN(new_n1550_));
  AOI21_X1   g1501(.A1(new_n663_), .A2(new_n1222_), .B(new_n1550_), .ZN(new_n1551_));
  NOR2_X1    g1502(.A1(new_n1551_), .A2(new_n1549_), .ZN(new_n1552_));
  INV_X1     g1503(.I(new_n1552_), .ZN(new_n1553_));
  NAND2_X1   g1504(.A1(new_n1546_), .A2(new_n1553_), .ZN(new_n1554_));
  NAND2_X1   g1505(.A1(new_n941_), .A2(new_n843_), .ZN(new_n1555_));
  NAND2_X1   g1506(.A1(new_n945_), .A2(new_n842_), .ZN(new_n1556_));
  NAND2_X1   g1507(.A1(new_n947_), .A2(new_n845_), .ZN(new_n1557_));
  NAND2_X1   g1508(.A1(new_n949_), .A2(new_n846_), .ZN(new_n1558_));
  AOI22_X1   g1509(.A1(new_n1556_), .A2(new_n1555_), .B1(new_n1557_), .B2(new_n1558_), .ZN(new_n1559_));
  NAND2_X1   g1510(.A1(new_n1545_), .A2(new_n1552_), .ZN(new_n1560_));
  INV_X1     g1511(.I(new_n1560_), .ZN(new_n1561_));
  OAI21_X1   g1512(.A1(new_n1559_), .A2(new_n1561_), .B(new_n1554_), .ZN(new_n1562_));
  NOR2_X1    g1513(.A1(new_n1539_), .A2(new_n1562_), .ZN(new_n1563_));
  NOR3_X1    g1514(.A1(new_n1531_), .A2(new_n1533_), .A3(new_n1529_), .ZN(new_n1564_));
  NOR2_X1    g1515(.A1(new_n1563_), .A2(new_n1564_), .ZN(new_n1565_));
  INV_X1     g1516(.I(new_n1362_), .ZN(new_n1566_));
  NAND2_X1   g1517(.A1(new_n1566_), .A2(new_n1363_), .ZN(new_n1567_));
  XOR2_X1    g1518(.A1(new_n1567_), .A2(new_n1356_), .Z(new_n1568_));
  NOR2_X1    g1519(.A1(new_n1565_), .A2(new_n1568_), .ZN(new_n1569_));
  INV_X1     g1520(.I(new_n1569_), .ZN(new_n1570_));
  NAND2_X1   g1521(.A1(new_n1570_), .A2(new_n1502_), .ZN(new_n1571_));
  NAND2_X1   g1522(.A1(new_n1565_), .A2(new_n1568_), .ZN(new_n1572_));
  NAND2_X1   g1523(.A1(new_n1571_), .A2(new_n1572_), .ZN(new_n1573_));
  NAND2_X1   g1524(.A1(new_n1365_), .A2(new_n1384_), .ZN(new_n1574_));
  XOR2_X1    g1525(.A1(new_n1574_), .A2(new_n1383_), .Z(new_n1575_));
  NAND2_X1   g1526(.A1(new_n1573_), .A2(new_n1575_), .ZN(new_n1576_));
  INV_X1     g1527(.I(new_n1576_), .ZN(new_n1577_));
  NOR2_X1    g1528(.A1(new_n1573_), .A2(new_n1575_), .ZN(new_n1578_));
  NOR2_X1    g1529(.A1(new_n1420_), .A2(new_n1417_), .ZN(new_n1579_));
  XOR2_X1    g1530(.A1(new_n1579_), .A2(new_n1485_), .Z(new_n1580_));
  NOR2_X1    g1531(.A1(new_n1578_), .A2(new_n1580_), .ZN(new_n1581_));
  OAI21_X1   g1532(.A1(new_n1581_), .A2(new_n1577_), .B(new_n1498_), .ZN(new_n1582_));
  NOR2_X1    g1533(.A1(new_n1581_), .A2(new_n1577_), .ZN(new_n1583_));
  NAND2_X1   g1534(.A1(new_n1583_), .A2(new_n1490_), .ZN(new_n1584_));
  INV_X1     g1535(.I(new_n1491_), .ZN(new_n1585_));
  NOR2_X1    g1536(.A1(new_n1585_), .A2(new_n1488_), .ZN(new_n1586_));
  NAND3_X1   g1537(.A1(new_n1582_), .A2(new_n1584_), .A3(new_n1586_), .ZN(new_n1587_));
  NOR2_X1    g1538(.A1(new_n1583_), .A2(new_n1490_), .ZN(new_n1588_));
  NOR3_X1    g1539(.A1(new_n1498_), .A2(new_n1577_), .A3(new_n1581_), .ZN(new_n1589_));
  INV_X1     g1540(.I(new_n1586_), .ZN(new_n1590_));
  OAI21_X1   g1541(.A1(new_n1588_), .A2(new_n1589_), .B(new_n1590_), .ZN(new_n1591_));
  NAND2_X1   g1542(.A1(new_n1587_), .A2(new_n1591_), .ZN(new_n1592_));
  NAND2_X1   g1543(.A1(new_n1473_), .A2(new_n1481_), .ZN(new_n1593_));
  NAND2_X1   g1544(.A1(new_n1593_), .A2(new_n1480_), .ZN(new_n1594_));
  INV_X1     g1545(.I(new_n1480_), .ZN(new_n1595_));
  NAND3_X1   g1546(.A1(new_n1473_), .A2(new_n1595_), .A3(new_n1481_), .ZN(new_n1596_));
  NOR2_X1    g1547(.A1(new_n1455_), .A2(new_n1448_), .ZN(new_n1597_));
  XOR2_X1    g1548(.A1(new_n1597_), .A2(new_n1454_), .Z(new_n1598_));
  AOI21_X1   g1549(.A1(new_n1594_), .A2(new_n1596_), .B(new_n1598_), .ZN(new_n1599_));
  XOR2_X1    g1550(.A1(new_n1504_), .A2(new_n1525_), .Z(new_n1600_));
  AOI21_X1   g1551(.A1(new_n1344_), .A2(new_n1343_), .B(new_n1032_), .ZN(new_n1601_));
  NOR2_X1    g1552(.A1(new_n1601_), .A2(new_n477_), .ZN(new_n1602_));
  NOR2_X1    g1553(.A1(new_n1345_), .A2(new_n478_), .ZN(new_n1603_));
  NOR2_X1    g1554(.A1(new_n1350_), .A2(new_n474_), .ZN(new_n1604_));
  NAND2_X1   g1555(.A1(new_n1344_), .A2(new_n1343_), .ZN(new_n1605_));
  NOR2_X1    g1556(.A1(new_n1605_), .A2(new_n1248_), .ZN(new_n1606_));
  NOR2_X1    g1557(.A1(new_n1606_), .A2(new_n473_), .ZN(new_n1607_));
  OAI22_X1   g1558(.A1(new_n1607_), .A2(new_n1604_), .B1(new_n1602_), .B2(new_n1603_), .ZN(new_n1608_));
  NAND2_X1   g1559(.A1(new_n1600_), .A2(new_n1608_), .ZN(new_n1609_));
  NAND2_X1   g1560(.A1(new_n618_), .A2(new_n1452_), .ZN(new_n1610_));
  NAND2_X1   g1561(.A1(new_n621_), .A2(new_n1453_), .ZN(new_n1611_));
  NAND2_X1   g1562(.A1(new_n625_), .A2(new_n1359_), .ZN(new_n1612_));
  NAND2_X1   g1563(.A1(new_n628_), .A2(new_n1360_), .ZN(new_n1613_));
  AOI22_X1   g1564(.A1(new_n1612_), .A2(new_n1613_), .B1(new_n1610_), .B2(new_n1611_), .ZN(new_n1614_));
  NOR2_X1    g1565(.A1(new_n1600_), .A2(new_n1608_), .ZN(new_n1615_));
  OAI21_X1   g1566(.A1(new_n1614_), .A2(new_n1615_), .B(new_n1609_), .ZN(new_n1616_));
  NAND3_X1   g1567(.A1(new_n1598_), .A2(new_n1594_), .A3(new_n1596_), .ZN(new_n1617_));
  AOI21_X1   g1568(.A1(new_n1616_), .A2(new_n1617_), .B(new_n1599_), .ZN(new_n1618_));
  INV_X1     g1569(.I(new_n1618_), .ZN(new_n1619_));
  INV_X1     g1570(.I(new_n1484_), .ZN(new_n1620_));
  NOR2_X1    g1571(.A1(new_n1620_), .A2(new_n1458_), .ZN(new_n1621_));
  XOR2_X1    g1572(.A1(new_n1621_), .A2(new_n1483_), .Z(new_n1622_));
  NAND2_X1   g1573(.A1(new_n1622_), .A2(new_n1619_), .ZN(new_n1623_));
  NOR2_X1    g1574(.A1(new_n1622_), .A2(new_n1619_), .ZN(new_n1624_));
  NAND2_X1   g1575(.A1(new_n1570_), .A2(new_n1572_), .ZN(new_n1625_));
  XOR2_X1    g1576(.A1(new_n1625_), .A2(new_n1502_), .Z(new_n1626_));
  OAI21_X1   g1577(.A1(new_n1626_), .A2(new_n1624_), .B(new_n1623_), .ZN(new_n1627_));
  INV_X1     g1578(.I(new_n1578_), .ZN(new_n1628_));
  AOI21_X1   g1579(.A1(new_n1628_), .A2(new_n1576_), .B(new_n1580_), .ZN(new_n1629_));
  INV_X1     g1580(.I(new_n1580_), .ZN(new_n1630_));
  NOR3_X1    g1581(.A1(new_n1577_), .A2(new_n1630_), .A3(new_n1578_), .ZN(new_n1631_));
  NOR3_X1    g1582(.A1(new_n1631_), .A2(new_n1629_), .A3(new_n1627_), .ZN(new_n1632_));
  XOR2_X1    g1583(.A1(new_n1539_), .A2(new_n1562_), .Z(new_n1633_));
  NAND2_X1   g1584(.A1(new_n1594_), .A2(new_n1596_), .ZN(new_n1634_));
  INV_X1     g1585(.I(new_n1598_), .ZN(new_n1635_));
  NAND2_X1   g1586(.A1(new_n1634_), .A2(new_n1635_), .ZN(new_n1636_));
  INV_X1     g1587(.I(new_n1616_), .ZN(new_n1637_));
  NAND3_X1   g1588(.A1(new_n1636_), .A2(new_n1637_), .A3(new_n1617_), .ZN(new_n1638_));
  INV_X1     g1589(.I(new_n1617_), .ZN(new_n1639_));
  OAI21_X1   g1590(.A1(new_n1639_), .A2(new_n1599_), .B(new_n1616_), .ZN(new_n1640_));
  AOI21_X1   g1591(.A1(new_n1640_), .A2(new_n1638_), .B(new_n1633_), .ZN(new_n1641_));
  NOR2_X1    g1592(.A1(new_n1345_), .A2(new_n474_), .ZN(new_n1642_));
  AOI21_X1   g1593(.A1(new_n474_), .A2(new_n1342_), .B(new_n1642_), .ZN(new_n1643_));
  NOR2_X1    g1594(.A1(new_n1350_), .A2(new_n671_), .ZN(new_n1644_));
  AOI21_X1   g1595(.A1(new_n671_), .A2(new_n1354_), .B(new_n1644_), .ZN(new_n1645_));
  NOR2_X1    g1596(.A1(new_n1645_), .A2(new_n1643_), .ZN(new_n1646_));
  NAND2_X1   g1597(.A1(new_n1446_), .A2(new_n478_), .ZN(new_n1647_));
  OAI21_X1   g1598(.A1(new_n462_), .A2(new_n1446_), .B(new_n1647_), .ZN(new_n1648_));
  AOI22_X1   g1599(.A1(new_n1648_), .A2(new_n1096_), .B1(new_n462_), .B2(new_n1523_), .ZN(new_n1649_));
  INV_X1     g1600(.I(new_n1649_), .ZN(new_n1650_));
  NOR2_X1    g1601(.A1(new_n1646_), .A2(new_n1650_), .ZN(new_n1651_));
  NOR2_X1    g1602(.A1(new_n812_), .A2(new_n1288_), .ZN(new_n1652_));
  NOR2_X1    g1603(.A1(new_n814_), .A2(new_n1287_), .ZN(new_n1653_));
  AOI21_X1   g1604(.A1(new_n423_), .A2(new_n1360_), .B(new_n538_), .ZN(new_n1654_));
  AOI21_X1   g1605(.A1(new_n422_), .A2(new_n1359_), .B(new_n636_), .ZN(new_n1655_));
  OAI21_X1   g1606(.A1(new_n1654_), .A2(new_n1655_), .B(new_n1462_), .ZN(new_n1656_));
  OAI21_X1   g1607(.A1(new_n1653_), .A2(new_n1652_), .B(new_n1656_), .ZN(new_n1657_));
  NAND2_X1   g1608(.A1(new_n1646_), .A2(new_n1650_), .ZN(new_n1658_));
  AOI21_X1   g1609(.A1(new_n1657_), .A2(new_n1658_), .B(new_n1651_), .ZN(new_n1659_));
  NOR2_X1    g1610(.A1(new_n1545_), .A2(new_n1552_), .ZN(new_n1660_));
  NOR2_X1    g1611(.A1(new_n1561_), .A2(new_n1660_), .ZN(new_n1661_));
  NOR2_X1    g1612(.A1(new_n1661_), .A2(new_n1559_), .ZN(new_n1662_));
  INV_X1     g1613(.I(new_n1559_), .ZN(new_n1663_));
  NAND2_X1   g1614(.A1(new_n1554_), .A2(new_n1560_), .ZN(new_n1664_));
  NOR2_X1    g1615(.A1(new_n1664_), .A2(new_n1663_), .ZN(new_n1665_));
  NOR2_X1    g1616(.A1(new_n1662_), .A2(new_n1665_), .ZN(new_n1666_));
  NOR2_X1    g1617(.A1(new_n1666_), .A2(new_n1659_), .ZN(new_n1667_));
  NAND2_X1   g1618(.A1(new_n1157_), .A2(new_n1519_), .ZN(new_n1668_));
  NOR2_X1    g1619(.A1(new_n1519_), .A2(new_n473_), .ZN(new_n1669_));
  NOR2_X1    g1620(.A1(new_n1446_), .A2(new_n477_), .ZN(new_n1670_));
  NOR2_X1    g1621(.A1(new_n1669_), .A2(new_n1670_), .ZN(new_n1671_));
  OAI22_X1   g1622(.A1(new_n1671_), .A2(new_n1157_), .B1(new_n478_), .B2(new_n1668_), .ZN(new_n1672_));
  NOR2_X1    g1623(.A1(new_n758_), .A2(new_n1453_), .ZN(new_n1673_));
  NOR2_X1    g1624(.A1(new_n594_), .A2(new_n1673_), .ZN(new_n1674_));
  NAND2_X1   g1625(.A1(new_n1674_), .A2(new_n1672_), .ZN(new_n1675_));
  NOR2_X1    g1626(.A1(new_n1311_), .A2(new_n663_), .ZN(new_n1676_));
  NOR2_X1    g1627(.A1(new_n1547_), .A2(new_n664_), .ZN(new_n1677_));
  NOR2_X1    g1628(.A1(new_n1316_), .A2(new_n845_), .ZN(new_n1678_));
  AOI22_X1   g1629(.A1(new_n1314_), .A2(new_n1315_), .B1(new_n804_), .B2(new_n1032_), .ZN(new_n1679_));
  NOR2_X1    g1630(.A1(new_n1679_), .A2(new_n846_), .ZN(new_n1680_));
  OAI22_X1   g1631(.A1(new_n1680_), .A2(new_n1678_), .B1(new_n1676_), .B2(new_n1677_), .ZN(new_n1681_));
  NAND2_X1   g1632(.A1(new_n1675_), .A2(new_n1681_), .ZN(new_n1682_));
  NAND2_X1   g1633(.A1(new_n941_), .A2(new_n1162_), .ZN(new_n1683_));
  NAND2_X1   g1634(.A1(new_n945_), .A2(new_n1161_), .ZN(new_n1684_));
  NAND2_X1   g1635(.A1(new_n947_), .A2(new_n842_), .ZN(new_n1685_));
  NAND2_X1   g1636(.A1(new_n949_), .A2(new_n843_), .ZN(new_n1686_));
  AOI22_X1   g1637(.A1(new_n1684_), .A2(new_n1683_), .B1(new_n1685_), .B2(new_n1686_), .ZN(new_n1687_));
  NOR2_X1    g1638(.A1(new_n1675_), .A2(new_n1681_), .ZN(new_n1688_));
  OAI21_X1   g1639(.A1(new_n1687_), .A2(new_n1688_), .B(new_n1682_), .ZN(new_n1689_));
  NAND2_X1   g1640(.A1(new_n1666_), .A2(new_n1659_), .ZN(new_n1690_));
  AOI21_X1   g1641(.A1(new_n1689_), .A2(new_n1690_), .B(new_n1667_), .ZN(new_n1691_));
  INV_X1     g1642(.I(new_n1691_), .ZN(new_n1692_));
  NAND3_X1   g1643(.A1(new_n1640_), .A2(new_n1638_), .A3(new_n1633_), .ZN(new_n1693_));
  AOI21_X1   g1644(.A1(new_n1692_), .A2(new_n1693_), .B(new_n1641_), .ZN(new_n1694_));
  INV_X1     g1645(.I(new_n1689_), .ZN(new_n1695_));
  INV_X1     g1646(.I(new_n1659_), .ZN(new_n1696_));
  NAND2_X1   g1647(.A1(new_n1664_), .A2(new_n1663_), .ZN(new_n1697_));
  NAND2_X1   g1648(.A1(new_n1661_), .A2(new_n1559_), .ZN(new_n1698_));
  AOI21_X1   g1649(.A1(new_n1698_), .A2(new_n1697_), .B(new_n1696_), .ZN(new_n1699_));
  NOR3_X1    g1650(.A1(new_n1662_), .A2(new_n1665_), .A3(new_n1659_), .ZN(new_n1700_));
  OAI21_X1   g1651(.A1(new_n1699_), .A2(new_n1700_), .B(new_n1695_), .ZN(new_n1701_));
  OAI21_X1   g1652(.A1(new_n1662_), .A2(new_n1665_), .B(new_n1659_), .ZN(new_n1702_));
  NAND3_X1   g1653(.A1(new_n1698_), .A2(new_n1697_), .A3(new_n1696_), .ZN(new_n1703_));
  NAND3_X1   g1654(.A1(new_n1702_), .A2(new_n1703_), .A3(new_n1689_), .ZN(new_n1704_));
  INV_X1     g1655(.I(new_n1615_), .ZN(new_n1705_));
  AOI21_X1   g1656(.A1(new_n1705_), .A2(new_n1609_), .B(new_n1614_), .ZN(new_n1706_));
  INV_X1     g1657(.I(new_n1614_), .ZN(new_n1707_));
  NAND2_X1   g1658(.A1(new_n1705_), .A2(new_n1609_), .ZN(new_n1708_));
  NOR2_X1    g1659(.A1(new_n1708_), .A2(new_n1707_), .ZN(new_n1709_));
  NOR2_X1    g1660(.A1(new_n1709_), .A2(new_n1706_), .ZN(new_n1710_));
  AOI21_X1   g1661(.A1(new_n1701_), .A2(new_n1704_), .B(new_n1710_), .ZN(new_n1711_));
  XOR2_X1    g1662(.A1(new_n1675_), .A2(new_n1681_), .Z(new_n1712_));
  XOR2_X1    g1663(.A1(new_n1712_), .A2(new_n1687_), .Z(new_n1713_));
  NAND2_X1   g1664(.A1(new_n627_), .A2(new_n1452_), .ZN(new_n1714_));
  INV_X1     g1665(.I(new_n1714_), .ZN(new_n1715_));
  NOR2_X1    g1666(.A1(new_n1713_), .A2(new_n1715_), .ZN(new_n1716_));
  NAND2_X1   g1667(.A1(new_n1216_), .A2(new_n845_), .ZN(new_n1717_));
  OAI21_X1   g1668(.A1(new_n845_), .A2(new_n1311_), .B(new_n1717_), .ZN(new_n1718_));
  NAND2_X1   g1669(.A1(new_n1222_), .A2(new_n842_), .ZN(new_n1719_));
  OAI21_X1   g1670(.A1(new_n842_), .A2(new_n1316_), .B(new_n1719_), .ZN(new_n1720_));
  NAND2_X1   g1671(.A1(new_n1720_), .A2(new_n1718_), .ZN(new_n1721_));
  NOR2_X1    g1672(.A1(new_n1601_), .A2(new_n670_), .ZN(new_n1722_));
  NOR2_X1    g1673(.A1(new_n1345_), .A2(new_n671_), .ZN(new_n1723_));
  NOR2_X1    g1674(.A1(new_n1350_), .A2(new_n664_), .ZN(new_n1724_));
  NOR2_X1    g1675(.A1(new_n1606_), .A2(new_n663_), .ZN(new_n1725_));
  OAI22_X1   g1676(.A1(new_n1725_), .A2(new_n1724_), .B1(new_n1722_), .B2(new_n1723_), .ZN(new_n1726_));
  NAND2_X1   g1677(.A1(new_n941_), .A2(new_n1288_), .ZN(new_n1727_));
  NAND2_X1   g1678(.A1(new_n945_), .A2(new_n1287_), .ZN(new_n1728_));
  NAND2_X1   g1679(.A1(new_n947_), .A2(new_n1161_), .ZN(new_n1729_));
  NAND2_X1   g1680(.A1(new_n949_), .A2(new_n1162_), .ZN(new_n1730_));
  AOI22_X1   g1681(.A1(new_n1728_), .A2(new_n1727_), .B1(new_n1729_), .B2(new_n1730_), .ZN(new_n1731_));
  NOR2_X1    g1682(.A1(new_n1721_), .A2(new_n1726_), .ZN(new_n1732_));
  NOR2_X1    g1683(.A1(new_n1732_), .A2(new_n1731_), .ZN(new_n1733_));
  AOI21_X1   g1684(.A1(new_n1721_), .A2(new_n1726_), .B(new_n1733_), .ZN(new_n1734_));
  INV_X1     g1685(.I(new_n1734_), .ZN(new_n1735_));
  NAND2_X1   g1686(.A1(new_n1713_), .A2(new_n1715_), .ZN(new_n1736_));
  AOI21_X1   g1687(.A1(new_n1735_), .A2(new_n1736_), .B(new_n1716_), .ZN(new_n1737_));
  INV_X1     g1688(.I(new_n1737_), .ZN(new_n1738_));
  NAND3_X1   g1689(.A1(new_n1701_), .A2(new_n1704_), .A3(new_n1710_), .ZN(new_n1739_));
  AOI21_X1   g1690(.A1(new_n1738_), .A2(new_n1739_), .B(new_n1711_), .ZN(new_n1740_));
  XNOR2_X1   g1691(.A1(new_n1539_), .A2(new_n1562_), .ZN(new_n1741_));
  NOR3_X1    g1692(.A1(new_n1639_), .A2(new_n1599_), .A3(new_n1616_), .ZN(new_n1742_));
  AOI21_X1   g1693(.A1(new_n1636_), .A2(new_n1617_), .B(new_n1637_), .ZN(new_n1743_));
  OAI21_X1   g1694(.A1(new_n1742_), .A2(new_n1743_), .B(new_n1741_), .ZN(new_n1744_));
  NAND3_X1   g1695(.A1(new_n1744_), .A2(new_n1693_), .A3(new_n1691_), .ZN(new_n1745_));
  NOR3_X1    g1696(.A1(new_n1742_), .A2(new_n1743_), .A3(new_n1741_), .ZN(new_n1746_));
  OAI21_X1   g1697(.A1(new_n1746_), .A2(new_n1641_), .B(new_n1692_), .ZN(new_n1747_));
  NAND3_X1   g1698(.A1(new_n1747_), .A2(new_n1745_), .A3(new_n1740_), .ZN(new_n1748_));
  AOI21_X1   g1699(.A1(new_n1702_), .A2(new_n1703_), .B(new_n1689_), .ZN(new_n1749_));
  NOR3_X1    g1700(.A1(new_n1699_), .A2(new_n1700_), .A3(new_n1695_), .ZN(new_n1750_));
  XOR2_X1    g1701(.A1(new_n1708_), .A2(new_n1614_), .Z(new_n1751_));
  OAI21_X1   g1702(.A1(new_n1749_), .A2(new_n1750_), .B(new_n1751_), .ZN(new_n1752_));
  NAND3_X1   g1703(.A1(new_n1752_), .A2(new_n1738_), .A3(new_n1739_), .ZN(new_n1753_));
  NOR3_X1    g1704(.A1(new_n1751_), .A2(new_n1750_), .A3(new_n1749_), .ZN(new_n1754_));
  OAI21_X1   g1705(.A1(new_n1754_), .A2(new_n1711_), .B(new_n1737_), .ZN(new_n1755_));
  NOR2_X1    g1706(.A1(new_n1601_), .A2(new_n663_), .ZN(new_n1756_));
  NOR2_X1    g1707(.A1(new_n1345_), .A2(new_n664_), .ZN(new_n1757_));
  NOR2_X1    g1708(.A1(new_n1350_), .A2(new_n846_), .ZN(new_n1758_));
  NOR2_X1    g1709(.A1(new_n1606_), .A2(new_n845_), .ZN(new_n1759_));
  OAI22_X1   g1710(.A1(new_n1759_), .A2(new_n1758_), .B1(new_n1756_), .B2(new_n1757_), .ZN(new_n1760_));
  NAND2_X1   g1711(.A1(new_n1446_), .A2(new_n671_), .ZN(new_n1761_));
  OAI21_X1   g1712(.A1(new_n473_), .A2(new_n1446_), .B(new_n1761_), .ZN(new_n1762_));
  AOI22_X1   g1713(.A1(new_n1762_), .A2(new_n1096_), .B1(new_n473_), .B2(new_n1523_), .ZN(new_n1763_));
  NAND2_X1   g1714(.A1(new_n1760_), .A2(new_n1763_), .ZN(new_n1764_));
  NAND2_X1   g1715(.A1(new_n1214_), .A2(new_n843_), .ZN(new_n1765_));
  NAND2_X1   g1716(.A1(new_n1216_), .A2(new_n842_), .ZN(new_n1766_));
  NAND2_X1   g1717(.A1(new_n1220_), .A2(new_n1162_), .ZN(new_n1767_));
  NAND2_X1   g1718(.A1(new_n1222_), .A2(new_n1161_), .ZN(new_n1768_));
  AOI22_X1   g1719(.A1(new_n1767_), .A2(new_n1768_), .B1(new_n1765_), .B2(new_n1766_), .ZN(new_n1769_));
  NOR2_X1    g1720(.A1(new_n1760_), .A2(new_n1763_), .ZN(new_n1770_));
  OAI21_X1   g1721(.A1(new_n1769_), .A2(new_n1770_), .B(new_n1764_), .ZN(new_n1771_));
  XNOR2_X1   g1722(.A1(new_n1674_), .A2(new_n1672_), .ZN(new_n1772_));
  NAND2_X1   g1723(.A1(new_n1771_), .A2(new_n1772_), .ZN(new_n1773_));
  INV_X1     g1724(.I(new_n1773_), .ZN(new_n1774_));
  NAND2_X1   g1725(.A1(new_n763_), .A2(new_n1453_), .ZN(new_n1775_));
  NAND2_X1   g1726(.A1(new_n767_), .A2(new_n1452_), .ZN(new_n1776_));
  NAND2_X1   g1727(.A1(new_n769_), .A2(new_n1359_), .ZN(new_n1777_));
  NAND2_X1   g1728(.A1(new_n771_), .A2(new_n1360_), .ZN(new_n1778_));
  AOI22_X1   g1729(.A1(new_n1776_), .A2(new_n1775_), .B1(new_n1777_), .B2(new_n1778_), .ZN(new_n1779_));
  INV_X1     g1730(.I(new_n1779_), .ZN(new_n1780_));
  OR2_X2     g1731(.A1(new_n1771_), .A2(new_n1772_), .Z(new_n1781_));
  AOI21_X1   g1732(.A1(new_n1780_), .A2(new_n1781_), .B(new_n1774_), .ZN(new_n1782_));
  INV_X1     g1733(.I(new_n1651_), .ZN(new_n1783_));
  NAND2_X1   g1734(.A1(new_n1783_), .A2(new_n1658_), .ZN(new_n1784_));
  XOR2_X1    g1735(.A1(new_n1784_), .A2(new_n1657_), .Z(new_n1785_));
  NOR2_X1    g1736(.A1(new_n1782_), .A2(new_n1785_), .ZN(new_n1786_));
  INV_X1     g1737(.I(new_n1786_), .ZN(new_n1787_));
  NAND2_X1   g1738(.A1(new_n1782_), .A2(new_n1785_), .ZN(new_n1788_));
  XNOR2_X1   g1739(.A1(new_n1712_), .A2(new_n1687_), .ZN(new_n1789_));
  NOR2_X1    g1740(.A1(new_n1789_), .A2(new_n1714_), .ZN(new_n1790_));
  NOR2_X1    g1741(.A1(new_n1790_), .A2(new_n1716_), .ZN(new_n1791_));
  NOR2_X1    g1742(.A1(new_n1791_), .A2(new_n1734_), .ZN(new_n1792_));
  NAND2_X1   g1743(.A1(new_n1789_), .A2(new_n1714_), .ZN(new_n1793_));
  NAND2_X1   g1744(.A1(new_n1793_), .A2(new_n1736_), .ZN(new_n1794_));
  NOR2_X1    g1745(.A1(new_n1794_), .A2(new_n1735_), .ZN(new_n1795_));
  OAI21_X1   g1746(.A1(new_n1792_), .A2(new_n1795_), .B(new_n1788_), .ZN(new_n1796_));
  NAND2_X1   g1747(.A1(new_n1796_), .A2(new_n1787_), .ZN(new_n1797_));
  AOI21_X1   g1748(.A1(new_n1753_), .A2(new_n1755_), .B(new_n1797_), .ZN(new_n1798_));
  NAND2_X1   g1749(.A1(new_n1214_), .A2(new_n1162_), .ZN(new_n1799_));
  NAND2_X1   g1750(.A1(new_n1216_), .A2(new_n1161_), .ZN(new_n1800_));
  NAND2_X1   g1751(.A1(new_n1799_), .A2(new_n1800_), .ZN(new_n1801_));
  NAND2_X1   g1752(.A1(new_n1220_), .A2(new_n1288_), .ZN(new_n1802_));
  NAND2_X1   g1753(.A1(new_n1222_), .A2(new_n1287_), .ZN(new_n1803_));
  NAND2_X1   g1754(.A1(new_n1802_), .A2(new_n1803_), .ZN(new_n1804_));
  NAND2_X1   g1755(.A1(new_n1342_), .A2(new_n846_), .ZN(new_n1805_));
  OAI21_X1   g1756(.A1(new_n1340_), .A2(new_n1341_), .B(new_n1032_), .ZN(new_n1806_));
  NAND2_X1   g1757(.A1(new_n1806_), .A2(new_n845_), .ZN(new_n1807_));
  NAND2_X1   g1758(.A1(new_n1805_), .A2(new_n1807_), .ZN(new_n1808_));
  NAND3_X1   g1759(.A1(new_n1349_), .A2(new_n1348_), .A3(new_n842_), .ZN(new_n1809_));
  OAI21_X1   g1760(.A1(new_n1606_), .A2(new_n842_), .B(new_n1809_), .ZN(new_n1810_));
  AOI22_X1   g1761(.A1(new_n1804_), .A2(new_n1801_), .B1(new_n1808_), .B2(new_n1810_), .ZN(new_n1811_));
  NAND2_X1   g1762(.A1(new_n947_), .A2(new_n1359_), .ZN(new_n1812_));
  INV_X1     g1763(.I(new_n1812_), .ZN(new_n1813_));
  NOR2_X1    g1764(.A1(new_n1044_), .A2(new_n1359_), .ZN(new_n1814_));
  NAND2_X1   g1765(.A1(new_n785_), .A2(new_n749_), .ZN(new_n1815_));
  NOR2_X1    g1766(.A1(new_n636_), .A2(new_n1452_), .ZN(new_n1816_));
  NOR2_X1    g1767(.A1(new_n592_), .A2(new_n1453_), .ZN(new_n1817_));
  OAI22_X1   g1768(.A1(new_n1816_), .A2(new_n705_), .B1(new_n804_), .B2(new_n1817_), .ZN(new_n1818_));
  NAND2_X1   g1769(.A1(new_n1818_), .A2(new_n1815_), .ZN(new_n1819_));
  OAI21_X1   g1770(.A1(new_n1813_), .A2(new_n1814_), .B(new_n1819_), .ZN(new_n1820_));
  NAND4_X1   g1771(.A1(new_n1804_), .A2(new_n1801_), .A3(new_n1808_), .A4(new_n1810_), .ZN(new_n1821_));
  AOI21_X1   g1772(.A1(new_n1820_), .A2(new_n1821_), .B(new_n1811_), .ZN(new_n1822_));
  INV_X1     g1773(.I(new_n1822_), .ZN(new_n1823_));
  INV_X1     g1774(.I(new_n1769_), .ZN(new_n1824_));
  NOR2_X1    g1775(.A1(new_n1756_), .A2(new_n1757_), .ZN(new_n1825_));
  AOI21_X1   g1776(.A1(new_n846_), .A2(new_n1354_), .B(new_n1758_), .ZN(new_n1826_));
  NOR2_X1    g1777(.A1(new_n1826_), .A2(new_n1825_), .ZN(new_n1827_));
  INV_X1     g1778(.I(new_n1763_), .ZN(new_n1828_));
  NAND2_X1   g1779(.A1(new_n1827_), .A2(new_n1828_), .ZN(new_n1829_));
  NAND2_X1   g1780(.A1(new_n1829_), .A2(new_n1764_), .ZN(new_n1830_));
  NOR2_X1    g1781(.A1(new_n1830_), .A2(new_n1824_), .ZN(new_n1831_));
  NOR2_X1    g1782(.A1(new_n1827_), .A2(new_n1828_), .ZN(new_n1832_));
  NOR2_X1    g1783(.A1(new_n1832_), .A2(new_n1770_), .ZN(new_n1833_));
  NOR2_X1    g1784(.A1(new_n1833_), .A2(new_n1769_), .ZN(new_n1834_));
  OAI21_X1   g1785(.A1(new_n1834_), .A2(new_n1831_), .B(new_n1823_), .ZN(new_n1835_));
  INV_X1     g1786(.I(new_n1835_), .ZN(new_n1836_));
  NOR2_X1    g1787(.A1(new_n760_), .A2(new_n1453_), .ZN(new_n1837_));
  NAND2_X1   g1788(.A1(new_n941_), .A2(new_n1360_), .ZN(new_n1838_));
  NAND2_X1   g1789(.A1(new_n945_), .A2(new_n1359_), .ZN(new_n1839_));
  NAND2_X1   g1790(.A1(new_n947_), .A2(new_n1287_), .ZN(new_n1840_));
  NAND2_X1   g1791(.A1(new_n949_), .A2(new_n1288_), .ZN(new_n1841_));
  AOI22_X1   g1792(.A1(new_n1839_), .A2(new_n1838_), .B1(new_n1840_), .B2(new_n1841_), .ZN(new_n1842_));
  NAND2_X1   g1793(.A1(new_n1446_), .A2(new_n664_), .ZN(new_n1843_));
  NAND2_X1   g1794(.A1(new_n1519_), .A2(new_n671_), .ZN(new_n1844_));
  AOI21_X1   g1795(.A1(new_n1844_), .A2(new_n1843_), .B(new_n1157_), .ZN(new_n1845_));
  NOR2_X1    g1796(.A1(new_n1668_), .A2(new_n671_), .ZN(new_n1846_));
  NOR2_X1    g1797(.A1(new_n1845_), .A2(new_n1846_), .ZN(new_n1847_));
  NOR2_X1    g1798(.A1(new_n940_), .A2(new_n1453_), .ZN(new_n1848_));
  NOR3_X1    g1799(.A1(new_n1847_), .A2(new_n751_), .A3(new_n1848_), .ZN(new_n1849_));
  NAND2_X1   g1800(.A1(new_n1842_), .A2(new_n1849_), .ZN(new_n1850_));
  INV_X1     g1801(.I(new_n1850_), .ZN(new_n1851_));
  NOR2_X1    g1802(.A1(new_n1842_), .A2(new_n1849_), .ZN(new_n1852_));
  NOR3_X1    g1803(.A1(new_n1851_), .A2(new_n1837_), .A3(new_n1852_), .ZN(new_n1853_));
  INV_X1     g1804(.I(new_n1837_), .ZN(new_n1854_));
  INV_X1     g1805(.I(new_n1852_), .ZN(new_n1855_));
  AOI21_X1   g1806(.A1(new_n1855_), .A2(new_n1850_), .B(new_n1854_), .ZN(new_n1856_));
  NOR2_X1    g1807(.A1(new_n1856_), .A2(new_n1853_), .ZN(new_n1857_));
  NAND2_X1   g1808(.A1(new_n1833_), .A2(new_n1769_), .ZN(new_n1858_));
  NAND2_X1   g1809(.A1(new_n1830_), .A2(new_n1824_), .ZN(new_n1859_));
  NAND3_X1   g1810(.A1(new_n1858_), .A2(new_n1859_), .A3(new_n1822_), .ZN(new_n1860_));
  AOI21_X1   g1811(.A1(new_n1857_), .A2(new_n1860_), .B(new_n1836_), .ZN(new_n1861_));
  INV_X1     g1812(.I(new_n1861_), .ZN(new_n1862_));
  NOR2_X1    g1813(.A1(new_n1311_), .A2(new_n1359_), .ZN(new_n1863_));
  NAND2_X1   g1814(.A1(new_n1310_), .A2(new_n1309_), .ZN(new_n1864_));
  AOI21_X1   g1815(.A1(new_n1864_), .A2(new_n749_), .B(new_n1360_), .ZN(new_n1865_));
  NAND3_X1   g1816(.A1(new_n998_), .A2(new_n804_), .A3(new_n1452_), .ZN(new_n1866_));
  NAND3_X1   g1817(.A1(new_n749_), .A2(new_n884_), .A3(new_n1453_), .ZN(new_n1867_));
  NAND4_X1   g1818(.A1(new_n1867_), .A2(new_n1866_), .A3(new_n1310_), .A4(new_n1309_), .ZN(new_n1868_));
  OAI21_X1   g1819(.A1(new_n1863_), .A2(new_n1865_), .B(new_n1868_), .ZN(new_n1869_));
  NOR2_X1    g1820(.A1(new_n1519_), .A2(new_n842_), .ZN(new_n1870_));
  NOR2_X1    g1821(.A1(new_n1446_), .A2(new_n845_), .ZN(new_n1871_));
  OAI21_X1   g1822(.A1(new_n1870_), .A2(new_n1871_), .B(new_n1096_), .ZN(new_n1872_));
  NOR3_X1    g1823(.A1(new_n1446_), .A2(new_n1096_), .A3(new_n846_), .ZN(new_n1873_));
  INV_X1     g1824(.I(new_n1873_), .ZN(new_n1874_));
  OAI21_X1   g1825(.A1(new_n998_), .A2(new_n1032_), .B(new_n1452_), .ZN(new_n1875_));
  AOI22_X1   g1826(.A1(new_n1872_), .A2(new_n1874_), .B1(new_n1050_), .B2(new_n1875_), .ZN(new_n1876_));
  NOR4_X1    g1827(.A1(new_n343_), .A2(new_n346_), .A3(new_n345_), .A4(new_n269_), .ZN(new_n1877_));
  NAND4_X1   g1828(.A1(new_n1877_), .A2(new_n1444_), .A3(new_n526_), .A4(new_n342_), .ZN(new_n1878_));
  NOR4_X1    g1829(.A1(new_n1878_), .A2(new_n1508_), .A3(new_n1505_), .A4(new_n1516_), .ZN(new_n1879_));
  NAND4_X1   g1830(.A1(new_n1879_), .A2(new_n843_), .A3(new_n1510_), .A4(new_n1514_), .ZN(new_n1880_));
  NAND2_X1   g1831(.A1(new_n1519_), .A2(new_n846_), .ZN(new_n1881_));
  AOI21_X1   g1832(.A1(new_n1881_), .A2(new_n1880_), .B(new_n1157_), .ZN(new_n1882_));
  AOI21_X1   g1833(.A1(new_n884_), .A2(new_n929_), .B(new_n1453_), .ZN(new_n1883_));
  NOR4_X1    g1834(.A1(new_n1882_), .A2(new_n930_), .A3(new_n1873_), .A4(new_n1883_), .ZN(new_n1884_));
  NOR2_X1    g1835(.A1(new_n1876_), .A2(new_n1884_), .ZN(new_n1885_));
  NAND2_X1   g1836(.A1(new_n1869_), .A2(new_n1885_), .ZN(new_n1886_));
  NOR2_X1    g1837(.A1(new_n1601_), .A2(new_n1161_), .ZN(new_n1887_));
  NOR2_X1    g1838(.A1(new_n1345_), .A2(new_n1162_), .ZN(new_n1888_));
  NOR2_X1    g1839(.A1(new_n1887_), .A2(new_n1888_), .ZN(new_n1889_));
  NOR2_X1    g1840(.A1(new_n1132_), .A2(new_n1096_), .ZN(new_n1890_));
  NOR3_X1    g1841(.A1(new_n1157_), .A2(new_n1275_), .A3(new_n929_), .ZN(new_n1891_));
  NOR3_X1    g1842(.A1(new_n1891_), .A2(new_n1890_), .A3(new_n1288_), .ZN(new_n1892_));
  AOI21_X1   g1843(.A1(new_n1354_), .A2(new_n1288_), .B(new_n1892_), .ZN(new_n1893_));
  OAI22_X1   g1844(.A1(new_n1869_), .A2(new_n1885_), .B1(new_n1889_), .B2(new_n1893_), .ZN(new_n1894_));
  NAND2_X1   g1845(.A1(new_n1848_), .A2(new_n750_), .ZN(new_n1895_));
  INV_X1     g1846(.I(new_n1895_), .ZN(new_n1896_));
  AOI21_X1   g1847(.A1(new_n1894_), .A2(new_n1886_), .B(new_n1896_), .ZN(new_n1897_));
  NAND2_X1   g1848(.A1(new_n1214_), .A2(new_n1360_), .ZN(new_n1898_));
  NAND2_X1   g1849(.A1(new_n1216_), .A2(new_n1359_), .ZN(new_n1899_));
  NOR3_X1    g1850(.A1(new_n749_), .A2(new_n884_), .A3(new_n1453_), .ZN(new_n1900_));
  NOR3_X1    g1851(.A1(new_n998_), .A2(new_n804_), .A3(new_n1452_), .ZN(new_n1901_));
  NOR4_X1    g1852(.A1(new_n1900_), .A2(new_n1901_), .A3(new_n1212_), .A4(new_n1213_), .ZN(new_n1902_));
  AOI21_X1   g1853(.A1(new_n1898_), .A2(new_n1899_), .B(new_n1902_), .ZN(new_n1903_));
  OAI22_X1   g1854(.A1(new_n1882_), .A2(new_n1873_), .B1(new_n930_), .B2(new_n1883_), .ZN(new_n1904_));
  NAND4_X1   g1855(.A1(new_n1872_), .A2(new_n1050_), .A3(new_n1874_), .A4(new_n1875_), .ZN(new_n1905_));
  NAND2_X1   g1856(.A1(new_n1905_), .A2(new_n1904_), .ZN(new_n1906_));
  NOR2_X1    g1857(.A1(new_n1903_), .A2(new_n1906_), .ZN(new_n1907_));
  NAND2_X1   g1858(.A1(new_n1342_), .A2(new_n1162_), .ZN(new_n1908_));
  NAND2_X1   g1859(.A1(new_n1806_), .A2(new_n1161_), .ZN(new_n1909_));
  NAND2_X1   g1860(.A1(new_n1908_), .A2(new_n1909_), .ZN(new_n1910_));
  NAND3_X1   g1861(.A1(new_n1349_), .A2(new_n1348_), .A3(new_n1287_), .ZN(new_n1911_));
  OAI21_X1   g1862(.A1(new_n1606_), .A2(new_n1287_), .B(new_n1911_), .ZN(new_n1912_));
  AOI22_X1   g1863(.A1(new_n1903_), .A2(new_n1906_), .B1(new_n1910_), .B2(new_n1912_), .ZN(new_n1913_));
  NOR3_X1    g1864(.A1(new_n1913_), .A2(new_n1907_), .A3(new_n1895_), .ZN(new_n1914_));
  NOR2_X1    g1865(.A1(new_n930_), .A2(new_n1883_), .ZN(new_n1915_));
  OAI21_X1   g1866(.A1(new_n1882_), .A2(new_n1873_), .B(new_n1915_), .ZN(new_n1916_));
  OAI21_X1   g1867(.A1(new_n1914_), .A2(new_n1897_), .B(new_n1916_), .ZN(new_n1917_));
  OAI21_X1   g1868(.A1(new_n1913_), .A2(new_n1907_), .B(new_n1895_), .ZN(new_n1918_));
  NAND3_X1   g1869(.A1(new_n1894_), .A2(new_n1886_), .A3(new_n1896_), .ZN(new_n1919_));
  INV_X1     g1870(.I(new_n1916_), .ZN(new_n1920_));
  NAND3_X1   g1871(.A1(new_n1918_), .A2(new_n1919_), .A3(new_n1920_), .ZN(new_n1921_));
  NAND2_X1   g1872(.A1(new_n1214_), .A2(new_n1288_), .ZN(new_n1922_));
  NAND2_X1   g1873(.A1(new_n1216_), .A2(new_n1287_), .ZN(new_n1923_));
  NAND2_X1   g1874(.A1(new_n1922_), .A2(new_n1923_), .ZN(new_n1924_));
  NAND2_X1   g1875(.A1(new_n1220_), .A2(new_n1360_), .ZN(new_n1925_));
  NAND2_X1   g1876(.A1(new_n1222_), .A2(new_n1359_), .ZN(new_n1926_));
  NAND2_X1   g1877(.A1(new_n1925_), .A2(new_n1926_), .ZN(new_n1927_));
  NAND2_X1   g1878(.A1(new_n1927_), .A2(new_n1924_), .ZN(new_n1928_));
  NOR2_X1    g1879(.A1(new_n1601_), .A2(new_n842_), .ZN(new_n1929_));
  NOR2_X1    g1880(.A1(new_n1345_), .A2(new_n843_), .ZN(new_n1930_));
  NAND3_X1   g1881(.A1(new_n1349_), .A2(new_n1348_), .A3(new_n1161_), .ZN(new_n1931_));
  INV_X1     g1882(.I(new_n1931_), .ZN(new_n1932_));
  AOI21_X1   g1883(.A1(new_n1353_), .A2(new_n1352_), .B(new_n1161_), .ZN(new_n1933_));
  OAI22_X1   g1884(.A1(new_n1929_), .A2(new_n1930_), .B1(new_n1933_), .B2(new_n1932_), .ZN(new_n1934_));
  NAND2_X1   g1885(.A1(new_n1446_), .A2(new_n846_), .ZN(new_n1935_));
  OAI21_X1   g1886(.A1(new_n663_), .A2(new_n1446_), .B(new_n1935_), .ZN(new_n1936_));
  AOI22_X1   g1887(.A1(new_n1936_), .A2(new_n1096_), .B1(new_n663_), .B2(new_n1523_), .ZN(new_n1937_));
  NOR2_X1    g1888(.A1(new_n1934_), .A2(new_n1937_), .ZN(new_n1938_));
  NAND2_X1   g1889(.A1(new_n1342_), .A2(new_n843_), .ZN(new_n1939_));
  NAND2_X1   g1890(.A1(new_n1806_), .A2(new_n842_), .ZN(new_n1940_));
  OAI21_X1   g1891(.A1(new_n1605_), .A2(new_n1248_), .B(new_n1162_), .ZN(new_n1941_));
  AOI22_X1   g1892(.A1(new_n1939_), .A2(new_n1940_), .B1(new_n1941_), .B2(new_n1931_), .ZN(new_n1942_));
  INV_X1     g1893(.I(new_n1937_), .ZN(new_n1943_));
  NOR2_X1    g1894(.A1(new_n1942_), .A2(new_n1943_), .ZN(new_n1944_));
  NOR3_X1    g1895(.A1(new_n1938_), .A2(new_n1944_), .A3(new_n1928_), .ZN(new_n1945_));
  AOI22_X1   g1896(.A1(new_n1925_), .A2(new_n1926_), .B1(new_n1922_), .B2(new_n1923_), .ZN(new_n1946_));
  NAND2_X1   g1897(.A1(new_n1942_), .A2(new_n1943_), .ZN(new_n1947_));
  NAND2_X1   g1898(.A1(new_n1934_), .A2(new_n1937_), .ZN(new_n1948_));
  AOI21_X1   g1899(.A1(new_n1948_), .A2(new_n1947_), .B(new_n1946_), .ZN(new_n1949_));
  NOR2_X1    g1900(.A1(new_n1949_), .A2(new_n1945_), .ZN(new_n1950_));
  AOI21_X1   g1901(.A1(new_n1917_), .A2(new_n1921_), .B(new_n1950_), .ZN(new_n1951_));
  NOR2_X1    g1902(.A1(new_n1889_), .A2(new_n1893_), .ZN(new_n1952_));
  NAND2_X1   g1903(.A1(new_n1903_), .A2(new_n1906_), .ZN(new_n1953_));
  AOI21_X1   g1904(.A1(new_n1953_), .A2(new_n1886_), .B(new_n1952_), .ZN(new_n1954_));
  NAND2_X1   g1905(.A1(new_n1910_), .A2(new_n1912_), .ZN(new_n1955_));
  NOR2_X1    g1906(.A1(new_n1869_), .A2(new_n1885_), .ZN(new_n1956_));
  NOR3_X1    g1907(.A1(new_n1907_), .A2(new_n1956_), .A3(new_n1955_), .ZN(new_n1957_));
  MUX2_X1    g1908(.I0(new_n1345_), .I1(new_n1601_), .S(new_n1288_), .Z(new_n1958_));
  NOR3_X1    g1909(.A1(new_n1032_), .A2(new_n1157_), .A3(new_n1360_), .ZN(new_n1959_));
  NOR3_X1    g1910(.A1(new_n929_), .A2(new_n1096_), .A3(new_n1359_), .ZN(new_n1960_));
  NOR3_X1    g1911(.A1(new_n1605_), .A2(new_n1960_), .A3(new_n1959_), .ZN(new_n1961_));
  NOR2_X1    g1912(.A1(new_n1519_), .A2(new_n1161_), .ZN(new_n1962_));
  NOR2_X1    g1913(.A1(new_n1446_), .A2(new_n842_), .ZN(new_n1963_));
  NOR2_X1    g1914(.A1(new_n1962_), .A2(new_n1963_), .ZN(new_n1964_));
  NOR2_X1    g1915(.A1(new_n1964_), .A2(new_n1157_), .ZN(new_n1965_));
  NOR2_X1    g1916(.A1(new_n1668_), .A2(new_n843_), .ZN(new_n1966_));
  NOR2_X1    g1917(.A1(new_n1965_), .A2(new_n1966_), .ZN(new_n1967_));
  OAI21_X1   g1918(.A1(new_n1958_), .A2(new_n1961_), .B(new_n1967_), .ZN(new_n1968_));
  NAND2_X1   g1919(.A1(new_n1446_), .A2(new_n1288_), .ZN(new_n1969_));
  NAND2_X1   g1920(.A1(new_n1519_), .A2(new_n1162_), .ZN(new_n1970_));
  AOI21_X1   g1921(.A1(new_n1970_), .A2(new_n1969_), .B(new_n1157_), .ZN(new_n1971_));
  NOR2_X1    g1922(.A1(new_n1668_), .A2(new_n1162_), .ZN(new_n1972_));
  NOR2_X1    g1923(.A1(new_n1971_), .A2(new_n1972_), .ZN(new_n1973_));
  NAND2_X1   g1924(.A1(new_n1348_), .A2(new_n1452_), .ZN(new_n1974_));
  NAND3_X1   g1925(.A1(new_n1974_), .A2(new_n1032_), .A3(new_n1133_), .ZN(new_n1975_));
  NOR2_X1    g1926(.A1(new_n1975_), .A2(new_n1973_), .ZN(new_n1976_));
  NOR3_X1    g1927(.A1(new_n1958_), .A2(new_n1967_), .A3(new_n1961_), .ZN(new_n1977_));
  OAI21_X1   g1928(.A1(new_n1976_), .A2(new_n1977_), .B(new_n1968_), .ZN(new_n1978_));
  OAI21_X1   g1929(.A1(new_n1954_), .A2(new_n1957_), .B(new_n1978_), .ZN(new_n1979_));
  NOR2_X1    g1930(.A1(new_n1519_), .A2(new_n1359_), .ZN(new_n1980_));
  NOR2_X1    g1931(.A1(new_n1446_), .A2(new_n1287_), .ZN(new_n1981_));
  OAI21_X1   g1932(.A1(new_n1980_), .A2(new_n1981_), .B(new_n1096_), .ZN(new_n1982_));
  NAND2_X1   g1933(.A1(new_n1523_), .A2(new_n1287_), .ZN(new_n1983_));
  NAND2_X1   g1934(.A1(new_n1519_), .A2(new_n1359_), .ZN(new_n1984_));
  NAND3_X1   g1935(.A1(new_n1984_), .A2(new_n1096_), .A3(new_n1453_), .ZN(new_n1985_));
  NAND3_X1   g1936(.A1(new_n1982_), .A2(new_n1985_), .A3(new_n1983_), .ZN(new_n1986_));
  AOI21_X1   g1937(.A1(new_n1982_), .A2(new_n1983_), .B(new_n1985_), .ZN(new_n1987_));
  NOR2_X1    g1938(.A1(new_n1353_), .A2(new_n1453_), .ZN(new_n1988_));
  OAI21_X1   g1939(.A1(new_n1987_), .A2(new_n1988_), .B(new_n1986_), .ZN(new_n1989_));
  NAND3_X1   g1940(.A1(new_n929_), .A2(new_n1096_), .A3(new_n1452_), .ZN(new_n1990_));
  NAND3_X1   g1941(.A1(new_n1032_), .A2(new_n1157_), .A3(new_n1453_), .ZN(new_n1991_));
  NAND3_X1   g1942(.A1(new_n1353_), .A2(new_n1990_), .A3(new_n1991_), .ZN(new_n1992_));
  XOR2_X1    g1943(.A1(new_n929_), .A2(new_n1359_), .Z(new_n1993_));
  NAND2_X1   g1944(.A1(new_n1993_), .A2(new_n1605_), .ZN(new_n1994_));
  NAND2_X1   g1945(.A1(new_n1994_), .A2(new_n1992_), .ZN(new_n1995_));
  NAND2_X1   g1946(.A1(new_n1989_), .A2(new_n1995_), .ZN(new_n1996_));
  NOR2_X1    g1947(.A1(new_n1890_), .A2(new_n1453_), .ZN(new_n1997_));
  NOR2_X1    g1948(.A1(new_n1997_), .A2(new_n1134_), .ZN(new_n1998_));
  NOR3_X1    g1949(.A1(new_n1998_), .A2(new_n1971_), .A3(new_n1972_), .ZN(new_n1999_));
  OAI22_X1   g1950(.A1(new_n1989_), .A2(new_n1995_), .B1(new_n1999_), .B2(new_n1976_), .ZN(new_n2000_));
  NOR3_X1    g1951(.A1(new_n1219_), .A2(new_n1218_), .A3(new_n1453_), .ZN(new_n2001_));
  AOI21_X1   g1952(.A1(new_n2000_), .A2(new_n1996_), .B(new_n2001_), .ZN(new_n2002_));
  MUX2_X1    g1953(.I0(new_n1806_), .I1(new_n1342_), .S(new_n1288_), .Z(new_n2003_));
  INV_X1     g1954(.I(new_n1961_), .ZN(new_n2004_));
  OAI22_X1   g1955(.A1(new_n1964_), .A2(new_n1157_), .B1(new_n843_), .B2(new_n1668_), .ZN(new_n2005_));
  AOI21_X1   g1956(.A1(new_n2003_), .A2(new_n2004_), .B(new_n2005_), .ZN(new_n2006_));
  OAI21_X1   g1957(.A1(new_n1971_), .A2(new_n1972_), .B(new_n1998_), .ZN(new_n2007_));
  OAI21_X1   g1958(.A1(new_n2006_), .A2(new_n1977_), .B(new_n2007_), .ZN(new_n2008_));
  NAND3_X1   g1959(.A1(new_n2003_), .A2(new_n2004_), .A3(new_n2005_), .ZN(new_n2009_));
  NAND3_X1   g1960(.A1(new_n1968_), .A2(new_n2009_), .A3(new_n1976_), .ZN(new_n2010_));
  NAND2_X1   g1961(.A1(new_n2008_), .A2(new_n2010_), .ZN(new_n2011_));
  NAND3_X1   g1962(.A1(new_n2000_), .A2(new_n1996_), .A3(new_n2001_), .ZN(new_n2012_));
  AOI21_X1   g1963(.A1(new_n2011_), .A2(new_n2012_), .B(new_n2002_), .ZN(new_n2013_));
  NOR3_X1    g1964(.A1(new_n1954_), .A2(new_n1957_), .A3(new_n1978_), .ZN(new_n2014_));
  OAI21_X1   g1965(.A1(new_n2013_), .A2(new_n2014_), .B(new_n1979_), .ZN(new_n2015_));
  NAND3_X1   g1966(.A1(new_n1917_), .A2(new_n1921_), .A3(new_n1950_), .ZN(new_n2016_));
  AOI21_X1   g1967(.A1(new_n2015_), .A2(new_n2016_), .B(new_n1951_), .ZN(new_n2017_));
  AOI21_X1   g1968(.A1(new_n1919_), .A2(new_n1916_), .B(new_n1897_), .ZN(new_n2018_));
  NOR2_X1    g1969(.A1(new_n1311_), .A2(new_n1161_), .ZN(new_n2019_));
  NOR2_X1    g1970(.A1(new_n1547_), .A2(new_n1162_), .ZN(new_n2020_));
  NOR2_X1    g1971(.A1(new_n2019_), .A2(new_n2020_), .ZN(new_n2021_));
  NOR2_X1    g1972(.A1(new_n1316_), .A2(new_n1287_), .ZN(new_n2022_));
  NOR2_X1    g1973(.A1(new_n1679_), .A2(new_n1288_), .ZN(new_n2023_));
  NOR2_X1    g1974(.A1(new_n2023_), .A2(new_n2022_), .ZN(new_n2024_));
  NOR2_X1    g1975(.A1(new_n1601_), .A2(new_n845_), .ZN(new_n2025_));
  NOR2_X1    g1976(.A1(new_n1345_), .A2(new_n846_), .ZN(new_n2026_));
  NOR2_X1    g1977(.A1(new_n2025_), .A2(new_n2026_), .ZN(new_n2027_));
  NOR3_X1    g1978(.A1(new_n1891_), .A2(new_n1890_), .A3(new_n843_), .ZN(new_n2028_));
  AOI21_X1   g1979(.A1(new_n1354_), .A2(new_n843_), .B(new_n2028_), .ZN(new_n2029_));
  NOR4_X1    g1980(.A1(new_n2024_), .A2(new_n2021_), .A3(new_n2027_), .A4(new_n2029_), .ZN(new_n2030_));
  OAI21_X1   g1981(.A1(new_n2030_), .A2(new_n1811_), .B(new_n1820_), .ZN(new_n2031_));
  OAI22_X1   g1982(.A1(new_n2024_), .A2(new_n2021_), .B1(new_n2027_), .B2(new_n2029_), .ZN(new_n2032_));
  NAND2_X1   g1983(.A1(new_n949_), .A2(new_n1360_), .ZN(new_n2033_));
  AOI22_X1   g1984(.A1(new_n1812_), .A2(new_n2033_), .B1(new_n1815_), .B2(new_n1818_), .ZN(new_n2034_));
  NAND3_X1   g1985(.A1(new_n2032_), .A2(new_n2034_), .A3(new_n1821_), .ZN(new_n2035_));
  NAND2_X1   g1986(.A1(new_n2031_), .A2(new_n2035_), .ZN(new_n2036_));
  AOI21_X1   g1987(.A1(new_n1942_), .A2(new_n1943_), .B(new_n1946_), .ZN(new_n2037_));
  NAND2_X1   g1988(.A1(new_n943_), .A2(new_n1452_), .ZN(new_n2038_));
  NOR4_X1    g1989(.A1(new_n939_), .A2(new_n592_), .A3(new_n940_), .A4(new_n1453_), .ZN(new_n2039_));
  OAI21_X1   g1990(.A1(new_n2039_), .A2(new_n2038_), .B(new_n752_), .ZN(new_n2040_));
  AOI21_X1   g1991(.A1(new_n2040_), .A2(new_n1847_), .B(new_n1849_), .ZN(new_n2041_));
  NOR3_X1    g1992(.A1(new_n2037_), .A2(new_n1944_), .A3(new_n2041_), .ZN(new_n2042_));
  NAND2_X1   g1993(.A1(new_n1947_), .A2(new_n1928_), .ZN(new_n2043_));
  INV_X1     g1994(.I(new_n1847_), .ZN(new_n2044_));
  INV_X1     g1995(.I(new_n1849_), .ZN(new_n2045_));
  NAND4_X1   g1996(.A1(new_n943_), .A2(new_n636_), .A3(new_n750_), .A4(new_n1452_), .ZN(new_n2046_));
  AOI21_X1   g1997(.A1(new_n2046_), .A2(new_n1848_), .B(new_n751_), .ZN(new_n2047_));
  OAI21_X1   g1998(.A1(new_n2044_), .A2(new_n2047_), .B(new_n2045_), .ZN(new_n2048_));
  AOI21_X1   g1999(.A1(new_n2043_), .A2(new_n1948_), .B(new_n2048_), .ZN(new_n2049_));
  NOR2_X1    g2000(.A1(new_n2049_), .A2(new_n2042_), .ZN(new_n2050_));
  NOR2_X1    g2001(.A1(new_n2050_), .A2(new_n2036_), .ZN(new_n2051_));
  AOI21_X1   g2002(.A1(new_n2032_), .A2(new_n1821_), .B(new_n2034_), .ZN(new_n2052_));
  NOR3_X1    g2003(.A1(new_n1820_), .A2(new_n2030_), .A3(new_n1811_), .ZN(new_n2053_));
  NOR2_X1    g2004(.A1(new_n2053_), .A2(new_n2052_), .ZN(new_n2054_));
  NOR3_X1    g2005(.A1(new_n2054_), .A2(new_n2042_), .A3(new_n2049_), .ZN(new_n2055_));
  NOR2_X1    g2006(.A1(new_n2051_), .A2(new_n2055_), .ZN(new_n2056_));
  AOI21_X1   g2007(.A1(new_n2017_), .A2(new_n2018_), .B(new_n2056_), .ZN(new_n2057_));
  NOR2_X1    g2008(.A1(new_n2017_), .A2(new_n2018_), .ZN(new_n2058_));
  NOR2_X1    g2009(.A1(new_n2037_), .A2(new_n1944_), .ZN(new_n2059_));
  NOR2_X1    g2010(.A1(new_n2059_), .A2(new_n2041_), .ZN(new_n2060_));
  NAND2_X1   g2011(.A1(new_n2059_), .A2(new_n2041_), .ZN(new_n2061_));
  AOI21_X1   g2012(.A1(new_n2036_), .A2(new_n2061_), .B(new_n2060_), .ZN(new_n2062_));
  INV_X1     g2013(.I(new_n2062_), .ZN(new_n2063_));
  NOR3_X1    g2014(.A1(new_n2057_), .A2(new_n2058_), .A3(new_n2063_), .ZN(new_n2064_));
  NAND2_X1   g2015(.A1(new_n1835_), .A2(new_n1860_), .ZN(new_n2065_));
  XOR2_X1    g2016(.A1(new_n2065_), .A2(new_n1857_), .Z(new_n2066_));
  OAI21_X1   g2017(.A1(new_n2057_), .A2(new_n2058_), .B(new_n2063_), .ZN(new_n2067_));
  OAI21_X1   g2018(.A1(new_n2064_), .A2(new_n2066_), .B(new_n2067_), .ZN(new_n2068_));
  NAND2_X1   g2019(.A1(new_n2068_), .A2(new_n1862_), .ZN(new_n2069_));
  XOR2_X1    g2020(.A1(new_n1721_), .A2(new_n1726_), .Z(new_n2070_));
  XNOR2_X1   g2021(.A1(new_n2070_), .A2(new_n1731_), .ZN(new_n2071_));
  AOI21_X1   g2022(.A1(new_n1854_), .A2(new_n1850_), .B(new_n1852_), .ZN(new_n2072_));
  INV_X1     g2023(.I(new_n2072_), .ZN(new_n2073_));
  NAND2_X1   g2024(.A1(new_n2071_), .A2(new_n2073_), .ZN(new_n2074_));
  XOR2_X1    g2025(.A1(new_n2070_), .A2(new_n1731_), .Z(new_n2075_));
  NAND2_X1   g2026(.A1(new_n2075_), .A2(new_n2072_), .ZN(new_n2076_));
  NAND2_X1   g2027(.A1(new_n1781_), .A2(new_n1773_), .ZN(new_n2077_));
  INV_X1     g2028(.I(new_n2077_), .ZN(new_n2078_));
  NAND2_X1   g2029(.A1(new_n2078_), .A2(new_n1779_), .ZN(new_n2079_));
  NAND2_X1   g2030(.A1(new_n2077_), .A2(new_n1780_), .ZN(new_n2080_));
  NAND4_X1   g2031(.A1(new_n2079_), .A2(new_n2074_), .A3(new_n2076_), .A4(new_n2080_), .ZN(new_n2081_));
  NOR2_X1    g2032(.A1(new_n2075_), .A2(new_n2072_), .ZN(new_n2082_));
  NOR2_X1    g2033(.A1(new_n2071_), .A2(new_n2073_), .ZN(new_n2083_));
  NOR2_X1    g2034(.A1(new_n2077_), .A2(new_n1780_), .ZN(new_n2084_));
  NOR2_X1    g2035(.A1(new_n2078_), .A2(new_n1779_), .ZN(new_n2085_));
  OAI22_X1   g2036(.A1(new_n2085_), .A2(new_n2084_), .B1(new_n2083_), .B2(new_n2082_), .ZN(new_n2086_));
  NAND2_X1   g2037(.A1(new_n2086_), .A2(new_n2081_), .ZN(new_n2087_));
  OAI21_X1   g2038(.A1(new_n2068_), .A2(new_n1862_), .B(new_n2087_), .ZN(new_n2088_));
  NAND2_X1   g2039(.A1(new_n2079_), .A2(new_n2080_), .ZN(new_n2089_));
  AOI21_X1   g2040(.A1(new_n2089_), .A2(new_n2076_), .B(new_n2082_), .ZN(new_n2090_));
  AOI21_X1   g2041(.A1(new_n2088_), .A2(new_n2069_), .B(new_n2090_), .ZN(new_n2091_));
  NAND3_X1   g2042(.A1(new_n2088_), .A2(new_n2069_), .A3(new_n2090_), .ZN(new_n2092_));
  NAND2_X1   g2043(.A1(new_n1794_), .A2(new_n1735_), .ZN(new_n2093_));
  NAND2_X1   g2044(.A1(new_n1791_), .A2(new_n1734_), .ZN(new_n2094_));
  NAND2_X1   g2045(.A1(new_n2094_), .A2(new_n2093_), .ZN(new_n2095_));
  NAND2_X1   g2046(.A1(new_n1787_), .A2(new_n1788_), .ZN(new_n2096_));
  NAND2_X1   g2047(.A1(new_n2095_), .A2(new_n2096_), .ZN(new_n2097_));
  NAND4_X1   g2048(.A1(new_n2094_), .A2(new_n2093_), .A3(new_n1787_), .A4(new_n1788_), .ZN(new_n2098_));
  NAND2_X1   g2049(.A1(new_n2097_), .A2(new_n2098_), .ZN(new_n2099_));
  AOI21_X1   g2050(.A1(new_n2092_), .A2(new_n2099_), .B(new_n2091_), .ZN(new_n2100_));
  NAND3_X1   g2051(.A1(new_n1753_), .A2(new_n1797_), .A3(new_n1755_), .ZN(new_n2101_));
  AOI21_X1   g2052(.A1(new_n2100_), .A2(new_n2101_), .B(new_n1798_), .ZN(new_n2102_));
  OAI21_X1   g2053(.A1(new_n1737_), .A2(new_n1754_), .B(new_n1752_), .ZN(new_n2103_));
  NOR3_X1    g2054(.A1(new_n1641_), .A2(new_n1746_), .A3(new_n1692_), .ZN(new_n2104_));
  AOI21_X1   g2055(.A1(new_n1744_), .A2(new_n1693_), .B(new_n1691_), .ZN(new_n2105_));
  OAI21_X1   g2056(.A1(new_n2104_), .A2(new_n2105_), .B(new_n2103_), .ZN(new_n2106_));
  NAND2_X1   g2057(.A1(new_n2106_), .A2(new_n1748_), .ZN(new_n2107_));
  OAI21_X1   g2058(.A1(new_n2102_), .A2(new_n2107_), .B(new_n1748_), .ZN(new_n2108_));
  INV_X1     g2059(.I(new_n1623_), .ZN(new_n2109_));
  NOR2_X1    g2060(.A1(new_n2109_), .A2(new_n1624_), .ZN(new_n2110_));
  XOR2_X1    g2061(.A1(new_n1626_), .A2(new_n2110_), .Z(new_n2111_));
  AOI21_X1   g2062(.A1(new_n2108_), .A2(new_n1694_), .B(new_n2111_), .ZN(new_n2112_));
  NOR3_X1    g2063(.A1(new_n2104_), .A2(new_n2105_), .A3(new_n2103_), .ZN(new_n2113_));
  INV_X1     g2064(.I(new_n1798_), .ZN(new_n2114_));
  AOI21_X1   g2065(.A1(new_n1918_), .A2(new_n1919_), .B(new_n1920_), .ZN(new_n2115_));
  NOR3_X1    g2066(.A1(new_n1914_), .A2(new_n1897_), .A3(new_n1916_), .ZN(new_n2116_));
  NAND3_X1   g2067(.A1(new_n1948_), .A2(new_n1947_), .A3(new_n1946_), .ZN(new_n2117_));
  OAI21_X1   g2068(.A1(new_n1938_), .A2(new_n1944_), .B(new_n1928_), .ZN(new_n2118_));
  NAND2_X1   g2069(.A1(new_n2118_), .A2(new_n2117_), .ZN(new_n2119_));
  OAI21_X1   g2070(.A1(new_n2116_), .A2(new_n2115_), .B(new_n2119_), .ZN(new_n2120_));
  OAI21_X1   g2071(.A1(new_n1907_), .A2(new_n1956_), .B(new_n1955_), .ZN(new_n2121_));
  NAND3_X1   g2072(.A1(new_n1953_), .A2(new_n1886_), .A3(new_n1952_), .ZN(new_n2122_));
  AOI21_X1   g2073(.A1(new_n2007_), .A2(new_n2009_), .B(new_n2006_), .ZN(new_n2123_));
  AOI21_X1   g2074(.A1(new_n2121_), .A2(new_n2122_), .B(new_n2123_), .ZN(new_n2124_));
  NAND2_X1   g2075(.A1(new_n1446_), .A2(new_n1360_), .ZN(new_n2125_));
  NAND2_X1   g2076(.A1(new_n1519_), .A2(new_n1288_), .ZN(new_n2126_));
  AOI21_X1   g2077(.A1(new_n2126_), .A2(new_n2125_), .B(new_n1157_), .ZN(new_n2127_));
  NOR2_X1    g2078(.A1(new_n1668_), .A2(new_n1288_), .ZN(new_n2128_));
  OAI21_X1   g2079(.A1(new_n1446_), .A2(new_n1360_), .B(new_n1453_), .ZN(new_n2129_));
  NOR2_X1    g2080(.A1(new_n2129_), .A2(new_n1157_), .ZN(new_n2130_));
  NOR3_X1    g2081(.A1(new_n2127_), .A2(new_n2130_), .A3(new_n2128_), .ZN(new_n2131_));
  OAI21_X1   g2082(.A1(new_n2127_), .A2(new_n2128_), .B(new_n2130_), .ZN(new_n2132_));
  NAND2_X1   g2083(.A1(new_n1605_), .A2(new_n1452_), .ZN(new_n2133_));
  AOI21_X1   g2084(.A1(new_n2132_), .A2(new_n2133_), .B(new_n2131_), .ZN(new_n2134_));
  AND3_X2    g2085(.A1(new_n1344_), .A2(new_n1990_), .A3(new_n1343_), .Z(new_n2135_));
  AOI22_X1   g2086(.A1(new_n2135_), .A2(new_n1991_), .B1(new_n1605_), .B2(new_n1993_), .ZN(new_n2136_));
  NOR2_X1    g2087(.A1(new_n2134_), .A2(new_n2136_), .ZN(new_n2137_));
  NAND2_X1   g2088(.A1(new_n1975_), .A2(new_n1973_), .ZN(new_n2138_));
  AOI22_X1   g2089(.A1(new_n2134_), .A2(new_n2136_), .B1(new_n2007_), .B2(new_n2138_), .ZN(new_n2139_));
  INV_X1     g2090(.I(new_n2001_), .ZN(new_n2140_));
  OAI21_X1   g2091(.A1(new_n2139_), .A2(new_n2137_), .B(new_n2140_), .ZN(new_n2141_));
  AOI21_X1   g2092(.A1(new_n1968_), .A2(new_n2009_), .B(new_n1976_), .ZN(new_n2142_));
  NOR3_X1    g2093(.A1(new_n2006_), .A2(new_n1977_), .A3(new_n2007_), .ZN(new_n2143_));
  NOR2_X1    g2094(.A1(new_n2143_), .A2(new_n2142_), .ZN(new_n2144_));
  NOR3_X1    g2095(.A1(new_n2139_), .A2(new_n2137_), .A3(new_n2140_), .ZN(new_n2145_));
  OAI21_X1   g2096(.A1(new_n2144_), .A2(new_n2145_), .B(new_n2141_), .ZN(new_n2146_));
  NAND3_X1   g2097(.A1(new_n2121_), .A2(new_n2122_), .A3(new_n2123_), .ZN(new_n2147_));
  AOI21_X1   g2098(.A1(new_n2146_), .A2(new_n2147_), .B(new_n2124_), .ZN(new_n2148_));
  NOR3_X1    g2099(.A1(new_n2116_), .A2(new_n2115_), .A3(new_n2119_), .ZN(new_n2149_));
  OAI21_X1   g2100(.A1(new_n2148_), .A2(new_n2149_), .B(new_n2120_), .ZN(new_n2150_));
  INV_X1     g2101(.I(new_n2018_), .ZN(new_n2151_));
  OAI21_X1   g2102(.A1(new_n2042_), .A2(new_n2049_), .B(new_n2054_), .ZN(new_n2152_));
  NAND2_X1   g2103(.A1(new_n2050_), .A2(new_n2036_), .ZN(new_n2153_));
  NAND2_X1   g2104(.A1(new_n2152_), .A2(new_n2153_), .ZN(new_n2154_));
  OAI21_X1   g2105(.A1(new_n2150_), .A2(new_n2151_), .B(new_n2154_), .ZN(new_n2155_));
  NAND2_X1   g2106(.A1(new_n2150_), .A2(new_n2151_), .ZN(new_n2156_));
  NAND3_X1   g2107(.A1(new_n2155_), .A2(new_n2156_), .A3(new_n2062_), .ZN(new_n2157_));
  NAND2_X1   g2108(.A1(new_n2065_), .A2(new_n1857_), .ZN(new_n2158_));
  NAND3_X1   g2109(.A1(new_n1855_), .A2(new_n1854_), .A3(new_n1850_), .ZN(new_n2159_));
  OAI21_X1   g2110(.A1(new_n1851_), .A2(new_n1852_), .B(new_n1837_), .ZN(new_n2160_));
  NAND2_X1   g2111(.A1(new_n2160_), .A2(new_n2159_), .ZN(new_n2161_));
  NAND3_X1   g2112(.A1(new_n2161_), .A2(new_n1835_), .A3(new_n1860_), .ZN(new_n2162_));
  NAND2_X1   g2113(.A1(new_n2158_), .A2(new_n2162_), .ZN(new_n2163_));
  NAND2_X1   g2114(.A1(new_n2157_), .A2(new_n2163_), .ZN(new_n2164_));
  AOI21_X1   g2115(.A1(new_n2164_), .A2(new_n2067_), .B(new_n1861_), .ZN(new_n2165_));
  AOI21_X1   g2116(.A1(new_n2155_), .A2(new_n2156_), .B(new_n2062_), .ZN(new_n2166_));
  AOI21_X1   g2117(.A1(new_n2157_), .A2(new_n2163_), .B(new_n2166_), .ZN(new_n2167_));
  NOR4_X1    g2118(.A1(new_n2085_), .A2(new_n2083_), .A3(new_n2082_), .A4(new_n2084_), .ZN(new_n2168_));
  AOI22_X1   g2119(.A1(new_n2079_), .A2(new_n2080_), .B1(new_n2074_), .B2(new_n2076_), .ZN(new_n2169_));
  NOR2_X1    g2120(.A1(new_n2169_), .A2(new_n2168_), .ZN(new_n2170_));
  AOI21_X1   g2121(.A1(new_n2167_), .A2(new_n1861_), .B(new_n2170_), .ZN(new_n2171_));
  INV_X1     g2122(.I(new_n2090_), .ZN(new_n2172_));
  OAI21_X1   g2123(.A1(new_n2171_), .A2(new_n2165_), .B(new_n2172_), .ZN(new_n2173_));
  NAND2_X1   g2124(.A1(new_n2092_), .A2(new_n2099_), .ZN(new_n2174_));
  NAND3_X1   g2125(.A1(new_n2174_), .A2(new_n2173_), .A3(new_n2101_), .ZN(new_n2175_));
  AOI21_X1   g2126(.A1(new_n2175_), .A2(new_n2114_), .B(new_n2107_), .ZN(new_n2176_));
  NOR3_X1    g2127(.A1(new_n2176_), .A2(new_n1694_), .A3(new_n2113_), .ZN(new_n2177_));
  INV_X1     g2128(.I(new_n1627_), .ZN(new_n2178_));
  INV_X1     g2129(.I(new_n1629_), .ZN(new_n2179_));
  NAND3_X1   g2130(.A1(new_n1628_), .A2(new_n1576_), .A3(new_n1580_), .ZN(new_n2180_));
  AOI21_X1   g2131(.A1(new_n2179_), .A2(new_n2180_), .B(new_n2178_), .ZN(new_n2181_));
  NOR3_X1    g2132(.A1(new_n2112_), .A2(new_n2177_), .A3(new_n2181_), .ZN(new_n2182_));
  OAI21_X1   g2133(.A1(new_n2182_), .A2(new_n1632_), .B(new_n1592_), .ZN(new_n2183_));
  INV_X1     g2134(.I(new_n1583_), .ZN(new_n2184_));
  XOR2_X1    g2135(.A1(new_n1490_), .A2(new_n1586_), .Z(new_n2185_));
  NOR2_X1    g2136(.A1(new_n2185_), .A2(new_n2184_), .ZN(new_n2186_));
  INV_X1     g2137(.I(new_n2186_), .ZN(new_n2187_));
  NAND3_X1   g2138(.A1(new_n2183_), .A2(new_n1497_), .A3(new_n2187_), .ZN(new_n2188_));
  NAND3_X1   g2139(.A1(new_n2188_), .A2(new_n1398_), .A3(new_n1494_), .ZN(new_n2189_));
  AOI21_X1   g2140(.A1(new_n2189_), .A2(new_n1397_), .B(new_n1243_), .ZN(new_n2190_));
  OAI21_X1   g2141(.A1(new_n2190_), .A2(new_n1240_), .B(new_n1191_), .ZN(new_n2191_));
  NAND2_X1   g2142(.A1(new_n2191_), .A2(new_n1188_), .ZN(new_n2192_));
  INV_X1     g2143(.I(new_n1243_), .ZN(new_n2193_));
  INV_X1     g2144(.I(new_n1398_), .ZN(new_n2194_));
  AOI21_X1   g2145(.A1(new_n1495_), .A2(new_n1496_), .B(new_n1492_), .ZN(new_n2195_));
  NOR3_X1    g2146(.A1(new_n1406_), .A2(new_n1403_), .A3(new_n1493_), .ZN(new_n2196_));
  NOR3_X1    g2147(.A1(new_n1588_), .A2(new_n1589_), .A3(new_n1590_), .ZN(new_n2197_));
  AOI21_X1   g2148(.A1(new_n1582_), .A2(new_n1584_), .B(new_n1586_), .ZN(new_n2198_));
  NOR2_X1    g2149(.A1(new_n2198_), .A2(new_n2197_), .ZN(new_n2199_));
  INV_X1     g2150(.I(new_n1632_), .ZN(new_n2200_));
  INV_X1     g2151(.I(new_n1694_), .ZN(new_n2201_));
  NOR3_X1    g2152(.A1(new_n2171_), .A2(new_n2165_), .A3(new_n2172_), .ZN(new_n2202_));
  AOI22_X1   g2153(.A1(new_n2094_), .A2(new_n2093_), .B1(new_n1787_), .B2(new_n1788_), .ZN(new_n2203_));
  NOR3_X1    g2154(.A1(new_n2096_), .A2(new_n1792_), .A3(new_n1795_), .ZN(new_n2204_));
  NOR2_X1    g2155(.A1(new_n2203_), .A2(new_n2204_), .ZN(new_n2205_));
  OAI21_X1   g2156(.A1(new_n2202_), .A2(new_n2205_), .B(new_n2173_), .ZN(new_n2206_));
  NOR3_X1    g2157(.A1(new_n1754_), .A2(new_n1711_), .A3(new_n1737_), .ZN(new_n2207_));
  INV_X1     g2158(.I(new_n1755_), .ZN(new_n2208_));
  AOI21_X1   g2159(.A1(new_n2095_), .A2(new_n1788_), .B(new_n1786_), .ZN(new_n2209_));
  NOR3_X1    g2160(.A1(new_n2208_), .A2(new_n2209_), .A3(new_n2207_), .ZN(new_n2210_));
  OAI21_X1   g2161(.A1(new_n2206_), .A2(new_n2210_), .B(new_n2114_), .ZN(new_n2211_));
  AOI21_X1   g2162(.A1(new_n1747_), .A2(new_n1745_), .B(new_n1740_), .ZN(new_n2212_));
  NOR2_X1    g2163(.A1(new_n2113_), .A2(new_n2212_), .ZN(new_n2213_));
  AOI21_X1   g2164(.A1(new_n2211_), .A2(new_n2213_), .B(new_n2113_), .ZN(new_n2214_));
  XNOR2_X1   g2165(.A1(new_n1626_), .A2(new_n2110_), .ZN(new_n2215_));
  OAI21_X1   g2166(.A1(new_n2214_), .A2(new_n2201_), .B(new_n2215_), .ZN(new_n2216_));
  NAND3_X1   g2167(.A1(new_n2164_), .A2(new_n1861_), .A3(new_n2067_), .ZN(new_n2217_));
  AOI21_X1   g2168(.A1(new_n2217_), .A2(new_n2087_), .B(new_n2165_), .ZN(new_n2218_));
  AOI21_X1   g2169(.A1(new_n2218_), .A2(new_n2090_), .B(new_n2205_), .ZN(new_n2219_));
  NOR3_X1    g2170(.A1(new_n2219_), .A2(new_n2091_), .A3(new_n2210_), .ZN(new_n2220_));
  OAI21_X1   g2171(.A1(new_n2220_), .A2(new_n1798_), .B(new_n2213_), .ZN(new_n2221_));
  NAND3_X1   g2172(.A1(new_n2221_), .A2(new_n2201_), .A3(new_n1748_), .ZN(new_n2222_));
  OAI21_X1   g2173(.A1(new_n1631_), .A2(new_n1629_), .B(new_n1627_), .ZN(new_n2223_));
  NAND3_X1   g2174(.A1(new_n2216_), .A2(new_n2222_), .A3(new_n2223_), .ZN(new_n2224_));
  AOI21_X1   g2175(.A1(new_n2224_), .A2(new_n2200_), .B(new_n2199_), .ZN(new_n2225_));
  NOR3_X1    g2176(.A1(new_n2225_), .A2(new_n2196_), .A3(new_n2186_), .ZN(new_n2226_));
  NOR3_X1    g2177(.A1(new_n2226_), .A2(new_n2194_), .A3(new_n2195_), .ZN(new_n2227_));
  OAI21_X1   g2178(.A1(new_n2227_), .A2(new_n1396_), .B(new_n2193_), .ZN(new_n2228_));
  NAND3_X1   g2179(.A1(new_n2228_), .A2(new_n1190_), .A3(new_n1241_), .ZN(new_n2229_));
  NOR2_X1    g2180(.A1(new_n964_), .A2(new_n967_), .ZN(new_n2230_));
  INV_X1     g2181(.I(new_n2230_), .ZN(new_n2231_));
  NAND3_X1   g2182(.A1(new_n2192_), .A2(new_n2229_), .A3(new_n2231_), .ZN(new_n2232_));
  AOI21_X1   g2183(.A1(new_n2232_), .A2(new_n970_), .B(new_n827_), .ZN(new_n2233_));
  INV_X1     g2184(.I(new_n826_), .ZN(new_n2234_));
  NAND2_X1   g2185(.A1(new_n824_), .A2(new_n2234_), .ZN(new_n2235_));
  INV_X1     g2186(.I(new_n2235_), .ZN(new_n2236_));
  NOR3_X1    g2187(.A1(new_n2233_), .A2(new_n657_), .A3(new_n2236_), .ZN(new_n2237_));
  OAI21_X1   g2188(.A1(new_n2237_), .A2(new_n655_), .B(new_n612_), .ZN(new_n2238_));
  INV_X1     g2189(.I(new_n612_), .ZN(new_n2239_));
  INV_X1     g2190(.I(new_n655_), .ZN(new_n2240_));
  INV_X1     g2191(.I(new_n827_), .ZN(new_n2241_));
  AOI21_X1   g2192(.A1(new_n2228_), .A2(new_n1241_), .B(new_n1190_), .ZN(new_n2242_));
  NOR2_X1    g2193(.A1(new_n2242_), .A2(new_n1187_), .ZN(new_n2243_));
  NOR3_X1    g2194(.A1(new_n2190_), .A2(new_n1191_), .A3(new_n1240_), .ZN(new_n2244_));
  NOR3_X1    g2195(.A1(new_n2243_), .A2(new_n2244_), .A3(new_n2230_), .ZN(new_n2245_));
  OAI21_X1   g2196(.A1(new_n2245_), .A2(new_n969_), .B(new_n2241_), .ZN(new_n2246_));
  NAND3_X1   g2197(.A1(new_n2246_), .A2(new_n656_), .A3(new_n2235_), .ZN(new_n2247_));
  NAND3_X1   g2198(.A1(new_n2247_), .A2(new_n2239_), .A3(new_n2240_), .ZN(new_n2248_));
  INV_X1     g2199(.I(new_n559_), .ZN(new_n2249_));
  INV_X1     g2200(.I(new_n1100_), .ZN(new_n2250_));
  NOR4_X1    g2201(.A1(new_n168_), .A2(new_n253_), .A3(new_n330_), .A4(new_n285_), .ZN(new_n2251_));
  NOR2_X1    g2202(.A1(new_n139_), .A2(new_n269_), .ZN(new_n2252_));
  INV_X1     g2203(.I(new_n2252_), .ZN(new_n2253_));
  NOR3_X1    g2204(.A1(new_n2253_), .A2(new_n210_), .A3(new_n271_), .ZN(new_n2254_));
  INV_X1     g2205(.I(new_n2254_), .ZN(new_n2255_));
  NOR2_X1    g2206(.A1(new_n2255_), .A2(new_n527_), .ZN(new_n2256_));
  NAND4_X1   g2207(.A1(new_n2256_), .A2(new_n2250_), .A3(new_n2249_), .A4(new_n2251_), .ZN(new_n2257_));
  OR3_X2     g2208(.A1(new_n2257_), .A2(new_n245_), .A3(new_n567_), .Z(new_n2258_));
  NOR2_X1    g2209(.A1(new_n164_), .A2(new_n332_), .ZN(new_n2259_));
  NAND4_X1   g2210(.A1(new_n2259_), .A2(new_n743_), .A3(new_n300_), .A4(new_n351_), .ZN(new_n2260_));
  NOR2_X1    g2211(.A1(new_n691_), .A2(new_n722_), .ZN(new_n2261_));
  NOR2_X1    g2212(.A1(new_n312_), .A2(new_n156_), .ZN(new_n2262_));
  INV_X1     g2213(.I(new_n508_), .ZN(new_n2263_));
  NOR4_X1    g2214(.A1(new_n2263_), .A2(new_n1120_), .A3(new_n413_), .A4(new_n718_), .ZN(new_n2264_));
  NAND4_X1   g2215(.A1(new_n2264_), .A2(new_n887_), .A3(new_n2261_), .A4(new_n2262_), .ZN(new_n2265_));
  NOR3_X1    g2216(.A1(new_n267_), .A2(new_n202_), .A3(new_n272_), .ZN(new_n2266_));
  NAND4_X1   g2217(.A1(new_n2266_), .A2(new_n849_), .A3(new_n1271_), .A4(new_n386_), .ZN(new_n2267_));
  OR3_X2     g2218(.A1(new_n2265_), .A2(new_n2260_), .A3(new_n2267_), .Z(new_n2268_));
  NOR4_X1    g2219(.A1(new_n2258_), .A2(new_n1018_), .A3(new_n1138_), .A4(new_n2268_), .ZN(new_n2269_));
  INV_X1     g2220(.I(new_n2269_), .ZN(new_n2270_));
  AOI21_X1   g2221(.A1(new_n2248_), .A2(new_n2238_), .B(new_n2270_), .ZN(new_n2271_));
  NOR2_X1    g2222(.A1(new_n249_), .A2(new_n126_), .ZN(new_n2272_));
  INV_X1     g2223(.I(new_n2272_), .ZN(new_n2273_));
  NOR4_X1    g2224(.A1(new_n254_), .A2(new_n437_), .A3(new_n580_), .A4(new_n536_), .ZN(new_n2274_));
  NAND4_X1   g2225(.A1(new_n2274_), .A2(new_n679_), .A3(new_n563_), .A4(new_n2273_), .ZN(new_n2275_));
  NOR4_X1    g2226(.A1(new_n313_), .A2(new_n201_), .A3(new_n296_), .A4(new_n450_), .ZN(new_n2276_));
  NOR2_X1    g2227(.A1(new_n193_), .A2(new_n265_), .ZN(new_n2277_));
  NAND4_X1   g2228(.A1(new_n2277_), .A2(new_n512_), .A3(new_n275_), .A4(new_n447_), .ZN(new_n2278_));
  INV_X1     g2229(.I(new_n2278_), .ZN(new_n2279_));
  NOR3_X1    g2230(.A1(new_n552_), .A2(new_n736_), .A3(new_n327_), .ZN(new_n2280_));
  NAND4_X1   g2231(.A1(new_n2279_), .A2(new_n1249_), .A3(new_n2276_), .A4(new_n2280_), .ZN(new_n2281_));
  INV_X1     g2232(.I(new_n731_), .ZN(new_n2282_));
  NOR3_X1    g2233(.A1(new_n241_), .A2(new_n729_), .A3(new_n435_), .ZN(new_n2283_));
  NOR3_X1    g2234(.A1(new_n974_), .A2(new_n304_), .A3(new_n735_), .ZN(new_n2284_));
  NOR4_X1    g2235(.A1(new_n505_), .A2(new_n360_), .A3(new_n381_), .A4(new_n695_), .ZN(new_n2285_));
  AND3_X2    g2236(.A1(new_n2284_), .A2(new_n2283_), .A3(new_n2285_), .Z(new_n2286_));
  NAND4_X1   g2237(.A1(new_n2286_), .A2(new_n565_), .A3(new_n574_), .A4(new_n2282_), .ZN(new_n2287_));
  NOR4_X1    g2238(.A1(new_n210_), .A2(new_n272_), .A3(new_n426_), .A4(new_n561_), .ZN(new_n2288_));
  NOR3_X1    g2239(.A1(new_n345_), .A2(new_n156_), .A3(new_n919_), .ZN(new_n2289_));
  NOR2_X1    g2240(.A1(new_n109_), .A2(new_n126_), .ZN(new_n2290_));
  NOR3_X1    g2241(.A1(new_n185_), .A2(new_n188_), .A3(new_n2290_), .ZN(new_n2291_));
  NAND4_X1   g2242(.A1(new_n2291_), .A2(new_n322_), .A3(new_n1266_), .A4(new_n699_), .ZN(new_n2292_));
  INV_X1     g2243(.I(new_n2292_), .ZN(new_n2293_));
  NAND4_X1   g2244(.A1(new_n2293_), .A2(new_n707_), .A3(new_n2288_), .A4(new_n2289_), .ZN(new_n2294_));
  NOR4_X1    g2245(.A1(new_n2287_), .A2(new_n2275_), .A3(new_n2281_), .A4(new_n2294_), .ZN(new_n2295_));
  NOR2_X1    g2246(.A1(new_n657_), .A2(new_n655_), .ZN(new_n2296_));
  OAI21_X1   g2247(.A1(new_n2233_), .A2(new_n2236_), .B(new_n2296_), .ZN(new_n2297_));
  INV_X1     g2248(.I(new_n2296_), .ZN(new_n2298_));
  NAND3_X1   g2249(.A1(new_n2246_), .A2(new_n2235_), .A3(new_n2298_), .ZN(new_n2299_));
  AOI21_X1   g2250(.A1(new_n2299_), .A2(new_n2297_), .B(new_n2295_), .ZN(new_n2300_));
  OAI21_X1   g2251(.A1(new_n2245_), .A2(new_n969_), .B(new_n827_), .ZN(new_n2301_));
  NAND3_X1   g2252(.A1(new_n2232_), .A2(new_n2241_), .A3(new_n970_), .ZN(new_n2302_));
  INV_X1     g2253(.I(new_n493_), .ZN(new_n2303_));
  NOR3_X1    g2254(.A1(new_n448_), .A2(new_n536_), .A3(new_n695_), .ZN(new_n2304_));
  NAND4_X1   g2255(.A1(new_n680_), .A2(new_n2304_), .A3(new_n737_), .A4(new_n1016_), .ZN(new_n2305_));
  NOR3_X1    g2256(.A1(new_n387_), .A2(new_n569_), .A3(new_n587_), .ZN(new_n2306_));
  INV_X1     g2257(.I(new_n2306_), .ZN(new_n2307_));
  NOR4_X1    g2258(.A1(new_n2305_), .A2(new_n876_), .A3(new_n2307_), .A4(new_n2303_), .ZN(new_n2308_));
  NAND4_X1   g2259(.A1(new_n2308_), .A2(new_n533_), .A3(new_n973_), .A4(new_n1083_), .ZN(new_n2309_));
  AOI21_X1   g2260(.A1(new_n2301_), .A2(new_n2302_), .B(new_n2309_), .ZN(new_n2310_));
  NOR2_X1    g2261(.A1(new_n969_), .A2(new_n2230_), .ZN(new_n2311_));
  OAI21_X1   g2262(.A1(new_n2243_), .A2(new_n2244_), .B(new_n2311_), .ZN(new_n2312_));
  INV_X1     g2263(.I(new_n2311_), .ZN(new_n2313_));
  NAND3_X1   g2264(.A1(new_n2192_), .A2(new_n2229_), .A3(new_n2313_), .ZN(new_n2314_));
  NAND2_X1   g2265(.A1(new_n2312_), .A2(new_n2314_), .ZN(new_n2315_));
  INV_X1     g2266(.I(new_n547_), .ZN(new_n2316_));
  INV_X1     g2267(.I(new_n567_), .ZN(new_n2317_));
  NAND4_X1   g2268(.A1(new_n2316_), .A2(new_n486_), .A3(new_n278_), .A4(new_n2317_), .ZN(new_n2318_));
  NOR3_X1    g2269(.A1(new_n723_), .A2(new_n310_), .A3(new_n494_), .ZN(new_n2319_));
  NOR3_X1    g2270(.A1(new_n261_), .A2(new_n159_), .A3(new_n745_), .ZN(new_n2320_));
  NOR2_X1    g2271(.A1(new_n250_), .A2(new_n1015_), .ZN(new_n2321_));
  NAND4_X1   g2272(.A1(new_n2320_), .A2(new_n2319_), .A3(new_n351_), .A4(new_n2321_), .ZN(new_n2322_));
  NOR2_X1    g2273(.A1(new_n452_), .A2(new_n382_), .ZN(new_n2323_));
  INV_X1     g2274(.I(new_n2323_), .ZN(new_n2324_));
  NOR4_X1    g2275(.A1(new_n559_), .A2(new_n2303_), .A3(new_n1069_), .A4(new_n2324_), .ZN(new_n2325_));
  NOR2_X1    g2276(.A1(new_n262_), .A2(new_n346_), .ZN(new_n2326_));
  AND4_X2    g2277(.A1(new_n293_), .A2(new_n2266_), .A3(new_n451_), .A4(new_n2326_), .Z(new_n2327_));
  NAND4_X1   g2278(.A1(new_n2325_), .A2(new_n2283_), .A3(new_n2327_), .A4(new_n2289_), .ZN(new_n2328_));
  NOR2_X1    g2279(.A1(new_n110_), .A2(new_n356_), .ZN(new_n2329_));
  INV_X1     g2280(.I(new_n2329_), .ZN(new_n2330_));
  NOR2_X1    g2281(.A1(new_n2330_), .A2(new_n208_), .ZN(new_n2331_));
  INV_X1     g2282(.I(new_n401_), .ZN(new_n2332_));
  NOR3_X1    g2283(.A1(new_n854_), .A2(new_n265_), .A3(new_n573_), .ZN(new_n2333_));
  NAND4_X1   g2284(.A1(new_n2333_), .A2(new_n563_), .A3(new_n1012_), .A4(new_n2332_), .ZN(new_n2334_));
  NOR2_X1    g2285(.A1(new_n2334_), .A2(new_n542_), .ZN(new_n2335_));
  NAND4_X1   g2286(.A1(new_n2335_), .A2(new_n506_), .A3(new_n685_), .A4(new_n2331_), .ZN(new_n2336_));
  NOR4_X1    g2287(.A1(new_n2336_), .A2(new_n2328_), .A3(new_n2318_), .A4(new_n2322_), .ZN(new_n2337_));
  INV_X1     g2288(.I(new_n2275_), .ZN(new_n2338_));
  NOR4_X1    g2289(.A1(new_n210_), .A2(new_n454_), .A3(new_n396_), .A4(new_n509_), .ZN(new_n2339_));
  NOR4_X1    g2290(.A1(new_n164_), .A2(new_n177_), .A3(new_n361_), .A4(new_n299_), .ZN(new_n2340_));
  NAND4_X1   g2291(.A1(new_n2339_), .A2(new_n318_), .A3(new_n2320_), .A4(new_n2340_), .ZN(new_n2341_));
  INV_X1     g2292(.I(new_n2341_), .ZN(new_n2342_));
  NOR4_X1    g2293(.A1(new_n2328_), .A2(new_n185_), .A3(new_n2290_), .A4(new_n389_), .ZN(new_n2343_));
  INV_X1     g2294(.I(new_n247_), .ZN(new_n2344_));
  NOR3_X1    g2295(.A1(new_n256_), .A2(new_n854_), .A3(new_n587_), .ZN(new_n2345_));
  INV_X1     g2296(.I(new_n2345_), .ZN(new_n2346_));
  NOR2_X1    g2297(.A1(new_n200_), .A2(new_n545_), .ZN(new_n2347_));
  NAND2_X1   g2298(.A1(new_n2347_), .A2(new_n909_), .ZN(new_n2348_));
  NAND4_X1   g2299(.A1(new_n887_), .A2(new_n1111_), .A3(new_n1073_), .A4(new_n871_), .ZN(new_n2349_));
  NOR4_X1    g2300(.A1(new_n2346_), .A2(new_n2348_), .A3(new_n2349_), .A4(new_n2344_), .ZN(new_n2350_));
  NAND4_X1   g2301(.A1(new_n2343_), .A2(new_n2338_), .A3(new_n2342_), .A4(new_n2350_), .ZN(new_n2351_));
  INV_X1     g2302(.I(new_n2351_), .ZN(new_n2352_));
  NAND3_X1   g2303(.A1(new_n2229_), .A2(new_n2191_), .A3(new_n1187_), .ZN(new_n2353_));
  OAI21_X1   g2304(.A1(new_n2242_), .A2(new_n2244_), .B(new_n1188_), .ZN(new_n2354_));
  AOI21_X1   g2305(.A1(new_n2354_), .A2(new_n2353_), .B(new_n2352_), .ZN(new_n2355_));
  INV_X1     g2306(.I(new_n1261_), .ZN(new_n2356_));
  NOR4_X1    g2307(.A1(new_n2356_), .A2(new_n205_), .A3(new_n345_), .A4(new_n695_), .ZN(new_n2357_));
  NOR4_X1    g2308(.A1(new_n549_), .A2(new_n127_), .A3(new_n723_), .A4(new_n272_), .ZN(new_n2358_));
  NAND2_X1   g2309(.A1(new_n1068_), .A2(new_n393_), .ZN(new_n2359_));
  NOR4_X1    g2310(.A1(new_n2359_), .A2(new_n197_), .A3(new_n561_), .A4(new_n377_), .ZN(new_n2360_));
  NAND4_X1   g2311(.A1(new_n1023_), .A2(new_n438_), .A3(new_n483_), .A4(new_n556_), .ZN(new_n2361_));
  NOR4_X1    g2312(.A1(new_n2361_), .A2(new_n2330_), .A3(new_n376_), .A4(new_n387_), .ZN(new_n2362_));
  NAND4_X1   g2313(.A1(new_n2362_), .A2(new_n2357_), .A3(new_n2358_), .A4(new_n2360_), .ZN(new_n2363_));
  NOR3_X1    g2314(.A1(new_n918_), .A2(new_n193_), .A3(new_n373_), .ZN(new_n2364_));
  INV_X1     g2315(.I(new_n2364_), .ZN(new_n2365_));
  NOR4_X1    g2316(.A1(new_n854_), .A2(new_n536_), .A3(new_n548_), .A4(new_n207_), .ZN(new_n2366_));
  NOR4_X1    g2317(.A1(new_n2253_), .A2(new_n231_), .A3(new_n317_), .A4(new_n1153_), .ZN(new_n2367_));
  NAND3_X1   g2318(.A1(new_n2367_), .A2(new_n894_), .A3(new_n2366_), .ZN(new_n2368_));
  NOR3_X1    g2319(.A1(new_n2365_), .A2(new_n2363_), .A3(new_n2368_), .ZN(new_n2369_));
  INV_X1     g2320(.I(new_n2369_), .ZN(new_n2370_));
  NOR3_X1    g2321(.A1(new_n2227_), .A2(new_n2193_), .A3(new_n1396_), .ZN(new_n2371_));
  OAI21_X1   g2322(.A1(new_n2371_), .A2(new_n2190_), .B(new_n2370_), .ZN(new_n2372_));
  NOR3_X1    g2323(.A1(new_n2371_), .A2(new_n2190_), .A3(new_n2370_), .ZN(new_n2373_));
  NAND2_X1   g2324(.A1(new_n1397_), .A2(new_n1398_), .ZN(new_n2374_));
  INV_X1     g2325(.I(new_n2374_), .ZN(new_n2375_));
  NOR3_X1    g2326(.A1(new_n2226_), .A2(new_n2195_), .A3(new_n2375_), .ZN(new_n2376_));
  AOI21_X1   g2327(.A1(new_n2188_), .A2(new_n1494_), .B(new_n2374_), .ZN(new_n2377_));
  NOR3_X1    g2328(.A1(new_n981_), .A2(new_n974_), .A3(new_n976_), .ZN(new_n2378_));
  NOR2_X1    g2329(.A1(new_n353_), .A2(new_n285_), .ZN(new_n2379_));
  INV_X1     g2330(.I(new_n2379_), .ZN(new_n2380_));
  NOR4_X1    g2331(.A1(new_n2263_), .A2(new_n234_), .A3(new_n2380_), .A4(new_n1265_), .ZN(new_n2381_));
  NOR4_X1    g2332(.A1(new_n440_), .A2(new_n400_), .A3(new_n736_), .A4(new_n718_), .ZN(new_n2382_));
  INV_X1     g2333(.I(new_n2382_), .ZN(new_n2383_));
  NAND4_X1   g2334(.A1(new_n1119_), .A2(new_n301_), .A3(new_n902_), .A4(new_n555_), .ZN(new_n2384_));
  NOR3_X1    g2335(.A1(new_n373_), .A2(new_n515_), .A3(new_n573_), .ZN(new_n2385_));
  INV_X1     g2336(.I(new_n2385_), .ZN(new_n2386_));
  NOR4_X1    g2337(.A1(new_n2383_), .A2(new_n199_), .A3(new_n2384_), .A4(new_n2386_), .ZN(new_n2387_));
  NAND4_X1   g2338(.A1(new_n2387_), .A2(new_n2378_), .A3(new_n923_), .A4(new_n2381_), .ZN(new_n2388_));
  INV_X1     g2339(.I(new_n2388_), .ZN(new_n2389_));
  OAI21_X1   g2340(.A1(new_n2376_), .A2(new_n2377_), .B(new_n2389_), .ZN(new_n2390_));
  NOR4_X1    g2341(.A1(new_n854_), .A2(new_n296_), .A3(new_n313_), .A4(new_n495_), .ZN(new_n2391_));
  NOR4_X1    g2342(.A1(new_n485_), .A2(new_n294_), .A3(new_n262_), .A4(new_n548_), .ZN(new_n2392_));
  NAND4_X1   g2343(.A1(new_n581_), .A2(new_n674_), .A3(new_n909_), .A4(new_n329_), .ZN(new_n2393_));
  NOR4_X1    g2344(.A1(new_n2393_), .A2(new_n317_), .A3(new_n382_), .A4(new_n415_), .ZN(new_n2394_));
  NAND4_X1   g2345(.A1(new_n2394_), .A2(new_n2282_), .A3(new_n2391_), .A4(new_n2392_), .ZN(new_n2395_));
  NOR4_X1    g2346(.A1(new_n179_), .A2(new_n202_), .A3(new_n515_), .A4(new_n497_), .ZN(new_n2396_));
  NOR3_X1    g2347(.A1(new_n250_), .A2(new_n267_), .A3(new_n205_), .ZN(new_n2397_));
  NOR2_X1    g2348(.A1(new_n587_), .A2(new_n2356_), .ZN(new_n2398_));
  INV_X1     g2349(.I(new_n2398_), .ZN(new_n2399_));
  NOR3_X1    g2350(.A1(new_n2399_), .A2(new_n164_), .A3(new_n378_), .ZN(new_n2400_));
  NAND4_X1   g2351(.A1(new_n2400_), .A2(new_n907_), .A3(new_n2396_), .A4(new_n2397_), .ZN(new_n2401_));
  NOR3_X1    g2352(.A1(new_n2258_), .A2(new_n2395_), .A3(new_n2401_), .ZN(new_n2402_));
  INV_X1     g2353(.I(new_n2402_), .ZN(new_n2403_));
  NAND2_X1   g2354(.A1(new_n1494_), .A2(new_n1497_), .ZN(new_n2404_));
  AOI21_X1   g2355(.A1(new_n2183_), .A2(new_n2187_), .B(new_n2404_), .ZN(new_n2405_));
  NOR2_X1    g2356(.A1(new_n2195_), .A2(new_n2196_), .ZN(new_n2406_));
  NOR3_X1    g2357(.A1(new_n2225_), .A2(new_n2186_), .A3(new_n2406_), .ZN(new_n2407_));
  OAI21_X1   g2358(.A1(new_n2407_), .A2(new_n2405_), .B(new_n2403_), .ZN(new_n2408_));
  AOI21_X1   g2359(.A1(new_n2224_), .A2(new_n2200_), .B(new_n1592_), .ZN(new_n2409_));
  NOR3_X1    g2360(.A1(new_n2182_), .A2(new_n2199_), .A3(new_n1632_), .ZN(new_n2410_));
  INV_X1     g2361(.I(new_n327_), .ZN(new_n2411_));
  NAND4_X1   g2362(.A1(new_n553_), .A2(new_n292_), .A3(new_n2411_), .A4(new_n677_), .ZN(new_n2412_));
  NOR2_X1    g2363(.A1(new_n267_), .A2(new_n360_), .ZN(new_n2413_));
  NOR3_X1    g2364(.A1(new_n549_), .A2(new_n415_), .A3(new_n444_), .ZN(new_n2414_));
  NAND4_X1   g2365(.A1(new_n2414_), .A2(new_n372_), .A3(new_n2413_), .A4(new_n380_), .ZN(new_n2415_));
  NOR4_X1    g2366(.A1(new_n389_), .A2(new_n691_), .A3(new_n452_), .A4(new_n561_), .ZN(new_n2416_));
  NAND4_X1   g2367(.A1(new_n2416_), .A2(new_n531_), .A3(new_n275_), .A4(new_n351_), .ZN(new_n2417_));
  NOR4_X1    g2368(.A1(new_n2417_), .A2(new_n2412_), .A3(new_n2415_), .A4(new_n974_), .ZN(new_n2418_));
  INV_X1     g2369(.I(new_n2418_), .ZN(new_n2419_));
  NAND2_X1   g2370(.A1(new_n354_), .A2(new_n589_), .ZN(new_n2420_));
  INV_X1     g2371(.I(new_n2420_), .ZN(new_n2421_));
  NOR4_X1    g2372(.A1(new_n193_), .A2(new_n253_), .A3(new_n545_), .A4(new_n196_), .ZN(new_n2422_));
  NAND4_X1   g2373(.A1(new_n2421_), .A2(new_n1012_), .A3(new_n2319_), .A4(new_n2422_), .ZN(new_n2423_));
  NOR3_X1    g2374(.A1(new_n2419_), .A2(new_n803_), .A3(new_n2423_), .ZN(new_n2424_));
  NOR3_X1    g2375(.A1(new_n2409_), .A2(new_n2410_), .A3(new_n2424_), .ZN(new_n2425_));
  NAND3_X1   g2376(.A1(new_n2175_), .A2(new_n2114_), .A3(new_n2107_), .ZN(new_n2426_));
  INV_X1     g2377(.I(new_n1141_), .ZN(new_n2427_));
  NOR2_X1    g2378(.A1(new_n738_), .A2(new_n789_), .ZN(new_n2428_));
  NAND3_X1   g2379(.A1(new_n1092_), .A2(new_n674_), .A3(new_n447_), .ZN(new_n2429_));
  NOR4_X1    g2380(.A1(new_n527_), .A2(new_n296_), .A3(new_n557_), .A4(new_n2429_), .ZN(new_n2430_));
  NAND4_X1   g2381(.A1(new_n2430_), .A2(new_n917_), .A3(new_n2428_), .A4(new_n2427_), .ZN(new_n2431_));
  NOR3_X1    g2382(.A1(new_n2287_), .A2(new_n2423_), .A3(new_n2431_), .ZN(new_n2432_));
  NAND3_X1   g2383(.A1(new_n2221_), .A2(new_n2426_), .A3(new_n2432_), .ZN(new_n2433_));
  NOR3_X1    g2384(.A1(new_n256_), .A2(new_n536_), .A3(new_n454_), .ZN(new_n2434_));
  NOR2_X1    g2385(.A1(new_n250_), .A2(new_n110_), .ZN(new_n2435_));
  INV_X1     g2386(.I(new_n2435_), .ZN(new_n2436_));
  NOR4_X1    g2387(.A1(new_n2436_), .A2(new_n2290_), .A3(new_n548_), .A4(new_n1154_), .ZN(new_n2437_));
  NOR2_X1    g2388(.A1(new_n516_), .A2(new_n200_), .ZN(new_n2438_));
  NAND2_X1   g2389(.A1(new_n436_), .A2(new_n408_), .ZN(new_n2439_));
  NOR4_X1    g2390(.A1(new_n2439_), .A2(new_n259_), .A3(new_n492_), .A4(new_n339_), .ZN(new_n2440_));
  NAND4_X1   g2391(.A1(new_n2437_), .A2(new_n2440_), .A3(new_n2434_), .A4(new_n2438_), .ZN(new_n2441_));
  NOR4_X1    g2392(.A1(new_n312_), .A2(new_n356_), .A3(new_n156_), .A4(new_n557_), .ZN(new_n2442_));
  NOR4_X1    g2393(.A1(new_n723_), .A2(new_n437_), .A3(new_n207_), .A4(new_n415_), .ZN(new_n2443_));
  NOR2_X1    g2394(.A1(new_n389_), .A2(new_n205_), .ZN(new_n2444_));
  INV_X1     g2395(.I(new_n2444_), .ZN(new_n2445_));
  NOR4_X1    g2396(.A1(new_n2445_), .A2(new_n265_), .A3(new_n267_), .A4(new_n876_), .ZN(new_n2446_));
  NAND4_X1   g2397(.A1(new_n2446_), .A2(new_n688_), .A3(new_n2442_), .A4(new_n2443_), .ZN(new_n2447_));
  NOR3_X1    g2398(.A1(new_n2447_), .A2(new_n2441_), .A3(new_n199_), .ZN(new_n2448_));
  INV_X1     g2399(.I(new_n2448_), .ZN(new_n2449_));
  NOR2_X1    g2400(.A1(new_n2433_), .A2(new_n2449_), .ZN(new_n2450_));
  INV_X1     g2401(.I(new_n2450_), .ZN(new_n2451_));
  NAND2_X1   g2402(.A1(new_n2433_), .A2(new_n2449_), .ZN(new_n2452_));
  OAI21_X1   g2403(.A1(new_n2176_), .A2(new_n2113_), .B(new_n1694_), .ZN(new_n2453_));
  NAND3_X1   g2404(.A1(new_n2222_), .A2(new_n2453_), .A3(new_n2111_), .ZN(new_n2454_));
  AOI21_X1   g2405(.A1(new_n2221_), .A2(new_n1748_), .B(new_n2201_), .ZN(new_n2455_));
  OAI21_X1   g2406(.A1(new_n2455_), .A2(new_n2177_), .B(new_n2215_), .ZN(new_n2456_));
  NAND3_X1   g2407(.A1(new_n2456_), .A2(new_n2454_), .A3(new_n2452_), .ZN(new_n2457_));
  INV_X1     g2408(.I(new_n571_), .ZN(new_n2458_));
  NOR3_X1    g2409(.A1(new_n545_), .A2(new_n722_), .A3(new_n272_), .ZN(new_n2459_));
  NAND4_X1   g2410(.A1(new_n2459_), .A2(new_n224_), .A3(new_n887_), .A4(new_n740_), .ZN(new_n2460_));
  NOR2_X1    g2411(.A1(new_n426_), .A2(new_n524_), .ZN(new_n2461_));
  NAND3_X1   g2412(.A1(new_n702_), .A2(new_n2461_), .A3(new_n318_), .ZN(new_n2462_));
  NOR4_X1    g2413(.A1(new_n2415_), .A2(new_n2460_), .A3(new_n2462_), .A4(new_n1074_), .ZN(new_n2463_));
  INV_X1     g2414(.I(new_n851_), .ZN(new_n2464_));
  NOR3_X1    g2415(.A1(new_n2464_), .A2(new_n527_), .A3(new_n2445_), .ZN(new_n2465_));
  NOR2_X1    g2416(.A1(new_n509_), .A2(new_n580_), .ZN(new_n2466_));
  INV_X1     g2417(.I(new_n2466_), .ZN(new_n2467_));
  NOR4_X1    g2418(.A1(new_n2467_), .A2(new_n277_), .A3(new_n299_), .A4(new_n401_), .ZN(new_n2468_));
  NOR2_X1    g2419(.A1(new_n454_), .A2(new_n485_), .ZN(new_n2469_));
  NAND3_X1   g2420(.A1(new_n2469_), .A2(new_n368_), .A3(new_n447_), .ZN(new_n2470_));
  NOR3_X1    g2421(.A1(new_n2346_), .A2(new_n2470_), .A3(new_n863_), .ZN(new_n2471_));
  NAND4_X1   g2422(.A1(new_n2471_), .A2(new_n2382_), .A3(new_n2465_), .A4(new_n2468_), .ZN(new_n2472_));
  INV_X1     g2423(.I(new_n2472_), .ZN(new_n2473_));
  NAND4_X1   g2424(.A1(new_n2473_), .A2(new_n2458_), .A3(new_n2463_), .A4(new_n915_), .ZN(new_n2474_));
  AOI21_X1   g2425(.A1(new_n2457_), .A2(new_n2451_), .B(new_n2474_), .ZN(new_n2475_));
  NOR2_X1    g2426(.A1(new_n2181_), .A2(new_n1632_), .ZN(new_n2476_));
  OAI21_X1   g2427(.A1(new_n2112_), .A2(new_n2177_), .B(new_n2476_), .ZN(new_n2477_));
  NOR2_X1    g2428(.A1(new_n2112_), .A2(new_n2177_), .ZN(new_n2478_));
  NAND2_X1   g2429(.A1(new_n2200_), .A2(new_n2223_), .ZN(new_n2479_));
  NAND2_X1   g2430(.A1(new_n2478_), .A2(new_n2479_), .ZN(new_n2480_));
  NAND2_X1   g2431(.A1(new_n2480_), .A2(new_n2477_), .ZN(new_n2481_));
  NAND3_X1   g2432(.A1(new_n2457_), .A2(new_n2451_), .A3(new_n2474_), .ZN(new_n2482_));
  AOI21_X1   g2433(.A1(new_n2481_), .A2(new_n2482_), .B(new_n2475_), .ZN(new_n2483_));
  OAI21_X1   g2434(.A1(new_n2409_), .A2(new_n2410_), .B(new_n2424_), .ZN(new_n2484_));
  AOI21_X1   g2435(.A1(new_n2483_), .A2(new_n2484_), .B(new_n2425_), .ZN(new_n2485_));
  NOR3_X1    g2436(.A1(new_n2407_), .A2(new_n2405_), .A3(new_n2403_), .ZN(new_n2486_));
  OAI21_X1   g2437(.A1(new_n2485_), .A2(new_n2486_), .B(new_n2408_), .ZN(new_n2487_));
  NOR3_X1    g2438(.A1(new_n2376_), .A2(new_n2377_), .A3(new_n2389_), .ZN(new_n2488_));
  OAI21_X1   g2439(.A1(new_n2487_), .A2(new_n2488_), .B(new_n2390_), .ZN(new_n2489_));
  OAI21_X1   g2440(.A1(new_n2489_), .A2(new_n2373_), .B(new_n2372_), .ZN(new_n2490_));
  NAND3_X1   g2441(.A1(new_n2354_), .A2(new_n2353_), .A3(new_n2352_), .ZN(new_n2491_));
  AOI21_X1   g2442(.A1(new_n2490_), .A2(new_n2491_), .B(new_n2355_), .ZN(new_n2492_));
  OAI21_X1   g2443(.A1(new_n2492_), .A2(new_n2337_), .B(new_n2315_), .ZN(new_n2493_));
  NAND2_X1   g2444(.A1(new_n2492_), .A2(new_n2337_), .ZN(new_n2494_));
  AOI21_X1   g2445(.A1(new_n2232_), .A2(new_n970_), .B(new_n2241_), .ZN(new_n2495_));
  NOR3_X1    g2446(.A1(new_n2245_), .A2(new_n827_), .A3(new_n969_), .ZN(new_n2496_));
  INV_X1     g2447(.I(new_n2309_), .ZN(new_n2497_));
  NOR3_X1    g2448(.A1(new_n2496_), .A2(new_n2495_), .A3(new_n2497_), .ZN(new_n2498_));
  AOI21_X1   g2449(.A1(new_n2493_), .A2(new_n2494_), .B(new_n2498_), .ZN(new_n2499_));
  INV_X1     g2450(.I(new_n2295_), .ZN(new_n2500_));
  AOI21_X1   g2451(.A1(new_n2246_), .A2(new_n2235_), .B(new_n2298_), .ZN(new_n2501_));
  NOR3_X1    g2452(.A1(new_n2233_), .A2(new_n2236_), .A3(new_n2296_), .ZN(new_n2502_));
  NOR3_X1    g2453(.A1(new_n2501_), .A2(new_n2502_), .A3(new_n2500_), .ZN(new_n2503_));
  NOR4_X1    g2454(.A1(new_n2499_), .A2(new_n2300_), .A3(new_n2310_), .A4(new_n2503_), .ZN(new_n2504_));
  NOR2_X1    g2455(.A1(new_n2504_), .A2(new_n2300_), .ZN(new_n2505_));
  NAND3_X1   g2456(.A1(new_n2248_), .A2(new_n2238_), .A3(new_n2270_), .ZN(new_n2506_));
  AOI21_X1   g2457(.A1(new_n2505_), .A2(new_n2506_), .B(new_n2271_), .ZN(new_n2507_));
  NOR2_X1    g2458(.A1(new_n2507_), .A2(new_n308_), .ZN(new_n2508_));
  INV_X1     g2459(.I(new_n2271_), .ZN(new_n2509_));
  OAI21_X1   g2460(.A1(new_n2501_), .A2(new_n2502_), .B(new_n2500_), .ZN(new_n2510_));
  OAI21_X1   g2461(.A1(new_n2496_), .A2(new_n2495_), .B(new_n2497_), .ZN(new_n2511_));
  AOI21_X1   g2462(.A1(new_n2192_), .A2(new_n2229_), .B(new_n2313_), .ZN(new_n2512_));
  NOR3_X1    g2463(.A1(new_n2243_), .A2(new_n2244_), .A3(new_n2311_), .ZN(new_n2513_));
  NOR2_X1    g2464(.A1(new_n2513_), .A2(new_n2512_), .ZN(new_n2514_));
  INV_X1     g2465(.I(new_n2337_), .ZN(new_n2515_));
  NOR3_X1    g2466(.A1(new_n2242_), .A2(new_n2244_), .A3(new_n1188_), .ZN(new_n2516_));
  AOI21_X1   g2467(.A1(new_n2229_), .A2(new_n2191_), .B(new_n1187_), .ZN(new_n2517_));
  OAI21_X1   g2468(.A1(new_n2517_), .A2(new_n2516_), .B(new_n2351_), .ZN(new_n2518_));
  NAND3_X1   g2469(.A1(new_n2189_), .A2(new_n1243_), .A3(new_n1397_), .ZN(new_n2519_));
  AOI21_X1   g2470(.A1(new_n2228_), .A2(new_n2519_), .B(new_n2369_), .ZN(new_n2520_));
  NAND3_X1   g2471(.A1(new_n2228_), .A2(new_n2519_), .A3(new_n2369_), .ZN(new_n2521_));
  NAND3_X1   g2472(.A1(new_n2188_), .A2(new_n1494_), .A3(new_n2374_), .ZN(new_n2522_));
  OAI21_X1   g2473(.A1(new_n2226_), .A2(new_n2195_), .B(new_n2375_), .ZN(new_n2523_));
  AOI21_X1   g2474(.A1(new_n2523_), .A2(new_n2522_), .B(new_n2388_), .ZN(new_n2524_));
  OAI21_X1   g2475(.A1(new_n2225_), .A2(new_n2186_), .B(new_n2406_), .ZN(new_n2525_));
  NAND3_X1   g2476(.A1(new_n2183_), .A2(new_n2187_), .A3(new_n2404_), .ZN(new_n2526_));
  AOI21_X1   g2477(.A1(new_n2525_), .A2(new_n2526_), .B(new_n2402_), .ZN(new_n2527_));
  INV_X1     g2478(.I(new_n2425_), .ZN(new_n2528_));
  NOR3_X1    g2479(.A1(new_n2220_), .A2(new_n1798_), .A3(new_n2213_), .ZN(new_n2529_));
  NOR2_X1    g2480(.A1(new_n2529_), .A2(new_n2176_), .ZN(new_n2530_));
  AOI21_X1   g2481(.A1(new_n2530_), .A2(new_n2432_), .B(new_n2448_), .ZN(new_n2531_));
  NOR3_X1    g2482(.A1(new_n2455_), .A2(new_n2177_), .A3(new_n2215_), .ZN(new_n2532_));
  AOI21_X1   g2483(.A1(new_n2222_), .A2(new_n2453_), .B(new_n2111_), .ZN(new_n2533_));
  NOR3_X1    g2484(.A1(new_n2532_), .A2(new_n2533_), .A3(new_n2531_), .ZN(new_n2534_));
  INV_X1     g2485(.I(new_n2474_), .ZN(new_n2535_));
  OAI21_X1   g2486(.A1(new_n2534_), .A2(new_n2450_), .B(new_n2535_), .ZN(new_n2536_));
  NOR2_X1    g2487(.A1(new_n2478_), .A2(new_n2479_), .ZN(new_n2537_));
  NOR3_X1    g2488(.A1(new_n2476_), .A2(new_n2112_), .A3(new_n2177_), .ZN(new_n2538_));
  NOR2_X1    g2489(.A1(new_n2537_), .A2(new_n2538_), .ZN(new_n2539_));
  NOR3_X1    g2490(.A1(new_n2534_), .A2(new_n2450_), .A3(new_n2535_), .ZN(new_n2540_));
  OAI21_X1   g2491(.A1(new_n2539_), .A2(new_n2540_), .B(new_n2536_), .ZN(new_n2541_));
  INV_X1     g2492(.I(new_n2484_), .ZN(new_n2542_));
  OAI21_X1   g2493(.A1(new_n2541_), .A2(new_n2542_), .B(new_n2528_), .ZN(new_n2543_));
  NAND3_X1   g2494(.A1(new_n2525_), .A2(new_n2526_), .A3(new_n2402_), .ZN(new_n2544_));
  AOI21_X1   g2495(.A1(new_n2543_), .A2(new_n2544_), .B(new_n2527_), .ZN(new_n2545_));
  NAND3_X1   g2496(.A1(new_n2523_), .A2(new_n2522_), .A3(new_n2388_), .ZN(new_n2546_));
  AOI21_X1   g2497(.A1(new_n2545_), .A2(new_n2546_), .B(new_n2524_), .ZN(new_n2547_));
  AOI21_X1   g2498(.A1(new_n2547_), .A2(new_n2521_), .B(new_n2520_), .ZN(new_n2548_));
  NOR3_X1    g2499(.A1(new_n2517_), .A2(new_n2516_), .A3(new_n2351_), .ZN(new_n2549_));
  OAI21_X1   g2500(.A1(new_n2548_), .A2(new_n2549_), .B(new_n2518_), .ZN(new_n2550_));
  AOI21_X1   g2501(.A1(new_n2550_), .A2(new_n2515_), .B(new_n2514_), .ZN(new_n2551_));
  NOR2_X1    g2502(.A1(new_n2550_), .A2(new_n2515_), .ZN(new_n2552_));
  NAND3_X1   g2503(.A1(new_n2301_), .A2(new_n2302_), .A3(new_n2309_), .ZN(new_n2553_));
  OAI21_X1   g2504(.A1(new_n2551_), .A2(new_n2552_), .B(new_n2553_), .ZN(new_n2554_));
  NAND3_X1   g2505(.A1(new_n2299_), .A2(new_n2297_), .A3(new_n2295_), .ZN(new_n2555_));
  NAND4_X1   g2506(.A1(new_n2554_), .A2(new_n2510_), .A3(new_n2511_), .A4(new_n2555_), .ZN(new_n2556_));
  NAND2_X1   g2507(.A1(new_n2556_), .A2(new_n2510_), .ZN(new_n2557_));
  AOI21_X1   g2508(.A1(new_n2247_), .A2(new_n2240_), .B(new_n2239_), .ZN(new_n2558_));
  NOR3_X1    g2509(.A1(new_n2237_), .A2(new_n612_), .A3(new_n655_), .ZN(new_n2559_));
  NOR3_X1    g2510(.A1(new_n2558_), .A2(new_n2559_), .A3(new_n2269_), .ZN(new_n2560_));
  OAI21_X1   g2511(.A1(new_n2557_), .A2(new_n2560_), .B(new_n2509_), .ZN(new_n2561_));
  NOR2_X1    g2512(.A1(new_n2561_), .A2(new_n307_), .ZN(new_n2562_));
  NOR2_X1    g2513(.A1(new_n2508_), .A2(new_n2562_), .ZN(new_n2563_));
  NOR2_X1    g2514(.A1(new_n2563_), .A2(new_n56_), .ZN(new_n2564_));
  NAND3_X1   g2515(.A1(new_n899_), .A2(new_n530_), .A3(new_n871_), .ZN(new_n2565_));
  NOR4_X1    g2516(.A1(new_n277_), .A2(new_n110_), .A3(new_n435_), .A4(new_n402_), .ZN(new_n2566_));
  NOR3_X1    g2517(.A1(new_n312_), .A2(new_n321_), .A3(new_n450_), .ZN(new_n2567_));
  NAND4_X1   g2518(.A1(new_n802_), .A2(new_n2567_), .A3(new_n2397_), .A4(new_n2566_), .ZN(new_n2568_));
  NOR4_X1    g2519(.A1(new_n2568_), .A2(new_n1120_), .A3(new_n567_), .A4(new_n2565_), .ZN(new_n2569_));
  NOR4_X1    g2520(.A1(new_n854_), .A2(new_n448_), .A3(new_n271_), .A4(new_n360_), .ZN(new_n2570_));
  NAND3_X1   g2521(.A1(new_n699_), .A2(new_n1271_), .A3(new_n491_), .ZN(new_n2571_));
  INV_X1     g2522(.I(new_n2571_), .ZN(new_n2572_));
  NOR2_X1    g2523(.A1(new_n276_), .A2(new_n299_), .ZN(new_n2573_));
  INV_X1     g2524(.I(new_n2573_), .ZN(new_n2574_));
  NOR3_X1    g2525(.A1(new_n2574_), .A2(new_n400_), .A3(new_n327_), .ZN(new_n2575_));
  NAND2_X1   g2526(.A1(new_n890_), .A2(new_n900_), .ZN(new_n2576_));
  NOR4_X1    g2527(.A1(new_n2576_), .A2(new_n296_), .A3(new_n378_), .A4(new_n2356_), .ZN(new_n2577_));
  NAND4_X1   g2528(.A1(new_n2575_), .A2(new_n429_), .A3(new_n374_), .A4(new_n2577_), .ZN(new_n2578_));
  INV_X1     g2529(.I(new_n2578_), .ZN(new_n2579_));
  NAND4_X1   g2530(.A1(new_n2579_), .A2(new_n2289_), .A3(new_n2570_), .A4(new_n2572_), .ZN(new_n2580_));
  INV_X1     g2531(.I(new_n2580_), .ZN(new_n2581_));
  NAND3_X1   g2532(.A1(new_n2581_), .A2(new_n734_), .A3(new_n2569_), .ZN(new_n2582_));
  OAI21_X1   g2533(.A1(new_n2507_), .A2(new_n308_), .B(new_n2582_), .ZN(new_n2583_));
  INV_X1     g2534(.I(new_n2582_), .ZN(new_n2584_));
  NAND3_X1   g2535(.A1(new_n2561_), .A2(new_n307_), .A3(new_n2584_), .ZN(new_n2585_));
  AND2_X2    g2536(.A1(new_n2583_), .A2(new_n2585_), .Z(new_n2586_));
  NOR2_X1    g2537(.A1(new_n1449_), .A2(\a[0] ), .ZN(new_n2587_));
  INV_X1     g2538(.I(new_n2587_), .ZN(new_n2588_));
  NOR2_X1    g2539(.A1(new_n2586_), .A2(new_n2588_), .ZN(new_n2589_));
  NAND4_X1   g2540(.A1(new_n1000_), .A2(new_n1431_), .A3(new_n739_), .A4(new_n797_), .ZN(new_n2590_));
  OR3_X2     g2541(.A1(new_n2467_), .A2(new_n2590_), .A3(new_n881_), .Z(new_n2591_));
  NOR4_X1    g2542(.A1(new_n2591_), .A2(new_n544_), .A3(new_n587_), .A4(new_n1511_), .ZN(new_n2592_));
  NOR4_X1    g2543(.A1(new_n2383_), .A2(new_n375_), .A3(new_n384_), .A4(new_n2334_), .ZN(new_n2593_));
  NAND3_X1   g2544(.A1(new_n364_), .A2(new_n2593_), .A3(new_n2592_), .ZN(new_n2594_));
  INV_X1     g2545(.I(new_n2594_), .ZN(new_n2595_));
  NAND2_X1   g2546(.A1(new_n2585_), .A2(new_n2595_), .ZN(new_n2596_));
  NAND3_X1   g2547(.A1(new_n2508_), .A2(new_n2584_), .A3(new_n2594_), .ZN(new_n2597_));
  NAND2_X1   g2548(.A1(new_n2597_), .A2(new_n2596_), .ZN(new_n2598_));
  NOR2_X1    g2549(.A1(new_n1449_), .A2(new_n53_), .ZN(new_n2599_));
  NOR2_X1    g2550(.A1(\a[1] ), .A2(\a[2] ), .ZN(new_n2600_));
  OAI21_X1   g2551(.A1(new_n2599_), .A2(new_n2600_), .B(\a[0] ), .ZN(new_n2601_));
  NOR2_X1    g2552(.A1(new_n2598_), .A2(new_n2601_), .ZN(new_n2602_));
  NOR3_X1    g2553(.A1(new_n2602_), .A2(new_n2589_), .A3(new_n2564_), .ZN(new_n2603_));
  NAND2_X1   g2554(.A1(new_n2583_), .A2(new_n2585_), .ZN(new_n2604_));
  NAND2_X1   g2555(.A1(new_n2561_), .A2(new_n307_), .ZN(new_n2605_));
  NAND2_X1   g2556(.A1(new_n2507_), .A2(new_n308_), .ZN(new_n2606_));
  NOR2_X1    g2557(.A1(new_n2560_), .A2(new_n2271_), .ZN(new_n2607_));
  NAND2_X1   g2558(.A1(new_n2557_), .A2(new_n2607_), .ZN(new_n2608_));
  NAND2_X1   g2559(.A1(new_n2509_), .A2(new_n2506_), .ZN(new_n2609_));
  NAND2_X1   g2560(.A1(new_n2505_), .A2(new_n2609_), .ZN(new_n2610_));
  NAND2_X1   g2561(.A1(new_n2610_), .A2(new_n2608_), .ZN(new_n2611_));
  AOI22_X1   g2562(.A1(new_n2554_), .A2(new_n2511_), .B1(new_n2510_), .B2(new_n2555_), .ZN(new_n2612_));
  NOR2_X1    g2563(.A1(new_n2612_), .A2(new_n2504_), .ZN(new_n2613_));
  NAND3_X1   g2564(.A1(new_n2312_), .A2(new_n2314_), .A3(new_n2337_), .ZN(new_n2614_));
  OAI21_X1   g2565(.A1(new_n2513_), .A2(new_n2512_), .B(new_n2515_), .ZN(new_n2615_));
  NAND2_X1   g2566(.A1(new_n2615_), .A2(new_n2614_), .ZN(new_n2616_));
  NOR2_X1    g2567(.A1(new_n2616_), .A2(new_n2492_), .ZN(new_n2617_));
  AOI21_X1   g2568(.A1(new_n2614_), .A2(new_n2615_), .B(new_n2550_), .ZN(new_n2618_));
  NOR3_X1    g2569(.A1(new_n2549_), .A2(new_n2355_), .A3(new_n2548_), .ZN(new_n2619_));
  AOI21_X1   g2570(.A1(new_n2518_), .A2(new_n2491_), .B(new_n2490_), .ZN(new_n2620_));
  NOR2_X1    g2571(.A1(new_n2373_), .A2(new_n2520_), .ZN(new_n2621_));
  NAND2_X1   g2572(.A1(new_n2621_), .A2(new_n2547_), .ZN(new_n2622_));
  NAND2_X1   g2573(.A1(new_n2372_), .A2(new_n2521_), .ZN(new_n2623_));
  NAND2_X1   g2574(.A1(new_n2623_), .A2(new_n2489_), .ZN(new_n2624_));
  NAND3_X1   g2575(.A1(new_n2523_), .A2(new_n2522_), .A3(new_n974_), .ZN(new_n2625_));
  NAND3_X1   g2576(.A1(new_n2390_), .A2(new_n2546_), .A3(new_n2625_), .ZN(new_n2626_));
  NOR2_X1    g2577(.A1(new_n2626_), .A2(new_n2545_), .ZN(new_n2627_));
  NOR2_X1    g2578(.A1(new_n2488_), .A2(new_n2524_), .ZN(new_n2628_));
  NOR2_X1    g2579(.A1(new_n2628_), .A2(new_n2487_), .ZN(new_n2629_));
  NOR2_X1    g2580(.A1(new_n2627_), .A2(new_n2629_), .ZN(new_n2630_));
  NAND3_X1   g2581(.A1(new_n2485_), .A2(new_n2408_), .A3(new_n2544_), .ZN(new_n2631_));
  NAND2_X1   g2582(.A1(new_n2408_), .A2(new_n2544_), .ZN(new_n2632_));
  NAND2_X1   g2583(.A1(new_n2632_), .A2(new_n2543_), .ZN(new_n2633_));
  NAND2_X1   g2584(.A1(new_n2482_), .A2(new_n2481_), .ZN(new_n2634_));
  OAI21_X1   g2585(.A1(new_n2182_), .A2(new_n1632_), .B(new_n2199_), .ZN(new_n2635_));
  NAND3_X1   g2586(.A1(new_n2224_), .A2(new_n1592_), .A3(new_n2200_), .ZN(new_n2636_));
  NAND3_X1   g2587(.A1(new_n2636_), .A2(new_n2635_), .A3(new_n2424_), .ZN(new_n2637_));
  INV_X1     g2588(.I(new_n2424_), .ZN(new_n2638_));
  OAI21_X1   g2589(.A1(new_n2409_), .A2(new_n2410_), .B(new_n2638_), .ZN(new_n2639_));
  NAND4_X1   g2590(.A1(new_n2634_), .A2(new_n2536_), .A3(new_n2639_), .A4(new_n2637_), .ZN(new_n2640_));
  NOR2_X1    g2591(.A1(new_n2540_), .A2(new_n2539_), .ZN(new_n2641_));
  NOR3_X1    g2592(.A1(new_n2409_), .A2(new_n2410_), .A3(new_n2638_), .ZN(new_n2642_));
  AOI21_X1   g2593(.A1(new_n2636_), .A2(new_n2635_), .B(new_n2424_), .ZN(new_n2643_));
  OAI22_X1   g2594(.A1(new_n2641_), .A2(new_n2475_), .B1(new_n2642_), .B2(new_n2643_), .ZN(new_n2644_));
  NAND2_X1   g2595(.A1(new_n2644_), .A2(new_n2640_), .ZN(new_n2645_));
  AOI21_X1   g2596(.A1(new_n2536_), .A2(new_n2482_), .B(new_n2539_), .ZN(new_n2646_));
  NOR3_X1    g2597(.A1(new_n2540_), .A2(new_n2475_), .A3(new_n2481_), .ZN(new_n2647_));
  NAND2_X1   g2598(.A1(new_n2433_), .A2(new_n2448_), .ZN(new_n2648_));
  NAND3_X1   g2599(.A1(new_n2530_), .A2(new_n2432_), .A3(new_n2449_), .ZN(new_n2649_));
  NAND4_X1   g2600(.A1(new_n2454_), .A2(new_n2456_), .A3(new_n2649_), .A4(new_n2648_), .ZN(new_n2650_));
  NAND2_X1   g2601(.A1(new_n2456_), .A2(new_n2454_), .ZN(new_n2651_));
  NAND2_X1   g2602(.A1(new_n2649_), .A2(new_n2648_), .ZN(new_n2652_));
  NAND2_X1   g2603(.A1(new_n2651_), .A2(new_n2652_), .ZN(new_n2653_));
  NAND2_X1   g2604(.A1(new_n2653_), .A2(new_n2650_), .ZN(new_n2654_));
  INV_X1     g2605(.I(new_n2433_), .ZN(new_n2655_));
  NOR2_X1    g2606(.A1(new_n2530_), .A2(new_n2432_), .ZN(new_n2656_));
  NOR2_X1    g2607(.A1(new_n2656_), .A2(new_n2655_), .ZN(new_n2657_));
  OAI22_X1   g2608(.A1(new_n2647_), .A2(new_n2646_), .B1(new_n2654_), .B2(new_n2657_), .ZN(new_n2658_));
  NAND2_X1   g2609(.A1(new_n2645_), .A2(new_n2658_), .ZN(new_n2659_));
  NAND3_X1   g2610(.A1(new_n2659_), .A2(new_n2631_), .A3(new_n2633_), .ZN(new_n2660_));
  AOI22_X1   g2611(.A1(new_n2622_), .A2(new_n2624_), .B1(new_n2630_), .B2(new_n2660_), .ZN(new_n2661_));
  NOR3_X1    g2612(.A1(new_n2661_), .A2(new_n2619_), .A3(new_n2620_), .ZN(new_n2662_));
  NOR3_X1    g2613(.A1(new_n2617_), .A2(new_n2618_), .A3(new_n2662_), .ZN(new_n2663_));
  NAND4_X1   g2614(.A1(new_n2493_), .A2(new_n2494_), .A3(new_n2511_), .A4(new_n2553_), .ZN(new_n2664_));
  OAI22_X1   g2615(.A1(new_n2551_), .A2(new_n2552_), .B1(new_n2310_), .B2(new_n2498_), .ZN(new_n2665_));
  NAND2_X1   g2616(.A1(new_n2665_), .A2(new_n2664_), .ZN(new_n2666_));
  OAI22_X1   g2617(.A1(new_n2612_), .A2(new_n2504_), .B1(new_n2666_), .B2(new_n2663_), .ZN(new_n2667_));
  NAND3_X1   g2618(.A1(new_n2550_), .A2(new_n2614_), .A3(new_n2615_), .ZN(new_n2668_));
  NAND2_X1   g2619(.A1(new_n2616_), .A2(new_n2492_), .ZN(new_n2669_));
  NAND2_X1   g2620(.A1(new_n2669_), .A2(new_n2668_), .ZN(new_n2670_));
  NOR2_X1    g2621(.A1(new_n2619_), .A2(new_n2620_), .ZN(new_n2671_));
  NOR2_X1    g2622(.A1(new_n2623_), .A2(new_n2489_), .ZN(new_n2672_));
  NOR2_X1    g2623(.A1(new_n2621_), .A2(new_n2547_), .ZN(new_n2673_));
  NAND3_X1   g2624(.A1(new_n2628_), .A2(new_n2487_), .A3(new_n2625_), .ZN(new_n2674_));
  NAND2_X1   g2625(.A1(new_n2390_), .A2(new_n2546_), .ZN(new_n2675_));
  NAND2_X1   g2626(.A1(new_n2545_), .A2(new_n2675_), .ZN(new_n2676_));
  NOR4_X1    g2627(.A1(new_n2641_), .A2(new_n2475_), .A3(new_n2642_), .A4(new_n2643_), .ZN(new_n2677_));
  AOI22_X1   g2628(.A1(new_n2634_), .A2(new_n2536_), .B1(new_n2639_), .B2(new_n2637_), .ZN(new_n2678_));
  NOR2_X1    g2629(.A1(new_n2677_), .A2(new_n2678_), .ZN(new_n2679_));
  OAI21_X1   g2630(.A1(new_n2540_), .A2(new_n2475_), .B(new_n2481_), .ZN(new_n2680_));
  NAND3_X1   g2631(.A1(new_n2536_), .A2(new_n2482_), .A3(new_n2539_), .ZN(new_n2681_));
  XOR2_X1    g2632(.A1(new_n2651_), .A2(new_n2652_), .Z(new_n2682_));
  NAND3_X1   g2633(.A1(new_n2680_), .A2(new_n2681_), .A3(new_n2682_), .ZN(new_n2683_));
  AOI22_X1   g2634(.A1(new_n2633_), .A2(new_n2631_), .B1(new_n2679_), .B2(new_n2683_), .ZN(new_n2684_));
  AOI21_X1   g2635(.A1(new_n2674_), .A2(new_n2676_), .B(new_n2684_), .ZN(new_n2685_));
  NOR3_X1    g2636(.A1(new_n2685_), .A2(new_n2673_), .A3(new_n2672_), .ZN(new_n2686_));
  NOR2_X1    g2637(.A1(new_n2671_), .A2(new_n2686_), .ZN(new_n2687_));
  NOR2_X1    g2638(.A1(new_n2663_), .A2(new_n2687_), .ZN(new_n2688_));
  NAND2_X1   g2639(.A1(new_n2688_), .A2(new_n2670_), .ZN(new_n2689_));
  NAND2_X1   g2640(.A1(new_n2689_), .A2(new_n2666_), .ZN(new_n2690_));
  NAND3_X1   g2641(.A1(new_n2690_), .A2(new_n2613_), .A3(new_n2667_), .ZN(new_n2691_));
  AOI22_X1   g2642(.A1(new_n2605_), .A2(new_n2606_), .B1(new_n2691_), .B2(new_n2611_), .ZN(new_n2692_));
  OAI22_X1   g2643(.A1(new_n2499_), .A2(new_n2310_), .B1(new_n2300_), .B2(new_n2503_), .ZN(new_n2693_));
  NAND2_X1   g2644(.A1(new_n2693_), .A2(new_n2556_), .ZN(new_n2694_));
  NAND3_X1   g2645(.A1(new_n2518_), .A2(new_n2491_), .A3(new_n2490_), .ZN(new_n2695_));
  OAI21_X1   g2646(.A1(new_n2549_), .A2(new_n2355_), .B(new_n2548_), .ZN(new_n2696_));
  NAND2_X1   g2647(.A1(new_n2622_), .A2(new_n2624_), .ZN(new_n2697_));
  NAND3_X1   g2648(.A1(new_n2660_), .A2(new_n2674_), .A3(new_n2676_), .ZN(new_n2698_));
  NAND2_X1   g2649(.A1(new_n2697_), .A2(new_n2698_), .ZN(new_n2699_));
  NAND3_X1   g2650(.A1(new_n2699_), .A2(new_n2695_), .A3(new_n2696_), .ZN(new_n2700_));
  NAND3_X1   g2651(.A1(new_n2669_), .A2(new_n2700_), .A3(new_n2668_), .ZN(new_n2701_));
  NOR4_X1    g2652(.A1(new_n2551_), .A2(new_n2552_), .A3(new_n2310_), .A4(new_n2498_), .ZN(new_n2702_));
  AOI22_X1   g2653(.A1(new_n2493_), .A2(new_n2494_), .B1(new_n2511_), .B2(new_n2553_), .ZN(new_n2703_));
  NOR2_X1    g2654(.A1(new_n2702_), .A2(new_n2703_), .ZN(new_n2704_));
  AOI22_X1   g2655(.A1(new_n2556_), .A2(new_n2693_), .B1(new_n2704_), .B2(new_n2701_), .ZN(new_n2705_));
  AOI21_X1   g2656(.A1(new_n2688_), .A2(new_n2670_), .B(new_n2704_), .ZN(new_n2706_));
  NOR3_X1    g2657(.A1(new_n2705_), .A2(new_n2706_), .A3(new_n2694_), .ZN(new_n2707_));
  NAND3_X1   g2658(.A1(new_n2610_), .A2(new_n2608_), .A3(new_n2667_), .ZN(new_n2708_));
  NAND3_X1   g2659(.A1(new_n2708_), .A2(new_n2606_), .A3(new_n2605_), .ZN(new_n2709_));
  OAI21_X1   g2660(.A1(new_n2692_), .A2(new_n2604_), .B(new_n2709_), .ZN(new_n2710_));
  NAND3_X1   g2661(.A1(new_n2583_), .A2(new_n2585_), .A3(new_n2595_), .ZN(new_n2711_));
  NAND3_X1   g2662(.A1(new_n2604_), .A2(new_n2597_), .A3(new_n2596_), .ZN(new_n2712_));
  AOI21_X1   g2663(.A1(new_n2711_), .A2(new_n2712_), .B(new_n2710_), .ZN(new_n2713_));
  NOR2_X1    g2664(.A1(new_n2505_), .A2(new_n2609_), .ZN(new_n2714_));
  NOR2_X1    g2665(.A1(new_n2557_), .A2(new_n2607_), .ZN(new_n2715_));
  NOR2_X1    g2666(.A1(new_n2714_), .A2(new_n2715_), .ZN(new_n2716_));
  OAI22_X1   g2667(.A1(new_n2508_), .A2(new_n2562_), .B1(new_n2716_), .B2(new_n2707_), .ZN(new_n2717_));
  AOI22_X1   g2668(.A1(new_n2586_), .A2(new_n2717_), .B1(new_n2563_), .B2(new_n2708_), .ZN(new_n2718_));
  NAND2_X1   g2669(.A1(new_n2712_), .A2(new_n2711_), .ZN(new_n2719_));
  NOR2_X1    g2670(.A1(new_n2719_), .A2(new_n2718_), .ZN(new_n2720_));
  XOR2_X1    g2671(.A1(\a[1] ), .A2(\a[2] ), .Z(new_n2721_));
  AND2_X2    g2672(.A1(new_n2721_), .A2(\a[0] ), .Z(new_n2722_));
  OAI21_X1   g2673(.A1(new_n2720_), .A2(new_n2713_), .B(new_n2722_), .ZN(new_n2723_));
  NAND3_X1   g2674(.A1(new_n2723_), .A2(new_n52_), .A3(new_n2603_), .ZN(new_n2724_));
  INV_X1     g2675(.I(new_n52_), .ZN(new_n2725_));
  INV_X1     g2676(.I(new_n2603_), .ZN(new_n2726_));
  NAND2_X1   g2677(.A1(new_n2719_), .A2(new_n2718_), .ZN(new_n2727_));
  NAND3_X1   g2678(.A1(new_n2710_), .A2(new_n2711_), .A3(new_n2712_), .ZN(new_n2728_));
  INV_X1     g2679(.I(new_n2722_), .ZN(new_n2729_));
  AOI21_X1   g2680(.A1(new_n2727_), .A2(new_n2728_), .B(new_n2729_), .ZN(new_n2730_));
  OAI21_X1   g2681(.A1(new_n2730_), .A2(new_n2726_), .B(new_n2725_), .ZN(new_n2731_));
  NAND2_X1   g2682(.A1(new_n2731_), .A2(new_n2724_), .ZN(new_n2732_));
  XOR2_X1    g2683(.A1(new_n663_), .A2(new_n846_), .Z(new_n2733_));
  XOR2_X1    g2684(.A1(new_n473_), .A2(new_n670_), .Z(new_n2734_));
  NOR2_X1    g2685(.A1(new_n2734_), .A2(new_n2733_), .ZN(new_n2735_));
  INV_X1     g2686(.I(new_n2735_), .ZN(new_n2736_));
  INV_X1     g2687(.I(new_n2733_), .ZN(new_n2737_));
  NOR2_X1    g2688(.A1(new_n2737_), .A2(new_n831_), .ZN(new_n2738_));
  INV_X1     g2689(.I(new_n2738_), .ZN(new_n2739_));
  OAI22_X1   g2690(.A1(new_n2654_), .A2(new_n2736_), .B1(new_n2657_), .B2(new_n2739_), .ZN(new_n2740_));
  INV_X1     g2691(.I(new_n2657_), .ZN(new_n2741_));
  XOR2_X1    g2692(.A1(new_n2654_), .A2(new_n2741_), .Z(new_n2742_));
  NAND2_X1   g2693(.A1(new_n2734_), .A2(new_n2737_), .ZN(new_n2743_));
  NOR2_X1    g2694(.A1(new_n2742_), .A2(new_n2743_), .ZN(new_n2744_));
  NOR2_X1    g2695(.A1(new_n2744_), .A2(new_n2740_), .ZN(new_n2745_));
  NOR2_X1    g2696(.A1(new_n2657_), .A2(new_n2733_), .ZN(new_n2746_));
  INV_X1     g2697(.I(new_n2746_), .ZN(new_n2747_));
  INV_X1     g2698(.I(new_n2743_), .ZN(new_n2748_));
  INV_X1     g2699(.I(new_n753_), .ZN(new_n2749_));
  NAND2_X1   g2700(.A1(new_n474_), .A2(new_n845_), .ZN(new_n2750_));
  NAND2_X1   g2701(.A1(new_n473_), .A2(new_n846_), .ZN(new_n2751_));
  OAI22_X1   g2702(.A1(new_n673_), .A2(new_n2750_), .B1(new_n2749_), .B2(new_n2751_), .ZN(new_n2752_));
  AOI22_X1   g2703(.A1(new_n2682_), .A2(new_n2738_), .B1(new_n2741_), .B2(new_n2752_), .ZN(new_n2753_));
  NOR2_X1    g2704(.A1(new_n2647_), .A2(new_n2646_), .ZN(new_n2754_));
  NAND2_X1   g2705(.A1(new_n2754_), .A2(new_n2735_), .ZN(new_n2755_));
  NAND2_X1   g2706(.A1(new_n2755_), .A2(new_n2753_), .ZN(new_n2756_));
  NAND2_X1   g2707(.A1(new_n2680_), .A2(new_n2681_), .ZN(new_n2757_));
  NAND2_X1   g2708(.A1(new_n2682_), .A2(new_n2657_), .ZN(new_n2758_));
  NOR2_X1    g2709(.A1(new_n2757_), .A2(new_n2758_), .ZN(new_n2759_));
  NOR2_X1    g2710(.A1(new_n2654_), .A2(new_n2741_), .ZN(new_n2760_));
  AOI21_X1   g2711(.A1(new_n2680_), .A2(new_n2681_), .B(new_n2760_), .ZN(new_n2761_));
  NOR2_X1    g2712(.A1(new_n2759_), .A2(new_n2761_), .ZN(new_n2762_));
  AOI21_X1   g2713(.A1(new_n2762_), .A2(new_n2748_), .B(new_n2756_), .ZN(new_n2763_));
  NAND4_X1   g2714(.A1(new_n2763_), .A2(new_n473_), .A3(new_n2745_), .A4(new_n2747_), .ZN(new_n2764_));
  NOR2_X1    g2715(.A1(new_n2657_), .A2(new_n631_), .ZN(new_n2765_));
  INV_X1     g2716(.I(new_n2765_), .ZN(new_n2766_));
  NOR2_X1    g2717(.A1(new_n2764_), .A2(new_n2766_), .ZN(new_n2767_));
  INV_X1     g2718(.I(new_n2752_), .ZN(new_n2768_));
  OAI22_X1   g2719(.A1(new_n2757_), .A2(new_n2739_), .B1(new_n2654_), .B2(new_n2768_), .ZN(new_n2769_));
  AOI21_X1   g2720(.A1(new_n2645_), .A2(new_n2735_), .B(new_n2769_), .ZN(new_n2770_));
  NAND3_X1   g2721(.A1(new_n2645_), .A2(new_n2658_), .A3(new_n2683_), .ZN(new_n2771_));
  NAND2_X1   g2722(.A1(new_n2658_), .A2(new_n2683_), .ZN(new_n2772_));
  NAND2_X1   g2723(.A1(new_n2772_), .A2(new_n2679_), .ZN(new_n2773_));
  NAND3_X1   g2724(.A1(new_n2773_), .A2(new_n2771_), .A3(new_n2748_), .ZN(new_n2774_));
  AOI21_X1   g2725(.A1(new_n2774_), .A2(new_n2770_), .B(new_n473_), .ZN(new_n2775_));
  INV_X1     g2726(.I(new_n2775_), .ZN(new_n2776_));
  NAND3_X1   g2727(.A1(new_n2774_), .A2(new_n473_), .A3(new_n2770_), .ZN(new_n2777_));
  NAND2_X1   g2728(.A1(new_n2764_), .A2(new_n2765_), .ZN(new_n2778_));
  INV_X1     g2729(.I(new_n2745_), .ZN(new_n2779_));
  NAND3_X1   g2730(.A1(new_n2760_), .A2(new_n2680_), .A3(new_n2681_), .ZN(new_n2780_));
  NAND2_X1   g2731(.A1(new_n2757_), .A2(new_n2758_), .ZN(new_n2781_));
  NAND3_X1   g2732(.A1(new_n2781_), .A2(new_n2748_), .A3(new_n2780_), .ZN(new_n2782_));
  NAND3_X1   g2733(.A1(new_n2782_), .A2(new_n2753_), .A3(new_n2755_), .ZN(new_n2783_));
  NOR4_X1    g2734(.A1(new_n2779_), .A2(new_n2783_), .A3(new_n474_), .A4(new_n2746_), .ZN(new_n2784_));
  NAND2_X1   g2735(.A1(new_n2784_), .A2(new_n2766_), .ZN(new_n2785_));
  AOI22_X1   g2736(.A1(new_n2785_), .A2(new_n2778_), .B1(new_n2776_), .B2(new_n2777_), .ZN(new_n2786_));
  NOR2_X1    g2737(.A1(new_n2786_), .A2(new_n2767_), .ZN(new_n2787_));
  OAI22_X1   g2738(.A1(new_n2679_), .A2(new_n2739_), .B1(new_n2757_), .B2(new_n2768_), .ZN(new_n2788_));
  NOR2_X1    g2739(.A1(new_n2632_), .A2(new_n2543_), .ZN(new_n2789_));
  NOR2_X1    g2740(.A1(new_n2486_), .A2(new_n2527_), .ZN(new_n2790_));
  NOR2_X1    g2741(.A1(new_n2790_), .A2(new_n2485_), .ZN(new_n2791_));
  NOR2_X1    g2742(.A1(new_n2789_), .A2(new_n2791_), .ZN(new_n2792_));
  NOR2_X1    g2743(.A1(new_n2792_), .A2(new_n2736_), .ZN(new_n2793_));
  NOR2_X1    g2744(.A1(new_n2793_), .A2(new_n2788_), .ZN(new_n2794_));
  INV_X1     g2745(.I(new_n2794_), .ZN(new_n2795_));
  NOR3_X1    g2746(.A1(new_n2645_), .A2(new_n2757_), .A3(new_n2654_), .ZN(new_n2796_));
  AOI21_X1   g2747(.A1(new_n2757_), .A2(new_n2657_), .B(new_n2654_), .ZN(new_n2797_));
  NOR3_X1    g2748(.A1(new_n2797_), .A2(new_n2679_), .A3(new_n2754_), .ZN(new_n2798_));
  OAI21_X1   g2749(.A1(new_n2796_), .A2(new_n2798_), .B(new_n2792_), .ZN(new_n2799_));
  NAND2_X1   g2750(.A1(new_n2633_), .A2(new_n2631_), .ZN(new_n2800_));
  NAND3_X1   g2751(.A1(new_n2679_), .A2(new_n2754_), .A3(new_n2682_), .ZN(new_n2801_));
  OAI21_X1   g2752(.A1(new_n2754_), .A2(new_n2741_), .B(new_n2682_), .ZN(new_n2802_));
  NAND3_X1   g2753(.A1(new_n2802_), .A2(new_n2645_), .A3(new_n2757_), .ZN(new_n2803_));
  NAND3_X1   g2754(.A1(new_n2800_), .A2(new_n2803_), .A3(new_n2801_), .ZN(new_n2804_));
  AOI21_X1   g2755(.A1(new_n2799_), .A2(new_n2804_), .B(new_n2743_), .ZN(new_n2805_));
  OAI21_X1   g2756(.A1(new_n2795_), .A2(new_n2805_), .B(new_n474_), .ZN(new_n2806_));
  AOI21_X1   g2757(.A1(new_n2801_), .A2(new_n2803_), .B(new_n2800_), .ZN(new_n2807_));
  NOR3_X1    g2758(.A1(new_n2792_), .A2(new_n2798_), .A3(new_n2796_), .ZN(new_n2808_));
  OAI21_X1   g2759(.A1(new_n2807_), .A2(new_n2808_), .B(new_n2748_), .ZN(new_n2809_));
  NAND3_X1   g2760(.A1(new_n2809_), .A2(new_n473_), .A3(new_n2794_), .ZN(new_n2810_));
  NAND2_X1   g2761(.A1(new_n2806_), .A2(new_n2810_), .ZN(new_n2811_));
  NOR2_X1    g2762(.A1(new_n631_), .A2(new_n466_), .ZN(new_n2812_));
  NOR2_X1    g2763(.A1(new_n477_), .A2(new_n473_), .ZN(new_n2813_));
  NOR2_X1    g2764(.A1(new_n480_), .A2(new_n462_), .ZN(new_n2814_));
  AOI21_X1   g2765(.A1(new_n462_), .A2(new_n2813_), .B(new_n2814_), .ZN(new_n2815_));
  INV_X1     g2766(.I(new_n2815_), .ZN(new_n2816_));
  AOI22_X1   g2767(.A1(new_n2682_), .A2(new_n2812_), .B1(new_n2741_), .B2(new_n2816_), .ZN(new_n2817_));
  INV_X1     g2768(.I(new_n466_), .ZN(new_n2818_));
  NOR2_X1    g2769(.A1(new_n631_), .A2(new_n2818_), .ZN(new_n2819_));
  INV_X1     g2770(.I(new_n2819_), .ZN(new_n2820_));
  OAI21_X1   g2771(.A1(new_n2742_), .A2(new_n2820_), .B(new_n2817_), .ZN(new_n2821_));
  NAND2_X1   g2772(.A1(new_n2821_), .A2(new_n465_), .ZN(new_n2822_));
  INV_X1     g2773(.I(new_n2821_), .ZN(new_n2823_));
  NAND2_X1   g2774(.A1(new_n2823_), .A2(new_n598_), .ZN(new_n2824_));
  NAND2_X1   g2775(.A1(new_n2824_), .A2(new_n2822_), .ZN(new_n2825_));
  NOR2_X1    g2776(.A1(new_n2765_), .A2(new_n598_), .ZN(new_n2826_));
  OAI22_X1   g2777(.A1(new_n2825_), .A2(new_n2826_), .B1(new_n2765_), .B2(new_n2822_), .ZN(new_n2827_));
  INV_X1     g2778(.I(new_n2827_), .ZN(new_n2828_));
  NOR2_X1    g2779(.A1(new_n2811_), .A2(new_n2828_), .ZN(new_n2829_));
  AOI21_X1   g2780(.A1(new_n2809_), .A2(new_n2794_), .B(new_n473_), .ZN(new_n2830_));
  NOR3_X1    g2781(.A1(new_n2795_), .A2(new_n2805_), .A3(new_n474_), .ZN(new_n2831_));
  NOR2_X1    g2782(.A1(new_n2831_), .A2(new_n2830_), .ZN(new_n2832_));
  NOR2_X1    g2783(.A1(new_n2832_), .A2(new_n2827_), .ZN(new_n2833_));
  NOR3_X1    g2784(.A1(new_n2833_), .A2(new_n2829_), .A3(new_n2787_), .ZN(new_n2834_));
  INV_X1     g2785(.I(new_n2767_), .ZN(new_n2835_));
  INV_X1     g2786(.I(new_n2777_), .ZN(new_n2836_));
  NOR2_X1    g2787(.A1(new_n2784_), .A2(new_n2766_), .ZN(new_n2837_));
  NOR2_X1    g2788(.A1(new_n2764_), .A2(new_n2765_), .ZN(new_n2838_));
  OAI22_X1   g2789(.A1(new_n2837_), .A2(new_n2838_), .B1(new_n2836_), .B2(new_n2775_), .ZN(new_n2839_));
  NAND2_X1   g2790(.A1(new_n2839_), .A2(new_n2835_), .ZN(new_n2840_));
  NAND2_X1   g2791(.A1(new_n2832_), .A2(new_n2827_), .ZN(new_n2841_));
  NAND2_X1   g2792(.A1(new_n2811_), .A2(new_n2828_), .ZN(new_n2842_));
  AOI21_X1   g2793(.A1(new_n2841_), .A2(new_n2842_), .B(new_n2840_), .ZN(new_n2843_));
  OR2_X2     g2794(.A1(new_n2843_), .A2(new_n2834_), .Z(new_n2844_));
  NAND2_X1   g2795(.A1(new_n2674_), .A2(new_n2676_), .ZN(new_n2845_));
  NOR2_X1    g2796(.A1(new_n1161_), .A2(new_n1288_), .ZN(new_n2846_));
  NOR2_X1    g2797(.A1(new_n1162_), .A2(new_n1287_), .ZN(new_n2847_));
  NOR2_X1    g2798(.A1(new_n2847_), .A2(new_n2846_), .ZN(new_n2848_));
  INV_X1     g2799(.I(new_n2848_), .ZN(new_n2849_));
  XNOR2_X1   g2800(.A1(new_n842_), .A2(new_n1287_), .ZN(new_n2850_));
  NOR2_X1    g2801(.A1(new_n2849_), .A2(new_n2850_), .ZN(new_n2851_));
  INV_X1     g2802(.I(new_n2851_), .ZN(new_n2852_));
  NOR2_X1    g2803(.A1(new_n1052_), .A2(new_n1287_), .ZN(new_n2853_));
  NOR2_X1    g2804(.A1(new_n1051_), .A2(new_n1288_), .ZN(new_n2854_));
  NOR3_X1    g2805(.A1(new_n2849_), .A2(new_n2854_), .A3(new_n2853_), .ZN(new_n2855_));
  INV_X1     g2806(.I(new_n2855_), .ZN(new_n2856_));
  OAI22_X1   g2807(.A1(new_n2697_), .A2(new_n2852_), .B1(new_n2845_), .B2(new_n2856_), .ZN(new_n2857_));
  NAND2_X1   g2808(.A1(new_n2696_), .A2(new_n2695_), .ZN(new_n2858_));
  NOR2_X1    g2809(.A1(new_n2848_), .A2(new_n1056_), .ZN(new_n2859_));
  INV_X1     g2810(.I(new_n2859_), .ZN(new_n2860_));
  NOR2_X1    g2811(.A1(new_n2858_), .A2(new_n2860_), .ZN(new_n2861_));
  NOR2_X1    g2812(.A1(new_n2861_), .A2(new_n2857_), .ZN(new_n2862_));
  NOR2_X1    g2813(.A1(new_n2848_), .A2(new_n1053_), .ZN(new_n2863_));
  NOR2_X1    g2814(.A1(new_n2686_), .A2(new_n2661_), .ZN(new_n2864_));
  NAND2_X1   g2815(.A1(new_n2864_), .A2(new_n2858_), .ZN(new_n2865_));
  NOR3_X1    g2816(.A1(new_n2647_), .A2(new_n2646_), .A3(new_n2654_), .ZN(new_n2866_));
  OAI22_X1   g2817(.A1(new_n2789_), .A2(new_n2791_), .B1(new_n2645_), .B2(new_n2866_), .ZN(new_n2867_));
  OAI21_X1   g2818(.A1(new_n2627_), .A2(new_n2629_), .B(new_n2867_), .ZN(new_n2868_));
  NAND3_X1   g2819(.A1(new_n2868_), .A2(new_n2622_), .A3(new_n2624_), .ZN(new_n2869_));
  NAND2_X1   g2820(.A1(new_n2699_), .A2(new_n2869_), .ZN(new_n2870_));
  NAND2_X1   g2821(.A1(new_n2870_), .A2(new_n2671_), .ZN(new_n2871_));
  NAND2_X1   g2822(.A1(new_n2871_), .A2(new_n2865_), .ZN(new_n2872_));
  NAND2_X1   g2823(.A1(new_n2872_), .A2(new_n2863_), .ZN(new_n2873_));
  AOI21_X1   g2824(.A1(new_n2873_), .A2(new_n2862_), .B(new_n846_), .ZN(new_n2874_));
  INV_X1     g2825(.I(new_n2874_), .ZN(new_n2875_));
  NAND3_X1   g2826(.A1(new_n2873_), .A2(new_n846_), .A3(new_n2862_), .ZN(new_n2876_));
  AOI21_X1   g2827(.A1(new_n2875_), .A2(new_n2876_), .B(new_n2844_), .ZN(new_n2877_));
  AOI22_X1   g2828(.A1(new_n2630_), .A2(new_n2851_), .B1(new_n2800_), .B2(new_n2855_), .ZN(new_n2878_));
  OAI21_X1   g2829(.A1(new_n2697_), .A2(new_n2860_), .B(new_n2878_), .ZN(new_n2879_));
  INV_X1     g2830(.I(new_n2863_), .ZN(new_n2880_));
  NOR2_X1    g2831(.A1(new_n2673_), .A2(new_n2672_), .ZN(new_n2881_));
  NAND2_X1   g2832(.A1(new_n2868_), .A2(new_n2698_), .ZN(new_n2882_));
  NAND2_X1   g2833(.A1(new_n2882_), .A2(new_n2881_), .ZN(new_n2883_));
  NAND3_X1   g2834(.A1(new_n2697_), .A2(new_n2698_), .A3(new_n2868_), .ZN(new_n2884_));
  AOI21_X1   g2835(.A1(new_n2883_), .A2(new_n2884_), .B(new_n2880_), .ZN(new_n2885_));
  OAI21_X1   g2836(.A1(new_n2885_), .A2(new_n2879_), .B(new_n846_), .ZN(new_n2886_));
  INV_X1     g2837(.I(new_n2886_), .ZN(new_n2887_));
  NOR3_X1    g2838(.A1(new_n2885_), .A2(new_n2879_), .A3(new_n846_), .ZN(new_n2888_));
  NOR4_X1    g2839(.A1(new_n2837_), .A2(new_n2838_), .A3(new_n2836_), .A4(new_n2775_), .ZN(new_n2889_));
  NOR2_X1    g2840(.A1(new_n2786_), .A2(new_n2889_), .ZN(new_n2890_));
  NOR3_X1    g2841(.A1(new_n2887_), .A2(new_n2888_), .A3(new_n2890_), .ZN(new_n2891_));
  INV_X1     g2842(.I(new_n2891_), .ZN(new_n2892_));
  OAI22_X1   g2843(.A1(new_n2792_), .A2(new_n2852_), .B1(new_n2679_), .B2(new_n2856_), .ZN(new_n2893_));
  NOR2_X1    g2844(.A1(new_n2845_), .A2(new_n2860_), .ZN(new_n2894_));
  NOR2_X1    g2845(.A1(new_n2894_), .A2(new_n2893_), .ZN(new_n2895_));
  INV_X1     g2846(.I(new_n2895_), .ZN(new_n2896_));
  AOI22_X1   g2847(.A1(new_n2680_), .A2(new_n2681_), .B1(new_n2682_), .B2(new_n2741_), .ZN(new_n2897_));
  AOI21_X1   g2848(.A1(new_n2640_), .A2(new_n2644_), .B(new_n2897_), .ZN(new_n2898_));
  NOR3_X1    g2849(.A1(new_n2898_), .A2(new_n2789_), .A3(new_n2791_), .ZN(new_n2899_));
  NOR2_X1    g2850(.A1(new_n2899_), .A2(new_n2684_), .ZN(new_n2900_));
  NAND2_X1   g2851(.A1(new_n2900_), .A2(new_n2845_), .ZN(new_n2901_));
  OAI21_X1   g2852(.A1(new_n2899_), .A2(new_n2684_), .B(new_n2630_), .ZN(new_n2902_));
  AOI21_X1   g2853(.A1(new_n2902_), .A2(new_n2901_), .B(new_n2880_), .ZN(new_n2903_));
  OAI21_X1   g2854(.A1(new_n2896_), .A2(new_n2903_), .B(new_n845_), .ZN(new_n2904_));
  NOR3_X1    g2855(.A1(new_n2896_), .A2(new_n2903_), .A3(new_n845_), .ZN(new_n2905_));
  INV_X1     g2856(.I(new_n2905_), .ZN(new_n2906_));
  NAND3_X1   g2857(.A1(new_n2745_), .A2(new_n473_), .A3(new_n2747_), .ZN(new_n2907_));
  INV_X1     g2858(.I(new_n2907_), .ZN(new_n2908_));
  XOR2_X1    g2859(.A1(new_n2783_), .A2(new_n473_), .Z(new_n2909_));
  NOR2_X1    g2860(.A1(new_n2909_), .A2(new_n2908_), .ZN(new_n2910_));
  NOR2_X1    g2861(.A1(new_n2910_), .A2(new_n2784_), .ZN(new_n2911_));
  AOI21_X1   g2862(.A1(new_n2906_), .A2(new_n2904_), .B(new_n2911_), .ZN(new_n2912_));
  AOI22_X1   g2863(.A1(new_n2645_), .A2(new_n2851_), .B1(new_n2754_), .B2(new_n2855_), .ZN(new_n2913_));
  OAI21_X1   g2864(.A1(new_n2792_), .A2(new_n2860_), .B(new_n2913_), .ZN(new_n2914_));
  AOI21_X1   g2865(.A1(new_n2799_), .A2(new_n2804_), .B(new_n2880_), .ZN(new_n2915_));
  OAI21_X1   g2866(.A1(new_n2915_), .A2(new_n2914_), .B(new_n846_), .ZN(new_n2916_));
  NOR3_X1    g2867(.A1(new_n2915_), .A2(new_n846_), .A3(new_n2914_), .ZN(new_n2917_));
  INV_X1     g2868(.I(new_n2917_), .ZN(new_n2918_));
  XOR2_X1    g2869(.A1(new_n2745_), .A2(new_n473_), .Z(new_n2919_));
  NOR2_X1    g2870(.A1(new_n2746_), .A2(new_n474_), .ZN(new_n2920_));
  INV_X1     g2871(.I(new_n2920_), .ZN(new_n2921_));
  NAND2_X1   g2872(.A1(new_n2919_), .A2(new_n2921_), .ZN(new_n2922_));
  NAND2_X1   g2873(.A1(new_n2922_), .A2(new_n2907_), .ZN(new_n2923_));
  NAND3_X1   g2874(.A1(new_n2918_), .A2(new_n2923_), .A3(new_n2916_), .ZN(new_n2924_));
  AOI21_X1   g2875(.A1(new_n2918_), .A2(new_n2916_), .B(new_n2923_), .ZN(new_n2925_));
  OAI22_X1   g2876(.A1(new_n2757_), .A2(new_n2852_), .B1(new_n2654_), .B2(new_n2856_), .ZN(new_n2926_));
  AOI21_X1   g2877(.A1(new_n2645_), .A2(new_n2859_), .B(new_n2926_), .ZN(new_n2927_));
  INV_X1     g2878(.I(new_n2927_), .ZN(new_n2928_));
  NOR3_X1    g2879(.A1(new_n2679_), .A2(new_n2897_), .A3(new_n2866_), .ZN(new_n2929_));
  NOR2_X1    g2880(.A1(new_n2897_), .A2(new_n2866_), .ZN(new_n2930_));
  NOR2_X1    g2881(.A1(new_n2930_), .A2(new_n2645_), .ZN(new_n2931_));
  NOR3_X1    g2882(.A1(new_n2931_), .A2(new_n2929_), .A3(new_n2880_), .ZN(new_n2932_));
  OAI21_X1   g2883(.A1(new_n2928_), .A2(new_n2932_), .B(new_n845_), .ZN(new_n2933_));
  NAND3_X1   g2884(.A1(new_n2773_), .A2(new_n2771_), .A3(new_n2863_), .ZN(new_n2934_));
  NAND3_X1   g2885(.A1(new_n2934_), .A2(new_n846_), .A3(new_n2927_), .ZN(new_n2935_));
  AOI21_X1   g2886(.A1(new_n2933_), .A2(new_n2935_), .B(new_n2746_), .ZN(new_n2936_));
  NAND2_X1   g2887(.A1(new_n2781_), .A2(new_n2780_), .ZN(new_n2937_));
  OAI22_X1   g2888(.A1(new_n2654_), .A2(new_n2852_), .B1(new_n2657_), .B2(new_n2856_), .ZN(new_n2938_));
  AOI21_X1   g2889(.A1(new_n2754_), .A2(new_n2859_), .B(new_n2938_), .ZN(new_n2939_));
  OAI21_X1   g2890(.A1(new_n2937_), .A2(new_n2880_), .B(new_n2939_), .ZN(new_n2940_));
  AOI22_X1   g2891(.A1(new_n2682_), .A2(new_n2859_), .B1(new_n2741_), .B2(new_n2851_), .ZN(new_n2941_));
  OAI21_X1   g2892(.A1(new_n2742_), .A2(new_n2880_), .B(new_n2941_), .ZN(new_n2942_));
  NOR2_X1    g2893(.A1(new_n2657_), .A2(new_n2848_), .ZN(new_n2943_));
  NOR4_X1    g2894(.A1(new_n2940_), .A2(new_n846_), .A3(new_n2942_), .A4(new_n2943_), .ZN(new_n2944_));
  INV_X1     g2895(.I(new_n2944_), .ZN(new_n2945_));
  NAND3_X1   g2896(.A1(new_n2933_), .A2(new_n2935_), .A3(new_n2746_), .ZN(new_n2946_));
  AOI21_X1   g2897(.A1(new_n2945_), .A2(new_n2946_), .B(new_n2936_), .ZN(new_n2947_));
  OAI21_X1   g2898(.A1(new_n2925_), .A2(new_n2947_), .B(new_n2924_), .ZN(new_n2948_));
  NAND3_X1   g2899(.A1(new_n2906_), .A2(new_n2904_), .A3(new_n2911_), .ZN(new_n2949_));
  AOI21_X1   g2900(.A1(new_n2948_), .A2(new_n2949_), .B(new_n2912_), .ZN(new_n2950_));
  OAI21_X1   g2901(.A1(new_n2887_), .A2(new_n2888_), .B(new_n2890_), .ZN(new_n2951_));
  INV_X1     g2902(.I(new_n2951_), .ZN(new_n2952_));
  OAI21_X1   g2903(.A1(new_n2950_), .A2(new_n2952_), .B(new_n2892_), .ZN(new_n2953_));
  NAND3_X1   g2904(.A1(new_n2844_), .A2(new_n2875_), .A3(new_n2876_), .ZN(new_n2954_));
  AOI21_X1   g2905(.A1(new_n2953_), .A2(new_n2954_), .B(new_n2877_), .ZN(new_n2955_));
  NOR2_X1    g2906(.A1(new_n2617_), .A2(new_n2618_), .ZN(new_n2956_));
  NOR2_X1    g2907(.A1(new_n2956_), .A2(new_n2860_), .ZN(new_n2957_));
  NOR2_X1    g2908(.A1(new_n2697_), .A2(new_n2856_), .ZN(new_n2958_));
  NOR2_X1    g2909(.A1(new_n2858_), .A2(new_n2852_), .ZN(new_n2959_));
  NOR3_X1    g2910(.A1(new_n2957_), .A2(new_n2958_), .A3(new_n2959_), .ZN(new_n2960_));
  INV_X1     g2911(.I(new_n2960_), .ZN(new_n2961_));
  OAI21_X1   g2912(.A1(new_n2617_), .A2(new_n2618_), .B(new_n2881_), .ZN(new_n2962_));
  NAND3_X1   g2913(.A1(new_n2669_), .A2(new_n2668_), .A3(new_n2869_), .ZN(new_n2963_));
  NAND3_X1   g2914(.A1(new_n2962_), .A2(new_n2963_), .A3(new_n2858_), .ZN(new_n2964_));
  NAND2_X1   g2915(.A1(new_n2699_), .A2(new_n2868_), .ZN(new_n2965_));
  NAND4_X1   g2916(.A1(new_n2669_), .A2(new_n2965_), .A3(new_n2668_), .A4(new_n2697_), .ZN(new_n2966_));
  NAND2_X1   g2917(.A1(new_n2962_), .A2(new_n2966_), .ZN(new_n2967_));
  AOI22_X1   g2918(.A1(new_n2967_), .A2(new_n2671_), .B1(new_n2670_), .B2(new_n2864_), .ZN(new_n2968_));
  AOI21_X1   g2919(.A1(new_n2968_), .A2(new_n2964_), .B(new_n2880_), .ZN(new_n2969_));
  OAI21_X1   g2920(.A1(new_n2969_), .A2(new_n2961_), .B(new_n846_), .ZN(new_n2970_));
  AOI21_X1   g2921(.A1(new_n2669_), .A2(new_n2668_), .B(new_n2697_), .ZN(new_n2971_));
  NOR2_X1    g2922(.A1(new_n2661_), .A2(new_n2685_), .ZN(new_n2972_));
  NOR4_X1    g2923(.A1(new_n2617_), .A2(new_n2618_), .A3(new_n2881_), .A4(new_n2972_), .ZN(new_n2973_));
  OAI21_X1   g2924(.A1(new_n2973_), .A2(new_n2971_), .B(new_n2671_), .ZN(new_n2974_));
  NAND2_X1   g2925(.A1(new_n2670_), .A2(new_n2864_), .ZN(new_n2975_));
  NAND3_X1   g2926(.A1(new_n2974_), .A2(new_n2964_), .A3(new_n2975_), .ZN(new_n2976_));
  NAND2_X1   g2927(.A1(new_n2976_), .A2(new_n2863_), .ZN(new_n2977_));
  NAND3_X1   g2928(.A1(new_n2977_), .A2(new_n845_), .A3(new_n2960_), .ZN(new_n2978_));
  NAND3_X1   g2929(.A1(new_n2839_), .A2(new_n2835_), .A3(new_n2828_), .ZN(new_n2979_));
  OAI21_X1   g2930(.A1(new_n2786_), .A2(new_n2767_), .B(new_n2827_), .ZN(new_n2980_));
  NAND2_X1   g2931(.A1(new_n2980_), .A2(new_n2832_), .ZN(new_n2981_));
  OAI22_X1   g2932(.A1(new_n2792_), .A2(new_n2739_), .B1(new_n2679_), .B2(new_n2768_), .ZN(new_n2982_));
  NOR2_X1    g2933(.A1(new_n2845_), .A2(new_n2736_), .ZN(new_n2983_));
  NOR2_X1    g2934(.A1(new_n2983_), .A2(new_n2982_), .ZN(new_n2984_));
  INV_X1     g2935(.I(new_n2984_), .ZN(new_n2985_));
  AOI21_X1   g2936(.A1(new_n2902_), .A2(new_n2901_), .B(new_n2743_), .ZN(new_n2986_));
  OAI21_X1   g2937(.A1(new_n2985_), .A2(new_n2986_), .B(new_n474_), .ZN(new_n2987_));
  NOR3_X1    g2938(.A1(new_n2630_), .A2(new_n2899_), .A3(new_n2684_), .ZN(new_n2988_));
  NOR2_X1    g2939(.A1(new_n2900_), .A2(new_n2845_), .ZN(new_n2989_));
  OAI21_X1   g2940(.A1(new_n2989_), .A2(new_n2988_), .B(new_n2748_), .ZN(new_n2990_));
  NAND3_X1   g2941(.A1(new_n2990_), .A2(new_n473_), .A3(new_n2984_), .ZN(new_n2991_));
  NAND2_X1   g2942(.A1(new_n2987_), .A2(new_n2991_), .ZN(new_n2992_));
  NAND3_X1   g2943(.A1(new_n2981_), .A2(new_n2979_), .A3(new_n2992_), .ZN(new_n2993_));
  AOI21_X1   g2944(.A1(new_n2839_), .A2(new_n2835_), .B(new_n2828_), .ZN(new_n2994_));
  OAI21_X1   g2945(.A1(new_n2811_), .A2(new_n2994_), .B(new_n2979_), .ZN(new_n2995_));
  INV_X1     g2946(.I(new_n2992_), .ZN(new_n2996_));
  NAND2_X1   g2947(.A1(new_n2995_), .A2(new_n2996_), .ZN(new_n2997_));
  NOR2_X1    g2948(.A1(new_n2813_), .A2(new_n598_), .ZN(new_n2998_));
  NOR2_X1    g2949(.A1(new_n479_), .A2(new_n465_), .ZN(new_n2999_));
  NOR3_X1    g2950(.A1(new_n2999_), .A2(new_n2818_), .A3(new_n2998_), .ZN(new_n3000_));
  INV_X1     g2951(.I(new_n3000_), .ZN(new_n3001_));
  OAI22_X1   g2952(.A1(new_n2654_), .A2(new_n2815_), .B1(new_n2657_), .B2(new_n3001_), .ZN(new_n3002_));
  INV_X1     g2953(.I(new_n2812_), .ZN(new_n3003_));
  NOR2_X1    g2954(.A1(new_n2757_), .A2(new_n3003_), .ZN(new_n3004_));
  NOR2_X1    g2955(.A1(new_n3004_), .A2(new_n3002_), .ZN(new_n3005_));
  OAI21_X1   g2956(.A1(new_n2937_), .A2(new_n2820_), .B(new_n3005_), .ZN(new_n3006_));
  NOR4_X1    g2957(.A1(new_n3006_), .A2(new_n598_), .A3(new_n2765_), .A4(new_n2821_), .ZN(new_n3007_));
  XOR2_X1    g2958(.A1(new_n3006_), .A2(new_n465_), .Z(new_n3008_));
  NOR3_X1    g2959(.A1(new_n2821_), .A2(new_n598_), .A3(new_n2765_), .ZN(new_n3009_));
  NOR2_X1    g2960(.A1(new_n3008_), .A2(new_n3009_), .ZN(new_n3010_));
  NOR2_X1    g2961(.A1(new_n3010_), .A2(new_n3007_), .ZN(new_n3011_));
  INV_X1     g2962(.I(new_n3011_), .ZN(new_n3012_));
  AOI21_X1   g2963(.A1(new_n2997_), .A2(new_n2993_), .B(new_n3012_), .ZN(new_n3013_));
  NOR2_X1    g2964(.A1(new_n2995_), .A2(new_n2996_), .ZN(new_n3014_));
  NOR3_X1    g2965(.A1(new_n2786_), .A2(new_n2767_), .A3(new_n2827_), .ZN(new_n3015_));
  AOI21_X1   g2966(.A1(new_n2832_), .A2(new_n2980_), .B(new_n3015_), .ZN(new_n3016_));
  NOR2_X1    g2967(.A1(new_n3016_), .A2(new_n2992_), .ZN(new_n3017_));
  NOR3_X1    g2968(.A1(new_n3017_), .A2(new_n3014_), .A3(new_n3011_), .ZN(new_n3018_));
  NOR2_X1    g2969(.A1(new_n3018_), .A2(new_n3013_), .ZN(new_n3019_));
  NAND3_X1   g2970(.A1(new_n2970_), .A2(new_n3019_), .A3(new_n2978_), .ZN(new_n3020_));
  AOI21_X1   g2971(.A1(new_n2977_), .A2(new_n2960_), .B(new_n845_), .ZN(new_n3021_));
  NOR3_X1    g2972(.A1(new_n2969_), .A2(new_n846_), .A3(new_n2961_), .ZN(new_n3022_));
  OAI21_X1   g2973(.A1(new_n3017_), .A2(new_n3014_), .B(new_n3011_), .ZN(new_n3023_));
  NAND3_X1   g2974(.A1(new_n2997_), .A2(new_n2993_), .A3(new_n3012_), .ZN(new_n3024_));
  NAND2_X1   g2975(.A1(new_n3023_), .A2(new_n3024_), .ZN(new_n3025_));
  OAI21_X1   g2976(.A1(new_n3022_), .A2(new_n3021_), .B(new_n3025_), .ZN(new_n3026_));
  NAND3_X1   g2977(.A1(new_n2955_), .A2(new_n3026_), .A3(new_n3020_), .ZN(new_n3027_));
  NOR2_X1    g2978(.A1(new_n2843_), .A2(new_n2834_), .ZN(new_n3028_));
  INV_X1     g2979(.I(new_n2876_), .ZN(new_n3029_));
  OAI21_X1   g2980(.A1(new_n3029_), .A2(new_n2874_), .B(new_n3028_), .ZN(new_n3030_));
  INV_X1     g2981(.I(new_n2904_), .ZN(new_n3031_));
  INV_X1     g2982(.I(new_n2911_), .ZN(new_n3032_));
  OAI21_X1   g2983(.A1(new_n3031_), .A2(new_n2905_), .B(new_n3032_), .ZN(new_n3033_));
  INV_X1     g2984(.I(new_n2916_), .ZN(new_n3034_));
  INV_X1     g2985(.I(new_n2923_), .ZN(new_n3035_));
  NOR3_X1    g2986(.A1(new_n3035_), .A2(new_n3034_), .A3(new_n2917_), .ZN(new_n3036_));
  INV_X1     g2987(.I(new_n2925_), .ZN(new_n3037_));
  INV_X1     g2988(.I(new_n2947_), .ZN(new_n3038_));
  AOI21_X1   g2989(.A1(new_n3037_), .A2(new_n3038_), .B(new_n3036_), .ZN(new_n3039_));
  NOR3_X1    g2990(.A1(new_n3031_), .A2(new_n3032_), .A3(new_n2905_), .ZN(new_n3040_));
  OAI21_X1   g2991(.A1(new_n3039_), .A2(new_n3040_), .B(new_n3033_), .ZN(new_n3041_));
  AOI21_X1   g2992(.A1(new_n3041_), .A2(new_n2951_), .B(new_n2891_), .ZN(new_n3042_));
  NOR3_X1    g2993(.A1(new_n3029_), .A2(new_n3028_), .A3(new_n2874_), .ZN(new_n3043_));
  OAI21_X1   g2994(.A1(new_n3042_), .A2(new_n3043_), .B(new_n3030_), .ZN(new_n3044_));
  NOR3_X1    g2995(.A1(new_n3022_), .A2(new_n3025_), .A3(new_n3021_), .ZN(new_n3045_));
  AOI21_X1   g2996(.A1(new_n2970_), .A2(new_n2978_), .B(new_n3019_), .ZN(new_n3046_));
  OAI21_X1   g2997(.A1(new_n3046_), .A2(new_n3045_), .B(new_n3044_), .ZN(new_n3047_));
  AND2_X2    g2998(.A1(new_n3027_), .A2(new_n3047_), .Z(new_n3048_));
  NOR2_X1    g2999(.A1(new_n1453_), .A2(new_n2725_), .ZN(new_n3049_));
  NOR3_X1    g3000(.A1(new_n1360_), .A2(new_n52_), .A3(new_n1452_), .ZN(new_n3050_));
  AOI21_X1   g3001(.A1(new_n1360_), .A2(new_n3049_), .B(new_n3050_), .ZN(new_n3051_));
  XOR2_X1    g3002(.A1(new_n1287_), .A2(new_n1359_), .Z(new_n3052_));
  INV_X1     g3003(.I(new_n3052_), .ZN(new_n3053_));
  NOR2_X1    g3004(.A1(new_n3049_), .A2(new_n1360_), .ZN(new_n3054_));
  AOI21_X1   g3005(.A1(new_n1453_), .A2(new_n2725_), .B(new_n1359_), .ZN(new_n3055_));
  NOR3_X1    g3006(.A1(new_n3053_), .A2(new_n3054_), .A3(new_n3055_), .ZN(new_n3056_));
  INV_X1     g3007(.I(new_n3056_), .ZN(new_n3057_));
  OAI22_X1   g3008(.A1(new_n2694_), .A2(new_n3051_), .B1(new_n2666_), .B2(new_n3057_), .ZN(new_n3058_));
  XNOR2_X1   g3009(.A1(new_n1452_), .A2(new_n52_), .ZN(new_n3059_));
  NOR2_X1    g3010(.A1(new_n3052_), .A2(new_n3059_), .ZN(new_n3060_));
  INV_X1     g3011(.I(new_n3060_), .ZN(new_n3061_));
  NOR2_X1    g3012(.A1(new_n2611_), .A2(new_n3061_), .ZN(new_n3062_));
  NOR2_X1    g3013(.A1(new_n3062_), .A2(new_n3058_), .ZN(new_n3063_));
  INV_X1     g3014(.I(new_n3063_), .ZN(new_n3064_));
  NOR2_X1    g3015(.A1(new_n2705_), .A2(new_n2706_), .ZN(new_n3065_));
  NAND3_X1   g3016(.A1(new_n2610_), .A2(new_n2608_), .A3(new_n2694_), .ZN(new_n3066_));
  OAI21_X1   g3017(.A1(new_n2714_), .A2(new_n2715_), .B(new_n2613_), .ZN(new_n3067_));
  NAND3_X1   g3018(.A1(new_n3067_), .A2(new_n3066_), .A3(new_n3065_), .ZN(new_n3068_));
  NAND2_X1   g3019(.A1(new_n2690_), .A2(new_n2667_), .ZN(new_n3069_));
  NOR3_X1    g3020(.A1(new_n2714_), .A2(new_n2715_), .A3(new_n2613_), .ZN(new_n3070_));
  AOI21_X1   g3021(.A1(new_n2610_), .A2(new_n2608_), .B(new_n2694_), .ZN(new_n3071_));
  OAI21_X1   g3022(.A1(new_n3070_), .A2(new_n3071_), .B(new_n3069_), .ZN(new_n3072_));
  NOR2_X1    g3023(.A1(new_n3053_), .A2(new_n3059_), .ZN(new_n3073_));
  INV_X1     g3024(.I(new_n3073_), .ZN(new_n3074_));
  AOI21_X1   g3025(.A1(new_n3072_), .A2(new_n3068_), .B(new_n3074_), .ZN(new_n3075_));
  OAI21_X1   g3026(.A1(new_n3075_), .A2(new_n3064_), .B(new_n1288_), .ZN(new_n3076_));
  NOR3_X1    g3027(.A1(new_n3070_), .A2(new_n3071_), .A3(new_n3069_), .ZN(new_n3077_));
  AOI21_X1   g3028(.A1(new_n3067_), .A2(new_n3066_), .B(new_n3065_), .ZN(new_n3078_));
  OAI21_X1   g3029(.A1(new_n3077_), .A2(new_n3078_), .B(new_n3073_), .ZN(new_n3079_));
  NAND3_X1   g3030(.A1(new_n3079_), .A2(new_n1287_), .A3(new_n3063_), .ZN(new_n3080_));
  NAND2_X1   g3031(.A1(new_n3076_), .A2(new_n3080_), .ZN(new_n3081_));
  NAND2_X1   g3032(.A1(new_n3048_), .A2(new_n3081_), .ZN(new_n3082_));
  NAND2_X1   g3033(.A1(new_n3027_), .A2(new_n3047_), .ZN(new_n3083_));
  NAND3_X1   g3034(.A1(new_n3083_), .A2(new_n3076_), .A3(new_n3080_), .ZN(new_n3084_));
  AOI21_X1   g3035(.A1(new_n2954_), .A2(new_n3030_), .B(new_n3042_), .ZN(new_n3085_));
  NOR3_X1    g3036(.A1(new_n2877_), .A2(new_n2953_), .A3(new_n3043_), .ZN(new_n3086_));
  NOR2_X1    g3037(.A1(new_n3086_), .A2(new_n3085_), .ZN(new_n3087_));
  NOR2_X1    g3038(.A1(new_n2956_), .A2(new_n3057_), .ZN(new_n3088_));
  NOR2_X1    g3039(.A1(new_n2694_), .A2(new_n3061_), .ZN(new_n3089_));
  NOR2_X1    g3040(.A1(new_n3089_), .A2(new_n3088_), .ZN(new_n3090_));
  OAI21_X1   g3041(.A1(new_n2666_), .A2(new_n3051_), .B(new_n3090_), .ZN(new_n3091_));
  NAND3_X1   g3042(.A1(new_n2693_), .A2(new_n2556_), .A3(new_n2670_), .ZN(new_n3092_));
  NAND2_X1   g3043(.A1(new_n2694_), .A2(new_n2689_), .ZN(new_n3093_));
  NAND3_X1   g3044(.A1(new_n3093_), .A2(new_n2666_), .A3(new_n3092_), .ZN(new_n3094_));
  OAI21_X1   g3045(.A1(new_n2612_), .A2(new_n2504_), .B(new_n2956_), .ZN(new_n3095_));
  OAI21_X1   g3046(.A1(new_n3095_), .A2(new_n2688_), .B(new_n3092_), .ZN(new_n3096_));
  OAI21_X1   g3047(.A1(new_n2956_), .A2(new_n2687_), .B(new_n2701_), .ZN(new_n3097_));
  NOR2_X1    g3048(.A1(new_n2694_), .A2(new_n3097_), .ZN(new_n3098_));
  AOI21_X1   g3049(.A1(new_n3096_), .A2(new_n2704_), .B(new_n3098_), .ZN(new_n3099_));
  AOI21_X1   g3050(.A1(new_n3099_), .A2(new_n3094_), .B(new_n3074_), .ZN(new_n3100_));
  OAI21_X1   g3051(.A1(new_n3100_), .A2(new_n3091_), .B(new_n1288_), .ZN(new_n3101_));
  INV_X1     g3052(.I(new_n3101_), .ZN(new_n3102_));
  NOR3_X1    g3053(.A1(new_n3100_), .A2(new_n1288_), .A3(new_n3091_), .ZN(new_n3103_));
  NOR3_X1    g3054(.A1(new_n3102_), .A2(new_n3103_), .A3(new_n3087_), .ZN(new_n3104_));
  OAI22_X1   g3055(.A1(new_n2956_), .A2(new_n3051_), .B1(new_n2858_), .B2(new_n3057_), .ZN(new_n3105_));
  NOR2_X1    g3056(.A1(new_n2666_), .A2(new_n3061_), .ZN(new_n3106_));
  NOR2_X1    g3057(.A1(new_n3106_), .A2(new_n3105_), .ZN(new_n3107_));
  INV_X1     g3058(.I(new_n3107_), .ZN(new_n3108_));
  AOI22_X1   g3059(.A1(new_n2669_), .A2(new_n2668_), .B1(new_n2858_), .B2(new_n2869_), .ZN(new_n3109_));
  NOR2_X1    g3060(.A1(new_n3109_), .A2(new_n2663_), .ZN(new_n3110_));
  NAND2_X1   g3061(.A1(new_n3110_), .A2(new_n2666_), .ZN(new_n3111_));
  NAND2_X1   g3062(.A1(new_n3097_), .A2(new_n2704_), .ZN(new_n3112_));
  AOI21_X1   g3063(.A1(new_n3112_), .A2(new_n3111_), .B(new_n3074_), .ZN(new_n3113_));
  OAI21_X1   g3064(.A1(new_n3108_), .A2(new_n3113_), .B(new_n1288_), .ZN(new_n3114_));
  INV_X1     g3065(.I(new_n3114_), .ZN(new_n3115_));
  NOR3_X1    g3066(.A1(new_n3108_), .A2(new_n3113_), .A3(new_n1288_), .ZN(new_n3116_));
  NOR3_X1    g3067(.A1(new_n3041_), .A2(new_n2952_), .A3(new_n2891_), .ZN(new_n3117_));
  AOI21_X1   g3068(.A1(new_n2892_), .A2(new_n2951_), .B(new_n2950_), .ZN(new_n3118_));
  NOR2_X1    g3069(.A1(new_n3117_), .A2(new_n3118_), .ZN(new_n3119_));
  OAI21_X1   g3070(.A1(new_n3115_), .A2(new_n3116_), .B(new_n3119_), .ZN(new_n3120_));
  INV_X1     g3071(.I(new_n3120_), .ZN(new_n3121_));
  INV_X1     g3072(.I(new_n3116_), .ZN(new_n3122_));
  NAND3_X1   g3073(.A1(new_n2892_), .A2(new_n2950_), .A3(new_n2951_), .ZN(new_n3123_));
  OAI21_X1   g3074(.A1(new_n2891_), .A2(new_n2952_), .B(new_n3041_), .ZN(new_n3124_));
  NAND2_X1   g3075(.A1(new_n3124_), .A2(new_n3123_), .ZN(new_n3125_));
  NAND3_X1   g3076(.A1(new_n3125_), .A2(new_n3122_), .A3(new_n3114_), .ZN(new_n3126_));
  NOR2_X1    g3077(.A1(new_n2956_), .A2(new_n3061_), .ZN(new_n3127_));
  NOR2_X1    g3078(.A1(new_n2697_), .A2(new_n3057_), .ZN(new_n3128_));
  NOR2_X1    g3079(.A1(new_n2858_), .A2(new_n3051_), .ZN(new_n3129_));
  NOR3_X1    g3080(.A1(new_n3127_), .A2(new_n3128_), .A3(new_n3129_), .ZN(new_n3130_));
  NAND2_X1   g3081(.A1(new_n2976_), .A2(new_n3073_), .ZN(new_n3131_));
  AOI21_X1   g3082(.A1(new_n3131_), .A2(new_n3130_), .B(new_n1287_), .ZN(new_n3132_));
  NAND3_X1   g3083(.A1(new_n3131_), .A2(new_n1287_), .A3(new_n3130_), .ZN(new_n3133_));
  INV_X1     g3084(.I(new_n3133_), .ZN(new_n3134_));
  OAI21_X1   g3085(.A1(new_n2912_), .A2(new_n3040_), .B(new_n2948_), .ZN(new_n3135_));
  NAND3_X1   g3086(.A1(new_n3039_), .A2(new_n3033_), .A3(new_n2949_), .ZN(new_n3136_));
  NAND2_X1   g3087(.A1(new_n3136_), .A2(new_n3135_), .ZN(new_n3137_));
  INV_X1     g3088(.I(new_n3137_), .ZN(new_n3138_));
  OAI21_X1   g3089(.A1(new_n3134_), .A2(new_n3132_), .B(new_n3138_), .ZN(new_n3139_));
  NOR3_X1    g3090(.A1(new_n3134_), .A2(new_n3138_), .A3(new_n3132_), .ZN(new_n3140_));
  INV_X1     g3091(.I(new_n3051_), .ZN(new_n3141_));
  NAND2_X1   g3092(.A1(new_n2630_), .A2(new_n3141_), .ZN(new_n3142_));
  NAND2_X1   g3093(.A1(new_n2800_), .A2(new_n3056_), .ZN(new_n3143_));
  NAND2_X1   g3094(.A1(new_n3142_), .A2(new_n3143_), .ZN(new_n3144_));
  AOI21_X1   g3095(.A1(new_n2881_), .A2(new_n3060_), .B(new_n3144_), .ZN(new_n3145_));
  AOI21_X1   g3096(.A1(new_n2698_), .A2(new_n2868_), .B(new_n2697_), .ZN(new_n3146_));
  NOR2_X1    g3097(.A1(new_n2882_), .A2(new_n2881_), .ZN(new_n3147_));
  OAI21_X1   g3098(.A1(new_n3147_), .A2(new_n3146_), .B(new_n3073_), .ZN(new_n3148_));
  AOI21_X1   g3099(.A1(new_n3148_), .A2(new_n3145_), .B(new_n1287_), .ZN(new_n3149_));
  NAND2_X1   g3100(.A1(new_n2881_), .A2(new_n3060_), .ZN(new_n3150_));
  NAND3_X1   g3101(.A1(new_n3150_), .A2(new_n3142_), .A3(new_n3143_), .ZN(new_n3151_));
  AOI21_X1   g3102(.A1(new_n2883_), .A2(new_n2884_), .B(new_n3074_), .ZN(new_n3152_));
  NOR3_X1    g3103(.A1(new_n3152_), .A2(new_n1288_), .A3(new_n3151_), .ZN(new_n3153_));
  AOI21_X1   g3104(.A1(new_n2934_), .A2(new_n2927_), .B(new_n846_), .ZN(new_n3154_));
  NOR3_X1    g3105(.A1(new_n2928_), .A2(new_n2932_), .A3(new_n845_), .ZN(new_n3155_));
  NOR3_X1    g3106(.A1(new_n3155_), .A2(new_n3154_), .A3(new_n2747_), .ZN(new_n3156_));
  NOR3_X1    g3107(.A1(new_n2936_), .A2(new_n3156_), .A3(new_n2945_), .ZN(new_n3157_));
  OAI21_X1   g3108(.A1(new_n3155_), .A2(new_n3154_), .B(new_n2747_), .ZN(new_n3158_));
  AOI21_X1   g3109(.A1(new_n3158_), .A2(new_n2946_), .B(new_n2944_), .ZN(new_n3159_));
  NOR2_X1    g3110(.A1(new_n3157_), .A2(new_n3159_), .ZN(new_n3160_));
  NOR3_X1    g3111(.A1(new_n3149_), .A2(new_n3153_), .A3(new_n3160_), .ZN(new_n3161_));
  INV_X1     g3112(.I(new_n3161_), .ZN(new_n3162_));
  XOR2_X1    g3113(.A1(new_n2942_), .A2(new_n845_), .Z(new_n3163_));
  NOR2_X1    g3114(.A1(new_n2943_), .A2(new_n846_), .ZN(new_n3164_));
  INV_X1     g3115(.I(new_n3164_), .ZN(new_n3165_));
  NAND2_X1   g3116(.A1(new_n2942_), .A2(new_n845_), .ZN(new_n3166_));
  NOR2_X1    g3117(.A1(new_n3166_), .A2(new_n2943_), .ZN(new_n3167_));
  AOI21_X1   g3118(.A1(new_n3163_), .A2(new_n3165_), .B(new_n3167_), .ZN(new_n3168_));
  INV_X1     g3119(.I(new_n3168_), .ZN(new_n3169_));
  OAI22_X1   g3120(.A1(new_n2654_), .A2(new_n3061_), .B1(new_n2657_), .B2(new_n3051_), .ZN(new_n3170_));
  INV_X1     g3121(.I(new_n3170_), .ZN(new_n3171_));
  OAI21_X1   g3122(.A1(new_n2742_), .A2(new_n3074_), .B(new_n3171_), .ZN(new_n3172_));
  NOR2_X1    g3123(.A1(new_n2657_), .A2(new_n3059_), .ZN(new_n3173_));
  AOI22_X1   g3124(.A1(new_n2682_), .A2(new_n3141_), .B1(new_n2741_), .B2(new_n3056_), .ZN(new_n3174_));
  NAND2_X1   g3125(.A1(new_n2754_), .A2(new_n3060_), .ZN(new_n3175_));
  NAND3_X1   g3126(.A1(new_n2781_), .A2(new_n2780_), .A3(new_n3073_), .ZN(new_n3176_));
  NAND3_X1   g3127(.A1(new_n3176_), .A2(new_n3174_), .A3(new_n3175_), .ZN(new_n3177_));
  NOR4_X1    g3128(.A1(new_n3177_), .A2(new_n1288_), .A3(new_n3172_), .A4(new_n3173_), .ZN(new_n3178_));
  NAND2_X1   g3129(.A1(new_n3178_), .A2(new_n2943_), .ZN(new_n3179_));
  OAI22_X1   g3130(.A1(new_n2757_), .A2(new_n3051_), .B1(new_n2654_), .B2(new_n3057_), .ZN(new_n3180_));
  AOI21_X1   g3131(.A1(new_n2645_), .A2(new_n3060_), .B(new_n3180_), .ZN(new_n3181_));
  NAND3_X1   g3132(.A1(new_n2773_), .A2(new_n2771_), .A3(new_n3073_), .ZN(new_n3182_));
  AOI21_X1   g3133(.A1(new_n3182_), .A2(new_n3181_), .B(new_n1287_), .ZN(new_n3183_));
  AOI22_X1   g3134(.A1(new_n2754_), .A2(new_n3141_), .B1(new_n2682_), .B2(new_n3056_), .ZN(new_n3184_));
  OAI21_X1   g3135(.A1(new_n2679_), .A2(new_n3061_), .B(new_n3184_), .ZN(new_n3185_));
  NOR3_X1    g3136(.A1(new_n2931_), .A2(new_n2929_), .A3(new_n3074_), .ZN(new_n3186_));
  NOR3_X1    g3137(.A1(new_n3186_), .A2(new_n1288_), .A3(new_n3185_), .ZN(new_n3187_));
  NOR2_X1    g3138(.A1(new_n3187_), .A2(new_n3183_), .ZN(new_n3188_));
  NOR2_X1    g3139(.A1(new_n3178_), .A2(new_n2943_), .ZN(new_n3189_));
  OAI21_X1   g3140(.A1(new_n3188_), .A2(new_n3189_), .B(new_n3179_), .ZN(new_n3190_));
  NOR2_X1    g3141(.A1(new_n3190_), .A2(new_n3169_), .ZN(new_n3191_));
  OAI22_X1   g3142(.A1(new_n2679_), .A2(new_n3051_), .B1(new_n2757_), .B2(new_n3057_), .ZN(new_n3192_));
  NOR2_X1    g3143(.A1(new_n2792_), .A2(new_n3061_), .ZN(new_n3193_));
  NOR2_X1    g3144(.A1(new_n3193_), .A2(new_n3192_), .ZN(new_n3194_));
  AOI21_X1   g3145(.A1(new_n2799_), .A2(new_n2804_), .B(new_n3074_), .ZN(new_n3195_));
  INV_X1     g3146(.I(new_n3195_), .ZN(new_n3196_));
  AOI21_X1   g3147(.A1(new_n3196_), .A2(new_n3194_), .B(new_n1287_), .ZN(new_n3197_));
  INV_X1     g3148(.I(new_n3194_), .ZN(new_n3198_));
  NOR3_X1    g3149(.A1(new_n3198_), .A2(new_n3195_), .A3(new_n1288_), .ZN(new_n3199_));
  NOR2_X1    g3150(.A1(new_n3197_), .A2(new_n3199_), .ZN(new_n3200_));
  NAND2_X1   g3151(.A1(new_n3190_), .A2(new_n3169_), .ZN(new_n3201_));
  AOI21_X1   g3152(.A1(new_n3200_), .A2(new_n3201_), .B(new_n3191_), .ZN(new_n3202_));
  OAI22_X1   g3153(.A1(new_n2792_), .A2(new_n3051_), .B1(new_n2679_), .B2(new_n3057_), .ZN(new_n3203_));
  NOR2_X1    g3154(.A1(new_n2845_), .A2(new_n3061_), .ZN(new_n3204_));
  NOR2_X1    g3155(.A1(new_n3204_), .A2(new_n3203_), .ZN(new_n3205_));
  OAI21_X1   g3156(.A1(new_n2989_), .A2(new_n2988_), .B(new_n3073_), .ZN(new_n3206_));
  AOI21_X1   g3157(.A1(new_n3206_), .A2(new_n3205_), .B(new_n1287_), .ZN(new_n3207_));
  INV_X1     g3158(.I(new_n3207_), .ZN(new_n3208_));
  NAND3_X1   g3159(.A1(new_n3206_), .A2(new_n1287_), .A3(new_n3205_), .ZN(new_n3209_));
  NAND2_X1   g3160(.A1(new_n3208_), .A2(new_n3209_), .ZN(new_n3210_));
  NOR2_X1    g3161(.A1(new_n3202_), .A2(new_n3210_), .ZN(new_n3211_));
  XOR2_X1    g3162(.A1(new_n2940_), .A2(new_n845_), .Z(new_n3212_));
  AOI21_X1   g3163(.A1(new_n3163_), .A2(new_n3164_), .B(new_n3212_), .ZN(new_n3213_));
  NOR2_X1    g3164(.A1(new_n3213_), .A2(new_n2944_), .ZN(new_n3214_));
  AOI21_X1   g3165(.A1(new_n3202_), .A2(new_n3210_), .B(new_n3214_), .ZN(new_n3215_));
  OAI21_X1   g3166(.A1(new_n3149_), .A2(new_n3153_), .B(new_n3160_), .ZN(new_n3216_));
  OAI21_X1   g3167(.A1(new_n3215_), .A2(new_n3211_), .B(new_n3216_), .ZN(new_n3217_));
  AOI22_X1   g3168(.A1(new_n2881_), .A2(new_n3141_), .B1(new_n2630_), .B2(new_n3056_), .ZN(new_n3218_));
  NAND2_X1   g3169(.A1(new_n2671_), .A2(new_n3060_), .ZN(new_n3219_));
  NAND2_X1   g3170(.A1(new_n3219_), .A2(new_n3218_), .ZN(new_n3220_));
  AOI21_X1   g3171(.A1(new_n2871_), .A2(new_n2865_), .B(new_n3074_), .ZN(new_n3221_));
  OAI21_X1   g3172(.A1(new_n3221_), .A2(new_n3220_), .B(new_n1288_), .ZN(new_n3222_));
  INV_X1     g3173(.I(new_n3220_), .ZN(new_n3223_));
  NOR2_X1    g3174(.A1(new_n2870_), .A2(new_n2671_), .ZN(new_n3224_));
  NOR2_X1    g3175(.A1(new_n2864_), .A2(new_n2858_), .ZN(new_n3225_));
  OAI21_X1   g3176(.A1(new_n3224_), .A2(new_n3225_), .B(new_n3073_), .ZN(new_n3226_));
  NAND3_X1   g3177(.A1(new_n3223_), .A2(new_n3226_), .A3(new_n1287_), .ZN(new_n3227_));
  NAND2_X1   g3178(.A1(new_n3227_), .A2(new_n3222_), .ZN(new_n3228_));
  AOI21_X1   g3179(.A1(new_n3217_), .A2(new_n3162_), .B(new_n3228_), .ZN(new_n3229_));
  NAND3_X1   g3180(.A1(new_n3217_), .A2(new_n3162_), .A3(new_n3228_), .ZN(new_n3230_));
  NOR3_X1    g3181(.A1(new_n3036_), .A2(new_n2925_), .A3(new_n3038_), .ZN(new_n3231_));
  AOI21_X1   g3182(.A1(new_n3037_), .A2(new_n2924_), .B(new_n2947_), .ZN(new_n3232_));
  NOR2_X1    g3183(.A1(new_n3232_), .A2(new_n3231_), .ZN(new_n3233_));
  INV_X1     g3184(.I(new_n3233_), .ZN(new_n3234_));
  AOI21_X1   g3185(.A1(new_n3230_), .A2(new_n3234_), .B(new_n3229_), .ZN(new_n3235_));
  INV_X1     g3186(.I(new_n3235_), .ZN(new_n3236_));
  OAI21_X1   g3187(.A1(new_n3236_), .A2(new_n3140_), .B(new_n3139_), .ZN(new_n3237_));
  AOI21_X1   g3188(.A1(new_n3237_), .A2(new_n3126_), .B(new_n3121_), .ZN(new_n3238_));
  OAI21_X1   g3189(.A1(new_n3102_), .A2(new_n3103_), .B(new_n3087_), .ZN(new_n3239_));
  AOI21_X1   g3190(.A1(new_n3238_), .A2(new_n3239_), .B(new_n3104_), .ZN(new_n3240_));
  NAND3_X1   g3191(.A1(new_n3240_), .A2(new_n3082_), .A3(new_n3084_), .ZN(new_n3241_));
  AOI21_X1   g3192(.A1(new_n3076_), .A2(new_n3080_), .B(new_n3083_), .ZN(new_n3242_));
  NOR2_X1    g3193(.A1(new_n3048_), .A2(new_n3081_), .ZN(new_n3243_));
  OR2_X2     g3194(.A1(new_n3086_), .A2(new_n3085_), .Z(new_n3244_));
  INV_X1     g3195(.I(new_n3103_), .ZN(new_n3245_));
  NAND3_X1   g3196(.A1(new_n3245_), .A2(new_n3244_), .A3(new_n3101_), .ZN(new_n3246_));
  NAND2_X1   g3197(.A1(new_n3120_), .A2(new_n3126_), .ZN(new_n3247_));
  INV_X1     g3198(.I(new_n3132_), .ZN(new_n3248_));
  AOI21_X1   g3199(.A1(new_n3248_), .A2(new_n3133_), .B(new_n3137_), .ZN(new_n3249_));
  NAND3_X1   g3200(.A1(new_n3248_), .A2(new_n3133_), .A3(new_n3137_), .ZN(new_n3250_));
  AOI21_X1   g3201(.A1(new_n3250_), .A2(new_n3235_), .B(new_n3249_), .ZN(new_n3251_));
  OAI21_X1   g3202(.A1(new_n3251_), .A2(new_n3247_), .B(new_n3120_), .ZN(new_n3252_));
  AOI21_X1   g3203(.A1(new_n3245_), .A2(new_n3101_), .B(new_n3244_), .ZN(new_n3253_));
  OAI21_X1   g3204(.A1(new_n3252_), .A2(new_n3253_), .B(new_n3246_), .ZN(new_n3254_));
  OAI21_X1   g3205(.A1(new_n3242_), .A2(new_n3243_), .B(new_n3254_), .ZN(new_n3255_));
  NAND3_X1   g3206(.A1(new_n2732_), .A2(new_n3255_), .A3(new_n3241_), .ZN(new_n3256_));
  INV_X1     g3207(.I(new_n3256_), .ZN(new_n3257_));
  OAI22_X1   g3208(.A1(new_n2563_), .A2(new_n2588_), .B1(new_n56_), .B2(new_n2611_), .ZN(new_n3258_));
  NOR2_X1    g3209(.A1(new_n2586_), .A2(new_n2601_), .ZN(new_n3259_));
  NOR2_X1    g3210(.A1(new_n3259_), .A2(new_n3258_), .ZN(new_n3260_));
  INV_X1     g3211(.I(new_n3260_), .ZN(new_n3261_));
  AOI21_X1   g3212(.A1(new_n2691_), .A2(new_n2611_), .B(new_n2705_), .ZN(new_n3262_));
  OAI21_X1   g3213(.A1(new_n3262_), .A2(new_n2563_), .B(new_n2708_), .ZN(new_n3263_));
  OAI21_X1   g3214(.A1(new_n2508_), .A2(new_n2562_), .B(new_n2716_), .ZN(new_n3264_));
  NAND2_X1   g3215(.A1(new_n2586_), .A2(new_n3264_), .ZN(new_n3265_));
  AOI21_X1   g3216(.A1(new_n2605_), .A2(new_n2606_), .B(new_n2611_), .ZN(new_n3266_));
  NAND2_X1   g3217(.A1(new_n3266_), .A2(new_n2604_), .ZN(new_n3267_));
  NAND2_X1   g3218(.A1(new_n3265_), .A2(new_n3267_), .ZN(new_n3268_));
  NAND2_X1   g3219(.A1(new_n3268_), .A2(new_n3263_), .ZN(new_n3269_));
  INV_X1     g3220(.I(new_n3263_), .ZN(new_n3270_));
  NAND3_X1   g3221(.A1(new_n3270_), .A2(new_n3265_), .A3(new_n3267_), .ZN(new_n3271_));
  AOI21_X1   g3222(.A1(new_n3269_), .A2(new_n3271_), .B(new_n2729_), .ZN(new_n3272_));
  OAI21_X1   g3223(.A1(new_n3272_), .A2(new_n3261_), .B(new_n52_), .ZN(new_n3273_));
  AOI21_X1   g3224(.A1(new_n3265_), .A2(new_n3267_), .B(new_n3270_), .ZN(new_n3274_));
  NOR2_X1    g3225(.A1(new_n3268_), .A2(new_n3263_), .ZN(new_n3275_));
  OAI21_X1   g3226(.A1(new_n3275_), .A2(new_n3274_), .B(new_n2722_), .ZN(new_n3276_));
  NAND3_X1   g3227(.A1(new_n3276_), .A2(new_n2725_), .A3(new_n3260_), .ZN(new_n3277_));
  NAND2_X1   g3228(.A1(new_n3277_), .A2(new_n3273_), .ZN(new_n3278_));
  NOR3_X1    g3229(.A1(new_n3252_), .A2(new_n3253_), .A3(new_n3104_), .ZN(new_n3279_));
  AOI21_X1   g3230(.A1(new_n3246_), .A2(new_n3239_), .B(new_n3238_), .ZN(new_n3280_));
  NOR2_X1    g3231(.A1(new_n3280_), .A2(new_n3279_), .ZN(new_n3281_));
  NAND2_X1   g3232(.A1(new_n3278_), .A2(new_n3281_), .ZN(new_n3282_));
  INV_X1     g3233(.I(new_n3282_), .ZN(new_n3283_));
  NOR2_X1    g3234(.A1(new_n2956_), .A2(new_n56_), .ZN(new_n3284_));
  NOR2_X1    g3235(.A1(new_n2694_), .A2(new_n2601_), .ZN(new_n3285_));
  NOR2_X1    g3236(.A1(new_n2666_), .A2(new_n2588_), .ZN(new_n3286_));
  NOR3_X1    g3237(.A1(new_n3285_), .A2(new_n3284_), .A3(new_n3286_), .ZN(new_n3287_));
  NOR3_X1    g3238(.A1(new_n2612_), .A2(new_n2504_), .A3(new_n2956_), .ZN(new_n3288_));
  AOI21_X1   g3239(.A1(new_n2670_), .A2(new_n2688_), .B(new_n2613_), .ZN(new_n3289_));
  NOR3_X1    g3240(.A1(new_n3289_), .A2(new_n2704_), .A3(new_n3288_), .ZN(new_n3290_));
  INV_X1     g3241(.I(new_n2688_), .ZN(new_n3291_));
  AOI21_X1   g3242(.A1(new_n2693_), .A2(new_n2556_), .B(new_n2670_), .ZN(new_n3292_));
  AOI21_X1   g3243(.A1(new_n3291_), .A2(new_n3292_), .B(new_n3288_), .ZN(new_n3293_));
  NAND2_X1   g3244(.A1(new_n2613_), .A2(new_n3110_), .ZN(new_n3294_));
  OAI21_X1   g3245(.A1(new_n3293_), .A2(new_n2666_), .B(new_n3294_), .ZN(new_n3295_));
  OAI21_X1   g3246(.A1(new_n3295_), .A2(new_n3290_), .B(new_n2722_), .ZN(new_n3296_));
  AOI21_X1   g3247(.A1(new_n3296_), .A2(new_n3287_), .B(new_n52_), .ZN(new_n3297_));
  INV_X1     g3248(.I(new_n3287_), .ZN(new_n3298_));
  AOI21_X1   g3249(.A1(new_n3099_), .A2(new_n3094_), .B(new_n2729_), .ZN(new_n3299_));
  NOR3_X1    g3250(.A1(new_n3299_), .A2(new_n2725_), .A3(new_n3298_), .ZN(new_n3300_));
  INV_X1     g3251(.I(new_n2943_), .ZN(new_n3301_));
  XOR2_X1    g3252(.A1(new_n2654_), .A2(new_n2657_), .Z(new_n3302_));
  AOI21_X1   g3253(.A1(new_n3302_), .A2(new_n3073_), .B(new_n3170_), .ZN(new_n3303_));
  INV_X1     g3254(.I(new_n3173_), .ZN(new_n3304_));
  OAI21_X1   g3255(.A1(new_n2757_), .A2(new_n3061_), .B(new_n3174_), .ZN(new_n3305_));
  AOI21_X1   g3256(.A1(new_n2762_), .A2(new_n3073_), .B(new_n3305_), .ZN(new_n3306_));
  NAND4_X1   g3257(.A1(new_n3306_), .A2(new_n1287_), .A3(new_n3303_), .A4(new_n3304_), .ZN(new_n3307_));
  NOR2_X1    g3258(.A1(new_n3307_), .A2(new_n3301_), .ZN(new_n3308_));
  OAI21_X1   g3259(.A1(new_n3186_), .A2(new_n3185_), .B(new_n1288_), .ZN(new_n3309_));
  NAND3_X1   g3260(.A1(new_n3182_), .A2(new_n1287_), .A3(new_n3181_), .ZN(new_n3310_));
  NAND2_X1   g3261(.A1(new_n3309_), .A2(new_n3310_), .ZN(new_n3311_));
  NAND2_X1   g3262(.A1(new_n3307_), .A2(new_n3301_), .ZN(new_n3312_));
  AOI21_X1   g3263(.A1(new_n3311_), .A2(new_n3312_), .B(new_n3308_), .ZN(new_n3313_));
  NAND2_X1   g3264(.A1(new_n3313_), .A2(new_n3168_), .ZN(new_n3314_));
  OAI21_X1   g3265(.A1(new_n3198_), .A2(new_n3195_), .B(new_n1288_), .ZN(new_n3315_));
  NAND3_X1   g3266(.A1(new_n3196_), .A2(new_n1287_), .A3(new_n3194_), .ZN(new_n3316_));
  NAND2_X1   g3267(.A1(new_n3316_), .A2(new_n3315_), .ZN(new_n3317_));
  NOR2_X1    g3268(.A1(new_n3313_), .A2(new_n3168_), .ZN(new_n3318_));
  OAI21_X1   g3269(.A1(new_n3317_), .A2(new_n3318_), .B(new_n3314_), .ZN(new_n3319_));
  AND3_X2    g3270(.A1(new_n3206_), .A2(new_n1287_), .A3(new_n3205_), .Z(new_n3320_));
  NOR2_X1    g3271(.A1(new_n3320_), .A2(new_n3207_), .ZN(new_n3321_));
  NAND2_X1   g3272(.A1(new_n3319_), .A2(new_n3321_), .ZN(new_n3322_));
  INV_X1     g3273(.I(new_n3214_), .ZN(new_n3323_));
  OAI21_X1   g3274(.A1(new_n3319_), .A2(new_n3321_), .B(new_n3323_), .ZN(new_n3324_));
  OAI21_X1   g3275(.A1(new_n3152_), .A2(new_n3151_), .B(new_n1288_), .ZN(new_n3325_));
  NAND3_X1   g3276(.A1(new_n3148_), .A2(new_n1287_), .A3(new_n3145_), .ZN(new_n3326_));
  NAND3_X1   g3277(.A1(new_n3158_), .A2(new_n2946_), .A3(new_n2944_), .ZN(new_n3327_));
  OAI21_X1   g3278(.A1(new_n2936_), .A2(new_n3156_), .B(new_n2945_), .ZN(new_n3328_));
  NAND2_X1   g3279(.A1(new_n3328_), .A2(new_n3327_), .ZN(new_n3329_));
  AOI21_X1   g3280(.A1(new_n3326_), .A2(new_n3325_), .B(new_n3329_), .ZN(new_n3330_));
  AOI21_X1   g3281(.A1(new_n3324_), .A2(new_n3322_), .B(new_n3330_), .ZN(new_n3331_));
  AOI21_X1   g3282(.A1(new_n3223_), .A2(new_n3226_), .B(new_n1287_), .ZN(new_n3332_));
  NOR3_X1    g3283(.A1(new_n3221_), .A2(new_n1288_), .A3(new_n3220_), .ZN(new_n3333_));
  NOR2_X1    g3284(.A1(new_n3332_), .A2(new_n3333_), .ZN(new_n3334_));
  NOR3_X1    g3285(.A1(new_n3331_), .A2(new_n3334_), .A3(new_n3161_), .ZN(new_n3335_));
  OAI21_X1   g3286(.A1(new_n3229_), .A2(new_n3335_), .B(new_n3233_), .ZN(new_n3336_));
  OAI21_X1   g3287(.A1(new_n3331_), .A2(new_n3161_), .B(new_n3334_), .ZN(new_n3337_));
  NAND3_X1   g3288(.A1(new_n3230_), .A2(new_n3337_), .A3(new_n3234_), .ZN(new_n3338_));
  NAND2_X1   g3289(.A1(new_n3336_), .A2(new_n3338_), .ZN(new_n3339_));
  NOR3_X1    g3290(.A1(new_n3297_), .A2(new_n3300_), .A3(new_n3339_), .ZN(new_n3340_));
  INV_X1     g3291(.I(new_n3340_), .ZN(new_n3341_));
  NOR2_X1    g3292(.A1(new_n2697_), .A2(new_n56_), .ZN(new_n3342_));
  NOR2_X1    g3293(.A1(new_n2858_), .A2(new_n2588_), .ZN(new_n3343_));
  NOR2_X1    g3294(.A1(new_n2956_), .A2(new_n2601_), .ZN(new_n3344_));
  NOR3_X1    g3295(.A1(new_n3344_), .A2(new_n3342_), .A3(new_n3343_), .ZN(new_n3345_));
  NAND2_X1   g3296(.A1(new_n2976_), .A2(new_n2722_), .ZN(new_n3346_));
  AOI21_X1   g3297(.A1(new_n3346_), .A2(new_n3345_), .B(new_n52_), .ZN(new_n3347_));
  INV_X1     g3298(.I(new_n3345_), .ZN(new_n3348_));
  AOI21_X1   g3299(.A1(new_n2968_), .A2(new_n2964_), .B(new_n2729_), .ZN(new_n3349_));
  NOR3_X1    g3300(.A1(new_n3349_), .A2(new_n2725_), .A3(new_n3348_), .ZN(new_n3350_));
  NOR2_X1    g3301(.A1(new_n3319_), .A2(new_n3321_), .ZN(new_n3351_));
  OAI21_X1   g3302(.A1(new_n3211_), .A2(new_n3351_), .B(new_n3214_), .ZN(new_n3352_));
  NAND2_X1   g3303(.A1(new_n3202_), .A2(new_n3210_), .ZN(new_n3353_));
  NAND3_X1   g3304(.A1(new_n3353_), .A2(new_n3322_), .A3(new_n3323_), .ZN(new_n3354_));
  NAND2_X1   g3305(.A1(new_n3352_), .A2(new_n3354_), .ZN(new_n3355_));
  NOR3_X1    g3306(.A1(new_n3350_), .A2(new_n3347_), .A3(new_n3355_), .ZN(new_n3356_));
  AOI22_X1   g3307(.A1(new_n2682_), .A2(new_n2587_), .B1(new_n55_), .B2(new_n2741_), .ZN(new_n3357_));
  INV_X1     g3308(.I(new_n2601_), .ZN(new_n3358_));
  NAND2_X1   g3309(.A1(new_n2754_), .A2(new_n3358_), .ZN(new_n3359_));
  AOI21_X1   g3310(.A1(new_n3359_), .A2(new_n3357_), .B(new_n2725_), .ZN(new_n3360_));
  OAI21_X1   g3311(.A1(new_n2657_), .A2(new_n50_), .B(new_n52_), .ZN(new_n3361_));
  NOR2_X1    g3312(.A1(new_n2654_), .A2(new_n2601_), .ZN(new_n3362_));
  NOR2_X1    g3313(.A1(new_n3362_), .A2(new_n3361_), .ZN(new_n3363_));
  NOR2_X1    g3314(.A1(new_n2725_), .A2(new_n2729_), .ZN(new_n3364_));
  INV_X1     g3315(.I(new_n3364_), .ZN(new_n3365_));
  AOI21_X1   g3316(.A1(new_n2781_), .A2(new_n2780_), .B(new_n3302_), .ZN(new_n3366_));
  OAI21_X1   g3317(.A1(new_n3366_), .A2(new_n3365_), .B(new_n3363_), .ZN(new_n3367_));
  NOR3_X1    g3318(.A1(new_n3367_), .A2(new_n3304_), .A3(new_n3360_), .ZN(new_n3368_));
  INV_X1     g3319(.I(new_n3360_), .ZN(new_n3369_));
  INV_X1     g3320(.I(new_n3363_), .ZN(new_n3370_));
  OAI21_X1   g3321(.A1(new_n2759_), .A2(new_n2761_), .B(new_n2742_), .ZN(new_n3371_));
  AOI21_X1   g3322(.A1(new_n3371_), .A2(new_n3364_), .B(new_n3370_), .ZN(new_n3372_));
  AOI21_X1   g3323(.A1(new_n3372_), .A2(new_n3369_), .B(new_n3173_), .ZN(new_n3373_));
  NOR3_X1    g3324(.A1(new_n2931_), .A2(new_n2929_), .A3(new_n2729_), .ZN(new_n3374_));
  AOI22_X1   g3325(.A1(new_n2754_), .A2(new_n2587_), .B1(new_n55_), .B2(new_n2682_), .ZN(new_n3375_));
  OAI21_X1   g3326(.A1(new_n2601_), .A2(new_n2679_), .B(new_n3375_), .ZN(new_n3376_));
  OAI21_X1   g3327(.A1(new_n3374_), .A2(new_n3376_), .B(new_n2725_), .ZN(new_n3377_));
  NAND3_X1   g3328(.A1(new_n2773_), .A2(new_n2771_), .A3(new_n2722_), .ZN(new_n3378_));
  OAI22_X1   g3329(.A1(new_n2757_), .A2(new_n2588_), .B1(new_n56_), .B2(new_n2654_), .ZN(new_n3379_));
  AOI21_X1   g3330(.A1(new_n3358_), .A2(new_n2645_), .B(new_n3379_), .ZN(new_n3380_));
  NAND3_X1   g3331(.A1(new_n3378_), .A2(new_n52_), .A3(new_n3380_), .ZN(new_n3381_));
  AOI21_X1   g3332(.A1(new_n3377_), .A2(new_n3381_), .B(new_n3373_), .ZN(new_n3382_));
  NOR3_X1    g3333(.A1(new_n3172_), .A2(new_n1288_), .A3(new_n3173_), .ZN(new_n3383_));
  NOR2_X1    g3334(.A1(new_n3303_), .A2(new_n1287_), .ZN(new_n3384_));
  NOR2_X1    g3335(.A1(new_n3172_), .A2(new_n1288_), .ZN(new_n3385_));
  NOR2_X1    g3336(.A1(new_n3173_), .A2(new_n1288_), .ZN(new_n3386_));
  NOR3_X1    g3337(.A1(new_n3384_), .A2(new_n3385_), .A3(new_n3386_), .ZN(new_n3387_));
  NOR2_X1    g3338(.A1(new_n3387_), .A2(new_n3383_), .ZN(new_n3388_));
  NOR3_X1    g3339(.A1(new_n3382_), .A2(new_n3368_), .A3(new_n3388_), .ZN(new_n3389_));
  AOI22_X1   g3340(.A1(new_n2645_), .A2(new_n2587_), .B1(new_n55_), .B2(new_n2754_), .ZN(new_n3390_));
  NAND2_X1   g3341(.A1(new_n2800_), .A2(new_n3358_), .ZN(new_n3391_));
  NAND2_X1   g3342(.A1(new_n3391_), .A2(new_n3390_), .ZN(new_n3392_));
  INV_X1     g3343(.I(new_n3392_), .ZN(new_n3393_));
  OAI21_X1   g3344(.A1(new_n2807_), .A2(new_n2808_), .B(new_n2722_), .ZN(new_n3394_));
  AOI21_X1   g3345(.A1(new_n3393_), .A2(new_n3394_), .B(new_n52_), .ZN(new_n3395_));
  AOI21_X1   g3346(.A1(new_n2799_), .A2(new_n2804_), .B(new_n2729_), .ZN(new_n3396_));
  NOR3_X1    g3347(.A1(new_n3396_), .A2(new_n2725_), .A3(new_n3392_), .ZN(new_n3397_));
  NOR2_X1    g3348(.A1(new_n3395_), .A2(new_n3397_), .ZN(new_n3398_));
  OAI21_X1   g3349(.A1(new_n3382_), .A2(new_n3368_), .B(new_n3388_), .ZN(new_n3399_));
  AOI21_X1   g3350(.A1(new_n3398_), .A2(new_n3399_), .B(new_n3389_), .ZN(new_n3400_));
  OAI22_X1   g3351(.A1(new_n2792_), .A2(new_n2588_), .B1(new_n56_), .B2(new_n2679_), .ZN(new_n3401_));
  AOI21_X1   g3352(.A1(new_n3358_), .A2(new_n2630_), .B(new_n3401_), .ZN(new_n3402_));
  OAI21_X1   g3353(.A1(new_n2989_), .A2(new_n2988_), .B(new_n2722_), .ZN(new_n3403_));
  AOI21_X1   g3354(.A1(new_n3403_), .A2(new_n3402_), .B(new_n2725_), .ZN(new_n3404_));
  AOI22_X1   g3355(.A1(new_n2800_), .A2(new_n2587_), .B1(new_n55_), .B2(new_n2645_), .ZN(new_n3405_));
  OAI21_X1   g3356(.A1(new_n2845_), .A2(new_n2601_), .B(new_n3405_), .ZN(new_n3406_));
  AOI21_X1   g3357(.A1(new_n2902_), .A2(new_n2901_), .B(new_n2729_), .ZN(new_n3407_));
  NOR3_X1    g3358(.A1(new_n3407_), .A2(new_n52_), .A3(new_n3406_), .ZN(new_n3408_));
  NOR2_X1    g3359(.A1(new_n3408_), .A2(new_n3404_), .ZN(new_n3409_));
  NOR2_X1    g3360(.A1(new_n3400_), .A2(new_n3409_), .ZN(new_n3410_));
  INV_X1     g3361(.I(new_n3383_), .ZN(new_n3411_));
  XOR2_X1    g3362(.A1(new_n3306_), .A2(new_n1287_), .Z(new_n3412_));
  NAND2_X1   g3363(.A1(new_n3412_), .A2(new_n3411_), .ZN(new_n3413_));
  NAND2_X1   g3364(.A1(new_n3413_), .A2(new_n3307_), .ZN(new_n3414_));
  INV_X1     g3365(.I(new_n3414_), .ZN(new_n3415_));
  AOI21_X1   g3366(.A1(new_n3400_), .A2(new_n3409_), .B(new_n3415_), .ZN(new_n3416_));
  NOR2_X1    g3367(.A1(new_n3416_), .A2(new_n3410_), .ZN(new_n3417_));
  OAI22_X1   g3368(.A1(new_n2845_), .A2(new_n2588_), .B1(new_n56_), .B2(new_n2792_), .ZN(new_n3418_));
  NOR2_X1    g3369(.A1(new_n2697_), .A2(new_n2601_), .ZN(new_n3419_));
  NOR2_X1    g3370(.A1(new_n3419_), .A2(new_n3418_), .ZN(new_n3420_));
  INV_X1     g3371(.I(new_n3420_), .ZN(new_n3421_));
  AOI21_X1   g3372(.A1(new_n2883_), .A2(new_n2884_), .B(new_n2729_), .ZN(new_n3422_));
  OAI21_X1   g3373(.A1(new_n3421_), .A2(new_n3422_), .B(new_n2725_), .ZN(new_n3423_));
  NOR3_X1    g3374(.A1(new_n3421_), .A2(new_n3422_), .A3(new_n2725_), .ZN(new_n3424_));
  INV_X1     g3375(.I(new_n3424_), .ZN(new_n3425_));
  NAND2_X1   g3376(.A1(new_n3425_), .A2(new_n3423_), .ZN(new_n3426_));
  NOR2_X1    g3377(.A1(new_n3417_), .A2(new_n3426_), .ZN(new_n3427_));
  NAND2_X1   g3378(.A1(new_n3179_), .A2(new_n3312_), .ZN(new_n3428_));
  XOR2_X1    g3379(.A1(new_n3428_), .A2(new_n3188_), .Z(new_n3429_));
  AOI21_X1   g3380(.A1(new_n3417_), .A2(new_n3426_), .B(new_n3429_), .ZN(new_n3430_));
  OAI22_X1   g3381(.A1(new_n2697_), .A2(new_n2588_), .B1(new_n56_), .B2(new_n2845_), .ZN(new_n3431_));
  NOR2_X1    g3382(.A1(new_n2858_), .A2(new_n2601_), .ZN(new_n3432_));
  NOR2_X1    g3383(.A1(new_n3432_), .A2(new_n3431_), .ZN(new_n3433_));
  INV_X1     g3384(.I(new_n3433_), .ZN(new_n3434_));
  AOI21_X1   g3385(.A1(new_n2871_), .A2(new_n2865_), .B(new_n2729_), .ZN(new_n3435_));
  OAI21_X1   g3386(.A1(new_n3434_), .A2(new_n3435_), .B(new_n52_), .ZN(new_n3436_));
  NAND2_X1   g3387(.A1(new_n2872_), .A2(new_n2722_), .ZN(new_n3437_));
  NAND3_X1   g3388(.A1(new_n3437_), .A2(new_n2725_), .A3(new_n3433_), .ZN(new_n3438_));
  NAND2_X1   g3389(.A1(new_n3438_), .A2(new_n3436_), .ZN(new_n3439_));
  NOR3_X1    g3390(.A1(new_n3430_), .A2(new_n3427_), .A3(new_n3439_), .ZN(new_n3440_));
  XOR2_X1    g3391(.A1(new_n3317_), .A2(new_n3168_), .Z(new_n3441_));
  XOR2_X1    g3392(.A1(new_n3441_), .A2(new_n3313_), .Z(new_n3442_));
  OAI21_X1   g3393(.A1(new_n3430_), .A2(new_n3427_), .B(new_n3439_), .ZN(new_n3443_));
  OAI21_X1   g3394(.A1(new_n3440_), .A2(new_n3442_), .B(new_n3443_), .ZN(new_n3444_));
  OAI21_X1   g3395(.A1(new_n3350_), .A2(new_n3347_), .B(new_n3355_), .ZN(new_n3445_));
  AOI21_X1   g3396(.A1(new_n3444_), .A2(new_n3445_), .B(new_n3356_), .ZN(new_n3446_));
  OAI22_X1   g3397(.A1(new_n2956_), .A2(new_n2588_), .B1(new_n56_), .B2(new_n2858_), .ZN(new_n3447_));
  NOR2_X1    g3398(.A1(new_n2666_), .A2(new_n2601_), .ZN(new_n3448_));
  NOR2_X1    g3399(.A1(new_n3448_), .A2(new_n3447_), .ZN(new_n3449_));
  NAND2_X1   g3400(.A1(new_n3112_), .A2(new_n3111_), .ZN(new_n3450_));
  NAND2_X1   g3401(.A1(new_n3450_), .A2(new_n2722_), .ZN(new_n3451_));
  AOI21_X1   g3402(.A1(new_n3451_), .A2(new_n3449_), .B(new_n52_), .ZN(new_n3452_));
  NOR2_X1    g3403(.A1(new_n3097_), .A2(new_n2704_), .ZN(new_n3453_));
  NOR2_X1    g3404(.A1(new_n3110_), .A2(new_n2666_), .ZN(new_n3454_));
  NOR2_X1    g3405(.A1(new_n3453_), .A2(new_n3454_), .ZN(new_n3455_));
  NOR2_X1    g3406(.A1(new_n3455_), .A2(new_n2729_), .ZN(new_n3456_));
  NOR4_X1    g3407(.A1(new_n3456_), .A2(new_n2725_), .A3(new_n3447_), .A4(new_n3448_), .ZN(new_n3457_));
  OR2_X2     g3408(.A1(new_n3457_), .A2(new_n3452_), .Z(new_n3458_));
  NOR2_X1    g3409(.A1(new_n3446_), .A2(new_n3458_), .ZN(new_n3459_));
  AOI22_X1   g3410(.A1(new_n3324_), .A2(new_n3322_), .B1(new_n3162_), .B2(new_n3216_), .ZN(new_n3460_));
  NOR4_X1    g3411(.A1(new_n3215_), .A2(new_n3211_), .A3(new_n3161_), .A4(new_n3330_), .ZN(new_n3461_));
  NOR2_X1    g3412(.A1(new_n3460_), .A2(new_n3461_), .ZN(new_n3462_));
  AOI21_X1   g3413(.A1(new_n3446_), .A2(new_n3458_), .B(new_n3462_), .ZN(new_n3463_));
  OAI21_X1   g3414(.A1(new_n3297_), .A2(new_n3300_), .B(new_n3339_), .ZN(new_n3464_));
  OAI21_X1   g3415(.A1(new_n3463_), .A2(new_n3459_), .B(new_n3464_), .ZN(new_n3465_));
  NAND3_X1   g3416(.A1(new_n3250_), .A2(new_n3139_), .A3(new_n3235_), .ZN(new_n3466_));
  INV_X1     g3417(.I(new_n3466_), .ZN(new_n3467_));
  AOI21_X1   g3418(.A1(new_n3250_), .A2(new_n3139_), .B(new_n3235_), .ZN(new_n3468_));
  NOR2_X1    g3419(.A1(new_n3467_), .A2(new_n3468_), .ZN(new_n3469_));
  NAND3_X1   g3420(.A1(new_n3465_), .A2(new_n3341_), .A3(new_n3469_), .ZN(new_n3470_));
  AOI22_X1   g3421(.A1(new_n2613_), .A2(new_n2587_), .B1(new_n55_), .B2(new_n2704_), .ZN(new_n3471_));
  OAI21_X1   g3422(.A1(new_n2611_), .A2(new_n2601_), .B(new_n3471_), .ZN(new_n3472_));
  NOR2_X1    g3423(.A1(new_n3077_), .A2(new_n3078_), .ZN(new_n3473_));
  NOR2_X1    g3424(.A1(new_n3473_), .A2(new_n2729_), .ZN(new_n3474_));
  OAI21_X1   g3425(.A1(new_n3474_), .A2(new_n3472_), .B(new_n2725_), .ZN(new_n3475_));
  OR3_X2     g3426(.A1(new_n3474_), .A2(new_n2725_), .A3(new_n3472_), .Z(new_n3476_));
  NAND2_X1   g3427(.A1(new_n3476_), .A2(new_n3475_), .ZN(new_n3477_));
  OAI21_X1   g3428(.A1(new_n3349_), .A2(new_n3348_), .B(new_n2725_), .ZN(new_n3478_));
  NAND3_X1   g3429(.A1(new_n3346_), .A2(new_n52_), .A3(new_n3345_), .ZN(new_n3479_));
  AOI21_X1   g3430(.A1(new_n3353_), .A2(new_n3322_), .B(new_n3323_), .ZN(new_n3480_));
  NOR3_X1    g3431(.A1(new_n3211_), .A2(new_n3351_), .A3(new_n3214_), .ZN(new_n3481_));
  NOR2_X1    g3432(.A1(new_n3480_), .A2(new_n3481_), .ZN(new_n3482_));
  NAND3_X1   g3433(.A1(new_n3478_), .A2(new_n3479_), .A3(new_n3482_), .ZN(new_n3483_));
  INV_X1     g3434(.I(new_n3368_), .ZN(new_n3484_));
  NOR2_X1    g3435(.A1(new_n3367_), .A2(new_n3360_), .ZN(new_n3485_));
  AOI21_X1   g3436(.A1(new_n3378_), .A2(new_n3380_), .B(new_n52_), .ZN(new_n3486_));
  NOR3_X1    g3437(.A1(new_n3374_), .A2(new_n2725_), .A3(new_n3376_), .ZN(new_n3487_));
  OAI22_X1   g3438(.A1(new_n3487_), .A2(new_n3486_), .B1(new_n3173_), .B2(new_n3485_), .ZN(new_n3488_));
  INV_X1     g3439(.I(new_n3388_), .ZN(new_n3489_));
  NAND3_X1   g3440(.A1(new_n3488_), .A2(new_n3489_), .A3(new_n3484_), .ZN(new_n3490_));
  OAI21_X1   g3441(.A1(new_n3396_), .A2(new_n3392_), .B(new_n2725_), .ZN(new_n3491_));
  NAND3_X1   g3442(.A1(new_n3393_), .A2(new_n3394_), .A3(new_n52_), .ZN(new_n3492_));
  NAND2_X1   g3443(.A1(new_n3492_), .A2(new_n3491_), .ZN(new_n3493_));
  AOI21_X1   g3444(.A1(new_n3488_), .A2(new_n3484_), .B(new_n3489_), .ZN(new_n3494_));
  OAI21_X1   g3445(.A1(new_n3493_), .A2(new_n3494_), .B(new_n3490_), .ZN(new_n3495_));
  OAI21_X1   g3446(.A1(new_n3407_), .A2(new_n3406_), .B(new_n52_), .ZN(new_n3496_));
  NAND3_X1   g3447(.A1(new_n3403_), .A2(new_n2725_), .A3(new_n3402_), .ZN(new_n3497_));
  NAND2_X1   g3448(.A1(new_n3496_), .A2(new_n3497_), .ZN(new_n3498_));
  NAND2_X1   g3449(.A1(new_n3495_), .A2(new_n3498_), .ZN(new_n3499_));
  OAI21_X1   g3450(.A1(new_n3495_), .A2(new_n3498_), .B(new_n3414_), .ZN(new_n3500_));
  NAND2_X1   g3451(.A1(new_n3500_), .A2(new_n3499_), .ZN(new_n3501_));
  INV_X1     g3452(.I(new_n3423_), .ZN(new_n3502_));
  NOR2_X1    g3453(.A1(new_n3502_), .A2(new_n3424_), .ZN(new_n3503_));
  NAND2_X1   g3454(.A1(new_n3501_), .A2(new_n3503_), .ZN(new_n3504_));
  INV_X1     g3455(.I(new_n3429_), .ZN(new_n3505_));
  OAI21_X1   g3456(.A1(new_n3501_), .A2(new_n3503_), .B(new_n3505_), .ZN(new_n3506_));
  AOI21_X1   g3457(.A1(new_n3437_), .A2(new_n3433_), .B(new_n2725_), .ZN(new_n3507_));
  NOR3_X1    g3458(.A1(new_n3434_), .A2(new_n3435_), .A3(new_n52_), .ZN(new_n3508_));
  NOR2_X1    g3459(.A1(new_n3507_), .A2(new_n3508_), .ZN(new_n3509_));
  NAND3_X1   g3460(.A1(new_n3506_), .A2(new_n3504_), .A3(new_n3509_), .ZN(new_n3510_));
  XOR2_X1    g3461(.A1(new_n3441_), .A2(new_n3190_), .Z(new_n3511_));
  AOI21_X1   g3462(.A1(new_n3506_), .A2(new_n3504_), .B(new_n3509_), .ZN(new_n3512_));
  AOI21_X1   g3463(.A1(new_n3510_), .A2(new_n3511_), .B(new_n3512_), .ZN(new_n3513_));
  AOI21_X1   g3464(.A1(new_n3478_), .A2(new_n3479_), .B(new_n3482_), .ZN(new_n3514_));
  OAI21_X1   g3465(.A1(new_n3513_), .A2(new_n3514_), .B(new_n3483_), .ZN(new_n3515_));
  NOR2_X1    g3466(.A1(new_n3457_), .A2(new_n3452_), .ZN(new_n3516_));
  NAND2_X1   g3467(.A1(new_n3515_), .A2(new_n3516_), .ZN(new_n3517_));
  INV_X1     g3468(.I(new_n3462_), .ZN(new_n3518_));
  OAI21_X1   g3469(.A1(new_n3515_), .A2(new_n3516_), .B(new_n3518_), .ZN(new_n3519_));
  OAI21_X1   g3470(.A1(new_n3299_), .A2(new_n3298_), .B(new_n2725_), .ZN(new_n3520_));
  NAND3_X1   g3471(.A1(new_n3296_), .A2(new_n52_), .A3(new_n3287_), .ZN(new_n3521_));
  AOI21_X1   g3472(.A1(new_n3230_), .A2(new_n3337_), .B(new_n3234_), .ZN(new_n3522_));
  NOR3_X1    g3473(.A1(new_n3229_), .A2(new_n3335_), .A3(new_n3233_), .ZN(new_n3523_));
  NOR2_X1    g3474(.A1(new_n3522_), .A2(new_n3523_), .ZN(new_n3524_));
  AOI21_X1   g3475(.A1(new_n3521_), .A2(new_n3520_), .B(new_n3524_), .ZN(new_n3525_));
  AOI21_X1   g3476(.A1(new_n3519_), .A2(new_n3517_), .B(new_n3525_), .ZN(new_n3526_));
  INV_X1     g3477(.I(new_n3468_), .ZN(new_n3527_));
  NAND2_X1   g3478(.A1(new_n3527_), .A2(new_n3466_), .ZN(new_n3528_));
  OAI21_X1   g3479(.A1(new_n3526_), .A2(new_n3340_), .B(new_n3528_), .ZN(new_n3529_));
  NAND2_X1   g3480(.A1(new_n3529_), .A2(new_n3477_), .ZN(new_n3530_));
  XOR2_X1    g3481(.A1(new_n3251_), .A2(new_n3247_), .Z(new_n3531_));
  INV_X1     g3482(.I(new_n3531_), .ZN(new_n3532_));
  NAND3_X1   g3483(.A1(new_n3530_), .A2(new_n3470_), .A3(new_n3532_), .ZN(new_n3533_));
  NOR3_X1    g3484(.A1(new_n3526_), .A2(new_n3340_), .A3(new_n3528_), .ZN(new_n3534_));
  AOI21_X1   g3485(.A1(new_n3477_), .A2(new_n3529_), .B(new_n3534_), .ZN(new_n3535_));
  NOR2_X1    g3486(.A1(new_n2611_), .A2(new_n2588_), .ZN(new_n3536_));
  INV_X1     g3487(.I(new_n3536_), .ZN(new_n3537_));
  INV_X1     g3488(.I(new_n2563_), .ZN(new_n3538_));
  AOI22_X1   g3489(.A1(new_n3538_), .A2(new_n3358_), .B1(new_n55_), .B2(new_n2613_), .ZN(new_n3539_));
  INV_X1     g3490(.I(new_n3539_), .ZN(new_n3540_));
  NOR3_X1    g3491(.A1(new_n2508_), .A2(new_n2562_), .A3(new_n2716_), .ZN(new_n3541_));
  OAI21_X1   g3492(.A1(new_n3541_), .A2(new_n3266_), .B(new_n3262_), .ZN(new_n3542_));
  OR3_X2     g3493(.A1(new_n3541_), .A2(new_n3266_), .A3(new_n3262_), .Z(new_n3543_));
  NAND2_X1   g3494(.A1(new_n3543_), .A2(new_n3542_), .ZN(new_n3544_));
  AOI21_X1   g3495(.A1(new_n3544_), .A2(new_n2722_), .B(new_n3540_), .ZN(new_n3545_));
  NAND3_X1   g3496(.A1(new_n3545_), .A2(new_n2725_), .A3(new_n3537_), .ZN(new_n3546_));
  NAND2_X1   g3497(.A1(new_n3544_), .A2(new_n2722_), .ZN(new_n3547_));
  NAND3_X1   g3498(.A1(new_n3547_), .A2(new_n3537_), .A3(new_n3539_), .ZN(new_n3548_));
  NAND2_X1   g3499(.A1(new_n3548_), .A2(new_n52_), .ZN(new_n3549_));
  NAND2_X1   g3500(.A1(new_n3549_), .A2(new_n3546_), .ZN(new_n3550_));
  OAI21_X1   g3501(.A1(new_n3535_), .A2(new_n3532_), .B(new_n3550_), .ZN(new_n3551_));
  NOR2_X1    g3502(.A1(new_n3278_), .A2(new_n3281_), .ZN(new_n3552_));
  AOI21_X1   g3503(.A1(new_n3551_), .A2(new_n3533_), .B(new_n3552_), .ZN(new_n3553_));
  AOI22_X1   g3504(.A1(new_n3255_), .A2(new_n3241_), .B1(new_n2724_), .B2(new_n2731_), .ZN(new_n3554_));
  NOR3_X1    g3505(.A1(new_n3254_), .A2(new_n3243_), .A3(new_n3242_), .ZN(new_n3555_));
  AOI21_X1   g3506(.A1(new_n3082_), .A2(new_n3084_), .B(new_n3240_), .ZN(new_n3556_));
  NOR3_X1    g3507(.A1(new_n3556_), .A2(new_n2732_), .A3(new_n3555_), .ZN(new_n3557_));
  NOR2_X1    g3508(.A1(new_n3554_), .A2(new_n3557_), .ZN(new_n3558_));
  NOR3_X1    g3509(.A1(new_n3553_), .A2(new_n3283_), .A3(new_n3558_), .ZN(new_n3559_));
  OAI22_X1   g3510(.A1(new_n2598_), .A2(new_n2588_), .B1(new_n2586_), .B2(new_n56_), .ZN(new_n3560_));
  INV_X1     g3511(.I(new_n456_), .ZN(new_n3561_));
  NAND3_X1   g3512(.A1(new_n3561_), .A2(new_n349_), .A3(new_n385_), .ZN(new_n3562_));
  NOR2_X1    g3513(.A1(new_n156_), .A2(new_n357_), .ZN(new_n3563_));
  INV_X1     g3514(.I(new_n3563_), .ZN(new_n3564_));
  NOR3_X1    g3515(.A1(new_n323_), .A2(new_n3564_), .A3(new_n413_), .ZN(new_n3565_));
  NAND4_X1   g3516(.A1(new_n3565_), .A2(new_n311_), .A3(new_n2273_), .A4(new_n1102_), .ZN(new_n3566_));
  NOR4_X1    g3517(.A1(new_n3562_), .A2(new_n334_), .A3(new_n399_), .A4(new_n3566_), .ZN(new_n3567_));
  NOR2_X1    g3518(.A1(new_n2585_), .A2(new_n2594_), .ZN(new_n3568_));
  NOR2_X1    g3519(.A1(new_n3568_), .A2(new_n3567_), .ZN(new_n3569_));
  INV_X1     g3520(.I(new_n3567_), .ZN(new_n3570_));
  NAND3_X1   g3521(.A1(new_n2508_), .A2(new_n2584_), .A3(new_n2595_), .ZN(new_n3571_));
  NOR2_X1    g3522(.A1(new_n3571_), .A2(new_n3570_), .ZN(new_n3572_));
  NOR2_X1    g3523(.A1(new_n3572_), .A2(new_n3569_), .ZN(new_n3573_));
  NOR2_X1    g3524(.A1(new_n3573_), .A2(new_n2601_), .ZN(new_n3574_));
  NOR2_X1    g3525(.A1(new_n3574_), .A2(new_n3560_), .ZN(new_n3575_));
  AOI21_X1   g3526(.A1(new_n2508_), .A2(new_n2584_), .B(new_n2594_), .ZN(new_n3576_));
  NOR2_X1    g3527(.A1(new_n2585_), .A2(new_n2595_), .ZN(new_n3577_));
  NOR2_X1    g3528(.A1(new_n3576_), .A2(new_n3577_), .ZN(new_n3578_));
  OAI21_X1   g3529(.A1(new_n3569_), .A2(new_n3572_), .B(new_n3578_), .ZN(new_n3579_));
  NAND2_X1   g3530(.A1(new_n3571_), .A2(new_n3570_), .ZN(new_n3580_));
  NAND2_X1   g3531(.A1(new_n3568_), .A2(new_n3567_), .ZN(new_n3581_));
  NAND3_X1   g3532(.A1(new_n2598_), .A2(new_n3580_), .A3(new_n3581_), .ZN(new_n3582_));
  NAND2_X1   g3533(.A1(new_n2718_), .A2(new_n2711_), .ZN(new_n3583_));
  AOI22_X1   g3534(.A1(new_n3583_), .A2(new_n2712_), .B1(new_n3579_), .B2(new_n3582_), .ZN(new_n3584_));
  NAND2_X1   g3535(.A1(new_n3579_), .A2(new_n3582_), .ZN(new_n3585_));
  INV_X1     g3536(.I(new_n2711_), .ZN(new_n3586_));
  OAI21_X1   g3537(.A1(new_n2710_), .A2(new_n3586_), .B(new_n2712_), .ZN(new_n3587_));
  NOR2_X1    g3538(.A1(new_n3585_), .A2(new_n3587_), .ZN(new_n3588_));
  OAI21_X1   g3539(.A1(new_n3584_), .A2(new_n3588_), .B(new_n2722_), .ZN(new_n3589_));
  AOI21_X1   g3540(.A1(new_n3589_), .A2(new_n3575_), .B(new_n52_), .ZN(new_n3590_));
  INV_X1     g3541(.I(new_n3575_), .ZN(new_n3591_));
  NAND2_X1   g3542(.A1(new_n3585_), .A2(new_n3587_), .ZN(new_n3592_));
  NAND4_X1   g3543(.A1(new_n3583_), .A2(new_n2712_), .A3(new_n3579_), .A4(new_n3582_), .ZN(new_n3593_));
  AOI21_X1   g3544(.A1(new_n3592_), .A2(new_n3593_), .B(new_n2729_), .ZN(new_n3594_));
  NOR3_X1    g3545(.A1(new_n3594_), .A2(new_n2725_), .A3(new_n3591_), .ZN(new_n3595_));
  NOR2_X1    g3546(.A1(new_n3590_), .A2(new_n3595_), .ZN(new_n3596_));
  INV_X1     g3547(.I(new_n3542_), .ZN(new_n3597_));
  NOR3_X1    g3548(.A1(new_n3541_), .A2(new_n3266_), .A3(new_n3262_), .ZN(new_n3598_));
  NOR2_X1    g3549(.A1(new_n3597_), .A2(new_n3598_), .ZN(new_n3599_));
  NOR2_X1    g3550(.A1(new_n2563_), .A2(new_n3061_), .ZN(new_n3600_));
  NOR2_X1    g3551(.A1(new_n2694_), .A2(new_n3057_), .ZN(new_n3601_));
  NOR2_X1    g3552(.A1(new_n2611_), .A2(new_n3051_), .ZN(new_n3602_));
  NOR3_X1    g3553(.A1(new_n3600_), .A2(new_n3601_), .A3(new_n3602_), .ZN(new_n3603_));
  OAI21_X1   g3554(.A1(new_n3599_), .A2(new_n3074_), .B(new_n3603_), .ZN(new_n3604_));
  OAI22_X1   g3555(.A1(new_n2956_), .A2(new_n2852_), .B1(new_n2858_), .B2(new_n2856_), .ZN(new_n3605_));
  NOR2_X1    g3556(.A1(new_n2666_), .A2(new_n2860_), .ZN(new_n3606_));
  NOR2_X1    g3557(.A1(new_n3606_), .A2(new_n3605_), .ZN(new_n3607_));
  INV_X1     g3558(.I(new_n3607_), .ZN(new_n3608_));
  AOI21_X1   g3559(.A1(new_n3112_), .A2(new_n3111_), .B(new_n2880_), .ZN(new_n3609_));
  OAI21_X1   g3560(.A1(new_n3608_), .A2(new_n3609_), .B(new_n846_), .ZN(new_n3610_));
  OAI21_X1   g3561(.A1(new_n3453_), .A2(new_n3454_), .B(new_n2863_), .ZN(new_n3611_));
  NAND3_X1   g3562(.A1(new_n3611_), .A2(new_n845_), .A3(new_n3607_), .ZN(new_n3612_));
  AOI21_X1   g3563(.A1(new_n3016_), .A2(new_n2992_), .B(new_n3011_), .ZN(new_n3613_));
  NOR2_X1    g3564(.A1(new_n3613_), .A2(new_n3017_), .ZN(new_n3614_));
  NAND2_X1   g3565(.A1(new_n2630_), .A2(new_n2738_), .ZN(new_n3615_));
  NAND2_X1   g3566(.A1(new_n2800_), .A2(new_n2752_), .ZN(new_n3616_));
  NAND2_X1   g3567(.A1(new_n2881_), .A2(new_n2735_), .ZN(new_n3617_));
  NAND3_X1   g3568(.A1(new_n3617_), .A2(new_n3615_), .A3(new_n3616_), .ZN(new_n3618_));
  AOI21_X1   g3569(.A1(new_n2883_), .A2(new_n2884_), .B(new_n2743_), .ZN(new_n3619_));
  OAI21_X1   g3570(.A1(new_n3619_), .A2(new_n3618_), .B(new_n474_), .ZN(new_n3620_));
  NOR3_X1    g3571(.A1(new_n3619_), .A2(new_n474_), .A3(new_n3618_), .ZN(new_n3621_));
  INV_X1     g3572(.I(new_n3621_), .ZN(new_n3622_));
  NOR2_X1    g3573(.A1(new_n2657_), .A2(new_n598_), .ZN(new_n3623_));
  INV_X1     g3574(.I(new_n3623_), .ZN(new_n3624_));
  OAI22_X1   g3575(.A1(new_n2757_), .A2(new_n2815_), .B1(new_n2654_), .B2(new_n3001_), .ZN(new_n3625_));
  AOI21_X1   g3576(.A1(new_n2645_), .A2(new_n2812_), .B(new_n3625_), .ZN(new_n3626_));
  INV_X1     g3577(.I(new_n3626_), .ZN(new_n3627_));
  NOR3_X1    g3578(.A1(new_n2931_), .A2(new_n2929_), .A3(new_n2820_), .ZN(new_n3628_));
  OAI21_X1   g3579(.A1(new_n3627_), .A2(new_n3628_), .B(new_n465_), .ZN(new_n3629_));
  NAND3_X1   g3580(.A1(new_n2773_), .A2(new_n2771_), .A3(new_n2819_), .ZN(new_n3630_));
  NAND3_X1   g3581(.A1(new_n3630_), .A2(new_n598_), .A3(new_n3626_), .ZN(new_n3631_));
  NAND2_X1   g3582(.A1(new_n3629_), .A2(new_n3631_), .ZN(new_n3632_));
  NAND2_X1   g3583(.A1(new_n3632_), .A2(new_n3007_), .ZN(new_n3633_));
  INV_X1     g3584(.I(new_n3007_), .ZN(new_n3634_));
  NAND3_X1   g3585(.A1(new_n3634_), .A2(new_n3629_), .A3(new_n3631_), .ZN(new_n3635_));
  NAND3_X1   g3586(.A1(new_n3633_), .A2(new_n3635_), .A3(new_n3624_), .ZN(new_n3636_));
  AOI21_X1   g3587(.A1(new_n3629_), .A2(new_n3631_), .B(new_n3634_), .ZN(new_n3637_));
  NOR2_X1    g3588(.A1(new_n3632_), .A2(new_n3007_), .ZN(new_n3638_));
  OAI21_X1   g3589(.A1(new_n3637_), .A2(new_n3638_), .B(new_n3623_), .ZN(new_n3639_));
  NAND2_X1   g3590(.A1(new_n3639_), .A2(new_n3636_), .ZN(new_n3640_));
  NAND3_X1   g3591(.A1(new_n3622_), .A2(new_n3620_), .A3(new_n3640_), .ZN(new_n3641_));
  INV_X1     g3592(.I(new_n3618_), .ZN(new_n3642_));
  OAI21_X1   g3593(.A1(new_n3147_), .A2(new_n3146_), .B(new_n2748_), .ZN(new_n3643_));
  AOI21_X1   g3594(.A1(new_n3642_), .A2(new_n3643_), .B(new_n473_), .ZN(new_n3644_));
  NOR3_X1    g3595(.A1(new_n3637_), .A2(new_n3638_), .A3(new_n3623_), .ZN(new_n3645_));
  AOI21_X1   g3596(.A1(new_n3633_), .A2(new_n3635_), .B(new_n3624_), .ZN(new_n3646_));
  NOR2_X1    g3597(.A1(new_n3645_), .A2(new_n3646_), .ZN(new_n3647_));
  OAI21_X1   g3598(.A1(new_n3644_), .A2(new_n3621_), .B(new_n3647_), .ZN(new_n3648_));
  NAND2_X1   g3599(.A1(new_n3641_), .A2(new_n3648_), .ZN(new_n3649_));
  NAND2_X1   g3600(.A1(new_n3614_), .A2(new_n3649_), .ZN(new_n3650_));
  OAI21_X1   g3601(.A1(new_n2995_), .A2(new_n2996_), .B(new_n3012_), .ZN(new_n3651_));
  NAND2_X1   g3602(.A1(new_n3651_), .A2(new_n2997_), .ZN(new_n3652_));
  NOR3_X1    g3603(.A1(new_n3647_), .A2(new_n3644_), .A3(new_n3621_), .ZN(new_n3653_));
  AOI21_X1   g3604(.A1(new_n3622_), .A2(new_n3620_), .B(new_n3640_), .ZN(new_n3654_));
  NOR2_X1    g3605(.A1(new_n3654_), .A2(new_n3653_), .ZN(new_n3655_));
  NAND2_X1   g3606(.A1(new_n3652_), .A2(new_n3655_), .ZN(new_n3656_));
  NAND4_X1   g3607(.A1(new_n3610_), .A2(new_n3612_), .A3(new_n3650_), .A4(new_n3656_), .ZN(new_n3657_));
  AOI21_X1   g3608(.A1(new_n3611_), .A2(new_n3607_), .B(new_n845_), .ZN(new_n3658_));
  NOR3_X1    g3609(.A1(new_n3608_), .A2(new_n3609_), .A3(new_n846_), .ZN(new_n3659_));
  NOR2_X1    g3610(.A1(new_n3652_), .A2(new_n3655_), .ZN(new_n3660_));
  NOR2_X1    g3611(.A1(new_n3614_), .A2(new_n3649_), .ZN(new_n3661_));
  OAI22_X1   g3612(.A1(new_n3659_), .A2(new_n3658_), .B1(new_n3661_), .B2(new_n3660_), .ZN(new_n3662_));
  NAND2_X1   g3613(.A1(new_n3662_), .A2(new_n3657_), .ZN(new_n3663_));
  AOI21_X1   g3614(.A1(new_n2955_), .A2(new_n3020_), .B(new_n3046_), .ZN(new_n3664_));
  NOR2_X1    g3615(.A1(new_n3664_), .A2(new_n3663_), .ZN(new_n3665_));
  NOR4_X1    g3616(.A1(new_n3659_), .A2(new_n3658_), .A3(new_n3661_), .A4(new_n3660_), .ZN(new_n3666_));
  AOI22_X1   g3617(.A1(new_n3610_), .A2(new_n3612_), .B1(new_n3650_), .B2(new_n3656_), .ZN(new_n3667_));
  NOR2_X1    g3618(.A1(new_n3666_), .A2(new_n3667_), .ZN(new_n3668_));
  OAI21_X1   g3619(.A1(new_n3044_), .A2(new_n3045_), .B(new_n3026_), .ZN(new_n3669_));
  NOR2_X1    g3620(.A1(new_n3669_), .A2(new_n3668_), .ZN(new_n3670_));
  OAI21_X1   g3621(.A1(new_n3670_), .A2(new_n3665_), .B(new_n1288_), .ZN(new_n3671_));
  NAND2_X1   g3622(.A1(new_n3669_), .A2(new_n3668_), .ZN(new_n3672_));
  NAND2_X1   g3623(.A1(new_n3664_), .A2(new_n3663_), .ZN(new_n3673_));
  NAND3_X1   g3624(.A1(new_n3672_), .A2(new_n3673_), .A3(new_n1287_), .ZN(new_n3674_));
  NAND3_X1   g3625(.A1(new_n3671_), .A2(new_n3674_), .A3(new_n3604_), .ZN(new_n3675_));
  INV_X1     g3626(.I(new_n3603_), .ZN(new_n3676_));
  AOI21_X1   g3627(.A1(new_n3544_), .A2(new_n3073_), .B(new_n3676_), .ZN(new_n3677_));
  AOI21_X1   g3628(.A1(new_n3672_), .A2(new_n3673_), .B(new_n1287_), .ZN(new_n3678_));
  NOR3_X1    g3629(.A1(new_n3670_), .A2(new_n3665_), .A3(new_n1288_), .ZN(new_n3679_));
  OAI21_X1   g3630(.A1(new_n3678_), .A2(new_n3679_), .B(new_n3677_), .ZN(new_n3680_));
  OAI21_X1   g3631(.A1(new_n3254_), .A2(new_n3243_), .B(new_n3082_), .ZN(new_n3681_));
  NAND3_X1   g3632(.A1(new_n3681_), .A2(new_n3680_), .A3(new_n3675_), .ZN(new_n3682_));
  NAND2_X1   g3633(.A1(new_n3680_), .A2(new_n3675_), .ZN(new_n3683_));
  AOI21_X1   g3634(.A1(new_n3240_), .A2(new_n3084_), .B(new_n3242_), .ZN(new_n3684_));
  NAND2_X1   g3635(.A1(new_n3683_), .A2(new_n3684_), .ZN(new_n3685_));
  AOI21_X1   g3636(.A1(new_n3682_), .A2(new_n3685_), .B(new_n3596_), .ZN(new_n3686_));
  OAI21_X1   g3637(.A1(new_n3594_), .A2(new_n3591_), .B(new_n2725_), .ZN(new_n3687_));
  NAND3_X1   g3638(.A1(new_n3589_), .A2(new_n52_), .A3(new_n3575_), .ZN(new_n3688_));
  NAND2_X1   g3639(.A1(new_n3687_), .A2(new_n3688_), .ZN(new_n3689_));
  NOR3_X1    g3640(.A1(new_n3678_), .A2(new_n3679_), .A3(new_n3677_), .ZN(new_n3690_));
  AOI21_X1   g3641(.A1(new_n3671_), .A2(new_n3674_), .B(new_n3604_), .ZN(new_n3691_));
  NOR3_X1    g3642(.A1(new_n3684_), .A2(new_n3690_), .A3(new_n3691_), .ZN(new_n3692_));
  NOR2_X1    g3643(.A1(new_n3690_), .A2(new_n3691_), .ZN(new_n3693_));
  NOR2_X1    g3644(.A1(new_n3693_), .A2(new_n3681_), .ZN(new_n3694_));
  NOR3_X1    g3645(.A1(new_n3694_), .A2(new_n3689_), .A3(new_n3692_), .ZN(new_n3695_));
  NOR2_X1    g3646(.A1(new_n3686_), .A2(new_n3695_), .ZN(new_n3696_));
  OAI21_X1   g3647(.A1(new_n3559_), .A2(new_n3257_), .B(new_n3696_), .ZN(new_n3697_));
  INV_X1     g3648(.I(new_n3477_), .ZN(new_n3698_));
  AOI21_X1   g3649(.A1(new_n3465_), .A2(new_n3341_), .B(new_n3469_), .ZN(new_n3699_));
  OAI21_X1   g3650(.A1(new_n3698_), .A2(new_n3699_), .B(new_n3470_), .ZN(new_n3700_));
  NOR2_X1    g3651(.A1(new_n3700_), .A2(new_n3531_), .ZN(new_n3701_));
  NOR2_X1    g3652(.A1(new_n3599_), .A2(new_n2729_), .ZN(new_n3702_));
  NOR4_X1    g3653(.A1(new_n3702_), .A2(new_n52_), .A3(new_n3536_), .A4(new_n3540_), .ZN(new_n3703_));
  AOI21_X1   g3654(.A1(new_n3545_), .A2(new_n3537_), .B(new_n2725_), .ZN(new_n3704_));
  NOR2_X1    g3655(.A1(new_n3703_), .A2(new_n3704_), .ZN(new_n3705_));
  AOI21_X1   g3656(.A1(new_n3700_), .A2(new_n3531_), .B(new_n3705_), .ZN(new_n3706_));
  NAND3_X1   g3657(.A1(new_n3238_), .A2(new_n3239_), .A3(new_n3246_), .ZN(new_n3707_));
  OAI21_X1   g3658(.A1(new_n3104_), .A2(new_n3253_), .B(new_n3252_), .ZN(new_n3708_));
  NAND2_X1   g3659(.A1(new_n3708_), .A2(new_n3707_), .ZN(new_n3709_));
  NAND3_X1   g3660(.A1(new_n3709_), .A2(new_n3277_), .A3(new_n3273_), .ZN(new_n3710_));
  OAI21_X1   g3661(.A1(new_n3706_), .A2(new_n3701_), .B(new_n3710_), .ZN(new_n3711_));
  OAI21_X1   g3662(.A1(new_n3555_), .A2(new_n3556_), .B(new_n2732_), .ZN(new_n3712_));
  NAND4_X1   g3663(.A1(new_n3255_), .A2(new_n3241_), .A3(new_n2724_), .A4(new_n2731_), .ZN(new_n3713_));
  NAND2_X1   g3664(.A1(new_n3712_), .A2(new_n3713_), .ZN(new_n3714_));
  NAND3_X1   g3665(.A1(new_n3711_), .A2(new_n3282_), .A3(new_n3714_), .ZN(new_n3715_));
  OAI21_X1   g3666(.A1(new_n3694_), .A2(new_n3692_), .B(new_n3689_), .ZN(new_n3716_));
  NAND3_X1   g3667(.A1(new_n3685_), .A2(new_n3596_), .A3(new_n3682_), .ZN(new_n3717_));
  NAND2_X1   g3668(.A1(new_n3716_), .A2(new_n3717_), .ZN(new_n3718_));
  NAND3_X1   g3669(.A1(new_n3715_), .A2(new_n3718_), .A3(new_n3256_), .ZN(new_n3719_));
  NAND2_X1   g3670(.A1(new_n3697_), .A2(new_n3719_), .ZN(new_n3720_));
  NOR4_X1    g3671(.A1(new_n168_), .A2(new_n201_), .A3(new_n345_), .A4(new_n1120_), .ZN(new_n3721_));
  NAND4_X1   g3672(.A1(new_n3721_), .A2(new_n714_), .A3(new_n431_), .A4(new_n912_), .ZN(new_n3722_));
  NAND4_X1   g3673(.A1(new_n508_), .A2(new_n2461_), .A3(new_n408_), .A4(new_n410_), .ZN(new_n3723_));
  NOR3_X1    g3674(.A1(new_n3722_), .A2(new_n3723_), .A3(new_n2445_), .ZN(new_n3724_));
  NAND3_X1   g3675(.A1(new_n692_), .A2(new_n690_), .A3(new_n694_), .ZN(new_n3725_));
  NOR4_X1    g3676(.A1(new_n3725_), .A2(new_n503_), .A3(new_n856_), .A4(new_n2260_), .ZN(new_n3726_));
  NOR4_X1    g3677(.A1(new_n277_), .A2(new_n263_), .A3(new_n381_), .A4(new_n497_), .ZN(new_n3727_));
  NAND4_X1   g3678(.A1(new_n2362_), .A2(new_n322_), .A3(new_n2345_), .A4(new_n3727_), .ZN(new_n3728_));
  INV_X1     g3679(.I(new_n3728_), .ZN(new_n3729_));
  NAND4_X1   g3680(.A1(new_n3729_), .A2(new_n2394_), .A3(new_n3724_), .A4(new_n3726_), .ZN(new_n3730_));
  NOR3_X1    g3681(.A1(new_n3553_), .A2(new_n3283_), .A3(new_n3714_), .ZN(new_n3731_));
  AOI21_X1   g3682(.A1(new_n3711_), .A2(new_n3282_), .B(new_n3558_), .ZN(new_n3732_));
  OAI21_X1   g3683(.A1(new_n3731_), .A2(new_n3732_), .B(new_n3730_), .ZN(new_n3733_));
  NOR4_X1    g3684(.A1(new_n185_), .A2(new_n267_), .A3(new_n723_), .A4(new_n377_), .ZN(new_n3734_));
  NOR4_X1    g3685(.A1(new_n2255_), .A2(new_n261_), .A3(new_n443_), .A4(new_n580_), .ZN(new_n3735_));
  NAND4_X1   g3686(.A1(new_n3735_), .A2(new_n427_), .A3(new_n1269_), .A4(new_n3734_), .ZN(new_n3736_));
  INV_X1     g3687(.I(new_n3736_), .ZN(new_n3737_));
  NAND4_X1   g3688(.A1(new_n3737_), .A2(new_n674_), .A3(new_n432_), .A4(new_n688_), .ZN(new_n3738_));
  INV_X1     g3689(.I(new_n2437_), .ZN(new_n3739_));
  NOR4_X1    g3690(.A1(new_n179_), .A2(new_n265_), .A3(new_n695_), .A4(new_n402_), .ZN(new_n3740_));
  NAND4_X1   g3691(.A1(new_n3740_), .A2(new_n393_), .A3(new_n350_), .A4(new_n1073_), .ZN(new_n3741_));
  NOR4_X1    g3692(.A1(new_n373_), .A2(new_n177_), .A3(new_n330_), .A4(new_n729_), .ZN(new_n3742_));
  NAND2_X1   g3693(.A1(new_n565_), .A2(new_n429_), .ZN(new_n3743_));
  NOR4_X1    g3694(.A1(new_n3743_), .A2(new_n389_), .A3(new_n745_), .A4(new_n736_), .ZN(new_n3744_));
  NOR4_X1    g3695(.A1(new_n454_), .A2(new_n310_), .A3(new_n341_), .A4(new_n1120_), .ZN(new_n3745_));
  NAND4_X1   g3696(.A1(new_n3744_), .A2(new_n3742_), .A3(new_n3745_), .A4(new_n702_), .ZN(new_n3746_));
  NOR3_X1    g3697(.A1(new_n3739_), .A2(new_n3741_), .A3(new_n3746_), .ZN(new_n3747_));
  INV_X1     g3698(.I(new_n3747_), .ZN(new_n3748_));
  NOR4_X1    g3699(.A1(new_n3738_), .A2(new_n388_), .A3(new_n2574_), .A4(new_n3748_), .ZN(new_n3749_));
  NOR2_X1    g3700(.A1(new_n3733_), .A2(new_n3749_), .ZN(new_n3750_));
  NOR2_X1    g3701(.A1(new_n3750_), .A2(new_n3720_), .ZN(new_n3751_));
  NAND2_X1   g3702(.A1(new_n3733_), .A2(new_n3749_), .ZN(new_n3752_));
  INV_X1     g3703(.I(new_n3752_), .ZN(new_n3753_));
  INV_X1     g3704(.I(new_n2567_), .ZN(new_n3754_));
  NOR4_X1    g3705(.A1(new_n3754_), .A2(new_n269_), .A3(new_n356_), .A4(new_n361_), .ZN(new_n3755_));
  NOR4_X1    g3706(.A1(new_n373_), .A2(new_n196_), .A3(new_n401_), .A4(new_n444_), .ZN(new_n3756_));
  NAND4_X1   g3707(.A1(new_n3755_), .A2(new_n268_), .A3(new_n2261_), .A4(new_n3756_), .ZN(new_n3757_));
  NOR2_X1    g3708(.A1(new_n587_), .A2(new_n573_), .ZN(new_n3758_));
  INV_X1     g3709(.I(new_n3758_), .ZN(new_n3759_));
  NOR2_X1    g3710(.A1(new_n3759_), .A2(new_n2324_), .ZN(new_n3760_));
  NOR4_X1    g3711(.A1(new_n185_), .A2(new_n201_), .A3(new_n377_), .A4(new_n425_), .ZN(new_n3761_));
  NOR2_X1    g3712(.A1(new_n253_), .A2(new_n415_), .ZN(new_n3762_));
  NAND4_X1   g3713(.A1(new_n328_), .A2(new_n3762_), .A3(new_n316_), .A4(new_n788_), .ZN(new_n3763_));
  INV_X1     g3714(.I(new_n3763_), .ZN(new_n3764_));
  NOR4_X1    g3715(.A1(new_n244_), .A2(new_n262_), .A3(new_n345_), .A4(new_n338_), .ZN(new_n3765_));
  NAND4_X1   g3716(.A1(new_n3764_), .A2(new_n3760_), .A3(new_n3761_), .A4(new_n3765_), .ZN(new_n3766_));
  INV_X1     g3717(.I(new_n3766_), .ZN(new_n3767_));
  NOR4_X1    g3718(.A1(new_n187_), .A2(new_n544_), .A3(new_n337_), .A4(new_n400_), .ZN(new_n3768_));
  NAND2_X1   g3719(.A1(new_n3767_), .A2(new_n3768_), .ZN(new_n3769_));
  NOR4_X1    g3720(.A1(new_n586_), .A2(new_n313_), .A3(new_n1440_), .A4(new_n687_), .ZN(new_n3770_));
  NAND2_X1   g3721(.A1(new_n3770_), .A2(new_n2577_), .ZN(new_n3771_));
  NOR4_X1    g3722(.A1(new_n3769_), .A2(new_n571_), .A3(new_n3771_), .A4(new_n3757_), .ZN(new_n3772_));
  NOR3_X1    g3723(.A1(new_n3751_), .A2(new_n3753_), .A3(new_n3772_), .ZN(new_n3773_));
  NOR2_X1    g3724(.A1(new_n3694_), .A2(new_n3692_), .ZN(new_n3774_));
  NAND3_X1   g3725(.A1(new_n3715_), .A2(new_n3256_), .A3(new_n3596_), .ZN(new_n3775_));
  AOI21_X1   g3726(.A1(new_n3715_), .A2(new_n3256_), .B(new_n3596_), .ZN(new_n3776_));
  OAI21_X1   g3727(.A1(new_n3774_), .A2(new_n3776_), .B(new_n3775_), .ZN(new_n3777_));
  NOR2_X1    g3728(.A1(new_n3670_), .A2(new_n3665_), .ZN(new_n3778_));
  NOR2_X1    g3729(.A1(new_n3677_), .A2(new_n1287_), .ZN(new_n3779_));
  NOR2_X1    g3730(.A1(new_n3604_), .A2(new_n1288_), .ZN(new_n3780_));
  OAI21_X1   g3731(.A1(new_n3780_), .A2(new_n3779_), .B(new_n3778_), .ZN(new_n3781_));
  NAND2_X1   g3732(.A1(new_n3682_), .A2(new_n3781_), .ZN(new_n3782_));
  OAI22_X1   g3733(.A1(new_n2563_), .A2(new_n3051_), .B1(new_n2611_), .B2(new_n3057_), .ZN(new_n3783_));
  NOR2_X1    g3734(.A1(new_n2586_), .A2(new_n3061_), .ZN(new_n3784_));
  NOR2_X1    g3735(.A1(new_n3784_), .A2(new_n3783_), .ZN(new_n3785_));
  INV_X1     g3736(.I(new_n3785_), .ZN(new_n3786_));
  AOI21_X1   g3737(.A1(new_n3269_), .A2(new_n3271_), .B(new_n3074_), .ZN(new_n3787_));
  OAI21_X1   g3738(.A1(new_n3787_), .A2(new_n3786_), .B(new_n1288_), .ZN(new_n3788_));
  OAI21_X1   g3739(.A1(new_n3275_), .A2(new_n3274_), .B(new_n3073_), .ZN(new_n3789_));
  NAND3_X1   g3740(.A1(new_n3789_), .A2(new_n1287_), .A3(new_n3785_), .ZN(new_n3790_));
  NAND2_X1   g3741(.A1(new_n3790_), .A2(new_n3788_), .ZN(new_n3791_));
  NOR2_X1    g3742(.A1(new_n2956_), .A2(new_n2856_), .ZN(new_n3792_));
  NOR2_X1    g3743(.A1(new_n2694_), .A2(new_n2860_), .ZN(new_n3793_));
  NOR2_X1    g3744(.A1(new_n2666_), .A2(new_n2852_), .ZN(new_n3794_));
  NOR3_X1    g3745(.A1(new_n3793_), .A2(new_n3792_), .A3(new_n3794_), .ZN(new_n3795_));
  INV_X1     g3746(.I(new_n3795_), .ZN(new_n3796_));
  AOI21_X1   g3747(.A1(new_n3099_), .A2(new_n3094_), .B(new_n2880_), .ZN(new_n3797_));
  OAI21_X1   g3748(.A1(new_n3797_), .A2(new_n3796_), .B(new_n846_), .ZN(new_n3798_));
  OAI21_X1   g3749(.A1(new_n3295_), .A2(new_n3290_), .B(new_n2863_), .ZN(new_n3799_));
  NAND3_X1   g3750(.A1(new_n3799_), .A2(new_n845_), .A3(new_n3795_), .ZN(new_n3800_));
  NAND2_X1   g3751(.A1(new_n3800_), .A2(new_n3798_), .ZN(new_n3801_));
  AOI21_X1   g3752(.A1(new_n3669_), .A2(new_n3657_), .B(new_n3667_), .ZN(new_n3802_));
  OAI21_X1   g3753(.A1(new_n3614_), .A2(new_n3654_), .B(new_n3641_), .ZN(new_n3803_));
  OAI22_X1   g3754(.A1(new_n2697_), .A2(new_n2739_), .B1(new_n2845_), .B2(new_n2768_), .ZN(new_n3804_));
  NOR2_X1    g3755(.A1(new_n2858_), .A2(new_n2736_), .ZN(new_n3805_));
  NOR2_X1    g3756(.A1(new_n3805_), .A2(new_n3804_), .ZN(new_n3806_));
  NAND2_X1   g3757(.A1(new_n2872_), .A2(new_n2748_), .ZN(new_n3807_));
  AOI21_X1   g3758(.A1(new_n3807_), .A2(new_n3806_), .B(new_n473_), .ZN(new_n3808_));
  NAND3_X1   g3759(.A1(new_n3807_), .A2(new_n473_), .A3(new_n3806_), .ZN(new_n3809_));
  INV_X1     g3760(.I(new_n3809_), .ZN(new_n3810_));
  AOI21_X1   g3761(.A1(new_n3629_), .A2(new_n3631_), .B(new_n3623_), .ZN(new_n3811_));
  NAND3_X1   g3762(.A1(new_n3629_), .A2(new_n3631_), .A3(new_n3623_), .ZN(new_n3812_));
  OAI21_X1   g3763(.A1(new_n3811_), .A2(new_n3634_), .B(new_n3812_), .ZN(new_n3813_));
  OAI22_X1   g3764(.A1(new_n2679_), .A2(new_n2815_), .B1(new_n2757_), .B2(new_n3001_), .ZN(new_n3814_));
  AOI21_X1   g3765(.A1(new_n2800_), .A2(new_n2812_), .B(new_n3814_), .ZN(new_n3815_));
  OAI21_X1   g3766(.A1(new_n2807_), .A2(new_n2808_), .B(new_n2819_), .ZN(new_n3816_));
  NAND2_X1   g3767(.A1(new_n3816_), .A2(new_n3815_), .ZN(new_n3817_));
  NOR2_X1    g3768(.A1(new_n3813_), .A2(new_n3817_), .ZN(new_n3818_));
  INV_X1     g3769(.I(new_n3818_), .ZN(new_n3819_));
  NAND2_X1   g3770(.A1(new_n3813_), .A2(new_n3817_), .ZN(new_n3820_));
  NOR2_X1    g3771(.A1(new_n2682_), .A2(new_n598_), .ZN(new_n3821_));
  AOI21_X1   g3772(.A1(new_n3819_), .A2(new_n3820_), .B(new_n3821_), .ZN(new_n3822_));
  INV_X1     g3773(.I(new_n3820_), .ZN(new_n3823_));
  INV_X1     g3774(.I(new_n3821_), .ZN(new_n3824_));
  NOR3_X1    g3775(.A1(new_n3823_), .A2(new_n3818_), .A3(new_n3824_), .ZN(new_n3825_));
  NOR2_X1    g3776(.A1(new_n3822_), .A2(new_n3825_), .ZN(new_n3826_));
  NOR3_X1    g3777(.A1(new_n3826_), .A2(new_n3810_), .A3(new_n3808_), .ZN(new_n3827_));
  INV_X1     g3778(.I(new_n3808_), .ZN(new_n3828_));
  OR2_X2     g3779(.A1(new_n3822_), .A2(new_n3825_), .Z(new_n3829_));
  AOI21_X1   g3780(.A1(new_n3828_), .A2(new_n3809_), .B(new_n3829_), .ZN(new_n3830_));
  NOR3_X1    g3781(.A1(new_n3830_), .A2(new_n3803_), .A3(new_n3827_), .ZN(new_n3831_));
  AOI21_X1   g3782(.A1(new_n3652_), .A2(new_n3648_), .B(new_n3653_), .ZN(new_n3832_));
  NAND3_X1   g3783(.A1(new_n3829_), .A2(new_n3828_), .A3(new_n3809_), .ZN(new_n3833_));
  OAI21_X1   g3784(.A1(new_n3810_), .A2(new_n3808_), .B(new_n3826_), .ZN(new_n3834_));
  AOI21_X1   g3785(.A1(new_n3833_), .A2(new_n3834_), .B(new_n3832_), .ZN(new_n3835_));
  NOR2_X1    g3786(.A1(new_n3831_), .A2(new_n3835_), .ZN(new_n3836_));
  INV_X1     g3787(.I(new_n3836_), .ZN(new_n3837_));
  NOR2_X1    g3788(.A1(new_n3802_), .A2(new_n3837_), .ZN(new_n3838_));
  OAI21_X1   g3789(.A1(new_n3664_), .A2(new_n3663_), .B(new_n3662_), .ZN(new_n3839_));
  NOR2_X1    g3790(.A1(new_n3839_), .A2(new_n3836_), .ZN(new_n3840_));
  NOR3_X1    g3791(.A1(new_n3840_), .A2(new_n3838_), .A3(new_n3801_), .ZN(new_n3841_));
  INV_X1     g3792(.I(new_n3801_), .ZN(new_n3842_));
  NAND2_X1   g3793(.A1(new_n3839_), .A2(new_n3836_), .ZN(new_n3843_));
  NAND2_X1   g3794(.A1(new_n3802_), .A2(new_n3837_), .ZN(new_n3844_));
  AOI21_X1   g3795(.A1(new_n3843_), .A2(new_n3844_), .B(new_n3842_), .ZN(new_n3845_));
  NOR2_X1    g3796(.A1(new_n3845_), .A2(new_n3841_), .ZN(new_n3846_));
  XOR2_X1    g3797(.A1(new_n3846_), .A2(new_n3791_), .Z(new_n3847_));
  NAND2_X1   g3798(.A1(new_n3847_), .A2(new_n3782_), .ZN(new_n3848_));
  INV_X1     g3799(.I(new_n3778_), .ZN(new_n3849_));
  NAND2_X1   g3800(.A1(new_n3604_), .A2(new_n1288_), .ZN(new_n3850_));
  NAND2_X1   g3801(.A1(new_n3677_), .A2(new_n1287_), .ZN(new_n3851_));
  AOI21_X1   g3802(.A1(new_n3850_), .A2(new_n3851_), .B(new_n3849_), .ZN(new_n3852_));
  NOR2_X1    g3803(.A1(new_n3692_), .A2(new_n3852_), .ZN(new_n3853_));
  NAND3_X1   g3804(.A1(new_n3843_), .A2(new_n3844_), .A3(new_n3842_), .ZN(new_n3854_));
  OAI21_X1   g3805(.A1(new_n3840_), .A2(new_n3838_), .B(new_n3801_), .ZN(new_n3855_));
  NAND2_X1   g3806(.A1(new_n3855_), .A2(new_n3854_), .ZN(new_n3856_));
  XOR2_X1    g3807(.A1(new_n3791_), .A2(new_n3856_), .Z(new_n3857_));
  NAND2_X1   g3808(.A1(new_n3857_), .A2(new_n3853_), .ZN(new_n3858_));
  NAND2_X1   g3809(.A1(new_n3580_), .A2(new_n3581_), .ZN(new_n3859_));
  AOI22_X1   g3810(.A1(new_n3859_), .A2(new_n2587_), .B1(new_n55_), .B2(new_n3578_), .ZN(new_n3860_));
  NOR4_X1    g3811(.A1(new_n326_), .A2(new_n164_), .A3(new_n345_), .A4(new_n415_), .ZN(new_n3861_));
  AND3_X2    g3812(.A1(new_n358_), .A2(new_n385_), .A3(new_n441_), .Z(new_n3862_));
  NOR2_X1    g3813(.A1(new_n456_), .A2(new_n727_), .ZN(new_n3863_));
  AND3_X2    g3814(.A1(new_n3861_), .A2(new_n3862_), .A3(new_n3863_), .Z(new_n3864_));
  INV_X1     g3815(.I(new_n3864_), .ZN(new_n3865_));
  NOR2_X1    g3816(.A1(new_n3572_), .A2(new_n3865_), .ZN(new_n3866_));
  NOR2_X1    g3817(.A1(new_n3581_), .A2(new_n3864_), .ZN(new_n3867_));
  NOR2_X1    g3818(.A1(new_n3866_), .A2(new_n3867_), .ZN(new_n3868_));
  INV_X1     g3819(.I(new_n3868_), .ZN(new_n3869_));
  OAI21_X1   g3820(.A1(new_n3869_), .A2(new_n2601_), .B(new_n3860_), .ZN(new_n3870_));
  INV_X1     g3821(.I(new_n3870_), .ZN(new_n3871_));
  NAND2_X1   g3822(.A1(new_n2586_), .A2(new_n2717_), .ZN(new_n3872_));
  NAND2_X1   g3823(.A1(new_n3872_), .A2(new_n3578_), .ZN(new_n3873_));
  NAND2_X1   g3824(.A1(new_n3873_), .A2(new_n3573_), .ZN(new_n3874_));
  OAI21_X1   g3825(.A1(new_n2710_), .A2(new_n2586_), .B(new_n2598_), .ZN(new_n3875_));
  NAND2_X1   g3826(.A1(new_n3875_), .A2(new_n3859_), .ZN(new_n3876_));
  NAND2_X1   g3827(.A1(new_n3876_), .A2(new_n3874_), .ZN(new_n3877_));
  NOR2_X1    g3828(.A1(new_n3877_), .A2(new_n3868_), .ZN(new_n3878_));
  INV_X1     g3829(.I(new_n3878_), .ZN(new_n3879_));
  NAND2_X1   g3830(.A1(new_n3877_), .A2(new_n3868_), .ZN(new_n3880_));
  NAND2_X1   g3831(.A1(new_n3879_), .A2(new_n3880_), .ZN(new_n3881_));
  NAND2_X1   g3832(.A1(new_n3881_), .A2(new_n2722_), .ZN(new_n3882_));
  AOI21_X1   g3833(.A1(new_n3882_), .A2(new_n3871_), .B(new_n52_), .ZN(new_n3883_));
  INV_X1     g3834(.I(new_n3880_), .ZN(new_n3884_));
  NOR2_X1    g3835(.A1(new_n3884_), .A2(new_n3878_), .ZN(new_n3885_));
  NOR2_X1    g3836(.A1(new_n3885_), .A2(new_n2729_), .ZN(new_n3886_));
  NOR3_X1    g3837(.A1(new_n3886_), .A2(new_n2725_), .A3(new_n3870_), .ZN(new_n3887_));
  NOR2_X1    g3838(.A1(new_n3887_), .A2(new_n3883_), .ZN(new_n3888_));
  NAND3_X1   g3839(.A1(new_n3888_), .A2(new_n3848_), .A3(new_n3858_), .ZN(new_n3889_));
  NOR2_X1    g3840(.A1(new_n3857_), .A2(new_n3853_), .ZN(new_n3890_));
  NOR2_X1    g3841(.A1(new_n3847_), .A2(new_n3782_), .ZN(new_n3891_));
  OAI21_X1   g3842(.A1(new_n3886_), .A2(new_n3870_), .B(new_n2725_), .ZN(new_n3892_));
  NAND3_X1   g3843(.A1(new_n3882_), .A2(new_n52_), .A3(new_n3871_), .ZN(new_n3893_));
  NAND2_X1   g3844(.A1(new_n3892_), .A2(new_n3893_), .ZN(new_n3894_));
  OAI21_X1   g3845(.A1(new_n3891_), .A2(new_n3890_), .B(new_n3894_), .ZN(new_n3895_));
  NAND2_X1   g3846(.A1(new_n3895_), .A2(new_n3889_), .ZN(new_n3896_));
  XOR2_X1    g3847(.A1(new_n3777_), .A2(new_n3896_), .Z(new_n3897_));
  OAI21_X1   g3848(.A1(new_n3751_), .A2(new_n3753_), .B(new_n3772_), .ZN(new_n3898_));
  OAI21_X1   g3849(.A1(new_n3897_), .A2(new_n3773_), .B(new_n3898_), .ZN(new_n3899_));
  NOR2_X1    g3850(.A1(new_n2563_), .A2(new_n3057_), .ZN(new_n3900_));
  NOR2_X1    g3851(.A1(new_n2586_), .A2(new_n3051_), .ZN(new_n3901_));
  NOR2_X1    g3852(.A1(new_n2598_), .A2(new_n3061_), .ZN(new_n3902_));
  NOR3_X1    g3853(.A1(new_n3902_), .A2(new_n3901_), .A3(new_n3900_), .ZN(new_n3903_));
  NAND2_X1   g3854(.A1(new_n2727_), .A2(new_n2728_), .ZN(new_n3904_));
  NAND2_X1   g3855(.A1(new_n3904_), .A2(new_n3073_), .ZN(new_n3905_));
  AOI21_X1   g3856(.A1(new_n3905_), .A2(new_n3903_), .B(new_n1287_), .ZN(new_n3906_));
  INV_X1     g3857(.I(new_n3903_), .ZN(new_n3907_));
  NOR2_X1    g3858(.A1(new_n2720_), .A2(new_n2713_), .ZN(new_n3908_));
  NOR2_X1    g3859(.A1(new_n3908_), .A2(new_n3074_), .ZN(new_n3909_));
  NOR3_X1    g3860(.A1(new_n3909_), .A2(new_n1288_), .A3(new_n3907_), .ZN(new_n3910_));
  NOR2_X1    g3861(.A1(new_n3910_), .A2(new_n3906_), .ZN(new_n3911_));
  OAI22_X1   g3862(.A1(new_n2694_), .A2(new_n2852_), .B1(new_n2666_), .B2(new_n2856_), .ZN(new_n3912_));
  NOR2_X1    g3863(.A1(new_n2611_), .A2(new_n2860_), .ZN(new_n3913_));
  NOR2_X1    g3864(.A1(new_n3913_), .A2(new_n3912_), .ZN(new_n3914_));
  INV_X1     g3865(.I(new_n3914_), .ZN(new_n3915_));
  AOI21_X1   g3866(.A1(new_n3072_), .A2(new_n3068_), .B(new_n2880_), .ZN(new_n3916_));
  OAI21_X1   g3867(.A1(new_n3916_), .A2(new_n3915_), .B(new_n845_), .ZN(new_n3917_));
  OAI21_X1   g3868(.A1(new_n3077_), .A2(new_n3078_), .B(new_n2863_), .ZN(new_n3918_));
  NAND3_X1   g3869(.A1(new_n3918_), .A2(new_n846_), .A3(new_n3914_), .ZN(new_n3919_));
  NOR2_X1    g3870(.A1(new_n2956_), .A2(new_n2736_), .ZN(new_n3920_));
  NOR2_X1    g3871(.A1(new_n2697_), .A2(new_n2768_), .ZN(new_n3921_));
  NOR2_X1    g3872(.A1(new_n2858_), .A2(new_n2739_), .ZN(new_n3922_));
  NOR3_X1    g3873(.A1(new_n3920_), .A2(new_n3921_), .A3(new_n3922_), .ZN(new_n3923_));
  INV_X1     g3874(.I(new_n3923_), .ZN(new_n3924_));
  AOI21_X1   g3875(.A1(new_n2968_), .A2(new_n2964_), .B(new_n2743_), .ZN(new_n3925_));
  OAI21_X1   g3876(.A1(new_n3925_), .A2(new_n3924_), .B(new_n474_), .ZN(new_n3926_));
  NAND2_X1   g3877(.A1(new_n2976_), .A2(new_n2748_), .ZN(new_n3927_));
  NAND3_X1   g3878(.A1(new_n3927_), .A2(new_n473_), .A3(new_n3923_), .ZN(new_n3928_));
  OAI22_X1   g3879(.A1(new_n2792_), .A2(new_n2815_), .B1(new_n2679_), .B2(new_n3001_), .ZN(new_n3929_));
  NOR2_X1    g3880(.A1(new_n2845_), .A2(new_n3003_), .ZN(new_n3930_));
  NOR2_X1    g3881(.A1(new_n3930_), .A2(new_n3929_), .ZN(new_n3931_));
  OAI21_X1   g3882(.A1(new_n2989_), .A2(new_n2988_), .B(new_n2819_), .ZN(new_n3932_));
  NOR2_X1    g3883(.A1(new_n2754_), .A2(new_n598_), .ZN(new_n3933_));
  AOI21_X1   g3884(.A1(new_n3932_), .A2(new_n3931_), .B(new_n3933_), .ZN(new_n3934_));
  NAND3_X1   g3885(.A1(new_n3932_), .A2(new_n3931_), .A3(new_n3933_), .ZN(new_n3935_));
  INV_X1     g3886(.I(new_n3935_), .ZN(new_n3936_));
  NOR2_X1    g3887(.A1(new_n3936_), .A2(new_n3934_), .ZN(new_n3937_));
  INV_X1     g3888(.I(new_n3817_), .ZN(new_n3938_));
  AOI21_X1   g3889(.A1(new_n3813_), .A2(new_n3938_), .B(new_n3824_), .ZN(new_n3939_));
  NAND3_X1   g3890(.A1(new_n3816_), .A2(new_n465_), .A3(new_n3815_), .ZN(new_n3940_));
  INV_X1     g3891(.I(new_n3940_), .ZN(new_n3941_));
  AOI21_X1   g3892(.A1(new_n3813_), .A2(new_n3817_), .B(new_n3941_), .ZN(new_n3942_));
  NOR3_X1    g3893(.A1(new_n3937_), .A2(new_n3942_), .A3(new_n3939_), .ZN(new_n3943_));
  INV_X1     g3894(.I(new_n3934_), .ZN(new_n3944_));
  NAND2_X1   g3895(.A1(new_n3944_), .A2(new_n3935_), .ZN(new_n3945_));
  NOR2_X1    g3896(.A1(new_n3942_), .A2(new_n3939_), .ZN(new_n3946_));
  NOR2_X1    g3897(.A1(new_n3946_), .A2(new_n3945_), .ZN(new_n3947_));
  NOR2_X1    g3898(.A1(new_n3947_), .A2(new_n3943_), .ZN(new_n3948_));
  INV_X1     g3899(.I(new_n3948_), .ZN(new_n3949_));
  NAND3_X1   g3900(.A1(new_n3926_), .A2(new_n3928_), .A3(new_n3949_), .ZN(new_n3950_));
  AOI21_X1   g3901(.A1(new_n3927_), .A2(new_n3923_), .B(new_n473_), .ZN(new_n3951_));
  INV_X1     g3902(.I(new_n3928_), .ZN(new_n3952_));
  OAI21_X1   g3903(.A1(new_n3952_), .A2(new_n3951_), .B(new_n3948_), .ZN(new_n3953_));
  AOI21_X1   g3904(.A1(new_n3803_), .A2(new_n3834_), .B(new_n3827_), .ZN(new_n3954_));
  NAND3_X1   g3905(.A1(new_n3953_), .A2(new_n3950_), .A3(new_n3954_), .ZN(new_n3955_));
  INV_X1     g3906(.I(new_n3950_), .ZN(new_n3956_));
  AOI21_X1   g3907(.A1(new_n3926_), .A2(new_n3928_), .B(new_n3949_), .ZN(new_n3957_));
  OAI21_X1   g3908(.A1(new_n3830_), .A2(new_n3832_), .B(new_n3833_), .ZN(new_n3958_));
  OAI21_X1   g3909(.A1(new_n3956_), .A2(new_n3957_), .B(new_n3958_), .ZN(new_n3959_));
  NAND4_X1   g3910(.A1(new_n3917_), .A2(new_n3959_), .A3(new_n3919_), .A4(new_n3955_), .ZN(new_n3960_));
  AOI21_X1   g3911(.A1(new_n3918_), .A2(new_n3914_), .B(new_n846_), .ZN(new_n3961_));
  NOR3_X1    g3912(.A1(new_n3916_), .A2(new_n3915_), .A3(new_n845_), .ZN(new_n3962_));
  NOR3_X1    g3913(.A1(new_n3956_), .A2(new_n3958_), .A3(new_n3957_), .ZN(new_n3963_));
  AOI21_X1   g3914(.A1(new_n3953_), .A2(new_n3950_), .B(new_n3954_), .ZN(new_n3964_));
  OAI22_X1   g3915(.A1(new_n3962_), .A2(new_n3961_), .B1(new_n3963_), .B2(new_n3964_), .ZN(new_n3965_));
  NAND2_X1   g3916(.A1(new_n3965_), .A2(new_n3960_), .ZN(new_n3966_));
  OAI21_X1   g3917(.A1(new_n3801_), .A2(new_n3838_), .B(new_n3844_), .ZN(new_n3967_));
  NOR2_X1    g3918(.A1(new_n3967_), .A2(new_n3966_), .ZN(new_n3968_));
  NOR4_X1    g3919(.A1(new_n3962_), .A2(new_n3961_), .A3(new_n3963_), .A4(new_n3964_), .ZN(new_n3969_));
  AOI22_X1   g3920(.A1(new_n3917_), .A2(new_n3919_), .B1(new_n3959_), .B2(new_n3955_), .ZN(new_n3970_));
  NOR2_X1    g3921(.A1(new_n3970_), .A2(new_n3969_), .ZN(new_n3971_));
  AOI21_X1   g3922(.A1(new_n3839_), .A2(new_n3836_), .B(new_n3801_), .ZN(new_n3972_));
  NOR2_X1    g3923(.A1(new_n3972_), .A2(new_n3840_), .ZN(new_n3973_));
  NOR2_X1    g3924(.A1(new_n3973_), .A2(new_n3971_), .ZN(new_n3974_));
  OAI21_X1   g3925(.A1(new_n3968_), .A2(new_n3974_), .B(new_n3911_), .ZN(new_n3975_));
  OAI21_X1   g3926(.A1(new_n3909_), .A2(new_n3907_), .B(new_n1288_), .ZN(new_n3976_));
  NAND3_X1   g3927(.A1(new_n3905_), .A2(new_n1287_), .A3(new_n3903_), .ZN(new_n3977_));
  NAND2_X1   g3928(.A1(new_n3976_), .A2(new_n3977_), .ZN(new_n3978_));
  NOR2_X1    g3929(.A1(new_n3968_), .A2(new_n3974_), .ZN(new_n3979_));
  NAND2_X1   g3930(.A1(new_n3979_), .A2(new_n3978_), .ZN(new_n3980_));
  NAND3_X1   g3931(.A1(new_n3980_), .A2(new_n3975_), .A3(new_n2725_), .ZN(new_n3981_));
  NOR2_X1    g3932(.A1(new_n3979_), .A2(new_n3978_), .ZN(new_n3982_));
  NOR3_X1    g3933(.A1(new_n3911_), .A2(new_n3968_), .A3(new_n3974_), .ZN(new_n3983_));
  OAI21_X1   g3934(.A1(new_n3982_), .A2(new_n3983_), .B(new_n52_), .ZN(new_n3984_));
  NAND2_X1   g3935(.A1(new_n3981_), .A2(new_n3984_), .ZN(new_n3985_));
  AOI22_X1   g3936(.A1(new_n3868_), .A2(new_n2587_), .B1(new_n55_), .B2(new_n3859_), .ZN(new_n3986_));
  NOR4_X1    g3937(.A1(new_n197_), .A2(new_n310_), .A3(new_n723_), .A4(new_n245_), .ZN(new_n3987_));
  NOR3_X1    g3938(.A1(new_n3759_), .A2(new_n321_), .A3(new_n356_), .ZN(new_n3988_));
  NAND3_X1   g3939(.A1(new_n3988_), .A2(new_n553_), .A3(new_n3987_), .ZN(new_n3989_));
  INV_X1     g3940(.I(new_n3989_), .ZN(new_n3990_));
  INV_X1     g3941(.I(new_n558_), .ZN(new_n3991_));
  INV_X1     g3942(.I(new_n259_), .ZN(new_n3992_));
  NOR4_X1    g3943(.A1(new_n187_), .A2(new_n201_), .A3(new_n253_), .A4(new_n338_), .ZN(new_n3993_));
  NAND4_X1   g3944(.A1(new_n3993_), .A2(new_n889_), .A3(new_n3992_), .A4(new_n2466_), .ZN(new_n3994_));
  NAND2_X1   g3945(.A1(new_n2321_), .A2(new_n369_), .ZN(new_n3995_));
  NOR4_X1    g3946(.A1(new_n3994_), .A2(new_n2267_), .A3(new_n3991_), .A4(new_n3995_), .ZN(new_n3996_));
  NAND3_X1   g3947(.A1(new_n3990_), .A2(new_n1118_), .A3(new_n3996_), .ZN(new_n3997_));
  OAI21_X1   g3948(.A1(new_n3581_), .A2(new_n3865_), .B(new_n3997_), .ZN(new_n3998_));
  INV_X1     g3949(.I(new_n3997_), .ZN(new_n3999_));
  NAND3_X1   g3950(.A1(new_n3572_), .A2(new_n3864_), .A3(new_n3999_), .ZN(new_n4000_));
  NAND2_X1   g3951(.A1(new_n4000_), .A2(new_n3998_), .ZN(new_n4001_));
  INV_X1     g3952(.I(new_n4001_), .ZN(new_n4002_));
  OAI21_X1   g3953(.A1(new_n2601_), .A2(new_n4002_), .B(new_n3986_), .ZN(new_n4003_));
  NAND2_X1   g3954(.A1(new_n4001_), .A2(new_n3859_), .ZN(new_n4004_));
  NAND2_X1   g3955(.A1(new_n4002_), .A2(new_n3876_), .ZN(new_n4005_));
  NAND3_X1   g3956(.A1(new_n4005_), .A2(new_n3869_), .A3(new_n4004_), .ZN(new_n4006_));
  AOI21_X1   g3957(.A1(new_n3578_), .A2(new_n3872_), .B(new_n3859_), .ZN(new_n4007_));
  AOI21_X1   g3958(.A1(new_n3859_), .A2(new_n3875_), .B(new_n4007_), .ZN(new_n4008_));
  AOI21_X1   g3959(.A1(new_n2718_), .A2(new_n2604_), .B(new_n3578_), .ZN(new_n4009_));
  NOR2_X1    g3960(.A1(new_n4007_), .A2(new_n4009_), .ZN(new_n4010_));
  NAND3_X1   g3961(.A1(new_n3573_), .A2(new_n4000_), .A3(new_n3998_), .ZN(new_n4011_));
  OAI21_X1   g3962(.A1(new_n4010_), .A2(new_n4011_), .B(new_n4004_), .ZN(new_n4012_));
  AOI22_X1   g3963(.A1(new_n4012_), .A2(new_n3868_), .B1(new_n4008_), .B2(new_n4001_), .ZN(new_n4013_));
  AOI21_X1   g3964(.A1(new_n4013_), .A2(new_n4006_), .B(new_n2729_), .ZN(new_n4014_));
  NOR2_X1    g3965(.A1(new_n4014_), .A2(new_n4003_), .ZN(new_n4015_));
  INV_X1     g3966(.I(new_n3791_), .ZN(new_n4016_));
  NOR3_X1    g3967(.A1(new_n3692_), .A2(new_n3852_), .A3(new_n3856_), .ZN(new_n4017_));
  OAI21_X1   g3968(.A1(new_n3692_), .A2(new_n3852_), .B(new_n3856_), .ZN(new_n4018_));
  AOI21_X1   g3969(.A1(new_n4016_), .A2(new_n4018_), .B(new_n4017_), .ZN(new_n4019_));
  NOR2_X1    g3970(.A1(new_n4019_), .A2(new_n4015_), .ZN(new_n4020_));
  INV_X1     g3971(.I(new_n4015_), .ZN(new_n4021_));
  NAND3_X1   g3972(.A1(new_n3682_), .A2(new_n3781_), .A3(new_n3846_), .ZN(new_n4022_));
  AOI21_X1   g3973(.A1(new_n3682_), .A2(new_n3781_), .B(new_n3846_), .ZN(new_n4023_));
  OAI21_X1   g3974(.A1(new_n3791_), .A2(new_n4023_), .B(new_n4022_), .ZN(new_n4024_));
  NOR2_X1    g3975(.A1(new_n4024_), .A2(new_n4021_), .ZN(new_n4025_));
  OAI21_X1   g3976(.A1(new_n4020_), .A2(new_n4025_), .B(new_n3985_), .ZN(new_n4026_));
  NOR3_X1    g3977(.A1(new_n3982_), .A2(new_n3983_), .A3(new_n52_), .ZN(new_n4027_));
  AOI21_X1   g3978(.A1(new_n3980_), .A2(new_n3975_), .B(new_n2725_), .ZN(new_n4028_));
  NOR2_X1    g3979(.A1(new_n4028_), .A2(new_n4027_), .ZN(new_n4029_));
  NAND2_X1   g3980(.A1(new_n4024_), .A2(new_n4021_), .ZN(new_n4030_));
  NAND2_X1   g3981(.A1(new_n4019_), .A2(new_n4015_), .ZN(new_n4031_));
  NAND3_X1   g3982(.A1(new_n4029_), .A2(new_n4031_), .A3(new_n4030_), .ZN(new_n4032_));
  NAND2_X1   g3983(.A1(new_n4026_), .A2(new_n4032_), .ZN(new_n4033_));
  NOR3_X1    g3984(.A1(new_n3891_), .A2(new_n3894_), .A3(new_n3890_), .ZN(new_n4034_));
  OAI21_X1   g3985(.A1(new_n3777_), .A2(new_n4034_), .B(new_n3895_), .ZN(new_n4035_));
  NOR2_X1    g3986(.A1(new_n4035_), .A2(new_n4033_), .ZN(new_n4036_));
  AOI21_X1   g3987(.A1(new_n4030_), .A2(new_n4031_), .B(new_n4029_), .ZN(new_n4037_));
  NOR3_X1    g3988(.A1(new_n3985_), .A2(new_n4020_), .A3(new_n4025_), .ZN(new_n4038_));
  NOR2_X1    g3989(.A1(new_n4037_), .A2(new_n4038_), .ZN(new_n4039_));
  INV_X1     g3990(.I(new_n3774_), .ZN(new_n4040_));
  OAI21_X1   g3991(.A1(new_n3559_), .A2(new_n3257_), .B(new_n3689_), .ZN(new_n4041_));
  NAND2_X1   g3992(.A1(new_n4041_), .A2(new_n4040_), .ZN(new_n4042_));
  NAND3_X1   g3993(.A1(new_n4042_), .A2(new_n3775_), .A3(new_n3889_), .ZN(new_n4043_));
  AOI21_X1   g3994(.A1(new_n4043_), .A2(new_n3895_), .B(new_n4039_), .ZN(new_n4044_));
  NOR2_X1    g3995(.A1(new_n4036_), .A2(new_n4044_), .ZN(new_n4045_));
  INV_X1     g3996(.I(new_n2368_), .ZN(new_n4046_));
  NOR2_X1    g3997(.A1(new_n718_), .A2(new_n267_), .ZN(new_n4047_));
  NAND4_X1   g3998(.A1(new_n4047_), .A2(new_n3758_), .A3(new_n563_), .A4(new_n702_), .ZN(new_n4048_));
  NAND2_X1   g3999(.A1(new_n2567_), .A2(new_n1077_), .ZN(new_n4049_));
  NOR4_X1    g4000(.A1(new_n4048_), .A2(new_n499_), .A3(new_n2344_), .A4(new_n4049_), .ZN(new_n4050_));
  NAND3_X1   g4001(.A1(new_n4046_), .A2(new_n523_), .A3(new_n4050_), .ZN(new_n4051_));
  NAND2_X1   g4002(.A1(new_n4045_), .A2(new_n4051_), .ZN(new_n4052_));
  INV_X1     g4003(.I(new_n4051_), .ZN(new_n4053_));
  OAI21_X1   g4004(.A1(new_n4036_), .A2(new_n4044_), .B(new_n4053_), .ZN(new_n4054_));
  NAND2_X1   g4005(.A1(new_n4052_), .A2(new_n4054_), .ZN(new_n4055_));
  INV_X1     g4006(.I(new_n3772_), .ZN(new_n4056_));
  XOR2_X1    g4007(.A1(new_n3896_), .A2(new_n4056_), .Z(new_n4057_));
  NOR3_X1    g4008(.A1(new_n3559_), .A2(new_n3257_), .A3(new_n3689_), .ZN(new_n4058_));
  AOI21_X1   g4009(.A1(new_n4040_), .A2(new_n4041_), .B(new_n4058_), .ZN(new_n4059_));
  NOR3_X1    g4010(.A1(new_n3751_), .A2(new_n3753_), .A3(new_n4059_), .ZN(new_n4060_));
  NAND3_X1   g4011(.A1(new_n3711_), .A2(new_n3282_), .A3(new_n3558_), .ZN(new_n4061_));
  OAI21_X1   g4012(.A1(new_n3553_), .A2(new_n3283_), .B(new_n3714_), .ZN(new_n4062_));
  NAND2_X1   g4013(.A1(new_n4062_), .A2(new_n4061_), .ZN(new_n4063_));
  INV_X1     g4014(.I(new_n3749_), .ZN(new_n4064_));
  NAND3_X1   g4015(.A1(new_n4063_), .A2(new_n3730_), .A3(new_n4064_), .ZN(new_n4065_));
  NAND3_X1   g4016(.A1(new_n4065_), .A2(new_n3697_), .A3(new_n3719_), .ZN(new_n4066_));
  AOI21_X1   g4017(.A1(new_n4066_), .A2(new_n3752_), .B(new_n3777_), .ZN(new_n4067_));
  NOR2_X1    g4018(.A1(new_n4060_), .A2(new_n4067_), .ZN(new_n4068_));
  XOR2_X1    g4019(.A1(new_n4068_), .A2(new_n4057_), .Z(new_n4069_));
  XOR2_X1    g4020(.A1(new_n4069_), .A2(new_n4055_), .Z(new_n4070_));
  XOR2_X1    g4021(.A1(new_n4070_), .A2(new_n3899_), .Z(new_n4071_));
  INV_X1     g4022(.I(new_n4071_), .ZN(\sin[0] ));
  XOR2_X1    g4023(.A1(\a[22] ), .A2(\a[23] ), .Z(new_n4073_));
  INV_X1     g4024(.I(new_n4073_), .ZN(new_n4074_));
  NOR2_X1    g4025(.A1(new_n4071_), .A2(new_n4074_), .ZN(new_n4075_));
  NAND3_X1   g4026(.A1(new_n4066_), .A2(new_n3752_), .A3(new_n4056_), .ZN(new_n4076_));
  XNOR2_X1   g4027(.A1(new_n3777_), .A2(new_n3896_), .ZN(new_n4077_));
  AOI21_X1   g4028(.A1(new_n4066_), .A2(new_n3752_), .B(new_n4056_), .ZN(new_n4078_));
  AOI21_X1   g4029(.A1(new_n4077_), .A2(new_n4076_), .B(new_n4078_), .ZN(new_n4079_));
  AOI21_X1   g4030(.A1(new_n4052_), .A2(new_n4054_), .B(new_n4079_), .ZN(new_n4080_));
  NOR2_X1    g4031(.A1(new_n4055_), .A2(new_n3899_), .ZN(new_n4081_));
  OAI21_X1   g4032(.A1(new_n4081_), .A2(new_n4080_), .B(new_n4069_), .ZN(new_n4082_));
  NOR2_X1    g4033(.A1(new_n3982_), .A2(new_n3983_), .ZN(new_n4083_));
  XOR2_X1    g4034(.A1(new_n4024_), .A2(new_n4083_), .Z(new_n4084_));
  XOR2_X1    g4035(.A1(new_n4015_), .A2(new_n52_), .Z(new_n4085_));
  NOR2_X1    g4036(.A1(new_n4084_), .A2(new_n4085_), .ZN(new_n4086_));
  AOI21_X1   g4037(.A1(new_n4035_), .A2(new_n4039_), .B(new_n4086_), .ZN(new_n4087_));
  AOI22_X1   g4038(.A1(new_n4001_), .A2(new_n2587_), .B1(new_n3868_), .B2(new_n55_), .ZN(new_n4088_));
  NOR4_X1    g4039(.A1(new_n193_), .A2(new_n210_), .A3(new_n388_), .A4(new_n443_), .ZN(new_n4089_));
  NAND4_X1   g4040(.A1(new_n4089_), .A2(new_n574_), .A3(new_n995_), .A4(new_n1017_), .ZN(new_n4090_));
  NOR4_X1    g4041(.A1(new_n387_), .A2(new_n191_), .A3(new_n444_), .A4(new_n687_), .ZN(new_n4091_));
  NOR2_X1    g4042(.A1(new_n2324_), .A2(new_n731_), .ZN(new_n4092_));
  NAND4_X1   g4043(.A1(new_n4092_), .A2(new_n418_), .A3(new_n2461_), .A4(new_n4091_), .ZN(new_n4093_));
  NOR4_X1    g4044(.A1(new_n4093_), .A2(new_n697_), .A3(new_n1436_), .A4(new_n4090_), .ZN(new_n4094_));
  NAND2_X1   g4045(.A1(new_n2473_), .A2(new_n4094_), .ZN(new_n4095_));
  NAND4_X1   g4046(.A1(new_n3572_), .A2(new_n3864_), .A3(new_n3999_), .A4(new_n4095_), .ZN(new_n4096_));
  NAND3_X1   g4047(.A1(new_n4000_), .A2(new_n2473_), .A3(new_n4094_), .ZN(new_n4097_));
  NAND2_X1   g4048(.A1(new_n4097_), .A2(new_n4096_), .ZN(new_n4098_));
  OAI21_X1   g4049(.A1(new_n2601_), .A2(new_n4098_), .B(new_n4088_), .ZN(new_n4099_));
  INV_X1     g4050(.I(new_n4099_), .ZN(new_n4100_));
  AOI21_X1   g4051(.A1(new_n3874_), .A2(new_n3868_), .B(new_n4001_), .ZN(new_n4101_));
  INV_X1     g4052(.I(new_n4101_), .ZN(new_n4102_));
  NAND2_X1   g4053(.A1(new_n3876_), .A2(new_n3869_), .ZN(new_n4103_));
  NAND2_X1   g4054(.A1(new_n4102_), .A2(new_n4103_), .ZN(new_n4104_));
  NAND3_X1   g4055(.A1(new_n4000_), .A2(new_n3998_), .A3(new_n4095_), .ZN(new_n4105_));
  NAND2_X1   g4056(.A1(new_n4098_), .A2(new_n4001_), .ZN(new_n4106_));
  NAND2_X1   g4057(.A1(new_n4106_), .A2(new_n4105_), .ZN(new_n4107_));
  NOR2_X1    g4058(.A1(new_n4104_), .A2(new_n4107_), .ZN(new_n4108_));
  AOI21_X1   g4059(.A1(new_n3869_), .A2(new_n3876_), .B(new_n4101_), .ZN(new_n4109_));
  AOI21_X1   g4060(.A1(new_n4105_), .A2(new_n4106_), .B(new_n4109_), .ZN(new_n4110_));
  OAI21_X1   g4061(.A1(new_n4110_), .A2(new_n4108_), .B(new_n2722_), .ZN(new_n4111_));
  AOI21_X1   g4062(.A1(new_n4111_), .A2(new_n4100_), .B(new_n2725_), .ZN(new_n4112_));
  NAND3_X1   g4063(.A1(new_n4109_), .A2(new_n4105_), .A3(new_n4106_), .ZN(new_n4113_));
  NAND2_X1   g4064(.A1(new_n4104_), .A2(new_n4107_), .ZN(new_n4114_));
  AOI21_X1   g4065(.A1(new_n4114_), .A2(new_n4113_), .B(new_n2729_), .ZN(new_n4115_));
  NOR3_X1    g4066(.A1(new_n4115_), .A2(new_n52_), .A3(new_n4099_), .ZN(new_n4116_));
  NOR2_X1    g4067(.A1(new_n4112_), .A2(new_n4116_), .ZN(new_n4117_));
  OAI22_X1   g4068(.A1(new_n2598_), .A2(new_n3051_), .B1(new_n2586_), .B2(new_n3057_), .ZN(new_n4118_));
  NOR2_X1    g4069(.A1(new_n3573_), .A2(new_n3061_), .ZN(new_n4119_));
  NOR2_X1    g4070(.A1(new_n4119_), .A2(new_n4118_), .ZN(new_n4120_));
  INV_X1     g4071(.I(new_n4120_), .ZN(new_n4121_));
  AOI21_X1   g4072(.A1(new_n3592_), .A2(new_n3593_), .B(new_n3074_), .ZN(new_n4122_));
  OAI21_X1   g4073(.A1(new_n4122_), .A2(new_n4121_), .B(new_n1288_), .ZN(new_n4123_));
  OAI21_X1   g4074(.A1(new_n3584_), .A2(new_n3588_), .B(new_n3073_), .ZN(new_n4124_));
  NAND3_X1   g4075(.A1(new_n4124_), .A2(new_n1287_), .A3(new_n4120_), .ZN(new_n4125_));
  NAND2_X1   g4076(.A1(new_n4123_), .A2(new_n4125_), .ZN(new_n4126_));
  NOR2_X1    g4077(.A1(new_n2563_), .A2(new_n2860_), .ZN(new_n4127_));
  NOR2_X1    g4078(.A1(new_n2694_), .A2(new_n2856_), .ZN(new_n4128_));
  NOR2_X1    g4079(.A1(new_n2611_), .A2(new_n2852_), .ZN(new_n4129_));
  NOR3_X1    g4080(.A1(new_n4127_), .A2(new_n4128_), .A3(new_n4129_), .ZN(new_n4130_));
  OAI21_X1   g4081(.A1(new_n3599_), .A2(new_n2880_), .B(new_n4130_), .ZN(new_n4131_));
  OAI22_X1   g4082(.A1(new_n2956_), .A2(new_n2739_), .B1(new_n2858_), .B2(new_n2768_), .ZN(new_n4132_));
  NOR2_X1    g4083(.A1(new_n2666_), .A2(new_n2736_), .ZN(new_n4133_));
  NOR2_X1    g4084(.A1(new_n4133_), .A2(new_n4132_), .ZN(new_n4134_));
  INV_X1     g4085(.I(new_n4134_), .ZN(new_n4135_));
  AOI21_X1   g4086(.A1(new_n3112_), .A2(new_n3111_), .B(new_n2743_), .ZN(new_n4136_));
  OAI21_X1   g4087(.A1(new_n4135_), .A2(new_n4136_), .B(new_n474_), .ZN(new_n4137_));
  NOR3_X1    g4088(.A1(new_n4135_), .A2(new_n4136_), .A3(new_n474_), .ZN(new_n4138_));
  INV_X1     g4089(.I(new_n4138_), .ZN(new_n4139_));
  NOR2_X1    g4090(.A1(new_n2645_), .A2(new_n598_), .ZN(new_n4140_));
  INV_X1     g4091(.I(new_n4140_), .ZN(new_n4141_));
  NAND4_X1   g4092(.A1(new_n3932_), .A2(new_n465_), .A3(new_n2754_), .A4(new_n3931_), .ZN(new_n4142_));
  INV_X1     g4093(.I(new_n4142_), .ZN(new_n4143_));
  OAI22_X1   g4094(.A1(new_n2845_), .A2(new_n2815_), .B1(new_n2792_), .B2(new_n3001_), .ZN(new_n4144_));
  AOI21_X1   g4095(.A1(new_n2881_), .A2(new_n2812_), .B(new_n4144_), .ZN(new_n4145_));
  OAI21_X1   g4096(.A1(new_n3147_), .A2(new_n3146_), .B(new_n2819_), .ZN(new_n4146_));
  NAND2_X1   g4097(.A1(new_n4146_), .A2(new_n4145_), .ZN(new_n4147_));
  INV_X1     g4098(.I(new_n4147_), .ZN(new_n4148_));
  OAI21_X1   g4099(.A1(new_n3943_), .A2(new_n4143_), .B(new_n4148_), .ZN(new_n4149_));
  AOI21_X1   g4100(.A1(new_n3630_), .A2(new_n3626_), .B(new_n598_), .ZN(new_n4150_));
  NOR3_X1    g4101(.A1(new_n3627_), .A2(new_n3628_), .A3(new_n465_), .ZN(new_n4151_));
  OAI21_X1   g4102(.A1(new_n4151_), .A2(new_n4150_), .B(new_n3624_), .ZN(new_n4152_));
  NOR3_X1    g4103(.A1(new_n4151_), .A2(new_n4150_), .A3(new_n3624_), .ZN(new_n4153_));
  AOI21_X1   g4104(.A1(new_n4152_), .A2(new_n3007_), .B(new_n4153_), .ZN(new_n4154_));
  OAI21_X1   g4105(.A1(new_n4154_), .A2(new_n3817_), .B(new_n3821_), .ZN(new_n4155_));
  OAI21_X1   g4106(.A1(new_n4154_), .A2(new_n3938_), .B(new_n3940_), .ZN(new_n4156_));
  NAND3_X1   g4107(.A1(new_n3945_), .A2(new_n4156_), .A3(new_n4155_), .ZN(new_n4157_));
  NAND3_X1   g4108(.A1(new_n4157_), .A2(new_n4142_), .A3(new_n4147_), .ZN(new_n4158_));
  NAND3_X1   g4109(.A1(new_n4149_), .A2(new_n4158_), .A3(new_n4141_), .ZN(new_n4159_));
  AOI21_X1   g4110(.A1(new_n4157_), .A2(new_n4142_), .B(new_n4147_), .ZN(new_n4160_));
  NOR3_X1    g4111(.A1(new_n3943_), .A2(new_n4143_), .A3(new_n4148_), .ZN(new_n4161_));
  OAI21_X1   g4112(.A1(new_n4161_), .A2(new_n4160_), .B(new_n4140_), .ZN(new_n4162_));
  NAND2_X1   g4113(.A1(new_n4162_), .A2(new_n4159_), .ZN(new_n4163_));
  NAND3_X1   g4114(.A1(new_n4139_), .A2(new_n4163_), .A3(new_n4137_), .ZN(new_n4164_));
  INV_X1     g4115(.I(new_n4137_), .ZN(new_n4165_));
  NOR3_X1    g4116(.A1(new_n4161_), .A2(new_n4160_), .A3(new_n4140_), .ZN(new_n4166_));
  AOI21_X1   g4117(.A1(new_n4149_), .A2(new_n4158_), .B(new_n4141_), .ZN(new_n4167_));
  NOR2_X1    g4118(.A1(new_n4166_), .A2(new_n4167_), .ZN(new_n4168_));
  OAI21_X1   g4119(.A1(new_n4165_), .A2(new_n4138_), .B(new_n4168_), .ZN(new_n4169_));
  NAND2_X1   g4120(.A1(new_n4169_), .A2(new_n4164_), .ZN(new_n4170_));
  AOI21_X1   g4121(.A1(new_n3950_), .A2(new_n3954_), .B(new_n3957_), .ZN(new_n4171_));
  NOR2_X1    g4122(.A1(new_n4170_), .A2(new_n4171_), .ZN(new_n4172_));
  NOR3_X1    g4123(.A1(new_n4168_), .A2(new_n4165_), .A3(new_n4138_), .ZN(new_n4173_));
  AOI21_X1   g4124(.A1(new_n4137_), .A2(new_n4139_), .B(new_n4163_), .ZN(new_n4174_));
  NOR2_X1    g4125(.A1(new_n4174_), .A2(new_n4173_), .ZN(new_n4175_));
  OAI21_X1   g4126(.A1(new_n3956_), .A2(new_n3958_), .B(new_n3953_), .ZN(new_n4176_));
  NOR2_X1    g4127(.A1(new_n4175_), .A2(new_n4176_), .ZN(new_n4177_));
  OAI21_X1   g4128(.A1(new_n4177_), .A2(new_n4172_), .B(new_n846_), .ZN(new_n4178_));
  NAND2_X1   g4129(.A1(new_n4175_), .A2(new_n4176_), .ZN(new_n4179_));
  NAND2_X1   g4130(.A1(new_n4170_), .A2(new_n4171_), .ZN(new_n4180_));
  NAND3_X1   g4131(.A1(new_n4179_), .A2(new_n4180_), .A3(new_n845_), .ZN(new_n4181_));
  NAND3_X1   g4132(.A1(new_n4178_), .A2(new_n4181_), .A3(new_n4131_), .ZN(new_n4182_));
  INV_X1     g4133(.I(new_n4130_), .ZN(new_n4183_));
  AOI21_X1   g4134(.A1(new_n3544_), .A2(new_n2863_), .B(new_n4183_), .ZN(new_n4184_));
  AOI21_X1   g4135(.A1(new_n4179_), .A2(new_n4180_), .B(new_n845_), .ZN(new_n4185_));
  NOR3_X1    g4136(.A1(new_n4177_), .A2(new_n4172_), .A3(new_n846_), .ZN(new_n4186_));
  OAI21_X1   g4137(.A1(new_n4185_), .A2(new_n4186_), .B(new_n4184_), .ZN(new_n4187_));
  OAI21_X1   g4138(.A1(new_n3967_), .A2(new_n3966_), .B(new_n3960_), .ZN(new_n4188_));
  NAND3_X1   g4139(.A1(new_n4188_), .A2(new_n4182_), .A3(new_n4187_), .ZN(new_n4189_));
  NAND2_X1   g4140(.A1(new_n4187_), .A2(new_n4182_), .ZN(new_n4190_));
  AOI21_X1   g4141(.A1(new_n3973_), .A2(new_n3971_), .B(new_n3969_), .ZN(new_n4191_));
  NAND2_X1   g4142(.A1(new_n4190_), .A2(new_n4191_), .ZN(new_n4192_));
  AOI21_X1   g4143(.A1(new_n4192_), .A2(new_n4189_), .B(new_n4126_), .ZN(new_n4193_));
  AOI21_X1   g4144(.A1(new_n4124_), .A2(new_n4120_), .B(new_n1287_), .ZN(new_n4194_));
  NOR3_X1    g4145(.A1(new_n4122_), .A2(new_n1288_), .A3(new_n4121_), .ZN(new_n4195_));
  NOR2_X1    g4146(.A1(new_n4194_), .A2(new_n4195_), .ZN(new_n4196_));
  NOR2_X1    g4147(.A1(new_n4190_), .A2(new_n4191_), .ZN(new_n4197_));
  AOI21_X1   g4148(.A1(new_n4182_), .A2(new_n4187_), .B(new_n4188_), .ZN(new_n4198_));
  NOR3_X1    g4149(.A1(new_n4198_), .A2(new_n4197_), .A3(new_n4196_), .ZN(new_n4199_));
  NOR2_X1    g4150(.A1(new_n4199_), .A2(new_n4193_), .ZN(new_n4200_));
  AOI21_X1   g4151(.A1(new_n3782_), .A2(new_n3856_), .B(new_n3791_), .ZN(new_n4201_));
  OAI21_X1   g4152(.A1(new_n4201_), .A2(new_n4017_), .B(new_n3980_), .ZN(new_n4202_));
  NAND3_X1   g4153(.A1(new_n4202_), .A2(new_n4200_), .A3(new_n3975_), .ZN(new_n4203_));
  OAI21_X1   g4154(.A1(new_n4198_), .A2(new_n4197_), .B(new_n4196_), .ZN(new_n4204_));
  NAND3_X1   g4155(.A1(new_n4192_), .A2(new_n4189_), .A3(new_n4126_), .ZN(new_n4205_));
  NAND2_X1   g4156(.A1(new_n4204_), .A2(new_n4205_), .ZN(new_n4206_));
  NAND2_X1   g4157(.A1(new_n4018_), .A2(new_n4016_), .ZN(new_n4207_));
  AOI21_X1   g4158(.A1(new_n4207_), .A2(new_n4022_), .B(new_n3983_), .ZN(new_n4208_));
  OAI21_X1   g4159(.A1(new_n4208_), .A2(new_n3982_), .B(new_n4206_), .ZN(new_n4209_));
  NAND3_X1   g4160(.A1(new_n4209_), .A2(new_n4203_), .A3(new_n4117_), .ZN(new_n4210_));
  INV_X1     g4161(.I(new_n4117_), .ZN(new_n4211_));
  NOR3_X1    g4162(.A1(new_n4208_), .A2(new_n4206_), .A3(new_n3982_), .ZN(new_n4212_));
  AOI21_X1   g4163(.A1(new_n4024_), .A2(new_n3980_), .B(new_n3982_), .ZN(new_n4213_));
  NOR2_X1    g4164(.A1(new_n4213_), .A2(new_n4200_), .ZN(new_n4214_));
  OAI21_X1   g4165(.A1(new_n4214_), .A2(new_n4212_), .B(new_n4211_), .ZN(new_n4215_));
  NOR3_X1    g4166(.A1(new_n2303_), .A2(new_n444_), .A3(new_n856_), .ZN(new_n4216_));
  NOR4_X1    g4167(.A1(new_n691_), .A2(new_n2272_), .A3(new_n435_), .A4(new_n357_), .ZN(new_n4217_));
  NOR4_X1    g4168(.A1(new_n179_), .A2(new_n723_), .A3(new_n332_), .A4(new_n378_), .ZN(new_n4218_));
  NAND4_X1   g4169(.A1(new_n2572_), .A2(new_n2567_), .A3(new_n4217_), .A4(new_n4218_), .ZN(new_n4219_));
  NOR3_X1    g4170(.A1(new_n4219_), .A2(new_n731_), .A3(new_n2380_), .ZN(new_n4220_));
  NAND4_X1   g4171(.A1(new_n4220_), .A2(new_n3767_), .A3(new_n2342_), .A4(new_n4216_), .ZN(new_n4221_));
  INV_X1     g4172(.I(new_n4221_), .ZN(new_n4222_));
  NAND3_X1   g4173(.A1(new_n4215_), .A2(new_n4210_), .A3(new_n4222_), .ZN(new_n4223_));
  NOR3_X1    g4174(.A1(new_n4214_), .A2(new_n4212_), .A3(new_n4211_), .ZN(new_n4224_));
  AOI21_X1   g4175(.A1(new_n4209_), .A2(new_n4203_), .B(new_n4117_), .ZN(new_n4225_));
  OAI21_X1   g4176(.A1(new_n4224_), .A2(new_n4225_), .B(new_n4221_), .ZN(new_n4226_));
  NAND2_X1   g4177(.A1(new_n4226_), .A2(new_n4223_), .ZN(new_n4227_));
  NOR2_X1    g4178(.A1(new_n4227_), .A2(new_n4087_), .ZN(new_n4228_));
  AOI21_X1   g4179(.A1(new_n3848_), .A2(new_n3858_), .B(new_n3888_), .ZN(new_n4229_));
  AOI21_X1   g4180(.A1(new_n4059_), .A2(new_n3889_), .B(new_n4229_), .ZN(new_n4230_));
  INV_X1     g4181(.I(new_n4086_), .ZN(new_n4231_));
  OAI21_X1   g4182(.A1(new_n4230_), .A2(new_n4033_), .B(new_n4231_), .ZN(new_n4232_));
  NOR3_X1    g4183(.A1(new_n4224_), .A2(new_n4225_), .A3(new_n4221_), .ZN(new_n4233_));
  AOI21_X1   g4184(.A1(new_n4215_), .A2(new_n4210_), .B(new_n4222_), .ZN(new_n4234_));
  NOR2_X1    g4185(.A1(new_n4233_), .A2(new_n4234_), .ZN(new_n4235_));
  NOR2_X1    g4186(.A1(new_n4235_), .A2(new_n4232_), .ZN(new_n4236_));
  NOR2_X1    g4187(.A1(new_n4236_), .A2(new_n4228_), .ZN(new_n4237_));
  OAI21_X1   g4188(.A1(new_n4036_), .A2(new_n4044_), .B(new_n4051_), .ZN(new_n4238_));
  NOR3_X1    g4189(.A1(new_n4036_), .A2(new_n4044_), .A3(new_n4051_), .ZN(new_n4239_));
  OAI21_X1   g4190(.A1(new_n3899_), .A2(new_n4239_), .B(new_n4238_), .ZN(new_n4240_));
  XOR2_X1    g4191(.A1(new_n4240_), .A2(new_n4237_), .Z(new_n4241_));
  NOR2_X1    g4192(.A1(new_n4241_), .A2(new_n4082_), .ZN(new_n4242_));
  INV_X1     g4193(.I(new_n4242_), .ZN(new_n4243_));
  NAND2_X1   g4194(.A1(new_n4241_), .A2(new_n4082_), .ZN(new_n4244_));
  NAND2_X1   g4195(.A1(new_n4243_), .A2(new_n4244_), .ZN(new_n4245_));
  XNOR2_X1   g4196(.A1(new_n4075_), .A2(new_n4245_), .ZN(\sin[1] ));
  NAND2_X1   g4197(.A1(new_n4071_), .A2(new_n4245_), .ZN(new_n4247_));
  NAND2_X1   g4198(.A1(new_n4247_), .A2(new_n4073_), .ZN(new_n4248_));
  NAND3_X1   g4199(.A1(new_n4043_), .A2(new_n4039_), .A3(new_n3895_), .ZN(new_n4249_));
  NAND2_X1   g4200(.A1(new_n4035_), .A2(new_n4033_), .ZN(new_n4250_));
  AOI21_X1   g4201(.A1(new_n4250_), .A2(new_n4249_), .B(new_n4053_), .ZN(new_n4251_));
  NAND3_X1   g4202(.A1(new_n4250_), .A2(new_n4249_), .A3(new_n4053_), .ZN(new_n4252_));
  AOI21_X1   g4203(.A1(new_n4079_), .A2(new_n4252_), .B(new_n4251_), .ZN(new_n4253_));
  NAND2_X1   g4204(.A1(new_n4215_), .A2(new_n4210_), .ZN(new_n4254_));
  INV_X1     g4205(.I(new_n4254_), .ZN(new_n4255_));
  NOR2_X1    g4206(.A1(new_n4087_), .A2(new_n4255_), .ZN(new_n4256_));
  AOI21_X1   g4207(.A1(new_n4043_), .A2(new_n3895_), .B(new_n4033_), .ZN(new_n4257_));
  NOR3_X1    g4208(.A1(new_n4257_), .A2(new_n4086_), .A3(new_n4254_), .ZN(new_n4258_));
  NOR2_X1    g4209(.A1(new_n4256_), .A2(new_n4258_), .ZN(new_n4259_));
  OAI22_X1   g4210(.A1(new_n4253_), .A2(new_n4237_), .B1(new_n4222_), .B2(new_n4259_), .ZN(new_n4260_));
  AOI21_X1   g4211(.A1(new_n4087_), .A2(new_n4210_), .B(new_n4225_), .ZN(new_n4261_));
  AOI22_X1   g4212(.A1(new_n3859_), .A2(new_n3141_), .B1(new_n3578_), .B2(new_n3056_), .ZN(new_n4262_));
  OAI21_X1   g4213(.A1(new_n3869_), .A2(new_n3061_), .B(new_n4262_), .ZN(new_n4263_));
  NOR2_X1    g4214(.A1(new_n3885_), .A2(new_n3074_), .ZN(new_n4264_));
  OAI21_X1   g4215(.A1(new_n4264_), .A2(new_n4263_), .B(new_n1288_), .ZN(new_n4265_));
  INV_X1     g4216(.I(new_n4263_), .ZN(new_n4266_));
  NAND2_X1   g4217(.A1(new_n3881_), .A2(new_n3073_), .ZN(new_n4267_));
  NAND3_X1   g4218(.A1(new_n4267_), .A2(new_n1287_), .A3(new_n4266_), .ZN(new_n4268_));
  AND2_X2    g4219(.A1(new_n4265_), .A2(new_n4268_), .Z(new_n4269_));
  OAI22_X1   g4220(.A1(new_n2563_), .A2(new_n2852_), .B1(new_n2611_), .B2(new_n2856_), .ZN(new_n4270_));
  NOR2_X1    g4221(.A1(new_n2586_), .A2(new_n2860_), .ZN(new_n4271_));
  NOR2_X1    g4222(.A1(new_n4271_), .A2(new_n4270_), .ZN(new_n4272_));
  NAND2_X1   g4223(.A1(new_n3269_), .A2(new_n3271_), .ZN(new_n4273_));
  NAND2_X1   g4224(.A1(new_n4273_), .A2(new_n2863_), .ZN(new_n4274_));
  AOI21_X1   g4225(.A1(new_n4274_), .A2(new_n4272_), .B(new_n846_), .ZN(new_n4275_));
  AND3_X2    g4226(.A1(new_n4274_), .A2(new_n846_), .A3(new_n4272_), .Z(new_n4276_));
  NOR2_X1    g4227(.A1(new_n4276_), .A2(new_n4275_), .ZN(new_n4277_));
  INV_X1     g4228(.I(new_n4277_), .ZN(new_n4278_));
  OAI22_X1   g4229(.A1(new_n2694_), .A2(new_n2736_), .B1(new_n2956_), .B2(new_n2768_), .ZN(new_n4279_));
  AOI21_X1   g4230(.A1(new_n2704_), .A2(new_n2738_), .B(new_n4279_), .ZN(new_n4280_));
  OAI21_X1   g4231(.A1(new_n3295_), .A2(new_n3290_), .B(new_n2748_), .ZN(new_n4281_));
  AOI21_X1   g4232(.A1(new_n4281_), .A2(new_n4280_), .B(new_n473_), .ZN(new_n4282_));
  NAND2_X1   g4233(.A1(new_n4281_), .A2(new_n4280_), .ZN(new_n4283_));
  NOR2_X1    g4234(.A1(new_n4283_), .A2(new_n474_), .ZN(new_n4284_));
  NOR2_X1    g4235(.A1(new_n4284_), .A2(new_n4282_), .ZN(new_n4285_));
  NOR2_X1    g4236(.A1(new_n2800_), .A2(new_n598_), .ZN(new_n4286_));
  INV_X1     g4237(.I(new_n4286_), .ZN(new_n4287_));
  OAI22_X1   g4238(.A1(new_n2697_), .A2(new_n2815_), .B1(new_n2845_), .B2(new_n3001_), .ZN(new_n4288_));
  AOI21_X1   g4239(.A1(new_n2671_), .A2(new_n2812_), .B(new_n4288_), .ZN(new_n4289_));
  NAND2_X1   g4240(.A1(new_n2872_), .A2(new_n2819_), .ZN(new_n4290_));
  NAND2_X1   g4241(.A1(new_n4290_), .A2(new_n4289_), .ZN(new_n4291_));
  INV_X1     g4242(.I(new_n4291_), .ZN(new_n4292_));
  NAND2_X1   g4243(.A1(new_n4149_), .A2(new_n4140_), .ZN(new_n4293_));
  AOI21_X1   g4244(.A1(new_n598_), .A2(new_n4148_), .B(new_n4161_), .ZN(new_n4294_));
  NAND2_X1   g4245(.A1(new_n4294_), .A2(new_n4293_), .ZN(new_n4295_));
  NAND2_X1   g4246(.A1(new_n4295_), .A2(new_n4292_), .ZN(new_n4296_));
  INV_X1     g4247(.I(new_n4296_), .ZN(new_n4297_));
  NOR2_X1    g4248(.A1(new_n4295_), .A2(new_n4292_), .ZN(new_n4298_));
  OAI21_X1   g4249(.A1(new_n4297_), .A2(new_n4298_), .B(new_n4287_), .ZN(new_n4299_));
  INV_X1     g4250(.I(new_n4298_), .ZN(new_n4300_));
  NOR2_X1    g4251(.A1(new_n4158_), .A2(new_n4291_), .ZN(new_n4301_));
  INV_X1     g4252(.I(new_n4301_), .ZN(new_n4302_));
  NAND4_X1   g4253(.A1(new_n4300_), .A2(new_n4286_), .A3(new_n4296_), .A4(new_n4302_), .ZN(new_n4303_));
  NAND2_X1   g4254(.A1(new_n4303_), .A2(new_n4299_), .ZN(new_n4304_));
  NAND2_X1   g4255(.A1(new_n4304_), .A2(new_n4285_), .ZN(new_n4305_));
  INV_X1     g4256(.I(new_n4305_), .ZN(new_n4306_));
  NOR2_X1    g4257(.A1(new_n4304_), .A2(new_n4285_), .ZN(new_n4307_));
  AOI21_X1   g4258(.A1(new_n4176_), .A2(new_n4164_), .B(new_n4174_), .ZN(new_n4308_));
  OAI21_X1   g4259(.A1(new_n4306_), .A2(new_n4307_), .B(new_n4308_), .ZN(new_n4309_));
  INV_X1     g4260(.I(new_n4307_), .ZN(new_n4310_));
  INV_X1     g4261(.I(new_n4308_), .ZN(new_n4311_));
  NAND3_X1   g4262(.A1(new_n4310_), .A2(new_n4305_), .A3(new_n4311_), .ZN(new_n4312_));
  NAND2_X1   g4263(.A1(new_n4309_), .A2(new_n4312_), .ZN(new_n4313_));
  XOR2_X1    g4264(.A1(new_n4184_), .A2(new_n846_), .Z(new_n4314_));
  NAND3_X1   g4265(.A1(new_n4314_), .A2(new_n4179_), .A3(new_n4180_), .ZN(new_n4315_));
  AOI21_X1   g4266(.A1(new_n4189_), .A2(new_n4315_), .B(new_n4313_), .ZN(new_n4316_));
  AOI21_X1   g4267(.A1(new_n4310_), .A2(new_n4305_), .B(new_n4311_), .ZN(new_n4317_));
  NOR3_X1    g4268(.A1(new_n4306_), .A2(new_n4307_), .A3(new_n4308_), .ZN(new_n4318_));
  NOR2_X1    g4269(.A1(new_n4317_), .A2(new_n4318_), .ZN(new_n4319_));
  INV_X1     g4270(.I(new_n4315_), .ZN(new_n4320_));
  NOR3_X1    g4271(.A1(new_n4320_), .A2(new_n4319_), .A3(new_n4197_), .ZN(new_n4321_));
  NOR3_X1    g4272(.A1(new_n4316_), .A2(new_n4321_), .A3(new_n4278_), .ZN(new_n4322_));
  OAI21_X1   g4273(.A1(new_n4320_), .A2(new_n4197_), .B(new_n4319_), .ZN(new_n4323_));
  NAND3_X1   g4274(.A1(new_n4313_), .A2(new_n4189_), .A3(new_n4315_), .ZN(new_n4324_));
  AOI21_X1   g4275(.A1(new_n4323_), .A2(new_n4324_), .B(new_n4277_), .ZN(new_n4325_));
  OAI21_X1   g4276(.A1(new_n4322_), .A2(new_n4325_), .B(new_n4269_), .ZN(new_n4326_));
  NAND2_X1   g4277(.A1(new_n4265_), .A2(new_n4268_), .ZN(new_n4327_));
  NAND3_X1   g4278(.A1(new_n4323_), .A2(new_n4277_), .A3(new_n4324_), .ZN(new_n4328_));
  OAI21_X1   g4279(.A1(new_n4316_), .A2(new_n4321_), .B(new_n4278_), .ZN(new_n4329_));
  NAND3_X1   g4280(.A1(new_n4329_), .A2(new_n4328_), .A3(new_n4327_), .ZN(new_n4330_));
  OAI21_X1   g4281(.A1(new_n4019_), .A2(new_n3983_), .B(new_n3975_), .ZN(new_n4331_));
  OAI21_X1   g4282(.A1(new_n4331_), .A2(new_n4206_), .B(new_n4205_), .ZN(new_n4332_));
  NAND3_X1   g4283(.A1(new_n4326_), .A2(new_n4332_), .A3(new_n4330_), .ZN(new_n4333_));
  AOI21_X1   g4284(.A1(new_n4329_), .A2(new_n4328_), .B(new_n4327_), .ZN(new_n4334_));
  NOR3_X1    g4285(.A1(new_n4269_), .A2(new_n4322_), .A3(new_n4325_), .ZN(new_n4335_));
  AOI21_X1   g4286(.A1(new_n4213_), .A2(new_n4204_), .B(new_n4199_), .ZN(new_n4336_));
  OAI21_X1   g4287(.A1(new_n4335_), .A2(new_n4334_), .B(new_n4336_), .ZN(new_n4337_));
  OAI22_X1   g4288(.A1(new_n4098_), .A2(new_n2588_), .B1(new_n4002_), .B2(new_n56_), .ZN(new_n4338_));
  NOR2_X1    g4289(.A1(new_n4104_), .A2(new_n4106_), .ZN(new_n4339_));
  NOR2_X1    g4290(.A1(new_n4109_), .A2(new_n4105_), .ZN(new_n4340_));
  NOR2_X1    g4291(.A1(new_n4339_), .A2(new_n4340_), .ZN(new_n4341_));
  NOR2_X1    g4292(.A1(new_n4341_), .A2(new_n2729_), .ZN(new_n4342_));
  NOR2_X1    g4293(.A1(new_n4342_), .A2(new_n4338_), .ZN(new_n4343_));
  XOR2_X1    g4294(.A1(new_n4343_), .A2(new_n2725_), .Z(new_n4344_));
  AOI21_X1   g4295(.A1(new_n4337_), .A2(new_n4333_), .B(new_n4344_), .ZN(new_n4345_));
  NOR3_X1    g4296(.A1(new_n4335_), .A2(new_n4336_), .A3(new_n4334_), .ZN(new_n4346_));
  AOI21_X1   g4297(.A1(new_n4326_), .A2(new_n4330_), .B(new_n4332_), .ZN(new_n4347_));
  INV_X1     g4298(.I(new_n4344_), .ZN(new_n4348_));
  NOR3_X1    g4299(.A1(new_n4347_), .A2(new_n4346_), .A3(new_n4348_), .ZN(new_n4349_));
  NOR2_X1    g4300(.A1(new_n4349_), .A2(new_n4345_), .ZN(new_n4350_));
  NOR2_X1    g4301(.A1(new_n4261_), .A2(new_n4350_), .ZN(new_n4351_));
  OAI21_X1   g4302(.A1(new_n4232_), .A2(new_n4224_), .B(new_n4215_), .ZN(new_n4352_));
  OAI21_X1   g4303(.A1(new_n4347_), .A2(new_n4346_), .B(new_n4348_), .ZN(new_n4353_));
  NAND3_X1   g4304(.A1(new_n4337_), .A2(new_n4333_), .A3(new_n4344_), .ZN(new_n4354_));
  NAND2_X1   g4305(.A1(new_n4353_), .A2(new_n4354_), .ZN(new_n4355_));
  NOR2_X1    g4306(.A1(new_n4352_), .A2(new_n4355_), .ZN(new_n4356_));
  NOR2_X1    g4307(.A1(new_n4356_), .A2(new_n4351_), .ZN(new_n4357_));
  NAND2_X1   g4308(.A1(new_n3729_), .A2(new_n683_), .ZN(new_n4358_));
  NOR2_X1    g4309(.A1(new_n718_), .A2(new_n1120_), .ZN(new_n4359_));
  NOR3_X1    g4310(.A1(new_n127_), .A2(new_n729_), .A3(new_n561_), .ZN(new_n4360_));
  NAND4_X1   g4311(.A1(new_n4359_), .A2(new_n3992_), .A3(new_n4360_), .A4(new_n578_), .ZN(new_n4361_));
  NOR4_X1    g4312(.A1(new_n549_), .A2(new_n193_), .A3(new_n285_), .A4(new_n310_), .ZN(new_n4362_));
  NOR3_X1    g4313(.A1(new_n426_), .A2(new_n536_), .A3(new_n745_), .ZN(new_n4363_));
  NAND4_X1   g4314(.A1(new_n4362_), .A2(new_n2413_), .A3(new_n507_), .A4(new_n4363_), .ZN(new_n4364_));
  NOR3_X1    g4315(.A1(new_n4358_), .A2(new_n4361_), .A3(new_n4364_), .ZN(new_n4365_));
  OAI21_X1   g4316(.A1(new_n4356_), .A2(new_n4351_), .B(new_n4365_), .ZN(new_n4366_));
  NAND2_X1   g4317(.A1(new_n4352_), .A2(new_n4355_), .ZN(new_n4367_));
  NAND2_X1   g4318(.A1(new_n4261_), .A2(new_n4350_), .ZN(new_n4368_));
  INV_X1     g4319(.I(new_n4365_), .ZN(new_n4369_));
  NAND3_X1   g4320(.A1(new_n4367_), .A2(new_n4368_), .A3(new_n4369_), .ZN(new_n4370_));
  NAND2_X1   g4321(.A1(new_n4366_), .A2(new_n4370_), .ZN(new_n4371_));
  AOI21_X1   g4322(.A1(new_n4357_), .A2(new_n4358_), .B(new_n4371_), .ZN(new_n4372_));
  NAND2_X1   g4323(.A1(new_n4372_), .A2(new_n4260_), .ZN(new_n4373_));
  NAND2_X1   g4324(.A1(new_n4235_), .A2(new_n4232_), .ZN(new_n4374_));
  NAND2_X1   g4325(.A1(new_n4227_), .A2(new_n4087_), .ZN(new_n4375_));
  NAND2_X1   g4326(.A1(new_n4374_), .A2(new_n4375_), .ZN(new_n4376_));
  OAI21_X1   g4327(.A1(new_n4257_), .A2(new_n4086_), .B(new_n4254_), .ZN(new_n4377_));
  NAND2_X1   g4328(.A1(new_n4087_), .A2(new_n4255_), .ZN(new_n4378_));
  AOI21_X1   g4329(.A1(new_n4378_), .A2(new_n4377_), .B(new_n4222_), .ZN(new_n4379_));
  AOI21_X1   g4330(.A1(new_n4240_), .A2(new_n4376_), .B(new_n4379_), .ZN(new_n4380_));
  NAND2_X1   g4331(.A1(new_n4371_), .A2(new_n4380_), .ZN(new_n4381_));
  NAND2_X1   g4332(.A1(new_n4373_), .A2(new_n4381_), .ZN(new_n4382_));
  NAND2_X1   g4333(.A1(new_n4382_), .A2(new_n4243_), .ZN(new_n4383_));
  NOR2_X1    g4334(.A1(new_n4382_), .A2(new_n4243_), .ZN(new_n4384_));
  INV_X1     g4335(.I(new_n4384_), .ZN(new_n4385_));
  NAND2_X1   g4336(.A1(new_n4385_), .A2(new_n4383_), .ZN(new_n4386_));
  XOR2_X1    g4337(.A1(new_n4386_), .A2(new_n4248_), .Z(\sin[2] ));
  NAND4_X1   g4338(.A1(new_n1000_), .A2(new_n408_), .A3(new_n740_), .A4(new_n912_), .ZN(new_n4388_));
  NOR4_X1    g4339(.A1(new_n323_), .A2(new_n2380_), .A3(new_n332_), .A4(new_n401_), .ZN(new_n4389_));
  NAND3_X1   g4340(.A1(new_n2338_), .A2(new_n897_), .A3(new_n4389_), .ZN(new_n4390_));
  NOR3_X1    g4341(.A1(new_n4390_), .A2(new_n720_), .A3(new_n4388_), .ZN(new_n4391_));
  NAND4_X1   g4342(.A1(new_n4391_), .A2(new_n1509_), .A3(new_n2249_), .A4(new_n3744_), .ZN(new_n4392_));
  INV_X1     g4343(.I(new_n4392_), .ZN(new_n4393_));
  AOI21_X1   g4344(.A1(new_n4261_), .A2(new_n4353_), .B(new_n4349_), .ZN(new_n4394_));
  NAND2_X1   g4345(.A1(new_n4333_), .A2(new_n4330_), .ZN(new_n4395_));
  NOR2_X1    g4346(.A1(new_n2563_), .A2(new_n2856_), .ZN(new_n4396_));
  NOR2_X1    g4347(.A1(new_n2586_), .A2(new_n2852_), .ZN(new_n4397_));
  NOR2_X1    g4348(.A1(new_n2598_), .A2(new_n2860_), .ZN(new_n4398_));
  NOR3_X1    g4349(.A1(new_n4398_), .A2(new_n4397_), .A3(new_n4396_), .ZN(new_n4399_));
  INV_X1     g4350(.I(new_n4399_), .ZN(new_n4400_));
  NOR2_X1    g4351(.A1(new_n3908_), .A2(new_n2880_), .ZN(new_n4401_));
  NOR2_X1    g4352(.A1(new_n4401_), .A2(new_n4400_), .ZN(new_n4402_));
  NOR2_X1    g4353(.A1(new_n4402_), .A2(new_n846_), .ZN(new_n4403_));
  NOR3_X1    g4354(.A1(new_n4401_), .A2(new_n845_), .A3(new_n4400_), .ZN(new_n4404_));
  NOR2_X1    g4355(.A1(new_n4403_), .A2(new_n4404_), .ZN(new_n4405_));
  INV_X1     g4356(.I(new_n4405_), .ZN(new_n4406_));
  AOI22_X1   g4357(.A1(new_n2613_), .A2(new_n2738_), .B1(new_n2704_), .B2(new_n2752_), .ZN(new_n4407_));
  OAI21_X1   g4358(.A1(new_n2611_), .A2(new_n2736_), .B(new_n4407_), .ZN(new_n4408_));
  NOR2_X1    g4359(.A1(new_n3473_), .A2(new_n2743_), .ZN(new_n4409_));
  OAI21_X1   g4360(.A1(new_n4409_), .A2(new_n4408_), .B(new_n474_), .ZN(new_n4410_));
  INV_X1     g4361(.I(new_n4410_), .ZN(new_n4411_));
  NOR3_X1    g4362(.A1(new_n4409_), .A2(new_n474_), .A3(new_n4408_), .ZN(new_n4412_));
  NOR2_X1    g4363(.A1(new_n4411_), .A2(new_n4412_), .ZN(new_n4413_));
  INV_X1     g4364(.I(new_n2976_), .ZN(new_n4414_));
  OAI22_X1   g4365(.A1(new_n2956_), .A2(new_n3003_), .B1(new_n2697_), .B2(new_n3001_), .ZN(new_n4415_));
  AOI21_X1   g4366(.A1(new_n2671_), .A2(new_n2816_), .B(new_n4415_), .ZN(new_n4416_));
  OAI21_X1   g4367(.A1(new_n4414_), .A2(new_n2820_), .B(new_n4416_), .ZN(new_n4417_));
  INV_X1     g4368(.I(new_n4417_), .ZN(new_n4418_));
  NOR2_X1    g4369(.A1(new_n4295_), .A2(new_n4291_), .ZN(new_n4419_));
  NOR2_X1    g4370(.A1(new_n4291_), .A2(new_n598_), .ZN(new_n4420_));
  OAI22_X1   g4371(.A1(new_n4287_), .A2(new_n4419_), .B1(new_n4298_), .B2(new_n4420_), .ZN(new_n4421_));
  NAND2_X1   g4372(.A1(new_n4421_), .A2(new_n4418_), .ZN(new_n4422_));
  NOR2_X1    g4373(.A1(new_n4419_), .A2(new_n4287_), .ZN(new_n4423_));
  NOR2_X1    g4374(.A1(new_n4298_), .A2(new_n4420_), .ZN(new_n4424_));
  NOR2_X1    g4375(.A1(new_n4423_), .A2(new_n4424_), .ZN(new_n4425_));
  NAND2_X1   g4376(.A1(new_n4425_), .A2(new_n4417_), .ZN(new_n4426_));
  NOR2_X1    g4377(.A1(new_n2630_), .A2(new_n598_), .ZN(new_n4427_));
  AOI21_X1   g4378(.A1(new_n4426_), .A2(new_n4422_), .B(new_n4427_), .ZN(new_n4428_));
  INV_X1     g4379(.I(new_n4422_), .ZN(new_n4429_));
  NOR2_X1    g4380(.A1(new_n4421_), .A2(new_n4418_), .ZN(new_n4430_));
  INV_X1     g4381(.I(new_n4427_), .ZN(new_n4431_));
  NOR3_X1    g4382(.A1(new_n4429_), .A2(new_n4430_), .A3(new_n4431_), .ZN(new_n4432_));
  NOR2_X1    g4383(.A1(new_n4432_), .A2(new_n4428_), .ZN(new_n4433_));
  OAI21_X1   g4384(.A1(new_n4318_), .A2(new_n4307_), .B(new_n4433_), .ZN(new_n4434_));
  OR2_X2     g4385(.A1(new_n4432_), .A2(new_n4428_), .Z(new_n4435_));
  AOI21_X1   g4386(.A1(new_n4305_), .A2(new_n4311_), .B(new_n4307_), .ZN(new_n4436_));
  NAND2_X1   g4387(.A1(new_n4435_), .A2(new_n4436_), .ZN(new_n4437_));
  NAND3_X1   g4388(.A1(new_n4437_), .A2(new_n4434_), .A3(new_n4413_), .ZN(new_n4438_));
  INV_X1     g4389(.I(new_n4413_), .ZN(new_n4439_));
  NOR2_X1    g4390(.A1(new_n4435_), .A2(new_n4436_), .ZN(new_n4440_));
  NOR3_X1    g4391(.A1(new_n4318_), .A2(new_n4307_), .A3(new_n4433_), .ZN(new_n4441_));
  OAI21_X1   g4392(.A1(new_n4440_), .A2(new_n4441_), .B(new_n4439_), .ZN(new_n4442_));
  NAND3_X1   g4393(.A1(new_n4442_), .A2(new_n4438_), .A3(new_n4406_), .ZN(new_n4443_));
  NOR3_X1    g4394(.A1(new_n4440_), .A2(new_n4441_), .A3(new_n4439_), .ZN(new_n4444_));
  AOI21_X1   g4395(.A1(new_n4437_), .A2(new_n4434_), .B(new_n4413_), .ZN(new_n4445_));
  OAI21_X1   g4396(.A1(new_n4445_), .A2(new_n4444_), .B(new_n4405_), .ZN(new_n4446_));
  NAND2_X1   g4397(.A1(new_n4446_), .A2(new_n4443_), .ZN(new_n4447_));
  NAND2_X1   g4398(.A1(new_n4323_), .A2(new_n4278_), .ZN(new_n4448_));
  OAI22_X1   g4399(.A1(new_n3869_), .A2(new_n3051_), .B1(new_n3057_), .B2(new_n3573_), .ZN(new_n4449_));
  NOR2_X1    g4400(.A1(new_n4002_), .A2(new_n3061_), .ZN(new_n4450_));
  NOR2_X1    g4401(.A1(new_n4449_), .A2(new_n4450_), .ZN(new_n4451_));
  INV_X1     g4402(.I(new_n4451_), .ZN(new_n4452_));
  AOI21_X1   g4403(.A1(new_n4013_), .A2(new_n4006_), .B(new_n3074_), .ZN(new_n4453_));
  OAI21_X1   g4404(.A1(new_n4453_), .A2(new_n4452_), .B(new_n1288_), .ZN(new_n4454_));
  INV_X1     g4405(.I(new_n4004_), .ZN(new_n4455_));
  AOI21_X1   g4406(.A1(new_n3874_), .A2(new_n3875_), .B(new_n4011_), .ZN(new_n4456_));
  OAI21_X1   g4407(.A1(new_n4456_), .A2(new_n4455_), .B(new_n3868_), .ZN(new_n4457_));
  NAND2_X1   g4408(.A1(new_n4008_), .A2(new_n4001_), .ZN(new_n4458_));
  NAND3_X1   g4409(.A1(new_n4457_), .A2(new_n4006_), .A3(new_n4458_), .ZN(new_n4459_));
  NAND2_X1   g4410(.A1(new_n4459_), .A2(new_n3073_), .ZN(new_n4460_));
  NAND3_X1   g4411(.A1(new_n4460_), .A2(new_n1287_), .A3(new_n4451_), .ZN(new_n4461_));
  NAND2_X1   g4412(.A1(new_n4461_), .A2(new_n4454_), .ZN(new_n4462_));
  NAND3_X1   g4413(.A1(new_n4448_), .A2(new_n4462_), .A3(new_n4324_), .ZN(new_n4463_));
  NOR2_X1    g4414(.A1(new_n4316_), .A2(new_n4277_), .ZN(new_n4464_));
  AOI21_X1   g4415(.A1(new_n4460_), .A2(new_n4451_), .B(new_n1287_), .ZN(new_n4465_));
  NOR3_X1    g4416(.A1(new_n4453_), .A2(new_n1288_), .A3(new_n4452_), .ZN(new_n4466_));
  NOR2_X1    g4417(.A1(new_n4465_), .A2(new_n4466_), .ZN(new_n4467_));
  OAI21_X1   g4418(.A1(new_n4464_), .A2(new_n4321_), .B(new_n4467_), .ZN(new_n4468_));
  AOI21_X1   g4419(.A1(new_n4463_), .A2(new_n4468_), .B(new_n4447_), .ZN(new_n4469_));
  NOR3_X1    g4420(.A1(new_n4445_), .A2(new_n4444_), .A3(new_n4405_), .ZN(new_n4470_));
  AOI21_X1   g4421(.A1(new_n4442_), .A2(new_n4438_), .B(new_n4406_), .ZN(new_n4471_));
  NOR2_X1    g4422(.A1(new_n4470_), .A2(new_n4471_), .ZN(new_n4472_));
  NOR3_X1    g4423(.A1(new_n4464_), .A2(new_n4467_), .A3(new_n4321_), .ZN(new_n4473_));
  AOI21_X1   g4424(.A1(new_n4448_), .A2(new_n4324_), .B(new_n4462_), .ZN(new_n4474_));
  NOR3_X1    g4425(.A1(new_n4472_), .A2(new_n4473_), .A3(new_n4474_), .ZN(new_n4475_));
  INV_X1     g4426(.I(new_n4098_), .ZN(new_n4476_));
  NAND2_X1   g4427(.A1(new_n4102_), .A2(new_n4476_), .ZN(new_n4477_));
  OAI22_X1   g4428(.A1(new_n4477_), .A2(new_n2729_), .B1(new_n56_), .B2(new_n4098_), .ZN(new_n4478_));
  XOR2_X1    g4429(.A1(new_n4478_), .A2(new_n52_), .Z(new_n4479_));
  INV_X1     g4430(.I(new_n4479_), .ZN(new_n4480_));
  NOR3_X1    g4431(.A1(new_n4469_), .A2(new_n4475_), .A3(new_n4480_), .ZN(new_n4481_));
  OAI21_X1   g4432(.A1(new_n4473_), .A2(new_n4474_), .B(new_n4472_), .ZN(new_n4482_));
  NAND3_X1   g4433(.A1(new_n4447_), .A2(new_n4468_), .A3(new_n4463_), .ZN(new_n4483_));
  AOI21_X1   g4434(.A1(new_n4482_), .A2(new_n4483_), .B(new_n4479_), .ZN(new_n4484_));
  OAI21_X1   g4435(.A1(new_n4484_), .A2(new_n4481_), .B(new_n4395_), .ZN(new_n4485_));
  NOR2_X1    g4436(.A1(new_n4346_), .A2(new_n4335_), .ZN(new_n4486_));
  NAND3_X1   g4437(.A1(new_n4482_), .A2(new_n4483_), .A3(new_n4479_), .ZN(new_n4487_));
  OAI21_X1   g4438(.A1(new_n4469_), .A2(new_n4475_), .B(new_n4480_), .ZN(new_n4488_));
  NAND3_X1   g4439(.A1(new_n4486_), .A2(new_n4488_), .A3(new_n4487_), .ZN(new_n4489_));
  NAND2_X1   g4440(.A1(new_n4489_), .A2(new_n4485_), .ZN(new_n4490_));
  NOR2_X1    g4441(.A1(new_n4394_), .A2(new_n4490_), .ZN(new_n4491_));
  OAI21_X1   g4442(.A1(new_n4352_), .A2(new_n4345_), .B(new_n4354_), .ZN(new_n4492_));
  AOI21_X1   g4443(.A1(new_n4487_), .A2(new_n4488_), .B(new_n4486_), .ZN(new_n4493_));
  NOR3_X1    g4444(.A1(new_n4481_), .A2(new_n4484_), .A3(new_n4395_), .ZN(new_n4494_));
  NOR2_X1    g4445(.A1(new_n4493_), .A2(new_n4494_), .ZN(new_n4495_));
  NOR2_X1    g4446(.A1(new_n4492_), .A2(new_n4495_), .ZN(new_n4496_));
  OAI21_X1   g4447(.A1(new_n4496_), .A2(new_n4491_), .B(new_n4393_), .ZN(new_n4497_));
  NOR3_X1    g4448(.A1(new_n4257_), .A2(new_n4086_), .A3(new_n4224_), .ZN(new_n4498_));
  NOR3_X1    g4449(.A1(new_n4498_), .A2(new_n4225_), .A3(new_n4345_), .ZN(new_n4499_));
  OAI21_X1   g4450(.A1(new_n4499_), .A2(new_n4349_), .B(new_n4495_), .ZN(new_n4500_));
  NAND2_X1   g4451(.A1(new_n4394_), .A2(new_n4490_), .ZN(new_n4501_));
  NAND3_X1   g4452(.A1(new_n4501_), .A2(new_n4500_), .A3(new_n4392_), .ZN(new_n4502_));
  NAND2_X1   g4453(.A1(new_n4497_), .A2(new_n4502_), .ZN(new_n4503_));
  NOR3_X1    g4454(.A1(new_n4356_), .A2(new_n4351_), .A3(new_n4365_), .ZN(new_n4504_));
  OAI21_X1   g4455(.A1(new_n4260_), .A2(new_n4504_), .B(new_n4366_), .ZN(new_n4505_));
  NOR2_X1    g4456(.A1(new_n4503_), .A2(new_n4505_), .ZN(new_n4506_));
  AOI21_X1   g4457(.A1(new_n4367_), .A2(new_n4368_), .B(new_n4369_), .ZN(new_n4507_));
  AOI21_X1   g4458(.A1(new_n4380_), .A2(new_n4370_), .B(new_n4507_), .ZN(new_n4508_));
  AOI21_X1   g4459(.A1(new_n4497_), .A2(new_n4502_), .B(new_n4508_), .ZN(new_n4509_));
  NOR2_X1    g4460(.A1(new_n4506_), .A2(new_n4509_), .ZN(new_n4510_));
  XNOR2_X1   g4461(.A1(new_n4510_), .A2(new_n4385_), .ZN(new_n4511_));
  INV_X1     g4462(.I(new_n4386_), .ZN(new_n4512_));
  OAI21_X1   g4463(.A1(new_n4512_), .A2(new_n4247_), .B(new_n4073_), .ZN(new_n4513_));
  XNOR2_X1   g4464(.A1(new_n4513_), .A2(new_n4511_), .ZN(\sin[3] ));
  NOR3_X1    g4465(.A1(new_n4511_), .A2(new_n4512_), .A3(new_n4247_), .ZN(new_n4515_));
  NOR2_X1    g4466(.A1(new_n4515_), .A2(new_n4074_), .ZN(new_n4516_));
  NAND2_X1   g4467(.A1(new_n4384_), .A2(new_n4510_), .ZN(new_n4517_));
  AOI21_X1   g4468(.A1(new_n4492_), .A2(new_n4495_), .B(new_n4493_), .ZN(new_n4518_));
  NOR2_X1    g4469(.A1(new_n4462_), .A2(new_n4479_), .ZN(new_n4519_));
  NAND2_X1   g4470(.A1(new_n4448_), .A2(new_n4324_), .ZN(new_n4520_));
  NAND2_X1   g4471(.A1(new_n4447_), .A2(new_n4520_), .ZN(new_n4521_));
  NOR2_X1    g4472(.A1(new_n4464_), .A2(new_n4321_), .ZN(new_n4522_));
  NAND2_X1   g4473(.A1(new_n4472_), .A2(new_n4522_), .ZN(new_n4523_));
  NOR2_X1    g4474(.A1(new_n4480_), .A2(new_n4467_), .ZN(new_n4524_));
  AOI21_X1   g4475(.A1(new_n4523_), .A2(new_n4521_), .B(new_n4524_), .ZN(new_n4525_));
  AOI21_X1   g4476(.A1(new_n4520_), .A2(new_n4446_), .B(new_n4470_), .ZN(new_n4526_));
  AOI22_X1   g4477(.A1(new_n4001_), .A2(new_n3141_), .B1(new_n3868_), .B2(new_n3056_), .ZN(new_n4527_));
  OAI21_X1   g4478(.A1(new_n3061_), .A2(new_n4098_), .B(new_n4527_), .ZN(new_n4528_));
  INV_X1     g4479(.I(new_n4528_), .ZN(new_n4529_));
  OAI21_X1   g4480(.A1(new_n4110_), .A2(new_n4108_), .B(new_n3073_), .ZN(new_n4530_));
  AOI21_X1   g4481(.A1(new_n4530_), .A2(new_n4529_), .B(new_n1287_), .ZN(new_n4531_));
  AOI21_X1   g4482(.A1(new_n4114_), .A2(new_n4113_), .B(new_n3074_), .ZN(new_n4532_));
  NOR3_X1    g4483(.A1(new_n4532_), .A2(new_n1288_), .A3(new_n4528_), .ZN(new_n4533_));
  NOR2_X1    g4484(.A1(new_n4531_), .A2(new_n4533_), .ZN(new_n4534_));
  INV_X1     g4485(.I(new_n4534_), .ZN(new_n4535_));
  OAI21_X1   g4486(.A1(new_n4439_), .A2(new_n4440_), .B(new_n4437_), .ZN(new_n4536_));
  OAI22_X1   g4487(.A1(new_n2563_), .A2(new_n2736_), .B1(new_n2694_), .B2(new_n2768_), .ZN(new_n4537_));
  AOI21_X1   g4488(.A1(new_n2716_), .A2(new_n2738_), .B(new_n4537_), .ZN(new_n4538_));
  NAND2_X1   g4489(.A1(new_n3544_), .A2(new_n2748_), .ZN(new_n4539_));
  AOI21_X1   g4490(.A1(new_n4539_), .A2(new_n4538_), .B(new_n473_), .ZN(new_n4540_));
  NAND2_X1   g4491(.A1(new_n4539_), .A2(new_n4538_), .ZN(new_n4541_));
  NOR2_X1    g4492(.A1(new_n4541_), .A2(new_n474_), .ZN(new_n4542_));
  NOR2_X1    g4493(.A1(new_n4542_), .A2(new_n4540_), .ZN(new_n4543_));
  NOR2_X1    g4494(.A1(new_n2697_), .A2(new_n598_), .ZN(new_n4544_));
  AOI22_X1   g4495(.A1(new_n2670_), .A2(new_n2816_), .B1(new_n2671_), .B2(new_n3000_), .ZN(new_n4545_));
  OAI21_X1   g4496(.A1(new_n2666_), .A2(new_n3003_), .B(new_n4545_), .ZN(new_n4546_));
  NOR2_X1    g4497(.A1(new_n3455_), .A2(new_n2820_), .ZN(new_n4547_));
  OAI21_X1   g4498(.A1(new_n4547_), .A2(new_n4546_), .B(new_n465_), .ZN(new_n4548_));
  OR3_X2     g4499(.A1(new_n4547_), .A2(new_n465_), .A3(new_n4546_), .Z(new_n4549_));
  NAND2_X1   g4500(.A1(new_n4549_), .A2(new_n4548_), .ZN(new_n4550_));
  NOR2_X1    g4501(.A1(new_n4550_), .A2(new_n52_), .ZN(new_n4551_));
  NAND2_X1   g4502(.A1(new_n4550_), .A2(new_n52_), .ZN(new_n4552_));
  INV_X1     g4503(.I(new_n4552_), .ZN(new_n4553_));
  NOR3_X1    g4504(.A1(new_n4553_), .A2(new_n4544_), .A3(new_n4551_), .ZN(new_n4554_));
  INV_X1     g4505(.I(new_n4544_), .ZN(new_n4555_));
  INV_X1     g4506(.I(new_n4551_), .ZN(new_n4556_));
  AOI21_X1   g4507(.A1(new_n4556_), .A2(new_n4552_), .B(new_n4555_), .ZN(new_n4557_));
  OAI21_X1   g4508(.A1(new_n4421_), .A2(new_n4417_), .B(new_n4427_), .ZN(new_n4558_));
  INV_X1     g4509(.I(new_n4558_), .ZN(new_n4559_));
  NOR2_X1    g4510(.A1(new_n4417_), .A2(new_n598_), .ZN(new_n4560_));
  INV_X1     g4511(.I(new_n4560_), .ZN(new_n4561_));
  OAI21_X1   g4512(.A1(new_n4421_), .A2(new_n4418_), .B(new_n4561_), .ZN(new_n4562_));
  INV_X1     g4513(.I(new_n4562_), .ZN(new_n4563_));
  OAI22_X1   g4514(.A1(new_n4559_), .A2(new_n4563_), .B1(new_n4557_), .B2(new_n4554_), .ZN(new_n4564_));
  NAND3_X1   g4515(.A1(new_n4556_), .A2(new_n4555_), .A3(new_n4552_), .ZN(new_n4565_));
  OAI21_X1   g4516(.A1(new_n4553_), .A2(new_n4551_), .B(new_n4544_), .ZN(new_n4566_));
  NAND4_X1   g4517(.A1(new_n4566_), .A2(new_n4565_), .A3(new_n4558_), .A4(new_n4562_), .ZN(new_n4567_));
  NAND2_X1   g4518(.A1(new_n4564_), .A2(new_n4567_), .ZN(new_n4568_));
  NOR2_X1    g4519(.A1(new_n4568_), .A2(new_n4543_), .ZN(new_n4569_));
  INV_X1     g4520(.I(new_n4543_), .ZN(new_n4570_));
  AOI22_X1   g4521(.A1(new_n4566_), .A2(new_n4565_), .B1(new_n4558_), .B2(new_n4562_), .ZN(new_n4571_));
  INV_X1     g4522(.I(new_n4567_), .ZN(new_n4572_));
  NOR2_X1    g4523(.A1(new_n4572_), .A2(new_n4571_), .ZN(new_n4573_));
  NOR2_X1    g4524(.A1(new_n4573_), .A2(new_n4570_), .ZN(new_n4574_));
  OAI22_X1   g4525(.A1(new_n2598_), .A2(new_n2852_), .B1(new_n2586_), .B2(new_n2856_), .ZN(new_n4575_));
  AOI21_X1   g4526(.A1(new_n2859_), .A2(new_n3859_), .B(new_n4575_), .ZN(new_n4576_));
  OAI21_X1   g4527(.A1(new_n3584_), .A2(new_n3588_), .B(new_n2863_), .ZN(new_n4577_));
  NAND2_X1   g4528(.A1(new_n4577_), .A2(new_n4576_), .ZN(new_n4578_));
  NAND2_X1   g4529(.A1(new_n4578_), .A2(new_n845_), .ZN(new_n4579_));
  NAND3_X1   g4530(.A1(new_n4577_), .A2(new_n846_), .A3(new_n4576_), .ZN(new_n4580_));
  NAND2_X1   g4531(.A1(new_n4579_), .A2(new_n4580_), .ZN(new_n4581_));
  OAI21_X1   g4532(.A1(new_n4574_), .A2(new_n4569_), .B(new_n4581_), .ZN(new_n4582_));
  NAND2_X1   g4533(.A1(new_n4573_), .A2(new_n4570_), .ZN(new_n4583_));
  NAND2_X1   g4534(.A1(new_n4568_), .A2(new_n4543_), .ZN(new_n4584_));
  NAND4_X1   g4535(.A1(new_n4583_), .A2(new_n4584_), .A3(new_n4579_), .A4(new_n4580_), .ZN(new_n4585_));
  NAND3_X1   g4536(.A1(new_n4585_), .A2(new_n4582_), .A3(new_n4536_), .ZN(new_n4586_));
  INV_X1     g4537(.I(new_n4586_), .ZN(new_n4587_));
  AOI21_X1   g4538(.A1(new_n4585_), .A2(new_n4582_), .B(new_n4536_), .ZN(new_n4588_));
  OAI21_X1   g4539(.A1(new_n4587_), .A2(new_n4588_), .B(new_n4535_), .ZN(new_n4589_));
  AOI21_X1   g4540(.A1(new_n4413_), .A2(new_n4434_), .B(new_n4441_), .ZN(new_n4590_));
  INV_X1     g4541(.I(new_n4582_), .ZN(new_n4591_));
  NOR3_X1    g4542(.A1(new_n4574_), .A2(new_n4581_), .A3(new_n4569_), .ZN(new_n4592_));
  OAI21_X1   g4543(.A1(new_n4591_), .A2(new_n4592_), .B(new_n4590_), .ZN(new_n4593_));
  NAND3_X1   g4544(.A1(new_n4593_), .A2(new_n4534_), .A3(new_n4586_), .ZN(new_n4594_));
  NAND2_X1   g4545(.A1(new_n4589_), .A2(new_n4594_), .ZN(new_n4595_));
  NOR2_X1    g4546(.A1(new_n4595_), .A2(new_n4526_), .ZN(new_n4596_));
  INV_X1     g4547(.I(new_n4526_), .ZN(new_n4597_));
  AOI21_X1   g4548(.A1(new_n4593_), .A2(new_n4586_), .B(new_n4534_), .ZN(new_n4598_));
  NOR3_X1    g4549(.A1(new_n4587_), .A2(new_n4535_), .A3(new_n4588_), .ZN(new_n4599_));
  NOR2_X1    g4550(.A1(new_n4599_), .A2(new_n4598_), .ZN(new_n4600_));
  NOR2_X1    g4551(.A1(new_n4600_), .A2(new_n4597_), .ZN(new_n4601_));
  NOR4_X1    g4552(.A1(new_n4601_), .A2(new_n4596_), .A3(new_n4525_), .A4(new_n4519_), .ZN(new_n4602_));
  NOR2_X1    g4553(.A1(new_n4525_), .A2(new_n4519_), .ZN(new_n4603_));
  NAND2_X1   g4554(.A1(new_n4600_), .A2(new_n4597_), .ZN(new_n4604_));
  NAND2_X1   g4555(.A1(new_n4595_), .A2(new_n4526_), .ZN(new_n4605_));
  AOI21_X1   g4556(.A1(new_n4604_), .A2(new_n4605_), .B(new_n4603_), .ZN(new_n4606_));
  NOR2_X1    g4557(.A1(new_n2356_), .A2(new_n159_), .ZN(new_n4607_));
  NOR4_X1    g4558(.A1(new_n2467_), .A2(new_n231_), .A3(new_n1069_), .A4(new_n446_), .ZN(new_n4608_));
  NAND4_X1   g4559(.A1(new_n4608_), .A2(new_n551_), .A3(new_n4359_), .A4(new_n4607_), .ZN(new_n4609_));
  NOR4_X1    g4560(.A1(new_n2441_), .A2(new_n4609_), .A3(new_n803_), .A4(new_n853_), .ZN(new_n4610_));
  OAI21_X1   g4561(.A1(new_n4606_), .A2(new_n4602_), .B(new_n4610_), .ZN(new_n4611_));
  NAND3_X1   g4562(.A1(new_n4603_), .A2(new_n4604_), .A3(new_n4605_), .ZN(new_n4612_));
  OAI22_X1   g4563(.A1(new_n4601_), .A2(new_n4596_), .B1(new_n4525_), .B2(new_n4519_), .ZN(new_n4613_));
  INV_X1     g4564(.I(new_n4610_), .ZN(new_n4614_));
  NAND3_X1   g4565(.A1(new_n4613_), .A2(new_n4612_), .A3(new_n4614_), .ZN(new_n4615_));
  NAND3_X1   g4566(.A1(new_n4613_), .A2(new_n4612_), .A3(new_n1257_), .ZN(new_n4616_));
  NAND3_X1   g4567(.A1(new_n4611_), .A2(new_n4615_), .A3(new_n4616_), .ZN(new_n4617_));
  NOR2_X1    g4568(.A1(new_n4617_), .A2(new_n4518_), .ZN(new_n4618_));
  OAI21_X1   g4569(.A1(new_n4394_), .A2(new_n4490_), .B(new_n4485_), .ZN(new_n4619_));
  AOI21_X1   g4570(.A1(new_n4613_), .A2(new_n4612_), .B(new_n4614_), .ZN(new_n4620_));
  NOR3_X1    g4571(.A1(new_n4606_), .A2(new_n4602_), .A3(new_n4610_), .ZN(new_n4621_));
  NOR2_X1    g4572(.A1(new_n4621_), .A2(new_n4620_), .ZN(new_n4622_));
  NOR2_X1    g4573(.A1(new_n4622_), .A2(new_n4619_), .ZN(new_n4623_));
  NOR2_X1    g4574(.A1(new_n4618_), .A2(new_n4623_), .ZN(new_n4624_));
  NOR3_X1    g4575(.A1(new_n4496_), .A2(new_n4491_), .A3(new_n4393_), .ZN(new_n4625_));
  AOI21_X1   g4576(.A1(new_n4508_), .A2(new_n4497_), .B(new_n4625_), .ZN(new_n4626_));
  XNOR2_X1   g4577(.A1(new_n4626_), .A2(new_n4624_), .ZN(new_n4627_));
  NOR2_X1    g4578(.A1(new_n4517_), .A2(new_n4627_), .ZN(new_n4628_));
  INV_X1     g4579(.I(new_n4628_), .ZN(new_n4629_));
  NAND2_X1   g4580(.A1(new_n4517_), .A2(new_n4627_), .ZN(new_n4630_));
  NAND2_X1   g4581(.A1(new_n4629_), .A2(new_n4630_), .ZN(new_n4631_));
  INV_X1     g4582(.I(new_n4631_), .ZN(new_n4632_));
  XOR2_X1    g4583(.A1(new_n4516_), .A2(new_n4632_), .Z(\sin[4] ));
  NAND2_X1   g4584(.A1(new_n4515_), .A2(new_n4631_), .ZN(new_n4634_));
  NAND2_X1   g4585(.A1(new_n4634_), .A2(new_n4073_), .ZN(new_n4635_));
  INV_X1     g4586(.I(new_n4603_), .ZN(new_n4636_));
  NOR2_X1    g4587(.A1(new_n4601_), .A2(new_n4596_), .ZN(new_n4637_));
  OAI21_X1   g4588(.A1(new_n4518_), .A2(new_n4637_), .B(new_n4636_), .ZN(new_n4638_));
  NAND3_X1   g4589(.A1(new_n4500_), .A2(new_n4485_), .A3(new_n4637_), .ZN(new_n4639_));
  NAND2_X1   g4590(.A1(new_n4638_), .A2(new_n4639_), .ZN(new_n4640_));
  AOI21_X1   g4591(.A1(new_n4597_), .A2(new_n4589_), .B(new_n4599_), .ZN(new_n4641_));
  AOI22_X1   g4592(.A1(new_n4476_), .A2(new_n3141_), .B1(new_n3056_), .B2(new_n4001_), .ZN(new_n4642_));
  OAI21_X1   g4593(.A1(new_n4341_), .A2(new_n3074_), .B(new_n4642_), .ZN(new_n4643_));
  XOR2_X1    g4594(.A1(new_n4643_), .A2(new_n1288_), .Z(new_n4644_));
  AOI21_X1   g4595(.A1(new_n4536_), .A2(new_n4585_), .B(new_n4591_), .ZN(new_n4645_));
  OAI22_X1   g4596(.A1(new_n3573_), .A2(new_n2852_), .B1(new_n2598_), .B2(new_n2856_), .ZN(new_n4646_));
  AOI21_X1   g4597(.A1(new_n3868_), .A2(new_n2859_), .B(new_n4646_), .ZN(new_n4647_));
  OAI21_X1   g4598(.A1(new_n3885_), .A2(new_n2880_), .B(new_n4647_), .ZN(new_n4648_));
  XOR2_X1    g4599(.A1(new_n4648_), .A2(new_n846_), .Z(new_n4649_));
  AOI21_X1   g4600(.A1(new_n4543_), .A2(new_n4567_), .B(new_n4571_), .ZN(new_n4650_));
  INV_X1     g4601(.I(new_n4650_), .ZN(new_n4651_));
  NAND2_X1   g4602(.A1(new_n4544_), .A2(new_n52_), .ZN(new_n4652_));
  NOR2_X1    g4603(.A1(new_n4544_), .A2(new_n52_), .ZN(new_n4653_));
  OAI21_X1   g4604(.A1(new_n4550_), .A2(new_n4653_), .B(new_n4652_), .ZN(new_n4654_));
  NOR2_X1    g4605(.A1(new_n2858_), .A2(new_n598_), .ZN(new_n4655_));
  INV_X1     g4606(.I(new_n4655_), .ZN(new_n4656_));
  NAND2_X1   g4607(.A1(new_n4656_), .A2(new_n2725_), .ZN(new_n4657_));
  NOR2_X1    g4608(.A1(new_n4656_), .A2(new_n2725_), .ZN(new_n4658_));
  INV_X1     g4609(.I(new_n4658_), .ZN(new_n4659_));
  NAND2_X1   g4610(.A1(new_n4659_), .A2(new_n4657_), .ZN(new_n4660_));
  XNOR2_X1   g4611(.A1(new_n4654_), .A2(new_n4660_), .ZN(new_n4661_));
  OAI22_X1   g4612(.A1(new_n2563_), .A2(new_n2739_), .B1(new_n2611_), .B2(new_n2768_), .ZN(new_n4662_));
  AOI21_X1   g4613(.A1(new_n2604_), .A2(new_n2735_), .B(new_n4662_), .ZN(new_n4663_));
  NAND2_X1   g4614(.A1(new_n4273_), .A2(new_n2748_), .ZN(new_n4664_));
  NAND2_X1   g4615(.A1(new_n4664_), .A2(new_n4663_), .ZN(new_n4665_));
  XOR2_X1    g4616(.A1(new_n4665_), .A2(new_n473_), .Z(new_n4666_));
  OAI22_X1   g4617(.A1(new_n2694_), .A2(new_n3003_), .B1(new_n2956_), .B2(new_n3001_), .ZN(new_n4667_));
  AOI21_X1   g4618(.A1(new_n2704_), .A2(new_n2816_), .B(new_n4667_), .ZN(new_n4668_));
  OAI21_X1   g4619(.A1(new_n3295_), .A2(new_n3290_), .B(new_n2819_), .ZN(new_n4669_));
  NAND2_X1   g4620(.A1(new_n4669_), .A2(new_n4668_), .ZN(new_n4670_));
  XOR2_X1    g4621(.A1(new_n4670_), .A2(new_n598_), .Z(new_n4671_));
  NOR2_X1    g4622(.A1(new_n4666_), .A2(new_n4671_), .ZN(new_n4672_));
  XOR2_X1    g4623(.A1(new_n4665_), .A2(new_n474_), .Z(new_n4673_));
  INV_X1     g4624(.I(new_n4671_), .ZN(new_n4674_));
  NOR2_X1    g4625(.A1(new_n4673_), .A2(new_n4674_), .ZN(new_n4675_));
  OAI21_X1   g4626(.A1(new_n4672_), .A2(new_n4675_), .B(new_n4661_), .ZN(new_n4676_));
  OR3_X2     g4627(.A1(new_n4672_), .A2(new_n4675_), .A3(new_n4661_), .Z(new_n4677_));
  AOI21_X1   g4628(.A1(new_n4677_), .A2(new_n4676_), .B(new_n4651_), .ZN(new_n4678_));
  INV_X1     g4629(.I(new_n4678_), .ZN(new_n4679_));
  NAND3_X1   g4630(.A1(new_n4677_), .A2(new_n4651_), .A3(new_n4676_), .ZN(new_n4680_));
  NAND3_X1   g4631(.A1(new_n4679_), .A2(new_n4680_), .A3(new_n4649_), .ZN(new_n4681_));
  AOI21_X1   g4632(.A1(new_n4679_), .A2(new_n4680_), .B(new_n4649_), .ZN(new_n4682_));
  INV_X1     g4633(.I(new_n4682_), .ZN(new_n4683_));
  NAND3_X1   g4634(.A1(new_n4683_), .A2(new_n4681_), .A3(new_n4645_), .ZN(new_n4684_));
  INV_X1     g4635(.I(new_n4645_), .ZN(new_n4685_));
  INV_X1     g4636(.I(new_n4681_), .ZN(new_n4686_));
  OAI21_X1   g4637(.A1(new_n4686_), .A2(new_n4682_), .B(new_n4685_), .ZN(new_n4687_));
  NAND3_X1   g4638(.A1(new_n4684_), .A2(new_n4687_), .A3(new_n4644_), .ZN(new_n4688_));
  INV_X1     g4639(.I(new_n4644_), .ZN(new_n4689_));
  NOR3_X1    g4640(.A1(new_n4686_), .A2(new_n4682_), .A3(new_n4685_), .ZN(new_n4690_));
  AOI21_X1   g4641(.A1(new_n4683_), .A2(new_n4681_), .B(new_n4645_), .ZN(new_n4691_));
  OAI21_X1   g4642(.A1(new_n4691_), .A2(new_n4690_), .B(new_n4689_), .ZN(new_n4692_));
  NAND3_X1   g4643(.A1(new_n4692_), .A2(new_n4688_), .A3(new_n4641_), .ZN(new_n4693_));
  INV_X1     g4644(.I(new_n4641_), .ZN(new_n4694_));
  NOR3_X1    g4645(.A1(new_n4691_), .A2(new_n4690_), .A3(new_n4689_), .ZN(new_n4695_));
  AOI21_X1   g4646(.A1(new_n4684_), .A2(new_n4687_), .B(new_n4644_), .ZN(new_n4696_));
  OAI21_X1   g4647(.A1(new_n4696_), .A2(new_n4695_), .B(new_n4694_), .ZN(new_n4697_));
  NAND2_X1   g4648(.A1(new_n4697_), .A2(new_n4693_), .ZN(new_n4698_));
  NAND4_X1   g4649(.A1(new_n1024_), .A2(new_n160_), .A3(new_n674_), .A4(new_n989_), .ZN(new_n4699_));
  NAND2_X1   g4650(.A1(new_n2469_), .A2(new_n912_), .ZN(new_n4700_));
  INV_X1     g4651(.I(new_n4700_), .ZN(new_n4701_));
  AND4_X2    g4652(.A1(new_n342_), .A2(new_n2360_), .A3(new_n701_), .A4(new_n2252_), .Z(new_n4702_));
  NAND4_X1   g4653(.A1(new_n4702_), .A2(new_n311_), .A3(new_n4217_), .A4(new_n4701_), .ZN(new_n4703_));
  NOR4_X1    g4654(.A1(new_n2580_), .A2(new_n4093_), .A3(new_n4699_), .A4(new_n4703_), .ZN(new_n4704_));
  INV_X1     g4655(.I(new_n4704_), .ZN(new_n4705_));
  NOR2_X1    g4656(.A1(new_n4698_), .A2(new_n4705_), .ZN(new_n4706_));
  AOI21_X1   g4657(.A1(new_n4697_), .A2(new_n4693_), .B(new_n4704_), .ZN(new_n4707_));
  NOR2_X1    g4658(.A1(new_n4706_), .A2(new_n4707_), .ZN(new_n4708_));
  XOR2_X1    g4659(.A1(new_n4708_), .A2(new_n4640_), .Z(new_n4709_));
  NOR2_X1    g4660(.A1(new_n4606_), .A2(new_n4602_), .ZN(new_n4710_));
  INV_X1     g4661(.I(new_n4710_), .ZN(new_n4711_));
  NOR2_X1    g4662(.A1(new_n4518_), .A2(new_n4711_), .ZN(new_n4712_));
  NOR2_X1    g4663(.A1(new_n4619_), .A2(new_n4710_), .ZN(new_n4713_));
  OAI21_X1   g4664(.A1(new_n4712_), .A2(new_n4713_), .B(new_n4614_), .ZN(new_n4714_));
  OAI21_X1   g4665(.A1(new_n4626_), .A2(new_n4624_), .B(new_n4714_), .ZN(new_n4715_));
  XOR2_X1    g4666(.A1(new_n4709_), .A2(new_n4715_), .Z(new_n4716_));
  XOR2_X1    g4667(.A1(new_n4716_), .A2(new_n4629_), .Z(new_n4717_));
  XNOR2_X1   g4668(.A1(new_n4635_), .A2(new_n4717_), .ZN(\sin[5] ));
  NOR2_X1    g4669(.A1(new_n4634_), .A2(new_n4717_), .ZN(new_n4719_));
  NOR2_X1    g4670(.A1(new_n4719_), .A2(new_n4074_), .ZN(new_n4720_));
  NOR2_X1    g4671(.A1(new_n4716_), .A2(new_n4629_), .ZN(new_n4721_));
  NOR2_X1    g4672(.A1(new_n4640_), .A2(new_n4698_), .ZN(new_n4722_));
  AOI22_X1   g4673(.A1(new_n4638_), .A2(new_n4639_), .B1(new_n4693_), .B2(new_n4697_), .ZN(new_n4723_));
  NOR2_X1    g4674(.A1(new_n4722_), .A2(new_n4723_), .ZN(new_n4724_));
  INV_X1     g4675(.I(new_n4724_), .ZN(new_n4725_));
  NAND3_X1   g4676(.A1(new_n4622_), .A2(new_n4619_), .A3(new_n4616_), .ZN(new_n4726_));
  OAI21_X1   g4677(.A1(new_n4619_), .A2(new_n4622_), .B(new_n4726_), .ZN(new_n4727_));
  AOI21_X1   g4678(.A1(new_n4501_), .A2(new_n4500_), .B(new_n4392_), .ZN(new_n4728_));
  OAI21_X1   g4679(.A1(new_n4505_), .A2(new_n4728_), .B(new_n4502_), .ZN(new_n4729_));
  NAND2_X1   g4680(.A1(new_n4729_), .A2(new_n4727_), .ZN(new_n4730_));
  AOI21_X1   g4681(.A1(new_n4730_), .A2(new_n4714_), .B(new_n4704_), .ZN(new_n4731_));
  NAND3_X1   g4682(.A1(new_n4730_), .A2(new_n4704_), .A3(new_n4714_), .ZN(new_n4732_));
  OAI21_X1   g4683(.A1(new_n4725_), .A2(new_n4731_), .B(new_n4732_), .ZN(new_n4733_));
  AOI21_X1   g4684(.A1(new_n4644_), .A2(new_n4684_), .B(new_n4691_), .ZN(new_n4734_));
  NAND2_X1   g4685(.A1(new_n4677_), .A2(new_n4676_), .ZN(new_n4735_));
  NAND2_X1   g4686(.A1(new_n4735_), .A2(new_n4651_), .ZN(new_n4736_));
  OAI21_X1   g4687(.A1(new_n4735_), .A2(new_n4651_), .B(new_n4649_), .ZN(new_n4737_));
  NAND3_X1   g4688(.A1(new_n4737_), .A2(new_n4736_), .A3(new_n1288_), .ZN(new_n4738_));
  NAND2_X1   g4689(.A1(new_n4737_), .A2(new_n4736_), .ZN(new_n4739_));
  NAND2_X1   g4690(.A1(new_n4739_), .A2(new_n1287_), .ZN(new_n4740_));
  NAND2_X1   g4691(.A1(new_n4740_), .A2(new_n4738_), .ZN(new_n4741_));
  INV_X1     g4692(.I(new_n4741_), .ZN(new_n4742_));
  INV_X1     g4693(.I(new_n4477_), .ZN(new_n4743_));
  AOI22_X1   g4694(.A1(new_n4743_), .A2(new_n3073_), .B1(new_n3056_), .B2(new_n4476_), .ZN(new_n4744_));
  OAI22_X1   g4695(.A1(new_n3869_), .A2(new_n2852_), .B1(new_n2856_), .B2(new_n3573_), .ZN(new_n4745_));
  AOI21_X1   g4696(.A1(new_n2859_), .A2(new_n4001_), .B(new_n4745_), .ZN(new_n4746_));
  NAND2_X1   g4697(.A1(new_n4459_), .A2(new_n2863_), .ZN(new_n4747_));
  NAND2_X1   g4698(.A1(new_n4747_), .A2(new_n4746_), .ZN(new_n4748_));
  XOR2_X1    g4699(.A1(new_n4748_), .A2(new_n845_), .Z(new_n4749_));
  INV_X1     g4700(.I(new_n4661_), .ZN(new_n4750_));
  NOR2_X1    g4701(.A1(new_n4666_), .A2(new_n4674_), .ZN(new_n4751_));
  NAND2_X1   g4702(.A1(new_n4666_), .A2(new_n4674_), .ZN(new_n4752_));
  AOI21_X1   g4703(.A1(new_n4750_), .A2(new_n4752_), .B(new_n4751_), .ZN(new_n4753_));
  INV_X1     g4704(.I(new_n4753_), .ZN(new_n4754_));
  NAND2_X1   g4705(.A1(new_n3578_), .A2(new_n2735_), .ZN(new_n4755_));
  AOI22_X1   g4706(.A1(new_n3538_), .A2(new_n2752_), .B1(new_n2604_), .B2(new_n2738_), .ZN(new_n4756_));
  NAND2_X1   g4707(.A1(new_n3904_), .A2(new_n2748_), .ZN(new_n4757_));
  NAND3_X1   g4708(.A1(new_n4757_), .A2(new_n4755_), .A3(new_n4756_), .ZN(new_n4758_));
  XOR2_X1    g4709(.A1(new_n4758_), .A2(new_n474_), .Z(new_n4759_));
  NOR2_X1    g4710(.A1(new_n2956_), .A2(new_n598_), .ZN(new_n4760_));
  INV_X1     g4711(.I(new_n4760_), .ZN(new_n4761_));
  AOI21_X1   g4712(.A1(new_n4654_), .A2(new_n4657_), .B(new_n4658_), .ZN(new_n4762_));
  NOR2_X1    g4713(.A1(new_n4762_), .A2(new_n52_), .ZN(new_n4763_));
  INV_X1     g4714(.I(new_n4763_), .ZN(new_n4764_));
  NAND2_X1   g4715(.A1(new_n4762_), .A2(new_n52_), .ZN(new_n4765_));
  AND3_X2    g4716(.A1(new_n4764_), .A2(new_n4761_), .A3(new_n4765_), .Z(new_n4766_));
  AOI21_X1   g4717(.A1(new_n4764_), .A2(new_n4765_), .B(new_n4761_), .ZN(new_n4767_));
  AOI22_X1   g4718(.A1(new_n2613_), .A2(new_n2816_), .B1(new_n2704_), .B2(new_n3000_), .ZN(new_n4768_));
  OAI21_X1   g4719(.A1(new_n2611_), .A2(new_n3003_), .B(new_n4768_), .ZN(new_n4769_));
  NOR2_X1    g4720(.A1(new_n3473_), .A2(new_n2820_), .ZN(new_n4770_));
  NOR2_X1    g4721(.A1(new_n4770_), .A2(new_n4769_), .ZN(new_n4771_));
  XOR2_X1    g4722(.A1(new_n4771_), .A2(new_n465_), .Z(new_n4772_));
  OR3_X2     g4723(.A1(new_n4766_), .A2(new_n4767_), .A3(new_n4772_), .Z(new_n4773_));
  OAI21_X1   g4724(.A1(new_n4766_), .A2(new_n4767_), .B(new_n4772_), .ZN(new_n4774_));
  NAND3_X1   g4725(.A1(new_n4773_), .A2(new_n4759_), .A3(new_n4774_), .ZN(new_n4775_));
  INV_X1     g4726(.I(new_n4759_), .ZN(new_n4776_));
  NAND2_X1   g4727(.A1(new_n4773_), .A2(new_n4774_), .ZN(new_n4777_));
  NAND2_X1   g4728(.A1(new_n4777_), .A2(new_n4776_), .ZN(new_n4778_));
  NAND3_X1   g4729(.A1(new_n4754_), .A2(new_n4775_), .A3(new_n4778_), .ZN(new_n4779_));
  NAND2_X1   g4730(.A1(new_n4778_), .A2(new_n4775_), .ZN(new_n4780_));
  NAND2_X1   g4731(.A1(new_n4780_), .A2(new_n4753_), .ZN(new_n4781_));
  NAND2_X1   g4732(.A1(new_n4781_), .A2(new_n4779_), .ZN(new_n4782_));
  NAND2_X1   g4733(.A1(new_n4782_), .A2(new_n4749_), .ZN(new_n4783_));
  INV_X1     g4734(.I(new_n4749_), .ZN(new_n4784_));
  NAND3_X1   g4735(.A1(new_n4781_), .A2(new_n4784_), .A3(new_n4779_), .ZN(new_n4785_));
  AOI21_X1   g4736(.A1(new_n4783_), .A2(new_n4785_), .B(new_n4744_), .ZN(new_n4786_));
  INV_X1     g4737(.I(new_n4786_), .ZN(new_n4787_));
  NAND3_X1   g4738(.A1(new_n4783_), .A2(new_n4785_), .A3(new_n4744_), .ZN(new_n4788_));
  NAND3_X1   g4739(.A1(new_n4742_), .A2(new_n4787_), .A3(new_n4788_), .ZN(new_n4789_));
  INV_X1     g4740(.I(new_n4788_), .ZN(new_n4790_));
  OAI21_X1   g4741(.A1(new_n4790_), .A2(new_n4786_), .B(new_n4741_), .ZN(new_n4791_));
  NAND3_X1   g4742(.A1(new_n4789_), .A2(new_n4791_), .A3(new_n4734_), .ZN(new_n4792_));
  OAI21_X1   g4743(.A1(new_n4689_), .A2(new_n4690_), .B(new_n4687_), .ZN(new_n4793_));
  NOR3_X1    g4744(.A1(new_n4790_), .A2(new_n4741_), .A3(new_n4786_), .ZN(new_n4794_));
  AOI21_X1   g4745(.A1(new_n4787_), .A2(new_n4788_), .B(new_n4742_), .ZN(new_n4795_));
  OAI21_X1   g4746(.A1(new_n4795_), .A2(new_n4794_), .B(new_n4793_), .ZN(new_n4796_));
  NAND2_X1   g4747(.A1(new_n4796_), .A2(new_n4792_), .ZN(new_n4797_));
  AOI21_X1   g4748(.A1(new_n4692_), .A2(new_n4688_), .B(new_n4694_), .ZN(new_n4798_));
  INV_X1     g4749(.I(new_n4637_), .ZN(new_n4799_));
  AOI21_X1   g4750(.A1(new_n4619_), .A2(new_n4799_), .B(new_n4603_), .ZN(new_n4800_));
  NOR2_X1    g4751(.A1(new_n4619_), .A2(new_n4799_), .ZN(new_n4801_));
  NOR3_X1    g4752(.A1(new_n4696_), .A2(new_n4695_), .A3(new_n4641_), .ZN(new_n4802_));
  NOR3_X1    g4753(.A1(new_n4800_), .A2(new_n4801_), .A3(new_n4802_), .ZN(new_n4803_));
  NOR2_X1    g4754(.A1(new_n4803_), .A2(new_n4798_), .ZN(new_n4804_));
  NAND2_X1   g4755(.A1(new_n4804_), .A2(new_n4797_), .ZN(new_n4805_));
  NOR3_X1    g4756(.A1(new_n4795_), .A2(new_n4793_), .A3(new_n4794_), .ZN(new_n4806_));
  AOI21_X1   g4757(.A1(new_n4789_), .A2(new_n4791_), .B(new_n4734_), .ZN(new_n4807_));
  NOR2_X1    g4758(.A1(new_n4806_), .A2(new_n4807_), .ZN(new_n4808_));
  INV_X1     g4759(.I(new_n4798_), .ZN(new_n4809_));
  NAND3_X1   g4760(.A1(new_n4692_), .A2(new_n4688_), .A3(new_n4694_), .ZN(new_n4810_));
  NAND3_X1   g4761(.A1(new_n4638_), .A2(new_n4639_), .A3(new_n4810_), .ZN(new_n4811_));
  NAND2_X1   g4762(.A1(new_n4811_), .A2(new_n4809_), .ZN(new_n4812_));
  NAND2_X1   g4763(.A1(new_n4812_), .A2(new_n4808_), .ZN(new_n4813_));
  NOR4_X1    g4764(.A1(new_n854_), .A2(new_n191_), .A3(new_n207_), .A4(new_n376_), .ZN(new_n4814_));
  INV_X1     g4765(.I(new_n4814_), .ZN(new_n4815_));
  NOR4_X1    g4766(.A1(new_n2464_), .A2(new_n291_), .A3(new_n1120_), .A4(new_n3564_), .ZN(new_n4816_));
  INV_X1     g4767(.I(new_n4816_), .ZN(new_n4817_));
  NOR3_X1    g4768(.A1(new_n2380_), .A2(new_n881_), .A3(new_n1154_), .ZN(new_n4818_));
  NOR4_X1    g4769(.A1(new_n2253_), .A2(new_n437_), .A3(new_n567_), .A4(new_n914_), .ZN(new_n4819_));
  AND4_X2    g4770(.A1(new_n550_), .A2(new_n2468_), .A3(new_n4818_), .A4(new_n4819_), .Z(new_n4820_));
  NAND2_X1   g4771(.A1(new_n4820_), .A2(new_n2440_), .ZN(new_n4821_));
  NOR4_X1    g4772(.A1(new_n4821_), .A2(new_n3769_), .A3(new_n4815_), .A4(new_n4817_), .ZN(new_n4822_));
  NAND3_X1   g4773(.A1(new_n4813_), .A2(new_n4805_), .A3(new_n4822_), .ZN(new_n4823_));
  NOR2_X1    g4774(.A1(new_n4812_), .A2(new_n4808_), .ZN(new_n4824_));
  NOR2_X1    g4775(.A1(new_n4804_), .A2(new_n4797_), .ZN(new_n4825_));
  INV_X1     g4776(.I(new_n4822_), .ZN(new_n4826_));
  OAI21_X1   g4777(.A1(new_n4824_), .A2(new_n4825_), .B(new_n4826_), .ZN(new_n4827_));
  NAND2_X1   g4778(.A1(new_n4827_), .A2(new_n4823_), .ZN(new_n4828_));
  XOR2_X1    g4779(.A1(new_n4828_), .A2(new_n4733_), .Z(new_n4829_));
  NOR2_X1    g4780(.A1(new_n4721_), .A2(new_n4829_), .ZN(new_n4830_));
  NAND2_X1   g4781(.A1(new_n4721_), .A2(new_n4829_), .ZN(new_n4831_));
  INV_X1     g4782(.I(new_n4831_), .ZN(new_n4832_));
  NOR2_X1    g4783(.A1(new_n4832_), .A2(new_n4830_), .ZN(new_n4833_));
  XOR2_X1    g4784(.A1(new_n4720_), .A2(new_n4833_), .Z(\sin[6] ));
  INV_X1     g4785(.I(new_n4719_), .ZN(new_n4835_));
  OAI21_X1   g4786(.A1(new_n4835_), .A2(new_n4833_), .B(new_n4073_), .ZN(new_n4836_));
  OAI21_X1   g4787(.A1(new_n4803_), .A2(new_n4798_), .B(new_n4797_), .ZN(new_n4837_));
  AOI21_X1   g4788(.A1(new_n4789_), .A2(new_n4791_), .B(new_n4793_), .ZN(new_n4838_));
  INV_X1     g4789(.I(new_n4838_), .ZN(new_n4839_));
  NAND2_X1   g4790(.A1(new_n4837_), .A2(new_n4839_), .ZN(new_n4840_));
  INV_X1     g4791(.I(new_n4739_), .ZN(new_n4841_));
  NAND2_X1   g4792(.A1(new_n4783_), .A2(new_n4785_), .ZN(new_n4842_));
  NOR2_X1    g4793(.A1(new_n4842_), .A2(new_n4841_), .ZN(new_n4843_));
  XOR2_X1    g4794(.A1(new_n4744_), .A2(new_n1288_), .Z(new_n4844_));
  AOI21_X1   g4795(.A1(new_n4842_), .A2(new_n4841_), .B(new_n4844_), .ZN(new_n4845_));
  NOR2_X1    g4796(.A1(new_n4845_), .A2(new_n4843_), .ZN(new_n4846_));
  AOI21_X1   g4797(.A1(new_n4775_), .A2(new_n4778_), .B(new_n4754_), .ZN(new_n4847_));
  OAI21_X1   g4798(.A1(new_n4847_), .A2(new_n4749_), .B(new_n4779_), .ZN(new_n4848_));
  INV_X1     g4799(.I(new_n4848_), .ZN(new_n4849_));
  AOI22_X1   g4800(.A1(new_n4001_), .A2(new_n2851_), .B1(new_n3868_), .B2(new_n2855_), .ZN(new_n4850_));
  OAI21_X1   g4801(.A1(new_n2860_), .A2(new_n4098_), .B(new_n4850_), .ZN(new_n4851_));
  NOR2_X1    g4802(.A1(new_n4110_), .A2(new_n4108_), .ZN(new_n4852_));
  NOR2_X1    g4803(.A1(new_n4852_), .A2(new_n2880_), .ZN(new_n4853_));
  NOR2_X1    g4804(.A1(new_n4853_), .A2(new_n4851_), .ZN(new_n4854_));
  XOR2_X1    g4805(.A1(new_n4854_), .A2(new_n845_), .Z(new_n4855_));
  INV_X1     g4806(.I(new_n4855_), .ZN(new_n4856_));
  NAND2_X1   g4807(.A1(new_n4773_), .A2(new_n4759_), .ZN(new_n4857_));
  NAND2_X1   g4808(.A1(new_n4857_), .A2(new_n4774_), .ZN(new_n4858_));
  NOR2_X1    g4809(.A1(new_n3584_), .A2(new_n3588_), .ZN(new_n4859_));
  OAI22_X1   g4810(.A1(new_n2598_), .A2(new_n2739_), .B1(new_n2586_), .B2(new_n2768_), .ZN(new_n4860_));
  AOI21_X1   g4811(.A1(new_n2735_), .A2(new_n3859_), .B(new_n4860_), .ZN(new_n4861_));
  OAI21_X1   g4812(.A1(new_n4859_), .A2(new_n2743_), .B(new_n4861_), .ZN(new_n4862_));
  XOR2_X1    g4813(.A1(new_n4862_), .A2(new_n474_), .Z(new_n4863_));
  INV_X1     g4814(.I(new_n4863_), .ZN(new_n4864_));
  NOR2_X1    g4815(.A1(new_n4761_), .A2(new_n2725_), .ZN(new_n4865_));
  AOI21_X1   g4816(.A1(new_n2725_), .A2(new_n4761_), .B(new_n4762_), .ZN(new_n4866_));
  NOR2_X1    g4817(.A1(new_n4866_), .A2(new_n4865_), .ZN(new_n4867_));
  OAI22_X1   g4818(.A1(new_n2563_), .A2(new_n3003_), .B1(new_n2694_), .B2(new_n3001_), .ZN(new_n4868_));
  NOR2_X1    g4819(.A1(new_n2611_), .A2(new_n2815_), .ZN(new_n4869_));
  NOR2_X1    g4820(.A1(new_n3599_), .A2(new_n2820_), .ZN(new_n4870_));
  NOR3_X1    g4821(.A1(new_n4870_), .A2(new_n4868_), .A3(new_n4869_), .ZN(new_n4871_));
  XOR2_X1    g4822(.A1(new_n4871_), .A2(new_n598_), .Z(new_n4872_));
  NOR2_X1    g4823(.A1(new_n2666_), .A2(new_n598_), .ZN(new_n4873_));
  XOR2_X1    g4824(.A1(new_n1287_), .A2(new_n2725_), .Z(new_n4874_));
  XOR2_X1    g4825(.A1(new_n4873_), .A2(new_n4874_), .Z(new_n4875_));
  INV_X1     g4826(.I(new_n4875_), .ZN(new_n4876_));
  NAND2_X1   g4827(.A1(new_n4872_), .A2(new_n4876_), .ZN(new_n4877_));
  XOR2_X1    g4828(.A1(new_n4871_), .A2(new_n465_), .Z(new_n4878_));
  NAND2_X1   g4829(.A1(new_n4878_), .A2(new_n4875_), .ZN(new_n4879_));
  NAND3_X1   g4830(.A1(new_n4877_), .A2(new_n4879_), .A3(new_n4867_), .ZN(new_n4880_));
  NOR2_X1    g4831(.A1(new_n4878_), .A2(new_n4875_), .ZN(new_n4881_));
  NOR2_X1    g4832(.A1(new_n4872_), .A2(new_n4876_), .ZN(new_n4882_));
  OAI22_X1   g4833(.A1(new_n4881_), .A2(new_n4882_), .B1(new_n4865_), .B2(new_n4866_), .ZN(new_n4883_));
  NAND2_X1   g4834(.A1(new_n4883_), .A2(new_n4880_), .ZN(new_n4884_));
  NAND2_X1   g4835(.A1(new_n4884_), .A2(new_n4864_), .ZN(new_n4885_));
  NAND3_X1   g4836(.A1(new_n4883_), .A2(new_n4880_), .A3(new_n4863_), .ZN(new_n4886_));
  NAND2_X1   g4837(.A1(new_n4885_), .A2(new_n4886_), .ZN(new_n4887_));
  NOR2_X1    g4838(.A1(new_n4887_), .A2(new_n4858_), .ZN(new_n4888_));
  AOI22_X1   g4839(.A1(new_n4885_), .A2(new_n4886_), .B1(new_n4774_), .B2(new_n4857_), .ZN(new_n4889_));
  NOR2_X1    g4840(.A1(new_n4888_), .A2(new_n4889_), .ZN(new_n4890_));
  NOR2_X1    g4841(.A1(new_n4890_), .A2(new_n4856_), .ZN(new_n4891_));
  INV_X1     g4842(.I(new_n4891_), .ZN(new_n4892_));
  NAND2_X1   g4843(.A1(new_n4890_), .A2(new_n4856_), .ZN(new_n4893_));
  NAND3_X1   g4844(.A1(new_n4892_), .A2(new_n4849_), .A3(new_n4893_), .ZN(new_n4894_));
  INV_X1     g4845(.I(new_n4893_), .ZN(new_n4895_));
  OAI21_X1   g4846(.A1(new_n4895_), .A2(new_n4891_), .B(new_n4848_), .ZN(new_n4896_));
  NAND3_X1   g4847(.A1(new_n4846_), .A2(new_n4894_), .A3(new_n4896_), .ZN(new_n4897_));
  AOI21_X1   g4848(.A1(new_n4896_), .A2(new_n4894_), .B(new_n4846_), .ZN(new_n4898_));
  INV_X1     g4849(.I(new_n4898_), .ZN(new_n4899_));
  NOR4_X1    g4850(.A1(new_n387_), .A2(new_n2356_), .A3(new_n723_), .A4(new_n201_), .ZN(new_n4900_));
  NOR3_X1    g4851(.A1(new_n924_), .A2(new_n443_), .A3(new_n515_), .ZN(new_n4901_));
  NAND4_X1   g4852(.A1(new_n690_), .A2(new_n4901_), .A3(new_n350_), .A4(new_n578_), .ZN(new_n4902_));
  NAND2_X1   g4853(.A1(new_n2343_), .A2(new_n4820_), .ZN(new_n4903_));
  NOR2_X1    g4854(.A1(new_n4903_), .A2(new_n4902_), .ZN(new_n4904_));
  AND3_X2    g4855(.A1(new_n4904_), .A2(new_n4701_), .A3(new_n4900_), .Z(new_n4905_));
  NAND3_X1   g4856(.A1(new_n4899_), .A2(new_n4897_), .A3(new_n4905_), .ZN(new_n4906_));
  AOI21_X1   g4857(.A1(new_n4899_), .A2(new_n4897_), .B(new_n4905_), .ZN(new_n4907_));
  INV_X1     g4858(.I(new_n4907_), .ZN(new_n4908_));
  NAND2_X1   g4859(.A1(new_n4908_), .A2(new_n4906_), .ZN(new_n4909_));
  XOR2_X1    g4860(.A1(new_n4909_), .A2(new_n4840_), .Z(new_n4910_));
  NOR3_X1    g4861(.A1(new_n4824_), .A2(new_n4825_), .A3(new_n4826_), .ZN(new_n4911_));
  OAI21_X1   g4862(.A1(new_n4733_), .A2(new_n4911_), .B(new_n4827_), .ZN(new_n4912_));
  NAND2_X1   g4863(.A1(new_n4912_), .A2(new_n4910_), .ZN(new_n4913_));
  XNOR2_X1   g4864(.A1(new_n4909_), .A2(new_n4840_), .ZN(new_n4914_));
  NAND2_X1   g4865(.A1(new_n4715_), .A2(new_n4705_), .ZN(new_n4915_));
  NOR2_X1    g4866(.A1(new_n4715_), .A2(new_n4705_), .ZN(new_n4916_));
  AOI21_X1   g4867(.A1(new_n4724_), .A2(new_n4915_), .B(new_n4916_), .ZN(new_n4917_));
  AOI21_X1   g4868(.A1(new_n4813_), .A2(new_n4805_), .B(new_n4822_), .ZN(new_n4918_));
  AOI21_X1   g4869(.A1(new_n4917_), .A2(new_n4823_), .B(new_n4918_), .ZN(new_n4919_));
  NAND2_X1   g4870(.A1(new_n4919_), .A2(new_n4914_), .ZN(new_n4920_));
  NAND2_X1   g4871(.A1(new_n4913_), .A2(new_n4920_), .ZN(new_n4921_));
  XNOR2_X1   g4872(.A1(new_n4831_), .A2(new_n4921_), .ZN(new_n4922_));
  XOR2_X1    g4873(.A1(new_n4836_), .A2(new_n4922_), .Z(\sin[7] ));
  AND2_X2    g4874(.A1(new_n4830_), .A2(new_n4921_), .Z(new_n4924_));
  NAND4_X1   g4875(.A1(new_n4721_), .A2(new_n4829_), .A3(new_n4913_), .A4(new_n4920_), .ZN(new_n4925_));
  INV_X1     g4876(.I(new_n4925_), .ZN(new_n4926_));
  OAI21_X1   g4877(.A1(new_n4924_), .A2(new_n4926_), .B(new_n4719_), .ZN(new_n4927_));
  NAND2_X1   g4878(.A1(new_n4927_), .A2(new_n4073_), .ZN(new_n4928_));
  INV_X1     g4879(.I(new_n4905_), .ZN(new_n4929_));
  AOI21_X1   g4880(.A1(new_n4811_), .A2(new_n4809_), .B(new_n4808_), .ZN(new_n4930_));
  NOR2_X1    g4881(.A1(new_n4930_), .A2(new_n4838_), .ZN(new_n4931_));
  NAND2_X1   g4882(.A1(new_n4899_), .A2(new_n4897_), .ZN(new_n4932_));
  INV_X1     g4883(.I(new_n4932_), .ZN(new_n4933_));
  NOR2_X1    g4884(.A1(new_n4931_), .A2(new_n4933_), .ZN(new_n4934_));
  NOR2_X1    g4885(.A1(new_n4840_), .A2(new_n4932_), .ZN(new_n4935_));
  OAI21_X1   g4886(.A1(new_n4934_), .A2(new_n4935_), .B(new_n4929_), .ZN(new_n4936_));
  OAI21_X1   g4887(.A1(new_n4919_), .A2(new_n4914_), .B(new_n4936_), .ZN(new_n4937_));
  NOR2_X1    g4888(.A1(new_n193_), .A2(new_n415_), .ZN(new_n4938_));
  NOR3_X1    g4889(.A1(new_n197_), .A2(new_n127_), .A3(new_n435_), .ZN(new_n4939_));
  AND4_X2    g4890(.A1(new_n240_), .A2(new_n4939_), .A3(new_n911_), .A4(new_n4938_), .Z(new_n4940_));
  NAND4_X1   g4891(.A1(new_n4940_), .A2(new_n855_), .A3(new_n882_), .A4(new_n2385_), .ZN(new_n4941_));
  NAND2_X1   g4892(.A1(new_n2326_), .A2(new_n1433_), .ZN(new_n4942_));
  NAND3_X1   g4893(.A1(new_n1111_), .A2(new_n2332_), .A3(new_n1068_), .ZN(new_n4943_));
  NOR4_X1    g4894(.A1(new_n4942_), .A2(new_n345_), .A3(new_n4943_), .A4(new_n984_), .ZN(new_n4944_));
  NAND3_X1   g4895(.A1(new_n2458_), .A2(new_n4944_), .A3(new_n2285_), .ZN(new_n4945_));
  NOR3_X1    g4896(.A1(new_n3738_), .A2(new_n4941_), .A3(new_n4945_), .ZN(new_n4946_));
  INV_X1     g4897(.I(new_n4946_), .ZN(new_n4947_));
  NAND3_X1   g4898(.A1(new_n4837_), .A2(new_n4839_), .A3(new_n4897_), .ZN(new_n4948_));
  NAND2_X1   g4899(.A1(new_n4948_), .A2(new_n4899_), .ZN(new_n4949_));
  OAI21_X1   g4900(.A1(new_n4895_), .A2(new_n4849_), .B(new_n4892_), .ZN(new_n4950_));
  INV_X1     g4901(.I(new_n4950_), .ZN(new_n4951_));
  AOI22_X1   g4902(.A1(new_n4476_), .A2(new_n2851_), .B1(new_n2855_), .B2(new_n4001_), .ZN(new_n4952_));
  OAI21_X1   g4903(.A1(new_n4341_), .A2(new_n2880_), .B(new_n4952_), .ZN(new_n4953_));
  XOR2_X1    g4904(.A1(new_n4953_), .A2(new_n845_), .Z(new_n4954_));
  INV_X1     g4905(.I(new_n4954_), .ZN(new_n4955_));
  OAI22_X1   g4906(.A1(new_n3573_), .A2(new_n2739_), .B1(new_n2598_), .B2(new_n2768_), .ZN(new_n4956_));
  AOI21_X1   g4907(.A1(new_n3868_), .A2(new_n2735_), .B(new_n4956_), .ZN(new_n4957_));
  OAI21_X1   g4908(.A1(new_n3885_), .A2(new_n2743_), .B(new_n4957_), .ZN(new_n4958_));
  XOR2_X1    g4909(.A1(new_n4958_), .A2(new_n473_), .Z(new_n4959_));
  INV_X1     g4910(.I(new_n4959_), .ZN(new_n4960_));
  AOI21_X1   g4911(.A1(new_n4867_), .A2(new_n4877_), .B(new_n4882_), .ZN(new_n4961_));
  OAI22_X1   g4912(.A1(new_n2563_), .A2(new_n2815_), .B1(new_n2611_), .B2(new_n3001_), .ZN(new_n4962_));
  AOI21_X1   g4913(.A1(new_n2604_), .A2(new_n2812_), .B(new_n4962_), .ZN(new_n4963_));
  NAND2_X1   g4914(.A1(new_n4273_), .A2(new_n2819_), .ZN(new_n4964_));
  NAND2_X1   g4915(.A1(new_n4964_), .A2(new_n4963_), .ZN(new_n4965_));
  XOR2_X1    g4916(.A1(new_n4965_), .A2(new_n465_), .Z(new_n4966_));
  AOI21_X1   g4917(.A1(new_n2725_), .A2(new_n1288_), .B(new_n4873_), .ZN(new_n4967_));
  AOI21_X1   g4918(.A1(new_n52_), .A2(new_n1287_), .B(new_n4967_), .ZN(new_n4968_));
  NOR2_X1    g4919(.A1(new_n2694_), .A2(new_n598_), .ZN(new_n4969_));
  INV_X1     g4920(.I(new_n4969_), .ZN(new_n4970_));
  NOR2_X1    g4921(.A1(new_n4968_), .A2(new_n4970_), .ZN(new_n4971_));
  NAND2_X1   g4922(.A1(new_n4968_), .A2(new_n4970_), .ZN(new_n4972_));
  INV_X1     g4923(.I(new_n4972_), .ZN(new_n4973_));
  NOR2_X1    g4924(.A1(new_n4973_), .A2(new_n4971_), .ZN(new_n4974_));
  XOR2_X1    g4925(.A1(new_n4966_), .A2(new_n4974_), .Z(new_n4975_));
  NAND2_X1   g4926(.A1(new_n4975_), .A2(new_n4961_), .ZN(new_n4976_));
  OR2_X2     g4927(.A1(new_n4975_), .A2(new_n4961_), .Z(new_n4977_));
  NAND2_X1   g4928(.A1(new_n4977_), .A2(new_n4976_), .ZN(new_n4978_));
  XOR2_X1    g4929(.A1(new_n4978_), .A2(new_n4960_), .Z(new_n4979_));
  OAI21_X1   g4930(.A1(new_n4887_), .A2(new_n4858_), .B(new_n4885_), .ZN(new_n4980_));
  NAND2_X1   g4931(.A1(new_n4979_), .A2(new_n4980_), .ZN(new_n4981_));
  OR2_X2     g4932(.A1(new_n4979_), .A2(new_n4980_), .Z(new_n4982_));
  NAND2_X1   g4933(.A1(new_n4982_), .A2(new_n4981_), .ZN(new_n4983_));
  XOR2_X1    g4934(.A1(new_n4983_), .A2(new_n4955_), .Z(new_n4984_));
  NOR2_X1    g4935(.A1(new_n4984_), .A2(new_n4951_), .ZN(new_n4985_));
  NAND2_X1   g4936(.A1(new_n4984_), .A2(new_n4951_), .ZN(new_n4986_));
  INV_X1     g4937(.I(new_n4986_), .ZN(new_n4987_));
  NOR2_X1    g4938(.A1(new_n4987_), .A2(new_n4985_), .ZN(new_n4988_));
  NOR2_X1    g4939(.A1(new_n4949_), .A2(new_n4988_), .ZN(new_n4989_));
  NAND2_X1   g4940(.A1(new_n4949_), .A2(new_n4988_), .ZN(new_n4990_));
  INV_X1     g4941(.I(new_n4990_), .ZN(new_n4991_));
  NOR3_X1    g4942(.A1(new_n4991_), .A2(new_n4989_), .A3(new_n4947_), .ZN(new_n4992_));
  INV_X1     g4943(.I(new_n4897_), .ZN(new_n4993_));
  NOR3_X1    g4944(.A1(new_n4930_), .A2(new_n4838_), .A3(new_n4993_), .ZN(new_n4994_));
  NOR2_X1    g4945(.A1(new_n4994_), .A2(new_n4898_), .ZN(new_n4995_));
  INV_X1     g4946(.I(new_n4988_), .ZN(new_n4996_));
  NAND2_X1   g4947(.A1(new_n4996_), .A2(new_n4995_), .ZN(new_n4997_));
  AOI21_X1   g4948(.A1(new_n4997_), .A2(new_n4990_), .B(new_n4946_), .ZN(new_n4998_));
  OAI21_X1   g4949(.A1(new_n4992_), .A2(new_n4998_), .B(new_n4937_), .ZN(new_n4999_));
  NAND2_X1   g4950(.A1(new_n4840_), .A2(new_n4932_), .ZN(new_n5000_));
  NAND2_X1   g4951(.A1(new_n4931_), .A2(new_n4933_), .ZN(new_n5001_));
  AOI21_X1   g4952(.A1(new_n5001_), .A2(new_n5000_), .B(new_n4905_), .ZN(new_n5002_));
  AOI21_X1   g4953(.A1(new_n4912_), .A2(new_n4910_), .B(new_n5002_), .ZN(new_n5003_));
  NAND3_X1   g4954(.A1(new_n4997_), .A2(new_n4990_), .A3(new_n4946_), .ZN(new_n5004_));
  OAI21_X1   g4955(.A1(new_n4991_), .A2(new_n4989_), .B(new_n4947_), .ZN(new_n5005_));
  NAND3_X1   g4956(.A1(new_n5003_), .A2(new_n5005_), .A3(new_n5004_), .ZN(new_n5006_));
  NAND2_X1   g4957(.A1(new_n4999_), .A2(new_n5006_), .ZN(new_n5007_));
  NAND2_X1   g4958(.A1(new_n4926_), .A2(new_n5007_), .ZN(new_n5008_));
  NAND3_X1   g4959(.A1(new_n4925_), .A2(new_n4999_), .A3(new_n5006_), .ZN(new_n5009_));
  NAND2_X1   g4960(.A1(new_n5008_), .A2(new_n5009_), .ZN(new_n5010_));
  XOR2_X1    g4961(.A1(new_n4928_), .A2(new_n5010_), .Z(\sin[8] ));
  AOI21_X1   g4962(.A1(new_n5008_), .A2(new_n5009_), .B(new_n4927_), .ZN(new_n5012_));
  NOR2_X1    g4963(.A1(new_n5012_), .A2(new_n4074_), .ZN(new_n5013_));
  OAI21_X1   g4964(.A1(new_n5003_), .A2(new_n4992_), .B(new_n5005_), .ZN(new_n5014_));
  NOR4_X1    g4965(.A1(new_n452_), .A2(new_n346_), .A3(new_n330_), .A4(new_n425_), .ZN(new_n5015_));
  NOR4_X1    g4966(.A1(new_n2571_), .A2(new_n179_), .A3(new_n207_), .A4(new_n381_), .ZN(new_n5016_));
  NAND4_X1   g4967(.A1(new_n5016_), .A2(new_n690_), .A3(new_n3563_), .A4(new_n5015_), .ZN(new_n5017_));
  NOR3_X1    g4968(.A1(new_n3771_), .A2(new_n2472_), .A3(new_n5017_), .ZN(new_n5018_));
  AND2_X2    g4969(.A1(new_n5018_), .A2(new_n728_), .Z(new_n5019_));
  NAND2_X1   g4970(.A1(new_n4981_), .A2(new_n4955_), .ZN(new_n5020_));
  NAND2_X1   g4971(.A1(new_n5020_), .A2(new_n4982_), .ZN(new_n5021_));
  NAND2_X1   g4972(.A1(new_n4976_), .A2(new_n4960_), .ZN(new_n5022_));
  NAND2_X1   g4973(.A1(new_n5022_), .A2(new_n4977_), .ZN(new_n5023_));
  XOR2_X1    g4974(.A1(new_n5023_), .A2(new_n845_), .Z(new_n5024_));
  OAI22_X1   g4975(.A1(new_n3869_), .A2(new_n2739_), .B1(new_n2768_), .B2(new_n3573_), .ZN(new_n5025_));
  AOI21_X1   g4976(.A1(new_n2735_), .A2(new_n4001_), .B(new_n5025_), .ZN(new_n5026_));
  NAND2_X1   g4977(.A1(new_n4459_), .A2(new_n2748_), .ZN(new_n5027_));
  NAND2_X1   g4978(.A1(new_n5027_), .A2(new_n5026_), .ZN(new_n5028_));
  XOR2_X1    g4979(.A1(new_n5028_), .A2(new_n473_), .Z(new_n5029_));
  INV_X1     g4980(.I(new_n4971_), .ZN(new_n5030_));
  OAI21_X1   g4981(.A1(new_n4966_), .A2(new_n4973_), .B(new_n5030_), .ZN(new_n5031_));
  OAI22_X1   g4982(.A1(new_n2586_), .A2(new_n2815_), .B1(new_n2563_), .B2(new_n3001_), .ZN(new_n5032_));
  AOI21_X1   g4983(.A1(new_n3578_), .A2(new_n2812_), .B(new_n5032_), .ZN(new_n5033_));
  OAI21_X1   g4984(.A1(new_n3908_), .A2(new_n2820_), .B(new_n5033_), .ZN(new_n5034_));
  XOR2_X1    g4985(.A1(new_n5034_), .A2(new_n598_), .Z(new_n5035_));
  OAI21_X1   g4986(.A1(new_n3070_), .A2(new_n3071_), .B(new_n465_), .ZN(new_n5036_));
  XOR2_X1    g4987(.A1(new_n5035_), .A2(new_n5036_), .Z(new_n5037_));
  AND2_X2    g4988(.A1(new_n5037_), .A2(new_n5031_), .Z(new_n5038_));
  NOR2_X1    g4989(.A1(new_n5037_), .A2(new_n5031_), .ZN(new_n5039_));
  NOR2_X1    g4990(.A1(new_n5038_), .A2(new_n5039_), .ZN(new_n5040_));
  XOR2_X1    g4991(.A1(new_n5040_), .A2(new_n5029_), .Z(new_n5041_));
  AOI22_X1   g4992(.A1(new_n4743_), .A2(new_n2863_), .B1(new_n2855_), .B2(new_n4476_), .ZN(new_n5042_));
  XOR2_X1    g4993(.A1(new_n5041_), .A2(new_n5042_), .Z(new_n5043_));
  XNOR2_X1   g4994(.A1(new_n5043_), .A2(new_n5024_), .ZN(new_n5044_));
  NOR2_X1    g4995(.A1(new_n5044_), .A2(new_n5021_), .ZN(new_n5045_));
  INV_X1     g4996(.I(new_n5045_), .ZN(new_n5046_));
  NAND2_X1   g4997(.A1(new_n5044_), .A2(new_n5021_), .ZN(new_n5047_));
  NAND2_X1   g4998(.A1(new_n5046_), .A2(new_n5047_), .ZN(new_n5048_));
  INV_X1     g4999(.I(new_n4985_), .ZN(new_n5049_));
  NAND3_X1   g5000(.A1(new_n4948_), .A2(new_n4899_), .A3(new_n5049_), .ZN(new_n5050_));
  AOI21_X1   g5001(.A1(new_n5050_), .A2(new_n4986_), .B(new_n5048_), .ZN(new_n5051_));
  INV_X1     g5002(.I(new_n5048_), .ZN(new_n5052_));
  NOR3_X1    g5003(.A1(new_n4994_), .A2(new_n4898_), .A3(new_n4985_), .ZN(new_n5053_));
  NOR3_X1    g5004(.A1(new_n5053_), .A2(new_n4987_), .A3(new_n5052_), .ZN(new_n5054_));
  OAI21_X1   g5005(.A1(new_n5054_), .A2(new_n5051_), .B(new_n5019_), .ZN(new_n5055_));
  NOR3_X1    g5006(.A1(new_n5054_), .A2(new_n5051_), .A3(new_n5019_), .ZN(new_n5056_));
  INV_X1     g5007(.I(new_n5056_), .ZN(new_n5057_));
  NAND2_X1   g5008(.A1(new_n5057_), .A2(new_n5055_), .ZN(new_n5058_));
  NAND2_X1   g5009(.A1(new_n5058_), .A2(new_n5014_), .ZN(new_n5059_));
  AOI21_X1   g5010(.A1(new_n4937_), .A2(new_n5004_), .B(new_n4998_), .ZN(new_n5060_));
  NAND3_X1   g5011(.A1(new_n5060_), .A2(new_n5055_), .A3(new_n5057_), .ZN(new_n5061_));
  NAND2_X1   g5012(.A1(new_n5059_), .A2(new_n5061_), .ZN(new_n5062_));
  INV_X1     g5013(.I(new_n5062_), .ZN(new_n5063_));
  NAND2_X1   g5014(.A1(new_n5063_), .A2(new_n5008_), .ZN(new_n5064_));
  AOI21_X1   g5015(.A1(new_n4999_), .A2(new_n5006_), .B(new_n4925_), .ZN(new_n5065_));
  NAND2_X1   g5016(.A1(new_n5065_), .A2(new_n5062_), .ZN(new_n5066_));
  NAND2_X1   g5017(.A1(new_n5064_), .A2(new_n5066_), .ZN(new_n5067_));
  XNOR2_X1   g5018(.A1(new_n5013_), .A2(new_n5067_), .ZN(\sin[9] ));
  AOI21_X1   g5019(.A1(new_n5012_), .A2(new_n5067_), .B(new_n4074_), .ZN(new_n5069_));
  INV_X1     g5020(.I(new_n5055_), .ZN(new_n5070_));
  OAI21_X1   g5021(.A1(new_n5060_), .A2(new_n5070_), .B(new_n5057_), .ZN(new_n5071_));
  INV_X1     g5022(.I(new_n537_), .ZN(new_n5072_));
  NAND4_X1   g5023(.A1(new_n2567_), .A2(new_n676_), .A3(new_n329_), .A4(new_n890_), .ZN(new_n5073_));
  NOR4_X1    g5024(.A1(new_n5073_), .A2(new_n168_), .A3(new_n735_), .A4(new_n881_), .ZN(new_n5074_));
  NAND4_X1   g5025(.A1(new_n5074_), .A2(new_n427_), .A3(new_n2261_), .A4(new_n3563_), .ZN(new_n5075_));
  NOR4_X1    g5026(.A1(new_n5075_), .A2(new_n5072_), .A3(new_n1143_), .A4(new_n3746_), .ZN(new_n5076_));
  INV_X1     g5027(.I(new_n5023_), .ZN(new_n5077_));
  NOR2_X1    g5028(.A1(new_n5041_), .A2(new_n5077_), .ZN(new_n5078_));
  XOR2_X1    g5029(.A1(new_n5042_), .A2(new_n846_), .Z(new_n5079_));
  AOI21_X1   g5030(.A1(new_n5041_), .A2(new_n5077_), .B(new_n5079_), .ZN(new_n5080_));
  NOR2_X1    g5031(.A1(new_n5080_), .A2(new_n5078_), .ZN(new_n5081_));
  NOR2_X1    g5032(.A1(new_n2563_), .A2(new_n598_), .ZN(new_n5082_));
  NOR2_X1    g5033(.A1(new_n4970_), .A2(new_n845_), .ZN(new_n5083_));
  NOR2_X1    g5034(.A1(new_n4969_), .A2(new_n846_), .ZN(new_n5084_));
  OR2_X2     g5035(.A1(new_n5083_), .A2(new_n5084_), .Z(new_n5085_));
  XNOR2_X1   g5036(.A1(new_n5085_), .A2(new_n5082_), .ZN(new_n5086_));
  AOI21_X1   g5037(.A1(new_n2611_), .A2(new_n4969_), .B(new_n5035_), .ZN(new_n5087_));
  NOR2_X1    g5038(.A1(new_n3066_), .A2(new_n598_), .ZN(new_n5088_));
  OAI21_X1   g5039(.A1(new_n5087_), .A2(new_n5088_), .B(new_n5086_), .ZN(new_n5089_));
  OR3_X2     g5040(.A1(new_n5087_), .A2(new_n5086_), .A3(new_n5088_), .Z(new_n5090_));
  AND2_X2    g5041(.A1(new_n5090_), .A2(new_n5089_), .Z(new_n5091_));
  OAI22_X1   g5042(.A1(new_n2598_), .A2(new_n2815_), .B1(new_n2586_), .B2(new_n3001_), .ZN(new_n5092_));
  AOI21_X1   g5043(.A1(new_n2812_), .A2(new_n3859_), .B(new_n5092_), .ZN(new_n5093_));
  OAI21_X1   g5044(.A1(new_n4859_), .A2(new_n2820_), .B(new_n5093_), .ZN(new_n5094_));
  XOR2_X1    g5045(.A1(new_n5094_), .A2(new_n465_), .Z(new_n5095_));
  XOR2_X1    g5046(.A1(new_n5091_), .A2(new_n5095_), .Z(new_n5096_));
  NOR2_X1    g5047(.A1(new_n5029_), .A2(new_n5039_), .ZN(new_n5097_));
  NOR2_X1    g5048(.A1(new_n5097_), .A2(new_n5038_), .ZN(new_n5098_));
  AOI22_X1   g5049(.A1(new_n4001_), .A2(new_n2738_), .B1(new_n3868_), .B2(new_n2752_), .ZN(new_n5099_));
  OAI21_X1   g5050(.A1(new_n2736_), .A2(new_n4098_), .B(new_n5099_), .ZN(new_n5100_));
  NOR2_X1    g5051(.A1(new_n4852_), .A2(new_n2743_), .ZN(new_n5101_));
  NOR2_X1    g5052(.A1(new_n5101_), .A2(new_n5100_), .ZN(new_n5102_));
  XOR2_X1    g5053(.A1(new_n5102_), .A2(new_n474_), .Z(new_n5103_));
  NAND2_X1   g5054(.A1(new_n5098_), .A2(new_n5103_), .ZN(new_n5104_));
  NOR2_X1    g5055(.A1(new_n5098_), .A2(new_n5103_), .ZN(new_n5105_));
  INV_X1     g5056(.I(new_n5105_), .ZN(new_n5106_));
  NAND2_X1   g5057(.A1(new_n5106_), .A2(new_n5104_), .ZN(new_n5107_));
  XOR2_X1    g5058(.A1(new_n5107_), .A2(new_n5096_), .Z(new_n5108_));
  XOR2_X1    g5059(.A1(new_n5108_), .A2(new_n5081_), .Z(new_n5109_));
  OAI21_X1   g5060(.A1(new_n5051_), .A2(new_n5045_), .B(new_n5109_), .ZN(new_n5110_));
  OAI21_X1   g5061(.A1(new_n5053_), .A2(new_n4987_), .B(new_n5052_), .ZN(new_n5111_));
  INV_X1     g5062(.I(new_n5109_), .ZN(new_n5112_));
  NAND3_X1   g5063(.A1(new_n5111_), .A2(new_n5046_), .A3(new_n5112_), .ZN(new_n5113_));
  NAND3_X1   g5064(.A1(new_n5113_), .A2(new_n5110_), .A3(new_n5076_), .ZN(new_n5114_));
  INV_X1     g5065(.I(new_n5114_), .ZN(new_n5115_));
  AOI21_X1   g5066(.A1(new_n5113_), .A2(new_n5110_), .B(new_n5076_), .ZN(new_n5116_));
  NOR2_X1    g5067(.A1(new_n5115_), .A2(new_n5116_), .ZN(new_n5117_));
  NAND2_X1   g5068(.A1(new_n5117_), .A2(new_n5071_), .ZN(new_n5118_));
  AOI21_X1   g5069(.A1(new_n5014_), .A2(new_n5055_), .B(new_n5056_), .ZN(new_n5119_));
  INV_X1     g5070(.I(new_n5116_), .ZN(new_n5120_));
  NAND2_X1   g5071(.A1(new_n5120_), .A2(new_n5114_), .ZN(new_n5121_));
  NAND2_X1   g5072(.A1(new_n5121_), .A2(new_n5119_), .ZN(new_n5122_));
  NAND2_X1   g5073(.A1(new_n5122_), .A2(new_n5118_), .ZN(new_n5123_));
  XOR2_X1    g5074(.A1(new_n5123_), .A2(new_n5066_), .Z(new_n5124_));
  XOR2_X1    g5075(.A1(new_n5069_), .A2(new_n5124_), .Z(\sin[10] ));
  NAND3_X1   g5076(.A1(new_n5123_), .A2(new_n5008_), .A3(new_n5063_), .ZN(new_n5126_));
  NAND4_X1   g5077(.A1(new_n5065_), .A2(new_n5122_), .A3(new_n5118_), .A4(new_n5062_), .ZN(new_n5127_));
  NAND2_X1   g5078(.A1(new_n5126_), .A2(new_n5127_), .ZN(new_n5128_));
  AOI21_X1   g5079(.A1(new_n5128_), .A2(new_n5012_), .B(new_n4074_), .ZN(new_n5129_));
  INV_X1     g5080(.I(new_n5081_), .ZN(new_n5130_));
  INV_X1     g5081(.I(new_n5108_), .ZN(new_n5131_));
  OAI21_X1   g5082(.A1(new_n5051_), .A2(new_n5045_), .B(new_n5131_), .ZN(new_n5132_));
  NOR3_X1    g5083(.A1(new_n5051_), .A2(new_n5045_), .A3(new_n5131_), .ZN(new_n5133_));
  AOI21_X1   g5084(.A1(new_n5130_), .A2(new_n5132_), .B(new_n5133_), .ZN(new_n5134_));
  INV_X1     g5085(.I(new_n5096_), .ZN(new_n5135_));
  NAND2_X1   g5086(.A1(new_n5135_), .A2(new_n5104_), .ZN(new_n5136_));
  NAND2_X1   g5087(.A1(new_n5136_), .A2(new_n5106_), .ZN(new_n5137_));
  NAND2_X1   g5088(.A1(new_n5091_), .A2(new_n5095_), .ZN(new_n5138_));
  NAND2_X1   g5089(.A1(new_n5138_), .A2(new_n5089_), .ZN(new_n5139_));
  AOI22_X1   g5090(.A1(new_n4476_), .A2(new_n2738_), .B1(new_n2752_), .B2(new_n4001_), .ZN(new_n5140_));
  OAI21_X1   g5091(.A1(new_n4341_), .A2(new_n2743_), .B(new_n5140_), .ZN(new_n5141_));
  XOR2_X1    g5092(.A1(new_n5141_), .A2(new_n473_), .Z(new_n5142_));
  OAI22_X1   g5093(.A1(new_n3573_), .A2(new_n2815_), .B1(new_n2598_), .B2(new_n3001_), .ZN(new_n5143_));
  AOI21_X1   g5094(.A1(new_n3868_), .A2(new_n2812_), .B(new_n5143_), .ZN(new_n5144_));
  OAI21_X1   g5095(.A1(new_n3885_), .A2(new_n2820_), .B(new_n5144_), .ZN(new_n5145_));
  XOR2_X1    g5096(.A1(new_n5145_), .A2(new_n598_), .Z(new_n5146_));
  INV_X1     g5097(.I(new_n5084_), .ZN(new_n5147_));
  OAI21_X1   g5098(.A1(new_n5082_), .A2(new_n5083_), .B(new_n5147_), .ZN(new_n5148_));
  NOR2_X1    g5099(.A1(new_n2586_), .A2(new_n598_), .ZN(new_n5149_));
  XOR2_X1    g5100(.A1(new_n5148_), .A2(new_n5149_), .Z(new_n5150_));
  XNOR2_X1   g5101(.A1(new_n5146_), .A2(new_n5150_), .ZN(new_n5151_));
  XNOR2_X1   g5102(.A1(new_n5151_), .A2(new_n5142_), .ZN(new_n5152_));
  XOR2_X1    g5103(.A1(new_n5152_), .A2(new_n5139_), .Z(new_n5153_));
  XNOR2_X1   g5104(.A1(new_n5153_), .A2(new_n5137_), .ZN(new_n5154_));
  NOR4_X1    g5105(.A1(new_n399_), .A2(new_n698_), .A3(new_n1257_), .A4(new_n916_), .ZN(new_n5155_));
  NAND4_X1   g5106(.A1(new_n535_), .A2(new_n449_), .A3(new_n3990_), .A4(new_n5155_), .ZN(new_n5156_));
  INV_X1     g5107(.I(new_n5156_), .ZN(new_n5157_));
  XOR2_X1    g5108(.A1(new_n5154_), .A2(new_n5157_), .Z(new_n5158_));
  XNOR2_X1   g5109(.A1(new_n5134_), .A2(new_n5158_), .ZN(new_n5159_));
  OAI21_X1   g5110(.A1(new_n5119_), .A2(new_n5115_), .B(new_n5120_), .ZN(new_n5160_));
  NAND2_X1   g5111(.A1(new_n5160_), .A2(new_n5159_), .ZN(new_n5161_));
  INV_X1     g5112(.I(new_n5159_), .ZN(new_n5162_));
  AOI21_X1   g5113(.A1(new_n5071_), .A2(new_n5114_), .B(new_n5116_), .ZN(new_n5163_));
  NAND2_X1   g5114(.A1(new_n5162_), .A2(new_n5163_), .ZN(new_n5164_));
  NAND2_X1   g5115(.A1(new_n5164_), .A2(new_n5161_), .ZN(new_n5165_));
  XOR2_X1    g5116(.A1(new_n5165_), .A2(new_n5127_), .Z(new_n5166_));
  XNOR2_X1   g5117(.A1(new_n5166_), .A2(new_n5129_), .ZN(\sin[11] ));
  NAND3_X1   g5118(.A1(new_n5166_), .A2(new_n5012_), .A3(new_n5128_), .ZN(new_n5168_));
  NAND2_X1   g5119(.A1(new_n5168_), .A2(new_n4073_), .ZN(new_n5169_));
  INV_X1     g5120(.I(new_n5127_), .ZN(new_n5170_));
  NAND2_X1   g5121(.A1(new_n5165_), .A2(new_n5170_), .ZN(new_n5171_));
  NAND2_X1   g5122(.A1(new_n5134_), .A2(new_n5154_), .ZN(new_n5172_));
  AOI21_X1   g5123(.A1(new_n5111_), .A2(new_n5046_), .B(new_n5108_), .ZN(new_n5173_));
  NAND3_X1   g5124(.A1(new_n5111_), .A2(new_n5046_), .A3(new_n5108_), .ZN(new_n5174_));
  OAI21_X1   g5125(.A1(new_n5081_), .A2(new_n5173_), .B(new_n5174_), .ZN(new_n5175_));
  INV_X1     g5126(.I(new_n5154_), .ZN(new_n5176_));
  NAND2_X1   g5127(.A1(new_n5175_), .A2(new_n5176_), .ZN(new_n5177_));
  NAND2_X1   g5128(.A1(new_n5177_), .A2(new_n5172_), .ZN(new_n5178_));
  AOI21_X1   g5129(.A1(new_n5160_), .A2(new_n5156_), .B(new_n5178_), .ZN(new_n5179_));
  NOR2_X1    g5130(.A1(new_n5160_), .A2(new_n5156_), .ZN(new_n5180_));
  NOR2_X1    g5131(.A1(new_n5153_), .A2(new_n5137_), .ZN(new_n5181_));
  NOR2_X1    g5132(.A1(new_n5173_), .A2(new_n5081_), .ZN(new_n5182_));
  NAND2_X1   g5133(.A1(new_n5153_), .A2(new_n5137_), .ZN(new_n5183_));
  INV_X1     g5134(.I(new_n5183_), .ZN(new_n5184_));
  NOR3_X1    g5135(.A1(new_n5182_), .A2(new_n5133_), .A3(new_n5184_), .ZN(new_n5185_));
  NOR2_X1    g5136(.A1(new_n5139_), .A2(new_n5151_), .ZN(new_n5186_));
  AOI21_X1   g5137(.A1(new_n5139_), .A2(new_n5151_), .B(new_n5142_), .ZN(new_n5187_));
  NOR2_X1    g5138(.A1(new_n5187_), .A2(new_n5186_), .ZN(new_n5188_));
  OAI22_X1   g5139(.A1(new_n3869_), .A2(new_n2815_), .B1(new_n3001_), .B2(new_n3573_), .ZN(new_n5189_));
  AOI21_X1   g5140(.A1(new_n2812_), .A2(new_n4001_), .B(new_n5189_), .ZN(new_n5190_));
  NAND2_X1   g5141(.A1(new_n4459_), .A2(new_n2819_), .ZN(new_n5191_));
  NAND2_X1   g5142(.A1(new_n5191_), .A2(new_n5190_), .ZN(new_n5192_));
  XOR2_X1    g5143(.A1(new_n5192_), .A2(new_n465_), .Z(new_n5193_));
  XOR2_X1    g5144(.A1(new_n5193_), .A2(new_n474_), .Z(new_n5194_));
  OAI22_X1   g5145(.A1(new_n4477_), .A2(new_n2743_), .B1(new_n2768_), .B2(new_n4098_), .ZN(new_n5195_));
  INV_X1     g5146(.I(new_n5148_), .ZN(new_n5196_));
  INV_X1     g5147(.I(new_n5149_), .ZN(new_n5197_));
  OAI21_X1   g5148(.A1(new_n5148_), .A2(new_n5149_), .B(new_n5146_), .ZN(new_n5198_));
  OAI21_X1   g5149(.A1(new_n5196_), .A2(new_n5197_), .B(new_n5198_), .ZN(new_n5199_));
  NOR2_X1    g5150(.A1(new_n2719_), .A2(new_n598_), .ZN(new_n5200_));
  XOR2_X1    g5151(.A1(new_n5199_), .A2(new_n5200_), .Z(new_n5201_));
  XNOR2_X1   g5152(.A1(new_n5201_), .A2(new_n5195_), .ZN(new_n5202_));
  XOR2_X1    g5153(.A1(new_n5202_), .A2(new_n5194_), .Z(new_n5203_));
  NAND2_X1   g5154(.A1(new_n5203_), .A2(new_n5188_), .ZN(new_n5204_));
  INV_X1     g5155(.I(new_n5204_), .ZN(new_n5205_));
  NOR2_X1    g5156(.A1(new_n5203_), .A2(new_n5188_), .ZN(new_n5206_));
  NOR2_X1    g5157(.A1(new_n5205_), .A2(new_n5206_), .ZN(new_n5207_));
  INV_X1     g5158(.I(new_n5207_), .ZN(new_n5208_));
  NOR3_X1    g5159(.A1(new_n5185_), .A2(new_n5181_), .A3(new_n5208_), .ZN(new_n5209_));
  AOI21_X1   g5160(.A1(new_n5134_), .A2(new_n5183_), .B(new_n5181_), .ZN(new_n5210_));
  NOR2_X1    g5161(.A1(new_n5210_), .A2(new_n5207_), .ZN(new_n5211_));
  INV_X1     g5162(.I(new_n4361_), .ZN(new_n5212_));
  NAND2_X1   g5163(.A1(new_n889_), .A2(new_n899_), .ZN(new_n5213_));
  NOR4_X1    g5164(.A1(new_n5213_), .A2(new_n452_), .A3(new_n299_), .A4(new_n321_), .ZN(new_n5214_));
  NOR4_X1    g5165(.A1(new_n2399_), .A2(new_n156_), .A3(new_n177_), .A4(new_n187_), .ZN(new_n5215_));
  NAND4_X1   g5166(.A1(new_n5215_), .A2(new_n5212_), .A3(new_n897_), .A4(new_n5214_), .ZN(new_n5216_));
  NOR3_X1    g5167(.A1(new_n2257_), .A2(new_n2336_), .A3(new_n5216_), .ZN(new_n5217_));
  NOR3_X1    g5168(.A1(new_n5211_), .A2(new_n5209_), .A3(new_n5217_), .ZN(new_n5218_));
  NAND2_X1   g5169(.A1(new_n5210_), .A2(new_n5207_), .ZN(new_n5219_));
  OAI21_X1   g5170(.A1(new_n5185_), .A2(new_n5181_), .B(new_n5208_), .ZN(new_n5220_));
  INV_X1     g5171(.I(new_n5217_), .ZN(new_n5221_));
  AOI21_X1   g5172(.A1(new_n5220_), .A2(new_n5219_), .B(new_n5221_), .ZN(new_n5222_));
  OAI22_X1   g5173(.A1(new_n5179_), .A2(new_n5180_), .B1(new_n5222_), .B2(new_n5218_), .ZN(new_n5223_));
  NOR4_X1    g5174(.A1(new_n5179_), .A2(new_n5180_), .A3(new_n5218_), .A4(new_n5222_), .ZN(new_n5224_));
  INV_X1     g5175(.I(new_n5224_), .ZN(new_n5225_));
  NAND3_X1   g5176(.A1(new_n5171_), .A2(new_n5225_), .A3(new_n5223_), .ZN(new_n5226_));
  AOI21_X1   g5177(.A1(new_n5164_), .A2(new_n5161_), .B(new_n5127_), .ZN(new_n5227_));
  INV_X1     g5178(.I(new_n5223_), .ZN(new_n5228_));
  OAI21_X1   g5179(.A1(new_n5228_), .A2(new_n5224_), .B(new_n5227_), .ZN(new_n5229_));
  NAND2_X1   g5180(.A1(new_n5226_), .A2(new_n5229_), .ZN(new_n5230_));
  XOR2_X1    g5181(.A1(new_n5169_), .A2(new_n5230_), .Z(\sin[12] ));
  NOR2_X1    g5182(.A1(new_n5201_), .A2(new_n5193_), .ZN(new_n5232_));
  XOR2_X1    g5183(.A1(new_n5195_), .A2(new_n473_), .Z(new_n5233_));
  AOI21_X1   g5184(.A1(new_n5201_), .A2(new_n5193_), .B(new_n5233_), .ZN(new_n5234_));
  NOR2_X1    g5185(.A1(new_n5234_), .A2(new_n5232_), .ZN(new_n5235_));
  INV_X1     g5186(.I(new_n5235_), .ZN(new_n5236_));
  NOR2_X1    g5187(.A1(new_n2598_), .A2(new_n598_), .ZN(new_n5237_));
  INV_X1     g5188(.I(new_n5237_), .ZN(new_n5238_));
  OAI21_X1   g5189(.A1(new_n5197_), .A2(new_n5237_), .B(new_n5199_), .ZN(new_n5239_));
  OAI21_X1   g5190(.A1(new_n5149_), .A2(new_n5238_), .B(new_n5239_), .ZN(new_n5240_));
  AOI22_X1   g5191(.A1(new_n4001_), .A2(new_n2816_), .B1(new_n3868_), .B2(new_n3000_), .ZN(new_n5241_));
  OAI21_X1   g5192(.A1(new_n3003_), .A2(new_n4098_), .B(new_n5241_), .ZN(new_n5242_));
  NOR2_X1    g5193(.A1(new_n4852_), .A2(new_n2820_), .ZN(new_n5243_));
  NOR2_X1    g5194(.A1(new_n5243_), .A2(new_n5242_), .ZN(new_n5244_));
  XOR2_X1    g5195(.A1(new_n5244_), .A2(new_n598_), .Z(new_n5245_));
  NOR2_X1    g5196(.A1(new_n3585_), .A2(new_n598_), .ZN(new_n5246_));
  XOR2_X1    g5197(.A1(new_n5246_), .A2(new_n473_), .Z(new_n5247_));
  XNOR2_X1   g5198(.A1(new_n5245_), .A2(new_n5247_), .ZN(new_n5248_));
  XNOR2_X1   g5199(.A1(new_n5240_), .A2(new_n5248_), .ZN(new_n5249_));
  XOR2_X1    g5200(.A1(new_n5249_), .A2(new_n5236_), .Z(new_n5250_));
  OAI21_X1   g5201(.A1(new_n5210_), .A2(new_n5208_), .B(new_n5204_), .ZN(new_n5251_));
  XOR2_X1    g5202(.A1(new_n5251_), .A2(new_n5250_), .Z(new_n5252_));
  INV_X1     g5203(.I(new_n2281_), .ZN(new_n5253_));
  INV_X1     g5204(.I(new_n4217_), .ZN(new_n5254_));
  NOR4_X1    g5205(.A1(new_n5254_), .A2(new_n200_), .A3(new_n388_), .A4(new_n524_), .ZN(new_n5255_));
  NOR4_X1    g5206(.A1(new_n191_), .A2(new_n495_), .A3(new_n729_), .A4(new_n722_), .ZN(new_n5256_));
  NAND2_X1   g5207(.A1(new_n2317_), .A2(new_n5256_), .ZN(new_n5257_));
  NOR2_X1    g5208(.A1(new_n267_), .A2(new_n545_), .ZN(new_n5258_));
  NAND4_X1   g5209(.A1(new_n5258_), .A2(new_n293_), .A3(new_n1085_), .A4(new_n1261_), .ZN(new_n5259_));
  NOR4_X1    g5210(.A1(new_n1138_), .A2(new_n868_), .A3(new_n5257_), .A4(new_n5259_), .ZN(new_n5260_));
  NAND4_X1   g5211(.A1(new_n3729_), .A2(new_n5253_), .A3(new_n5255_), .A4(new_n5260_), .ZN(new_n5261_));
  INV_X1     g5212(.I(new_n5261_), .ZN(new_n5262_));
  NAND2_X1   g5213(.A1(new_n5252_), .A2(new_n5262_), .ZN(new_n5263_));
  INV_X1     g5214(.I(new_n5250_), .ZN(new_n5264_));
  XOR2_X1    g5215(.A1(new_n5251_), .A2(new_n5264_), .Z(new_n5265_));
  NAND2_X1   g5216(.A1(new_n5265_), .A2(new_n5261_), .ZN(new_n5266_));
  NAND2_X1   g5217(.A1(new_n5263_), .A2(new_n5266_), .ZN(new_n5267_));
  AOI21_X1   g5218(.A1(new_n5220_), .A2(new_n5219_), .B(new_n5217_), .ZN(new_n5268_));
  NOR3_X1    g5219(.A1(new_n5211_), .A2(new_n5209_), .A3(new_n5221_), .ZN(new_n5269_));
  NOR3_X1    g5220(.A1(new_n5179_), .A2(new_n5180_), .A3(new_n5269_), .ZN(new_n5270_));
  NOR2_X1    g5221(.A1(new_n5270_), .A2(new_n5268_), .ZN(new_n5271_));
  NAND2_X1   g5222(.A1(new_n5229_), .A2(new_n5271_), .ZN(new_n5272_));
  AOI21_X1   g5223(.A1(new_n5225_), .A2(new_n5223_), .B(new_n5171_), .ZN(new_n5273_));
  INV_X1     g5224(.I(new_n5268_), .ZN(new_n5274_));
  NOR3_X1    g5225(.A1(new_n5182_), .A2(new_n5133_), .A3(new_n5176_), .ZN(new_n5275_));
  NOR2_X1    g5226(.A1(new_n5134_), .A2(new_n5154_), .ZN(new_n5276_));
  NOR2_X1    g5227(.A1(new_n5276_), .A2(new_n5275_), .ZN(new_n5277_));
  OAI21_X1   g5228(.A1(new_n5163_), .A2(new_n5157_), .B(new_n5277_), .ZN(new_n5278_));
  NAND2_X1   g5229(.A1(new_n5163_), .A2(new_n5157_), .ZN(new_n5279_));
  NAND3_X1   g5230(.A1(new_n5220_), .A2(new_n5219_), .A3(new_n5217_), .ZN(new_n5280_));
  NAND3_X1   g5231(.A1(new_n5278_), .A2(new_n5279_), .A3(new_n5280_), .ZN(new_n5281_));
  NAND2_X1   g5232(.A1(new_n5281_), .A2(new_n5274_), .ZN(new_n5282_));
  NAND2_X1   g5233(.A1(new_n5273_), .A2(new_n5282_), .ZN(new_n5283_));
  NAND3_X1   g5234(.A1(new_n5283_), .A2(new_n5272_), .A3(new_n5267_), .ZN(new_n5284_));
  NAND2_X1   g5235(.A1(new_n5283_), .A2(new_n5272_), .ZN(new_n5285_));
  NAND3_X1   g5236(.A1(new_n5285_), .A2(new_n5263_), .A3(new_n5266_), .ZN(new_n5286_));
  NAND2_X1   g5237(.A1(new_n5286_), .A2(new_n5284_), .ZN(new_n5287_));
  AOI21_X1   g5238(.A1(new_n5226_), .A2(new_n5229_), .B(new_n5168_), .ZN(new_n5288_));
  NOR2_X1    g5239(.A1(new_n5288_), .A2(new_n4074_), .ZN(new_n5289_));
  XOR2_X1    g5240(.A1(new_n5287_), .A2(new_n5289_), .Z(\sin[13] ));
  NAND3_X1   g5241(.A1(new_n5286_), .A2(new_n5284_), .A3(new_n5288_), .ZN(new_n5291_));
  NAND2_X1   g5242(.A1(new_n5291_), .A2(new_n4073_), .ZN(new_n5292_));
  NAND3_X1   g5243(.A1(new_n5271_), .A2(new_n5263_), .A3(new_n5266_), .ZN(new_n5293_));
  NOR2_X1    g5244(.A1(new_n5265_), .A2(new_n5261_), .ZN(new_n5294_));
  NOR2_X1    g5245(.A1(new_n5252_), .A2(new_n5262_), .ZN(new_n5295_));
  OAI21_X1   g5246(.A1(new_n5294_), .A2(new_n5295_), .B(new_n5282_), .ZN(new_n5296_));
  NAND2_X1   g5247(.A1(new_n5296_), .A2(new_n5293_), .ZN(new_n5297_));
  NAND2_X1   g5248(.A1(new_n5297_), .A2(new_n5273_), .ZN(new_n5298_));
  XOR2_X1    g5249(.A1(new_n5250_), .A2(new_n5261_), .Z(new_n5299_));
  INV_X1     g5250(.I(new_n5299_), .ZN(new_n5300_));
  AOI21_X1   g5251(.A1(new_n2281_), .A2(new_n5250_), .B(new_n5300_), .ZN(new_n5301_));
  NAND2_X1   g5252(.A1(new_n5251_), .A2(new_n5301_), .ZN(new_n5302_));
  OAI21_X1   g5253(.A1(new_n5251_), .A2(new_n5299_), .B(new_n5302_), .ZN(new_n5303_));
  OAI21_X1   g5254(.A1(new_n5270_), .A2(new_n5268_), .B(new_n5303_), .ZN(new_n5304_));
  NAND2_X1   g5255(.A1(new_n5304_), .A2(new_n5266_), .ZN(new_n5305_));
  AOI21_X1   g5256(.A1(new_n5251_), .A2(new_n5235_), .B(new_n5249_), .ZN(new_n5306_));
  NOR2_X1    g5257(.A1(new_n5251_), .A2(new_n5235_), .ZN(new_n5307_));
  INV_X1     g5258(.I(new_n5245_), .ZN(new_n5308_));
  NAND2_X1   g5259(.A1(new_n5308_), .A2(new_n5247_), .ZN(new_n5309_));
  OAI21_X1   g5260(.A1(new_n5308_), .A2(new_n5247_), .B(new_n5240_), .ZN(new_n5310_));
  NAND2_X1   g5261(.A1(new_n5310_), .A2(new_n5309_), .ZN(new_n5311_));
  AOI22_X1   g5262(.A1(new_n4476_), .A2(new_n2816_), .B1(new_n3000_), .B2(new_n4001_), .ZN(new_n5312_));
  OAI21_X1   g5263(.A1(new_n4341_), .A2(new_n2820_), .B(new_n5312_), .ZN(new_n5313_));
  XOR2_X1    g5264(.A1(new_n5313_), .A2(new_n598_), .Z(new_n5314_));
  NAND2_X1   g5265(.A1(new_n3582_), .A2(new_n474_), .ZN(new_n5315_));
  AOI21_X1   g5266(.A1(new_n5315_), .A2(new_n3579_), .B(new_n598_), .ZN(new_n5316_));
  NOR3_X1    g5267(.A1(new_n5316_), .A2(new_n598_), .A3(new_n3869_), .ZN(new_n5317_));
  OAI21_X1   g5268(.A1(new_n598_), .A2(new_n3869_), .B(new_n5316_), .ZN(new_n5318_));
  INV_X1     g5269(.I(new_n5318_), .ZN(new_n5319_));
  NOR2_X1    g5270(.A1(new_n5319_), .A2(new_n5317_), .ZN(new_n5320_));
  XOR2_X1    g5271(.A1(new_n5314_), .A2(new_n5320_), .Z(new_n5321_));
  NOR2_X1    g5272(.A1(new_n5311_), .A2(new_n5321_), .ZN(new_n5322_));
  NAND2_X1   g5273(.A1(new_n5311_), .A2(new_n5321_), .ZN(new_n5323_));
  INV_X1     g5274(.I(new_n5323_), .ZN(new_n5324_));
  NOR2_X1    g5275(.A1(new_n5324_), .A2(new_n5322_), .ZN(new_n5325_));
  NOR3_X1    g5276(.A1(new_n5306_), .A2(new_n5307_), .A3(new_n5325_), .ZN(new_n5326_));
  INV_X1     g5277(.I(new_n5326_), .ZN(new_n5327_));
  OAI21_X1   g5278(.A1(new_n5306_), .A2(new_n5307_), .B(new_n5325_), .ZN(new_n5328_));
  NAND4_X1   g5279(.A1(new_n2398_), .A2(new_n380_), .A3(new_n2461_), .A4(new_n3563_), .ZN(new_n5329_));
  NOR4_X1    g5280(.A1(new_n353_), .A2(new_n339_), .A3(new_n698_), .A4(new_n269_), .ZN(new_n5330_));
  NAND4_X1   g5281(.A1(new_n5330_), .A2(new_n1079_), .A3(new_n408_), .A4(new_n439_), .ZN(new_n5331_));
  NOR3_X1    g5282(.A1(new_n5329_), .A2(new_n5331_), .A3(new_n1074_), .ZN(new_n5332_));
  INV_X1     g5283(.I(new_n5332_), .ZN(new_n5333_));
  NOR4_X1    g5284(.A1(new_n2287_), .A2(new_n859_), .A3(new_n1439_), .A4(new_n5333_), .ZN(new_n5334_));
  INV_X1     g5285(.I(new_n5334_), .ZN(new_n5335_));
  NAND3_X1   g5286(.A1(new_n5327_), .A2(new_n5328_), .A3(new_n5335_), .ZN(new_n5336_));
  INV_X1     g5287(.I(new_n5328_), .ZN(new_n5337_));
  OAI21_X1   g5288(.A1(new_n5337_), .A2(new_n5326_), .B(new_n5334_), .ZN(new_n5338_));
  NAND3_X1   g5289(.A1(new_n5305_), .A2(new_n5338_), .A3(new_n5336_), .ZN(new_n5339_));
  OAI21_X1   g5290(.A1(new_n5185_), .A2(new_n5181_), .B(new_n5207_), .ZN(new_n5340_));
  INV_X1     g5291(.I(new_n5301_), .ZN(new_n5341_));
  AOI21_X1   g5292(.A1(new_n5340_), .A2(new_n5204_), .B(new_n5341_), .ZN(new_n5342_));
  NOR2_X1    g5293(.A1(new_n5251_), .A2(new_n5299_), .ZN(new_n5343_));
  NOR2_X1    g5294(.A1(new_n5343_), .A2(new_n5342_), .ZN(new_n5344_));
  AOI21_X1   g5295(.A1(new_n5281_), .A2(new_n5274_), .B(new_n5344_), .ZN(new_n5345_));
  NOR2_X1    g5296(.A1(new_n5345_), .A2(new_n5295_), .ZN(new_n5346_));
  NOR3_X1    g5297(.A1(new_n5337_), .A2(new_n5326_), .A3(new_n5334_), .ZN(new_n5347_));
  AOI21_X1   g5298(.A1(new_n5327_), .A2(new_n5328_), .B(new_n5335_), .ZN(new_n5348_));
  OAI21_X1   g5299(.A1(new_n5347_), .A2(new_n5348_), .B(new_n5346_), .ZN(new_n5349_));
  NAND2_X1   g5300(.A1(new_n5349_), .A2(new_n5339_), .ZN(new_n5350_));
  NOR2_X1    g5301(.A1(new_n5350_), .A2(new_n5298_), .ZN(new_n5351_));
  AOI21_X1   g5302(.A1(new_n5293_), .A2(new_n5296_), .B(new_n5229_), .ZN(new_n5352_));
  AOI21_X1   g5303(.A1(new_n5339_), .A2(new_n5349_), .B(new_n5352_), .ZN(new_n5353_));
  NAND4_X1   g5304(.A1(new_n5346_), .A2(new_n5338_), .A3(new_n5336_), .A4(new_n5171_), .ZN(new_n5354_));
  OAI21_X1   g5305(.A1(new_n5351_), .A2(new_n5353_), .B(new_n5354_), .ZN(new_n5355_));
  XOR2_X1    g5306(.A1(new_n5292_), .A2(new_n5355_), .Z(\sin[14] ));
  NAND4_X1   g5307(.A1(new_n5355_), .A2(new_n5284_), .A3(new_n5286_), .A4(new_n5288_), .ZN(new_n5357_));
  NAND2_X1   g5308(.A1(new_n5357_), .A2(new_n4073_), .ZN(new_n5358_));
  NOR2_X1    g5309(.A1(new_n5337_), .A2(new_n5326_), .ZN(new_n5359_));
  OAI21_X1   g5310(.A1(new_n5345_), .A2(new_n5295_), .B(new_n5335_), .ZN(new_n5360_));
  NOR3_X1    g5311(.A1(new_n5345_), .A2(new_n5295_), .A3(new_n5335_), .ZN(new_n5361_));
  AOI21_X1   g5312(.A1(new_n5359_), .A2(new_n5360_), .B(new_n5361_), .ZN(new_n5362_));
  NOR4_X1    g5313(.A1(new_n2464_), .A2(new_n2263_), .A3(new_n269_), .A4(new_n377_), .ZN(new_n5363_));
  NOR4_X1    g5314(.A1(new_n736_), .A2(new_n327_), .A3(new_n745_), .A4(new_n381_), .ZN(new_n5364_));
  NAND4_X1   g5315(.A1(new_n5363_), .A2(new_n1067_), .A3(new_n5214_), .A4(new_n5364_), .ZN(new_n5365_));
  NOR4_X1    g5316(.A1(new_n1274_), .A2(new_n207_), .A3(new_n265_), .A4(new_n272_), .ZN(new_n5366_));
  INV_X1     g5317(.I(new_n5366_), .ZN(new_n5367_));
  NOR3_X1    g5318(.A1(new_n5367_), .A2(new_n2401_), .A3(new_n5365_), .ZN(new_n5368_));
  INV_X1     g5319(.I(new_n5368_), .ZN(new_n5369_));
  AOI22_X1   g5320(.A1(new_n4743_), .A2(new_n2819_), .B1(new_n3000_), .B2(new_n4476_), .ZN(new_n5370_));
  NOR2_X1    g5321(.A1(new_n4002_), .A2(new_n3868_), .ZN(new_n5371_));
  NOR2_X1    g5322(.A1(new_n3869_), .A2(new_n4001_), .ZN(new_n5372_));
  OR3_X2     g5323(.A1(new_n5371_), .A2(new_n598_), .A3(new_n5372_), .Z(new_n5373_));
  XNOR2_X1   g5324(.A1(new_n5370_), .A2(new_n5373_), .ZN(new_n5374_));
  INV_X1     g5325(.I(new_n5374_), .ZN(new_n5375_));
  AOI21_X1   g5326(.A1(new_n5314_), .A2(new_n5318_), .B(new_n5317_), .ZN(new_n5376_));
  XOR2_X1    g5327(.A1(new_n5376_), .A2(new_n5375_), .Z(new_n5377_));
  INV_X1     g5328(.I(new_n5377_), .ZN(new_n5378_));
  NOR3_X1    g5329(.A1(new_n5306_), .A2(new_n5307_), .A3(new_n5324_), .ZN(new_n5379_));
  OAI21_X1   g5330(.A1(new_n5379_), .A2(new_n5322_), .B(new_n5378_), .ZN(new_n5380_));
  INV_X1     g5331(.I(new_n5322_), .ZN(new_n5381_));
  INV_X1     g5332(.I(new_n5249_), .ZN(new_n5382_));
  INV_X1     g5333(.I(new_n5181_), .ZN(new_n5383_));
  OAI21_X1   g5334(.A1(new_n5175_), .A2(new_n5184_), .B(new_n5383_), .ZN(new_n5384_));
  AOI21_X1   g5335(.A1(new_n5384_), .A2(new_n5207_), .B(new_n5205_), .ZN(new_n5385_));
  OAI21_X1   g5336(.A1(new_n5385_), .A2(new_n5236_), .B(new_n5382_), .ZN(new_n5386_));
  NAND2_X1   g5337(.A1(new_n5385_), .A2(new_n5236_), .ZN(new_n5387_));
  NAND3_X1   g5338(.A1(new_n5386_), .A2(new_n5387_), .A3(new_n5323_), .ZN(new_n5388_));
  NAND3_X1   g5339(.A1(new_n5388_), .A2(new_n5381_), .A3(new_n5377_), .ZN(new_n5389_));
  AOI21_X1   g5340(.A1(new_n5389_), .A2(new_n5380_), .B(new_n5369_), .ZN(new_n5390_));
  AOI21_X1   g5341(.A1(new_n5388_), .A2(new_n5381_), .B(new_n5377_), .ZN(new_n5391_));
  NOR3_X1    g5342(.A1(new_n5379_), .A2(new_n5322_), .A3(new_n5378_), .ZN(new_n5392_));
  NOR3_X1    g5343(.A1(new_n5391_), .A2(new_n5392_), .A3(new_n5368_), .ZN(new_n5393_));
  NOR2_X1    g5344(.A1(new_n5390_), .A2(new_n5393_), .ZN(new_n5394_));
  NAND2_X1   g5345(.A1(new_n5362_), .A2(new_n5394_), .ZN(new_n5395_));
  INV_X1     g5346(.I(new_n5359_), .ZN(new_n5396_));
  AOI21_X1   g5347(.A1(new_n5304_), .A2(new_n5266_), .B(new_n5334_), .ZN(new_n5397_));
  NAND3_X1   g5348(.A1(new_n5304_), .A2(new_n5266_), .A3(new_n5334_), .ZN(new_n5398_));
  OAI21_X1   g5349(.A1(new_n5396_), .A2(new_n5397_), .B(new_n5398_), .ZN(new_n5399_));
  OAI21_X1   g5350(.A1(new_n5391_), .A2(new_n5392_), .B(new_n5368_), .ZN(new_n5400_));
  NAND3_X1   g5351(.A1(new_n5389_), .A2(new_n5380_), .A3(new_n5369_), .ZN(new_n5401_));
  NAND2_X1   g5352(.A1(new_n5400_), .A2(new_n5401_), .ZN(new_n5402_));
  NAND2_X1   g5353(.A1(new_n5399_), .A2(new_n5402_), .ZN(new_n5403_));
  NAND4_X1   g5354(.A1(new_n5403_), .A2(new_n5395_), .A3(new_n5350_), .A4(new_n5352_), .ZN(new_n5404_));
  NOR3_X1    g5355(.A1(new_n5346_), .A2(new_n5347_), .A3(new_n5348_), .ZN(new_n5405_));
  AOI21_X1   g5356(.A1(new_n5336_), .A2(new_n5338_), .B(new_n5305_), .ZN(new_n5406_));
  OAI21_X1   g5357(.A1(new_n5405_), .A2(new_n5406_), .B(new_n5352_), .ZN(new_n5407_));
  NOR2_X1    g5358(.A1(new_n5399_), .A2(new_n5402_), .ZN(new_n5408_));
  NOR2_X1    g5359(.A1(new_n5362_), .A2(new_n5394_), .ZN(new_n5409_));
  OAI21_X1   g5360(.A1(new_n5408_), .A2(new_n5409_), .B(new_n5407_), .ZN(new_n5410_));
  NAND2_X1   g5361(.A1(new_n5410_), .A2(new_n5404_), .ZN(new_n5411_));
  XOR2_X1    g5362(.A1(new_n5358_), .A2(new_n5411_), .Z(\sin[15] ));
  INV_X1     g5363(.I(new_n5355_), .ZN(new_n5413_));
  NOR2_X1    g5364(.A1(new_n5413_), .A2(new_n5291_), .ZN(new_n5414_));
  NAND2_X1   g5365(.A1(new_n5414_), .A2(new_n5411_), .ZN(new_n5415_));
  NAND2_X1   g5366(.A1(new_n5415_), .A2(new_n4073_), .ZN(new_n5416_));
  NOR3_X1    g5367(.A1(new_n5407_), .A2(new_n5408_), .A3(new_n5409_), .ZN(new_n5417_));
  AOI21_X1   g5368(.A1(new_n5399_), .A2(new_n5401_), .B(new_n5390_), .ZN(new_n5418_));
  AND2_X2    g5369(.A1(new_n5370_), .A2(new_n598_), .Z(new_n5419_));
  INV_X1     g5370(.I(new_n5372_), .ZN(new_n5420_));
  AOI21_X1   g5371(.A1(new_n5370_), .A2(new_n5420_), .B(new_n5371_), .ZN(new_n5421_));
  AOI21_X1   g5372(.A1(new_n5421_), .A2(new_n465_), .B(new_n5419_), .ZN(new_n5422_));
  INV_X1     g5373(.I(new_n5422_), .ZN(new_n5423_));
  NAND2_X1   g5374(.A1(new_n5376_), .A2(new_n5374_), .ZN(new_n5424_));
  AOI21_X1   g5375(.A1(new_n5380_), .A2(new_n5424_), .B(new_n5423_), .ZN(new_n5425_));
  INV_X1     g5376(.I(new_n5424_), .ZN(new_n5426_));
  NOR3_X1    g5377(.A1(new_n5391_), .A2(new_n5422_), .A3(new_n5426_), .ZN(new_n5427_));
  NOR2_X1    g5378(.A1(new_n4098_), .A2(new_n3868_), .ZN(new_n5428_));
  NOR2_X1    g5379(.A1(new_n4476_), .A2(new_n3869_), .ZN(new_n5429_));
  NOR3_X1    g5380(.A1(new_n5429_), .A2(new_n598_), .A3(new_n5428_), .ZN(new_n5430_));
  NOR3_X1    g5381(.A1(new_n5427_), .A2(new_n5425_), .A3(new_n5430_), .ZN(new_n5431_));
  OAI21_X1   g5382(.A1(new_n5391_), .A2(new_n5426_), .B(new_n5422_), .ZN(new_n5432_));
  NAND3_X1   g5383(.A1(new_n5380_), .A2(new_n5423_), .A3(new_n5424_), .ZN(new_n5433_));
  INV_X1     g5384(.I(new_n5430_), .ZN(new_n5434_));
  AOI21_X1   g5385(.A1(new_n5432_), .A2(new_n5433_), .B(new_n5434_), .ZN(new_n5435_));
  INV_X1     g5386(.I(new_n2320_), .ZN(new_n5436_));
  NOR2_X1    g5387(.A1(new_n854_), .A2(new_n312_), .ZN(new_n5437_));
  NAND4_X1   g5388(.A1(new_n5437_), .A2(new_n424_), .A3(new_n498_), .A4(new_n481_), .ZN(new_n5438_));
  NOR4_X1    g5389(.A1(new_n5438_), .A2(new_n5436_), .A3(new_n5259_), .A4(new_n3763_), .ZN(new_n5439_));
  NAND3_X1   g5390(.A1(new_n2364_), .A2(new_n3726_), .A3(new_n5439_), .ZN(new_n5440_));
  INV_X1     g5391(.I(new_n5440_), .ZN(new_n5441_));
  OAI21_X1   g5392(.A1(new_n5431_), .A2(new_n5435_), .B(new_n5441_), .ZN(new_n5442_));
  NAND3_X1   g5393(.A1(new_n5432_), .A2(new_n5433_), .A3(new_n5434_), .ZN(new_n5443_));
  OAI21_X1   g5394(.A1(new_n5427_), .A2(new_n5425_), .B(new_n5430_), .ZN(new_n5444_));
  NAND3_X1   g5395(.A1(new_n5444_), .A2(new_n5443_), .A3(new_n5440_), .ZN(new_n5445_));
  NAND3_X1   g5396(.A1(new_n5418_), .A2(new_n5442_), .A3(new_n5445_), .ZN(new_n5446_));
  OAI21_X1   g5397(.A1(new_n5362_), .A2(new_n5393_), .B(new_n5400_), .ZN(new_n5447_));
  AOI21_X1   g5398(.A1(new_n5444_), .A2(new_n5443_), .B(new_n5440_), .ZN(new_n5448_));
  NOR3_X1    g5399(.A1(new_n5431_), .A2(new_n5435_), .A3(new_n5441_), .ZN(new_n5449_));
  OAI21_X1   g5400(.A1(new_n5449_), .A2(new_n5448_), .B(new_n5447_), .ZN(new_n5450_));
  NAND3_X1   g5401(.A1(new_n5417_), .A2(new_n5450_), .A3(new_n5446_), .ZN(new_n5451_));
  NOR3_X1    g5402(.A1(new_n5447_), .A2(new_n5449_), .A3(new_n5448_), .ZN(new_n5452_));
  AOI21_X1   g5403(.A1(new_n5442_), .A2(new_n5445_), .B(new_n5418_), .ZN(new_n5453_));
  OAI21_X1   g5404(.A1(new_n5453_), .A2(new_n5452_), .B(new_n5404_), .ZN(new_n5454_));
  NAND2_X1   g5405(.A1(new_n5454_), .A2(new_n5451_), .ZN(new_n5455_));
  XOR2_X1    g5406(.A1(new_n5416_), .A2(new_n5455_), .Z(\sin[16] ));
  NOR2_X1    g5407(.A1(new_n906_), .A2(new_n868_), .ZN(new_n5457_));
  NOR4_X1    g5408(.A1(new_n691_), .A2(new_n177_), .A3(new_n321_), .A4(new_n722_), .ZN(new_n5458_));
  NOR3_X1    g5409(.A1(new_n185_), .A2(new_n139_), .A3(new_n695_), .ZN(new_n5459_));
  NAND4_X1   g5410(.A1(new_n5458_), .A2(new_n712_), .A3(new_n5459_), .A4(new_n5457_), .ZN(new_n5460_));
  INV_X1     g5411(.I(new_n5460_), .ZN(new_n5461_));
  NAND4_X1   g5412(.A1(new_n2581_), .A2(new_n568_), .A3(new_n591_), .A4(new_n5461_), .ZN(new_n5462_));
  INV_X1     g5413(.I(new_n5462_), .ZN(new_n5463_));
  OAI21_X1   g5414(.A1(new_n5447_), .A2(new_n5448_), .B(new_n5445_), .ZN(new_n5464_));
  NOR2_X1    g5415(.A1(new_n5464_), .A2(new_n5463_), .ZN(new_n5465_));
  AOI21_X1   g5416(.A1(new_n5418_), .A2(new_n5442_), .B(new_n5449_), .ZN(new_n5466_));
  NOR2_X1    g5417(.A1(new_n5466_), .A2(new_n5462_), .ZN(new_n5467_));
  NOR2_X1    g5418(.A1(new_n5467_), .A2(new_n5465_), .ZN(new_n5468_));
  NAND2_X1   g5419(.A1(new_n5468_), .A2(new_n5451_), .ZN(new_n5469_));
  NOR3_X1    g5420(.A1(new_n5453_), .A2(new_n5452_), .A3(new_n5404_), .ZN(new_n5470_));
  NAND2_X1   g5421(.A1(new_n5466_), .A2(new_n5462_), .ZN(new_n5471_));
  NAND2_X1   g5422(.A1(new_n5464_), .A2(new_n5463_), .ZN(new_n5472_));
  NAND2_X1   g5423(.A1(new_n5471_), .A2(new_n5472_), .ZN(new_n5473_));
  NAND2_X1   g5424(.A1(new_n5473_), .A2(new_n5470_), .ZN(new_n5474_));
  NAND2_X1   g5425(.A1(new_n5469_), .A2(new_n5474_), .ZN(new_n5475_));
  INV_X1     g5426(.I(new_n5411_), .ZN(new_n5476_));
  NOR2_X1    g5427(.A1(new_n5476_), .A2(new_n5357_), .ZN(new_n5477_));
  AOI21_X1   g5428(.A1(new_n5477_), .A2(new_n5455_), .B(new_n4074_), .ZN(new_n5478_));
  XNOR2_X1   g5429(.A1(new_n5478_), .A2(new_n5475_), .ZN(\sin[17] ));
  AOI21_X1   g5430(.A1(new_n5471_), .A2(new_n5472_), .B(new_n5451_), .ZN(new_n5480_));
  NOR2_X1    g5431(.A1(new_n5473_), .A2(new_n5454_), .ZN(new_n5481_));
  OAI21_X1   g5432(.A1(new_n5481_), .A2(new_n5480_), .B(new_n5477_), .ZN(new_n5482_));
  NAND2_X1   g5433(.A1(new_n5482_), .A2(new_n4073_), .ZN(new_n5483_));
  INV_X1     g5434(.I(new_n572_), .ZN(new_n5484_));
  NAND3_X1   g5435(.A1(new_n438_), .A2(new_n877_), .A3(new_n740_), .ZN(new_n5485_));
  NOR4_X1    g5436(.A1(new_n974_), .A2(new_n5485_), .A3(new_n321_), .A4(new_n339_), .ZN(new_n5486_));
  NAND4_X1   g5437(.A1(new_n5486_), .A2(new_n507_), .A3(new_n2279_), .A4(new_n1149_), .ZN(new_n5487_));
  NOR4_X1    g5438(.A1(new_n3736_), .A2(new_n5484_), .A3(new_n1117_), .A4(new_n5487_), .ZN(new_n5488_));
  INV_X1     g5439(.I(new_n5488_), .ZN(new_n5489_));
  AOI21_X1   g5440(.A1(new_n5464_), .A2(new_n5462_), .B(new_n5489_), .ZN(new_n5490_));
  OAI21_X1   g5441(.A1(new_n5468_), .A2(new_n5451_), .B(new_n5490_), .ZN(new_n5491_));
  NAND3_X1   g5442(.A1(new_n5464_), .A2(new_n5462_), .A3(new_n5489_), .ZN(new_n5492_));
  INV_X1     g5443(.I(new_n5490_), .ZN(new_n5493_));
  NAND3_X1   g5444(.A1(new_n5473_), .A2(new_n5493_), .A3(new_n5470_), .ZN(new_n5494_));
  NAND3_X1   g5445(.A1(new_n5491_), .A2(new_n5494_), .A3(new_n5492_), .ZN(new_n5495_));
  XOR2_X1    g5446(.A1(new_n5483_), .A2(new_n5495_), .Z(\sin[18] ));
  NOR4_X1    g5447(.A1(new_n2290_), .A2(new_n263_), .A3(new_n2272_), .A4(new_n450_), .ZN(new_n5497_));
  NOR4_X1    g5448(.A1(new_n4700_), .A2(new_n312_), .A3(new_n402_), .A4(new_n549_), .ZN(new_n5498_));
  NAND4_X1   g5449(.A1(new_n5498_), .A2(new_n169_), .A3(new_n526_), .A4(new_n5497_), .ZN(new_n5499_));
  NOR3_X1    g5450(.A1(new_n5367_), .A2(new_n928_), .A3(new_n5499_), .ZN(new_n5500_));
  INV_X1     g5451(.I(new_n5500_), .ZN(new_n5501_));
  NAND2_X1   g5452(.A1(new_n5492_), .A2(new_n5501_), .ZN(new_n5502_));
  NAND4_X1   g5453(.A1(new_n5464_), .A2(new_n5462_), .A3(new_n5489_), .A4(new_n5500_), .ZN(new_n5503_));
  NAND2_X1   g5454(.A1(new_n5502_), .A2(new_n5503_), .ZN(new_n5504_));
  NAND2_X1   g5455(.A1(new_n5494_), .A2(new_n5504_), .ZN(new_n5505_));
  NAND4_X1   g5456(.A1(new_n5480_), .A2(new_n5493_), .A3(new_n5502_), .A4(new_n5503_), .ZN(new_n5506_));
  NAND2_X1   g5457(.A1(new_n5506_), .A2(new_n5505_), .ZN(new_n5507_));
  OR3_X2     g5458(.A1(new_n5454_), .A2(new_n5465_), .A3(new_n5467_), .Z(new_n5508_));
  AOI21_X1   g5459(.A1(new_n5508_), .A2(new_n5474_), .B(new_n5415_), .ZN(new_n5509_));
  AOI21_X1   g5460(.A1(new_n5509_), .A2(new_n5495_), .B(new_n4074_), .ZN(new_n5510_));
  XOR2_X1    g5461(.A1(new_n5510_), .A2(new_n5507_), .Z(\sin[19] ));
  NOR4_X1    g5462(.A1(new_n2356_), .A2(new_n544_), .A3(new_n201_), .A4(new_n400_), .ZN(new_n5512_));
  NOR2_X1    g5463(.A1(new_n2436_), .A2(new_n492_), .ZN(new_n5513_));
  NAND4_X1   g5464(.A1(new_n5513_), .A2(new_n342_), .A3(new_n406_), .A4(new_n5512_), .ZN(new_n5514_));
  NOR2_X1    g5465(.A1(new_n5514_), .A2(new_n2253_), .ZN(new_n5515_));
  NOR2_X1    g5466(.A1(new_n4945_), .A2(new_n456_), .ZN(new_n5516_));
  NAND3_X1   g5467(.A1(new_n5516_), .A2(new_n982_), .A3(new_n5515_), .ZN(new_n5517_));
  INV_X1     g5468(.I(new_n5517_), .ZN(new_n5518_));
  NAND4_X1   g5469(.A1(new_n5464_), .A2(new_n5462_), .A3(new_n5489_), .A4(new_n5501_), .ZN(new_n5519_));
  NAND2_X1   g5470(.A1(new_n5519_), .A2(new_n5518_), .ZN(new_n5520_));
  NOR4_X1    g5471(.A1(new_n5466_), .A2(new_n5463_), .A3(new_n5488_), .A4(new_n5500_), .ZN(new_n5521_));
  NAND2_X1   g5472(.A1(new_n5521_), .A2(new_n5517_), .ZN(new_n5522_));
  AND2_X2    g5473(.A1(new_n5522_), .A2(new_n5520_), .Z(new_n5523_));
  NOR3_X1    g5474(.A1(new_n5466_), .A2(new_n5463_), .A3(new_n5488_), .ZN(new_n5524_));
  NOR2_X1    g5475(.A1(new_n5524_), .A2(new_n5500_), .ZN(new_n5525_));
  INV_X1     g5476(.I(new_n5503_), .ZN(new_n5526_));
  NOR2_X1    g5477(.A1(new_n5525_), .A2(new_n5526_), .ZN(new_n5527_));
  NOR2_X1    g5478(.A1(new_n5527_), .A2(new_n5494_), .ZN(new_n5528_));
  NAND4_X1   g5479(.A1(new_n5504_), .A2(new_n5480_), .A3(new_n5493_), .A4(new_n5520_), .ZN(new_n5529_));
  OAI21_X1   g5480(.A1(new_n5523_), .A2(new_n5528_), .B(new_n5529_), .ZN(new_n5530_));
  NAND4_X1   g5481(.A1(new_n5509_), .A2(new_n5495_), .A3(new_n5505_), .A4(new_n5506_), .ZN(new_n5531_));
  NAND2_X1   g5482(.A1(new_n5531_), .A2(new_n4073_), .ZN(new_n5532_));
  XOR2_X1    g5483(.A1(new_n5532_), .A2(new_n5530_), .Z(\sin[20] ));
  NOR3_X1    g5484(.A1(new_n5468_), .A2(new_n5451_), .A3(new_n5490_), .ZN(new_n5534_));
  AOI22_X1   g5485(.A1(new_n5534_), .A2(new_n5504_), .B1(new_n5520_), .B2(new_n5522_), .ZN(new_n5535_));
  INV_X1     g5486(.I(new_n5520_), .ZN(new_n5536_));
  NOR3_X1    g5487(.A1(new_n5527_), .A2(new_n5494_), .A3(new_n5536_), .ZN(new_n5537_));
  NOR2_X1    g5488(.A1(new_n5535_), .A2(new_n5537_), .ZN(new_n5538_));
  NOR2_X1    g5489(.A1(new_n5531_), .A2(new_n5538_), .ZN(new_n5539_));
  NOR2_X1    g5490(.A1(new_n5539_), .A2(new_n4074_), .ZN(new_n5540_));
  NAND4_X1   g5491(.A1(new_n469_), .A2(new_n391_), .A3(new_n2347_), .A4(new_n3863_), .ZN(new_n5541_));
  INV_X1     g5492(.I(new_n5541_), .ZN(new_n5542_));
  NOR3_X1    g5493(.A1(new_n5519_), .A2(new_n5518_), .A3(new_n5542_), .ZN(new_n5543_));
  AOI21_X1   g5494(.A1(new_n5521_), .A2(new_n5517_), .B(new_n5541_), .ZN(new_n5544_));
  NOR2_X1    g5495(.A1(new_n5544_), .A2(new_n5543_), .ZN(new_n5545_));
  NAND4_X1   g5496(.A1(new_n5545_), .A2(new_n5534_), .A3(new_n5504_), .A4(new_n5520_), .ZN(new_n5546_));
  NAND3_X1   g5497(.A1(new_n5521_), .A2(new_n5517_), .A3(new_n5541_), .ZN(new_n5547_));
  OAI21_X1   g5498(.A1(new_n5519_), .A2(new_n5518_), .B(new_n5542_), .ZN(new_n5548_));
  NAND2_X1   g5499(.A1(new_n5547_), .A2(new_n5548_), .ZN(new_n5549_));
  NAND2_X1   g5500(.A1(new_n5529_), .A2(new_n5549_), .ZN(new_n5550_));
  NAND2_X1   g5501(.A1(new_n5550_), .A2(new_n5546_), .ZN(new_n5551_));
  XNOR2_X1   g5502(.A1(new_n5540_), .A2(new_n5551_), .ZN(\sin[21] ));
  AOI21_X1   g5503(.A1(new_n5473_), .A2(new_n5470_), .B(new_n5493_), .ZN(new_n5553_));
  NOR3_X1    g5504(.A1(new_n5553_), .A2(new_n5534_), .A3(new_n5524_), .ZN(new_n5554_));
  NOR2_X1    g5505(.A1(new_n5534_), .A2(new_n5527_), .ZN(new_n5555_));
  NOR2_X1    g5506(.A1(new_n5494_), .A2(new_n5504_), .ZN(new_n5556_));
  NOR4_X1    g5507(.A1(new_n5482_), .A2(new_n5554_), .A3(new_n5555_), .A4(new_n5556_), .ZN(new_n5557_));
  NAND3_X1   g5508(.A1(new_n5551_), .A2(new_n5557_), .A3(new_n5530_), .ZN(new_n5558_));
  NAND2_X1   g5509(.A1(new_n5558_), .A2(new_n4073_), .ZN(new_n5559_));
  NOR4_X1    g5510(.A1(new_n5549_), .A2(new_n5494_), .A3(new_n5527_), .A4(new_n5536_), .ZN(new_n5560_));
  NAND2_X1   g5511(.A1(new_n469_), .A2(new_n442_), .ZN(new_n5561_));
  NAND2_X1   g5512(.A1(new_n5560_), .A2(new_n5561_), .ZN(new_n5562_));
  INV_X1     g5513(.I(new_n5561_), .ZN(new_n5563_));
  NOR2_X1    g5514(.A1(new_n5547_), .A2(new_n5563_), .ZN(new_n5564_));
  INV_X1     g5515(.I(new_n5564_), .ZN(new_n5565_));
  NAND3_X1   g5516(.A1(new_n5546_), .A2(new_n5547_), .A3(new_n5563_), .ZN(new_n5566_));
  NAND3_X1   g5517(.A1(new_n5566_), .A2(new_n5562_), .A3(new_n5565_), .ZN(new_n5567_));
  XOR2_X1    g5518(.A1(new_n5559_), .A2(new_n5567_), .Z(\sin[22] ));
  NOR2_X1    g5519(.A1(new_n128_), .A2(new_n89_), .ZN(new_n5569_));
  INV_X1     g5520(.I(new_n5569_), .ZN(new_n5570_));
  NOR2_X1    g5521(.A1(new_n5546_), .A2(new_n5565_), .ZN(new_n5571_));
  AOI21_X1   g5522(.A1(new_n5562_), .A2(new_n5565_), .B(new_n5571_), .ZN(new_n5572_));
  NAND3_X1   g5523(.A1(new_n5567_), .A2(new_n5539_), .A3(new_n5551_), .ZN(new_n5573_));
  AOI21_X1   g5524(.A1(new_n5573_), .A2(new_n4073_), .B(new_n5572_), .ZN(new_n5574_));
  INV_X1     g5525(.I(new_n5572_), .ZN(new_n5575_));
  NOR2_X1    g5526(.A1(new_n5546_), .A2(new_n5563_), .ZN(new_n5576_));
  NOR3_X1    g5527(.A1(new_n5560_), .A2(new_n5543_), .A3(new_n5561_), .ZN(new_n5577_));
  NOR3_X1    g5528(.A1(new_n5577_), .A2(new_n5576_), .A3(new_n5564_), .ZN(new_n5578_));
  OAI21_X1   g5529(.A1(new_n5558_), .A2(new_n5578_), .B(new_n4073_), .ZN(new_n5579_));
  NOR2_X1    g5530(.A1(new_n5579_), .A2(new_n5575_), .ZN(new_n5580_));
  OAI21_X1   g5531(.A1(new_n5580_), .A2(new_n5574_), .B(new_n5570_), .ZN(\sin[23] ));
  INV_X1     g5532(.I(new_n5571_), .ZN(new_n5582_));
  AOI21_X1   g5533(.A1(new_n5573_), .A2(new_n5582_), .B(new_n5569_), .ZN(new_n5583_));
  NAND2_X1   g5534(.A1(new_n5562_), .A2(new_n5565_), .ZN(new_n5584_));
  NAND4_X1   g5535(.A1(new_n5567_), .A2(new_n5539_), .A3(new_n5584_), .A4(new_n5551_), .ZN(new_n5585_));
  AOI21_X1   g5536(.A1(new_n5583_), .A2(new_n5585_), .B(new_n4074_), .ZN(\sin[24] ));
endmodule


