// Benchmark "source.pla" written by ABC on Sun Mar  6 13:13:10 2022

module pdc  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    \v16.0 , \v16.1 , \v16.2 , \v16.3 , \v16.4 , \v16.5 , \v16.6 , \v16.7 ,
    \v16.8 , \v16.9 , \v16.10 , \v16.11 , \v16.12 , \v16.13 , \v16.14 ,
    \v16.15 , \v16.16 , \v16.17 , \v16.18 , \v16.19 , \v16.20 , \v16.21 ,
    \v16.22 , \v16.23 , \v16.24 , \v16.25 , \v16.26 , \v16.27 , \v16.28 ,
    \v16.29 , \v16.30 , \v16.31 , \v16.32 , \v16.33 , \v16.34 , \v16.35 ,
    \v16.36 , \v16.37 , \v16.38 , \v16.39   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15;
  output \v16.0 , \v16.1 , \v16.2 , \v16.3 , \v16.4 , \v16.5 , \v16.6 ,
    \v16.7 , \v16.8 , \v16.9 , \v16.10 , \v16.11 , \v16.12 , \v16.13 ,
    \v16.14 , \v16.15 , \v16.16 , \v16.17 , \v16.18 , \v16.19 , \v16.20 ,
    \v16.21 , \v16.22 , \v16.23 , \v16.24 , \v16.25 , \v16.26 , \v16.27 ,
    \v16.28 , \v16.29 , \v16.30 , \v16.31 , \v16.32 , \v16.33 , \v16.34 ,
    \v16.35 , \v16.36 , \v16.37 , \v16.38 , \v16.39 ;
  assign \v16.0  = ~v3 & ~v4 & ((~v2 & (v0 ? ~v1 : (v1 & ~v5 & (v7 | (~v7 & ((~v11 & ~v12 & ((~v8 & v9 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) | (v8 & ~v9 & ~v13 & ~v14 & ~v15) | (~v8 & ~v9 & v10 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) | (~v13 & ~v14 & ~v15 & v8 & v9 & ~v10))) | (~v8 & ~v9 & ~v10))))))) | (v0 & ~v1 & v2));
  assign \v16.1  = ~v3 & v4 & ((v0 & ~v1 & v2) | (~v2 & (v0 ? ~v1 : (v1 & ~v5 & (v7 | (~v7 & ((~v8 & ~v9 & ~v10) | (~v11 & ~v12 & (((~v9 ^ ~v10) & ((~v8 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) | (~v14 & ~v15 & v8 & ~v13))) | (~v8 & v9 & v10 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))))))))));
  assign \v16.2  = ~v3 & ~v4 & ((~v2 & (v0 ? (~v1 & v5) : (v1 & ~v5 & v6 & (v7 | (~v7 & ((~v11 & ~v12 & ((~v8 & v9 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) | (v8 & ~v9 & ~v13 & ~v14 & ~v15) | (~v8 & ~v9 & v10 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) | (~v13 & ~v14 & ~v15 & v8 & v9 & ~v10))) | (~v8 & ~v9 & ~v10))))))) | (v0 & ~v1 & v2 & v5));
  assign \v16.3  = ~v3 & ((~v1 & ((v4 & ((v5 & (v0 | (~v0 & ~v2 & v10 & ~v11 & ~v12 & ~v13 & v14 & ~v15 & (~v8 ^ ~v9)) | (~v0 & ~v2 & (((~v8 ^ ~v9) & ((v6 & ((v12 & ((v14 & (((v13 ^ v15) & (v10 ^ v11)) | (v10 & ~v11 & ~v13 & ~v15))) | (v10 & ~v11 & ~v13 & ~v14))) | (v10 & ~v11 & ~v12 & v13 & v14 & ~v15))) | (~v6 & ~v10 & ~v11 & v14 & ~v15 & ~v12 & ~v13))) | (v6 & v10 & ~v11 & v12 & ~v13 & v14 & ~v15 & (~v8 ^ v9)))))) | (~v0 & ~v2 & ~v5 & ~v6 & ((v14 & (~v15 | (v12 & ~v13 & v15))) | (v12 & ~v13 & ~v14))))) | (~v0 & ~v2 & ~v4 & ~v5 & v6 & ((v14 & (~v15 | (v12 & ~v13 & v15)) & ((~v8 & (v9 ? (~v10 & ~v11) : (v10 ^ v11))) | (v8 & ~v9 & ~v10 & ~v11))) | (v12 & ~v13 & ~v14 & ((~v8 & (v9 ? (~v10 & ~v11) : (v10 ^ v11))) | (v8 & ~v9 & ~v10 & ~v11))))) | (~v0 & ~v2 & (((~v8 ^ ~v9) & ((v14 & ((~v15 & ((~v4 & ~v7 & (v5 ? ~v6 : (v6 & v11))) | (v4 & v5 & ~v6 & v7 & v11) | (v4 & v5 & v7 & (v6 ? (v11 & ~v12) : (~v11 & v12))) | (v4 & v5 & v7 & ((~v6 & ~v11 & ~v12 & v13) | (v6 & v11 & v12 & ~v13))))) | (v12 & ~v13 & v15 & (((v4 ? (v7 & ~v11) : (~v7 & v11)) & (~v5 ^ ~v6)) | (v5 & ~v6 & (v4 ? (v7 & v11) : (~v7 & ~v11))))))) | (v12 & ~v13 & ~v14 & ((v11 & ((v5 & (v4 ? v7 : (~v6 & ~v7))) | (~v4 & ~v5 & v6 & ~v7))) | (v5 & ~v6 & ~v11 & (~v4 ^ v7)))) | (~v4 & v5 & ~v6 & v7 & ~v11))) | (v14 & ((~v15 & ((v5 & ~v6 & (~v8 ^ v9) & (~v4 ^ v7)) | (~v4 & ~v5 & v6 & ~v7 & v8 & v9) | (v4 & v5 & v6 & v7 & ~v12 & (~v8 ^ v9)) | (v4 & v5 & v6 & v7 & v12 & v13 & (~v8 ^ v9)))) | (v12 & ~v13 & v15 & ((~v4 & ~v5 & v6 & ~v7 & v8 & v9) | (v5 & (~v8 ^ v9) & (v4 ? v7 : (~v6 & ~v7))))) | (v4 & v5 & v6 & v7 & v11 & v12 & ~v13 & ~v15 & (~v8 ^ v9)))) | (v12 & ~v13 & ~v14 & ((~v4 & ~v5 & v6 & ~v7 & v8 & v9) | (v5 & (~v8 ^ v9) & (v4 ? v7 : (~v6 & ~v7))))) | (v6 & (v12 ? (((v10 ^ ~v11) & ((v14 & (((v13 ^ v15) & ((v4 & v5 & v7 & (~v8 ^ ~v9)) | (~v4 & ~v5 & ~v7 & ~v8 & ~v9))) | (~v4 & ~v5 & ~v7 & ~v13 & ~v15 & ~v8 & ~v9))) | (~v4 & ~v5 & ~v7 & ~v8 & ~v9 & ~v13 & ~v14))) | (~v11 & (((~v8 ^ ~v9) & ((~v13 & ((~v4 & ~v5 & ~v7 & v10) | (v4 & v5 & v7 & ~v10 & ~v14) | (v4 & v5 & v7 & ~v10 & v14 & ~v15))) | (~v4 & ~v5 & ~v7 & v14 & ~v15 & v10 & v13))) | (v4 & v5 & v7 & ~v10 & ~v13 & v14 & ~v15 & (~v8 ^ v9))))) : (v14 & ~v15 & ((~v11 & (((~v8 ^ ~v9) & ((~v4 & ~v5 & ~v7 & v10) | (v4 & v5 & v7 & ~v10))) | (~v8 & ~v9 & ~v10 & ~v4 & ~v5 & ~v7))) | (~v4 & ~v5 & ~v7 & ~v8 & ~v9 & v10 & v11))))))))) | (~v0 & v1 & ~v2 & v4 & ~v5 & v6 & (v7 | (~v7 & ((~v8 & ~v9 & ~v10) | (~v11 & ~v12 & (((~v9 ^ ~v10) & ((~v8 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) | (~v14 & ~v15 & v8 & ~v13))) | (~v8 & v9 & v10 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))))))));
  assign \v16.4  = ~v0 & ~v1 & ~v2 & ~v3 & ((v12 & (((v10 ^ v11) & ((((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6)))) & (v13 | (~v13 & v14 & v15))) | (v6 & ((v14 & (((v13 ^ v15) & ((v4 & v5 & ~v7 & (~v8 ^ ~v9)) | (~v4 & ~v5 & v7 & ~v8 & ~v9))) | (~v4 & ~v5 & v7 & ~v8 & ~v9 & v13 & v15))) | (~v4 & ~v5 & v7 & ~v8 & ~v9 & v13 & ~v14))))) | ((~v8 ^ ~v9) & (((v10 ^ ~v11) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6)))) & (v13 | (~v13 & v14 & v15))) | (v6 & ((~v10 & ((~v5 & v7 & ((v14 & ((~v4 & ~v11 & (v13 | (~v13 & v15))) | (~v13 & v15 & v4 & v11))) | (~v4 & ~v11 & v13 & ~v14))) | (v4 & v5 & ~v7 & v11 & v13 & (~v14 | (v14 & v15))))) | (v4 & ~v5 & v7 & v10 & v14 & v15 & v11 & ~v13))))) | ((v10 ^ ~v11) & (~v8 ^ v9) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6)))) & (v13 | (~v13 & v14 & v15))) | (v4 & v5 & v6 & ~v7 & ~v10 & v11 & v13 & v14 & v15 & (~v8 ^ v9)))) | ((~v8 ^ ~v9) & ((~v12 & v14 & ((v15 & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))))) | (v4 & v5 & ~v6 & ~v13 & ~v15 & ~v7 & v11))) | (~v6 & v7 & v11 & ~v4 & v5))) | (~v12 & v14 & v15 & (~v8 ^ v9) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))))) | (v6 & ~v12 & v14 & v15 & ((~v10 & (((~v8 ^ ~v9) & ((v4 & v5 & ~v7 & v11) | (v7 & ~v11 & ~v4 & ~v5))) | (~v4 & ~v5 & v7 & ~v8 & ~v9 & v11))) | (~v4 & ~v5 & v7 & v10 & ~v11 & ~v8 & ~v9))));
  assign \v16.5  = ~v0 & ~v1 & ~v2 & ~v3 & (((~v8 ^ ~v9) & (((v14 ^ v15) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))))) | ((v14 ^ ~v15) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6)))) & (v12 ^ v13)) | (~v11 & ((v4 & ~v13 & v14 & ((~v5 & v6 & v7 & v12 & v15) | (v5 & ~v6 & ~v7 & ~v12 & ~v15))) | (~v4 & v5 & ~v6 & v7))))) | ((v14 ^ v15) & (~v8 ^ v9) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))))) | ((v14 ^ ~v15) & (~v8 ^ v9) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6)))) & (v12 ^ v13)) | (v6 & (((v14 ^ v15) & (((v10 ? (~v11 & ~v13) : (v11 & v13)) & ((v12 & ((v4 & v5 & ~v7 & (~v8 ^ ~v9)) | (~v4 & ~v5 & v7 & ~v8 & ~v9))) | (~v4 & ~v5 & v7 & ~v8 & ~v9 & ~v12))) | (~v4 & ~v5 & v7 & ((~v10 & ((~v11 & (~v8 ^ ~v9)) | (~v8 & ~v9 & v11 & ~v13))) | (~v8 & ~v9 & v10 & ~v11 & v13))))) | ((v12 ^ v13) & ((~v10 & (((~v8 ^ ~v9) & ((~v4 & ~v5 & v7 & ~v11 & (v14 ^ ~v15)) | (v4 & v5 & ~v7 & v11 & v14 & v15))) | (~v4 & ~v5 & v7 & ~v8 & ~v9 & v11 & (v14 ^ ~v15)))) | (~v4 & ~v5 & v7 & ~v8 & ~v9 & v10 & ~v11 & (v14 ^ ~v15)))) | (v4 & v5 & ~v7 & v10 & ~v11 & ((v12 & ~v13 & v14 & ~v15 & (~v8 ^ v9)) | ((~v8 ^ ~v9) & ((v14 & (v12 ? (v13 ^ v15) : ~v15)) | (~v14 & ~v15 & v12 & ~v13))))))));
  assign \v16.6  = ~v0 & ~v1 & v3;
  assign \v16.7  = ~v3 & ~v4 & ~v5 & ((v0 & ~v1 & v2) | (~v2 & (v0 ? ~v1 : (v1 & ~v6 & (v7 | (~v7 & ((~v11 & ~v12 & ((~v8 & v9 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) | (v8 & ~v9 & ~v13 & ~v14 & ~v15) | (~v8 & ~v9 & v10 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) | (~v13 & ~v14 & ~v15 & v8 & v9 & ~v10))) | (~v8 & ~v9 & ~v10))))))));
  assign \v16.8  = ~v3 & ((~v1 & ((~v5 & ((v4 & (v0 | (~v0 & ~v2 & ~v6 & ((~v14 & (v15 | (~v12 & v13 & ~v15))) | (~v12 & v13 & v14))))) | (~v0 & ~v2 & ~v4 & v6 & ((~v14 & ((~v8 & (v9 ? (~v10 & ~v11) : (v10 ^ v11))) | (v8 & ~v9 & ~v10 & ~v11)) & (v15 | (~v12 & v13 & ~v15))) | (~v12 & v13 & v14 & ((~v8 & (v9 ? (~v10 & ~v11) : (v10 ^ v11))) | (v8 & ~v9 & ~v10 & ~v11))))))) | (~v0 & ~v2 & v4 & v5 & v6 & (~v8 ^ ~v9) & (v10 ? (~v11 & ((~v14 & v15 & v12 & ~v13) | (v14 & ~v15 & ~v12 & v13))) : (v11 & v13 & v15 & (v12 ^ v14)))) | (~v0 & ~v2 & ((~v14 & (((v10 ^ ~v11) & (((~v8 ^ v9) & ((v5 & (v4 ? v7 : (~v6 & ~v7))) | (~v4 & ~v5 & v6 & ~v7)) & (v15 | (~v12 & v13 & ~v15))) | (v5 & (~v8 ^ ~v9) & (v4 ? v7 : (~v6 & ~v7)) & (v15 | (~v12 & v13 & ~v15))))) | ((((v10 ^ v11) & ((~v4 & ~v7 & (~v5 ^ ~v6)) | (v4 & v5 & ~v6 & v7))) | (~v4 & ~v5 & v6 & ~v7 & v10 & v11)) & (~v8 ^ ~v9) & (v15 | (~v12 & v13 & ~v15))) | ((v10 ^ v11) & ((v15 & ((~v4 & ~v5 & v6 & ~v7 & v8 & v9) | (v5 & (~v8 ^ v9) & (v4 ? v7 : (~v6 & ~v7))) | (v4 & v5 & v6 & v7 & ~v12 & (~v8 ^ ~v9)))) | (~v12 & v13 & ~v15 & ((~v4 & ~v5 & v6 & ~v7 & v8 & v9) | (v5 & (((~v8 ^ v9) & (v4 ? v7 : (~v6 & ~v7))) | (v4 & v6 & v7 & (~v8 ^ ~v9)))))))) | (v4 & v5 & v6 & v7 & v12 & v15 & (~v8 ^ ~v9) & (v10 ? (~v11 & v13) : (v11 & ~v13))))) | (~v12 & v13 & v14 & (((v10 ^ ~v11) & (((~v8 ^ v9) & ((v5 & (v4 ? v7 : (~v6 & ~v7))) | (~v4 & ~v5 & v6 & ~v7))) | (v5 & (~v8 ^ ~v9) & (v4 ? v7 : (~v6 & ~v7))))) | ((~v8 ^ ~v9) & (((v10 ^ v11) & ((~v4 & ~v7 & (~v5 ^ ~v6)) | (v4 & v5 & ~v6 & v7))) | (~v4 & ~v5 & v6 & ~v7 & v10 & v11))) | ((v10 ^ v11) & ((~v4 & ~v5 & v6 & ~v7 & v8 & v9) | (v5 & (~v8 ^ v9) & (v4 ? v7 : (~v6 & ~v7))))) | (v4 & v5 & v6 & v7 & (~v8 ^ ~v9) & (v10 ? (~v11 & v15) : (v11 & ~v15))))))))) | (~v0 & v1 & ~v2 & v4 & ~v5 & ~v6 & (v7 | (~v7 & ((~v8 & ~v9 & ~v10) | (~v11 & ~v12 & (((~v9 ^ ~v10) & ((~v8 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) | (~v14 & ~v15 & v8 & ~v13))) | (~v8 & v9 & v10 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))))))));
  assign \v16.9  = ~v0 & ~v1 & ~v2 & ~v3 & ((~v15 & (((v10 ^ v11) & ((((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6)))) & (~v14 | (~v12 & ~v13 & v14))) | (~v4 & ~v5 & v6 & v7 & ~v8 & ~v9 & (~v14 | (~v12 & ~v13 & v14))))) | ((~v8 ^ ~v9) & (((v10 ^ ~v11) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6)))) & (~v14 | (~v12 & ~v13 & v14))) | (v6 & ((~v11 & ((~v13 & (((v12 ^ v14) & ((v4 & v5 & ~v7 & v10) | (~v4 & ~v5 & v7 & ~v10))) | (~v4 & ~v5 & v7 & ~v10 & ~v12 & ~v14))) | (~v4 & ~v5 & v7 & ~v10 & v13 & ~v14))) | (v4 & v5 & ~v7 & ~v10 & v13 & ~v14 & v11 & v12))))) | ((v10 ^ ~v11) & (~v8 ^ v9) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6)))) & (~v14 | (~v12 & ~v13 & v14))))) | (~v12 & ~v13 & v15 & (((v10 ^ v11) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))) | (~v4 & ~v5 & v6 & v7 & ~v8 & ~v9))) | ((~v8 ^ ~v9) & (((v10 ^ ~v11) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))))) | (~v4 & ~v5 & v6 & v7 & ~v10 & ~v11))) | ((v10 ^ ~v11) & (~v8 ^ v9) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))))) | (v4 & v5 & v6 & ~v7 & ~v10 & v11 & v14 & (~v8 ^ ~v9)))));
  assign \v16.10  = ~v0 & ~v1 & ~v2 & ~v3 & v4 & v5 & (((~v8 ^ ~v9) & ((v6 & v7) | (~v6 & ~v7 & ~v12 & ~v13 & v14 & ~v15))) | (v6 & v7 & (~v8 ^ v9)));
  assign \v16.11  = ~v0 & ~v1 & ~v2 & ~v3 & ~v4 & ~v5 & v6 & v7 & ((~v8 & (v9 ? (~v10 & ~v11) : (v10 ^ v11))) | (v8 & ~v9 & ~v10 & ~v11));
  assign \v16.12  = ~v0 & ~v1 & ~v2 & ~v3 & v4 & ~v5 & ~v6 & ~v7;
  assign \v16.13  = ~v0 & ~v1 & ~v2 & ~v3 & v4 & ~v5 & ~v6 & v7;
  assign \v16.14  = v0 & ~v1;
  assign \v16.15  = (~v1 & (v0 ^ v2)) | (~v0 & v1 & v2);
  assign \v16.16  = ~v0 & ~v1 & ~v2 & ~v3 & v8 & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))) | (~v9 & ((v4 & ~v13 & v14 & ((~v5 & v6 & v7 & v12 & v15) | (v5 & ~v6 & ~v7 & ~v12 & ~v15))) | (~v4 & v5 & ~v6 & v7))) | (v6 & (v4 ? (v5 & ~v7 & ((((v10 & ~v11 & ~v13 & ~v15) | (~v10 & v11 & v13 & v15)) & (v9 ? (v12 & v14) : (v12 | (~v12 & v14)))) | (~v9 & ((v14 & ((~v13 & v15 & ~v10 & v11) | (v13 & ~v15 & v10 & ~v11) | (v12 & ((~v13 & v15 & v10 & ~v11) | (v13 & ~v15 & ~v10 & v11))))) | (v12 & ~v14 & ((~v13 & v15 & v10 & ~v11) | (v13 & ~v15 & ~v10 & v11))))))) : (~v5 & v7 & ~v9 & ~v10 & ~v11))));
  assign \v16.17  = ~v0 & ~v1 & ~v2 & ~v3 & v9 & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))) | (~v8 & ((v4 & ~v13 & v14 & ((~v5 & v6 & v7 & v12 & v15) | (v5 & ~v6 & ~v7 & ~v12 & ~v15))) | (~v4 & v5 & ~v6 & v7))) | (v6 & (v4 ? (v5 & ~v7 & ((((v10 & ~v11 & ~v13 & ~v15) | (~v10 & v11 & v13 & v15)) & (v8 ? (v12 & v14) : (v12 | (~v12 & v14)))) | (~v8 & ((v14 & ((~v13 & v15 & ~v10 & v11) | (v13 & ~v15 & v10 & ~v11) | (v12 & ((~v13 & v15 & v10 & ~v11) | (v13 & ~v15 & ~v10 & v11))))) | (v12 & ~v14 & ((~v13 & v15 & v10 & ~v11) | (v13 & ~v15 & ~v10 & v11))))))) : (~v5 & v7 & ~v8 & ~v10 & ~v11))));
  assign \v16.18  = ~v0 & ~v1 & ~v2 & ~v3 & v10 & (((~v8 ^ v9) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))))) | ((~v8 ^ ~v9) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))) | (v4 & ~v13 & v14 & ((~v5 & v6 & v7 & v12 & v15) | (v5 & ~v6 & ~v7 & ~v12 & ~v15))) | (~v4 & v5 & ~v6 & v7))) | (v6 & ~v11 & ((v14 & ((~v15 & ((v4 & v5 & ~v7 & (~v8 ^ ~v9)) | (~v4 & ~v5 & v7 & ~v8 & ~v9))) | (~v4 & ~v5 & v7 & ~v8 & ~v9 & v15))) | (~v4 & ~v5 & v7 & ~v8 & ~v9 & ~v14) | (v4 & v5 & ~v7 & v12 & ~v13 & (v8 ? (v14 ? (v9 ^ v15) : ~v9) : (v14 ? (~v9 ^ v15) : v9))))));
  assign \v16.19  = ~v0 & ~v1 & ~v2 & ~v3 & v11 & (((~v8 ^ v9) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))))) | ((~v8 ^ ~v9) & ((~v7 & (v4 ? (~v5 & ~v6) : (~v5 ^ ~v6))) | (v4 & v7 & (v5 | (~v5 & ~v6))) | (v4 & ~v13 & v14 & ((~v5 & v6 & v7 & v12 & v15) | (v5 & ~v6 & ~v7 & ~v12 & ~v15))) | (~v4 & v5 & ~v6 & v7))) | (v6 & ~v10 & ((~v4 & ~v5 & v7 & ~v8 & ~v9 & ~v14) | (v14 & ((v15 & ((v4 & v5 & ~v7 & (~v8 ^ ~v9)) | (~v4 & ~v5 & v7 & ~v8 & ~v9))) | (~v4 & ~v5 & v7 & ~v8 & ~v9 & ~v15))) | (v4 & v5 & ~v7 & v12 & v13 & (v8 ? (v14 ? (~v9 ^ v15) : ~v9) : (v14 ? (v9 ^ v15) : v9))))));
  assign \v16.20  = ~v0 & ~v1 & ~v2 & ~v3 & ~v4 & ((~v5 & v6 & v7 & ((~v8 & (v9 ? (~v10 & ~v11) : (v10 ^ v11))) | (v8 & ~v9 & ~v10 & ~v11))) | ((~v8 ^ ~v9) & ((~v7 & (~v5 ^ ~v6)) | (v5 & ~v6 & v7))) | (~v7 & (~v8 ^ v9) & (~v5 ^ ~v6)));
  assign \v16.21  = ~v0 & ~v1 & ~v2 & ~v3 & ~v4 & v5 & ~v6 & ((v8 & ~v9) | (~v8 & v9) | (~v7 & (~v8 ^ v9)));
  assign \v16.22  = ~v0 & ~v1 & ~v2 & ~v3 & v4 & ~v13 & v14 & (~v8 ^ ~v9) & ((~v5 & v6 & v7 & v12 & v15) | (v5 & ~v6 & ~v7 & ~v12 & ~v15));
  assign \v16.23  = ~v0 & ~v2 & ((~v3 & (((v14 ^ v15) & ((~v8 & ((v9 & ((v10 & ((~v11 & ((~v12 & ((v4 & ((~v13 & (v1 ? ~v7 : (v5 & v7))) | (~v1 & v5 & v7 & v13))) | (v1 & ~v4 & ~v5 & ~v7 & ~v13))) | (~v1 & v4 & v5 & v7 & v12))) | (~v1 & v4 & v5 & v7 & v11))) | (~v1 & v4 & v5 & v7 & ~v10))) | (~v1 & v4 & v5 & v7 & ~v9))) | (~v1 & v4 & v5 & v7 & v8) | (v1 & ~v4 & v5 & v6 & ~v7 & ~v8 & v9 & v10 & ~v11 & ~v12 & ~v13))) | (~v8 & ((v9 & ((v10 & ((~v11 & ((~v12 & ((v13 & ((v4 & ((~v14 & ~v15 & (v1 ? ~v7 : (v5 & v7))) | (~v1 & v5 & v7 & v14 & v15))) | (v1 & ~v4 & ~v5 & ~v7 & ~v14 & ~v15))) | (~v1 & v4 & v5 & v7 & ~v13 & (v14 ^ ~v15)))) | (~v1 & v4 & v5 & v7 & v12 & (v14 ^ ~v15)))) | (~v1 & v4 & v5 & v7 & v11 & (v14 ^ ~v15)))) | (~v1 & v4 & v5 & v7 & ~v10 & (v14 ^ ~v15)))) | (~v1 & v4 & v5 & v7 & ~v9 & (v14 ^ ~v15)))) | (~v1 & v4 & v5 & v7 & v8 & (v14 ^ ~v15)) | (v1 & ~v4 & v5 & v6 & ~v7 & ~v8 & v9 & v10 & ~v11 & ~v14 & ~v15 & ~v12 & v13))) | (v1 & v3 & v4 & v5 & ~v6 & ~v7));
  assign \v16.24  = ~v0 & v1 & ~v2 & ~v3 & ~v7 & ~v11 & ~v12 & ((~v13 & ((~v14 & ((~v9 & ((~v4 & ~v5 & v8 & ~v10 & ~v15) | (v4 & v5 & ~v6 & ~v8 & v10 & v15))) | (v4 & v5 & ~v6 & ~v8 & v9 & v15))) | (v4 & v5 & ~v6 & ~v8 & v14 & ~v15 & (v9 | (~v9 & v10))))) | (v4 & v5 & ~v6 & ~v8 & v13 & ~v14 & ~v15 & (v9 | (~v9 & v10))));
  assign \v16.25  = ~v0 & ~v1 & ~v2 & ~v3 & v4 & v5 & v7;
  assign \v16.26  = ~v0 & ~v1 & ~v2 & ~v3 & v4 & v5 & v6 & ~v7 & ((v14 & (((~v8 ^ ~v9) & (v10 ? (~v11 & ~v15) : (v11 & v15))) | (v12 & (((~v8 ^ v9) & ((v10 & ~v11 & ~v13 & ~v15) | (~v10 & v11 & v13 & v15))) | ((~v8 ^ ~v9) & ((~v13 & v15 & v10 & ~v11) | (v13 & ~v15 & ~v10 & v11))))))) | (v12 & ~v14 & (~v8 ^ ~v9) & (v10 ? (~v11 & ~v13) : (v11 & v13))));
  assign \v16.27  = v7 & v6 & v5 & ~v4 & ~v3 & ~v2 & v0 & v1;
  assign \v16.28  = (~v7 & ((~v2 & (v0 ? (~v1 & ~v3) : (v1 & ~v9 & ((~v5 & ((~v6 & (v3 ? (v8 ^ v10) : (~v8 & v10 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))) | (~v3 & v6 & ~v8 & v10 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))) | (~v3 & v5 & v6 & ~v8 & v10 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))))) | (v0 & ~v1 & v2 & ~v3))) | (~v0 & v1 & ~v2 & ~v3 & v5 & v6 & v7 & ~v8 & ~v9 & v10 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) | (~v0 & v1 & ~v2 & v4 & (v3 ? (~v5 & (v6 | (~v6 & v7))) : (v5 & ~v6 & ~v7 & ~v8 & ~v9 & v10 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15)))));
  assign \v16.29  = (~v2 & (v0 ? (~v1 & ~v3 & v7) : (v1 & ~v10 & ((~v7 & ((~v5 & ((~v6 & (v3 ? (~v8 ^ ~v9) : (~v8 & v9 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))) | (~v3 & v6 & ~v8 & v9 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))) | (~v3 & v5 & v6 & ~v8 & v9 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))) | (~v3 & v5 & v6 & v7 & ~v8 & v9 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))))) | (v0 & ~v1 & v2 & ~v3 & v7) | (~v0 & v1 & ~v2 & v4 & v5 & (v3 ? (v6 | (~v6 & v7)) : (~v6 & ~v7 & ~v8 & v9 & ~v10 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15)))));
  assign \v16.30  = ~v3 & ((v0 & ~v1 & v2) | (~v2 & (v0 ? ~v1 : (v1 & v5 & v6 & ~v8 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15)) & (~v9 ^ ~v10)))) | (~v0 & v1 & ~v2 & ((~v5 & (v7 | (~v7 & ~v8 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15)) & (~v9 ^ ~v10)))) | (v4 & v5 & ~v6 & ~v7 & ~v8 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15)) & (~v9 ^ ~v10)))));
  assign \v16.31  = ~v0 & v1 & ~v2 & ~v7 & ((~v8 & ((~v5 & ((~v4 & ((~v6 & (v3 ? (~v9 ^ ~v10) : (~v9 & ~v10))) | (~v9 & ~v10 & ~v3 & v6))) | (v3 & v4 & ~v6 & (~v9 ^ ~v10)))) | (~v3 & ~v4 & v5 & v6 & ~v9 & ~v10))) | (v3 & ~v5 & ~v6 & v8 & ~v9 & ~v10));
  assign \v16.32  = ~v0 & v1 & ~v2 & ((v7 & ((v4 & ((v6 & (v3 | (~v3 & ~v5))) | (~v3 & ~v5 & ~v6))) | (~v3 & ~v4 & ~v5))) | (v3 & v4 & v5 & ~v6 & ~v7));
  assign \v16.33  = ~v3 & ((~v2 & (v0 ? (~v1 & ~v6) : (v1 & v5 & v6 & ~v8 & ~v11 & ~v12 & ~v13 & ~v14 & v15 & (~v9 ^ ~v10)))) | (v0 & ~v1 & v2 & ~v6) | (~v0 & v1 & ~v2 & ~v7 & ~v8 & ((~v11 & ~v12 & ~v13 & ~v14 & v15 & ((~v5 & (v9 | (~v9 & v10))) | (v9 & v10 & v5 & v6) | (v4 & v5 & ~v6 & (v9 | (~v9 & v10))))) | (v4 & ~v5 & ~v9 & ~v10))));
  assign \v16.34  = ~v3 & ((v6 & ((v0 & ~v1 & v2) | (~v2 & (v0 ? ~v1 : (v1 & v5 & ~v8 & ~v11 & ~v12 & ~v13 & v14 & ~v15 & (~v9 ^ ~v10)))) | (~v0 & ~v2 & ((~v1 & v4 & v5 & v7 & v8) | (~v8 & ((~v1 & v4 & v5 & v7 & ~v9) | (v9 & ((~v1 & v4 & v5 & v7 & v11) | (~v11 & ((~v1 & v4 & v5 & v7 & v12) | (~v12 & ((~v13 & ((v14 & ((~v15 & ((v1 & ~v5 & ~v7) | (v5 & v7 & ~v1 & v4))) | (~v1 & v4 & v5 & v7 & v15))) | (~v1 & v4 & v5 & v7 & ~v14))) | (~v1 & v4 & v5 & v7 & v13))))))))) | (v1 & ~v7 & ~v8 & ((v10 & ~v11 & ~v12 & ~v13 & v14 & ~v15 & (~v5 ^ v9)) | (v4 & ~v9 & ~v10))))))) | (~v0 & ~v2 & ~v6 & ((~v1 & v4 & v5 & v7 & v8) | (~v8 & ((~v1 & v4 & v5 & v7 & ~v9) | (v9 & ((~v1 & v4 & v5 & v7 & v11) | (~v11 & ((~v1 & v4 & v5 & v7 & v12) | (~v12 & ((~v1 & v4 & v5 & v7 & v13) | (~v13 & ((~v1 & v4 & v5 & v7 & ~v14) | (v14 & ((v4 & ((~v15 & (v1 ? ~v7 : (v5 & v7))) | (~v1 & v5 & v7 & v15))) | (v1 & ~v4 & ~v5 & ~v7 & ~v15))))))))))))) | (v1 & ~v7 & ~v8 & ~v9 & v10 & ~v11 & ~v12 & ~v13 & v14 & ~v15 & (v4 | (~v4 & ~v5))))));
  assign \v16.35  = ~v0 & v1 & ~v2 & ~v3 & ~v8 & ((~v11 & ~v12 & v13 & ~v14 & ~v15 & (((~v9 ^ ~v10) & ((~v5 & ~v6 & ~v7) | (v6 & (v5 | (~v5 & ~v7))) | (v4 & v5 & ~v6 & ~v7))) | (~v7 & v9 & v10 & (v4 | (~v4 & ~v5) | (~v4 & v5 & v6))))) | (v4 & ~v5 & ~v6 & ~v7 & ~v9 & ~v10));
  assign \v16.36  = v4 & ((v0 & ~v1 & v2 & ~v3) | (~v2 & (v0 ? (~v1 & ~v3) : (((~v9 ^ ~v10) & ((~v3 & (((v14 ^ v15) & ((~v8 & ((~v11 & ((~v12 & ((~v13 & (v1 ? ~v7 : (v5 & v7))) | (~v1 & v5 & v7 & v13))) | (~v1 & v5 & v7 & v12))) | (~v1 & v5 & v7 & v11))) | (~v1 & v5 & v7 & v8))) | (~v8 & ((~v11 & ((~v12 & ((v13 & ((~v14 & ~v15 & (v1 ? ~v7 : (v5 & v7))) | (~v1 & v5 & v7 & v14 & v15))) | (~v1 & v5 & v7 & ~v13 & (v14 ^ ~v15)))) | (~v1 & v5 & v7 & v12 & (v14 ^ ~v15)))) | (~v1 & v5 & v7 & v11 & (v14 ^ ~v15)))) | (~v1 & v5 & v7 & v8 & (v14 ^ ~v15)) | (v1 & v5 & v6 & v7 & ~v8 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))) | (v1 & v3 & ~v5 & ~v6 & ~v7 & ~v8))) | (~v6 & (v1 ? ((~v7 & (v3 ? (v5 | (~v9 & ~v10 & ~v5 & v8)) : (~v8 & v9 & v10 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))))) | (~v3 & ~v5 & v7)) : (~v3 & v5 & v7 & (v9 ^ ~v10)))) | (~v3 & v6 & (((v14 ^ v15) & ((~v8 & ((v9 & v10 & ((~v11 & ((~v12 & ((~v13 & (v1 ? ~v7 : (v5 & v7))) | (~v1 & v5 & v7 & v13))) | (~v1 & v5 & v7 & v12))) | (~v1 & v5 & v7 & v11))) | (~v1 & v5 & v7 & ~v9 & ~v10))) | (~v1 & v5 & v7 & v8 & (v9 ^ ~v10)))) | (v1 & ((~v5 & (v7 | (v9 & v10 & ~v7 & ~v8 & v13 & ~v14 & ~v15 & ~v11 & ~v12))) | (v13 & ~v14 & ~v15 & ~v11 & ~v12 & v5 & ~v7 & ~v8 & v9 & v10))) | (~v1 & v5 & v7 & (v14 ^ ~v15) & (v9 ^ ~v10))))))));
  assign \v16.37  = ~v4 & ((v0 & ~v1 & v2 & ~v3) | (~v2 & (v0 ? (~v1 & ~v3) : (v1 & ((~v8 & (((~v9 ^ ~v10) & ((~v3 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15)) & ((~v5 & ~v6 & ~v7) | (v6 & (v5 | (~v5 & ~v7))))) | (~v6 & ~v7 & v3 & ~v5))) | (~v3 & ~v7 & (~v5 | (v5 & v6)) & (v9 ? (v10 & ~v11 & ~v12 & (v13 ? (~v14 & ~v15) : (v14 ^ v15))) : ~v10)))) | (~v5 & ((~v3 & v7) | (v8 & ~v9 & ~v10 & v3 & ~v6 & ~v7))))))));
  assign \v16.38  = ~v0 & v1 & ~v2 & v3 & v4 & ~v6 & v7;
  assign \v16.39  = ~v0 & v1 & ~v2 & v3 & v4 & v6 & ~v7;
endmodule


