// Benchmark "bar" written by ABC on Thu Sep 14 18:32:26 2023

module bar ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] , \shift[2] ,
    \shift[3] , \shift[4] , \shift[5] , \shift[6] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] ,
    \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ;
  wire new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n826_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n946_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n956_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n979_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n994_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1003_, new_n1004_, new_n1005_, new_n1007_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1037_, new_n1038_, new_n1039_,
    new_n1041_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1054_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1068_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1079_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1471_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1480_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1549_, new_n1550_, new_n1552_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1588_, new_n1589_, new_n1591_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1638_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1656_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1663_, new_n1664_, new_n1665_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1688_, new_n1689_,
    new_n1690_, new_n1692_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_,
    new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_,
    new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_,
    new_n1792_, new_n1793_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2192_, new_n2193_, new_n2194_,
    new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2274_, new_n2275_, new_n2276_, new_n2277_,
    new_n2278_, new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_,
    new_n2285_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2305_,
    new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_,
    new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_,
    new_n2318_, new_n2319_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_,
    new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_,
    new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_,
    new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2356_, new_n2357_,
    new_n2358_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2373_, new_n2374_, new_n2375_, new_n2377_, new_n2378_, new_n2379_,
    new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_,
    new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_,
    new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_,
    new_n2462_, new_n2463_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_,
    new_n2577_, new_n2578_, new_n2579_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2646_, new_n2647_,
    new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_,
    new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2660_,
    new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_,
    new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_,
    new_n2673_, new_n2674_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_,
    new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_,
    new_n2769_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2832_, new_n2833_, new_n2834_,
    new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_,
    new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2931_, new_n2932_,
    new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2970_, new_n2971_,
    new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_,
    new_n2979_, new_n2980_, new_n2982_, new_n2983_, new_n2985_, new_n2986_,
    new_n2988_, new_n2989_, new_n2991_, new_n2992_, new_n2994_, new_n2995_,
    new_n2997_, new_n2998_, new_n3000_, new_n3001_, new_n3003_, new_n3004_,
    new_n3006_, new_n3007_, new_n3009_, new_n3010_, new_n3012_, new_n3013_,
    new_n3015_, new_n3016_, new_n3018_, new_n3019_, new_n3021_, new_n3022_,
    new_n3024_, new_n3025_, new_n3027_, new_n3028_, new_n3030_, new_n3031_,
    new_n3033_, new_n3034_, new_n3036_, new_n3037_, new_n3039_, new_n3040_,
    new_n3042_, new_n3043_, new_n3045_, new_n3046_, new_n3048_, new_n3049_,
    new_n3051_, new_n3052_, new_n3054_, new_n3055_, new_n3057_, new_n3058_,
    new_n3060_, new_n3061_, new_n3063_, new_n3065_, new_n3067_, new_n3068_,
    new_n3070_, new_n3071_, new_n3073_, new_n3074_, new_n3076_, new_n3077_,
    new_n3079_, new_n3080_, new_n3082_, new_n3083_, new_n3085_, new_n3086_,
    new_n3088_, new_n3089_, new_n3091_, new_n3092_, new_n3094_, new_n3095_,
    new_n3097_, new_n3098_, new_n3100_, new_n3101_, new_n3103_, new_n3104_,
    new_n3106_, new_n3107_, new_n3109_, new_n3110_, new_n3112_, new_n3113_,
    new_n3115_, new_n3116_, new_n3118_, new_n3119_, new_n3121_, new_n3123_,
    new_n3124_, new_n3126_, new_n3127_, new_n3129_, new_n3130_, new_n3132_,
    new_n3133_, new_n3135_, new_n3136_, new_n3138_, new_n3139_, new_n3141_,
    new_n3142_, new_n3144_, new_n3145_, new_n3147_, new_n3148_, new_n3150_,
    new_n3151_, new_n3153_, new_n3154_, new_n3156_, new_n3158_, new_n3159_,
    new_n3161_, new_n3162_, new_n3164_, new_n3165_;
  INV_X1     g0000(.I(\shift[6] ), .ZN(new_n264_));
  INV_X1     g0001(.I(\shift[4] ), .ZN(new_n265_));
  INV_X1     g0002(.I(\shift[5] ), .ZN(new_n266_));
  NAND3_X1   g0003(.A1(\a[117] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n267_));
  NAND2_X1   g0004(.A1(\shift[0] ), .A2(\shift[1] ), .ZN(new_n268_));
  INV_X1     g0005(.I(\shift[1] ), .ZN(new_n269_));
  NOR2_X1    g0006(.A1(new_n269_), .A2(\a[117] ), .ZN(new_n270_));
  NAND2_X1   g0007(.A1(new_n270_), .A2(new_n268_), .ZN(new_n271_));
  NAND2_X1   g0008(.A1(new_n271_), .A2(new_n267_), .ZN(new_n272_));
  NAND3_X1   g0009(.A1(\a[119] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n273_));
  INV_X1     g0010(.I(\a[119] ), .ZN(new_n274_));
  NAND3_X1   g0011(.A1(new_n274_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n275_));
  OR2_X2     g0012(.A1(\shift[2] ), .A2(\shift[3] ), .Z(new_n276_));
  INV_X1     g0013(.I(\a[118] ), .ZN(new_n277_));
  INV_X1     g0014(.I(\a[120] ), .ZN(new_n278_));
  NOR2_X1    g0015(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1   g0016(.A1(new_n279_), .A2(new_n276_), .ZN(new_n280_));
  AOI21_X1   g0017(.A1(new_n273_), .A2(new_n275_), .B(new_n280_), .ZN(new_n281_));
  NAND3_X1   g0018(.A1(\a[121] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n282_));
  NOR2_X1    g0019(.A1(new_n269_), .A2(\a[121] ), .ZN(new_n283_));
  NAND2_X1   g0020(.A1(new_n283_), .A2(new_n268_), .ZN(new_n284_));
  NAND2_X1   g0021(.A1(new_n284_), .A2(new_n282_), .ZN(new_n285_));
  NAND3_X1   g0022(.A1(\a[123] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n286_));
  INV_X1     g0023(.I(\a[123] ), .ZN(new_n287_));
  NAND3_X1   g0024(.A1(new_n287_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n288_));
  NAND3_X1   g0025(.A1(new_n276_), .A2(\a[122] ), .A3(\a[124] ), .ZN(new_n289_));
  AOI21_X1   g0026(.A1(new_n286_), .A2(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND4_X1   g0027(.A1(new_n281_), .A2(new_n290_), .A3(new_n272_), .A4(new_n285_), .ZN(new_n291_));
  NAND3_X1   g0028(.A1(\a[125] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n292_));
  INV_X1     g0029(.I(\a[125] ), .ZN(new_n293_));
  INV_X1     g0030(.I(\shift[0] ), .ZN(new_n294_));
  NAND3_X1   g0031(.A1(new_n293_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n295_));
  NAND2_X1   g0032(.A1(new_n295_), .A2(new_n292_), .ZN(new_n296_));
  NAND3_X1   g0033(.A1(\a[0] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n297_));
  INV_X1     g0034(.I(new_n297_), .ZN(new_n298_));
  NOR3_X1    g0035(.A1(new_n294_), .A2(\a[0] ), .A3(\shift[1] ), .ZN(new_n299_));
  NOR2_X1    g0036(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1     g0037(.I(\a[126] ), .ZN(new_n301_));
  INV_X1     g0038(.I(\a[127] ), .ZN(new_n302_));
  NOR2_X1    g0039(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1   g0040(.A1(new_n303_), .A2(new_n276_), .ZN(new_n304_));
  NOR2_X1    g0041(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1   g0042(.A1(\a[113] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n306_));
  INV_X1     g0043(.I(\a[113] ), .ZN(new_n307_));
  NAND3_X1   g0044(.A1(new_n307_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n308_));
  NAND2_X1   g0045(.A1(new_n308_), .A2(new_n306_), .ZN(new_n309_));
  NAND3_X1   g0046(.A1(\a[115] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n310_));
  INV_X1     g0047(.I(new_n310_), .ZN(new_n311_));
  NOR3_X1    g0048(.A1(new_n294_), .A2(\a[115] ), .A3(\shift[1] ), .ZN(new_n312_));
  NOR2_X1    g0049(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1   g0050(.A1(new_n276_), .A2(\a[114] ), .A3(\a[116] ), .ZN(new_n314_));
  NOR2_X1    g0051(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND4_X1   g0052(.A1(new_n305_), .A2(new_n315_), .A3(new_n296_), .A4(new_n309_), .ZN(new_n316_));
  NOR4_X1    g0053(.A1(new_n291_), .A2(new_n316_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n317_));
  NAND2_X1   g0054(.A1(new_n275_), .A2(new_n273_), .ZN(new_n318_));
  NAND4_X1   g0055(.A1(new_n272_), .A2(new_n318_), .A3(new_n276_), .A4(new_n279_), .ZN(new_n319_));
  NAND2_X1   g0056(.A1(new_n288_), .A2(new_n286_), .ZN(new_n320_));
  INV_X1     g0057(.I(\a[122] ), .ZN(new_n321_));
  INV_X1     g0058(.I(\a[124] ), .ZN(new_n322_));
  NOR2_X1    g0059(.A1(\shift[2] ), .A2(\shift[3] ), .ZN(new_n323_));
  NOR3_X1    g0060(.A1(new_n323_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n324_));
  NAND3_X1   g0061(.A1(new_n285_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1     g0062(.I(\a[0] ), .ZN(new_n326_));
  NAND3_X1   g0063(.A1(new_n326_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n327_));
  NAND2_X1   g0064(.A1(new_n327_), .A2(new_n297_), .ZN(new_n328_));
  NAND4_X1   g0065(.A1(new_n296_), .A2(new_n328_), .A3(new_n276_), .A4(new_n303_), .ZN(new_n329_));
  INV_X1     g0066(.I(\a[115] ), .ZN(new_n330_));
  NAND3_X1   g0067(.A1(new_n330_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n331_));
  NAND2_X1   g0068(.A1(new_n331_), .A2(new_n310_), .ZN(new_n332_));
  AND2_X2    g0069(.A1(\a[114] ), .A2(\a[116] ), .Z(new_n333_));
  NAND4_X1   g0070(.A1(new_n309_), .A2(new_n332_), .A3(new_n276_), .A4(new_n333_), .ZN(new_n334_));
  NOR4_X1    g0071(.A1(new_n319_), .A2(new_n325_), .A3(new_n329_), .A4(new_n334_), .ZN(new_n335_));
  NOR3_X1    g0072(.A1(new_n335_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n336_));
  NOR2_X1    g0073(.A1(new_n336_), .A2(new_n317_), .ZN(new_n337_));
  NAND3_X1   g0074(.A1(\a[69] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n338_));
  NOR2_X1    g0075(.A1(new_n269_), .A2(\a[69] ), .ZN(new_n339_));
  NAND2_X1   g0076(.A1(new_n339_), .A2(new_n268_), .ZN(new_n340_));
  NAND2_X1   g0077(.A1(new_n340_), .A2(new_n338_), .ZN(new_n341_));
  INV_X1     g0078(.I(\a[71] ), .ZN(new_n342_));
  NOR3_X1    g0079(.A1(new_n342_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n343_));
  NOR3_X1    g0080(.A1(new_n294_), .A2(\a[71] ), .A3(\shift[1] ), .ZN(new_n344_));
  NOR2_X1    g0081(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1   g0082(.A1(new_n276_), .A2(\a[70] ), .A3(\a[72] ), .ZN(new_n346_));
  NOR2_X1    g0083(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1   g0084(.A1(\a[73] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n348_));
  NOR2_X1    g0085(.A1(new_n269_), .A2(\a[73] ), .ZN(new_n349_));
  NAND2_X1   g0086(.A1(new_n349_), .A2(new_n268_), .ZN(new_n350_));
  NAND2_X1   g0087(.A1(new_n350_), .A2(new_n348_), .ZN(new_n351_));
  NAND3_X1   g0088(.A1(\a[75] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n352_));
  INV_X1     g0089(.I(new_n352_), .ZN(new_n353_));
  NOR3_X1    g0090(.A1(new_n294_), .A2(\a[75] ), .A3(\shift[1] ), .ZN(new_n354_));
  NOR2_X1    g0091(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1     g0092(.I(\a[74] ), .ZN(new_n356_));
  INV_X1     g0093(.I(\a[76] ), .ZN(new_n357_));
  NOR2_X1    g0094(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1   g0095(.A1(new_n358_), .A2(new_n276_), .ZN(new_n359_));
  NOR2_X1    g0096(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1   g0097(.A1(new_n347_), .A2(new_n360_), .A3(new_n341_), .A4(new_n351_), .ZN(new_n361_));
  NAND3_X1   g0098(.A1(\a[77] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n362_));
  NOR2_X1    g0099(.A1(new_n269_), .A2(\a[77] ), .ZN(new_n363_));
  NAND2_X1   g0100(.A1(new_n363_), .A2(new_n268_), .ZN(new_n364_));
  NAND2_X1   g0101(.A1(new_n364_), .A2(new_n362_), .ZN(new_n365_));
  NAND3_X1   g0102(.A1(\a[79] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n366_));
  INV_X1     g0103(.I(new_n366_), .ZN(new_n367_));
  NOR3_X1    g0104(.A1(new_n294_), .A2(\a[79] ), .A3(\shift[1] ), .ZN(new_n368_));
  NOR2_X1    g0105(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1   g0106(.A1(new_n276_), .A2(\a[78] ), .A3(\a[80] ), .ZN(new_n370_));
  NOR2_X1    g0107(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1   g0108(.A1(\a[65] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n372_));
  NOR2_X1    g0109(.A1(new_n269_), .A2(\a[65] ), .ZN(new_n373_));
  NAND2_X1   g0110(.A1(new_n373_), .A2(new_n268_), .ZN(new_n374_));
  NAND2_X1   g0111(.A1(new_n374_), .A2(new_n372_), .ZN(new_n375_));
  NAND3_X1   g0112(.A1(\a[67] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n376_));
  INV_X1     g0113(.I(\a[67] ), .ZN(new_n377_));
  NAND3_X1   g0114(.A1(new_n377_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n378_));
  NAND3_X1   g0115(.A1(new_n276_), .A2(\a[66] ), .A3(\a[68] ), .ZN(new_n379_));
  AOI21_X1   g0116(.A1(new_n376_), .A2(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND4_X1   g0117(.A1(new_n380_), .A2(new_n371_), .A3(new_n365_), .A4(new_n375_), .ZN(new_n381_));
  NOR4_X1    g0118(.A1(new_n381_), .A2(new_n361_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n382_));
  NOR2_X1    g0119(.A1(new_n381_), .A2(new_n361_), .ZN(new_n383_));
  NOR3_X1    g0120(.A1(new_n383_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n384_));
  NAND3_X1   g0121(.A1(\a[85] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n385_));
  NOR2_X1    g0122(.A1(new_n269_), .A2(\a[85] ), .ZN(new_n386_));
  NAND2_X1   g0123(.A1(new_n386_), .A2(new_n268_), .ZN(new_n387_));
  NAND2_X1   g0124(.A1(new_n387_), .A2(new_n385_), .ZN(new_n388_));
  NAND3_X1   g0125(.A1(\a[87] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n389_));
  INV_X1     g0126(.I(\a[87] ), .ZN(new_n390_));
  NAND3_X1   g0127(.A1(new_n390_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n391_));
  NAND3_X1   g0128(.A1(new_n276_), .A2(\a[86] ), .A3(\a[88] ), .ZN(new_n392_));
  AOI21_X1   g0129(.A1(new_n389_), .A2(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND3_X1   g0130(.A1(\a[89] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n394_));
  INV_X1     g0131(.I(\a[89] ), .ZN(new_n395_));
  NAND3_X1   g0132(.A1(new_n395_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n396_));
  NAND2_X1   g0133(.A1(new_n396_), .A2(new_n394_), .ZN(new_n397_));
  NAND3_X1   g0134(.A1(\a[91] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n398_));
  INV_X1     g0135(.I(\a[91] ), .ZN(new_n399_));
  NAND3_X1   g0136(.A1(new_n399_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n400_));
  INV_X1     g0137(.I(\a[90] ), .ZN(new_n401_));
  INV_X1     g0138(.I(\a[92] ), .ZN(new_n402_));
  NOR2_X1    g0139(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1   g0140(.A1(new_n403_), .A2(new_n276_), .ZN(new_n404_));
  AOI21_X1   g0141(.A1(new_n398_), .A2(new_n400_), .B(new_n404_), .ZN(new_n405_));
  NAND4_X1   g0142(.A1(new_n405_), .A2(new_n393_), .A3(new_n388_), .A4(new_n397_), .ZN(new_n406_));
  NAND3_X1   g0143(.A1(\a[93] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n407_));
  NOR2_X1    g0144(.A1(new_n269_), .A2(\a[93] ), .ZN(new_n408_));
  NAND2_X1   g0145(.A1(new_n408_), .A2(new_n268_), .ZN(new_n409_));
  NAND2_X1   g0146(.A1(new_n409_), .A2(new_n407_), .ZN(new_n410_));
  INV_X1     g0147(.I(\a[95] ), .ZN(new_n411_));
  NOR3_X1    g0148(.A1(new_n411_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n412_));
  NOR3_X1    g0149(.A1(new_n294_), .A2(\a[95] ), .A3(\shift[1] ), .ZN(new_n413_));
  NOR2_X1    g0150(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1   g0151(.A1(new_n276_), .A2(\a[94] ), .A3(\a[96] ), .ZN(new_n415_));
  NOR2_X1    g0152(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1   g0153(.A1(\a[81] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n417_));
  INV_X1     g0154(.I(\a[81] ), .ZN(new_n418_));
  NAND3_X1   g0155(.A1(new_n418_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n419_));
  NAND2_X1   g0156(.A1(new_n419_), .A2(new_n417_), .ZN(new_n420_));
  NAND3_X1   g0157(.A1(\a[83] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n421_));
  INV_X1     g0158(.I(\a[83] ), .ZN(new_n422_));
  NAND3_X1   g0159(.A1(new_n422_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n423_));
  INV_X1     g0160(.I(\a[82] ), .ZN(new_n424_));
  INV_X1     g0161(.I(\a[84] ), .ZN(new_n425_));
  NOR2_X1    g0162(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1   g0163(.A1(new_n426_), .A2(new_n276_), .ZN(new_n427_));
  AOI21_X1   g0164(.A1(new_n421_), .A2(new_n423_), .B(new_n427_), .ZN(new_n428_));
  NAND4_X1   g0165(.A1(new_n428_), .A2(new_n416_), .A3(new_n410_), .A4(new_n420_), .ZN(new_n429_));
  NAND3_X1   g0166(.A1(\a[101] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n430_));
  NOR2_X1    g0167(.A1(new_n269_), .A2(\a[101] ), .ZN(new_n431_));
  NAND2_X1   g0168(.A1(new_n431_), .A2(new_n268_), .ZN(new_n432_));
  NAND2_X1   g0169(.A1(new_n432_), .A2(new_n430_), .ZN(new_n433_));
  NAND3_X1   g0170(.A1(\a[103] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n434_));
  INV_X1     g0171(.I(\a[103] ), .ZN(new_n435_));
  NAND3_X1   g0172(.A1(new_n435_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n436_));
  INV_X1     g0173(.I(\a[102] ), .ZN(new_n437_));
  INV_X1     g0174(.I(\a[104] ), .ZN(new_n438_));
  NOR2_X1    g0175(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1   g0176(.A1(new_n439_), .A2(new_n276_), .ZN(new_n440_));
  AOI21_X1   g0177(.A1(new_n434_), .A2(new_n436_), .B(new_n440_), .ZN(new_n441_));
  NAND3_X1   g0178(.A1(\a[105] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n442_));
  NOR2_X1    g0179(.A1(new_n269_), .A2(\a[105] ), .ZN(new_n443_));
  NAND2_X1   g0180(.A1(new_n443_), .A2(new_n268_), .ZN(new_n444_));
  NAND2_X1   g0181(.A1(new_n444_), .A2(new_n442_), .ZN(new_n445_));
  NAND3_X1   g0182(.A1(\a[107] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n446_));
  INV_X1     g0183(.I(new_n446_), .ZN(new_n447_));
  NOR3_X1    g0184(.A1(new_n294_), .A2(\a[107] ), .A3(\shift[1] ), .ZN(new_n448_));
  NOR2_X1    g0185(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1   g0186(.A1(new_n276_), .A2(\a[106] ), .A3(\a[108] ), .ZN(new_n450_));
  NOR2_X1    g0187(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1   g0188(.A1(new_n441_), .A2(new_n451_), .A3(new_n433_), .A4(new_n445_), .ZN(new_n452_));
  NAND3_X1   g0189(.A1(\a[109] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n453_));
  NOR2_X1    g0190(.A1(new_n269_), .A2(\a[109] ), .ZN(new_n454_));
  NAND2_X1   g0191(.A1(new_n454_), .A2(new_n268_), .ZN(new_n455_));
  NAND2_X1   g0192(.A1(new_n455_), .A2(new_n453_), .ZN(new_n456_));
  AND3_X2    g0193(.A1(\a[111] ), .A2(\shift[0] ), .A3(\shift[1] ), .Z(new_n457_));
  NOR3_X1    g0194(.A1(new_n294_), .A2(\a[111] ), .A3(\shift[1] ), .ZN(new_n458_));
  NOR2_X1    g0195(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1   g0196(.A1(new_n276_), .A2(\a[110] ), .A3(\a[112] ), .ZN(new_n460_));
  NOR2_X1    g0197(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1   g0198(.A1(\a[97] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n462_));
  INV_X1     g0199(.I(\a[97] ), .ZN(new_n463_));
  NAND3_X1   g0200(.A1(new_n463_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n464_));
  NAND2_X1   g0201(.A1(new_n464_), .A2(new_n462_), .ZN(new_n465_));
  NAND3_X1   g0202(.A1(\a[99] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n466_));
  INV_X1     g0203(.I(new_n466_), .ZN(new_n467_));
  NOR3_X1    g0204(.A1(new_n294_), .A2(\a[99] ), .A3(\shift[1] ), .ZN(new_n468_));
  NOR2_X1    g0205(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1     g0206(.I(\a[98] ), .ZN(new_n470_));
  INV_X1     g0207(.I(\a[100] ), .ZN(new_n471_));
  NOR2_X1    g0208(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1   g0209(.A1(new_n472_), .A2(new_n276_), .ZN(new_n473_));
  NOR2_X1    g0210(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1   g0211(.A1(new_n474_), .A2(new_n461_), .A3(new_n456_), .A4(new_n465_), .ZN(new_n475_));
  NOR4_X1    g0212(.A1(new_n406_), .A2(new_n452_), .A3(new_n429_), .A4(new_n475_), .ZN(new_n476_));
  OAI21_X1   g0213(.A1(new_n384_), .A2(new_n382_), .B(new_n476_), .ZN(new_n477_));
  OAI21_X1   g0214(.A1(new_n477_), .A2(new_n337_), .B(new_n264_), .ZN(new_n478_));
  NAND3_X1   g0215(.A1(\a[53] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n479_));
  NOR2_X1    g0216(.A1(new_n269_), .A2(\a[53] ), .ZN(new_n480_));
  NAND2_X1   g0217(.A1(new_n480_), .A2(new_n268_), .ZN(new_n481_));
  NAND2_X1   g0218(.A1(new_n481_), .A2(new_n479_), .ZN(new_n482_));
  INV_X1     g0219(.I(\a[55] ), .ZN(new_n483_));
  NOR3_X1    g0220(.A1(new_n483_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n484_));
  NOR3_X1    g0221(.A1(new_n294_), .A2(\a[55] ), .A3(\shift[1] ), .ZN(new_n485_));
  NOR2_X1    g0222(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1   g0223(.A1(\a[54] ), .A2(\a[56] ), .ZN(new_n487_));
  NOR3_X1    g0224(.A1(new_n486_), .A2(new_n323_), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1   g0225(.A1(\a[57] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n489_));
  NOR2_X1    g0226(.A1(new_n269_), .A2(\a[57] ), .ZN(new_n490_));
  NAND2_X1   g0227(.A1(new_n490_), .A2(new_n268_), .ZN(new_n491_));
  NAND2_X1   g0228(.A1(new_n491_), .A2(new_n489_), .ZN(new_n492_));
  NAND3_X1   g0229(.A1(\a[59] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n493_));
  INV_X1     g0230(.I(\a[59] ), .ZN(new_n494_));
  NAND3_X1   g0231(.A1(new_n494_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n495_));
  NAND3_X1   g0232(.A1(new_n276_), .A2(\a[58] ), .A3(\a[60] ), .ZN(new_n496_));
  AOI21_X1   g0233(.A1(new_n493_), .A2(new_n495_), .B(new_n496_), .ZN(new_n497_));
  NAND4_X1   g0234(.A1(new_n488_), .A2(new_n497_), .A3(new_n482_), .A4(new_n492_), .ZN(new_n498_));
  NAND3_X1   g0235(.A1(\a[61] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n499_));
  NOR2_X1    g0236(.A1(new_n269_), .A2(\a[61] ), .ZN(new_n500_));
  NAND2_X1   g0237(.A1(new_n500_), .A2(new_n268_), .ZN(new_n501_));
  NAND2_X1   g0238(.A1(new_n501_), .A2(new_n499_), .ZN(new_n502_));
  NAND3_X1   g0239(.A1(\a[63] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n503_));
  INV_X1     g0240(.I(new_n503_), .ZN(new_n504_));
  NOR3_X1    g0241(.A1(new_n294_), .A2(\a[63] ), .A3(\shift[1] ), .ZN(new_n505_));
  NOR2_X1    g0242(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1   g0243(.A1(new_n276_), .A2(\a[62] ), .A3(\a[64] ), .ZN(new_n507_));
  NOR2_X1    g0244(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1   g0245(.A1(\a[49] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n509_));
  INV_X1     g0246(.I(new_n509_), .ZN(new_n510_));
  NOR3_X1    g0247(.A1(new_n269_), .A2(\a[49] ), .A3(\shift[0] ), .ZN(new_n511_));
  NOR2_X1    g0248(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1   g0249(.A1(\a[51] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n513_));
  INV_X1     g0250(.I(new_n513_), .ZN(new_n514_));
  NOR3_X1    g0251(.A1(new_n294_), .A2(\a[51] ), .A3(\shift[1] ), .ZN(new_n515_));
  NOR2_X1    g0252(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1     g0253(.I(\a[50] ), .ZN(new_n517_));
  INV_X1     g0254(.I(\a[52] ), .ZN(new_n518_));
  NOR3_X1    g0255(.A1(new_n323_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1     g0256(.I(new_n519_), .ZN(new_n520_));
  NOR3_X1    g0257(.A1(new_n512_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n521_));
  NAND3_X1   g0258(.A1(new_n521_), .A2(new_n502_), .A3(new_n508_), .ZN(new_n522_));
  NOR4_X1    g0259(.A1(new_n498_), .A2(new_n522_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n523_));
  INV_X1     g0260(.I(new_n486_), .ZN(new_n524_));
  NOR2_X1    g0261(.A1(new_n323_), .A2(new_n487_), .ZN(new_n525_));
  NAND3_X1   g0262(.A1(new_n524_), .A2(new_n482_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1   g0263(.A1(new_n495_), .A2(new_n493_), .ZN(new_n527_));
  INV_X1     g0264(.I(new_n496_), .ZN(new_n528_));
  NAND3_X1   g0265(.A1(new_n528_), .A2(new_n492_), .A3(new_n527_), .ZN(new_n529_));
  INV_X1     g0266(.I(\a[63] ), .ZN(new_n530_));
  NAND3_X1   g0267(.A1(new_n530_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n531_));
  NAND2_X1   g0268(.A1(new_n531_), .A2(new_n503_), .ZN(new_n532_));
  INV_X1     g0269(.I(\a[62] ), .ZN(new_n533_));
  INV_X1     g0270(.I(\a[64] ), .ZN(new_n534_));
  NOR3_X1    g0271(.A1(new_n323_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  NAND3_X1   g0272(.A1(new_n502_), .A2(new_n532_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1     g0273(.I(new_n511_), .ZN(new_n537_));
  NAND2_X1   g0274(.A1(new_n537_), .A2(new_n509_), .ZN(new_n538_));
  INV_X1     g0275(.I(\a[51] ), .ZN(new_n539_));
  NAND3_X1   g0276(.A1(new_n539_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n540_));
  NAND2_X1   g0277(.A1(new_n540_), .A2(new_n513_), .ZN(new_n541_));
  NAND3_X1   g0278(.A1(new_n538_), .A2(new_n541_), .A3(new_n519_), .ZN(new_n542_));
  NOR4_X1    g0279(.A1(new_n526_), .A2(new_n529_), .A3(new_n542_), .A4(new_n536_), .ZN(new_n543_));
  NOR3_X1    g0280(.A1(new_n543_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n544_));
  NOR2_X1    g0281(.A1(new_n544_), .A2(new_n523_), .ZN(new_n545_));
  NAND3_X1   g0282(.A1(\a[5] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n546_));
  NOR2_X1    g0283(.A1(new_n269_), .A2(\a[5] ), .ZN(new_n547_));
  NAND2_X1   g0284(.A1(new_n547_), .A2(new_n268_), .ZN(new_n548_));
  NAND2_X1   g0285(.A1(new_n548_), .A2(new_n546_), .ZN(new_n549_));
  NAND3_X1   g0286(.A1(\a[7] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n550_));
  INV_X1     g0287(.I(new_n550_), .ZN(new_n551_));
  NOR3_X1    g0288(.A1(new_n294_), .A2(\a[7] ), .A3(\shift[1] ), .ZN(new_n552_));
  NOR2_X1    g0289(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1     g0290(.I(\a[6] ), .ZN(new_n554_));
  INV_X1     g0291(.I(\a[8] ), .ZN(new_n555_));
  NOR2_X1    g0292(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1   g0293(.A1(new_n556_), .A2(new_n276_), .ZN(new_n557_));
  NOR2_X1    g0294(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1   g0295(.A1(\a[9] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n559_));
  INV_X1     g0296(.I(\a[9] ), .ZN(new_n560_));
  NAND3_X1   g0297(.A1(new_n560_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n561_));
  NAND2_X1   g0298(.A1(new_n561_), .A2(new_n559_), .ZN(new_n562_));
  NAND3_X1   g0299(.A1(\a[11] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n563_));
  INV_X1     g0300(.I(\a[11] ), .ZN(new_n564_));
  NAND3_X1   g0301(.A1(new_n564_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n565_));
  INV_X1     g0302(.I(\a[10] ), .ZN(new_n566_));
  INV_X1     g0303(.I(\a[12] ), .ZN(new_n567_));
  NOR2_X1    g0304(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1   g0305(.A1(new_n568_), .A2(new_n276_), .ZN(new_n569_));
  AOI21_X1   g0306(.A1(new_n563_), .A2(new_n565_), .B(new_n569_), .ZN(new_n570_));
  NAND4_X1   g0307(.A1(new_n570_), .A2(new_n558_), .A3(new_n549_), .A4(new_n562_), .ZN(new_n571_));
  NAND3_X1   g0308(.A1(\a[13] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n572_));
  NOR2_X1    g0309(.A1(new_n269_), .A2(\a[13] ), .ZN(new_n573_));
  NAND2_X1   g0310(.A1(new_n573_), .A2(new_n268_), .ZN(new_n574_));
  NAND2_X1   g0311(.A1(new_n574_), .A2(new_n572_), .ZN(new_n575_));
  INV_X1     g0312(.I(\a[15] ), .ZN(new_n576_));
  NOR3_X1    g0313(.A1(new_n576_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n577_));
  NOR3_X1    g0314(.A1(new_n294_), .A2(\a[15] ), .A3(\shift[1] ), .ZN(new_n578_));
  NOR2_X1    g0315(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1   g0316(.A1(new_n276_), .A2(\a[14] ), .A3(\a[16] ), .ZN(new_n580_));
  NOR2_X1    g0317(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1   g0318(.A1(\a[1] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n582_));
  INV_X1     g0319(.I(\a[1] ), .ZN(new_n583_));
  NAND3_X1   g0320(.A1(new_n583_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n584_));
  NAND2_X1   g0321(.A1(new_n584_), .A2(new_n582_), .ZN(new_n585_));
  AND3_X2    g0322(.A1(\a[3] ), .A2(\shift[0] ), .A3(\shift[1] ), .Z(new_n586_));
  NOR3_X1    g0323(.A1(new_n294_), .A2(\a[3] ), .A3(\shift[1] ), .ZN(new_n587_));
  NOR2_X1    g0324(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1     g0325(.I(\a[2] ), .ZN(new_n589_));
  INV_X1     g0326(.I(\a[4] ), .ZN(new_n590_));
  NOR2_X1    g0327(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1   g0328(.A1(new_n591_), .A2(new_n276_), .ZN(new_n592_));
  NOR2_X1    g0329(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  NAND4_X1   g0330(.A1(new_n581_), .A2(new_n593_), .A3(new_n575_), .A4(new_n585_), .ZN(new_n594_));
  NOR4_X1    g0331(.A1(new_n571_), .A2(new_n594_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n595_));
  NOR2_X1    g0332(.A1(new_n571_), .A2(new_n594_), .ZN(new_n596_));
  NOR3_X1    g0333(.A1(new_n596_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n597_));
  NAND3_X1   g0334(.A1(\a[21] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n598_));
  NOR2_X1    g0335(.A1(new_n269_), .A2(\a[21] ), .ZN(new_n599_));
  NAND2_X1   g0336(.A1(new_n599_), .A2(new_n268_), .ZN(new_n600_));
  NAND2_X1   g0337(.A1(new_n600_), .A2(new_n598_), .ZN(new_n601_));
  INV_X1     g0338(.I(\a[23] ), .ZN(new_n602_));
  NOR3_X1    g0339(.A1(new_n602_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n603_));
  NOR3_X1    g0340(.A1(new_n294_), .A2(\a[23] ), .A3(\shift[1] ), .ZN(new_n604_));
  NOR2_X1    g0341(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1   g0342(.A1(new_n276_), .A2(\a[22] ), .A3(\a[24] ), .ZN(new_n606_));
  NOR2_X1    g0343(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1   g0344(.A1(\a[25] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n608_));
  INV_X1     g0345(.I(new_n608_), .ZN(new_n609_));
  NOR3_X1    g0346(.A1(new_n269_), .A2(\a[25] ), .A3(\shift[0] ), .ZN(new_n610_));
  NOR2_X1    g0347(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1   g0348(.A1(\a[27] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n612_));
  INV_X1     g0349(.I(new_n612_), .ZN(new_n613_));
  NOR3_X1    g0350(.A1(new_n294_), .A2(\a[27] ), .A3(\shift[1] ), .ZN(new_n614_));
  NOR2_X1    g0351(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X2    g0352(.A1(\a[26] ), .A2(\a[28] ), .Z(new_n616_));
  NAND2_X1   g0353(.A1(new_n276_), .A2(new_n616_), .ZN(new_n617_));
  NOR3_X1    g0354(.A1(new_n611_), .A2(new_n615_), .A3(new_n617_), .ZN(new_n618_));
  NAND3_X1   g0355(.A1(new_n618_), .A2(new_n601_), .A3(new_n607_), .ZN(new_n619_));
  NAND3_X1   g0356(.A1(\a[29] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n620_));
  INV_X1     g0357(.I(new_n620_), .ZN(new_n621_));
  NOR3_X1    g0358(.A1(new_n269_), .A2(\a[29] ), .A3(\shift[0] ), .ZN(new_n622_));
  NOR2_X1    g0359(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1   g0360(.A1(\a[31] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n624_));
  INV_X1     g0361(.I(new_n624_), .ZN(new_n625_));
  NOR3_X1    g0362(.A1(new_n294_), .A2(\a[31] ), .A3(\shift[1] ), .ZN(new_n626_));
  NOR2_X1    g0363(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1   g0364(.A1(\a[30] ), .A2(\a[32] ), .ZN(new_n628_));
  NOR4_X1    g0365(.A1(new_n623_), .A2(new_n627_), .A3(new_n323_), .A4(new_n628_), .ZN(new_n629_));
  NAND3_X1   g0366(.A1(\a[17] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n630_));
  INV_X1     g0367(.I(\a[17] ), .ZN(new_n631_));
  NAND3_X1   g0368(.A1(new_n631_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n632_));
  NAND2_X1   g0369(.A1(new_n632_), .A2(new_n630_), .ZN(new_n633_));
  NAND3_X1   g0370(.A1(\a[19] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n634_));
  INV_X1     g0371(.I(\a[19] ), .ZN(new_n635_));
  NAND3_X1   g0372(.A1(new_n635_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n636_));
  NAND2_X1   g0373(.A1(new_n636_), .A2(new_n634_), .ZN(new_n637_));
  NAND2_X1   g0374(.A1(\a[18] ), .A2(\a[20] ), .ZN(new_n638_));
  NOR2_X1    g0375(.A1(new_n323_), .A2(new_n638_), .ZN(new_n639_));
  AND3_X2    g0376(.A1(new_n633_), .A2(new_n637_), .A3(new_n639_), .Z(new_n640_));
  NAND2_X1   g0377(.A1(new_n640_), .A2(new_n629_), .ZN(new_n641_));
  INV_X1     g0378(.I(\a[37] ), .ZN(new_n642_));
  NOR2_X1    g0379(.A1(new_n642_), .A2(new_n294_), .ZN(new_n643_));
  NOR4_X1    g0380(.A1(new_n643_), .A2(\a[40] ), .A3(\shift[0] ), .A4(new_n269_), .ZN(new_n644_));
  NOR2_X1    g0381(.A1(\a[40] ), .A2(\shift[0] ), .ZN(new_n645_));
  NOR4_X1    g0382(.A1(new_n645_), .A2(new_n642_), .A3(new_n294_), .A4(new_n269_), .ZN(new_n646_));
  INV_X1     g0383(.I(\a[39] ), .ZN(new_n647_));
  INV_X1     g0384(.I(\a[38] ), .ZN(new_n648_));
  NAND3_X1   g0385(.A1(new_n647_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n650_));
  NAND3_X1   g0386(.A1(\a[38] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n652_));
  AOI21_X1   g0387(.A1(new_n650_), .A2(new_n652_), .B(new_n323_), .ZN(new_n653_));
  OAI21_X1   g0388(.A1(new_n644_), .A2(new_n646_), .B(new_n653_), .ZN(new_n654_));
  NAND3_X1   g0389(.A1(\a[33] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n655_));
  INV_X1     g0390(.I(new_n655_), .ZN(new_n656_));
  NOR3_X1    g0391(.A1(new_n269_), .A2(\a[33] ), .A3(\shift[0] ), .ZN(new_n657_));
  NOR2_X1    g0392(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1   g0393(.A1(\a[35] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n659_));
  INV_X1     g0394(.I(new_n659_), .ZN(new_n660_));
  NOR3_X1    g0395(.A1(new_n294_), .A2(\a[35] ), .A3(\shift[1] ), .ZN(new_n661_));
  NOR2_X1    g0396(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1     g0397(.I(\a[34] ), .ZN(new_n663_));
  INV_X1     g0398(.I(\a[36] ), .ZN(new_n664_));
  NOR3_X1    g0399(.A1(new_n323_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1     g0400(.I(new_n665_), .ZN(new_n666_));
  NOR3_X1    g0401(.A1(new_n658_), .A2(new_n662_), .A3(new_n666_), .ZN(new_n667_));
  NAND3_X1   g0402(.A1(\a[41] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n668_));
  INV_X1     g0403(.I(new_n668_), .ZN(new_n669_));
  NOR3_X1    g0404(.A1(new_n269_), .A2(\a[41] ), .A3(\shift[0] ), .ZN(new_n670_));
  NOR2_X1    g0405(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1   g0406(.A1(\a[43] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n672_));
  INV_X1     g0407(.I(new_n672_), .ZN(new_n673_));
  NOR3_X1    g0408(.A1(new_n294_), .A2(\a[43] ), .A3(\shift[1] ), .ZN(new_n674_));
  NOR2_X1    g0409(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1     g0410(.I(\a[42] ), .ZN(new_n676_));
  INV_X1     g0411(.I(\a[44] ), .ZN(new_n677_));
  NOR2_X1    g0412(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1     g0413(.I(new_n678_), .ZN(new_n679_));
  NOR4_X1    g0414(.A1(new_n671_), .A2(new_n675_), .A3(new_n323_), .A4(new_n679_), .ZN(new_n680_));
  NAND3_X1   g0415(.A1(\a[45] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n681_));
  INV_X1     g0416(.I(new_n681_), .ZN(new_n682_));
  NOR3_X1    g0417(.A1(new_n269_), .A2(\a[45] ), .A3(\shift[0] ), .ZN(new_n683_));
  NOR2_X1    g0418(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1   g0419(.A1(\a[47] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n685_));
  INV_X1     g0420(.I(new_n685_), .ZN(new_n686_));
  NOR3_X1    g0421(.A1(new_n294_), .A2(\a[47] ), .A3(\shift[1] ), .ZN(new_n687_));
  NOR2_X1    g0422(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1     g0423(.I(\a[46] ), .ZN(new_n689_));
  INV_X1     g0424(.I(\a[48] ), .ZN(new_n690_));
  NOR2_X1    g0425(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1   g0426(.A1(new_n691_), .A2(new_n276_), .ZN(new_n692_));
  NOR3_X1    g0427(.A1(new_n684_), .A2(new_n688_), .A3(new_n692_), .ZN(new_n693_));
  NAND3_X1   g0428(.A1(new_n680_), .A2(new_n667_), .A3(new_n693_), .ZN(new_n694_));
  NOR4_X1    g0429(.A1(new_n694_), .A2(new_n641_), .A3(new_n619_), .A4(new_n654_), .ZN(new_n695_));
  OAI21_X1   g0430(.A1(new_n597_), .A2(new_n595_), .B(new_n695_), .ZN(new_n696_));
  OAI21_X1   g0431(.A1(new_n696_), .A2(new_n545_), .B(\shift[6] ), .ZN(new_n697_));
  NAND2_X1   g0432(.A1(new_n478_), .A2(new_n697_), .ZN(\result[0] ));
  INV_X1     g0433(.I(\a[121] ), .ZN(new_n699_));
  NAND2_X1   g0434(.A1(\a[118] ), .A2(\shift[0] ), .ZN(new_n700_));
  NAND4_X1   g0435(.A1(new_n700_), .A2(new_n699_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n701_));
  NAND3_X1   g0436(.A1(\a[118] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n702_));
  NAND2_X1   g0437(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1   g0438(.A1(new_n278_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n705_));
  NAND3_X1   g0439(.A1(\a[119] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n707_));
  AOI21_X1   g0440(.A1(new_n705_), .A2(new_n707_), .B(new_n323_), .ZN(new_n708_));
  NAND2_X1   g0441(.A1(\a[122] ), .A2(\shift[0] ), .ZN(new_n709_));
  NAND4_X1   g0442(.A1(new_n709_), .A2(new_n293_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n710_));
  NAND3_X1   g0443(.A1(\a[122] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n712_));
  NAND2_X1   g0444(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1   g0445(.A1(new_n322_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n715_));
  NAND3_X1   g0446(.A1(\a[123] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n717_));
  AOI21_X1   g0447(.A1(new_n715_), .A2(new_n717_), .B(new_n323_), .ZN(new_n718_));
  NAND4_X1   g0448(.A1(new_n703_), .A2(new_n713_), .A3(new_n708_), .A4(new_n718_), .ZN(new_n719_));
  NAND3_X1   g0449(.A1(\a[1] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n720_));
  NOR3_X1    g0450(.A1(new_n269_), .A2(\a[126] ), .A3(\shift[0] ), .ZN(new_n721_));
  NAND2_X1   g0451(.A1(new_n721_), .A2(new_n720_), .ZN(new_n722_));
  NAND2_X1   g0452(.A1(new_n301_), .A2(new_n294_), .ZN(new_n723_));
  NAND4_X1   g0453(.A1(new_n723_), .A2(\a[1] ), .A3(\shift[0] ), .A4(\shift[1] ), .ZN(new_n724_));
  NAND2_X1   g0454(.A1(new_n724_), .A2(new_n722_), .ZN(new_n725_));
  NAND3_X1   g0455(.A1(\a[0] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n726_));
  NOR3_X1    g0456(.A1(new_n269_), .A2(\a[127] ), .A3(\shift[0] ), .ZN(new_n727_));
  NAND2_X1   g0457(.A1(new_n727_), .A2(new_n726_), .ZN(new_n728_));
  INV_X1     g0458(.I(new_n726_), .ZN(new_n729_));
  NAND3_X1   g0459(.A1(new_n302_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n730_));
  NAND2_X1   g0460(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  AOI21_X1   g0461(.A1(new_n731_), .A2(new_n728_), .B(new_n323_), .ZN(new_n732_));
  INV_X1     g0462(.I(\a[117] ), .ZN(new_n733_));
  NAND2_X1   g0463(.A1(\a[114] ), .A2(\shift[0] ), .ZN(new_n734_));
  NAND4_X1   g0464(.A1(new_n734_), .A2(new_n733_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n735_));
  NAND3_X1   g0465(.A1(\a[114] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n736_));
  NAND2_X1   g0466(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1     g0467(.I(\a[116] ), .ZN(new_n738_));
  NAND3_X1   g0468(.A1(new_n738_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n740_));
  NAND3_X1   g0469(.A1(\a[115] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n742_));
  AOI21_X1   g0470(.A1(new_n740_), .A2(new_n742_), .B(new_n323_), .ZN(new_n743_));
  NAND4_X1   g0471(.A1(new_n732_), .A2(new_n725_), .A3(new_n737_), .A4(new_n743_), .ZN(new_n744_));
  NOR4_X1    g0472(.A1(new_n744_), .A2(new_n265_), .A3(new_n266_), .A4(new_n719_), .ZN(new_n745_));
  NOR2_X1    g0473(.A1(new_n744_), .A2(new_n719_), .ZN(new_n746_));
  NOR3_X1    g0474(.A1(new_n746_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n747_));
  NOR2_X1    g0475(.A1(new_n747_), .A2(new_n745_), .ZN(new_n748_));
  INV_X1     g0476(.I(\a[73] ), .ZN(new_n749_));
  NAND2_X1   g0477(.A1(\a[70] ), .A2(\shift[0] ), .ZN(new_n750_));
  NAND4_X1   g0478(.A1(new_n750_), .A2(new_n749_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n751_));
  NAND3_X1   g0479(.A1(\a[70] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n752_));
  NAND2_X1   g0480(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1     g0481(.I(\a[72] ), .ZN(new_n754_));
  NAND3_X1   g0482(.A1(new_n754_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n756_));
  NAND3_X1   g0483(.A1(\a[71] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n758_));
  AOI21_X1   g0484(.A1(new_n756_), .A2(new_n758_), .B(new_n323_), .ZN(new_n759_));
  INV_X1     g0485(.I(\a[77] ), .ZN(new_n760_));
  NAND2_X1   g0486(.A1(\a[74] ), .A2(\shift[0] ), .ZN(new_n761_));
  NAND4_X1   g0487(.A1(new_n761_), .A2(new_n760_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n762_));
  NAND3_X1   g0488(.A1(\a[74] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n763_));
  NAND2_X1   g0489(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1     g0490(.I(\a[75] ), .ZN(new_n765_));
  NAND3_X1   g0491(.A1(new_n357_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n767_));
  NAND3_X1   g0492(.A1(\a[75] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n769_));
  AOI21_X1   g0493(.A1(new_n767_), .A2(new_n769_), .B(new_n323_), .ZN(new_n770_));
  NAND4_X1   g0494(.A1(new_n753_), .A2(new_n764_), .A3(new_n759_), .A4(new_n770_), .ZN(new_n771_));
  NAND2_X1   g0495(.A1(\a[78] ), .A2(\shift[0] ), .ZN(new_n772_));
  NAND4_X1   g0496(.A1(new_n772_), .A2(new_n418_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n773_));
  NAND3_X1   g0497(.A1(\a[78] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n775_));
  NAND2_X1   g0498(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1     g0499(.I(\a[80] ), .ZN(new_n777_));
  INV_X1     g0500(.I(\a[79] ), .ZN(new_n778_));
  NAND3_X1   g0501(.A1(new_n777_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n780_));
  NAND3_X1   g0502(.A1(\a[79] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n782_));
  AOI21_X1   g0503(.A1(new_n780_), .A2(new_n782_), .B(new_n323_), .ZN(new_n783_));
  INV_X1     g0504(.I(\a[69] ), .ZN(new_n784_));
  NAND2_X1   g0505(.A1(\a[66] ), .A2(\shift[0] ), .ZN(new_n785_));
  NAND4_X1   g0506(.A1(new_n785_), .A2(new_n784_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n786_));
  NAND3_X1   g0507(.A1(\a[66] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n787_));
  NAND2_X1   g0508(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1     g0509(.I(\a[68] ), .ZN(new_n789_));
  NAND3_X1   g0510(.A1(new_n789_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n791_));
  NAND3_X1   g0511(.A1(\a[67] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n793_));
  AOI21_X1   g0512(.A1(new_n791_), .A2(new_n793_), .B(new_n323_), .ZN(new_n794_));
  NAND4_X1   g0513(.A1(new_n776_), .A2(new_n788_), .A3(new_n783_), .A4(new_n794_), .ZN(new_n795_));
  NOR4_X1    g0514(.A1(new_n771_), .A2(new_n795_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n796_));
  NOR2_X1    g0515(.A1(new_n771_), .A2(new_n795_), .ZN(new_n797_));
  NOR3_X1    g0516(.A1(new_n797_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n798_));
  NAND2_X1   g0517(.A1(\a[86] ), .A2(\shift[0] ), .ZN(new_n799_));
  NAND4_X1   g0518(.A1(new_n799_), .A2(new_n395_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n800_));
  NAND3_X1   g0519(.A1(\a[86] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n802_));
  NAND2_X1   g0520(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1     g0521(.I(\a[88] ), .ZN(new_n804_));
  NAND3_X1   g0522(.A1(new_n804_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n806_));
  NAND3_X1   g0523(.A1(\a[87] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n808_));
  AOI21_X1   g0524(.A1(new_n806_), .A2(new_n808_), .B(new_n323_), .ZN(new_n809_));
  INV_X1     g0525(.I(\a[93] ), .ZN(new_n810_));
  NAND2_X1   g0526(.A1(\a[90] ), .A2(\shift[0] ), .ZN(new_n811_));
  NAND4_X1   g0527(.A1(new_n811_), .A2(new_n810_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n812_));
  NAND3_X1   g0528(.A1(\a[90] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n813_));
  NAND2_X1   g0529(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1   g0530(.A1(new_n402_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n816_));
  NAND3_X1   g0531(.A1(\a[91] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n818_));
  AOI21_X1   g0532(.A1(new_n816_), .A2(new_n818_), .B(new_n323_), .ZN(new_n819_));
  NAND4_X1   g0533(.A1(new_n803_), .A2(new_n814_), .A3(new_n809_), .A4(new_n819_), .ZN(new_n820_));
  NAND2_X1   g0534(.A1(\a[94] ), .A2(\shift[0] ), .ZN(new_n821_));
  NAND4_X1   g0535(.A1(new_n821_), .A2(new_n463_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n822_));
  NAND3_X1   g0536(.A1(\a[94] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n824_));
  NAND2_X1   g0537(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1     g0538(.I(\a[96] ), .ZN(new_n826_));
  NAND3_X1   g0539(.A1(new_n826_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n828_));
  NAND3_X1   g0540(.A1(\a[95] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n830_));
  AOI21_X1   g0541(.A1(new_n828_), .A2(new_n830_), .B(new_n323_), .ZN(new_n831_));
  INV_X1     g0542(.I(\a[85] ), .ZN(new_n832_));
  NAND2_X1   g0543(.A1(\a[82] ), .A2(\shift[0] ), .ZN(new_n833_));
  NAND4_X1   g0544(.A1(new_n833_), .A2(new_n832_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n834_));
  NAND3_X1   g0545(.A1(\a[82] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n835_));
  NAND2_X1   g0546(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1   g0547(.A1(new_n425_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n838_));
  NAND3_X1   g0548(.A1(\a[83] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n840_));
  AOI21_X1   g0549(.A1(new_n838_), .A2(new_n840_), .B(new_n323_), .ZN(new_n841_));
  NAND4_X1   g0550(.A1(new_n825_), .A2(new_n836_), .A3(new_n831_), .A4(new_n841_), .ZN(new_n842_));
  INV_X1     g0551(.I(\a[105] ), .ZN(new_n843_));
  NAND2_X1   g0552(.A1(\a[102] ), .A2(\shift[0] ), .ZN(new_n844_));
  NAND4_X1   g0553(.A1(new_n844_), .A2(new_n843_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n845_));
  NAND3_X1   g0554(.A1(\a[102] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n846_));
  NAND2_X1   g0555(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1   g0556(.A1(new_n438_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n849_));
  NAND3_X1   g0557(.A1(\a[103] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n851_));
  AOI21_X1   g0558(.A1(new_n849_), .A2(new_n851_), .B(new_n323_), .ZN(new_n852_));
  INV_X1     g0559(.I(\a[109] ), .ZN(new_n853_));
  NAND2_X1   g0560(.A1(\a[106] ), .A2(\shift[0] ), .ZN(new_n854_));
  NAND4_X1   g0561(.A1(new_n854_), .A2(new_n853_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n855_));
  NAND3_X1   g0562(.A1(\a[106] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n856_));
  NAND2_X1   g0563(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1     g0564(.I(\a[108] ), .ZN(new_n858_));
  INV_X1     g0565(.I(\a[107] ), .ZN(new_n859_));
  NAND3_X1   g0566(.A1(new_n858_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n861_));
  NAND3_X1   g0567(.A1(\a[107] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n863_));
  AOI21_X1   g0568(.A1(new_n861_), .A2(new_n863_), .B(new_n323_), .ZN(new_n864_));
  NAND4_X1   g0569(.A1(new_n847_), .A2(new_n857_), .A3(new_n852_), .A4(new_n864_), .ZN(new_n865_));
  NAND2_X1   g0570(.A1(\a[110] ), .A2(\shift[0] ), .ZN(new_n866_));
  NAND4_X1   g0571(.A1(new_n866_), .A2(new_n307_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n867_));
  NAND3_X1   g0572(.A1(\a[110] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n869_));
  NAND2_X1   g0573(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1     g0574(.I(\a[112] ), .ZN(new_n871_));
  INV_X1     g0575(.I(\a[111] ), .ZN(new_n872_));
  NAND3_X1   g0576(.A1(new_n871_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n874_));
  NAND3_X1   g0577(.A1(\a[111] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n876_));
  AOI21_X1   g0578(.A1(new_n874_), .A2(new_n876_), .B(new_n323_), .ZN(new_n877_));
  INV_X1     g0579(.I(\a[101] ), .ZN(new_n878_));
  NAND2_X1   g0580(.A1(\a[98] ), .A2(\shift[0] ), .ZN(new_n879_));
  NAND4_X1   g0581(.A1(new_n879_), .A2(new_n878_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n880_));
  NAND3_X1   g0582(.A1(\a[98] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n881_));
  NAND2_X1   g0583(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1     g0584(.I(\a[99] ), .ZN(new_n883_));
  NAND3_X1   g0585(.A1(new_n471_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n885_));
  NAND3_X1   g0586(.A1(\a[99] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n887_));
  AOI21_X1   g0587(.A1(new_n885_), .A2(new_n887_), .B(new_n323_), .ZN(new_n888_));
  NAND4_X1   g0588(.A1(new_n870_), .A2(new_n882_), .A3(new_n877_), .A4(new_n888_), .ZN(new_n889_));
  NOR4_X1    g0589(.A1(new_n820_), .A2(new_n842_), .A3(new_n865_), .A4(new_n889_), .ZN(new_n890_));
  OAI21_X1   g0590(.A1(new_n798_), .A2(new_n796_), .B(new_n890_), .ZN(new_n891_));
  OAI21_X1   g0591(.A1(new_n748_), .A2(new_n891_), .B(new_n264_), .ZN(new_n892_));
  NAND2_X1   g0592(.A1(\shift[4] ), .A2(\shift[5] ), .ZN(new_n893_));
  INV_X1     g0593(.I(\a[57] ), .ZN(new_n894_));
  NAND2_X1   g0594(.A1(\a[54] ), .A2(\shift[0] ), .ZN(new_n895_));
  NAND4_X1   g0595(.A1(new_n895_), .A2(new_n894_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n896_));
  NAND3_X1   g0596(.A1(\a[54] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n897_));
  NAND2_X1   g0597(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1     g0598(.I(\a[56] ), .ZN(new_n899_));
  NAND3_X1   g0599(.A1(new_n899_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n901_));
  NAND3_X1   g0600(.A1(\a[55] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n903_));
  AOI21_X1   g0601(.A1(new_n901_), .A2(new_n903_), .B(new_n323_), .ZN(new_n904_));
  INV_X1     g0602(.I(\a[61] ), .ZN(new_n905_));
  NAND2_X1   g0603(.A1(\a[58] ), .A2(\shift[0] ), .ZN(new_n906_));
  NAND4_X1   g0604(.A1(new_n906_), .A2(new_n905_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n907_));
  NAND3_X1   g0605(.A1(\a[58] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n908_));
  NAND2_X1   g0606(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1     g0607(.I(\a[60] ), .ZN(new_n910_));
  NAND3_X1   g0608(.A1(new_n910_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n912_));
  NAND3_X1   g0609(.A1(\a[59] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n914_));
  AOI21_X1   g0610(.A1(new_n912_), .A2(new_n914_), .B(new_n323_), .ZN(new_n915_));
  NAND4_X1   g0611(.A1(new_n898_), .A2(new_n909_), .A3(new_n904_), .A4(new_n915_), .ZN(new_n916_));
  INV_X1     g0612(.I(\a[65] ), .ZN(new_n917_));
  NAND2_X1   g0613(.A1(\a[62] ), .A2(\shift[0] ), .ZN(new_n918_));
  NAND4_X1   g0614(.A1(new_n918_), .A2(new_n917_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n919_));
  NAND3_X1   g0615(.A1(\a[62] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n920_));
  NAND2_X1   g0616(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NAND3_X1   g0617(.A1(new_n534_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n923_));
  NAND3_X1   g0618(.A1(\a[63] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n925_));
  AOI21_X1   g0619(.A1(new_n923_), .A2(new_n925_), .B(new_n323_), .ZN(new_n926_));
  INV_X1     g0620(.I(\a[53] ), .ZN(new_n927_));
  NAND2_X1   g0621(.A1(\a[50] ), .A2(\shift[0] ), .ZN(new_n928_));
  NAND4_X1   g0622(.A1(new_n928_), .A2(new_n927_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n929_));
  NAND3_X1   g0623(.A1(\a[50] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n930_));
  NAND2_X1   g0624(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NAND3_X1   g0625(.A1(new_n518_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n933_));
  NAND3_X1   g0626(.A1(\a[51] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n935_));
  AOI21_X1   g0627(.A1(new_n933_), .A2(new_n935_), .B(new_n323_), .ZN(new_n936_));
  NAND4_X1   g0628(.A1(new_n921_), .A2(new_n931_), .A3(new_n926_), .A4(new_n936_), .ZN(new_n937_));
  NOR3_X1    g0629(.A1(new_n916_), .A2(new_n937_), .A3(new_n893_), .ZN(new_n938_));
  NAND2_X1   g0630(.A1(\a[6] ), .A2(\shift[0] ), .ZN(new_n939_));
  NAND4_X1   g0631(.A1(new_n939_), .A2(new_n560_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n940_));
  NAND3_X1   g0632(.A1(\a[6] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n942_));
  NAND2_X1   g0633(.A1(new_n940_), .A2(new_n942_), .ZN(new_n943_));
  INV_X1     g0634(.I(\a[7] ), .ZN(new_n944_));
  NAND3_X1   g0635(.A1(new_n555_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n946_));
  NAND3_X1   g0636(.A1(\a[7] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n948_));
  AOI21_X1   g0637(.A1(new_n946_), .A2(new_n948_), .B(new_n323_), .ZN(new_n949_));
  INV_X1     g0638(.I(\a[13] ), .ZN(new_n950_));
  NAND2_X1   g0639(.A1(\a[10] ), .A2(\shift[0] ), .ZN(new_n951_));
  NAND4_X1   g0640(.A1(new_n951_), .A2(new_n950_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n952_));
  NAND3_X1   g0641(.A1(\a[10] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n953_));
  NAND2_X1   g0642(.A1(new_n952_), .A2(new_n953_), .ZN(new_n954_));
  NAND3_X1   g0643(.A1(new_n567_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n956_));
  NAND3_X1   g0644(.A1(\a[11] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n958_));
  AOI21_X1   g0645(.A1(new_n956_), .A2(new_n958_), .B(new_n323_), .ZN(new_n959_));
  NAND4_X1   g0646(.A1(new_n943_), .A2(new_n954_), .A3(new_n949_), .A4(new_n959_), .ZN(new_n960_));
  NAND2_X1   g0647(.A1(\a[14] ), .A2(\shift[0] ), .ZN(new_n961_));
  NAND4_X1   g0648(.A1(new_n961_), .A2(new_n631_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n962_));
  NAND3_X1   g0649(.A1(\a[14] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n964_));
  NAND2_X1   g0650(.A1(new_n962_), .A2(new_n964_), .ZN(new_n965_));
  INV_X1     g0651(.I(\a[16] ), .ZN(new_n966_));
  NAND3_X1   g0652(.A1(new_n966_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n968_));
  NAND3_X1   g0653(.A1(\a[15] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n970_));
  AOI21_X1   g0654(.A1(new_n968_), .A2(new_n970_), .B(new_n323_), .ZN(new_n971_));
  INV_X1     g0655(.I(\a[5] ), .ZN(new_n972_));
  NAND2_X1   g0656(.A1(\a[2] ), .A2(\shift[0] ), .ZN(new_n973_));
  NAND4_X1   g0657(.A1(new_n973_), .A2(new_n972_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n974_));
  NAND3_X1   g0658(.A1(\a[2] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n975_));
  NAND2_X1   g0659(.A1(new_n974_), .A2(new_n975_), .ZN(new_n976_));
  INV_X1     g0660(.I(\a[3] ), .ZN(new_n977_));
  NAND3_X1   g0661(.A1(new_n590_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n979_));
  NAND3_X1   g0662(.A1(\a[3] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n981_));
  AOI21_X1   g0663(.A1(new_n979_), .A2(new_n981_), .B(new_n323_), .ZN(new_n982_));
  NAND4_X1   g0664(.A1(new_n965_), .A2(new_n976_), .A3(new_n971_), .A4(new_n982_), .ZN(new_n983_));
  NOR2_X1    g0665(.A1(new_n266_), .A2(\shift[4] ), .ZN(new_n984_));
  OAI21_X1   g0666(.A1(new_n960_), .A2(new_n983_), .B(new_n984_), .ZN(new_n985_));
  XOR2_X1    g0667(.A1(new_n985_), .A2(new_n938_), .Z(new_n986_));
  INV_X1     g0668(.I(new_n893_), .ZN(new_n987_));
  NAND3_X1   g0669(.A1(\a[34] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n988_));
  NOR2_X1    g0670(.A1(\a[37] ), .A2(\shift[0] ), .ZN(new_n989_));
  AND3_X2    g0671(.A1(new_n988_), .A2(\shift[1] ), .A3(new_n989_), .Z(new_n990_));
  AOI21_X1   g0672(.A1(\shift[1] ), .A2(new_n989_), .B(new_n988_), .ZN(new_n991_));
  INV_X1     g0673(.I(\a[35] ), .ZN(new_n992_));
  NAND3_X1   g0674(.A1(new_n664_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n994_));
  NAND3_X1   g0675(.A1(\a[35] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n996_));
  AOI21_X1   g0676(.A1(new_n994_), .A2(new_n996_), .B(new_n323_), .ZN(new_n997_));
  OAI21_X1   g0677(.A1(new_n990_), .A2(new_n991_), .B(new_n997_), .ZN(new_n998_));
  INV_X1     g0678(.I(\a[49] ), .ZN(new_n999_));
  NAND2_X1   g0679(.A1(\a[46] ), .A2(\shift[0] ), .ZN(new_n1000_));
  NAND4_X1   g0680(.A1(new_n1000_), .A2(new_n999_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1001_));
  NAND3_X1   g0681(.A1(\a[46] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1003_));
  NAND2_X1   g0682(.A1(new_n1001_), .A2(new_n1003_), .ZN(new_n1004_));
  INV_X1     g0683(.I(\a[47] ), .ZN(new_n1005_));
  NAND3_X1   g0684(.A1(new_n690_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1007_));
  NAND3_X1   g0685(.A1(\a[47] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1009_));
  AOI21_X1   g0686(.A1(new_n1007_), .A2(new_n1009_), .B(new_n323_), .ZN(new_n1010_));
  NAND2_X1   g0687(.A1(new_n1004_), .A2(new_n1010_), .ZN(new_n1011_));
  NAND3_X1   g0688(.A1(\a[40] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1012_));
  INV_X1     g0689(.I(\a[40] ), .ZN(new_n1013_));
  NAND3_X1   g0690(.A1(new_n1013_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1014_));
  NAND2_X1   g0691(.A1(new_n1014_), .A2(new_n1012_), .ZN(new_n1015_));
  NAND3_X1   g0692(.A1(\a[38] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1016_));
  NAND3_X1   g0693(.A1(new_n648_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n1017_));
  NAND2_X1   g0694(.A1(new_n1017_), .A2(new_n1016_), .ZN(new_n1018_));
  INV_X1     g0695(.I(\a[41] ), .ZN(new_n1019_));
  NOR3_X1    g0696(.A1(new_n323_), .A2(new_n647_), .A3(new_n1019_), .ZN(new_n1020_));
  NAND3_X1   g0697(.A1(new_n1015_), .A2(new_n1018_), .A3(new_n1020_), .ZN(new_n1021_));
  NAND3_X1   g0698(.A1(\a[42] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1022_));
  NAND3_X1   g0699(.A1(new_n676_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n1023_));
  NAND2_X1   g0700(.A1(new_n1023_), .A2(new_n1022_), .ZN(new_n1024_));
  NAND3_X1   g0701(.A1(\a[44] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1025_));
  NAND3_X1   g0702(.A1(new_n677_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1026_));
  NAND2_X1   g0703(.A1(new_n1026_), .A2(new_n1025_), .ZN(new_n1027_));
  INV_X1     g0704(.I(\a[43] ), .ZN(new_n1028_));
  INV_X1     g0705(.I(\a[45] ), .ZN(new_n1029_));
  NOR2_X1    g0706(.A1(new_n1028_), .A2(new_n1029_), .ZN(new_n1030_));
  NAND4_X1   g0707(.A1(new_n1024_), .A2(new_n1027_), .A3(new_n276_), .A4(new_n1030_), .ZN(new_n1031_));
  NOR4_X1    g0708(.A1(new_n998_), .A2(new_n1031_), .A3(new_n1011_), .A4(new_n1021_), .ZN(new_n1032_));
  INV_X1     g0709(.I(\a[25] ), .ZN(new_n1033_));
  NAND2_X1   g0710(.A1(\a[22] ), .A2(\shift[0] ), .ZN(new_n1034_));
  NAND4_X1   g0711(.A1(new_n1034_), .A2(new_n1033_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1035_));
  NAND3_X1   g0712(.A1(\a[22] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1037_));
  NAND2_X1   g0713(.A1(new_n1035_), .A2(new_n1037_), .ZN(new_n1038_));
  INV_X1     g0714(.I(\a[24] ), .ZN(new_n1039_));
  NAND3_X1   g0715(.A1(new_n1039_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1041_));
  NAND3_X1   g0716(.A1(\a[23] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1043_));
  AOI21_X1   g0717(.A1(new_n1041_), .A2(new_n1043_), .B(new_n323_), .ZN(new_n1044_));
  INV_X1     g0718(.I(\a[29] ), .ZN(new_n1045_));
  NAND2_X1   g0719(.A1(\a[26] ), .A2(\shift[0] ), .ZN(new_n1046_));
  NAND4_X1   g0720(.A1(new_n1046_), .A2(new_n1045_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1047_));
  NAND3_X1   g0721(.A1(\a[26] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1049_));
  NAND2_X1   g0722(.A1(new_n1047_), .A2(new_n1049_), .ZN(new_n1050_));
  INV_X1     g0723(.I(\a[28] ), .ZN(new_n1051_));
  INV_X1     g0724(.I(\a[27] ), .ZN(new_n1052_));
  NAND3_X1   g0725(.A1(new_n1051_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1054_));
  NAND3_X1   g0726(.A1(\a[27] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1056_));
  AOI21_X1   g0727(.A1(new_n1054_), .A2(new_n1056_), .B(new_n323_), .ZN(new_n1057_));
  NAND4_X1   g0728(.A1(new_n1038_), .A2(new_n1050_), .A3(new_n1044_), .A4(new_n1057_), .ZN(new_n1058_));
  INV_X1     g0729(.I(\a[33] ), .ZN(new_n1059_));
  NAND2_X1   g0730(.A1(\a[30] ), .A2(\shift[0] ), .ZN(new_n1060_));
  NAND4_X1   g0731(.A1(new_n1060_), .A2(new_n1059_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1061_));
  NAND3_X1   g0732(.A1(\a[30] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1063_));
  NAND2_X1   g0733(.A1(new_n1061_), .A2(new_n1063_), .ZN(new_n1064_));
  INV_X1     g0734(.I(\a[32] ), .ZN(new_n1065_));
  INV_X1     g0735(.I(\a[31] ), .ZN(new_n1066_));
  NAND3_X1   g0736(.A1(new_n1065_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1068_));
  NAND3_X1   g0737(.A1(\a[31] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1070_));
  AOI21_X1   g0738(.A1(new_n1068_), .A2(new_n1070_), .B(new_n323_), .ZN(new_n1071_));
  INV_X1     g0739(.I(\a[21] ), .ZN(new_n1072_));
  NAND2_X1   g0740(.A1(\a[18] ), .A2(\shift[0] ), .ZN(new_n1073_));
  NAND4_X1   g0741(.A1(new_n1073_), .A2(new_n1072_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1074_));
  NAND3_X1   g0742(.A1(\a[18] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1075_));
  NAND2_X1   g0743(.A1(new_n1074_), .A2(new_n1075_), .ZN(new_n1076_));
  INV_X1     g0744(.I(\a[20] ), .ZN(new_n1077_));
  NAND3_X1   g0745(.A1(new_n1077_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1079_));
  NAND3_X1   g0746(.A1(\a[19] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1081_));
  AOI21_X1   g0747(.A1(new_n1079_), .A2(new_n1081_), .B(new_n323_), .ZN(new_n1082_));
  NAND4_X1   g0748(.A1(new_n1064_), .A2(new_n1076_), .A3(new_n1071_), .A4(new_n1082_), .ZN(new_n1083_));
  OAI21_X1   g0749(.A1(new_n1058_), .A2(new_n1083_), .B(new_n984_), .ZN(new_n1084_));
  AOI21_X1   g0750(.A1(new_n987_), .A2(new_n1032_), .B(new_n1084_), .ZN(new_n1085_));
  AND3_X2    g0751(.A1(new_n1084_), .A2(new_n987_), .A3(new_n1032_), .Z(new_n1086_));
  NOR2_X1    g0752(.A1(new_n1086_), .A2(new_n1085_), .ZN(new_n1087_));
  OAI21_X1   g0753(.A1(new_n1087_), .A2(new_n986_), .B(\shift[6] ), .ZN(new_n1088_));
  NAND2_X1   g0754(.A1(new_n1088_), .A2(new_n892_), .ZN(\result[1] ));
  NAND3_X1   g0755(.A1(\a[121] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1090_));
  NAND3_X1   g0756(.A1(new_n699_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1091_));
  NAND2_X1   g0757(.A1(new_n1091_), .A2(new_n1090_), .ZN(new_n1092_));
  NAND3_X1   g0758(.A1(\a[119] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1093_));
  NOR2_X1    g0759(.A1(new_n269_), .A2(\a[119] ), .ZN(new_n1094_));
  NAND2_X1   g0760(.A1(new_n1094_), .A2(new_n268_), .ZN(new_n1095_));
  NOR2_X1    g0761(.A1(new_n278_), .A2(new_n321_), .ZN(new_n1096_));
  NAND2_X1   g0762(.A1(new_n1096_), .A2(new_n276_), .ZN(new_n1097_));
  AOI21_X1   g0763(.A1(new_n1093_), .A2(new_n1095_), .B(new_n1097_), .ZN(new_n1098_));
  NAND3_X1   g0764(.A1(\a[125] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1099_));
  NAND3_X1   g0765(.A1(new_n293_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1100_));
  NAND2_X1   g0766(.A1(new_n1100_), .A2(new_n1099_), .ZN(new_n1101_));
  NAND3_X1   g0767(.A1(\a[123] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1102_));
  INV_X1     g0768(.I(new_n1102_), .ZN(new_n1103_));
  NOR3_X1    g0769(.A1(new_n269_), .A2(\a[123] ), .A3(\shift[0] ), .ZN(new_n1104_));
  NOR2_X1    g0770(.A1(new_n1103_), .A2(new_n1104_), .ZN(new_n1105_));
  NAND3_X1   g0771(.A1(new_n276_), .A2(\a[124] ), .A3(\a[126] ), .ZN(new_n1106_));
  NOR2_X1    g0772(.A1(new_n1105_), .A2(new_n1106_), .ZN(new_n1107_));
  NAND4_X1   g0773(.A1(new_n1098_), .A2(new_n1107_), .A3(new_n1092_), .A4(new_n1101_), .ZN(new_n1108_));
  NAND3_X1   g0774(.A1(\a[1] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1109_));
  NAND3_X1   g0775(.A1(new_n583_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1110_));
  NAND2_X1   g0776(.A1(new_n1110_), .A2(new_n1109_), .ZN(new_n1111_));
  NAND3_X1   g0777(.A1(\a[0] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1112_));
  INV_X1     g0778(.I(new_n1112_), .ZN(new_n1113_));
  NOR3_X1    g0779(.A1(new_n269_), .A2(\a[0] ), .A3(\shift[0] ), .ZN(new_n1114_));
  NOR2_X1    g0780(.A1(new_n1113_), .A2(new_n1114_), .ZN(new_n1115_));
  NOR2_X1    g0781(.A1(new_n589_), .A2(new_n302_), .ZN(new_n1116_));
  NAND2_X1   g0782(.A1(new_n1116_), .A2(new_n276_), .ZN(new_n1117_));
  NOR2_X1    g0783(.A1(new_n1115_), .A2(new_n1117_), .ZN(new_n1118_));
  NAND3_X1   g0784(.A1(\a[117] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1119_));
  NAND3_X1   g0785(.A1(new_n733_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1120_));
  NAND2_X1   g0786(.A1(new_n1120_), .A2(new_n1119_), .ZN(new_n1121_));
  NAND3_X1   g0787(.A1(\a[115] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1122_));
  INV_X1     g0788(.I(new_n1122_), .ZN(new_n1123_));
  NOR3_X1    g0789(.A1(new_n269_), .A2(\a[115] ), .A3(\shift[0] ), .ZN(new_n1124_));
  NOR2_X1    g0790(.A1(new_n1123_), .A2(new_n1124_), .ZN(new_n1125_));
  NOR2_X1    g0791(.A1(new_n738_), .A2(new_n277_), .ZN(new_n1126_));
  NAND2_X1   g0792(.A1(new_n1126_), .A2(new_n276_), .ZN(new_n1127_));
  NOR2_X1    g0793(.A1(new_n1125_), .A2(new_n1127_), .ZN(new_n1128_));
  NAND4_X1   g0794(.A1(new_n1118_), .A2(new_n1128_), .A3(new_n1111_), .A4(new_n1121_), .ZN(new_n1129_));
  NOR4_X1    g0795(.A1(new_n1108_), .A2(new_n1129_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1130_));
  NAND2_X1   g0796(.A1(new_n1095_), .A2(new_n1093_), .ZN(new_n1131_));
  NAND4_X1   g0797(.A1(new_n1131_), .A2(new_n276_), .A3(new_n1092_), .A4(new_n1096_), .ZN(new_n1132_));
  NAND2_X1   g0798(.A1(new_n1107_), .A2(new_n1101_), .ZN(new_n1133_));
  NAND3_X1   g0799(.A1(new_n326_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n1134_));
  NAND2_X1   g0800(.A1(new_n1134_), .A2(new_n1112_), .ZN(new_n1135_));
  NAND4_X1   g0801(.A1(new_n1111_), .A2(new_n1135_), .A3(new_n276_), .A4(new_n1116_), .ZN(new_n1136_));
  NAND3_X1   g0802(.A1(new_n330_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n1137_));
  NAND2_X1   g0803(.A1(new_n1137_), .A2(new_n1122_), .ZN(new_n1138_));
  NAND4_X1   g0804(.A1(new_n1121_), .A2(new_n1138_), .A3(new_n276_), .A4(new_n1126_), .ZN(new_n1139_));
  NOR4_X1    g0805(.A1(new_n1133_), .A2(new_n1132_), .A3(new_n1136_), .A4(new_n1139_), .ZN(new_n1140_));
  NOR3_X1    g0806(.A1(new_n1140_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1141_));
  NOR2_X1    g0807(.A1(new_n1141_), .A2(new_n1130_), .ZN(new_n1142_));
  NAND3_X1   g0808(.A1(\a[73] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1143_));
  NAND3_X1   g0809(.A1(new_n749_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1144_));
  NAND2_X1   g0810(.A1(new_n1144_), .A2(new_n1143_), .ZN(new_n1145_));
  NAND3_X1   g0811(.A1(\a[71] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1146_));
  NOR2_X1    g0812(.A1(new_n269_), .A2(\a[71] ), .ZN(new_n1147_));
  NAND2_X1   g0813(.A1(new_n1147_), .A2(new_n268_), .ZN(new_n1148_));
  NOR2_X1    g0814(.A1(new_n754_), .A2(new_n356_), .ZN(new_n1149_));
  NAND2_X1   g0815(.A1(new_n1149_), .A2(new_n276_), .ZN(new_n1150_));
  AOI21_X1   g0816(.A1(new_n1146_), .A2(new_n1148_), .B(new_n1150_), .ZN(new_n1151_));
  NAND3_X1   g0817(.A1(\a[77] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1152_));
  NAND3_X1   g0818(.A1(new_n760_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1153_));
  NAND2_X1   g0819(.A1(new_n1153_), .A2(new_n1152_), .ZN(new_n1154_));
  NAND3_X1   g0820(.A1(\a[75] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1155_));
  NOR2_X1    g0821(.A1(new_n269_), .A2(\a[75] ), .ZN(new_n1156_));
  NAND2_X1   g0822(.A1(new_n1156_), .A2(new_n268_), .ZN(new_n1157_));
  NAND3_X1   g0823(.A1(new_n276_), .A2(\a[76] ), .A3(\a[78] ), .ZN(new_n1158_));
  AOI21_X1   g0824(.A1(new_n1155_), .A2(new_n1157_), .B(new_n1158_), .ZN(new_n1159_));
  NAND4_X1   g0825(.A1(new_n1151_), .A2(new_n1159_), .A3(new_n1145_), .A4(new_n1154_), .ZN(new_n1160_));
  NAND3_X1   g0826(.A1(\a[81] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1161_));
  NAND3_X1   g0827(.A1(new_n418_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1162_));
  NAND2_X1   g0828(.A1(new_n1162_), .A2(new_n1161_), .ZN(new_n1163_));
  NAND3_X1   g0829(.A1(\a[79] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1164_));
  INV_X1     g0830(.I(new_n1164_), .ZN(new_n1165_));
  NOR3_X1    g0831(.A1(new_n269_), .A2(\a[79] ), .A3(\shift[0] ), .ZN(new_n1166_));
  NOR2_X1    g0832(.A1(new_n1165_), .A2(new_n1166_), .ZN(new_n1167_));
  NOR2_X1    g0833(.A1(new_n777_), .A2(new_n424_), .ZN(new_n1168_));
  NAND2_X1   g0834(.A1(new_n1168_), .A2(new_n276_), .ZN(new_n1169_));
  NOR2_X1    g0835(.A1(new_n1167_), .A2(new_n1169_), .ZN(new_n1170_));
  NAND3_X1   g0836(.A1(\a[69] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1171_));
  NAND3_X1   g0837(.A1(new_n784_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1172_));
  NAND2_X1   g0838(.A1(new_n1172_), .A2(new_n1171_), .ZN(new_n1173_));
  NAND3_X1   g0839(.A1(\a[67] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1174_));
  INV_X1     g0840(.I(new_n1174_), .ZN(new_n1175_));
  NOR3_X1    g0841(.A1(new_n269_), .A2(\a[67] ), .A3(\shift[0] ), .ZN(new_n1176_));
  NOR2_X1    g0842(.A1(new_n1175_), .A2(new_n1176_), .ZN(new_n1177_));
  INV_X1     g0843(.I(\a[70] ), .ZN(new_n1178_));
  NOR2_X1    g0844(.A1(new_n789_), .A2(new_n1178_), .ZN(new_n1179_));
  NAND2_X1   g0845(.A1(new_n1179_), .A2(new_n276_), .ZN(new_n1180_));
  NOR2_X1    g0846(.A1(new_n1177_), .A2(new_n1180_), .ZN(new_n1181_));
  NAND4_X1   g0847(.A1(new_n1170_), .A2(new_n1181_), .A3(new_n1163_), .A4(new_n1173_), .ZN(new_n1182_));
  NOR4_X1    g0848(.A1(new_n1160_), .A2(new_n1182_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1183_));
  NOR2_X1    g0849(.A1(new_n1160_), .A2(new_n1182_), .ZN(new_n1184_));
  NOR3_X1    g0850(.A1(new_n1184_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n1185_));
  NAND3_X1   g0851(.A1(\a[89] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1186_));
  NAND3_X1   g0852(.A1(new_n395_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1187_));
  NAND2_X1   g0853(.A1(new_n1187_), .A2(new_n1186_), .ZN(new_n1188_));
  NAND3_X1   g0854(.A1(\a[87] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1189_));
  NOR2_X1    g0855(.A1(new_n269_), .A2(\a[87] ), .ZN(new_n1190_));
  NAND2_X1   g0856(.A1(new_n1190_), .A2(new_n268_), .ZN(new_n1191_));
  NAND3_X1   g0857(.A1(new_n276_), .A2(\a[88] ), .A3(\a[90] ), .ZN(new_n1192_));
  AOI21_X1   g0858(.A1(new_n1189_), .A2(new_n1191_), .B(new_n1192_), .ZN(new_n1193_));
  NAND3_X1   g0859(.A1(\a[93] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1194_));
  NAND3_X1   g0860(.A1(new_n810_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1195_));
  NAND2_X1   g0861(.A1(new_n1195_), .A2(new_n1194_), .ZN(new_n1196_));
  NAND3_X1   g0862(.A1(\a[91] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1197_));
  NOR2_X1    g0863(.A1(new_n269_), .A2(\a[91] ), .ZN(new_n1198_));
  NAND2_X1   g0864(.A1(new_n1198_), .A2(new_n268_), .ZN(new_n1199_));
  AND2_X2    g0865(.A1(\a[92] ), .A2(\a[94] ), .Z(new_n1200_));
  NAND2_X1   g0866(.A1(new_n276_), .A2(new_n1200_), .ZN(new_n1201_));
  AOI21_X1   g0867(.A1(new_n1197_), .A2(new_n1199_), .B(new_n1201_), .ZN(new_n1202_));
  NAND4_X1   g0868(.A1(new_n1202_), .A2(new_n1193_), .A3(new_n1188_), .A4(new_n1196_), .ZN(new_n1203_));
  NAND3_X1   g0869(.A1(\a[97] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1204_));
  NAND3_X1   g0870(.A1(new_n463_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1205_));
  NAND2_X1   g0871(.A1(new_n1205_), .A2(new_n1204_), .ZN(new_n1206_));
  NAND3_X1   g0872(.A1(\a[95] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1207_));
  NOR2_X1    g0873(.A1(new_n269_), .A2(\a[95] ), .ZN(new_n1208_));
  NAND2_X1   g0874(.A1(new_n1208_), .A2(new_n268_), .ZN(new_n1209_));
  NOR2_X1    g0875(.A1(new_n826_), .A2(new_n470_), .ZN(new_n1210_));
  NAND2_X1   g0876(.A1(new_n1210_), .A2(new_n276_), .ZN(new_n1211_));
  AOI21_X1   g0877(.A1(new_n1207_), .A2(new_n1209_), .B(new_n1211_), .ZN(new_n1212_));
  NAND3_X1   g0878(.A1(\a[85] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1213_));
  NAND3_X1   g0879(.A1(new_n832_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1214_));
  NAND2_X1   g0880(.A1(new_n1214_), .A2(new_n1213_), .ZN(new_n1215_));
  NAND3_X1   g0881(.A1(\a[83] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1216_));
  INV_X1     g0882(.I(new_n1216_), .ZN(new_n1217_));
  NOR3_X1    g0883(.A1(new_n269_), .A2(\a[83] ), .A3(\shift[0] ), .ZN(new_n1218_));
  NOR2_X1    g0884(.A1(new_n1217_), .A2(new_n1218_), .ZN(new_n1219_));
  INV_X1     g0885(.I(\a[86] ), .ZN(new_n1220_));
  NOR2_X1    g0886(.A1(new_n425_), .A2(new_n1220_), .ZN(new_n1221_));
  NAND2_X1   g0887(.A1(new_n1221_), .A2(new_n276_), .ZN(new_n1222_));
  NOR2_X1    g0888(.A1(new_n1219_), .A2(new_n1222_), .ZN(new_n1223_));
  NAND4_X1   g0889(.A1(new_n1212_), .A2(new_n1223_), .A3(new_n1206_), .A4(new_n1215_), .ZN(new_n1224_));
  NAND3_X1   g0890(.A1(\a[105] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1225_));
  NAND3_X1   g0891(.A1(new_n843_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1226_));
  NAND2_X1   g0892(.A1(new_n1226_), .A2(new_n1225_), .ZN(new_n1227_));
  NAND3_X1   g0893(.A1(\a[103] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1228_));
  NOR2_X1    g0894(.A1(new_n269_), .A2(\a[103] ), .ZN(new_n1229_));
  NAND2_X1   g0895(.A1(new_n1229_), .A2(new_n268_), .ZN(new_n1230_));
  INV_X1     g0896(.I(\a[106] ), .ZN(new_n1231_));
  NOR2_X1    g0897(.A1(new_n438_), .A2(new_n1231_), .ZN(new_n1232_));
  NAND2_X1   g0898(.A1(new_n1232_), .A2(new_n276_), .ZN(new_n1233_));
  AOI21_X1   g0899(.A1(new_n1228_), .A2(new_n1230_), .B(new_n1233_), .ZN(new_n1234_));
  NAND3_X1   g0900(.A1(\a[109] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1235_));
  NAND3_X1   g0901(.A1(new_n853_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1236_));
  NAND2_X1   g0902(.A1(new_n1236_), .A2(new_n1235_), .ZN(new_n1237_));
  NOR3_X1    g0903(.A1(new_n859_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n1238_));
  NOR3_X1    g0904(.A1(new_n269_), .A2(\a[107] ), .A3(\shift[0] ), .ZN(new_n1239_));
  NOR2_X1    g0905(.A1(new_n1238_), .A2(new_n1239_), .ZN(new_n1240_));
  NAND3_X1   g0906(.A1(new_n276_), .A2(\a[108] ), .A3(\a[110] ), .ZN(new_n1241_));
  NOR2_X1    g0907(.A1(new_n1240_), .A2(new_n1241_), .ZN(new_n1242_));
  NAND4_X1   g0908(.A1(new_n1234_), .A2(new_n1242_), .A3(new_n1227_), .A4(new_n1237_), .ZN(new_n1243_));
  NAND3_X1   g0909(.A1(\a[113] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1244_));
  NAND3_X1   g0910(.A1(new_n307_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1245_));
  NAND2_X1   g0911(.A1(new_n1245_), .A2(new_n1244_), .ZN(new_n1246_));
  AND3_X2    g0912(.A1(\a[111] ), .A2(\shift[0] ), .A3(\shift[1] ), .Z(new_n1247_));
  NOR3_X1    g0913(.A1(new_n269_), .A2(\a[111] ), .A3(\shift[0] ), .ZN(new_n1248_));
  NOR2_X1    g0914(.A1(new_n1247_), .A2(new_n1248_), .ZN(new_n1249_));
  NAND3_X1   g0915(.A1(new_n276_), .A2(\a[112] ), .A3(\a[114] ), .ZN(new_n1250_));
  NOR2_X1    g0916(.A1(new_n1249_), .A2(new_n1250_), .ZN(new_n1251_));
  NAND3_X1   g0917(.A1(\a[101] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1252_));
  NAND3_X1   g0918(.A1(new_n878_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1253_));
  NAND2_X1   g0919(.A1(new_n1253_), .A2(new_n1252_), .ZN(new_n1254_));
  NAND3_X1   g0920(.A1(\a[99] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1255_));
  NOR2_X1    g0921(.A1(new_n269_), .A2(\a[99] ), .ZN(new_n1256_));
  NAND2_X1   g0922(.A1(new_n1256_), .A2(new_n268_), .ZN(new_n1257_));
  NOR2_X1    g0923(.A1(new_n471_), .A2(new_n437_), .ZN(new_n1258_));
  NAND2_X1   g0924(.A1(new_n1258_), .A2(new_n276_), .ZN(new_n1259_));
  AOI21_X1   g0925(.A1(new_n1255_), .A2(new_n1257_), .B(new_n1259_), .ZN(new_n1260_));
  NAND4_X1   g0926(.A1(new_n1260_), .A2(new_n1246_), .A3(new_n1251_), .A4(new_n1254_), .ZN(new_n1261_));
  NOR4_X1    g0927(.A1(new_n1203_), .A2(new_n1224_), .A3(new_n1243_), .A4(new_n1261_), .ZN(new_n1262_));
  OAI21_X1   g0928(.A1(new_n1185_), .A2(new_n1183_), .B(new_n1262_), .ZN(new_n1263_));
  OAI21_X1   g0929(.A1(new_n1263_), .A2(new_n1142_), .B(new_n264_), .ZN(new_n1264_));
  INV_X1     g0930(.I(new_n984_), .ZN(new_n1265_));
  NAND3_X1   g0931(.A1(\a[57] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1266_));
  NAND3_X1   g0932(.A1(new_n894_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1267_));
  NAND2_X1   g0933(.A1(new_n1267_), .A2(new_n1266_), .ZN(new_n1268_));
  NAND3_X1   g0934(.A1(\a[55] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1269_));
  NOR2_X1    g0935(.A1(new_n269_), .A2(\a[55] ), .ZN(new_n1270_));
  NAND2_X1   g0936(.A1(new_n1270_), .A2(new_n268_), .ZN(new_n1271_));
  AND2_X2    g0937(.A1(\a[56] ), .A2(\a[58] ), .Z(new_n1272_));
  NAND2_X1   g0938(.A1(new_n276_), .A2(new_n1272_), .ZN(new_n1273_));
  AOI21_X1   g0939(.A1(new_n1269_), .A2(new_n1271_), .B(new_n1273_), .ZN(new_n1274_));
  NAND3_X1   g0940(.A1(\a[61] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1275_));
  NAND3_X1   g0941(.A1(new_n905_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1276_));
  NAND2_X1   g0942(.A1(new_n1276_), .A2(new_n1275_), .ZN(new_n1277_));
  NAND3_X1   g0943(.A1(\a[59] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1278_));
  NOR2_X1    g0944(.A1(new_n269_), .A2(\a[59] ), .ZN(new_n1279_));
  NAND2_X1   g0945(.A1(new_n1279_), .A2(new_n268_), .ZN(new_n1280_));
  NOR2_X1    g0946(.A1(new_n910_), .A2(new_n533_), .ZN(new_n1281_));
  NAND2_X1   g0947(.A1(new_n1281_), .A2(new_n276_), .ZN(new_n1282_));
  AOI21_X1   g0948(.A1(new_n1278_), .A2(new_n1280_), .B(new_n1282_), .ZN(new_n1283_));
  NAND4_X1   g0949(.A1(new_n1283_), .A2(new_n1274_), .A3(new_n1268_), .A4(new_n1277_), .ZN(new_n1284_));
  NAND3_X1   g0950(.A1(\a[65] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1285_));
  NAND3_X1   g0951(.A1(new_n917_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1286_));
  NAND2_X1   g0952(.A1(new_n1286_), .A2(new_n1285_), .ZN(new_n1287_));
  NOR3_X1    g0953(.A1(new_n530_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n1288_));
  NOR3_X1    g0954(.A1(new_n269_), .A2(\a[63] ), .A3(\shift[0] ), .ZN(new_n1289_));
  NOR2_X1    g0955(.A1(new_n1288_), .A2(new_n1289_), .ZN(new_n1290_));
  NAND3_X1   g0956(.A1(new_n276_), .A2(\a[64] ), .A3(\a[66] ), .ZN(new_n1291_));
  NOR2_X1    g0957(.A1(new_n1290_), .A2(new_n1291_), .ZN(new_n1292_));
  NAND3_X1   g0958(.A1(\a[53] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1293_));
  NAND3_X1   g0959(.A1(new_n927_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1294_));
  NAND2_X1   g0960(.A1(new_n1294_), .A2(new_n1293_), .ZN(new_n1295_));
  NAND3_X1   g0961(.A1(\a[51] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1296_));
  INV_X1     g0962(.I(new_n1296_), .ZN(new_n1297_));
  NOR3_X1    g0963(.A1(new_n269_), .A2(\a[51] ), .A3(\shift[0] ), .ZN(new_n1298_));
  NOR2_X1    g0964(.A1(new_n1297_), .A2(new_n1298_), .ZN(new_n1299_));
  AND2_X2    g0965(.A1(\a[52] ), .A2(\a[54] ), .Z(new_n1300_));
  NAND2_X1   g0966(.A1(new_n276_), .A2(new_n1300_), .ZN(new_n1301_));
  NOR2_X1    g0967(.A1(new_n1299_), .A2(new_n1301_), .ZN(new_n1302_));
  NAND4_X1   g0968(.A1(new_n1292_), .A2(new_n1302_), .A3(new_n1287_), .A4(new_n1295_), .ZN(new_n1303_));
  NOR3_X1    g0969(.A1(new_n1284_), .A2(new_n1303_), .A3(new_n893_), .ZN(new_n1304_));
  NAND3_X1   g0970(.A1(\a[9] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1305_));
  NAND3_X1   g0971(.A1(new_n560_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1306_));
  NAND2_X1   g0972(.A1(new_n1306_), .A2(new_n1305_), .ZN(new_n1307_));
  NAND3_X1   g0973(.A1(\a[7] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1308_));
  NOR2_X1    g0974(.A1(new_n269_), .A2(\a[7] ), .ZN(new_n1309_));
  NAND2_X1   g0975(.A1(new_n1309_), .A2(new_n268_), .ZN(new_n1310_));
  NAND3_X1   g0976(.A1(new_n276_), .A2(\a[8] ), .A3(\a[10] ), .ZN(new_n1311_));
  AOI21_X1   g0977(.A1(new_n1308_), .A2(new_n1310_), .B(new_n1311_), .ZN(new_n1312_));
  NAND3_X1   g0978(.A1(\a[13] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1313_));
  NAND3_X1   g0979(.A1(new_n950_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1314_));
  NAND2_X1   g0980(.A1(new_n1314_), .A2(new_n1313_), .ZN(new_n1315_));
  NAND3_X1   g0981(.A1(\a[11] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1316_));
  NOR2_X1    g0982(.A1(new_n269_), .A2(\a[11] ), .ZN(new_n1317_));
  NAND2_X1   g0983(.A1(new_n1317_), .A2(new_n268_), .ZN(new_n1318_));
  NAND3_X1   g0984(.A1(new_n276_), .A2(\a[12] ), .A3(\a[14] ), .ZN(new_n1319_));
  AOI21_X1   g0985(.A1(new_n1316_), .A2(new_n1318_), .B(new_n1319_), .ZN(new_n1320_));
  NAND4_X1   g0986(.A1(new_n1312_), .A2(new_n1320_), .A3(new_n1307_), .A4(new_n1315_), .ZN(new_n1321_));
  NAND3_X1   g0987(.A1(\a[17] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1322_));
  NAND3_X1   g0988(.A1(new_n631_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1323_));
  NAND2_X1   g0989(.A1(new_n1323_), .A2(new_n1322_), .ZN(new_n1324_));
  NAND3_X1   g0990(.A1(\a[15] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1325_));
  NOR2_X1    g0991(.A1(new_n269_), .A2(\a[15] ), .ZN(new_n1326_));
  NAND2_X1   g0992(.A1(new_n1326_), .A2(new_n268_), .ZN(new_n1327_));
  NAND3_X1   g0993(.A1(new_n276_), .A2(\a[16] ), .A3(\a[18] ), .ZN(new_n1328_));
  AOI21_X1   g0994(.A1(new_n1325_), .A2(new_n1327_), .B(new_n1328_), .ZN(new_n1329_));
  NAND3_X1   g0995(.A1(\a[5] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1330_));
  NAND3_X1   g0996(.A1(new_n972_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1331_));
  NAND2_X1   g0997(.A1(new_n1331_), .A2(new_n1330_), .ZN(new_n1332_));
  AND3_X2    g0998(.A1(\a[3] ), .A2(\shift[0] ), .A3(\shift[1] ), .Z(new_n1333_));
  NOR3_X1    g0999(.A1(new_n269_), .A2(\a[3] ), .A3(\shift[0] ), .ZN(new_n1334_));
  NOR2_X1    g1000(.A1(new_n1333_), .A2(new_n1334_), .ZN(new_n1335_));
  NOR2_X1    g1001(.A1(new_n590_), .A2(new_n554_), .ZN(new_n1336_));
  NAND2_X1   g1002(.A1(new_n1336_), .A2(new_n276_), .ZN(new_n1337_));
  NOR2_X1    g1003(.A1(new_n1335_), .A2(new_n1337_), .ZN(new_n1338_));
  NAND4_X1   g1004(.A1(new_n1329_), .A2(new_n1324_), .A3(new_n1338_), .A4(new_n1332_), .ZN(new_n1339_));
  NOR2_X1    g1005(.A1(new_n1321_), .A2(new_n1339_), .ZN(new_n1340_));
  NOR3_X1    g1006(.A1(new_n1304_), .A2(new_n1340_), .A3(new_n1265_), .ZN(new_n1341_));
  NOR4_X1    g1007(.A1(new_n1284_), .A2(new_n1303_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1342_));
  NOR2_X1    g1008(.A1(new_n1341_), .A2(new_n1342_), .ZN(new_n1343_));
  NAND3_X1   g1009(.A1(\a[41] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1344_));
  NAND3_X1   g1010(.A1(new_n1019_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1345_));
  NAND2_X1   g1011(.A1(new_n1345_), .A2(new_n1344_), .ZN(new_n1346_));
  NAND3_X1   g1012(.A1(\a[39] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1347_));
  NOR2_X1    g1013(.A1(new_n269_), .A2(\a[39] ), .ZN(new_n1348_));
  NAND2_X1   g1014(.A1(new_n1348_), .A2(new_n268_), .ZN(new_n1349_));
  NAND3_X1   g1015(.A1(new_n276_), .A2(\a[40] ), .A3(\a[42] ), .ZN(new_n1350_));
  AOI21_X1   g1016(.A1(new_n1347_), .A2(new_n1349_), .B(new_n1350_), .ZN(new_n1351_));
  NAND3_X1   g1017(.A1(\a[43] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1352_));
  NOR2_X1    g1018(.A1(new_n269_), .A2(\a[43] ), .ZN(new_n1353_));
  NAND2_X1   g1019(.A1(new_n1353_), .A2(new_n268_), .ZN(new_n1354_));
  NAND2_X1   g1020(.A1(new_n1354_), .A2(new_n1352_), .ZN(new_n1355_));
  NAND3_X1   g1021(.A1(\a[45] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1356_));
  NAND3_X1   g1022(.A1(new_n1029_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1357_));
  NAND3_X1   g1023(.A1(new_n276_), .A2(\a[44] ), .A3(\a[46] ), .ZN(new_n1358_));
  AOI21_X1   g1024(.A1(new_n1356_), .A2(new_n1357_), .B(new_n1358_), .ZN(new_n1359_));
  NAND4_X1   g1025(.A1(new_n1351_), .A2(new_n1359_), .A3(new_n1346_), .A4(new_n1355_), .ZN(new_n1360_));
  NAND3_X1   g1026(.A1(\a[49] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1361_));
  NAND3_X1   g1027(.A1(new_n999_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1362_));
  NAND2_X1   g1028(.A1(new_n1362_), .A2(new_n1361_), .ZN(new_n1363_));
  NAND3_X1   g1029(.A1(\a[47] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1364_));
  INV_X1     g1030(.I(new_n1364_), .ZN(new_n1365_));
  NOR3_X1    g1031(.A1(new_n269_), .A2(\a[47] ), .A3(\shift[0] ), .ZN(new_n1366_));
  NOR2_X1    g1032(.A1(new_n1365_), .A2(new_n1366_), .ZN(new_n1367_));
  NOR2_X1    g1033(.A1(new_n690_), .A2(new_n517_), .ZN(new_n1368_));
  NAND2_X1   g1034(.A1(new_n1368_), .A2(new_n276_), .ZN(new_n1369_));
  NOR2_X1    g1035(.A1(new_n1367_), .A2(new_n1369_), .ZN(new_n1370_));
  NAND3_X1   g1036(.A1(\a[37] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1371_));
  NAND3_X1   g1037(.A1(new_n642_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1372_));
  NAND2_X1   g1038(.A1(new_n1372_), .A2(new_n1371_), .ZN(new_n1373_));
  NOR3_X1    g1039(.A1(new_n992_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n1374_));
  NOR3_X1    g1040(.A1(new_n269_), .A2(\a[35] ), .A3(\shift[0] ), .ZN(new_n1375_));
  NOR2_X1    g1041(.A1(new_n1374_), .A2(new_n1375_), .ZN(new_n1376_));
  NAND3_X1   g1042(.A1(new_n276_), .A2(\a[36] ), .A3(\a[38] ), .ZN(new_n1377_));
  NOR2_X1    g1043(.A1(new_n1376_), .A2(new_n1377_), .ZN(new_n1378_));
  NAND4_X1   g1044(.A1(new_n1378_), .A2(new_n1370_), .A3(new_n1363_), .A4(new_n1373_), .ZN(new_n1379_));
  NOR3_X1    g1045(.A1(new_n1360_), .A2(new_n1379_), .A3(new_n893_), .ZN(new_n1380_));
  NAND3_X1   g1046(.A1(\a[25] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1381_));
  NAND3_X1   g1047(.A1(new_n1033_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1382_));
  NAND2_X1   g1048(.A1(new_n1382_), .A2(new_n1381_), .ZN(new_n1383_));
  NOR3_X1    g1049(.A1(new_n602_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n1384_));
  NOR3_X1    g1050(.A1(new_n269_), .A2(\a[23] ), .A3(\shift[0] ), .ZN(new_n1385_));
  NOR2_X1    g1051(.A1(new_n1384_), .A2(new_n1385_), .ZN(new_n1386_));
  NAND3_X1   g1052(.A1(new_n276_), .A2(\a[24] ), .A3(\a[26] ), .ZN(new_n1387_));
  NOR2_X1    g1053(.A1(new_n1386_), .A2(new_n1387_), .ZN(new_n1388_));
  NAND3_X1   g1054(.A1(\a[29] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1389_));
  NAND3_X1   g1055(.A1(new_n1045_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1390_));
  NAND2_X1   g1056(.A1(new_n1390_), .A2(new_n1389_), .ZN(new_n1391_));
  NOR3_X1    g1057(.A1(new_n1052_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n1392_));
  NOR3_X1    g1058(.A1(new_n269_), .A2(\a[27] ), .A3(\shift[0] ), .ZN(new_n1393_));
  NOR2_X1    g1059(.A1(new_n1392_), .A2(new_n1393_), .ZN(new_n1394_));
  NAND3_X1   g1060(.A1(new_n276_), .A2(\a[28] ), .A3(\a[30] ), .ZN(new_n1395_));
  NOR2_X1    g1061(.A1(new_n1394_), .A2(new_n1395_), .ZN(new_n1396_));
  NAND4_X1   g1062(.A1(new_n1388_), .A2(new_n1396_), .A3(new_n1383_), .A4(new_n1391_), .ZN(new_n1397_));
  NAND3_X1   g1063(.A1(\a[33] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1398_));
  NAND3_X1   g1064(.A1(new_n1059_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1399_));
  NAND2_X1   g1065(.A1(new_n1399_), .A2(new_n1398_), .ZN(new_n1400_));
  AND3_X2    g1066(.A1(\a[31] ), .A2(\shift[0] ), .A3(\shift[1] ), .Z(new_n1401_));
  NOR3_X1    g1067(.A1(new_n269_), .A2(\a[31] ), .A3(\shift[0] ), .ZN(new_n1402_));
  NOR2_X1    g1068(.A1(new_n1401_), .A2(new_n1402_), .ZN(new_n1403_));
  NAND3_X1   g1069(.A1(new_n276_), .A2(\a[32] ), .A3(\a[34] ), .ZN(new_n1404_));
  NOR2_X1    g1070(.A1(new_n1403_), .A2(new_n1404_), .ZN(new_n1405_));
  NAND3_X1   g1071(.A1(\a[21] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1406_));
  NAND3_X1   g1072(.A1(new_n1072_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1407_));
  NAND2_X1   g1073(.A1(new_n1407_), .A2(new_n1406_), .ZN(new_n1408_));
  NOR3_X1    g1074(.A1(new_n635_), .A2(new_n294_), .A3(new_n269_), .ZN(new_n1409_));
  NOR3_X1    g1075(.A1(new_n269_), .A2(\a[19] ), .A3(\shift[0] ), .ZN(new_n1410_));
  NOR2_X1    g1076(.A1(new_n1409_), .A2(new_n1410_), .ZN(new_n1411_));
  NAND3_X1   g1077(.A1(new_n276_), .A2(\a[20] ), .A3(\a[22] ), .ZN(new_n1412_));
  NOR2_X1    g1078(.A1(new_n1411_), .A2(new_n1412_), .ZN(new_n1413_));
  NAND4_X1   g1079(.A1(new_n1413_), .A2(new_n1405_), .A3(new_n1400_), .A4(new_n1408_), .ZN(new_n1414_));
  NOR2_X1    g1080(.A1(new_n1397_), .A2(new_n1414_), .ZN(new_n1415_));
  NOR3_X1    g1081(.A1(new_n1380_), .A2(new_n1415_), .A3(new_n1265_), .ZN(new_n1416_));
  NOR4_X1    g1082(.A1(new_n1360_), .A2(new_n1379_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1417_));
  NOR2_X1    g1083(.A1(new_n1416_), .A2(new_n1417_), .ZN(new_n1418_));
  OAI21_X1   g1084(.A1(new_n1343_), .A2(new_n1418_), .B(\shift[6] ), .ZN(new_n1419_));
  NAND2_X1   g1085(.A1(new_n1419_), .A2(new_n1264_), .ZN(\result[2] ));
  NOR2_X1    g1086(.A1(new_n843_), .A2(new_n294_), .ZN(new_n1421_));
  NOR2_X1    g1087(.A1(new_n294_), .A2(\a[106] ), .ZN(new_n1422_));
  MUX2_X1    g1088(.I0(new_n1422_), .I1(new_n1421_), .S(\shift[1] ), .Z(new_n1423_));
  NAND2_X1   g1089(.A1(\a[104] ), .A2(\shift[0] ), .ZN(new_n1424_));
  NAND4_X1   g1090(.A1(new_n1424_), .A2(new_n859_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1425_));
  NAND3_X1   g1091(.A1(\a[104] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1427_));
  AOI21_X1   g1092(.A1(new_n1425_), .A2(new_n1427_), .B(new_n323_), .ZN(new_n1428_));
  NOR2_X1    g1093(.A1(new_n853_), .A2(new_n294_), .ZN(new_n1429_));
  NOR2_X1    g1094(.A1(new_n294_), .A2(\a[110] ), .ZN(new_n1430_));
  MUX2_X1    g1095(.I0(new_n1430_), .I1(new_n1429_), .S(\shift[1] ), .Z(new_n1431_));
  NAND2_X1   g1096(.A1(\a[108] ), .A2(\shift[0] ), .ZN(new_n1432_));
  NAND4_X1   g1097(.A1(new_n1432_), .A2(new_n872_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1433_));
  NAND3_X1   g1098(.A1(\a[108] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1435_));
  AOI21_X1   g1099(.A1(new_n1433_), .A2(new_n1435_), .B(new_n323_), .ZN(new_n1436_));
  NAND4_X1   g1100(.A1(new_n1423_), .A2(new_n1431_), .A3(new_n1428_), .A4(new_n1436_), .ZN(new_n1437_));
  NOR2_X1    g1101(.A1(new_n307_), .A2(new_n294_), .ZN(new_n1438_));
  NOR2_X1    g1102(.A1(new_n294_), .A2(\a[114] ), .ZN(new_n1439_));
  MUX2_X1    g1103(.I0(new_n1439_), .I1(new_n1438_), .S(\shift[1] ), .Z(new_n1440_));
  NAND2_X1   g1104(.A1(\a[112] ), .A2(\shift[0] ), .ZN(new_n1441_));
  NAND4_X1   g1105(.A1(new_n1441_), .A2(new_n330_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1442_));
  NAND3_X1   g1106(.A1(\a[112] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1444_));
  AOI21_X1   g1107(.A1(new_n1442_), .A2(new_n1444_), .B(new_n323_), .ZN(new_n1445_));
  NOR2_X1    g1108(.A1(new_n878_), .A2(new_n294_), .ZN(new_n1446_));
  NOR2_X1    g1109(.A1(new_n294_), .A2(\a[102] ), .ZN(new_n1447_));
  MUX2_X1    g1110(.I0(new_n1447_), .I1(new_n1446_), .S(\shift[1] ), .Z(new_n1448_));
  NAND2_X1   g1111(.A1(\a[100] ), .A2(\shift[0] ), .ZN(new_n1449_));
  NAND4_X1   g1112(.A1(new_n1449_), .A2(new_n435_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1450_));
  NAND3_X1   g1113(.A1(\a[100] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1451_));
  AOI21_X1   g1114(.A1(new_n1450_), .A2(new_n1451_), .B(new_n323_), .ZN(new_n1452_));
  NAND4_X1   g1115(.A1(new_n1440_), .A2(new_n1448_), .A3(new_n1445_), .A4(new_n1452_), .ZN(new_n1453_));
  NOR3_X1    g1116(.A1(new_n1437_), .A2(new_n1453_), .A3(new_n893_), .ZN(new_n1454_));
  NOR2_X1    g1117(.A1(new_n395_), .A2(new_n294_), .ZN(new_n1455_));
  NOR2_X1    g1118(.A1(new_n294_), .A2(\a[90] ), .ZN(new_n1456_));
  MUX2_X1    g1119(.I0(new_n1456_), .I1(new_n1455_), .S(\shift[1] ), .Z(new_n1457_));
  NAND2_X1   g1120(.A1(\a[88] ), .A2(\shift[0] ), .ZN(new_n1458_));
  NAND4_X1   g1121(.A1(new_n1458_), .A2(new_n399_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1459_));
  NAND3_X1   g1122(.A1(\a[88] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1460_));
  AOI21_X1   g1123(.A1(new_n1459_), .A2(new_n1460_), .B(new_n323_), .ZN(new_n1461_));
  NOR2_X1    g1124(.A1(new_n810_), .A2(new_n294_), .ZN(new_n1462_));
  NOR2_X1    g1125(.A1(new_n294_), .A2(\a[94] ), .ZN(new_n1463_));
  MUX2_X1    g1126(.I0(new_n1463_), .I1(new_n1462_), .S(\shift[1] ), .Z(new_n1464_));
  NAND2_X1   g1127(.A1(\a[92] ), .A2(\shift[0] ), .ZN(new_n1465_));
  NAND4_X1   g1128(.A1(new_n1465_), .A2(new_n411_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1466_));
  NAND3_X1   g1129(.A1(\a[92] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1467_));
  AOI21_X1   g1130(.A1(new_n1466_), .A2(new_n1467_), .B(new_n323_), .ZN(new_n1468_));
  NAND4_X1   g1131(.A1(new_n1457_), .A2(new_n1464_), .A3(new_n1461_), .A4(new_n1468_), .ZN(new_n1469_));
  NAND3_X1   g1132(.A1(new_n470_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1471_));
  NAND3_X1   g1133(.A1(\a[97] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1473_));
  NAND2_X1   g1134(.A1(new_n1471_), .A2(new_n1473_), .ZN(new_n1474_));
  NAND2_X1   g1135(.A1(\a[96] ), .A2(\shift[0] ), .ZN(new_n1475_));
  NAND4_X1   g1136(.A1(new_n1475_), .A2(new_n883_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1476_));
  NAND3_X1   g1137(.A1(\a[96] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1477_));
  AOI21_X1   g1138(.A1(new_n1476_), .A2(new_n1477_), .B(new_n323_), .ZN(new_n1478_));
  NAND3_X1   g1139(.A1(new_n1220_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1480_));
  NAND3_X1   g1140(.A1(\a[85] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1482_));
  NAND2_X1   g1141(.A1(new_n1480_), .A2(new_n1482_), .ZN(new_n1483_));
  NAND2_X1   g1142(.A1(\a[84] ), .A2(\shift[0] ), .ZN(new_n1484_));
  NAND4_X1   g1143(.A1(new_n1484_), .A2(new_n390_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1485_));
  NAND3_X1   g1144(.A1(\a[84] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1486_));
  AOI21_X1   g1145(.A1(new_n1485_), .A2(new_n1486_), .B(new_n323_), .ZN(new_n1487_));
  NAND4_X1   g1146(.A1(new_n1478_), .A2(new_n1487_), .A3(new_n1474_), .A4(new_n1483_), .ZN(new_n1488_));
  OAI21_X1   g1147(.A1(new_n1469_), .A2(new_n1488_), .B(\shift[5] ), .ZN(new_n1489_));
  NOR3_X1    g1148(.A1(new_n1454_), .A2(new_n1489_), .A3(\shift[4] ), .ZN(new_n1490_));
  NOR4_X1    g1149(.A1(new_n1437_), .A2(new_n1453_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1492_));
  NOR2_X1    g1150(.A1(new_n1490_), .A2(new_n1492_), .ZN(new_n1493_));
  NOR2_X1    g1151(.A1(new_n699_), .A2(new_n294_), .ZN(new_n1494_));
  NOR2_X1    g1152(.A1(new_n294_), .A2(\a[122] ), .ZN(new_n1495_));
  MUX2_X1    g1153(.I0(new_n1495_), .I1(new_n1494_), .S(\shift[1] ), .Z(new_n1496_));
  NAND2_X1   g1154(.A1(\a[120] ), .A2(\shift[0] ), .ZN(new_n1497_));
  NAND4_X1   g1155(.A1(new_n1497_), .A2(new_n287_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1498_));
  NAND3_X1   g1156(.A1(\a[120] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1500_));
  AOI21_X1   g1157(.A1(new_n1498_), .A2(new_n1500_), .B(new_n323_), .ZN(new_n1501_));
  NOR2_X1    g1158(.A1(new_n293_), .A2(new_n294_), .ZN(new_n1502_));
  NOR2_X1    g1159(.A1(new_n294_), .A2(\a[126] ), .ZN(new_n1503_));
  MUX2_X1    g1160(.I0(new_n1503_), .I1(new_n1502_), .S(\shift[1] ), .Z(new_n1504_));
  NAND3_X1   g1161(.A1(\a[124] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1505_));
  NAND2_X1   g1162(.A1(new_n727_), .A2(new_n1505_), .ZN(new_n1506_));
  NAND4_X1   g1163(.A1(new_n730_), .A2(\a[124] ), .A3(\shift[0] ), .A4(\shift[1] ), .ZN(new_n1507_));
  AOI21_X1   g1164(.A1(new_n1507_), .A2(new_n1506_), .B(new_n323_), .ZN(new_n1508_));
  NAND4_X1   g1165(.A1(new_n1508_), .A2(new_n1496_), .A3(new_n1501_), .A4(new_n1504_), .ZN(new_n1509_));
  NOR2_X1    g1166(.A1(new_n294_), .A2(\a[2] ), .ZN(new_n1510_));
  NAND3_X1   g1167(.A1(new_n1510_), .A2(new_n269_), .A3(new_n720_), .ZN(new_n1511_));
  NAND3_X1   g1168(.A1(\a[1] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1512_));
  NAND2_X1   g1169(.A1(new_n1511_), .A2(new_n1512_), .ZN(new_n1513_));
  NOR2_X1    g1170(.A1(new_n269_), .A2(\a[3] ), .ZN(new_n1514_));
  NAND3_X1   g1171(.A1(new_n1514_), .A2(new_n294_), .A3(new_n726_), .ZN(new_n1515_));
  NAND3_X1   g1172(.A1(\a[0] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1516_));
  AOI21_X1   g1173(.A1(new_n1515_), .A2(new_n1516_), .B(new_n323_), .ZN(new_n1517_));
  NOR2_X1    g1174(.A1(new_n733_), .A2(new_n294_), .ZN(new_n1518_));
  NOR2_X1    g1175(.A1(new_n294_), .A2(\a[118] ), .ZN(new_n1519_));
  MUX2_X1    g1176(.I0(new_n1519_), .I1(new_n1518_), .S(\shift[1] ), .Z(new_n1520_));
  NAND2_X1   g1177(.A1(\a[116] ), .A2(\shift[0] ), .ZN(new_n1521_));
  NAND4_X1   g1178(.A1(new_n1521_), .A2(new_n274_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1522_));
  NAND3_X1   g1179(.A1(\a[116] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1523_));
  AOI21_X1   g1180(.A1(new_n1522_), .A2(new_n1523_), .B(new_n323_), .ZN(new_n1524_));
  NAND4_X1   g1181(.A1(new_n1517_), .A2(new_n1520_), .A3(new_n1513_), .A4(new_n1524_), .ZN(new_n1525_));
  NOR3_X1    g1182(.A1(new_n1509_), .A2(new_n893_), .A3(new_n1525_), .ZN(new_n1526_));
  NOR2_X1    g1183(.A1(new_n749_), .A2(new_n294_), .ZN(new_n1527_));
  NOR2_X1    g1184(.A1(new_n294_), .A2(\a[74] ), .ZN(new_n1528_));
  MUX2_X1    g1185(.I0(new_n1528_), .I1(new_n1527_), .S(\shift[1] ), .Z(new_n1529_));
  NAND2_X1   g1186(.A1(\a[72] ), .A2(\shift[0] ), .ZN(new_n1530_));
  NAND4_X1   g1187(.A1(new_n1530_), .A2(new_n765_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1531_));
  NAND3_X1   g1188(.A1(\a[72] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1532_));
  AOI21_X1   g1189(.A1(new_n1531_), .A2(new_n1532_), .B(new_n323_), .ZN(new_n1533_));
  NOR2_X1    g1190(.A1(new_n760_), .A2(new_n294_), .ZN(new_n1534_));
  NOR2_X1    g1191(.A1(new_n294_), .A2(\a[78] ), .ZN(new_n1535_));
  MUX2_X1    g1192(.I0(new_n1535_), .I1(new_n1534_), .S(\shift[1] ), .Z(new_n1536_));
  NAND2_X1   g1193(.A1(\a[76] ), .A2(\shift[0] ), .ZN(new_n1537_));
  NAND4_X1   g1194(.A1(new_n1537_), .A2(new_n778_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1538_));
  NAND3_X1   g1195(.A1(\a[76] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1540_));
  AOI21_X1   g1196(.A1(new_n1538_), .A2(new_n1540_), .B(new_n323_), .ZN(new_n1541_));
  NAND4_X1   g1197(.A1(new_n1529_), .A2(new_n1536_), .A3(new_n1533_), .A4(new_n1541_), .ZN(new_n1542_));
  NOR2_X1    g1198(.A1(new_n418_), .A2(new_n294_), .ZN(new_n1543_));
  NOR2_X1    g1199(.A1(new_n294_), .A2(\a[82] ), .ZN(new_n1544_));
  MUX2_X1    g1200(.I0(new_n1544_), .I1(new_n1543_), .S(\shift[1] ), .Z(new_n1545_));
  NAND2_X1   g1201(.A1(\a[80] ), .A2(\shift[0] ), .ZN(new_n1546_));
  NAND4_X1   g1202(.A1(new_n1546_), .A2(new_n422_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1547_));
  NAND3_X1   g1203(.A1(\a[80] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1549_));
  AOI21_X1   g1204(.A1(new_n1547_), .A2(new_n1549_), .B(new_n323_), .ZN(new_n1550_));
  NAND3_X1   g1205(.A1(new_n1178_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1552_));
  NAND3_X1   g1206(.A1(\a[69] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1554_));
  NAND2_X1   g1207(.A1(new_n1552_), .A2(new_n1554_), .ZN(new_n1555_));
  NAND2_X1   g1208(.A1(\a[68] ), .A2(\shift[0] ), .ZN(new_n1556_));
  NAND4_X1   g1209(.A1(new_n1556_), .A2(new_n342_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1557_));
  NAND3_X1   g1210(.A1(\a[68] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1558_));
  AOI21_X1   g1211(.A1(new_n1557_), .A2(new_n1558_), .B(new_n323_), .ZN(new_n1559_));
  NAND4_X1   g1212(.A1(new_n1545_), .A2(new_n1550_), .A3(new_n1559_), .A4(new_n1555_), .ZN(new_n1560_));
  OAI21_X1   g1213(.A1(new_n1542_), .A2(new_n1560_), .B(new_n984_), .ZN(new_n1561_));
  NOR2_X1    g1214(.A1(new_n1526_), .A2(new_n1561_), .ZN(new_n1562_));
  NOR2_X1    g1215(.A1(new_n1542_), .A2(new_n1560_), .ZN(new_n1563_));
  NOR4_X1    g1216(.A1(new_n1509_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1525_), .ZN(new_n1564_));
  NOR2_X1    g1217(.A1(new_n1562_), .A2(new_n1564_), .ZN(new_n1565_));
  OAI21_X1   g1218(.A1(new_n1565_), .A2(new_n1493_), .B(new_n264_), .ZN(new_n1566_));
  NOR2_X1    g1219(.A1(new_n560_), .A2(new_n294_), .ZN(new_n1567_));
  NOR2_X1    g1220(.A1(new_n294_), .A2(\a[10] ), .ZN(new_n1568_));
  MUX2_X1    g1221(.I0(new_n1568_), .I1(new_n1567_), .S(\shift[1] ), .Z(new_n1569_));
  NAND2_X1   g1222(.A1(\a[8] ), .A2(\shift[0] ), .ZN(new_n1570_));
  NAND4_X1   g1223(.A1(new_n1570_), .A2(new_n564_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1571_));
  NAND3_X1   g1224(.A1(\a[8] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1572_));
  AOI21_X1   g1225(.A1(new_n1571_), .A2(new_n1572_), .B(new_n323_), .ZN(new_n1573_));
  NOR2_X1    g1226(.A1(new_n950_), .A2(new_n294_), .ZN(new_n1574_));
  NOR2_X1    g1227(.A1(new_n294_), .A2(\a[14] ), .ZN(new_n1575_));
  MUX2_X1    g1228(.I0(new_n1575_), .I1(new_n1574_), .S(\shift[1] ), .Z(new_n1576_));
  NAND2_X1   g1229(.A1(\a[12] ), .A2(\shift[0] ), .ZN(new_n1577_));
  NAND4_X1   g1230(.A1(new_n1577_), .A2(new_n576_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1578_));
  NAND3_X1   g1231(.A1(\a[12] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1579_));
  AOI21_X1   g1232(.A1(new_n1578_), .A2(new_n1579_), .B(new_n323_), .ZN(new_n1580_));
  NAND4_X1   g1233(.A1(new_n1569_), .A2(new_n1576_), .A3(new_n1573_), .A4(new_n1580_), .ZN(new_n1581_));
  NOR2_X1    g1234(.A1(new_n631_), .A2(new_n294_), .ZN(new_n1582_));
  NOR2_X1    g1235(.A1(new_n294_), .A2(\a[18] ), .ZN(new_n1583_));
  MUX2_X1    g1236(.I0(new_n1583_), .I1(new_n1582_), .S(\shift[1] ), .Z(new_n1584_));
  NAND2_X1   g1237(.A1(\a[16] ), .A2(\shift[0] ), .ZN(new_n1585_));
  NAND4_X1   g1238(.A1(new_n1585_), .A2(new_n635_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1586_));
  NAND3_X1   g1239(.A1(\a[16] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1588_));
  AOI21_X1   g1240(.A1(new_n1586_), .A2(new_n1588_), .B(new_n323_), .ZN(new_n1589_));
  NAND3_X1   g1241(.A1(new_n554_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1591_));
  NAND3_X1   g1242(.A1(\a[5] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1593_));
  NAND2_X1   g1243(.A1(new_n1591_), .A2(new_n1593_), .ZN(new_n1594_));
  NAND2_X1   g1244(.A1(\a[4] ), .A2(\shift[0] ), .ZN(new_n1595_));
  NAND4_X1   g1245(.A1(new_n1595_), .A2(new_n944_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1596_));
  NAND3_X1   g1246(.A1(\a[4] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1597_));
  AOI21_X1   g1247(.A1(new_n1596_), .A2(new_n1597_), .B(new_n323_), .ZN(new_n1598_));
  NAND4_X1   g1248(.A1(new_n1584_), .A2(new_n1589_), .A3(new_n1598_), .A4(new_n1594_), .ZN(new_n1599_));
  OAI21_X1   g1249(.A1(new_n1581_), .A2(new_n1599_), .B(\shift[5] ), .ZN(new_n1600_));
  XOR2_X1    g1250(.A1(new_n1600_), .A2(new_n987_), .Z(new_n1601_));
  NOR2_X1    g1251(.A1(new_n894_), .A2(new_n294_), .ZN(new_n1602_));
  NOR2_X1    g1252(.A1(new_n294_), .A2(\a[58] ), .ZN(new_n1603_));
  MUX2_X1    g1253(.I0(new_n1603_), .I1(new_n1602_), .S(\shift[1] ), .Z(new_n1604_));
  NAND2_X1   g1254(.A1(\a[56] ), .A2(\shift[0] ), .ZN(new_n1605_));
  NAND4_X1   g1255(.A1(new_n1605_), .A2(new_n494_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1606_));
  NAND3_X1   g1256(.A1(\a[56] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1607_));
  AOI21_X1   g1257(.A1(new_n1606_), .A2(new_n1607_), .B(new_n323_), .ZN(new_n1608_));
  NOR2_X1    g1258(.A1(new_n905_), .A2(new_n294_), .ZN(new_n1609_));
  NOR2_X1    g1259(.A1(new_n294_), .A2(\a[62] ), .ZN(new_n1610_));
  MUX2_X1    g1260(.I0(new_n1610_), .I1(new_n1609_), .S(\shift[1] ), .Z(new_n1611_));
  NAND2_X1   g1261(.A1(\a[60] ), .A2(\shift[0] ), .ZN(new_n1612_));
  NAND4_X1   g1262(.A1(new_n1612_), .A2(new_n530_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1613_));
  NAND3_X1   g1263(.A1(\a[60] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1615_));
  AOI21_X1   g1264(.A1(new_n1613_), .A2(new_n1615_), .B(new_n323_), .ZN(new_n1616_));
  NAND4_X1   g1265(.A1(new_n1604_), .A2(new_n1611_), .A3(new_n1608_), .A4(new_n1616_), .ZN(new_n1617_));
  NOR2_X1    g1266(.A1(new_n917_), .A2(new_n294_), .ZN(new_n1618_));
  NOR2_X1    g1267(.A1(new_n294_), .A2(\a[66] ), .ZN(new_n1619_));
  MUX2_X1    g1268(.I0(new_n1619_), .I1(new_n1618_), .S(\shift[1] ), .Z(new_n1620_));
  NAND2_X1   g1269(.A1(\a[64] ), .A2(\shift[0] ), .ZN(new_n1621_));
  NAND4_X1   g1270(.A1(new_n1621_), .A2(new_n377_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1622_));
  NAND3_X1   g1271(.A1(\a[64] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1624_));
  AOI21_X1   g1272(.A1(new_n1622_), .A2(new_n1624_), .B(new_n323_), .ZN(new_n1625_));
  NOR2_X1    g1273(.A1(new_n927_), .A2(new_n294_), .ZN(new_n1626_));
  NOR2_X1    g1274(.A1(new_n294_), .A2(\a[54] ), .ZN(new_n1627_));
  MUX2_X1    g1275(.I0(new_n1627_), .I1(new_n1626_), .S(\shift[1] ), .Z(new_n1628_));
  NAND2_X1   g1276(.A1(\a[52] ), .A2(\shift[0] ), .ZN(new_n1629_));
  NAND4_X1   g1277(.A1(new_n1629_), .A2(new_n483_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1630_));
  NAND3_X1   g1278(.A1(\a[52] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1631_));
  AOI21_X1   g1279(.A1(new_n1630_), .A2(new_n1631_), .B(new_n323_), .ZN(new_n1632_));
  NAND4_X1   g1280(.A1(new_n1620_), .A2(new_n1628_), .A3(new_n1625_), .A4(new_n1632_), .ZN(new_n1633_));
  NOR4_X1    g1281(.A1(new_n1617_), .A2(new_n1633_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1634_));
  OAI21_X1   g1282(.A1(new_n1617_), .A2(new_n1633_), .B(\shift[4] ), .ZN(new_n1635_));
  NOR2_X1    g1283(.A1(new_n1635_), .A2(new_n987_), .ZN(new_n1636_));
  NAND3_X1   g1284(.A1(new_n676_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1638_));
  NAND3_X1   g1285(.A1(\a[41] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1640_));
  NAND2_X1   g1286(.A1(new_n1638_), .A2(new_n1640_), .ZN(new_n1641_));
  NAND2_X1   g1287(.A1(\a[40] ), .A2(\shift[0] ), .ZN(new_n1642_));
  NAND4_X1   g1288(.A1(new_n1642_), .A2(new_n1028_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1643_));
  NAND3_X1   g1289(.A1(\a[40] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1644_));
  AOI21_X1   g1290(.A1(new_n1643_), .A2(new_n1644_), .B(new_n323_), .ZN(new_n1645_));
  NAND3_X1   g1291(.A1(\a[44] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1646_));
  NAND3_X1   g1292(.A1(new_n677_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n1647_));
  NAND2_X1   g1293(.A1(new_n1647_), .A2(new_n1646_), .ZN(new_n1648_));
  NAND3_X1   g1294(.A1(\a[46] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1649_));
  NAND3_X1   g1295(.A1(new_n689_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1650_));
  NAND2_X1   g1296(.A1(new_n1650_), .A2(new_n1649_), .ZN(new_n1651_));
  NOR3_X1    g1297(.A1(new_n323_), .A2(new_n1029_), .A3(new_n1005_), .ZN(new_n1652_));
  AND2_X2    g1298(.A1(new_n1651_), .A2(new_n1652_), .Z(new_n1653_));
  NAND4_X1   g1299(.A1(new_n1653_), .A2(new_n1641_), .A3(new_n1645_), .A4(new_n1648_), .ZN(new_n1654_));
  NAND3_X1   g1300(.A1(new_n517_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1656_));
  NAND3_X1   g1301(.A1(\a[49] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1658_));
  NAND2_X1   g1302(.A1(new_n1656_), .A2(new_n1658_), .ZN(new_n1659_));
  NAND2_X1   g1303(.A1(\a[48] ), .A2(\shift[0] ), .ZN(new_n1660_));
  NAND4_X1   g1304(.A1(new_n1660_), .A2(new_n539_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1661_));
  NAND3_X1   g1305(.A1(\a[48] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1663_));
  AOI21_X1   g1306(.A1(new_n1661_), .A2(new_n1663_), .B(new_n323_), .ZN(new_n1664_));
  NAND3_X1   g1307(.A1(new_n648_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1665_));
  NAND3_X1   g1308(.A1(\a[37] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1667_));
  NAND2_X1   g1309(.A1(new_n1665_), .A2(new_n1667_), .ZN(new_n1668_));
  NAND2_X1   g1310(.A1(\a[36] ), .A2(\shift[0] ), .ZN(new_n1669_));
  NAND4_X1   g1311(.A1(new_n1669_), .A2(new_n647_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1670_));
  NAND3_X1   g1312(.A1(\a[36] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1671_));
  AOI21_X1   g1313(.A1(new_n1670_), .A2(new_n1671_), .B(new_n323_), .ZN(new_n1672_));
  NAND4_X1   g1314(.A1(new_n1664_), .A2(new_n1672_), .A3(new_n1659_), .A4(new_n1668_), .ZN(new_n1673_));
  NOR2_X1    g1315(.A1(new_n1033_), .A2(new_n294_), .ZN(new_n1674_));
  NOR2_X1    g1316(.A1(new_n294_), .A2(\a[26] ), .ZN(new_n1675_));
  MUX2_X1    g1317(.I0(new_n1675_), .I1(new_n1674_), .S(\shift[1] ), .Z(new_n1676_));
  NAND2_X1   g1318(.A1(\a[24] ), .A2(\shift[0] ), .ZN(new_n1677_));
  NAND4_X1   g1319(.A1(new_n1677_), .A2(new_n1052_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1678_));
  NAND3_X1   g1320(.A1(\a[24] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1680_));
  AOI21_X1   g1321(.A1(new_n1678_), .A2(new_n1680_), .B(new_n323_), .ZN(new_n1681_));
  NOR2_X1    g1322(.A1(new_n1045_), .A2(new_n294_), .ZN(new_n1682_));
  NOR2_X1    g1323(.A1(new_n294_), .A2(\a[30] ), .ZN(new_n1683_));
  MUX2_X1    g1324(.I0(new_n1683_), .I1(new_n1682_), .S(\shift[1] ), .Z(new_n1684_));
  NAND2_X1   g1325(.A1(\a[28] ), .A2(\shift[0] ), .ZN(new_n1685_));
  NAND4_X1   g1326(.A1(new_n1685_), .A2(new_n1066_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1686_));
  NAND3_X1   g1327(.A1(\a[28] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1688_));
  AOI21_X1   g1328(.A1(new_n1686_), .A2(new_n1688_), .B(new_n323_), .ZN(new_n1689_));
  NAND4_X1   g1329(.A1(new_n1676_), .A2(new_n1684_), .A3(new_n1681_), .A4(new_n1689_), .ZN(new_n1690_));
  NAND3_X1   g1330(.A1(new_n663_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1692_));
  NAND3_X1   g1331(.A1(\a[33] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1694_));
  NAND2_X1   g1332(.A1(new_n1692_), .A2(new_n1694_), .ZN(new_n1695_));
  NAND2_X1   g1333(.A1(\a[32] ), .A2(\shift[0] ), .ZN(new_n1696_));
  NAND4_X1   g1334(.A1(new_n1696_), .A2(new_n992_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1697_));
  NAND3_X1   g1335(.A1(\a[32] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1699_));
  AOI21_X1   g1336(.A1(new_n1697_), .A2(new_n1699_), .B(new_n323_), .ZN(new_n1700_));
  NOR2_X1    g1337(.A1(new_n1072_), .A2(new_n294_), .ZN(new_n1701_));
  NOR2_X1    g1338(.A1(new_n294_), .A2(\a[22] ), .ZN(new_n1702_));
  MUX2_X1    g1339(.I0(new_n1702_), .I1(new_n1701_), .S(\shift[1] ), .Z(new_n1703_));
  NAND2_X1   g1340(.A1(\a[20] ), .A2(\shift[0] ), .ZN(new_n1704_));
  NAND4_X1   g1341(.A1(new_n1704_), .A2(new_n602_), .A3(new_n294_), .A4(\shift[1] ), .ZN(new_n1705_));
  NAND3_X1   g1342(.A1(\a[20] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1707_));
  AOI21_X1   g1343(.A1(new_n1705_), .A2(new_n1707_), .B(new_n323_), .ZN(new_n1708_));
  NAND4_X1   g1344(.A1(new_n1703_), .A2(new_n1700_), .A3(new_n1708_), .A4(new_n1695_), .ZN(new_n1709_));
  NOR4_X1    g1345(.A1(new_n1654_), .A2(new_n1673_), .A3(new_n1690_), .A4(new_n1709_), .ZN(new_n1710_));
  OAI21_X1   g1346(.A1(new_n1636_), .A2(new_n1634_), .B(new_n1710_), .ZN(new_n1711_));
  OAI21_X1   g1347(.A1(new_n1601_), .A2(new_n1711_), .B(\shift[6] ), .ZN(new_n1712_));
  NAND2_X1   g1348(.A1(new_n1712_), .A2(new_n1566_), .ZN(\result[3] ));
  NAND4_X1   g1349(.A1(new_n305_), .A2(new_n593_), .A3(new_n296_), .A4(new_n585_), .ZN(new_n1714_));
  NOR4_X1    g1350(.A1(new_n291_), .A2(new_n1714_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1715_));
  NAND3_X1   g1351(.A1(\a[3] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1716_));
  NAND3_X1   g1352(.A1(new_n977_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1717_));
  NAND2_X1   g1353(.A1(new_n1717_), .A2(new_n1716_), .ZN(new_n1718_));
  NAND4_X1   g1354(.A1(new_n585_), .A2(new_n1718_), .A3(new_n276_), .A4(new_n591_), .ZN(new_n1719_));
  NOR4_X1    g1355(.A1(new_n319_), .A2(new_n325_), .A3(new_n329_), .A4(new_n1719_), .ZN(new_n1720_));
  NOR3_X1    g1356(.A1(new_n1720_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1721_));
  NOR2_X1    g1357(.A1(new_n1721_), .A2(new_n1715_), .ZN(new_n1722_));
  NAND4_X1   g1358(.A1(new_n428_), .A2(new_n347_), .A3(new_n341_), .A4(new_n420_), .ZN(new_n1723_));
  NAND4_X1   g1359(.A1(new_n360_), .A2(new_n371_), .A3(new_n351_), .A4(new_n365_), .ZN(new_n1724_));
  NOR4_X1    g1360(.A1(new_n1723_), .A2(new_n1724_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1725_));
  NOR2_X1    g1361(.A1(new_n1723_), .A2(new_n1724_), .ZN(new_n1726_));
  NOR3_X1    g1362(.A1(new_n1726_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n1727_));
  NAND4_X1   g1363(.A1(new_n416_), .A2(new_n474_), .A3(new_n410_), .A4(new_n465_), .ZN(new_n1728_));
  NAND4_X1   g1364(.A1(new_n315_), .A2(new_n461_), .A3(new_n309_), .A4(new_n456_), .ZN(new_n1729_));
  NOR4_X1    g1365(.A1(new_n406_), .A2(new_n452_), .A3(new_n1728_), .A4(new_n1729_), .ZN(new_n1730_));
  OAI21_X1   g1366(.A1(new_n1727_), .A2(new_n1725_), .B(new_n1730_), .ZN(new_n1731_));
  OAI21_X1   g1367(.A1(new_n1731_), .A2(new_n1722_), .B(new_n264_), .ZN(new_n1732_));
  NAND3_X1   g1368(.A1(new_n680_), .A2(new_n521_), .A3(new_n693_), .ZN(new_n1733_));
  NOR4_X1    g1369(.A1(new_n1733_), .A2(new_n265_), .A3(new_n266_), .A4(new_n654_), .ZN(new_n1734_));
  NAND3_X1   g1370(.A1(new_n1019_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n1735_));
  NAND2_X1   g1371(.A1(new_n1735_), .A2(new_n668_), .ZN(new_n1736_));
  NAND3_X1   g1372(.A1(new_n1028_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1737_));
  NAND2_X1   g1373(.A1(new_n1737_), .A2(new_n672_), .ZN(new_n1738_));
  NAND4_X1   g1374(.A1(new_n1736_), .A2(new_n1738_), .A3(new_n276_), .A4(new_n678_), .ZN(new_n1739_));
  NAND3_X1   g1375(.A1(new_n1029_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n1740_));
  NAND2_X1   g1376(.A1(new_n1740_), .A2(new_n681_), .ZN(new_n1741_));
  NAND3_X1   g1377(.A1(new_n1005_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n1742_));
  NAND2_X1   g1378(.A1(new_n1742_), .A2(new_n685_), .ZN(new_n1743_));
  NAND4_X1   g1379(.A1(new_n1741_), .A2(new_n1743_), .A3(new_n276_), .A4(new_n691_), .ZN(new_n1744_));
  NOR4_X1    g1380(.A1(new_n542_), .A2(new_n654_), .A3(new_n1739_), .A4(new_n1744_), .ZN(new_n1745_));
  NOR3_X1    g1381(.A1(new_n1745_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1746_));
  NOR2_X1    g1382(.A1(new_n1746_), .A2(new_n1734_), .ZN(new_n1747_));
  NAND2_X1   g1383(.A1(new_n629_), .A2(new_n667_), .ZN(new_n1748_));
  NOR4_X1    g1384(.A1(new_n1748_), .A2(new_n619_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1749_));
  NOR2_X1    g1385(.A1(new_n1748_), .A2(new_n619_), .ZN(new_n1750_));
  NOR3_X1    g1386(.A1(new_n1750_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n1751_));
  NAND4_X1   g1387(.A1(new_n488_), .A2(new_n380_), .A3(new_n375_), .A4(new_n482_), .ZN(new_n1752_));
  NAND4_X1   g1388(.A1(new_n497_), .A2(new_n508_), .A3(new_n492_), .A4(new_n502_), .ZN(new_n1753_));
  NAND3_X1   g1389(.A1(new_n640_), .A2(new_n549_), .A3(new_n558_), .ZN(new_n1754_));
  NAND4_X1   g1390(.A1(new_n570_), .A2(new_n581_), .A3(new_n562_), .A4(new_n575_), .ZN(new_n1755_));
  NOR4_X1    g1391(.A1(new_n1754_), .A2(new_n1752_), .A3(new_n1755_), .A4(new_n1753_), .ZN(new_n1756_));
  OAI21_X1   g1392(.A1(new_n1751_), .A2(new_n1749_), .B(new_n1756_), .ZN(new_n1757_));
  OAI21_X1   g1393(.A1(new_n1757_), .A2(new_n1747_), .B(\shift[6] ), .ZN(new_n1758_));
  NAND2_X1   g1394(.A1(new_n1758_), .A2(new_n1732_), .ZN(\result[4] ));
  NAND4_X1   g1395(.A1(new_n732_), .A2(new_n725_), .A3(new_n976_), .A4(new_n982_), .ZN(new_n1760_));
  NOR4_X1    g1396(.A1(new_n1760_), .A2(new_n265_), .A3(new_n266_), .A4(new_n719_), .ZN(new_n1761_));
  NOR2_X1    g1397(.A1(new_n1760_), .A2(new_n719_), .ZN(new_n1762_));
  NOR3_X1    g1398(.A1(new_n1762_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1763_));
  NOR2_X1    g1399(.A1(new_n1763_), .A2(new_n1761_), .ZN(new_n1764_));
  NAND4_X1   g1400(.A1(new_n753_), .A2(new_n836_), .A3(new_n759_), .A4(new_n841_), .ZN(new_n1765_));
  NAND4_X1   g1401(.A1(new_n764_), .A2(new_n776_), .A3(new_n770_), .A4(new_n783_), .ZN(new_n1766_));
  NOR4_X1    g1402(.A1(new_n1765_), .A2(new_n1766_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1767_));
  NOR2_X1    g1403(.A1(new_n1765_), .A2(new_n1766_), .ZN(new_n1768_));
  NOR3_X1    g1404(.A1(new_n1768_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n1769_));
  NAND4_X1   g1405(.A1(new_n825_), .A2(new_n882_), .A3(new_n831_), .A4(new_n888_), .ZN(new_n1770_));
  NAND4_X1   g1406(.A1(new_n737_), .A2(new_n870_), .A3(new_n743_), .A4(new_n877_), .ZN(new_n1771_));
  NOR4_X1    g1407(.A1(new_n820_), .A2(new_n865_), .A3(new_n1770_), .A4(new_n1771_), .ZN(new_n1772_));
  OAI21_X1   g1408(.A1(new_n1769_), .A2(new_n1767_), .B(new_n1772_), .ZN(new_n1773_));
  OAI21_X1   g1409(.A1(new_n1764_), .A2(new_n1773_), .B(new_n264_), .ZN(new_n1774_));
  NAND2_X1   g1410(.A1(new_n989_), .A2(\shift[1] ), .ZN(new_n1775_));
  XOR2_X1    g1411(.A1(new_n1775_), .A2(new_n988_), .Z(new_n1776_));
  NAND4_X1   g1412(.A1(new_n1776_), .A2(new_n997_), .A3(new_n1038_), .A4(new_n1044_), .ZN(new_n1777_));
  NAND4_X1   g1413(.A1(new_n1050_), .A2(new_n1064_), .A3(new_n1057_), .A4(new_n1071_), .ZN(new_n1778_));
  NOR4_X1    g1414(.A1(new_n1777_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1778_), .ZN(new_n1779_));
  NOR2_X1    g1415(.A1(new_n1777_), .A2(new_n1778_), .ZN(new_n1780_));
  NOR3_X1    g1416(.A1(new_n1780_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n1781_));
  NOR2_X1    g1417(.A1(new_n1781_), .A2(new_n1779_), .ZN(new_n1782_));
  NAND2_X1   g1418(.A1(new_n931_), .A2(new_n936_), .ZN(new_n1783_));
  OR3_X2     g1419(.A1(new_n1031_), .A2(new_n1011_), .A3(new_n1021_), .Z(new_n1784_));
  NOR4_X1    g1420(.A1(new_n1784_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1783_), .ZN(new_n1785_));
  NOR4_X1    g1421(.A1(new_n1783_), .A2(new_n1031_), .A3(new_n1011_), .A4(new_n1021_), .ZN(new_n1786_));
  NOR3_X1    g1422(.A1(new_n1786_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1787_));
  NAND4_X1   g1423(.A1(new_n788_), .A2(new_n898_), .A3(new_n794_), .A4(new_n904_), .ZN(new_n1788_));
  NAND4_X1   g1424(.A1(new_n909_), .A2(new_n921_), .A3(new_n915_), .A4(new_n926_), .ZN(new_n1789_));
  NAND4_X1   g1425(.A1(new_n965_), .A2(new_n1076_), .A3(new_n971_), .A4(new_n1082_), .ZN(new_n1790_));
  NOR4_X1    g1426(.A1(new_n960_), .A2(new_n1788_), .A3(new_n1789_), .A4(new_n1790_), .ZN(new_n1791_));
  OAI21_X1   g1427(.A1(new_n1785_), .A2(new_n1787_), .B(new_n1791_), .ZN(new_n1792_));
  OAI21_X1   g1428(.A1(new_n1782_), .A2(new_n1792_), .B(\shift[6] ), .ZN(new_n1793_));
  NAND2_X1   g1429(.A1(new_n1793_), .A2(new_n1774_), .ZN(\result[5] ));
  NAND4_X1   g1430(.A1(new_n1118_), .A2(new_n1338_), .A3(new_n1111_), .A4(new_n1332_), .ZN(new_n1795_));
  NOR4_X1    g1431(.A1(new_n1108_), .A2(new_n1795_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1796_));
  NOR2_X1    g1432(.A1(new_n1108_), .A2(new_n1795_), .ZN(new_n1797_));
  NOR3_X1    g1433(.A1(new_n1797_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1798_));
  NOR2_X1    g1434(.A1(new_n1798_), .A2(new_n1796_), .ZN(new_n1799_));
  NAND4_X1   g1435(.A1(new_n1151_), .A2(new_n1223_), .A3(new_n1145_), .A4(new_n1215_), .ZN(new_n1800_));
  NAND4_X1   g1436(.A1(new_n1159_), .A2(new_n1170_), .A3(new_n1154_), .A4(new_n1163_), .ZN(new_n1801_));
  NOR4_X1    g1437(.A1(new_n1800_), .A2(new_n1801_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1802_));
  NOR2_X1    g1438(.A1(new_n1800_), .A2(new_n1801_), .ZN(new_n1803_));
  NOR3_X1    g1439(.A1(new_n1803_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n1804_));
  NAND4_X1   g1440(.A1(new_n1212_), .A2(new_n1260_), .A3(new_n1206_), .A4(new_n1254_), .ZN(new_n1805_));
  NAND4_X1   g1441(.A1(new_n1128_), .A2(new_n1251_), .A3(new_n1121_), .A4(new_n1246_), .ZN(new_n1806_));
  NOR4_X1    g1442(.A1(new_n1805_), .A2(new_n1203_), .A3(new_n1243_), .A4(new_n1806_), .ZN(new_n1807_));
  OAI21_X1   g1443(.A1(new_n1804_), .A2(new_n1802_), .B(new_n1807_), .ZN(new_n1808_));
  OAI21_X1   g1444(.A1(new_n1808_), .A2(new_n1799_), .B(new_n264_), .ZN(new_n1809_));
  NAND4_X1   g1445(.A1(new_n1378_), .A2(new_n1388_), .A3(new_n1373_), .A4(new_n1383_), .ZN(new_n1810_));
  NAND4_X1   g1446(.A1(new_n1396_), .A2(new_n1405_), .A3(new_n1391_), .A4(new_n1400_), .ZN(new_n1811_));
  OAI21_X1   g1447(.A1(new_n1810_), .A2(new_n1811_), .B(\shift[5] ), .ZN(new_n1812_));
  XOR2_X1    g1448(.A1(new_n1812_), .A2(new_n987_), .Z(new_n1813_));
  NAND4_X1   g1449(.A1(new_n1351_), .A2(new_n1302_), .A3(new_n1295_), .A4(new_n1346_), .ZN(new_n1814_));
  NAND4_X1   g1450(.A1(new_n1359_), .A2(new_n1370_), .A3(new_n1355_), .A4(new_n1363_), .ZN(new_n1815_));
  NOR4_X1    g1451(.A1(new_n1814_), .A2(new_n1815_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1816_));
  NOR2_X1    g1452(.A1(new_n1814_), .A2(new_n1815_), .ZN(new_n1817_));
  NOR3_X1    g1453(.A1(new_n1817_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1818_));
  NAND4_X1   g1454(.A1(new_n1274_), .A2(new_n1181_), .A3(new_n1173_), .A4(new_n1268_), .ZN(new_n1819_));
  NAND4_X1   g1455(.A1(new_n1283_), .A2(new_n1292_), .A3(new_n1277_), .A4(new_n1287_), .ZN(new_n1820_));
  NAND4_X1   g1456(.A1(new_n1329_), .A2(new_n1413_), .A3(new_n1324_), .A4(new_n1408_), .ZN(new_n1821_));
  NOR4_X1    g1457(.A1(new_n1321_), .A2(new_n1819_), .A3(new_n1820_), .A4(new_n1821_), .ZN(new_n1822_));
  OAI21_X1   g1458(.A1(new_n1818_), .A2(new_n1816_), .B(new_n1822_), .ZN(new_n1823_));
  OAI21_X1   g1459(.A1(new_n1813_), .A2(new_n1823_), .B(\shift[6] ), .ZN(new_n1824_));
  NAND2_X1   g1460(.A1(new_n1824_), .A2(new_n1809_), .ZN(\result[6] ));
  NAND4_X1   g1461(.A1(new_n1517_), .A2(new_n1513_), .A3(new_n1594_), .A4(new_n1598_), .ZN(new_n1826_));
  NOR4_X1    g1462(.A1(new_n1509_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1826_), .ZN(new_n1827_));
  NOR2_X1    g1463(.A1(new_n1509_), .A2(new_n1826_), .ZN(new_n1828_));
  NOR3_X1    g1464(.A1(new_n1828_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1829_));
  NOR2_X1    g1465(.A1(new_n1829_), .A2(new_n1827_), .ZN(new_n1830_));
  NAND4_X1   g1466(.A1(new_n1529_), .A2(new_n1487_), .A3(new_n1533_), .A4(new_n1483_), .ZN(new_n1831_));
  NAND4_X1   g1467(.A1(new_n1536_), .A2(new_n1545_), .A3(new_n1541_), .A4(new_n1550_), .ZN(new_n1832_));
  NOR4_X1    g1468(.A1(new_n1832_), .A2(new_n1831_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1833_));
  OAI21_X1   g1469(.A1(new_n1832_), .A2(new_n1831_), .B(\shift[5] ), .ZN(new_n1834_));
  NOR2_X1    g1470(.A1(new_n1834_), .A2(new_n987_), .ZN(new_n1835_));
  NAND4_X1   g1471(.A1(new_n1448_), .A2(new_n1457_), .A3(new_n1452_), .A4(new_n1461_), .ZN(new_n1836_));
  NAND4_X1   g1472(.A1(new_n1464_), .A2(new_n1468_), .A3(new_n1478_), .A4(new_n1474_), .ZN(new_n1837_));
  NAND4_X1   g1473(.A1(new_n1440_), .A2(new_n1520_), .A3(new_n1445_), .A4(new_n1524_), .ZN(new_n1838_));
  NOR4_X1    g1474(.A1(new_n1437_), .A2(new_n1836_), .A3(new_n1838_), .A4(new_n1837_), .ZN(new_n1839_));
  OAI21_X1   g1475(.A1(new_n1835_), .A2(new_n1833_), .B(new_n1839_), .ZN(new_n1840_));
  OAI21_X1   g1476(.A1(new_n1830_), .A2(new_n1840_), .B(new_n264_), .ZN(new_n1841_));
  NAND4_X1   g1477(.A1(new_n1676_), .A2(new_n1672_), .A3(new_n1681_), .A4(new_n1668_), .ZN(new_n1842_));
  NAND4_X1   g1478(.A1(new_n1684_), .A2(new_n1689_), .A3(new_n1700_), .A4(new_n1695_), .ZN(new_n1843_));
  OAI21_X1   g1479(.A1(new_n1842_), .A2(new_n1843_), .B(\shift[5] ), .ZN(new_n1844_));
  XOR2_X1    g1480(.A1(new_n1844_), .A2(new_n987_), .Z(new_n1845_));
  NAND4_X1   g1481(.A1(new_n1628_), .A2(new_n1632_), .A3(new_n1664_), .A4(new_n1659_), .ZN(new_n1846_));
  NOR4_X1    g1482(.A1(new_n1654_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1846_), .ZN(new_n1847_));
  NAND2_X1   g1483(.A1(new_n1645_), .A2(new_n1641_), .ZN(new_n1848_));
  NAND3_X1   g1484(.A1(new_n1648_), .A2(new_n1651_), .A3(new_n1652_), .ZN(new_n1849_));
  NOR3_X1    g1485(.A1(new_n1846_), .A2(new_n1848_), .A3(new_n1849_), .ZN(new_n1850_));
  NOR3_X1    g1486(.A1(new_n1850_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1851_));
  NAND4_X1   g1487(.A1(new_n1604_), .A2(new_n1559_), .A3(new_n1608_), .A4(new_n1555_), .ZN(new_n1852_));
  NAND4_X1   g1488(.A1(new_n1611_), .A2(new_n1620_), .A3(new_n1616_), .A4(new_n1625_), .ZN(new_n1853_));
  NAND4_X1   g1489(.A1(new_n1569_), .A2(new_n1703_), .A3(new_n1573_), .A4(new_n1708_), .ZN(new_n1854_));
  NAND4_X1   g1490(.A1(new_n1576_), .A2(new_n1584_), .A3(new_n1580_), .A4(new_n1589_), .ZN(new_n1855_));
  NOR4_X1    g1491(.A1(new_n1853_), .A2(new_n1854_), .A3(new_n1855_), .A4(new_n1852_), .ZN(new_n1856_));
  OAI21_X1   g1492(.A1(new_n1851_), .A2(new_n1847_), .B(new_n1856_), .ZN(new_n1857_));
  OAI21_X1   g1493(.A1(new_n1845_), .A2(new_n1857_), .B(\shift[6] ), .ZN(new_n1858_));
  NAND2_X1   g1494(.A1(new_n1858_), .A2(new_n1841_), .ZN(\result[7] ));
  NAND4_X1   g1495(.A1(new_n290_), .A2(new_n305_), .A3(new_n285_), .A4(new_n296_), .ZN(new_n1860_));
  NAND4_X1   g1496(.A1(new_n558_), .A2(new_n593_), .A3(new_n549_), .A4(new_n585_), .ZN(new_n1861_));
  NOR4_X1    g1497(.A1(new_n1860_), .A2(new_n1861_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1862_));
  NOR2_X1    g1498(.A1(new_n1860_), .A2(new_n1861_), .ZN(new_n1863_));
  NOR3_X1    g1499(.A1(new_n1863_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1864_));
  NOR2_X1    g1500(.A1(new_n1864_), .A2(new_n1862_), .ZN(new_n1865_));
  NAND4_X1   g1501(.A1(new_n428_), .A2(new_n393_), .A3(new_n388_), .A4(new_n420_), .ZN(new_n1866_));
  NOR4_X1    g1502(.A1(new_n1866_), .A2(new_n1724_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1867_));
  NOR2_X1    g1503(.A1(new_n1866_), .A2(new_n1724_), .ZN(new_n1868_));
  NOR3_X1    g1504(.A1(new_n1868_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n1869_));
  NAND4_X1   g1505(.A1(new_n405_), .A2(new_n416_), .A3(new_n397_), .A4(new_n410_), .ZN(new_n1870_));
  NAND4_X1   g1506(.A1(new_n441_), .A2(new_n474_), .A3(new_n433_), .A4(new_n465_), .ZN(new_n1871_));
  NAND4_X1   g1507(.A1(new_n451_), .A2(new_n461_), .A3(new_n445_), .A4(new_n456_), .ZN(new_n1872_));
  NAND4_X1   g1508(.A1(new_n281_), .A2(new_n315_), .A3(new_n272_), .A4(new_n309_), .ZN(new_n1873_));
  NOR4_X1    g1509(.A1(new_n1871_), .A2(new_n1873_), .A3(new_n1870_), .A4(new_n1872_), .ZN(new_n1874_));
  OAI21_X1   g1510(.A1(new_n1869_), .A2(new_n1867_), .B(new_n1874_), .ZN(new_n1875_));
  OAI21_X1   g1511(.A1(new_n1875_), .A2(new_n1865_), .B(new_n264_), .ZN(new_n1876_));
  NAND3_X1   g1512(.A1(new_n629_), .A2(new_n667_), .A3(new_n618_), .ZN(new_n1877_));
  NOR4_X1    g1513(.A1(new_n1877_), .A2(new_n265_), .A3(new_n266_), .A4(new_n654_), .ZN(new_n1878_));
  OAI21_X1   g1514(.A1(new_n1877_), .A2(new_n654_), .B(\shift[5] ), .ZN(new_n1879_));
  NOR2_X1    g1515(.A1(new_n1879_), .A2(new_n987_), .ZN(new_n1880_));
  NOR2_X1    g1516(.A1(new_n1880_), .A2(new_n1878_), .ZN(new_n1881_));
  NAND2_X1   g1517(.A1(new_n680_), .A2(new_n693_), .ZN(new_n1882_));
  NAND3_X1   g1518(.A1(new_n521_), .A2(new_n488_), .A3(new_n482_), .ZN(new_n1883_));
  NOR4_X1    g1519(.A1(new_n1883_), .A2(new_n1882_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1884_));
  NOR4_X1    g1520(.A1(new_n526_), .A2(new_n542_), .A3(new_n1739_), .A4(new_n1744_), .ZN(new_n1885_));
  NOR3_X1    g1521(.A1(new_n1885_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1886_));
  NAND4_X1   g1522(.A1(new_n380_), .A2(new_n347_), .A3(new_n341_), .A4(new_n375_), .ZN(new_n1887_));
  INV_X1     g1523(.I(new_n634_), .ZN(new_n1888_));
  NOR3_X1    g1524(.A1(new_n294_), .A2(\a[19] ), .A3(\shift[1] ), .ZN(new_n1889_));
  NOR2_X1    g1525(.A1(new_n1888_), .A2(new_n1889_), .ZN(new_n1890_));
  INV_X1     g1526(.I(new_n639_), .ZN(new_n1891_));
  NOR2_X1    g1527(.A1(new_n1890_), .A2(new_n1891_), .ZN(new_n1892_));
  NAND4_X1   g1528(.A1(new_n1892_), .A2(new_n607_), .A3(new_n601_), .A4(new_n633_), .ZN(new_n1893_));
  NOR4_X1    g1529(.A1(new_n1753_), .A2(new_n1755_), .A3(new_n1887_), .A4(new_n1893_), .ZN(new_n1894_));
  OAI21_X1   g1530(.A1(new_n1886_), .A2(new_n1884_), .B(new_n1894_), .ZN(new_n1895_));
  OAI21_X1   g1531(.A1(new_n1881_), .A2(new_n1895_), .B(\shift[6] ), .ZN(new_n1896_));
  NAND2_X1   g1532(.A1(new_n1876_), .A2(new_n1896_), .ZN(\result[8] ));
  NAND4_X1   g1533(.A1(new_n732_), .A2(new_n725_), .A3(new_n713_), .A4(new_n718_), .ZN(new_n1898_));
  NAND4_X1   g1534(.A1(new_n943_), .A2(new_n976_), .A3(new_n949_), .A4(new_n982_), .ZN(new_n1899_));
  NOR4_X1    g1535(.A1(new_n1898_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1899_), .ZN(new_n1900_));
  NOR2_X1    g1536(.A1(new_n1898_), .A2(new_n1899_), .ZN(new_n1901_));
  NOR3_X1    g1537(.A1(new_n1901_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1902_));
  NOR2_X1    g1538(.A1(new_n1902_), .A2(new_n1900_), .ZN(new_n1903_));
  NAND4_X1   g1539(.A1(new_n803_), .A2(new_n836_), .A3(new_n809_), .A4(new_n841_), .ZN(new_n1904_));
  NOR4_X1    g1540(.A1(new_n1766_), .A2(new_n1904_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1905_));
  OAI21_X1   g1541(.A1(new_n1766_), .A2(new_n1904_), .B(\shift[5] ), .ZN(new_n1906_));
  NOR2_X1    g1542(.A1(new_n1906_), .A2(new_n987_), .ZN(new_n1907_));
  NAND4_X1   g1543(.A1(new_n814_), .A2(new_n825_), .A3(new_n819_), .A4(new_n831_), .ZN(new_n1908_));
  NAND4_X1   g1544(.A1(new_n847_), .A2(new_n882_), .A3(new_n852_), .A4(new_n888_), .ZN(new_n1909_));
  NAND4_X1   g1545(.A1(new_n857_), .A2(new_n870_), .A3(new_n864_), .A4(new_n877_), .ZN(new_n1910_));
  NAND4_X1   g1546(.A1(new_n703_), .A2(new_n737_), .A3(new_n708_), .A4(new_n743_), .ZN(new_n1911_));
  NOR4_X1    g1547(.A1(new_n1908_), .A2(new_n1909_), .A3(new_n1910_), .A4(new_n1911_), .ZN(new_n1912_));
  OAI21_X1   g1548(.A1(new_n1907_), .A2(new_n1905_), .B(new_n1912_), .ZN(new_n1913_));
  OAI21_X1   g1549(.A1(new_n1903_), .A2(new_n1913_), .B(new_n264_), .ZN(new_n1914_));
  OR2_X2     g1550(.A1(new_n998_), .A2(new_n1021_), .Z(new_n1915_));
  NOR4_X1    g1551(.A1(new_n1915_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1778_), .ZN(new_n1916_));
  NOR3_X1    g1552(.A1(new_n1778_), .A2(new_n998_), .A3(new_n1021_), .ZN(new_n1917_));
  NOR3_X1    g1553(.A1(new_n1917_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n1918_));
  NOR2_X1    g1554(.A1(new_n1916_), .A2(new_n1918_), .ZN(new_n1919_));
  NAND2_X1   g1555(.A1(new_n898_), .A2(new_n904_), .ZN(new_n1920_));
  OR2_X2     g1556(.A1(new_n1031_), .A2(new_n1920_), .Z(new_n1921_));
  NAND4_X1   g1557(.A1(new_n931_), .A2(new_n1004_), .A3(new_n936_), .A4(new_n1010_), .ZN(new_n1922_));
  NOR4_X1    g1558(.A1(new_n1921_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1922_), .ZN(new_n1923_));
  NOR3_X1    g1559(.A1(new_n1922_), .A2(new_n1920_), .A3(new_n1031_), .ZN(new_n1924_));
  NOR3_X1    g1560(.A1(new_n1924_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1925_));
  NAND4_X1   g1561(.A1(new_n753_), .A2(new_n788_), .A3(new_n759_), .A4(new_n794_), .ZN(new_n1926_));
  NAND4_X1   g1562(.A1(new_n954_), .A2(new_n965_), .A3(new_n959_), .A4(new_n971_), .ZN(new_n1927_));
  NAND4_X1   g1563(.A1(new_n1038_), .A2(new_n1076_), .A3(new_n1044_), .A4(new_n1082_), .ZN(new_n1928_));
  NOR4_X1    g1564(.A1(new_n1789_), .A2(new_n1926_), .A3(new_n1927_), .A4(new_n1928_), .ZN(new_n1929_));
  OAI21_X1   g1565(.A1(new_n1923_), .A2(new_n1925_), .B(new_n1929_), .ZN(new_n1930_));
  OAI21_X1   g1566(.A1(new_n1919_), .A2(new_n1930_), .B(\shift[6] ), .ZN(new_n1931_));
  NAND2_X1   g1567(.A1(new_n1931_), .A2(new_n1914_), .ZN(\result[9] ));
  NAND4_X1   g1568(.A1(new_n1107_), .A2(new_n1118_), .A3(new_n1101_), .A4(new_n1111_), .ZN(new_n1933_));
  NAND4_X1   g1569(.A1(new_n1312_), .A2(new_n1307_), .A3(new_n1338_), .A4(new_n1332_), .ZN(new_n1934_));
  NOR4_X1    g1570(.A1(new_n1934_), .A2(new_n1933_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1935_));
  NAND2_X1   g1571(.A1(new_n1310_), .A2(new_n1308_), .ZN(new_n1936_));
  INV_X1     g1572(.I(new_n1311_), .ZN(new_n1937_));
  NAND3_X1   g1573(.A1(new_n1937_), .A2(new_n1936_), .A3(new_n1307_), .ZN(new_n1938_));
  NAND3_X1   g1574(.A1(\a[3] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1939_));
  NAND3_X1   g1575(.A1(new_n977_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n1940_));
  NAND2_X1   g1576(.A1(new_n1940_), .A2(new_n1939_), .ZN(new_n1941_));
  NAND4_X1   g1577(.A1(new_n1332_), .A2(new_n1941_), .A3(new_n276_), .A4(new_n1336_), .ZN(new_n1942_));
  NOR4_X1    g1578(.A1(new_n1133_), .A2(new_n1938_), .A3(new_n1136_), .A4(new_n1942_), .ZN(new_n1943_));
  NOR3_X1    g1579(.A1(new_n1943_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1944_));
  NOR2_X1    g1580(.A1(new_n1944_), .A2(new_n1935_), .ZN(new_n1945_));
  NAND4_X1   g1581(.A1(new_n1193_), .A2(new_n1223_), .A3(new_n1188_), .A4(new_n1215_), .ZN(new_n1946_));
  NOR4_X1    g1582(.A1(new_n1801_), .A2(new_n1946_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1947_));
  NOR2_X1    g1583(.A1(new_n1801_), .A2(new_n1946_), .ZN(new_n1948_));
  NOR3_X1    g1584(.A1(new_n1948_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n1949_));
  NAND4_X1   g1585(.A1(new_n1212_), .A2(new_n1202_), .A3(new_n1196_), .A4(new_n1206_), .ZN(new_n1950_));
  NAND4_X1   g1586(.A1(new_n1234_), .A2(new_n1260_), .A3(new_n1227_), .A4(new_n1254_), .ZN(new_n1951_));
  NAND4_X1   g1587(.A1(new_n1242_), .A2(new_n1251_), .A3(new_n1237_), .A4(new_n1246_), .ZN(new_n1952_));
  NAND4_X1   g1588(.A1(new_n1098_), .A2(new_n1128_), .A3(new_n1092_), .A4(new_n1121_), .ZN(new_n1953_));
  NOR4_X1    g1589(.A1(new_n1951_), .A2(new_n1950_), .A3(new_n1953_), .A4(new_n1952_), .ZN(new_n1954_));
  OAI21_X1   g1590(.A1(new_n1949_), .A2(new_n1947_), .B(new_n1954_), .ZN(new_n1955_));
  OAI21_X1   g1591(.A1(new_n1955_), .A2(new_n1945_), .B(new_n264_), .ZN(new_n1956_));
  NAND4_X1   g1592(.A1(new_n1351_), .A2(new_n1378_), .A3(new_n1346_), .A4(new_n1373_), .ZN(new_n1957_));
  OAI21_X1   g1593(.A1(new_n1957_), .A2(new_n1811_), .B(\shift[5] ), .ZN(new_n1958_));
  XOR2_X1    g1594(.A1(new_n1958_), .A2(new_n987_), .Z(new_n1959_));
  NAND4_X1   g1595(.A1(new_n1274_), .A2(new_n1302_), .A3(new_n1268_), .A4(new_n1295_), .ZN(new_n1960_));
  NOR4_X1    g1596(.A1(new_n1960_), .A2(new_n1815_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1961_));
  NOR2_X1    g1597(.A1(new_n1960_), .A2(new_n1815_), .ZN(new_n1962_));
  NOR3_X1    g1598(.A1(new_n1962_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1963_));
  NAND4_X1   g1599(.A1(new_n1151_), .A2(new_n1181_), .A3(new_n1145_), .A4(new_n1173_), .ZN(new_n1964_));
  NAND4_X1   g1600(.A1(new_n1320_), .A2(new_n1329_), .A3(new_n1315_), .A4(new_n1324_), .ZN(new_n1965_));
  NAND4_X1   g1601(.A1(new_n1388_), .A2(new_n1413_), .A3(new_n1383_), .A4(new_n1408_), .ZN(new_n1966_));
  NOR4_X1    g1602(.A1(new_n1820_), .A2(new_n1965_), .A3(new_n1964_), .A4(new_n1966_), .ZN(new_n1967_));
  OAI21_X1   g1603(.A1(new_n1963_), .A2(new_n1961_), .B(new_n1967_), .ZN(new_n1968_));
  OAI21_X1   g1604(.A1(new_n1959_), .A2(new_n1968_), .B(\shift[6] ), .ZN(new_n1969_));
  NAND2_X1   g1605(.A1(new_n1969_), .A2(new_n1956_), .ZN(\result[10] ));
  NAND4_X1   g1606(.A1(new_n1508_), .A2(new_n1504_), .A3(new_n1513_), .A4(new_n1517_), .ZN(new_n1971_));
  NAND4_X1   g1607(.A1(new_n1569_), .A2(new_n1573_), .A3(new_n1598_), .A4(new_n1594_), .ZN(new_n1972_));
  NOR4_X1    g1608(.A1(new_n1971_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1972_), .ZN(new_n1973_));
  NOR2_X1    g1609(.A1(new_n1971_), .A2(new_n1972_), .ZN(new_n1974_));
  NOR3_X1    g1610(.A1(new_n1974_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1975_));
  NOR2_X1    g1611(.A1(new_n1975_), .A2(new_n1973_), .ZN(new_n1976_));
  NAND4_X1   g1612(.A1(new_n1457_), .A2(new_n1461_), .A3(new_n1487_), .A4(new_n1483_), .ZN(new_n1977_));
  NOR4_X1    g1613(.A1(new_n1832_), .A2(new_n1977_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n1978_));
  OAI21_X1   g1614(.A1(new_n1832_), .A2(new_n1977_), .B(\shift[5] ), .ZN(new_n1979_));
  NOR2_X1    g1615(.A1(new_n1979_), .A2(new_n987_), .ZN(new_n1980_));
  NAND4_X1   g1616(.A1(new_n1423_), .A2(new_n1448_), .A3(new_n1428_), .A4(new_n1452_), .ZN(new_n1981_));
  NAND4_X1   g1617(.A1(new_n1431_), .A2(new_n1440_), .A3(new_n1436_), .A4(new_n1445_), .ZN(new_n1982_));
  NAND4_X1   g1618(.A1(new_n1496_), .A2(new_n1520_), .A3(new_n1501_), .A4(new_n1524_), .ZN(new_n1983_));
  NOR4_X1    g1619(.A1(new_n1981_), .A2(new_n1982_), .A3(new_n1983_), .A4(new_n1837_), .ZN(new_n1984_));
  OAI21_X1   g1620(.A1(new_n1980_), .A2(new_n1978_), .B(new_n1984_), .ZN(new_n1985_));
  OAI21_X1   g1621(.A1(new_n1976_), .A2(new_n1985_), .B(new_n264_), .ZN(new_n1986_));
  NAND4_X1   g1622(.A1(new_n1645_), .A2(new_n1672_), .A3(new_n1641_), .A4(new_n1668_), .ZN(new_n1987_));
  OAI21_X1   g1623(.A1(new_n1843_), .A2(new_n1987_), .B(\shift[5] ), .ZN(new_n1988_));
  XOR2_X1    g1624(.A1(new_n1988_), .A2(new_n987_), .Z(new_n1989_));
  NAND4_X1   g1625(.A1(new_n1653_), .A2(new_n1648_), .A3(new_n1659_), .A4(new_n1664_), .ZN(new_n1990_));
  NAND4_X1   g1626(.A1(new_n1604_), .A2(new_n1628_), .A3(new_n1608_), .A4(new_n1632_), .ZN(new_n1991_));
  NOR4_X1    g1627(.A1(new_n1990_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1991_), .ZN(new_n1992_));
  NAND2_X1   g1628(.A1(new_n1664_), .A2(new_n1659_), .ZN(new_n1993_));
  NOR3_X1    g1629(.A1(new_n1991_), .A2(new_n1849_), .A3(new_n1993_), .ZN(new_n1994_));
  NOR3_X1    g1630(.A1(new_n1994_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n1995_));
  NAND4_X1   g1631(.A1(new_n1529_), .A2(new_n1533_), .A3(new_n1559_), .A4(new_n1555_), .ZN(new_n1996_));
  NAND4_X1   g1632(.A1(new_n1676_), .A2(new_n1703_), .A3(new_n1681_), .A4(new_n1708_), .ZN(new_n1997_));
  NOR4_X1    g1633(.A1(new_n1853_), .A2(new_n1855_), .A3(new_n1997_), .A4(new_n1996_), .ZN(new_n1998_));
  OAI21_X1   g1634(.A1(new_n1995_), .A2(new_n1992_), .B(new_n1998_), .ZN(new_n1999_));
  OAI21_X1   g1635(.A1(new_n1999_), .A2(new_n1989_), .B(\shift[6] ), .ZN(new_n2000_));
  NAND2_X1   g1636(.A1(new_n2000_), .A2(new_n1986_), .ZN(\result[11] ));
  NOR4_X1    g1637(.A1(new_n571_), .A2(new_n1714_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2002_));
  NAND2_X1   g1638(.A1(new_n558_), .A2(new_n549_), .ZN(new_n2003_));
  NAND2_X1   g1639(.A1(new_n565_), .A2(new_n563_), .ZN(new_n2004_));
  NAND4_X1   g1640(.A1(new_n562_), .A2(new_n2004_), .A3(new_n276_), .A4(new_n568_), .ZN(new_n2005_));
  NOR4_X1    g1641(.A1(new_n2003_), .A2(new_n329_), .A3(new_n2005_), .A4(new_n1719_), .ZN(new_n2006_));
  NOR3_X1    g1642(.A1(new_n2006_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2007_));
  NOR2_X1    g1643(.A1(new_n2007_), .A2(new_n2002_), .ZN(new_n2008_));
  NAND4_X1   g1644(.A1(new_n428_), .A2(new_n371_), .A3(new_n365_), .A4(new_n420_), .ZN(new_n2009_));
  NOR4_X1    g1645(.A1(new_n406_), .A2(new_n2009_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2010_));
  INV_X1     g1646(.I(new_n368_), .ZN(new_n2011_));
  NAND2_X1   g1647(.A1(new_n2011_), .A2(new_n366_), .ZN(new_n2012_));
  INV_X1     g1648(.I(new_n370_), .ZN(new_n2013_));
  NAND3_X1   g1649(.A1(new_n2012_), .A2(new_n2013_), .A3(new_n365_), .ZN(new_n2014_));
  NAND2_X1   g1650(.A1(new_n391_), .A2(new_n389_), .ZN(new_n2015_));
  NOR2_X1    g1651(.A1(new_n1220_), .A2(new_n804_), .ZN(new_n2016_));
  NAND4_X1   g1652(.A1(new_n388_), .A2(new_n276_), .A3(new_n2015_), .A4(new_n2016_), .ZN(new_n2017_));
  NAND2_X1   g1653(.A1(new_n400_), .A2(new_n398_), .ZN(new_n2018_));
  NAND4_X1   g1654(.A1(new_n397_), .A2(new_n2018_), .A3(new_n276_), .A4(new_n403_), .ZN(new_n2019_));
  NAND2_X1   g1655(.A1(new_n423_), .A2(new_n421_), .ZN(new_n2020_));
  NAND4_X1   g1656(.A1(new_n420_), .A2(new_n2020_), .A3(new_n276_), .A4(new_n426_), .ZN(new_n2021_));
  NOR4_X1    g1657(.A1(new_n2014_), .A2(new_n2017_), .A3(new_n2019_), .A4(new_n2021_), .ZN(new_n2022_));
  NOR3_X1    g1658(.A1(new_n2022_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2023_));
  NOR4_X1    g1659(.A1(new_n291_), .A2(new_n452_), .A3(new_n1728_), .A4(new_n1729_), .ZN(new_n2024_));
  OAI21_X1   g1660(.A1(new_n2023_), .A2(new_n2010_), .B(new_n2024_), .ZN(new_n2025_));
  OAI21_X1   g1661(.A1(new_n2025_), .A2(new_n2008_), .B(new_n264_), .ZN(new_n2026_));
  NAND3_X1   g1662(.A1(new_n629_), .A2(new_n680_), .A3(new_n667_), .ZN(new_n2027_));
  NOR4_X1    g1663(.A1(new_n2027_), .A2(new_n265_), .A3(new_n266_), .A4(new_n654_), .ZN(new_n2028_));
  INV_X1     g1664(.I(new_n622_), .ZN(new_n2029_));
  NAND2_X1   g1665(.A1(new_n2029_), .A2(new_n620_), .ZN(new_n2030_));
  NAND3_X1   g1666(.A1(new_n1066_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n2031_));
  NAND2_X1   g1667(.A1(new_n2031_), .A2(new_n624_), .ZN(new_n2032_));
  NOR2_X1    g1668(.A1(new_n323_), .A2(new_n628_), .ZN(new_n2033_));
  NAND3_X1   g1669(.A1(new_n2030_), .A2(new_n2032_), .A3(new_n2033_), .ZN(new_n2034_));
  INV_X1     g1670(.I(new_n657_), .ZN(new_n2035_));
  NAND2_X1   g1671(.A1(new_n2035_), .A2(new_n655_), .ZN(new_n2036_));
  NAND3_X1   g1672(.A1(new_n992_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n2037_));
  NAND2_X1   g1673(.A1(new_n2037_), .A2(new_n659_), .ZN(new_n2038_));
  NAND3_X1   g1674(.A1(new_n2036_), .A2(new_n2038_), .A3(new_n665_), .ZN(new_n2039_));
  NOR4_X1    g1675(.A1(new_n2034_), .A2(new_n2039_), .A3(new_n654_), .A4(new_n1739_), .ZN(new_n2040_));
  NOR3_X1    g1676(.A1(new_n2040_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2041_));
  NOR2_X1    g1677(.A1(new_n2041_), .A2(new_n2028_), .ZN(new_n2042_));
  NAND3_X1   g1678(.A1(new_n693_), .A2(new_n488_), .A3(new_n482_), .ZN(new_n2043_));
  NAND3_X1   g1679(.A1(new_n521_), .A2(new_n497_), .A3(new_n492_), .ZN(new_n2044_));
  NOR4_X1    g1680(.A1(new_n2044_), .A2(new_n2043_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2045_));
  NOR4_X1    g1681(.A1(new_n526_), .A2(new_n529_), .A3(new_n542_), .A4(new_n1744_), .ZN(new_n2046_));
  NOR3_X1    g1682(.A1(new_n2046_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2047_));
  NAND4_X1   g1683(.A1(new_n380_), .A2(new_n508_), .A3(new_n375_), .A4(new_n502_), .ZN(new_n2048_));
  NAND4_X1   g1684(.A1(new_n1892_), .A2(new_n581_), .A3(new_n575_), .A4(new_n633_), .ZN(new_n2049_));
  NOR4_X1    g1685(.A1(new_n619_), .A2(new_n2048_), .A3(new_n2049_), .A4(new_n361_), .ZN(new_n2050_));
  OAI21_X1   g1686(.A1(new_n2047_), .A2(new_n2045_), .B(new_n2050_), .ZN(new_n2051_));
  OAI21_X1   g1687(.A1(new_n2051_), .A2(new_n2042_), .B(\shift[6] ), .ZN(new_n2052_));
  NAND2_X1   g1688(.A1(new_n2052_), .A2(new_n2026_), .ZN(\result[12] ));
  NOR4_X1    g1689(.A1(new_n1760_), .A2(new_n265_), .A3(new_n266_), .A4(new_n960_), .ZN(new_n2054_));
  NOR2_X1    g1690(.A1(new_n1760_), .A2(new_n960_), .ZN(new_n2055_));
  NOR3_X1    g1691(.A1(new_n2055_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2056_));
  NOR2_X1    g1692(.A1(new_n2056_), .A2(new_n2054_), .ZN(new_n2057_));
  NAND4_X1   g1693(.A1(new_n776_), .A2(new_n836_), .A3(new_n783_), .A4(new_n841_), .ZN(new_n2058_));
  NOR4_X1    g1694(.A1(new_n820_), .A2(new_n2058_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2059_));
  OAI21_X1   g1695(.A1(new_n820_), .A2(new_n2058_), .B(\shift[5] ), .ZN(new_n2060_));
  NOR2_X1    g1696(.A1(new_n2060_), .A2(new_n987_), .ZN(new_n2061_));
  NOR4_X1    g1697(.A1(new_n719_), .A2(new_n865_), .A3(new_n1770_), .A4(new_n1771_), .ZN(new_n2062_));
  OAI21_X1   g1698(.A1(new_n2061_), .A2(new_n2059_), .B(new_n2062_), .ZN(new_n2063_));
  OAI21_X1   g1699(.A1(new_n2057_), .A2(new_n2063_), .B(new_n264_), .ZN(new_n2064_));
  NAND2_X1   g1700(.A1(new_n1064_), .A2(new_n1071_), .ZN(new_n2065_));
  NOR4_X1    g1701(.A1(new_n998_), .A2(new_n1031_), .A3(new_n2065_), .A4(new_n1021_), .ZN(new_n2066_));
  NOR2_X1    g1702(.A1(new_n2066_), .A2(new_n266_), .ZN(new_n2067_));
  NOR2_X1    g1703(.A1(new_n2067_), .A2(new_n893_), .ZN(new_n2068_));
  NOR3_X1    g1704(.A1(new_n2066_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2069_));
  NOR2_X1    g1705(.A1(new_n2068_), .A2(new_n2069_), .ZN(new_n2070_));
  NOR4_X1    g1706(.A1(new_n916_), .A2(new_n1922_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2071_));
  NOR2_X1    g1707(.A1(new_n916_), .A2(new_n1922_), .ZN(new_n2072_));
  NOR3_X1    g1708(.A1(new_n2072_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2073_));
  NAND4_X1   g1709(.A1(new_n788_), .A2(new_n921_), .A3(new_n794_), .A4(new_n926_), .ZN(new_n2074_));
  NOR4_X1    g1710(.A1(new_n771_), .A2(new_n1058_), .A3(new_n1790_), .A4(new_n2074_), .ZN(new_n2075_));
  OAI21_X1   g1711(.A1(new_n2073_), .A2(new_n2071_), .B(new_n2075_), .ZN(new_n2076_));
  OAI21_X1   g1712(.A1(new_n2070_), .A2(new_n2076_), .B(\shift[6] ), .ZN(new_n2077_));
  NAND2_X1   g1713(.A1(new_n2077_), .A2(new_n2064_), .ZN(\result[13] ));
  NOR4_X1    g1714(.A1(new_n1321_), .A2(new_n1795_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2079_));
  NAND2_X1   g1715(.A1(new_n1318_), .A2(new_n1316_), .ZN(new_n2080_));
  INV_X1     g1716(.I(new_n1319_), .ZN(new_n2081_));
  NAND3_X1   g1717(.A1(new_n2081_), .A2(new_n2080_), .A3(new_n1315_), .ZN(new_n2082_));
  NOR4_X1    g1718(.A1(new_n1938_), .A2(new_n2082_), .A3(new_n1136_), .A4(new_n1942_), .ZN(new_n2083_));
  NOR3_X1    g1719(.A1(new_n2083_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2084_));
  NOR2_X1    g1720(.A1(new_n2084_), .A2(new_n2079_), .ZN(new_n2085_));
  NAND4_X1   g1721(.A1(new_n1170_), .A2(new_n1223_), .A3(new_n1163_), .A4(new_n1215_), .ZN(new_n2086_));
  NOR4_X1    g1722(.A1(new_n1203_), .A2(new_n2086_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2087_));
  NAND2_X1   g1723(.A1(new_n1170_), .A2(new_n1163_), .ZN(new_n2088_));
  NAND2_X1   g1724(.A1(new_n1191_), .A2(new_n1189_), .ZN(new_n2089_));
  NOR2_X1    g1725(.A1(new_n804_), .A2(new_n401_), .ZN(new_n2090_));
  NAND4_X1   g1726(.A1(new_n2089_), .A2(new_n276_), .A3(new_n1188_), .A4(new_n2090_), .ZN(new_n2091_));
  NAND2_X1   g1727(.A1(new_n1199_), .A2(new_n1197_), .ZN(new_n2092_));
  NAND4_X1   g1728(.A1(new_n2092_), .A2(new_n276_), .A3(new_n1196_), .A4(new_n1200_), .ZN(new_n2093_));
  NAND3_X1   g1729(.A1(new_n422_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n2094_));
  NAND2_X1   g1730(.A1(new_n2094_), .A2(new_n1216_), .ZN(new_n2095_));
  NAND4_X1   g1731(.A1(new_n1215_), .A2(new_n2095_), .A3(new_n276_), .A4(new_n1221_), .ZN(new_n2096_));
  NOR4_X1    g1732(.A1(new_n2088_), .A2(new_n2091_), .A3(new_n2093_), .A4(new_n2096_), .ZN(new_n2097_));
  NOR3_X1    g1733(.A1(new_n2097_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2098_));
  NOR4_X1    g1734(.A1(new_n1805_), .A2(new_n1108_), .A3(new_n1243_), .A4(new_n1806_), .ZN(new_n2099_));
  OAI21_X1   g1735(.A1(new_n2098_), .A2(new_n2087_), .B(new_n2099_), .ZN(new_n2100_));
  OAI21_X1   g1736(.A1(new_n2100_), .A2(new_n2085_), .B(new_n264_), .ZN(new_n2101_));
  NAND4_X1   g1737(.A1(new_n1378_), .A2(new_n1405_), .A3(new_n1373_), .A4(new_n1400_), .ZN(new_n2102_));
  NOR4_X1    g1738(.A1(new_n1360_), .A2(new_n2102_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2103_));
  NOR2_X1    g1739(.A1(new_n1360_), .A2(new_n2102_), .ZN(new_n2104_));
  NOR3_X1    g1740(.A1(new_n2104_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2105_));
  NOR2_X1    g1741(.A1(new_n2105_), .A2(new_n2103_), .ZN(new_n2106_));
  NAND4_X1   g1742(.A1(new_n1302_), .A2(new_n1370_), .A3(new_n1295_), .A4(new_n1363_), .ZN(new_n2107_));
  NOR4_X1    g1743(.A1(new_n1284_), .A2(new_n2107_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2108_));
  NAND2_X1   g1744(.A1(new_n1274_), .A2(new_n1268_), .ZN(new_n2109_));
  NAND2_X1   g1745(.A1(new_n1280_), .A2(new_n1278_), .ZN(new_n2110_));
  NAND4_X1   g1746(.A1(new_n2110_), .A2(new_n276_), .A3(new_n1277_), .A4(new_n1281_), .ZN(new_n2111_));
  INV_X1     g1747(.I(new_n1298_), .ZN(new_n2112_));
  NAND2_X1   g1748(.A1(new_n2112_), .A2(new_n1296_), .ZN(new_n2113_));
  NAND4_X1   g1749(.A1(new_n2113_), .A2(new_n276_), .A3(new_n1295_), .A4(new_n1300_), .ZN(new_n2114_));
  NAND3_X1   g1750(.A1(new_n1005_), .A2(new_n294_), .A3(\shift[1] ), .ZN(new_n2115_));
  NAND2_X1   g1751(.A1(new_n2115_), .A2(new_n1364_), .ZN(new_n2116_));
  NAND4_X1   g1752(.A1(new_n1363_), .A2(new_n2116_), .A3(new_n276_), .A4(new_n1368_), .ZN(new_n2117_));
  NOR4_X1    g1753(.A1(new_n2109_), .A2(new_n2111_), .A3(new_n2114_), .A4(new_n2117_), .ZN(new_n2118_));
  NOR3_X1    g1754(.A1(new_n2118_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2119_));
  NAND4_X1   g1755(.A1(new_n1292_), .A2(new_n1181_), .A3(new_n1173_), .A4(new_n1287_), .ZN(new_n2120_));
  NOR4_X1    g1756(.A1(new_n1160_), .A2(new_n1397_), .A3(new_n1821_), .A4(new_n2120_), .ZN(new_n2121_));
  OAI21_X1   g1757(.A1(new_n2119_), .A2(new_n2108_), .B(new_n2121_), .ZN(new_n2122_));
  OAI21_X1   g1758(.A1(new_n2122_), .A2(new_n2106_), .B(\shift[6] ), .ZN(new_n2123_));
  NAND2_X1   g1759(.A1(new_n2123_), .A2(new_n2101_), .ZN(\result[14] ));
  NOR4_X1    g1760(.A1(new_n1826_), .A2(new_n1581_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2125_));
  NOR2_X1    g1761(.A1(new_n1826_), .A2(new_n1581_), .ZN(new_n2126_));
  NOR3_X1    g1762(.A1(new_n2126_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2127_));
  NOR2_X1    g1763(.A1(new_n2127_), .A2(new_n2125_), .ZN(new_n2128_));
  NAND4_X1   g1764(.A1(new_n1545_), .A2(new_n1487_), .A3(new_n1550_), .A4(new_n1483_), .ZN(new_n2129_));
  NOR4_X1    g1765(.A1(new_n1469_), .A2(new_n2129_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2130_));
  OAI21_X1   g1766(.A1(new_n1469_), .A2(new_n2129_), .B(\shift[5] ), .ZN(new_n2131_));
  NOR2_X1    g1767(.A1(new_n2131_), .A2(new_n987_), .ZN(new_n2132_));
  NAND4_X1   g1768(.A1(new_n1448_), .A2(new_n1452_), .A3(new_n1478_), .A4(new_n1474_), .ZN(new_n2133_));
  NOR4_X1    g1769(.A1(new_n1509_), .A2(new_n1437_), .A3(new_n1838_), .A4(new_n2133_), .ZN(new_n2134_));
  OAI21_X1   g1770(.A1(new_n2132_), .A2(new_n2130_), .B(new_n2134_), .ZN(new_n2135_));
  OAI21_X1   g1771(.A1(new_n2135_), .A2(new_n2128_), .B(new_n264_), .ZN(new_n2136_));
  NAND4_X1   g1772(.A1(new_n1672_), .A2(new_n1700_), .A3(new_n1668_), .A4(new_n1695_), .ZN(new_n2137_));
  NOR4_X1    g1773(.A1(new_n1654_), .A2(new_n265_), .A3(new_n266_), .A4(new_n2137_), .ZN(new_n2138_));
  NOR3_X1    g1774(.A1(new_n2137_), .A2(new_n1848_), .A3(new_n1849_), .ZN(new_n2139_));
  NOR3_X1    g1775(.A1(new_n2139_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2140_));
  NOR2_X1    g1776(.A1(new_n2140_), .A2(new_n2138_), .ZN(new_n2141_));
  NOR4_X1    g1777(.A1(new_n1617_), .A2(new_n1846_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2142_));
  NOR2_X1    g1778(.A1(new_n1617_), .A2(new_n1846_), .ZN(new_n2143_));
  NOR3_X1    g1779(.A1(new_n2143_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2144_));
  NAND4_X1   g1780(.A1(new_n1620_), .A2(new_n1559_), .A3(new_n1625_), .A4(new_n1555_), .ZN(new_n2145_));
  NAND4_X1   g1781(.A1(new_n1584_), .A2(new_n1703_), .A3(new_n1589_), .A4(new_n1708_), .ZN(new_n2146_));
  NOR4_X1    g1782(.A1(new_n1542_), .A2(new_n1690_), .A3(new_n2146_), .A4(new_n2145_), .ZN(new_n2147_));
  OAI21_X1   g1783(.A1(new_n2144_), .A2(new_n2142_), .B(new_n2147_), .ZN(new_n2148_));
  OAI21_X1   g1784(.A1(new_n2148_), .A2(new_n2141_), .B(\shift[6] ), .ZN(new_n2149_));
  NAND2_X1   g1785(.A1(new_n2136_), .A2(new_n2149_), .ZN(\result[15] ));
  NOR4_X1    g1786(.A1(new_n406_), .A2(new_n429_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2151_));
  NOR2_X1    g1787(.A1(new_n406_), .A2(new_n429_), .ZN(new_n2152_));
  NOR3_X1    g1788(.A1(new_n2152_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2153_));
  NOR2_X1    g1789(.A1(new_n2153_), .A2(new_n2151_), .ZN(new_n2154_));
  NOR4_X1    g1790(.A1(new_n452_), .A2(new_n571_), .A3(new_n475_), .A4(new_n594_), .ZN(new_n2155_));
  OAI21_X1   g1791(.A1(new_n336_), .A2(new_n317_), .B(new_n2155_), .ZN(new_n2156_));
  OAI21_X1   g1792(.A1(new_n2154_), .A2(new_n2156_), .B(new_n264_), .ZN(new_n2157_));
  NAND2_X1   g1793(.A1(new_n607_), .A2(new_n601_), .ZN(new_n2158_));
  INV_X1     g1794(.I(new_n610_), .ZN(new_n2159_));
  NAND2_X1   g1795(.A1(new_n2159_), .A2(new_n608_), .ZN(new_n2160_));
  NAND3_X1   g1796(.A1(new_n1052_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n2161_));
  NAND2_X1   g1797(.A1(new_n2161_), .A2(new_n612_), .ZN(new_n2162_));
  NAND4_X1   g1798(.A1(new_n2160_), .A2(new_n276_), .A3(new_n2162_), .A4(new_n616_), .ZN(new_n2163_));
  NAND3_X1   g1799(.A1(new_n633_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n2164_));
  NOR4_X1    g1800(.A1(new_n2158_), .A2(new_n2163_), .A3(new_n2034_), .A4(new_n2164_), .ZN(new_n2165_));
  NOR3_X1    g1801(.A1(new_n381_), .A2(new_n361_), .A3(new_n893_), .ZN(new_n2166_));
  NOR3_X1    g1802(.A1(new_n2166_), .A2(new_n2165_), .A3(new_n1265_), .ZN(new_n2167_));
  NOR4_X1    g1803(.A1(new_n381_), .A2(new_n361_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2168_));
  NOR2_X1    g1804(.A1(new_n2167_), .A2(new_n2168_), .ZN(new_n2169_));
  NOR2_X1    g1805(.A1(new_n694_), .A2(new_n654_), .ZN(new_n2170_));
  NOR3_X1    g1806(.A1(new_n498_), .A2(new_n522_), .A3(new_n893_), .ZN(new_n2171_));
  NOR3_X1    g1807(.A1(new_n2171_), .A2(new_n2170_), .A3(new_n1265_), .ZN(new_n2172_));
  NOR4_X1    g1808(.A1(new_n498_), .A2(new_n522_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2173_));
  NOR2_X1    g1809(.A1(new_n2172_), .A2(new_n2173_), .ZN(new_n2174_));
  OAI21_X1   g1810(.A1(new_n2174_), .A2(new_n2169_), .B(\shift[6] ), .ZN(new_n2175_));
  NAND2_X1   g1811(.A1(new_n2175_), .A2(new_n2157_), .ZN(\result[16] ));
  OAI21_X1   g1812(.A1(new_n820_), .A2(new_n842_), .B(\shift[5] ), .ZN(new_n2177_));
  XOR2_X1    g1813(.A1(new_n2177_), .A2(new_n987_), .Z(new_n2178_));
  NOR4_X1    g1814(.A1(new_n865_), .A2(new_n889_), .A3(new_n960_), .A4(new_n983_), .ZN(new_n2179_));
  OAI21_X1   g1815(.A1(new_n747_), .A2(new_n745_), .B(new_n2179_), .ZN(new_n2180_));
  OAI21_X1   g1816(.A1(new_n2180_), .A2(new_n2178_), .B(new_n264_), .ZN(new_n2181_));
  NOR2_X1    g1817(.A1(new_n1032_), .A2(new_n266_), .ZN(new_n2182_));
  NOR2_X1    g1818(.A1(new_n2182_), .A2(new_n893_), .ZN(new_n2183_));
  NOR3_X1    g1819(.A1(new_n1032_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2184_));
  NOR2_X1    g1820(.A1(new_n2183_), .A2(new_n2184_), .ZN(new_n2185_));
  NOR4_X1    g1821(.A1(new_n771_), .A2(new_n795_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2186_));
  NOR3_X1    g1822(.A1(new_n797_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2187_));
  NOR4_X1    g1823(.A1(new_n916_), .A2(new_n937_), .A3(new_n1058_), .A4(new_n1083_), .ZN(new_n2188_));
  OAI21_X1   g1824(.A1(new_n2187_), .A2(new_n2186_), .B(new_n2188_), .ZN(new_n2189_));
  OAI21_X1   g1825(.A1(new_n2185_), .A2(new_n2189_), .B(\shift[6] ), .ZN(new_n2190_));
  NAND2_X1   g1826(.A1(new_n2181_), .A2(new_n2190_), .ZN(\result[17] ));
  NOR4_X1    g1827(.A1(new_n1203_), .A2(new_n1224_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2192_));
  NOR2_X1    g1828(.A1(new_n1203_), .A2(new_n1224_), .ZN(new_n2193_));
  NOR3_X1    g1829(.A1(new_n2193_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2194_));
  NOR2_X1    g1830(.A1(new_n2194_), .A2(new_n2192_), .ZN(new_n2195_));
  NOR4_X1    g1831(.A1(new_n1243_), .A2(new_n1261_), .A3(new_n1321_), .A4(new_n1339_), .ZN(new_n2196_));
  OAI21_X1   g1832(.A1(new_n1141_), .A2(new_n1130_), .B(new_n2196_), .ZN(new_n2197_));
  OAI21_X1   g1833(.A1(new_n2195_), .A2(new_n2197_), .B(new_n264_), .ZN(new_n2198_));
  NOR4_X1    g1834(.A1(new_n1360_), .A2(new_n1379_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2199_));
  NOR2_X1    g1835(.A1(new_n1360_), .A2(new_n1379_), .ZN(new_n2200_));
  NOR3_X1    g1836(.A1(new_n2200_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2201_));
  NOR2_X1    g1837(.A1(new_n2201_), .A2(new_n2199_), .ZN(new_n2202_));
  NOR4_X1    g1838(.A1(new_n1160_), .A2(new_n1182_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2203_));
  NOR3_X1    g1839(.A1(new_n1184_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2204_));
  NOR4_X1    g1840(.A1(new_n1284_), .A2(new_n1303_), .A3(new_n1397_), .A4(new_n1414_), .ZN(new_n2205_));
  OAI21_X1   g1841(.A1(new_n2204_), .A2(new_n2203_), .B(new_n2205_), .ZN(new_n2206_));
  OAI21_X1   g1842(.A1(new_n2206_), .A2(new_n2202_), .B(\shift[6] ), .ZN(new_n2207_));
  NAND2_X1   g1843(.A1(new_n2207_), .A2(new_n2198_), .ZN(\result[18] ));
  NOR4_X1    g1844(.A1(new_n1509_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1525_), .ZN(new_n2209_));
  NOR2_X1    g1845(.A1(new_n1509_), .A2(new_n1525_), .ZN(new_n2210_));
  NOR3_X1    g1846(.A1(new_n2210_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2211_));
  NOR2_X1    g1847(.A1(new_n2211_), .A2(new_n2209_), .ZN(new_n2212_));
  NOR4_X1    g1848(.A1(new_n1437_), .A2(new_n1453_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2213_));
  OAI21_X1   g1849(.A1(new_n1437_), .A2(new_n1453_), .B(\shift[5] ), .ZN(new_n2214_));
  NOR2_X1    g1850(.A1(new_n2214_), .A2(new_n987_), .ZN(new_n2215_));
  NOR4_X1    g1851(.A1(new_n1469_), .A2(new_n1581_), .A3(new_n1599_), .A4(new_n1488_), .ZN(new_n2216_));
  OAI21_X1   g1852(.A1(new_n2215_), .A2(new_n2213_), .B(new_n2216_), .ZN(new_n2217_));
  OAI21_X1   g1853(.A1(new_n2212_), .A2(new_n2217_), .B(new_n264_), .ZN(new_n2218_));
  NOR4_X1    g1854(.A1(new_n1654_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1673_), .ZN(new_n2219_));
  NOR3_X1    g1855(.A1(new_n1673_), .A2(new_n1848_), .A3(new_n1849_), .ZN(new_n2220_));
  NOR3_X1    g1856(.A1(new_n2220_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2221_));
  NOR2_X1    g1857(.A1(new_n2221_), .A2(new_n2219_), .ZN(new_n2222_));
  NOR4_X1    g1858(.A1(new_n1542_), .A2(new_n1560_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2223_));
  NOR3_X1    g1859(.A1(new_n1563_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2224_));
  NOR4_X1    g1860(.A1(new_n1617_), .A2(new_n1690_), .A3(new_n1633_), .A4(new_n1709_), .ZN(new_n2225_));
  OAI21_X1   g1861(.A1(new_n2224_), .A2(new_n2223_), .B(new_n2225_), .ZN(new_n2226_));
  OAI21_X1   g1862(.A1(new_n2226_), .A2(new_n2222_), .B(\shift[6] ), .ZN(new_n2227_));
  NAND2_X1   g1863(.A1(new_n2218_), .A2(new_n2227_), .ZN(\result[19] ));
  NOR4_X1    g1864(.A1(new_n406_), .A2(new_n1728_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2229_));
  NOR2_X1    g1865(.A1(new_n406_), .A2(new_n1728_), .ZN(new_n2230_));
  NOR3_X1    g1866(.A1(new_n2230_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2231_));
  NOR2_X1    g1867(.A1(new_n2231_), .A2(new_n2229_), .ZN(new_n2232_));
  NOR4_X1    g1868(.A1(new_n1754_), .A2(new_n452_), .A3(new_n1755_), .A4(new_n1729_), .ZN(new_n2233_));
  OAI21_X1   g1869(.A1(new_n1721_), .A2(new_n1715_), .B(new_n2233_), .ZN(new_n2234_));
  OAI21_X1   g1870(.A1(new_n2232_), .A2(new_n2234_), .B(new_n264_), .ZN(new_n2235_));
  NOR4_X1    g1871(.A1(new_n1752_), .A2(new_n1753_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2236_));
  NOR2_X1    g1872(.A1(new_n1752_), .A2(new_n1753_), .ZN(new_n2237_));
  NOR3_X1    g1873(.A1(new_n2237_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2238_));
  NOR2_X1    g1874(.A1(new_n2238_), .A2(new_n2236_), .ZN(new_n2239_));
  NOR4_X1    g1875(.A1(new_n1733_), .A2(new_n1748_), .A3(new_n619_), .A4(new_n654_), .ZN(new_n2240_));
  OAI21_X1   g1876(.A1(new_n1727_), .A2(new_n1725_), .B(new_n2240_), .ZN(new_n2241_));
  OAI21_X1   g1877(.A1(new_n2241_), .A2(new_n2239_), .B(\shift[6] ), .ZN(new_n2242_));
  NAND2_X1   g1878(.A1(new_n2242_), .A2(new_n2235_), .ZN(\result[20] ));
  OAI21_X1   g1879(.A1(new_n820_), .A2(new_n1770_), .B(\shift[5] ), .ZN(new_n2244_));
  XOR2_X1    g1880(.A1(new_n2244_), .A2(new_n987_), .Z(new_n2245_));
  NOR4_X1    g1881(.A1(new_n865_), .A2(new_n960_), .A3(new_n1771_), .A4(new_n1790_), .ZN(new_n2246_));
  OAI21_X1   g1882(.A1(new_n1763_), .A2(new_n1761_), .B(new_n2246_), .ZN(new_n2247_));
  OAI21_X1   g1883(.A1(new_n2247_), .A2(new_n2245_), .B(new_n264_), .ZN(new_n2248_));
  OAI21_X1   g1884(.A1(new_n1788_), .A2(new_n1789_), .B(\shift[4] ), .ZN(new_n2249_));
  XOR2_X1    g1885(.A1(new_n2249_), .A2(new_n987_), .Z(new_n2250_));
  NOR4_X1    g1886(.A1(new_n1784_), .A2(new_n1783_), .A3(new_n1777_), .A4(new_n1778_), .ZN(new_n2251_));
  OAI21_X1   g1887(.A1(new_n1767_), .A2(new_n1769_), .B(new_n2251_), .ZN(new_n2252_));
  OAI21_X1   g1888(.A1(new_n2252_), .A2(new_n2250_), .B(\shift[6] ), .ZN(new_n2253_));
  NAND2_X1   g1889(.A1(new_n2253_), .A2(new_n2248_), .ZN(\result[21] ));
  NOR4_X1    g1890(.A1(new_n1805_), .A2(new_n1203_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2255_));
  NAND2_X1   g1891(.A1(new_n1209_), .A2(new_n1207_), .ZN(new_n2256_));
  NAND4_X1   g1892(.A1(new_n2256_), .A2(new_n276_), .A3(new_n1206_), .A4(new_n1210_), .ZN(new_n2257_));
  NAND2_X1   g1893(.A1(new_n1257_), .A2(new_n1255_), .ZN(new_n2258_));
  NAND4_X1   g1894(.A1(new_n2258_), .A2(new_n276_), .A3(new_n1254_), .A4(new_n1258_), .ZN(new_n2259_));
  NOR4_X1    g1895(.A1(new_n2091_), .A2(new_n2093_), .A3(new_n2257_), .A4(new_n2259_), .ZN(new_n2260_));
  NOR3_X1    g1896(.A1(new_n2260_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2261_));
  NOR2_X1    g1897(.A1(new_n2261_), .A2(new_n2255_), .ZN(new_n2262_));
  NOR4_X1    g1898(.A1(new_n1321_), .A2(new_n1243_), .A3(new_n1821_), .A4(new_n1806_), .ZN(new_n2263_));
  OAI21_X1   g1899(.A1(new_n1798_), .A2(new_n1796_), .B(new_n2263_), .ZN(new_n2264_));
  OAI21_X1   g1900(.A1(new_n2264_), .A2(new_n2262_), .B(new_n264_), .ZN(new_n2265_));
  NOR4_X1    g1901(.A1(new_n1820_), .A2(new_n1819_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2266_));
  NOR2_X1    g1902(.A1(new_n1820_), .A2(new_n1819_), .ZN(new_n2267_));
  NOR3_X1    g1903(.A1(new_n2267_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2268_));
  NOR2_X1    g1904(.A1(new_n2268_), .A2(new_n2266_), .ZN(new_n2269_));
  NOR4_X1    g1905(.A1(new_n1814_), .A2(new_n1815_), .A3(new_n1810_), .A4(new_n1811_), .ZN(new_n2270_));
  OAI21_X1   g1906(.A1(new_n1804_), .A2(new_n1802_), .B(new_n2270_), .ZN(new_n2271_));
  OAI21_X1   g1907(.A1(new_n2271_), .A2(new_n2269_), .B(\shift[6] ), .ZN(new_n2272_));
  NAND2_X1   g1908(.A1(new_n2272_), .A2(new_n2265_), .ZN(\result[22] ));
  NOR3_X1    g1909(.A1(new_n1836_), .A2(new_n1837_), .A3(new_n893_), .ZN(new_n2274_));
  OAI21_X1   g1910(.A1(new_n1854_), .A2(new_n1855_), .B(new_n984_), .ZN(new_n2275_));
  XOR2_X1    g1911(.A1(new_n2275_), .A2(new_n2274_), .Z(new_n2276_));
  OAI21_X1   g1912(.A1(new_n1437_), .A2(new_n1838_), .B(new_n984_), .ZN(new_n2277_));
  AOI21_X1   g1913(.A1(new_n1828_), .A2(new_n987_), .B(new_n2277_), .ZN(new_n2278_));
  NOR4_X1    g1914(.A1(new_n1509_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1826_), .ZN(new_n2280_));
  NOR2_X1    g1915(.A1(new_n2278_), .A2(new_n2280_), .ZN(new_n2281_));
  OAI21_X1   g1916(.A1(new_n2276_), .A2(new_n2281_), .B(new_n264_), .ZN(new_n2282_));
  NOR2_X1    g1917(.A1(new_n265_), .A2(\shift[5] ), .ZN(new_n2283_));
  OAI21_X1   g1918(.A1(new_n1853_), .A2(new_n1852_), .B(new_n2283_), .ZN(new_n2284_));
  AOI21_X1   g1919(.A1(new_n987_), .A2(new_n1850_), .B(new_n2284_), .ZN(new_n2285_));
  NOR4_X1    g1920(.A1(new_n1654_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1846_), .ZN(new_n2287_));
  NOR2_X1    g1921(.A1(new_n2285_), .A2(new_n2287_), .ZN(new_n2288_));
  NOR3_X1    g1922(.A1(new_n1832_), .A2(new_n1831_), .A3(new_n893_), .ZN(new_n2289_));
  NOR3_X1    g1923(.A1(new_n1844_), .A2(new_n2289_), .A3(\shift[4] ), .ZN(new_n2290_));
  NOR2_X1    g1924(.A1(new_n1842_), .A2(new_n1843_), .ZN(new_n2291_));
  NOR4_X1    g1925(.A1(new_n1832_), .A2(new_n1831_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2292_));
  NOR2_X1    g1926(.A1(new_n2290_), .A2(new_n2292_), .ZN(new_n2293_));
  OAI21_X1   g1927(.A1(new_n2288_), .A2(new_n2293_), .B(\shift[6] ), .ZN(new_n2294_));
  NAND2_X1   g1928(.A1(new_n2282_), .A2(new_n2294_), .ZN(\result[23] ));
  NOR2_X1    g1929(.A1(new_n1755_), .A2(new_n1893_), .ZN(new_n2296_));
  NOR3_X1    g1930(.A1(new_n1871_), .A2(new_n1870_), .A3(new_n893_), .ZN(new_n2297_));
  NOR3_X1    g1931(.A1(new_n2297_), .A2(new_n2296_), .A3(new_n1265_), .ZN(new_n2298_));
  NOR4_X1    g1932(.A1(new_n1871_), .A2(new_n1870_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2299_));
  NOR2_X1    g1933(.A1(new_n2298_), .A2(new_n2299_), .ZN(new_n2300_));
  NOR3_X1    g1934(.A1(new_n1860_), .A2(new_n1861_), .A3(new_n893_), .ZN(new_n2301_));
  OAI21_X1   g1935(.A1(new_n1873_), .A2(new_n1872_), .B(new_n984_), .ZN(new_n2302_));
  NOR2_X1    g1936(.A1(new_n2302_), .A2(new_n2301_), .ZN(new_n2303_));
  NOR4_X1    g1937(.A1(new_n1860_), .A2(new_n1861_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2305_));
  NOR2_X1    g1938(.A1(new_n2303_), .A2(new_n2305_), .ZN(new_n2306_));
  OAI21_X1   g1939(.A1(new_n2300_), .A2(new_n2306_), .B(new_n264_), .ZN(new_n2307_));
  NOR2_X1    g1940(.A1(new_n1753_), .A2(new_n1887_), .ZN(new_n2308_));
  INV_X1     g1941(.I(new_n2283_), .ZN(new_n2309_));
  NOR3_X1    g1942(.A1(new_n1883_), .A2(new_n1882_), .A3(new_n893_), .ZN(new_n2310_));
  NOR3_X1    g1943(.A1(new_n2310_), .A2(new_n2308_), .A3(new_n2309_), .ZN(new_n2311_));
  NOR4_X1    g1944(.A1(new_n1883_), .A2(new_n1882_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2312_));
  NOR2_X1    g1945(.A1(new_n2311_), .A2(new_n2312_), .ZN(new_n2313_));
  NOR3_X1    g1946(.A1(new_n1866_), .A2(new_n1724_), .A3(new_n893_), .ZN(new_n2314_));
  NOR3_X1    g1947(.A1(new_n1879_), .A2(new_n2314_), .A3(\shift[4] ), .ZN(new_n2315_));
  NOR2_X1    g1948(.A1(new_n1877_), .A2(new_n654_), .ZN(new_n2316_));
  NOR4_X1    g1949(.A1(new_n1866_), .A2(new_n1724_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2317_));
  NOR2_X1    g1950(.A1(new_n2315_), .A2(new_n2317_), .ZN(new_n2318_));
  OAI21_X1   g1951(.A1(new_n2318_), .A2(new_n2313_), .B(\shift[6] ), .ZN(new_n2319_));
  NAND2_X1   g1952(.A1(new_n2319_), .A2(new_n2307_), .ZN(\result[24] ));
  NOR3_X1    g1953(.A1(new_n1908_), .A2(new_n1909_), .A3(new_n893_), .ZN(new_n2321_));
  OAI21_X1   g1954(.A1(new_n1927_), .A2(new_n1928_), .B(new_n984_), .ZN(new_n2322_));
  XOR2_X1    g1955(.A1(new_n2322_), .A2(new_n2321_), .Z(new_n2323_));
  OAI21_X1   g1956(.A1(new_n1910_), .A2(new_n1911_), .B(new_n984_), .ZN(new_n2324_));
  AOI21_X1   g1957(.A1(new_n1901_), .A2(new_n987_), .B(new_n2324_), .ZN(new_n2325_));
  NOR4_X1    g1958(.A1(new_n1898_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1899_), .ZN(new_n2327_));
  NOR2_X1    g1959(.A1(new_n2325_), .A2(new_n2327_), .ZN(new_n2328_));
  OAI21_X1   g1960(.A1(new_n2323_), .A2(new_n2328_), .B(new_n264_), .ZN(new_n2329_));
  NOR4_X1    g1961(.A1(new_n1922_), .A2(new_n893_), .A3(new_n1920_), .A4(new_n1031_), .ZN(new_n2330_));
  OAI21_X1   g1962(.A1(new_n1789_), .A2(new_n1926_), .B(new_n2283_), .ZN(new_n2331_));
  XOR2_X1    g1963(.A1(new_n2330_), .A2(new_n2331_), .Z(new_n2332_));
  NOR3_X1    g1964(.A1(new_n1766_), .A2(new_n1904_), .A3(new_n893_), .ZN(new_n2333_));
  NOR4_X1    g1965(.A1(new_n2333_), .A2(new_n1917_), .A3(\shift[4] ), .A4(new_n266_), .ZN(new_n2334_));
  NOR4_X1    g1966(.A1(new_n1766_), .A2(new_n1904_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2335_));
  NOR2_X1    g1967(.A1(new_n2334_), .A2(new_n2335_), .ZN(new_n2336_));
  OAI21_X1   g1968(.A1(new_n2332_), .A2(new_n2336_), .B(\shift[6] ), .ZN(new_n2337_));
  NAND2_X1   g1969(.A1(new_n2329_), .A2(new_n2337_), .ZN(\result[25] ));
  NOR4_X1    g1970(.A1(new_n1951_), .A2(new_n1950_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2339_));
  NAND2_X1   g1971(.A1(new_n1230_), .A2(new_n1228_), .ZN(new_n2340_));
  NAND4_X1   g1972(.A1(new_n2340_), .A2(new_n276_), .A3(new_n1227_), .A4(new_n1232_), .ZN(new_n2341_));
  NOR4_X1    g1973(.A1(new_n2093_), .A2(new_n2257_), .A3(new_n2341_), .A4(new_n2259_), .ZN(new_n2342_));
  NOR3_X1    g1974(.A1(new_n2342_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2343_));
  NOR2_X1    g1975(.A1(new_n2343_), .A2(new_n2339_), .ZN(new_n2344_));
  NOR4_X1    g1976(.A1(new_n1965_), .A2(new_n1953_), .A3(new_n1966_), .A4(new_n1952_), .ZN(new_n2345_));
  OAI21_X1   g1977(.A1(new_n1944_), .A2(new_n1935_), .B(new_n2345_), .ZN(new_n2346_));
  OAI21_X1   g1978(.A1(new_n2344_), .A2(new_n2346_), .B(new_n264_), .ZN(new_n2347_));
  NOR2_X1    g1979(.A1(new_n1820_), .A2(new_n1964_), .ZN(new_n2348_));
  NOR3_X1    g1980(.A1(new_n1960_), .A2(new_n1815_), .A3(new_n893_), .ZN(new_n2349_));
  NOR3_X1    g1981(.A1(new_n2349_), .A2(new_n2348_), .A3(new_n2309_), .ZN(new_n2350_));
  NOR4_X1    g1982(.A1(new_n1960_), .A2(new_n1815_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2351_));
  NOR2_X1    g1983(.A1(new_n2350_), .A2(new_n2351_), .ZN(new_n2352_));
  NOR3_X1    g1984(.A1(new_n1801_), .A2(new_n1946_), .A3(new_n893_), .ZN(new_n2353_));
  NOR3_X1    g1985(.A1(new_n2353_), .A2(new_n1958_), .A3(\shift[4] ), .ZN(new_n2354_));
  NOR4_X1    g1986(.A1(new_n1801_), .A2(new_n1946_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2356_));
  NOR2_X1    g1987(.A1(new_n2354_), .A2(new_n2356_), .ZN(new_n2357_));
  OAI21_X1   g1988(.A1(new_n2357_), .A2(new_n2352_), .B(\shift[6] ), .ZN(new_n2358_));
  NAND2_X1   g1989(.A1(new_n2358_), .A2(new_n2347_), .ZN(\result[26] ));
  OAI21_X1   g1990(.A1(new_n1981_), .A2(new_n1837_), .B(\shift[5] ), .ZN(new_n2360_));
  XOR2_X1    g1991(.A1(new_n2360_), .A2(new_n987_), .Z(new_n2361_));
  NOR4_X1    g1992(.A1(new_n1855_), .A2(new_n1982_), .A3(new_n1983_), .A4(new_n1997_), .ZN(new_n2362_));
  OAI21_X1   g1993(.A1(new_n1975_), .A2(new_n1973_), .B(new_n2362_), .ZN(new_n2363_));
  OAI21_X1   g1994(.A1(new_n2363_), .A2(new_n2361_), .B(new_n264_), .ZN(new_n2364_));
  OAI21_X1   g1995(.A1(new_n1853_), .A2(new_n1996_), .B(new_n2283_), .ZN(new_n2365_));
  AOI21_X1   g1996(.A1(new_n987_), .A2(new_n1994_), .B(new_n2365_), .ZN(new_n2366_));
  NOR4_X1    g1997(.A1(new_n1990_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1991_), .ZN(new_n2368_));
  NOR2_X1    g1998(.A1(new_n2366_), .A2(new_n2368_), .ZN(new_n2369_));
  NOR3_X1    g1999(.A1(new_n1832_), .A2(new_n1977_), .A3(new_n893_), .ZN(new_n2370_));
  NOR3_X1    g2000(.A1(new_n2370_), .A2(new_n1988_), .A3(\shift[4] ), .ZN(new_n2371_));
  NOR4_X1    g2001(.A1(new_n1832_), .A2(new_n1977_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2373_));
  NOR2_X1    g2002(.A1(new_n2371_), .A2(new_n2373_), .ZN(new_n2374_));
  OAI21_X1   g2003(.A1(new_n2369_), .A2(new_n2374_), .B(\shift[6] ), .ZN(new_n2375_));
  NAND2_X1   g2004(.A1(new_n2364_), .A2(new_n2375_), .ZN(\result[27] ));
  NOR4_X1    g2005(.A1(new_n452_), .A2(new_n1728_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2377_));
  NAND2_X1   g2006(.A1(new_n416_), .A2(new_n410_), .ZN(new_n2378_));
  NAND2_X1   g2007(.A1(new_n436_), .A2(new_n434_), .ZN(new_n2379_));
  NAND4_X1   g2008(.A1(new_n433_), .A2(new_n276_), .A3(new_n2379_), .A4(new_n439_), .ZN(new_n2380_));
  NAND3_X1   g2009(.A1(new_n859_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n2381_));
  NAND2_X1   g2010(.A1(new_n2381_), .A2(new_n446_), .ZN(new_n2382_));
  NOR3_X1    g2011(.A1(new_n323_), .A2(new_n1231_), .A3(new_n858_), .ZN(new_n2383_));
  NAND3_X1   g2012(.A1(new_n445_), .A2(new_n2382_), .A3(new_n2383_), .ZN(new_n2384_));
  NAND3_X1   g2013(.A1(new_n883_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n2385_));
  NAND2_X1   g2014(.A1(new_n2385_), .A2(new_n466_), .ZN(new_n2386_));
  NAND4_X1   g2015(.A1(new_n465_), .A2(new_n2386_), .A3(new_n276_), .A4(new_n472_), .ZN(new_n2387_));
  NOR4_X1    g2016(.A1(new_n2378_), .A2(new_n2380_), .A3(new_n2384_), .A4(new_n2387_), .ZN(new_n2388_));
  NOR3_X1    g2017(.A1(new_n2388_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2389_));
  NOR2_X1    g2018(.A1(new_n2389_), .A2(new_n2377_), .ZN(new_n2390_));
  NOR4_X1    g2019(.A1(new_n291_), .A2(new_n619_), .A3(new_n2049_), .A4(new_n1729_), .ZN(new_n2391_));
  OAI21_X1   g2020(.A1(new_n2007_), .A2(new_n2002_), .B(new_n2391_), .ZN(new_n2392_));
  OAI21_X1   g2021(.A1(new_n2392_), .A2(new_n2390_), .B(new_n264_), .ZN(new_n2393_));
  NAND2_X1   g2022(.A1(new_n347_), .A2(new_n341_), .ZN(new_n2394_));
  NAND3_X1   g2023(.A1(new_n765_), .A2(new_n269_), .A3(\shift[0] ), .ZN(new_n2395_));
  NAND2_X1   g2024(.A1(new_n2395_), .A2(new_n352_), .ZN(new_n2396_));
  NAND4_X1   g2025(.A1(new_n351_), .A2(new_n276_), .A3(new_n2396_), .A4(new_n358_), .ZN(new_n2397_));
  NOR2_X1    g2026(.A1(new_n2394_), .A2(new_n2397_), .ZN(new_n2398_));
  NAND2_X1   g2027(.A1(new_n378_), .A2(new_n376_), .ZN(new_n2399_));
  NAND2_X1   g2028(.A1(\a[66] ), .A2(\a[68] ), .ZN(new_n2400_));
  NOR2_X1    g2029(.A1(new_n323_), .A2(new_n2400_), .ZN(new_n2401_));
  NAND3_X1   g2030(.A1(new_n375_), .A2(new_n2399_), .A3(new_n2401_), .ZN(new_n2402_));
  NOR2_X1    g2031(.A1(new_n2402_), .A2(new_n536_), .ZN(new_n2403_));
  NAND2_X1   g2032(.A1(new_n2398_), .A2(new_n2403_), .ZN(new_n2404_));
  NOR2_X1    g2033(.A1(new_n526_), .A2(new_n1744_), .ZN(new_n2405_));
  NOR2_X1    g2034(.A1(new_n529_), .A2(new_n542_), .ZN(new_n2406_));
  NAND3_X1   g2035(.A1(new_n2405_), .A2(new_n2406_), .A3(new_n987_), .ZN(new_n2407_));
  NAND3_X1   g2036(.A1(new_n2407_), .A2(new_n2404_), .A3(new_n2283_), .ZN(new_n2408_));
  NAND3_X1   g2037(.A1(new_n2046_), .A2(\shift[4] ), .A3(\shift[5] ), .ZN(new_n2410_));
  NOR2_X1    g2038(.A1(new_n2040_), .A2(new_n266_), .ZN(new_n2411_));
  NAND2_X1   g2039(.A1(new_n2022_), .A2(new_n987_), .ZN(new_n2412_));
  NAND3_X1   g2040(.A1(new_n2412_), .A2(new_n2411_), .A3(new_n265_), .ZN(new_n2413_));
  NAND3_X1   g2041(.A1(new_n2022_), .A2(\shift[4] ), .A3(\shift[5] ), .ZN(new_n2414_));
  AOI22_X1   g2042(.A1(new_n2413_), .A2(new_n2414_), .B1(new_n2408_), .B2(new_n2410_), .ZN(new_n2415_));
  OAI21_X1   g2043(.A1(new_n264_), .A2(new_n2415_), .B(new_n2393_), .ZN(\result[28] ));
  OAI21_X1   g2044(.A1(new_n865_), .A2(new_n1770_), .B(\shift[5] ), .ZN(new_n2417_));
  XOR2_X1    g2045(.A1(new_n2417_), .A2(new_n987_), .Z(new_n2418_));
  NOR4_X1    g2046(.A1(new_n719_), .A2(new_n1058_), .A3(new_n1771_), .A4(new_n1790_), .ZN(new_n2419_));
  OAI21_X1   g2047(.A1(new_n2056_), .A2(new_n2054_), .B(new_n2419_), .ZN(new_n2420_));
  NOR2_X1    g2048(.A1(new_n2420_), .A2(new_n2418_), .ZN(new_n2421_));
  NOR2_X1    g2049(.A1(new_n771_), .A2(new_n2074_), .ZN(new_n2422_));
  NOR3_X1    g2050(.A1(new_n916_), .A2(new_n1922_), .A3(new_n893_), .ZN(new_n2423_));
  NOR3_X1    g2051(.A1(new_n2423_), .A2(new_n2422_), .A3(new_n2309_), .ZN(new_n2424_));
  NOR4_X1    g2052(.A1(new_n916_), .A2(new_n1922_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2425_));
  NOR2_X1    g2053(.A1(new_n2424_), .A2(new_n2425_), .ZN(new_n2426_));
  NOR3_X1    g2054(.A1(new_n820_), .A2(new_n2058_), .A3(new_n893_), .ZN(new_n2427_));
  NOR4_X1    g2055(.A1(new_n2427_), .A2(new_n2066_), .A3(\shift[4] ), .A4(new_n266_), .ZN(new_n2428_));
  NOR4_X1    g2056(.A1(new_n820_), .A2(new_n2058_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2429_));
  NOR2_X1    g2057(.A1(new_n2428_), .A2(new_n2429_), .ZN(new_n2430_));
  OAI21_X1   g2058(.A1(new_n2430_), .A2(new_n2426_), .B(\shift[6] ), .ZN(new_n2431_));
  OAI21_X1   g2059(.A1(new_n2421_), .A2(\shift[6] ), .B(new_n2431_), .ZN(\result[29] ));
  NOR4_X1    g2060(.A1(new_n1805_), .A2(new_n1243_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2433_));
  NOR2_X1    g2061(.A1(new_n1805_), .A2(new_n1243_), .ZN(new_n2434_));
  NOR3_X1    g2062(.A1(new_n2434_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2435_));
  NOR2_X1    g2063(.A1(new_n2435_), .A2(new_n2433_), .ZN(new_n2436_));
  NOR4_X1    g2064(.A1(new_n1108_), .A2(new_n1821_), .A3(new_n1397_), .A4(new_n1806_), .ZN(new_n2437_));
  OAI21_X1   g2065(.A1(new_n2084_), .A2(new_n2079_), .B(new_n2437_), .ZN(new_n2438_));
  OAI21_X1   g2066(.A1(new_n2436_), .A2(new_n2438_), .B(new_n264_), .ZN(new_n2439_));
  NOR2_X1    g2067(.A1(new_n1160_), .A2(new_n2120_), .ZN(new_n2440_));
  NOR3_X1    g2068(.A1(new_n1284_), .A2(new_n2107_), .A3(new_n893_), .ZN(new_n2441_));
  NOR3_X1    g2069(.A1(new_n2441_), .A2(new_n2440_), .A3(new_n2309_), .ZN(new_n2442_));
  NOR4_X1    g2070(.A1(new_n1284_), .A2(new_n2107_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2443_));
  NOR2_X1    g2071(.A1(new_n2442_), .A2(new_n2443_), .ZN(new_n2444_));
  NOR3_X1    g2072(.A1(new_n1203_), .A2(new_n2086_), .A3(new_n893_), .ZN(new_n2445_));
  NOR4_X1    g2073(.A1(new_n2445_), .A2(new_n2104_), .A3(\shift[4] ), .A4(new_n266_), .ZN(new_n2446_));
  NOR4_X1    g2074(.A1(new_n1203_), .A2(new_n2086_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2447_));
  NOR2_X1    g2075(.A1(new_n2446_), .A2(new_n2447_), .ZN(new_n2448_));
  OAI21_X1   g2076(.A1(new_n2448_), .A2(new_n2444_), .B(\shift[6] ), .ZN(new_n2449_));
  NAND2_X1   g2077(.A1(new_n2449_), .A2(new_n2439_), .ZN(\result[30] ));
  OAI21_X1   g2078(.A1(new_n1437_), .A2(new_n2133_), .B(\shift[5] ), .ZN(new_n2451_));
  XOR2_X1    g2079(.A1(new_n2451_), .A2(new_n987_), .Z(new_n2452_));
  NOR4_X1    g2080(.A1(new_n1509_), .A2(new_n1690_), .A3(new_n1838_), .A4(new_n2146_), .ZN(new_n2453_));
  OAI21_X1   g2081(.A1(new_n2127_), .A2(new_n2125_), .B(new_n2453_), .ZN(new_n2454_));
  OAI21_X1   g2082(.A1(new_n2452_), .A2(new_n2454_), .B(new_n264_), .ZN(new_n2455_));
  NOR3_X1    g2083(.A1(new_n1617_), .A2(new_n1846_), .A3(new_n893_), .ZN(new_n2456_));
  OAI21_X1   g2084(.A1(new_n1542_), .A2(new_n2145_), .B(new_n2283_), .ZN(new_n2457_));
  XOR2_X1    g2085(.A1(new_n2457_), .A2(new_n2456_), .Z(new_n2458_));
  NOR3_X1    g2086(.A1(new_n1469_), .A2(new_n2129_), .A3(new_n893_), .ZN(new_n2459_));
  NOR4_X1    g2087(.A1(new_n2459_), .A2(\shift[4] ), .A3(new_n2139_), .A4(new_n266_), .ZN(new_n2460_));
  NOR4_X1    g2088(.A1(new_n1469_), .A2(new_n2129_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2461_));
  NOR2_X1    g2089(.A1(new_n2460_), .A2(new_n2461_), .ZN(new_n2462_));
  OAI21_X1   g2090(.A1(new_n2458_), .A2(new_n2462_), .B(\shift[6] ), .ZN(new_n2463_));
  NAND2_X1   g2091(.A1(new_n2463_), .A2(new_n2455_), .ZN(\result[31] ));
  NOR4_X1    g2092(.A1(new_n571_), .A2(new_n594_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2465_));
  NOR3_X1    g2093(.A1(new_n596_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2466_));
  NOR2_X1    g2094(.A1(new_n2466_), .A2(new_n2465_), .ZN(new_n2467_));
  NOR4_X1    g2095(.A1(new_n291_), .A2(new_n316_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2468_));
  NOR3_X1    g2096(.A1(new_n335_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2469_));
  NOR4_X1    g2097(.A1(new_n641_), .A2(new_n452_), .A3(new_n619_), .A4(new_n475_), .ZN(new_n2470_));
  OAI21_X1   g2098(.A1(new_n2469_), .A2(new_n2468_), .B(new_n2470_), .ZN(new_n2471_));
  OAI21_X1   g2099(.A1(new_n2467_), .A2(new_n2471_), .B(new_n264_), .ZN(new_n2472_));
  NOR4_X1    g2100(.A1(new_n498_), .A2(new_n522_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2473_));
  NOR3_X1    g2101(.A1(new_n543_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2474_));
  NOR2_X1    g2102(.A1(new_n2474_), .A2(new_n2473_), .ZN(new_n2475_));
  NOR4_X1    g2103(.A1(new_n381_), .A2(new_n361_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2476_));
  NOR3_X1    g2104(.A1(new_n383_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2477_));
  NOR4_X1    g2105(.A1(new_n694_), .A2(new_n406_), .A3(new_n429_), .A4(new_n654_), .ZN(new_n2478_));
  OAI21_X1   g2106(.A1(new_n2477_), .A2(new_n2476_), .B(new_n2478_), .ZN(new_n2479_));
  OAI21_X1   g2107(.A1(new_n2479_), .A2(new_n2475_), .B(\shift[6] ), .ZN(new_n2480_));
  NAND2_X1   g2108(.A1(new_n2480_), .A2(new_n2472_), .ZN(\result[32] ));
  OAI21_X1   g2109(.A1(new_n960_), .A2(new_n983_), .B(\shift[4] ), .ZN(new_n2482_));
  XOR2_X1    g2110(.A1(new_n2482_), .A2(new_n987_), .Z(new_n2483_));
  NOR4_X1    g2111(.A1(new_n744_), .A2(new_n265_), .A3(new_n266_), .A4(new_n719_), .ZN(new_n2484_));
  NOR3_X1    g2112(.A1(new_n746_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2485_));
  NOR4_X1    g2113(.A1(new_n865_), .A2(new_n889_), .A3(new_n1058_), .A4(new_n1083_), .ZN(new_n2486_));
  OAI21_X1   g2114(.A1(new_n2485_), .A2(new_n2484_), .B(new_n2486_), .ZN(new_n2487_));
  OAI21_X1   g2115(.A1(new_n2487_), .A2(new_n2483_), .B(new_n264_), .ZN(new_n2488_));
  NOR3_X1    g2116(.A1(new_n771_), .A2(new_n795_), .A3(new_n893_), .ZN(new_n2489_));
  OAI21_X1   g2117(.A1(new_n916_), .A2(new_n937_), .B(new_n984_), .ZN(new_n2490_));
  XOR2_X1    g2118(.A1(new_n2490_), .A2(new_n2489_), .Z(new_n2491_));
  NOR3_X1    g2119(.A1(new_n820_), .A2(new_n842_), .A3(new_n893_), .ZN(new_n2492_));
  NOR4_X1    g2120(.A1(new_n2492_), .A2(new_n1032_), .A3(\shift[4] ), .A4(new_n266_), .ZN(new_n2493_));
  NOR4_X1    g2121(.A1(new_n820_), .A2(new_n842_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2494_));
  NOR2_X1    g2122(.A1(new_n2493_), .A2(new_n2494_), .ZN(new_n2495_));
  OAI21_X1   g2123(.A1(new_n2491_), .A2(new_n2495_), .B(\shift[6] ), .ZN(new_n2496_));
  NAND2_X1   g2124(.A1(new_n2488_), .A2(new_n2496_), .ZN(\result[33] ));
  NOR4_X1    g2125(.A1(new_n1321_), .A2(new_n1339_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2498_));
  NOR3_X1    g2126(.A1(new_n1340_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2499_));
  NOR2_X1    g2127(.A1(new_n2499_), .A2(new_n2498_), .ZN(new_n2500_));
  NOR4_X1    g2128(.A1(new_n1108_), .A2(new_n1129_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2501_));
  NOR3_X1    g2129(.A1(new_n1140_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2502_));
  NOR4_X1    g2130(.A1(new_n1243_), .A2(new_n1261_), .A3(new_n1397_), .A4(new_n1414_), .ZN(new_n2503_));
  OAI21_X1   g2131(.A1(new_n2502_), .A2(new_n2501_), .B(new_n2503_), .ZN(new_n2504_));
  OAI21_X1   g2132(.A1(new_n2500_), .A2(new_n2504_), .B(new_n264_), .ZN(new_n2505_));
  NOR2_X1    g2133(.A1(new_n1284_), .A2(new_n1303_), .ZN(new_n2506_));
  NOR3_X1    g2134(.A1(new_n1160_), .A2(new_n1182_), .A3(new_n893_), .ZN(new_n2507_));
  NOR3_X1    g2135(.A1(new_n2507_), .A2(new_n2506_), .A3(new_n1265_), .ZN(new_n2508_));
  NOR4_X1    g2136(.A1(new_n1160_), .A2(new_n1182_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2509_));
  NOR2_X1    g2137(.A1(new_n2508_), .A2(new_n2509_), .ZN(new_n2510_));
  NOR3_X1    g2138(.A1(new_n1203_), .A2(new_n1224_), .A3(new_n893_), .ZN(new_n2511_));
  NOR4_X1    g2139(.A1(new_n2511_), .A2(new_n2200_), .A3(\shift[4] ), .A4(new_n266_), .ZN(new_n2512_));
  NOR4_X1    g2140(.A1(new_n1203_), .A2(new_n1224_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2513_));
  NOR2_X1    g2141(.A1(new_n2512_), .A2(new_n2513_), .ZN(new_n2514_));
  OAI21_X1   g2142(.A1(new_n2514_), .A2(new_n2510_), .B(\shift[6] ), .ZN(new_n2515_));
  NAND2_X1   g2143(.A1(new_n2515_), .A2(new_n2505_), .ZN(\result[34] ));
  OAI21_X1   g2144(.A1(new_n1690_), .A2(new_n1709_), .B(new_n984_), .ZN(new_n2517_));
  XOR2_X1    g2145(.A1(new_n1454_), .A2(new_n2517_), .Z(new_n2518_));
  NOR2_X1    g2146(.A1(new_n1581_), .A2(new_n1599_), .ZN(new_n2519_));
  NOR3_X1    g2147(.A1(new_n1526_), .A2(new_n2519_), .A3(new_n2309_), .ZN(new_n2520_));
  NOR4_X1    g2148(.A1(new_n1509_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1525_), .ZN(new_n2521_));
  NOR2_X1    g2149(.A1(new_n2520_), .A2(new_n2521_), .ZN(new_n2522_));
  OAI21_X1   g2150(.A1(new_n2522_), .A2(new_n2518_), .B(new_n264_), .ZN(new_n2523_));
  XOR2_X1    g2151(.A1(new_n1489_), .A2(new_n987_), .Z(new_n2524_));
  NOR4_X1    g2152(.A1(new_n1654_), .A2(new_n1617_), .A3(new_n1633_), .A4(new_n1673_), .ZN(new_n2525_));
  OAI21_X1   g2153(.A1(new_n2224_), .A2(new_n2223_), .B(new_n2525_), .ZN(new_n2526_));
  OAI21_X1   g2154(.A1(new_n2524_), .A2(new_n2526_), .B(\shift[6] ), .ZN(new_n2527_));
  NAND2_X1   g2155(.A1(new_n2523_), .A2(new_n2527_), .ZN(\result[35] ));
  NOR4_X1    g2156(.A1(new_n1748_), .A2(new_n619_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2529_));
  NOR3_X1    g2157(.A1(new_n1750_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2530_));
  NOR2_X1    g2158(.A1(new_n2530_), .A2(new_n2529_), .ZN(new_n2531_));
  NOR2_X1    g2159(.A1(new_n319_), .A2(new_n325_), .ZN(new_n2532_));
  NOR2_X1    g2160(.A1(new_n329_), .A2(new_n1719_), .ZN(new_n2533_));
  NAND2_X1   g2161(.A1(new_n2532_), .A2(new_n2533_), .ZN(new_n2534_));
  AOI21_X1   g2162(.A1(new_n2534_), .A2(\shift[5] ), .B(new_n893_), .ZN(new_n2535_));
  NOR3_X1    g2163(.A1(new_n1720_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2536_));
  OAI21_X1   g2164(.A1(new_n2535_), .A2(new_n2536_), .B(new_n2233_), .ZN(new_n2537_));
  OAI21_X1   g2165(.A1(new_n2537_), .A2(new_n2531_), .B(new_n264_), .ZN(new_n2538_));
  NOR4_X1    g2166(.A1(new_n1733_), .A2(new_n265_), .A3(new_n266_), .A4(new_n654_), .ZN(new_n2539_));
  NOR3_X1    g2167(.A1(new_n1745_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2540_));
  NOR2_X1    g2168(.A1(new_n2540_), .A2(new_n2539_), .ZN(new_n2541_));
  NOR4_X1    g2169(.A1(new_n1723_), .A2(new_n1724_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2542_));
  NOR3_X1    g2170(.A1(new_n1726_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2543_));
  NOR4_X1    g2171(.A1(new_n406_), .A2(new_n1752_), .A3(new_n1753_), .A4(new_n1728_), .ZN(new_n2544_));
  OAI21_X1   g2172(.A1(new_n2543_), .A2(new_n2542_), .B(new_n2544_), .ZN(new_n2545_));
  OAI21_X1   g2173(.A1(new_n2545_), .A2(new_n2541_), .B(\shift[6] ), .ZN(new_n2546_));
  NAND2_X1   g2174(.A1(new_n2538_), .A2(new_n2546_), .ZN(\result[36] ));
  NOR4_X1    g2175(.A1(new_n1777_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1778_), .ZN(new_n2548_));
  NOR3_X1    g2176(.A1(new_n1780_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2549_));
  NOR2_X1    g2177(.A1(new_n2549_), .A2(new_n2548_), .ZN(new_n2550_));
  NOR4_X1    g2178(.A1(new_n1760_), .A2(new_n265_), .A3(new_n266_), .A4(new_n719_), .ZN(new_n2551_));
  NOR3_X1    g2179(.A1(new_n1762_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2552_));
  OAI21_X1   g2180(.A1(new_n2552_), .A2(new_n2551_), .B(new_n2246_), .ZN(new_n2553_));
  OAI21_X1   g2181(.A1(new_n2550_), .A2(new_n2553_), .B(new_n264_), .ZN(new_n2554_));
  NOR2_X1    g2182(.A1(new_n1786_), .A2(new_n266_), .ZN(new_n2555_));
  NOR2_X1    g2183(.A1(new_n2555_), .A2(new_n893_), .ZN(new_n2556_));
  NOR3_X1    g2184(.A1(new_n1786_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2557_));
  NOR2_X1    g2185(.A1(new_n2556_), .A2(new_n2557_), .ZN(new_n2558_));
  NOR4_X1    g2186(.A1(new_n1765_), .A2(new_n1766_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2559_));
  NOR3_X1    g2187(.A1(new_n1768_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2560_));
  NOR4_X1    g2188(.A1(new_n820_), .A2(new_n1770_), .A3(new_n1788_), .A4(new_n1789_), .ZN(new_n2561_));
  OAI21_X1   g2189(.A1(new_n2560_), .A2(new_n2559_), .B(new_n2561_), .ZN(new_n2562_));
  OAI21_X1   g2190(.A1(new_n2558_), .A2(new_n2562_), .B(\shift[6] ), .ZN(new_n2563_));
  NAND2_X1   g2191(.A1(new_n2554_), .A2(new_n2563_), .ZN(\result[37] ));
  OAI21_X1   g2192(.A1(new_n1810_), .A2(new_n1811_), .B(\shift[4] ), .ZN(new_n2565_));
  XOR2_X1    g2193(.A1(new_n2565_), .A2(new_n987_), .Z(new_n2566_));
  NOR4_X1    g2194(.A1(new_n1108_), .A2(new_n1795_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2567_));
  NOR3_X1    g2195(.A1(new_n1797_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2568_));
  OAI21_X1   g2196(.A1(new_n2568_), .A2(new_n2567_), .B(new_n2263_), .ZN(new_n2569_));
  OAI21_X1   g2197(.A1(new_n2566_), .A2(new_n2569_), .B(new_n264_), .ZN(new_n2570_));
  NOR4_X1    g2198(.A1(new_n1814_), .A2(new_n1815_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2571_));
  OAI21_X1   g2199(.A1(new_n1814_), .A2(new_n1815_), .B(\shift[5] ), .ZN(new_n2572_));
  NOR2_X1    g2200(.A1(new_n2572_), .A2(new_n987_), .ZN(new_n2573_));
  NOR2_X1    g2201(.A1(new_n2573_), .A2(new_n2571_), .ZN(new_n2574_));
  NOR4_X1    g2202(.A1(new_n1800_), .A2(new_n1801_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2575_));
  NOR3_X1    g2203(.A1(new_n1803_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2576_));
  NOR4_X1    g2204(.A1(new_n1203_), .A2(new_n1805_), .A3(new_n1820_), .A4(new_n1819_), .ZN(new_n2577_));
  OAI21_X1   g2205(.A1(new_n2576_), .A2(new_n2575_), .B(new_n2577_), .ZN(new_n2578_));
  OAI21_X1   g2206(.A1(new_n2578_), .A2(new_n2574_), .B(\shift[6] ), .ZN(new_n2579_));
  NAND2_X1   g2207(.A1(new_n2570_), .A2(new_n2579_), .ZN(\result[38] ));
  NOR4_X1    g2208(.A1(new_n1509_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1826_), .ZN(new_n2581_));
  NOR3_X1    g2209(.A1(new_n1828_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2582_));
  NOR2_X1    g2210(.A1(new_n2582_), .A2(new_n2581_), .ZN(new_n2583_));
  NOR4_X1    g2211(.A1(new_n1842_), .A2(new_n1843_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2584_));
  NOR3_X1    g2212(.A1(new_n2291_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2585_));
  NOR4_X1    g2213(.A1(new_n1437_), .A2(new_n1838_), .A3(new_n1854_), .A4(new_n1855_), .ZN(new_n2586_));
  OAI21_X1   g2214(.A1(new_n2585_), .A2(new_n2584_), .B(new_n2586_), .ZN(new_n2587_));
  OAI21_X1   g2215(.A1(new_n2583_), .A2(new_n2587_), .B(new_n264_), .ZN(new_n2588_));
  OAI21_X1   g2216(.A1(new_n1832_), .A2(new_n1831_), .B(\shift[4] ), .ZN(new_n2589_));
  XOR2_X1    g2217(.A1(new_n2589_), .A2(new_n987_), .Z(new_n2590_));
  NOR4_X1    g2218(.A1(new_n1654_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1846_), .ZN(new_n2591_));
  NOR3_X1    g2219(.A1(new_n1850_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2592_));
  NOR4_X1    g2220(.A1(new_n1836_), .A2(new_n1853_), .A3(new_n1837_), .A4(new_n1852_), .ZN(new_n2593_));
  OAI21_X1   g2221(.A1(new_n2592_), .A2(new_n2591_), .B(new_n2593_), .ZN(new_n2594_));
  OAI21_X1   g2222(.A1(new_n2590_), .A2(new_n2594_), .B(\shift[6] ), .ZN(new_n2595_));
  NAND2_X1   g2223(.A1(new_n2595_), .A2(new_n2588_), .ZN(\result[39] ));
  NOR4_X1    g2224(.A1(new_n1877_), .A2(new_n265_), .A3(new_n266_), .A4(new_n654_), .ZN(new_n2597_));
  NOR3_X1    g2225(.A1(new_n2316_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2598_));
  NOR2_X1    g2226(.A1(new_n2598_), .A2(new_n2597_), .ZN(new_n2599_));
  NOR4_X1    g2227(.A1(new_n1860_), .A2(new_n1861_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2600_));
  NOR3_X1    g2228(.A1(new_n1863_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2601_));
  NOR4_X1    g2229(.A1(new_n1755_), .A2(new_n1873_), .A3(new_n1893_), .A4(new_n1872_), .ZN(new_n2602_));
  OAI21_X1   g2230(.A1(new_n2601_), .A2(new_n2600_), .B(new_n2602_), .ZN(new_n2603_));
  OAI21_X1   g2231(.A1(new_n2599_), .A2(new_n2603_), .B(new_n264_), .ZN(new_n2604_));
  NOR4_X1    g2232(.A1(new_n1866_), .A2(new_n1724_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2605_));
  NOR3_X1    g2233(.A1(new_n1868_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2606_));
  NOR2_X1    g2234(.A1(new_n2606_), .A2(new_n2605_), .ZN(new_n2607_));
  NOR4_X1    g2235(.A1(new_n1883_), .A2(new_n1882_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2608_));
  NOR3_X1    g2236(.A1(new_n1885_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2609_));
  NOR4_X1    g2237(.A1(new_n1753_), .A2(new_n1870_), .A3(new_n1871_), .A4(new_n1887_), .ZN(new_n2610_));
  OAI21_X1   g2238(.A1(new_n2609_), .A2(new_n2608_), .B(new_n2610_), .ZN(new_n2611_));
  OAI21_X1   g2239(.A1(new_n2607_), .A2(new_n2611_), .B(\shift[6] ), .ZN(new_n2612_));
  NAND2_X1   g2240(.A1(new_n2604_), .A2(new_n2612_), .ZN(\result[40] ));
  NOR4_X1    g2241(.A1(new_n1898_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1899_), .ZN(new_n2614_));
  NOR3_X1    g2242(.A1(new_n1901_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2615_));
  NOR2_X1    g2243(.A1(new_n2615_), .A2(new_n2614_), .ZN(new_n2616_));
  NOR4_X1    g2244(.A1(new_n1915_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1778_), .ZN(new_n2617_));
  NOR3_X1    g2245(.A1(new_n1917_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2618_));
  NOR4_X1    g2246(.A1(new_n1910_), .A2(new_n1911_), .A3(new_n1927_), .A4(new_n1928_), .ZN(new_n2619_));
  OAI21_X1   g2247(.A1(new_n2617_), .A2(new_n2618_), .B(new_n2619_), .ZN(new_n2620_));
  OAI21_X1   g2248(.A1(new_n2620_), .A2(new_n2616_), .B(new_n264_), .ZN(new_n2621_));
  OAI21_X1   g2249(.A1(new_n1766_), .A2(new_n1904_), .B(\shift[4] ), .ZN(new_n2622_));
  XOR2_X1    g2250(.A1(new_n2622_), .A2(new_n987_), .Z(new_n2623_));
  NOR4_X1    g2251(.A1(new_n1921_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1922_), .ZN(new_n2624_));
  NOR3_X1    g2252(.A1(new_n1924_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2625_));
  NOR4_X1    g2253(.A1(new_n1789_), .A2(new_n1908_), .A3(new_n1909_), .A4(new_n1926_), .ZN(new_n2626_));
  OAI21_X1   g2254(.A1(new_n2624_), .A2(new_n2625_), .B(new_n2626_), .ZN(new_n2627_));
  OAI21_X1   g2255(.A1(new_n2623_), .A2(new_n2627_), .B(\shift[6] ), .ZN(new_n2628_));
  NAND2_X1   g2256(.A1(new_n2621_), .A2(new_n2628_), .ZN(\result[41] ));
  OAI21_X1   g2257(.A1(new_n1957_), .A2(new_n1811_), .B(\shift[4] ), .ZN(new_n2630_));
  XOR2_X1    g2258(.A1(new_n2630_), .A2(new_n987_), .Z(new_n2631_));
  NOR4_X1    g2259(.A1(new_n1934_), .A2(new_n1933_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2632_));
  NOR3_X1    g2260(.A1(new_n1943_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2633_));
  OAI21_X1   g2261(.A1(new_n2633_), .A2(new_n2632_), .B(new_n2345_), .ZN(new_n2634_));
  OAI21_X1   g2262(.A1(new_n2631_), .A2(new_n2634_), .B(new_n264_), .ZN(new_n2635_));
  NOR4_X1    g2263(.A1(new_n1801_), .A2(new_n1946_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2636_));
  NOR3_X1    g2264(.A1(new_n1948_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2637_));
  NOR2_X1    g2265(.A1(new_n2637_), .A2(new_n2636_), .ZN(new_n2638_));
  NOR4_X1    g2266(.A1(new_n1960_), .A2(new_n1815_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2639_));
  OAI21_X1   g2267(.A1(new_n1960_), .A2(new_n1815_), .B(\shift[5] ), .ZN(new_n2640_));
  NOR2_X1    g2268(.A1(new_n2640_), .A2(new_n987_), .ZN(new_n2641_));
  NOR4_X1    g2269(.A1(new_n1820_), .A2(new_n1950_), .A3(new_n1951_), .A4(new_n1964_), .ZN(new_n2642_));
  OAI21_X1   g2270(.A1(new_n2641_), .A2(new_n2639_), .B(new_n2642_), .ZN(new_n2643_));
  OAI21_X1   g2271(.A1(new_n2643_), .A2(new_n2638_), .B(\shift[6] ), .ZN(new_n2644_));
  NAND2_X1   g2272(.A1(new_n2635_), .A2(new_n2644_), .ZN(\result[42] ));
  OAI21_X1   g2273(.A1(new_n1843_), .A2(new_n1987_), .B(\shift[4] ), .ZN(new_n2646_));
  XOR2_X1    g2274(.A1(new_n2646_), .A2(new_n987_), .Z(new_n2647_));
  NOR4_X1    g2275(.A1(new_n1971_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1972_), .ZN(new_n2648_));
  NOR3_X1    g2276(.A1(new_n1974_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2649_));
  OAI21_X1   g2277(.A1(new_n2649_), .A2(new_n2648_), .B(new_n2362_), .ZN(new_n2650_));
  OAI21_X1   g2278(.A1(new_n2650_), .A2(new_n2647_), .B(new_n264_), .ZN(new_n2651_));
  OAI21_X1   g2279(.A1(new_n1832_), .A2(new_n1977_), .B(\shift[4] ), .ZN(new_n2652_));
  XOR2_X1    g2280(.A1(new_n2652_), .A2(new_n987_), .Z(new_n2653_));
  NOR4_X1    g2281(.A1(new_n1990_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1991_), .ZN(new_n2654_));
  NOR3_X1    g2282(.A1(new_n1994_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2655_));
  NOR4_X1    g2283(.A1(new_n1853_), .A2(new_n1981_), .A3(new_n1837_), .A4(new_n1996_), .ZN(new_n2656_));
  OAI21_X1   g2284(.A1(new_n2655_), .A2(new_n2654_), .B(new_n2656_), .ZN(new_n2657_));
  OAI21_X1   g2285(.A1(new_n2653_), .A2(new_n2657_), .B(\shift[6] ), .ZN(new_n2658_));
  NAND2_X1   g2286(.A1(new_n2651_), .A2(new_n2658_), .ZN(\result[43] ));
  NOR4_X1    g2287(.A1(new_n2027_), .A2(new_n265_), .A3(new_n266_), .A4(new_n654_), .ZN(new_n2660_));
  NOR3_X1    g2288(.A1(new_n2040_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2661_));
  NOR2_X1    g2289(.A1(new_n2661_), .A2(new_n2660_), .ZN(new_n2662_));
  NOR4_X1    g2290(.A1(new_n571_), .A2(new_n1714_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2663_));
  NOR3_X1    g2291(.A1(new_n2006_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2664_));
  OAI21_X1   g2292(.A1(new_n2664_), .A2(new_n2663_), .B(new_n2391_), .ZN(new_n2665_));
  OAI21_X1   g2293(.A1(new_n2665_), .A2(new_n2662_), .B(new_n264_), .ZN(new_n2666_));
  NOR4_X1    g2294(.A1(new_n406_), .A2(new_n2009_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2667_));
  NOR3_X1    g2295(.A1(new_n2022_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2668_));
  NOR2_X1    g2296(.A1(new_n2668_), .A2(new_n2667_), .ZN(new_n2669_));
  NOR4_X1    g2297(.A1(new_n2044_), .A2(new_n2043_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2670_));
  NOR3_X1    g2298(.A1(new_n2046_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2671_));
  NOR4_X1    g2299(.A1(new_n361_), .A2(new_n452_), .A3(new_n2048_), .A4(new_n1728_), .ZN(new_n2672_));
  OAI21_X1   g2300(.A1(new_n2671_), .A2(new_n2670_), .B(new_n2672_), .ZN(new_n2673_));
  OAI21_X1   g2301(.A1(new_n2673_), .A2(new_n2669_), .B(\shift[6] ), .ZN(new_n2674_));
  NAND2_X1   g2302(.A1(new_n2666_), .A2(new_n2674_), .ZN(\result[44] ));
  AND3_X2    g2303(.A1(new_n2066_), .A2(\shift[4] ), .A3(\shift[5] ), .Z(new_n2676_));
  NOR3_X1    g2304(.A1(new_n2066_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2677_));
  NOR2_X1    g2305(.A1(new_n2676_), .A2(new_n2677_), .ZN(new_n2678_));
  NOR4_X1    g2306(.A1(new_n1760_), .A2(new_n265_), .A3(new_n266_), .A4(new_n960_), .ZN(new_n2679_));
  NOR3_X1    g2307(.A1(new_n2055_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2680_));
  OAI21_X1   g2308(.A1(new_n2680_), .A2(new_n2679_), .B(new_n2419_), .ZN(new_n2681_));
  OAI21_X1   g2309(.A1(new_n2681_), .A2(new_n2678_), .B(new_n264_), .ZN(new_n2682_));
  OAI21_X1   g2310(.A1(new_n820_), .A2(new_n2058_), .B(\shift[4] ), .ZN(new_n2683_));
  XOR2_X1    g2311(.A1(new_n2683_), .A2(new_n987_), .Z(new_n2684_));
  NOR4_X1    g2312(.A1(new_n916_), .A2(new_n1922_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2685_));
  OAI21_X1   g2313(.A1(new_n916_), .A2(new_n1922_), .B(\shift[5] ), .ZN(new_n2686_));
  NOR2_X1    g2314(.A1(new_n2686_), .A2(new_n987_), .ZN(new_n2687_));
  NOR4_X1    g2315(.A1(new_n771_), .A2(new_n865_), .A3(new_n1770_), .A4(new_n2074_), .ZN(new_n2688_));
  OAI21_X1   g2316(.A1(new_n2687_), .A2(new_n2685_), .B(new_n2688_), .ZN(new_n2689_));
  OAI21_X1   g2317(.A1(new_n2684_), .A2(new_n2689_), .B(\shift[6] ), .ZN(new_n2690_));
  NAND2_X1   g2318(.A1(new_n2682_), .A2(new_n2690_), .ZN(\result[45] ));
  NOR4_X1    g2319(.A1(new_n1360_), .A2(new_n2102_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2692_));
  NOR3_X1    g2320(.A1(new_n2104_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2693_));
  NOR2_X1    g2321(.A1(new_n2693_), .A2(new_n2692_), .ZN(new_n2694_));
  NOR4_X1    g2322(.A1(new_n1321_), .A2(new_n1795_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2695_));
  NOR3_X1    g2323(.A1(new_n2083_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2696_));
  OAI21_X1   g2324(.A1(new_n2696_), .A2(new_n2695_), .B(new_n2437_), .ZN(new_n2697_));
  OAI21_X1   g2325(.A1(new_n2694_), .A2(new_n2697_), .B(new_n264_), .ZN(new_n2698_));
  NOR4_X1    g2326(.A1(new_n1203_), .A2(new_n2086_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2699_));
  NOR3_X1    g2327(.A1(new_n2097_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2700_));
  NOR2_X1    g2328(.A1(new_n2700_), .A2(new_n2699_), .ZN(new_n2701_));
  NOR4_X1    g2329(.A1(new_n1284_), .A2(new_n2107_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2702_));
  NOR3_X1    g2330(.A1(new_n2118_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2703_));
  NOR4_X1    g2331(.A1(new_n1160_), .A2(new_n1805_), .A3(new_n1243_), .A4(new_n2120_), .ZN(new_n2704_));
  OAI21_X1   g2332(.A1(new_n2703_), .A2(new_n2702_), .B(new_n2704_), .ZN(new_n2705_));
  OAI21_X1   g2333(.A1(new_n2705_), .A2(new_n2701_), .B(\shift[6] ), .ZN(new_n2706_));
  NAND2_X1   g2334(.A1(new_n2706_), .A2(new_n2698_), .ZN(\result[46] ));
  NOR4_X1    g2335(.A1(new_n1654_), .A2(new_n265_), .A3(new_n266_), .A4(new_n2137_), .ZN(new_n2708_));
  NOR3_X1    g2336(.A1(new_n2139_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2709_));
  NOR2_X1    g2337(.A1(new_n2709_), .A2(new_n2708_), .ZN(new_n2710_));
  NOR4_X1    g2338(.A1(new_n1826_), .A2(new_n1581_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2711_));
  NOR3_X1    g2339(.A1(new_n2126_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2712_));
  OAI21_X1   g2340(.A1(new_n2712_), .A2(new_n2711_), .B(new_n2453_), .ZN(new_n2713_));
  OAI21_X1   g2341(.A1(new_n2713_), .A2(new_n2710_), .B(new_n264_), .ZN(new_n2714_));
  OAI21_X1   g2342(.A1(new_n1469_), .A2(new_n2129_), .B(\shift[4] ), .ZN(new_n2715_));
  XOR2_X1    g2343(.A1(new_n2715_), .A2(new_n987_), .Z(new_n2716_));
  NOR4_X1    g2344(.A1(new_n1617_), .A2(new_n1846_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2717_));
  OAI21_X1   g2345(.A1(new_n1617_), .A2(new_n1846_), .B(\shift[5] ), .ZN(new_n2718_));
  NOR2_X1    g2346(.A1(new_n2718_), .A2(new_n987_), .ZN(new_n2719_));
  NOR4_X1    g2347(.A1(new_n1437_), .A2(new_n1542_), .A3(new_n2133_), .A4(new_n2145_), .ZN(new_n2720_));
  OAI21_X1   g2348(.A1(new_n2719_), .A2(new_n2717_), .B(new_n2720_), .ZN(new_n2721_));
  OAI21_X1   g2349(.A1(new_n2716_), .A2(new_n2721_), .B(\shift[6] ), .ZN(new_n2722_));
  NAND2_X1   g2350(.A1(new_n2722_), .A2(new_n2714_), .ZN(\result[47] ));
  NOR4_X1    g2351(.A1(new_n641_), .A2(new_n619_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2724_));
  NOR3_X1    g2352(.A1(new_n2165_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2725_));
  NOR2_X1    g2353(.A1(new_n2725_), .A2(new_n2724_), .ZN(new_n2726_));
  NOR4_X1    g2354(.A1(new_n694_), .A2(new_n571_), .A3(new_n594_), .A4(new_n654_), .ZN(new_n2727_));
  OAI21_X1   g2355(.A1(new_n2469_), .A2(new_n2468_), .B(new_n2727_), .ZN(new_n2728_));
  OAI21_X1   g2356(.A1(new_n2728_), .A2(new_n2726_), .B(new_n264_), .ZN(new_n2729_));
  NOR2_X1    g2357(.A1(new_n2017_), .A2(new_n2019_), .ZN(new_n2730_));
  NOR2_X1    g2358(.A1(new_n2378_), .A2(new_n2021_), .ZN(new_n2731_));
  NAND2_X1   g2359(.A1(new_n2731_), .A2(new_n2730_), .ZN(new_n2732_));
  NOR2_X1    g2360(.A1(new_n2014_), .A2(new_n2402_), .ZN(new_n2733_));
  NAND3_X1   g2361(.A1(new_n2398_), .A2(new_n2733_), .A3(new_n987_), .ZN(new_n2734_));
  NAND3_X1   g2362(.A1(new_n2734_), .A2(new_n2732_), .A3(new_n2283_), .ZN(new_n2735_));
  NAND3_X1   g2363(.A1(new_n383_), .A2(\shift[4] ), .A3(\shift[5] ), .ZN(new_n2736_));
  NOR2_X1    g2364(.A1(new_n543_), .A2(new_n266_), .ZN(new_n2737_));
  NOR2_X1    g2365(.A1(new_n2380_), .A2(new_n2384_), .ZN(new_n2738_));
  NAND2_X1   g2366(.A1(new_n461_), .A2(new_n456_), .ZN(new_n2739_));
  NOR2_X1    g2367(.A1(new_n2739_), .A2(new_n2387_), .ZN(new_n2740_));
  NAND3_X1   g2368(.A1(new_n2740_), .A2(new_n2738_), .A3(new_n987_), .ZN(new_n2741_));
  NAND3_X1   g2369(.A1(new_n2737_), .A2(new_n265_), .A3(new_n2741_), .ZN(new_n2742_));
  NAND4_X1   g2370(.A1(new_n2740_), .A2(new_n2738_), .A3(\shift[4] ), .A4(\shift[5] ), .ZN(new_n2743_));
  AOI22_X1   g2371(.A1(new_n2742_), .A2(new_n2743_), .B1(new_n2735_), .B2(new_n2736_), .ZN(new_n2744_));
  OAI21_X1   g2372(.A1(new_n2744_), .A2(new_n264_), .B(new_n2729_), .ZN(\result[48] ));
  NOR4_X1    g2373(.A1(new_n1784_), .A2(new_n265_), .A3(new_n266_), .A4(new_n998_), .ZN(new_n2746_));
  NOR3_X1    g2374(.A1(new_n1032_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2747_));
  NOR2_X1    g2375(.A1(new_n2746_), .A2(new_n2747_), .ZN(new_n2748_));
  NOR4_X1    g2376(.A1(new_n960_), .A2(new_n983_), .A3(new_n1058_), .A4(new_n1083_), .ZN(new_n2749_));
  OAI21_X1   g2377(.A1(new_n2485_), .A2(new_n2484_), .B(new_n2749_), .ZN(new_n2750_));
  OAI21_X1   g2378(.A1(new_n2750_), .A2(new_n2748_), .B(new_n264_), .ZN(new_n2751_));
  OAI21_X1   g2379(.A1(new_n820_), .A2(new_n842_), .B(\shift[4] ), .ZN(new_n2752_));
  XOR2_X1    g2380(.A1(new_n2752_), .A2(new_n987_), .Z(new_n2753_));
  NOR4_X1    g2381(.A1(new_n865_), .A2(new_n889_), .A3(new_n916_), .A4(new_n937_), .ZN(new_n2754_));
  OAI21_X1   g2382(.A1(new_n798_), .A2(new_n796_), .B(new_n2754_), .ZN(new_n2755_));
  OAI21_X1   g2383(.A1(new_n2753_), .A2(new_n2755_), .B(\shift[6] ), .ZN(new_n2756_));
  NAND2_X1   g2384(.A1(new_n2751_), .A2(new_n2756_), .ZN(\result[49] ));
  NOR4_X1    g2385(.A1(new_n1360_), .A2(new_n1379_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2758_));
  NOR3_X1    g2386(.A1(new_n2200_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2759_));
  NOR2_X1    g2387(.A1(new_n2759_), .A2(new_n2758_), .ZN(new_n2760_));
  NOR4_X1    g2388(.A1(new_n1321_), .A2(new_n1339_), .A3(new_n1397_), .A4(new_n1414_), .ZN(new_n2761_));
  OAI21_X1   g2389(.A1(new_n2502_), .A2(new_n2501_), .B(new_n2761_), .ZN(new_n2762_));
  OAI21_X1   g2390(.A1(new_n2760_), .A2(new_n2762_), .B(new_n264_), .ZN(new_n2763_));
  NOR4_X1    g2391(.A1(new_n1203_), .A2(new_n1224_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2764_));
  NOR3_X1    g2392(.A1(new_n2193_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2765_));
  NOR2_X1    g2393(.A1(new_n2765_), .A2(new_n2764_), .ZN(new_n2766_));
  NOR4_X1    g2394(.A1(new_n1243_), .A2(new_n1284_), .A3(new_n1261_), .A4(new_n1303_), .ZN(new_n2767_));
  OAI21_X1   g2395(.A1(new_n1185_), .A2(new_n1183_), .B(new_n2767_), .ZN(new_n2768_));
  OAI21_X1   g2396(.A1(new_n2768_), .A2(new_n2766_), .B(\shift[6] ), .ZN(new_n2769_));
  NAND2_X1   g2397(.A1(new_n2769_), .A2(new_n2763_), .ZN(\result[50] ));
  NOR4_X1    g2398(.A1(new_n1509_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1525_), .ZN(new_n2771_));
  NOR3_X1    g2399(.A1(new_n2210_), .A2(\shift[4] ), .A3(new_n266_), .ZN(new_n2772_));
  NOR2_X1    g2400(.A1(new_n2772_), .A2(new_n2771_), .ZN(new_n2773_));
  NOR4_X1    g2401(.A1(new_n1654_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1673_), .ZN(new_n2774_));
  NOR3_X1    g2402(.A1(new_n2220_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2775_));
  NOR4_X1    g2403(.A1(new_n1581_), .A2(new_n1690_), .A3(new_n1599_), .A4(new_n1709_), .ZN(new_n2776_));
  OAI21_X1   g2404(.A1(new_n2775_), .A2(new_n2774_), .B(new_n2776_), .ZN(new_n2777_));
  OAI21_X1   g2405(.A1(new_n2773_), .A2(new_n2777_), .B(new_n264_), .ZN(new_n2778_));
  OAI21_X1   g2406(.A1(new_n1617_), .A2(new_n1633_), .B(new_n984_), .ZN(new_n2779_));
  XOR2_X1    g2407(.A1(new_n2779_), .A2(new_n1454_), .Z(new_n2780_));
  NOR3_X1    g2408(.A1(new_n1469_), .A2(new_n893_), .A3(new_n1488_), .ZN(new_n2781_));
  XOR2_X1    g2409(.A1(new_n1561_), .A2(new_n2781_), .Z(new_n2782_));
  OAI21_X1   g2410(.A1(new_n2780_), .A2(new_n2782_), .B(\shift[6] ), .ZN(new_n2783_));
  NAND2_X1   g2411(.A1(new_n2783_), .A2(new_n2778_), .ZN(\result[51] ));
  NOR3_X1    g2412(.A1(new_n291_), .A2(new_n1714_), .A3(new_n893_), .ZN(new_n2785_));
  NOR4_X1    g2413(.A1(new_n2785_), .A2(\shift[4] ), .A3(new_n266_), .A4(new_n1745_), .ZN(new_n2786_));
  NOR3_X1    g2414(.A1(new_n2534_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n2787_));
  NOR2_X1    g2415(.A1(new_n2786_), .A2(new_n2787_), .ZN(new_n2788_));
  NOR3_X1    g2416(.A1(new_n1748_), .A2(new_n619_), .A3(new_n893_), .ZN(new_n2789_));
  OAI21_X1   g2417(.A1(new_n1754_), .A2(new_n1755_), .B(new_n984_), .ZN(new_n2790_));
  NOR2_X1    g2418(.A1(new_n2790_), .A2(new_n2789_), .ZN(new_n2791_));
  NOR4_X1    g2419(.A1(new_n1748_), .A2(new_n619_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2793_));
  NOR2_X1    g2420(.A1(new_n2791_), .A2(new_n2793_), .ZN(new_n2794_));
  OAI21_X1   g2421(.A1(new_n2788_), .A2(new_n2794_), .B(new_n264_), .ZN(new_n2795_));
  NOR3_X1    g2422(.A1(new_n1723_), .A2(new_n1724_), .A3(new_n893_), .ZN(new_n2796_));
  NOR3_X1    g2423(.A1(new_n2796_), .A2(new_n2230_), .A3(new_n2309_), .ZN(new_n2797_));
  NOR4_X1    g2424(.A1(new_n1723_), .A2(new_n1724_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2798_));
  NOR2_X1    g2425(.A1(new_n2797_), .A2(new_n2798_), .ZN(new_n2799_));
  NOR3_X1    g2426(.A1(new_n452_), .A2(new_n1729_), .A3(new_n893_), .ZN(new_n2800_));
  OAI21_X1   g2427(.A1(new_n1752_), .A2(new_n1753_), .B(new_n984_), .ZN(new_n2801_));
  NOR2_X1    g2428(.A1(new_n2801_), .A2(new_n2800_), .ZN(new_n2802_));
  NOR4_X1    g2429(.A1(new_n452_), .A2(new_n1729_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2803_));
  NOR2_X1    g2430(.A1(new_n2802_), .A2(new_n2803_), .ZN(new_n2804_));
  OAI21_X1   g2431(.A1(new_n2799_), .A2(new_n2804_), .B(\shift[6] ), .ZN(new_n2805_));
  NAND2_X1   g2432(.A1(new_n2795_), .A2(new_n2805_), .ZN(\result[52] ));
  NOR3_X1    g2433(.A1(new_n1760_), .A2(new_n893_), .A3(new_n719_), .ZN(new_n2807_));
  NOR4_X1    g2434(.A1(new_n2807_), .A2(\shift[4] ), .A3(new_n266_), .A4(new_n1786_), .ZN(new_n2808_));
  NOR4_X1    g2435(.A1(new_n1760_), .A2(new_n265_), .A3(new_n266_), .A4(new_n719_), .ZN(new_n2809_));
  NOR2_X1    g2436(.A1(new_n2808_), .A2(new_n2809_), .ZN(new_n2810_));
  NAND2_X1   g2437(.A1(new_n1038_), .A2(new_n1044_), .ZN(new_n2811_));
  NOR4_X1    g2438(.A1(new_n1778_), .A2(new_n893_), .A3(new_n998_), .A4(new_n2811_), .ZN(new_n2812_));
  OAI21_X1   g2439(.A1(new_n960_), .A2(new_n1790_), .B(new_n984_), .ZN(new_n2813_));
  XOR2_X1    g2440(.A1(new_n2812_), .A2(new_n2813_), .Z(new_n2814_));
  OAI21_X1   g2441(.A1(new_n2810_), .A2(new_n2814_), .B(new_n264_), .ZN(new_n2815_));
  NOR3_X1    g2442(.A1(new_n1765_), .A2(new_n1766_), .A3(new_n893_), .ZN(new_n2816_));
  OAI21_X1   g2443(.A1(new_n820_), .A2(new_n1770_), .B(new_n2283_), .ZN(new_n2817_));
  XOR2_X1    g2444(.A1(new_n2817_), .A2(new_n2816_), .Z(new_n2818_));
  NOR3_X1    g2445(.A1(new_n865_), .A2(new_n1771_), .A3(new_n893_), .ZN(new_n2819_));
  OAI21_X1   g2446(.A1(new_n1788_), .A2(new_n1789_), .B(new_n984_), .ZN(new_n2820_));
  XOR2_X1    g2447(.A1(new_n2820_), .A2(new_n2819_), .Z(new_n2821_));
  OAI21_X1   g2448(.A1(new_n2818_), .A2(new_n2821_), .B(\shift[6] ), .ZN(new_n2822_));
  NAND2_X1   g2449(.A1(new_n2815_), .A2(new_n2822_), .ZN(\result[53] ));
  NOR3_X1    g2450(.A1(new_n1108_), .A2(new_n1795_), .A3(new_n893_), .ZN(new_n2824_));
  NOR3_X1    g2451(.A1(new_n2572_), .A2(new_n2824_), .A3(\shift[4] ), .ZN(new_n2825_));
  NOR4_X1    g2452(.A1(new_n1108_), .A2(new_n1795_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2826_));
  NOR2_X1    g2453(.A1(new_n2825_), .A2(new_n2826_), .ZN(new_n2827_));
  NOR3_X1    g2454(.A1(new_n1810_), .A2(new_n1811_), .A3(new_n893_), .ZN(new_n2828_));
  OAI21_X1   g2455(.A1(new_n1321_), .A2(new_n1821_), .B(new_n984_), .ZN(new_n2829_));
  NOR2_X1    g2456(.A1(new_n2829_), .A2(new_n2828_), .ZN(new_n2830_));
  NOR4_X1    g2457(.A1(new_n1810_), .A2(new_n1811_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2832_));
  NOR2_X1    g2458(.A1(new_n2830_), .A2(new_n2832_), .ZN(new_n2833_));
  OAI21_X1   g2459(.A1(new_n2827_), .A2(new_n2833_), .B(new_n264_), .ZN(new_n2834_));
  NOR3_X1    g2460(.A1(new_n1800_), .A2(new_n1801_), .A3(new_n893_), .ZN(new_n2835_));
  NOR3_X1    g2461(.A1(new_n2835_), .A2(new_n2260_), .A3(new_n2309_), .ZN(new_n2836_));
  NOR4_X1    g2462(.A1(new_n1800_), .A2(new_n1801_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2837_));
  NOR2_X1    g2463(.A1(new_n2836_), .A2(new_n2837_), .ZN(new_n2838_));
  NOR3_X1    g2464(.A1(new_n1243_), .A2(new_n1806_), .A3(new_n893_), .ZN(new_n2839_));
  OAI21_X1   g2465(.A1(new_n1820_), .A2(new_n1819_), .B(new_n984_), .ZN(new_n2840_));
  NOR2_X1    g2466(.A1(new_n2840_), .A2(new_n2839_), .ZN(new_n2841_));
  NOR4_X1    g2467(.A1(new_n1243_), .A2(new_n1806_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2842_));
  NOR2_X1    g2468(.A1(new_n2841_), .A2(new_n2842_), .ZN(new_n2843_));
  OAI21_X1   g2469(.A1(new_n2838_), .A2(new_n2843_), .B(\shift[6] ), .ZN(new_n2844_));
  NAND2_X1   g2470(.A1(new_n2834_), .A2(new_n2844_), .ZN(\result[54] ));
  NOR2_X1    g2471(.A1(new_n2592_), .A2(new_n2591_), .ZN(new_n2846_));
  NOR4_X1    g2472(.A1(new_n1854_), .A2(new_n1855_), .A3(new_n1842_), .A4(new_n1843_), .ZN(new_n2847_));
  OAI21_X1   g2473(.A1(new_n1829_), .A2(new_n1827_), .B(new_n2847_), .ZN(new_n2848_));
  OAI21_X1   g2474(.A1(new_n2848_), .A2(new_n2846_), .B(new_n264_), .ZN(new_n2849_));
  OAI21_X1   g2475(.A1(new_n1836_), .A2(new_n1837_), .B(\shift[4] ), .ZN(new_n2850_));
  XOR2_X1    g2476(.A1(new_n2850_), .A2(new_n987_), .Z(new_n2851_));
  NOR4_X1    g2477(.A1(new_n1437_), .A2(new_n1838_), .A3(new_n1853_), .A4(new_n1852_), .ZN(new_n2852_));
  OAI21_X1   g2478(.A1(new_n1835_), .A2(new_n1833_), .B(new_n2852_), .ZN(new_n2853_));
  OAI21_X1   g2479(.A1(new_n2851_), .A2(new_n2853_), .B(\shift[6] ), .ZN(new_n2854_));
  NAND2_X1   g2480(.A1(new_n2849_), .A2(new_n2854_), .ZN(\result[55] ));
  NOR2_X1    g2481(.A1(new_n2609_), .A2(new_n2608_), .ZN(new_n2856_));
  NOR4_X1    g2482(.A1(new_n1877_), .A2(new_n1755_), .A3(new_n1893_), .A4(new_n654_), .ZN(new_n2857_));
  OAI21_X1   g2483(.A1(new_n1864_), .A2(new_n1862_), .B(new_n2857_), .ZN(new_n2858_));
  OAI21_X1   g2484(.A1(new_n2858_), .A2(new_n2856_), .B(new_n264_), .ZN(new_n2859_));
  NOR4_X1    g2485(.A1(new_n1871_), .A2(new_n1870_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2860_));
  OAI21_X1   g2486(.A1(new_n1871_), .A2(new_n1870_), .B(\shift[4] ), .ZN(new_n2861_));
  NOR2_X1    g2487(.A1(new_n2861_), .A2(new_n987_), .ZN(new_n2862_));
  NOR2_X1    g2488(.A1(new_n2862_), .A2(new_n2860_), .ZN(new_n2863_));
  NOR4_X1    g2489(.A1(new_n1753_), .A2(new_n1873_), .A3(new_n1887_), .A4(new_n1872_), .ZN(new_n2864_));
  OAI21_X1   g2490(.A1(new_n1869_), .A2(new_n1867_), .B(new_n2864_), .ZN(new_n2865_));
  OAI21_X1   g2491(.A1(new_n2865_), .A2(new_n2863_), .B(\shift[6] ), .ZN(new_n2866_));
  NAND2_X1   g2492(.A1(new_n2866_), .A2(new_n2859_), .ZN(\result[56] ));
  NOR2_X1    g2493(.A1(new_n2624_), .A2(new_n2625_), .ZN(new_n2868_));
  NOR4_X1    g2494(.A1(new_n1915_), .A2(new_n1778_), .A3(new_n1927_), .A4(new_n1928_), .ZN(new_n2869_));
  OAI21_X1   g2495(.A1(new_n1902_), .A2(new_n1900_), .B(new_n2869_), .ZN(new_n2870_));
  OAI21_X1   g2496(.A1(new_n2870_), .A2(new_n2868_), .B(new_n264_), .ZN(new_n2871_));
  OAI21_X1   g2497(.A1(new_n1908_), .A2(new_n1909_), .B(\shift[4] ), .ZN(new_n2872_));
  XOR2_X1    g2498(.A1(new_n2872_), .A2(new_n987_), .Z(new_n2873_));
  NOR4_X1    g2499(.A1(new_n1789_), .A2(new_n1910_), .A3(new_n1911_), .A4(new_n1926_), .ZN(new_n2874_));
  OAI21_X1   g2500(.A1(new_n1907_), .A2(new_n1905_), .B(new_n2874_), .ZN(new_n2875_));
  OAI21_X1   g2501(.A1(new_n2873_), .A2(new_n2875_), .B(\shift[6] ), .ZN(new_n2876_));
  NAND2_X1   g2502(.A1(new_n2871_), .A2(new_n2876_), .ZN(\result[57] ));
  NOR3_X1    g2503(.A1(new_n1934_), .A2(new_n1933_), .A3(new_n893_), .ZN(new_n2878_));
  NOR3_X1    g2504(.A1(new_n2640_), .A2(new_n2878_), .A3(\shift[4] ), .ZN(new_n2879_));
  NOR4_X1    g2505(.A1(new_n1934_), .A2(new_n1933_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2880_));
  NOR2_X1    g2506(.A1(new_n2879_), .A2(new_n2880_), .ZN(new_n2881_));
  NOR2_X1    g2507(.A1(new_n1965_), .A2(new_n1966_), .ZN(new_n2882_));
  NOR3_X1    g2508(.A1(new_n1957_), .A2(new_n1811_), .A3(new_n893_), .ZN(new_n2883_));
  NOR3_X1    g2509(.A1(new_n2883_), .A2(new_n2882_), .A3(new_n1265_), .ZN(new_n2884_));
  NOR4_X1    g2510(.A1(new_n1957_), .A2(new_n1811_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2885_));
  NOR2_X1    g2511(.A1(new_n2884_), .A2(new_n2885_), .ZN(new_n2886_));
  OAI21_X1   g2512(.A1(new_n2881_), .A2(new_n2886_), .B(new_n264_), .ZN(new_n2887_));
  NOR4_X1    g2513(.A1(new_n1951_), .A2(new_n1950_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2888_));
  NOR3_X1    g2514(.A1(new_n2342_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2889_));
  NOR2_X1    g2515(.A1(new_n2889_), .A2(new_n2888_), .ZN(new_n2890_));
  NOR4_X1    g2516(.A1(new_n1820_), .A2(new_n1953_), .A3(new_n1964_), .A4(new_n1952_), .ZN(new_n2891_));
  OAI21_X1   g2517(.A1(new_n1949_), .A2(new_n1947_), .B(new_n2891_), .ZN(new_n2892_));
  OAI21_X1   g2518(.A1(new_n2892_), .A2(new_n2890_), .B(\shift[6] ), .ZN(new_n2893_));
  NAND2_X1   g2519(.A1(new_n2887_), .A2(new_n2893_), .ZN(\result[58] ));
  NAND2_X1   g2520(.A1(new_n1508_), .A2(new_n1504_), .ZN(new_n2895_));
  NAND2_X1   g2521(.A1(new_n1517_), .A2(new_n1513_), .ZN(new_n2896_));
  NOR4_X1    g2522(.A1(new_n2895_), .A2(new_n1972_), .A3(new_n893_), .A4(new_n2896_), .ZN(new_n2897_));
  NOR4_X1    g2523(.A1(new_n2897_), .A2(\shift[4] ), .A3(new_n1994_), .A4(new_n266_), .ZN(new_n2898_));
  NOR4_X1    g2524(.A1(new_n1971_), .A2(new_n265_), .A3(new_n266_), .A4(new_n1972_), .ZN(new_n2899_));
  NOR2_X1    g2525(.A1(new_n2898_), .A2(new_n2899_), .ZN(new_n2900_));
  NOR3_X1    g2526(.A1(new_n1843_), .A2(new_n1987_), .A3(new_n893_), .ZN(new_n2901_));
  OAI21_X1   g2527(.A1(new_n1855_), .A2(new_n1997_), .B(new_n984_), .ZN(new_n2902_));
  XOR2_X1    g2528(.A1(new_n2902_), .A2(new_n2901_), .Z(new_n2903_));
  OAI21_X1   g2529(.A1(new_n2900_), .A2(new_n2903_), .B(new_n264_), .ZN(new_n2904_));
  OAI21_X1   g2530(.A1(new_n1981_), .A2(new_n1837_), .B(\shift[4] ), .ZN(new_n2905_));
  XOR2_X1    g2531(.A1(new_n2905_), .A2(new_n987_), .Z(new_n2906_));
  NOR4_X1    g2532(.A1(new_n1853_), .A2(new_n1982_), .A3(new_n1983_), .A4(new_n1996_), .ZN(new_n2907_));
  OAI21_X1   g2533(.A1(new_n1980_), .A2(new_n1978_), .B(new_n2907_), .ZN(new_n2908_));
  OAI21_X1   g2534(.A1(new_n2906_), .A2(new_n2908_), .B(\shift[6] ), .ZN(new_n2909_));
  NAND2_X1   g2535(.A1(new_n2904_), .A2(new_n2909_), .ZN(\result[59] ));
  NOR2_X1    g2536(.A1(new_n2046_), .A2(new_n266_), .ZN(new_n2911_));
  NAND2_X1   g2537(.A1(new_n2006_), .A2(new_n987_), .ZN(new_n2912_));
  NAND3_X1   g2538(.A1(new_n2911_), .A2(new_n2912_), .A3(new_n265_), .ZN(new_n2913_));
  NAND3_X1   g2539(.A1(new_n2006_), .A2(\shift[4] ), .A3(\shift[5] ), .ZN(new_n2914_));
  AND2_X2    g2540(.A1(new_n581_), .A2(new_n575_), .Z(new_n2915_));
  INV_X1     g2541(.I(new_n601_), .ZN(new_n2916_));
  NOR3_X1    g2542(.A1(new_n2916_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n2917_));
  NAND4_X1   g2543(.A1(new_n2915_), .A2(new_n2917_), .A3(new_n618_), .A4(new_n640_), .ZN(new_n2918_));
  NAND2_X1   g2544(.A1(new_n2040_), .A2(new_n987_), .ZN(new_n2919_));
  NAND3_X1   g2545(.A1(new_n2919_), .A2(new_n2918_), .A3(new_n984_), .ZN(new_n2920_));
  NAND3_X1   g2546(.A1(new_n2040_), .A2(\shift[4] ), .A3(\shift[5] ), .ZN(new_n2922_));
  AOI22_X1   g2547(.A1(new_n2913_), .A2(new_n2914_), .B1(new_n2920_), .B2(new_n2922_), .ZN(new_n2923_));
  NOR4_X1    g2548(.A1(new_n452_), .A2(new_n1728_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2924_));
  NOR3_X1    g2549(.A1(new_n2388_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2925_));
  NOR2_X1    g2550(.A1(new_n2925_), .A2(new_n2924_), .ZN(new_n2926_));
  NOR4_X1    g2551(.A1(new_n291_), .A2(new_n2048_), .A3(new_n361_), .A4(new_n1729_), .ZN(new_n2927_));
  OAI21_X1   g2552(.A1(new_n2023_), .A2(new_n2010_), .B(new_n2927_), .ZN(new_n2928_));
  OAI21_X1   g2553(.A1(new_n2928_), .A2(new_n2926_), .B(\shift[6] ), .ZN(new_n2929_));
  OAI21_X1   g2554(.A1(new_n2923_), .A2(\shift[6] ), .B(new_n2929_), .ZN(\result[60] ));
  NOR3_X1    g2555(.A1(new_n1760_), .A2(new_n893_), .A3(new_n960_), .ZN(new_n2931_));
  NOR3_X1    g2556(.A1(new_n2931_), .A2(\shift[4] ), .A3(new_n2686_), .ZN(new_n2932_));
  NOR4_X1    g2557(.A1(new_n1760_), .A2(new_n265_), .A3(new_n266_), .A4(new_n960_), .ZN(new_n2933_));
  NOR2_X1    g2558(.A1(new_n2932_), .A2(new_n2933_), .ZN(new_n2934_));
  OAI21_X1   g2559(.A1(new_n1058_), .A2(new_n1790_), .B(new_n984_), .ZN(new_n2935_));
  AOI21_X1   g2560(.A1(new_n987_), .A2(new_n2066_), .B(new_n2935_), .ZN(new_n2936_));
  AND3_X2    g2561(.A1(new_n2935_), .A2(new_n987_), .A3(new_n2066_), .Z(new_n2937_));
  NOR2_X1    g2562(.A1(new_n2937_), .A2(new_n2936_), .ZN(new_n2938_));
  OAI21_X1   g2563(.A1(new_n2938_), .A2(new_n2934_), .B(new_n264_), .ZN(new_n2939_));
  OAI21_X1   g2564(.A1(new_n865_), .A2(new_n1770_), .B(\shift[4] ), .ZN(new_n2940_));
  XOR2_X1    g2565(.A1(new_n2940_), .A2(new_n987_), .Z(new_n2941_));
  NOR4_X1    g2566(.A1(new_n719_), .A2(new_n771_), .A3(new_n1771_), .A4(new_n2074_), .ZN(new_n2942_));
  OAI21_X1   g2567(.A1(new_n2061_), .A2(new_n2059_), .B(new_n2942_), .ZN(new_n2943_));
  OAI21_X1   g2568(.A1(new_n2941_), .A2(new_n2943_), .B(\shift[6] ), .ZN(new_n2944_));
  NAND2_X1   g2569(.A1(new_n2939_), .A2(new_n2944_), .ZN(\result[61] ));
  NOR3_X1    g2570(.A1(new_n1321_), .A2(new_n1795_), .A3(new_n893_), .ZN(new_n2946_));
  NOR4_X1    g2571(.A1(new_n2946_), .A2(\shift[4] ), .A3(new_n2118_), .A4(new_n266_), .ZN(new_n2947_));
  NOR4_X1    g2572(.A1(new_n1321_), .A2(new_n1795_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2948_));
  NOR2_X1    g2573(.A1(new_n2947_), .A2(new_n2948_), .ZN(new_n2949_));
  NOR2_X1    g2574(.A1(new_n1821_), .A2(new_n1397_), .ZN(new_n2950_));
  NOR3_X1    g2575(.A1(new_n1360_), .A2(new_n2102_), .A3(new_n893_), .ZN(new_n2951_));
  NOR3_X1    g2576(.A1(new_n2951_), .A2(new_n2950_), .A3(new_n1265_), .ZN(new_n2952_));
  NOR4_X1    g2577(.A1(new_n1360_), .A2(new_n2102_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2953_));
  NOR2_X1    g2578(.A1(new_n2952_), .A2(new_n2953_), .ZN(new_n2954_));
  OAI21_X1   g2579(.A1(new_n2949_), .A2(new_n2954_), .B(new_n264_), .ZN(new_n2955_));
  NOR4_X1    g2580(.A1(new_n1805_), .A2(new_n1243_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2956_));
  NOR3_X1    g2581(.A1(new_n2434_), .A2(new_n265_), .A3(\shift[5] ), .ZN(new_n2957_));
  NOR2_X1    g2582(.A1(new_n2957_), .A2(new_n2956_), .ZN(new_n2958_));
  NOR4_X1    g2583(.A1(new_n1160_), .A2(new_n1108_), .A3(new_n2120_), .A4(new_n1806_), .ZN(new_n2959_));
  OAI21_X1   g2584(.A1(new_n2098_), .A2(new_n2087_), .B(new_n2959_), .ZN(new_n2960_));
  OAI21_X1   g2585(.A1(new_n2958_), .A2(new_n2960_), .B(\shift[6] ), .ZN(new_n2961_));
  NAND2_X1   g2586(.A1(new_n2955_), .A2(new_n2961_), .ZN(\result[62] ));
  NOR3_X1    g2587(.A1(new_n1826_), .A2(new_n1581_), .A3(new_n893_), .ZN(new_n2963_));
  NOR3_X1    g2588(.A1(new_n2963_), .A2(new_n2718_), .A3(\shift[4] ), .ZN(new_n2964_));
  NOR4_X1    g2589(.A1(new_n1826_), .A2(new_n1581_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n2965_));
  NOR2_X1    g2590(.A1(new_n2964_), .A2(new_n2965_), .ZN(new_n2966_));
  OAI21_X1   g2591(.A1(new_n1690_), .A2(new_n2146_), .B(new_n984_), .ZN(new_n2967_));
  AOI21_X1   g2592(.A1(new_n987_), .A2(new_n2139_), .B(new_n2967_), .ZN(new_n2968_));
  NOR4_X1    g2593(.A1(new_n1654_), .A2(new_n265_), .A3(new_n266_), .A4(new_n2137_), .ZN(new_n2970_));
  NOR2_X1    g2594(.A1(new_n2968_), .A2(new_n2970_), .ZN(new_n2971_));
  OAI21_X1   g2595(.A1(new_n2971_), .A2(new_n2966_), .B(new_n264_), .ZN(new_n2972_));
  OAI21_X1   g2596(.A1(new_n1437_), .A2(new_n2133_), .B(\shift[4] ), .ZN(new_n2973_));
  XOR2_X1    g2597(.A1(new_n2973_), .A2(new_n987_), .Z(new_n2974_));
  NOR4_X1    g2598(.A1(new_n1509_), .A2(new_n1542_), .A3(new_n1838_), .A4(new_n2145_), .ZN(new_n2975_));
  OAI21_X1   g2599(.A1(new_n2132_), .A2(new_n2130_), .B(new_n2975_), .ZN(new_n2976_));
  OAI21_X1   g2600(.A1(new_n2974_), .A2(new_n2976_), .B(\shift[6] ), .ZN(new_n2977_));
  NAND2_X1   g2601(.A1(new_n2972_), .A2(new_n2977_), .ZN(\result[63] ));
  OAI21_X1   g2602(.A1(new_n696_), .A2(new_n545_), .B(new_n264_), .ZN(new_n2979_));
  OAI21_X1   g2603(.A1(new_n477_), .A2(new_n337_), .B(\shift[6] ), .ZN(new_n2980_));
  NAND2_X1   g2604(.A1(new_n2980_), .A2(new_n2979_), .ZN(\result[64] ));
  OAI21_X1   g2605(.A1(new_n1087_), .A2(new_n986_), .B(new_n264_), .ZN(new_n2982_));
  OAI21_X1   g2606(.A1(new_n748_), .A2(new_n891_), .B(\shift[6] ), .ZN(new_n2983_));
  NAND2_X1   g2607(.A1(new_n2982_), .A2(new_n2983_), .ZN(\result[65] ));
  OAI21_X1   g2608(.A1(new_n1343_), .A2(new_n1418_), .B(new_n264_), .ZN(new_n2985_));
  OAI21_X1   g2609(.A1(new_n1263_), .A2(new_n1142_), .B(\shift[6] ), .ZN(new_n2986_));
  NAND2_X1   g2610(.A1(new_n2985_), .A2(new_n2986_), .ZN(\result[66] ));
  OAI21_X1   g2611(.A1(new_n1601_), .A2(new_n1711_), .B(new_n264_), .ZN(new_n2988_));
  OAI21_X1   g2612(.A1(new_n1565_), .A2(new_n1493_), .B(\shift[6] ), .ZN(new_n2989_));
  NAND2_X1   g2613(.A1(new_n2988_), .A2(new_n2989_), .ZN(\result[67] ));
  OAI21_X1   g2614(.A1(new_n1757_), .A2(new_n1747_), .B(new_n264_), .ZN(new_n2991_));
  OAI21_X1   g2615(.A1(new_n1731_), .A2(new_n1722_), .B(\shift[6] ), .ZN(new_n2992_));
  NAND2_X1   g2616(.A1(new_n2991_), .A2(new_n2992_), .ZN(\result[68] ));
  OAI21_X1   g2617(.A1(new_n1782_), .A2(new_n1792_), .B(new_n264_), .ZN(new_n2994_));
  OAI21_X1   g2618(.A1(new_n1764_), .A2(new_n1773_), .B(\shift[6] ), .ZN(new_n2995_));
  NAND2_X1   g2619(.A1(new_n2994_), .A2(new_n2995_), .ZN(\result[69] ));
  OAI21_X1   g2620(.A1(new_n1813_), .A2(new_n1823_), .B(new_n264_), .ZN(new_n2997_));
  OAI21_X1   g2621(.A1(new_n1808_), .A2(new_n1799_), .B(\shift[6] ), .ZN(new_n2998_));
  NAND2_X1   g2622(.A1(new_n2997_), .A2(new_n2998_), .ZN(\result[70] ));
  OAI21_X1   g2623(.A1(new_n1845_), .A2(new_n1857_), .B(new_n264_), .ZN(new_n3000_));
  OAI21_X1   g2624(.A1(new_n1830_), .A2(new_n1840_), .B(\shift[6] ), .ZN(new_n3001_));
  NAND2_X1   g2625(.A1(new_n3000_), .A2(new_n3001_), .ZN(\result[71] ));
  OAI21_X1   g2626(.A1(new_n1881_), .A2(new_n1895_), .B(new_n264_), .ZN(new_n3003_));
  OAI21_X1   g2627(.A1(new_n1875_), .A2(new_n1865_), .B(\shift[6] ), .ZN(new_n3004_));
  NAND2_X1   g2628(.A1(new_n3004_), .A2(new_n3003_), .ZN(\result[72] ));
  OAI21_X1   g2629(.A1(new_n1919_), .A2(new_n1930_), .B(new_n264_), .ZN(new_n3006_));
  OAI21_X1   g2630(.A1(new_n1903_), .A2(new_n1913_), .B(\shift[6] ), .ZN(new_n3007_));
  NAND2_X1   g2631(.A1(new_n3006_), .A2(new_n3007_), .ZN(\result[73] ));
  OAI21_X1   g2632(.A1(new_n1959_), .A2(new_n1968_), .B(new_n264_), .ZN(new_n3009_));
  OAI21_X1   g2633(.A1(new_n1955_), .A2(new_n1945_), .B(\shift[6] ), .ZN(new_n3010_));
  NAND2_X1   g2634(.A1(new_n3009_), .A2(new_n3010_), .ZN(\result[74] ));
  OAI21_X1   g2635(.A1(new_n1999_), .A2(new_n1989_), .B(new_n264_), .ZN(new_n3012_));
  OAI21_X1   g2636(.A1(new_n1976_), .A2(new_n1985_), .B(\shift[6] ), .ZN(new_n3013_));
  NAND2_X1   g2637(.A1(new_n3012_), .A2(new_n3013_), .ZN(\result[75] ));
  OAI21_X1   g2638(.A1(new_n2051_), .A2(new_n2042_), .B(new_n264_), .ZN(new_n3015_));
  OAI21_X1   g2639(.A1(new_n2025_), .A2(new_n2008_), .B(\shift[6] ), .ZN(new_n3016_));
  NAND2_X1   g2640(.A1(new_n3015_), .A2(new_n3016_), .ZN(\result[76] ));
  OAI21_X1   g2641(.A1(new_n2070_), .A2(new_n2076_), .B(new_n264_), .ZN(new_n3018_));
  OAI21_X1   g2642(.A1(new_n2057_), .A2(new_n2063_), .B(\shift[6] ), .ZN(new_n3019_));
  NAND2_X1   g2643(.A1(new_n3018_), .A2(new_n3019_), .ZN(\result[77] ));
  OAI21_X1   g2644(.A1(new_n2122_), .A2(new_n2106_), .B(new_n264_), .ZN(new_n3021_));
  OAI21_X1   g2645(.A1(new_n2100_), .A2(new_n2085_), .B(\shift[6] ), .ZN(new_n3022_));
  NAND2_X1   g2646(.A1(new_n3021_), .A2(new_n3022_), .ZN(\result[78] ));
  OAI21_X1   g2647(.A1(new_n2148_), .A2(new_n2141_), .B(new_n264_), .ZN(new_n3024_));
  OAI21_X1   g2648(.A1(new_n2135_), .A2(new_n2128_), .B(\shift[6] ), .ZN(new_n3025_));
  NAND2_X1   g2649(.A1(new_n3025_), .A2(new_n3024_), .ZN(\result[79] ));
  OAI21_X1   g2650(.A1(new_n2174_), .A2(new_n2169_), .B(new_n264_), .ZN(new_n3027_));
  OAI21_X1   g2651(.A1(new_n2154_), .A2(new_n2156_), .B(\shift[6] ), .ZN(new_n3028_));
  NAND2_X1   g2652(.A1(new_n3027_), .A2(new_n3028_), .ZN(\result[80] ));
  OAI21_X1   g2653(.A1(new_n2185_), .A2(new_n2189_), .B(new_n264_), .ZN(new_n3030_));
  OAI21_X1   g2654(.A1(new_n2180_), .A2(new_n2178_), .B(\shift[6] ), .ZN(new_n3031_));
  NAND2_X1   g2655(.A1(new_n3031_), .A2(new_n3030_), .ZN(\result[81] ));
  OAI21_X1   g2656(.A1(new_n2206_), .A2(new_n2202_), .B(new_n264_), .ZN(new_n3033_));
  OAI21_X1   g2657(.A1(new_n2195_), .A2(new_n2197_), .B(\shift[6] ), .ZN(new_n3034_));
  NAND2_X1   g2658(.A1(new_n3033_), .A2(new_n3034_), .ZN(\result[82] ));
  OAI21_X1   g2659(.A1(new_n2226_), .A2(new_n2222_), .B(new_n264_), .ZN(new_n3036_));
  OAI21_X1   g2660(.A1(new_n2212_), .A2(new_n2217_), .B(\shift[6] ), .ZN(new_n3037_));
  NAND2_X1   g2661(.A1(new_n3037_), .A2(new_n3036_), .ZN(\result[83] ));
  OAI21_X1   g2662(.A1(new_n2241_), .A2(new_n2239_), .B(new_n264_), .ZN(new_n3039_));
  OAI21_X1   g2663(.A1(new_n2232_), .A2(new_n2234_), .B(\shift[6] ), .ZN(new_n3040_));
  NAND2_X1   g2664(.A1(new_n3039_), .A2(new_n3040_), .ZN(\result[84] ));
  OAI21_X1   g2665(.A1(new_n2252_), .A2(new_n2250_), .B(new_n264_), .ZN(new_n3042_));
  OAI21_X1   g2666(.A1(new_n2247_), .A2(new_n2245_), .B(\shift[6] ), .ZN(new_n3043_));
  NAND2_X1   g2667(.A1(new_n3042_), .A2(new_n3043_), .ZN(\result[85] ));
  OAI21_X1   g2668(.A1(new_n2271_), .A2(new_n2269_), .B(new_n264_), .ZN(new_n3045_));
  OAI21_X1   g2669(.A1(new_n2264_), .A2(new_n2262_), .B(\shift[6] ), .ZN(new_n3046_));
  NAND2_X1   g2670(.A1(new_n3045_), .A2(new_n3046_), .ZN(\result[86] ));
  OAI21_X1   g2671(.A1(new_n2288_), .A2(new_n2293_), .B(new_n264_), .ZN(new_n3048_));
  OAI21_X1   g2672(.A1(new_n2276_), .A2(new_n2281_), .B(\shift[6] ), .ZN(new_n3049_));
  NAND2_X1   g2673(.A1(new_n3049_), .A2(new_n3048_), .ZN(\result[87] ));
  OAI21_X1   g2674(.A1(new_n2318_), .A2(new_n2313_), .B(new_n264_), .ZN(new_n3051_));
  OAI21_X1   g2675(.A1(new_n2300_), .A2(new_n2306_), .B(\shift[6] ), .ZN(new_n3052_));
  NAND2_X1   g2676(.A1(new_n3051_), .A2(new_n3052_), .ZN(\result[88] ));
  OAI21_X1   g2677(.A1(new_n2332_), .A2(new_n2336_), .B(new_n264_), .ZN(new_n3054_));
  OAI21_X1   g2678(.A1(new_n2323_), .A2(new_n2328_), .B(\shift[6] ), .ZN(new_n3055_));
  NAND2_X1   g2679(.A1(new_n3055_), .A2(new_n3054_), .ZN(\result[89] ));
  OAI21_X1   g2680(.A1(new_n2357_), .A2(new_n2352_), .B(new_n264_), .ZN(new_n3057_));
  OAI21_X1   g2681(.A1(new_n2344_), .A2(new_n2346_), .B(\shift[6] ), .ZN(new_n3058_));
  NAND2_X1   g2682(.A1(new_n3057_), .A2(new_n3058_), .ZN(\result[90] ));
  OAI21_X1   g2683(.A1(new_n2369_), .A2(new_n2374_), .B(new_n264_), .ZN(new_n3060_));
  OAI21_X1   g2684(.A1(new_n2363_), .A2(new_n2361_), .B(\shift[6] ), .ZN(new_n3061_));
  NAND2_X1   g2685(.A1(new_n3061_), .A2(new_n3060_), .ZN(\result[91] ));
  OAI21_X1   g2686(.A1(new_n2392_), .A2(new_n2390_), .B(\shift[6] ), .ZN(new_n3063_));
  OAI21_X1   g2687(.A1(\shift[6] ), .A2(new_n2415_), .B(new_n3063_), .ZN(\result[92] ));
  OAI21_X1   g2688(.A1(new_n2430_), .A2(new_n2426_), .B(new_n264_), .ZN(new_n3065_));
  OAI21_X1   g2689(.A1(new_n2421_), .A2(new_n264_), .B(new_n3065_), .ZN(\result[93] ));
  OAI21_X1   g2690(.A1(new_n2448_), .A2(new_n2444_), .B(new_n264_), .ZN(new_n3067_));
  OAI21_X1   g2691(.A1(new_n2436_), .A2(new_n2438_), .B(\shift[6] ), .ZN(new_n3068_));
  NAND2_X1   g2692(.A1(new_n3067_), .A2(new_n3068_), .ZN(\result[94] ));
  OAI21_X1   g2693(.A1(new_n2458_), .A2(new_n2462_), .B(new_n264_), .ZN(new_n3070_));
  OAI21_X1   g2694(.A1(new_n2452_), .A2(new_n2454_), .B(\shift[6] ), .ZN(new_n3071_));
  NAND2_X1   g2695(.A1(new_n3070_), .A2(new_n3071_), .ZN(\result[95] ));
  OAI21_X1   g2696(.A1(new_n2479_), .A2(new_n2475_), .B(new_n264_), .ZN(new_n3073_));
  OAI21_X1   g2697(.A1(new_n2467_), .A2(new_n2471_), .B(\shift[6] ), .ZN(new_n3074_));
  NAND2_X1   g2698(.A1(new_n3073_), .A2(new_n3074_), .ZN(\result[96] ));
  OAI21_X1   g2699(.A1(new_n2491_), .A2(new_n2495_), .B(new_n264_), .ZN(new_n3076_));
  OAI21_X1   g2700(.A1(new_n2487_), .A2(new_n2483_), .B(\shift[6] ), .ZN(new_n3077_));
  NAND2_X1   g2701(.A1(new_n3077_), .A2(new_n3076_), .ZN(\result[97] ));
  OAI21_X1   g2702(.A1(new_n2514_), .A2(new_n2510_), .B(new_n264_), .ZN(new_n3079_));
  OAI21_X1   g2703(.A1(new_n2500_), .A2(new_n2504_), .B(\shift[6] ), .ZN(new_n3080_));
  NAND2_X1   g2704(.A1(new_n3079_), .A2(new_n3080_), .ZN(\result[98] ));
  OAI21_X1   g2705(.A1(new_n2524_), .A2(new_n2526_), .B(new_n264_), .ZN(new_n3082_));
  OAI21_X1   g2706(.A1(new_n2522_), .A2(new_n2518_), .B(\shift[6] ), .ZN(new_n3083_));
  NAND2_X1   g2707(.A1(new_n3083_), .A2(new_n3082_), .ZN(\result[99] ));
  OAI21_X1   g2708(.A1(new_n2545_), .A2(new_n2541_), .B(new_n264_), .ZN(new_n3085_));
  OAI21_X1   g2709(.A1(new_n2537_), .A2(new_n2531_), .B(\shift[6] ), .ZN(new_n3086_));
  NAND2_X1   g2710(.A1(new_n3086_), .A2(new_n3085_), .ZN(\result[100] ));
  OAI21_X1   g2711(.A1(new_n2558_), .A2(new_n2562_), .B(new_n264_), .ZN(new_n3088_));
  OAI21_X1   g2712(.A1(new_n2550_), .A2(new_n2553_), .B(\shift[6] ), .ZN(new_n3089_));
  NAND2_X1   g2713(.A1(new_n3089_), .A2(new_n3088_), .ZN(\result[101] ));
  OAI21_X1   g2714(.A1(new_n2578_), .A2(new_n2574_), .B(new_n264_), .ZN(new_n3091_));
  OAI21_X1   g2715(.A1(new_n2566_), .A2(new_n2569_), .B(\shift[6] ), .ZN(new_n3092_));
  NAND2_X1   g2716(.A1(new_n3092_), .A2(new_n3091_), .ZN(\result[102] ));
  OAI21_X1   g2717(.A1(new_n2590_), .A2(new_n2594_), .B(new_n264_), .ZN(new_n3094_));
  OAI21_X1   g2718(.A1(new_n2583_), .A2(new_n2587_), .B(\shift[6] ), .ZN(new_n3095_));
  NAND2_X1   g2719(.A1(new_n3094_), .A2(new_n3095_), .ZN(\result[103] ));
  OAI21_X1   g2720(.A1(new_n2607_), .A2(new_n2611_), .B(new_n264_), .ZN(new_n3097_));
  OAI21_X1   g2721(.A1(new_n2599_), .A2(new_n2603_), .B(\shift[6] ), .ZN(new_n3098_));
  NAND2_X1   g2722(.A1(new_n3098_), .A2(new_n3097_), .ZN(\result[104] ));
  OAI21_X1   g2723(.A1(new_n2623_), .A2(new_n2627_), .B(new_n264_), .ZN(new_n3100_));
  OAI21_X1   g2724(.A1(new_n2620_), .A2(new_n2616_), .B(\shift[6] ), .ZN(new_n3101_));
  NAND2_X1   g2725(.A1(new_n3101_), .A2(new_n3100_), .ZN(\result[105] ));
  OAI21_X1   g2726(.A1(new_n2643_), .A2(new_n2638_), .B(new_n264_), .ZN(new_n3103_));
  OAI21_X1   g2727(.A1(new_n2631_), .A2(new_n2634_), .B(\shift[6] ), .ZN(new_n3104_));
  NAND2_X1   g2728(.A1(new_n3104_), .A2(new_n3103_), .ZN(\result[106] ));
  OAI21_X1   g2729(.A1(new_n2653_), .A2(new_n2657_), .B(new_n264_), .ZN(new_n3106_));
  OAI21_X1   g2730(.A1(new_n2650_), .A2(new_n2647_), .B(\shift[6] ), .ZN(new_n3107_));
  NAND2_X1   g2731(.A1(new_n3107_), .A2(new_n3106_), .ZN(\result[107] ));
  OAI21_X1   g2732(.A1(new_n2673_), .A2(new_n2669_), .B(new_n264_), .ZN(new_n3109_));
  OAI21_X1   g2733(.A1(new_n2665_), .A2(new_n2662_), .B(\shift[6] ), .ZN(new_n3110_));
  NAND2_X1   g2734(.A1(new_n3110_), .A2(new_n3109_), .ZN(\result[108] ));
  OAI21_X1   g2735(.A1(new_n2684_), .A2(new_n2689_), .B(new_n264_), .ZN(new_n3112_));
  OAI21_X1   g2736(.A1(new_n2681_), .A2(new_n2678_), .B(\shift[6] ), .ZN(new_n3113_));
  NAND2_X1   g2737(.A1(new_n3113_), .A2(new_n3112_), .ZN(\result[109] ));
  OAI21_X1   g2738(.A1(new_n2705_), .A2(new_n2701_), .B(new_n264_), .ZN(new_n3115_));
  OAI21_X1   g2739(.A1(new_n2694_), .A2(new_n2697_), .B(\shift[6] ), .ZN(new_n3116_));
  NAND2_X1   g2740(.A1(new_n3115_), .A2(new_n3116_), .ZN(\result[110] ));
  OAI21_X1   g2741(.A1(new_n2716_), .A2(new_n2721_), .B(new_n264_), .ZN(new_n3118_));
  OAI21_X1   g2742(.A1(new_n2713_), .A2(new_n2710_), .B(\shift[6] ), .ZN(new_n3119_));
  NAND2_X1   g2743(.A1(new_n3118_), .A2(new_n3119_), .ZN(\result[111] ));
  OAI21_X1   g2744(.A1(new_n2728_), .A2(new_n2726_), .B(\shift[6] ), .ZN(new_n3121_));
  OAI21_X1   g2745(.A1(new_n2744_), .A2(\shift[6] ), .B(new_n3121_), .ZN(\result[112] ));
  OAI21_X1   g2746(.A1(new_n2753_), .A2(new_n2755_), .B(new_n264_), .ZN(new_n3123_));
  OAI21_X1   g2747(.A1(new_n2750_), .A2(new_n2748_), .B(\shift[6] ), .ZN(new_n3124_));
  NAND2_X1   g2748(.A1(new_n3124_), .A2(new_n3123_), .ZN(\result[113] ));
  OAI21_X1   g2749(.A1(new_n2768_), .A2(new_n2766_), .B(new_n264_), .ZN(new_n3126_));
  OAI21_X1   g2750(.A1(new_n2760_), .A2(new_n2762_), .B(\shift[6] ), .ZN(new_n3127_));
  NAND2_X1   g2751(.A1(new_n3126_), .A2(new_n3127_), .ZN(\result[114] ));
  OAI21_X1   g2752(.A1(new_n2780_), .A2(new_n2782_), .B(new_n264_), .ZN(new_n3129_));
  OAI21_X1   g2753(.A1(new_n2773_), .A2(new_n2777_), .B(\shift[6] ), .ZN(new_n3130_));
  NAND2_X1   g2754(.A1(new_n3129_), .A2(new_n3130_), .ZN(\result[115] ));
  OAI21_X1   g2755(.A1(new_n2799_), .A2(new_n2804_), .B(new_n264_), .ZN(new_n3132_));
  OAI21_X1   g2756(.A1(new_n2788_), .A2(new_n2794_), .B(\shift[6] ), .ZN(new_n3133_));
  NAND2_X1   g2757(.A1(new_n3133_), .A2(new_n3132_), .ZN(\result[116] ));
  OAI21_X1   g2758(.A1(new_n2818_), .A2(new_n2821_), .B(new_n264_), .ZN(new_n3135_));
  OAI21_X1   g2759(.A1(new_n2810_), .A2(new_n2814_), .B(\shift[6] ), .ZN(new_n3136_));
  NAND2_X1   g2760(.A1(new_n3136_), .A2(new_n3135_), .ZN(\result[117] ));
  OAI21_X1   g2761(.A1(new_n2838_), .A2(new_n2843_), .B(new_n264_), .ZN(new_n3138_));
  OAI21_X1   g2762(.A1(new_n2827_), .A2(new_n2833_), .B(\shift[6] ), .ZN(new_n3139_));
  NAND2_X1   g2763(.A1(new_n3138_), .A2(new_n3139_), .ZN(\result[118] ));
  OAI21_X1   g2764(.A1(new_n2851_), .A2(new_n2853_), .B(new_n264_), .ZN(new_n3141_));
  OAI21_X1   g2765(.A1(new_n2848_), .A2(new_n2846_), .B(\shift[6] ), .ZN(new_n3142_));
  NAND2_X1   g2766(.A1(new_n3142_), .A2(new_n3141_), .ZN(\result[119] ));
  OAI21_X1   g2767(.A1(new_n2865_), .A2(new_n2863_), .B(new_n264_), .ZN(new_n3144_));
  OAI21_X1   g2768(.A1(new_n2858_), .A2(new_n2856_), .B(\shift[6] ), .ZN(new_n3145_));
  NAND2_X1   g2769(.A1(new_n3144_), .A2(new_n3145_), .ZN(\result[120] ));
  OAI21_X1   g2770(.A1(new_n2873_), .A2(new_n2875_), .B(new_n264_), .ZN(new_n3147_));
  OAI21_X1   g2771(.A1(new_n2870_), .A2(new_n2868_), .B(\shift[6] ), .ZN(new_n3148_));
  NAND2_X1   g2772(.A1(new_n3148_), .A2(new_n3147_), .ZN(\result[121] ));
  OAI21_X1   g2773(.A1(new_n2892_), .A2(new_n2890_), .B(new_n264_), .ZN(new_n3150_));
  OAI21_X1   g2774(.A1(new_n2881_), .A2(new_n2886_), .B(\shift[6] ), .ZN(new_n3151_));
  NAND2_X1   g2775(.A1(new_n3151_), .A2(new_n3150_), .ZN(\result[122] ));
  OAI21_X1   g2776(.A1(new_n2906_), .A2(new_n2908_), .B(new_n264_), .ZN(new_n3153_));
  OAI21_X1   g2777(.A1(new_n2900_), .A2(new_n2903_), .B(\shift[6] ), .ZN(new_n3154_));
  NAND2_X1   g2778(.A1(new_n3154_), .A2(new_n3153_), .ZN(\result[123] ));
  OAI21_X1   g2779(.A1(new_n2928_), .A2(new_n2926_), .B(new_n264_), .ZN(new_n3156_));
  OAI21_X1   g2780(.A1(new_n2923_), .A2(new_n264_), .B(new_n3156_), .ZN(\result[124] ));
  OAI21_X1   g2781(.A1(new_n2941_), .A2(new_n2943_), .B(new_n264_), .ZN(new_n3158_));
  OAI21_X1   g2782(.A1(new_n2938_), .A2(new_n2934_), .B(\shift[6] ), .ZN(new_n3159_));
  NAND2_X1   g2783(.A1(new_n3159_), .A2(new_n3158_), .ZN(\result[125] ));
  OAI21_X1   g2784(.A1(new_n2958_), .A2(new_n2960_), .B(new_n264_), .ZN(new_n3161_));
  OAI21_X1   g2785(.A1(new_n2949_), .A2(new_n2954_), .B(\shift[6] ), .ZN(new_n3162_));
  NAND2_X1   g2786(.A1(new_n3162_), .A2(new_n3161_), .ZN(\result[126] ));
  OAI21_X1   g2787(.A1(new_n2974_), .A2(new_n2976_), .B(new_n264_), .ZN(new_n3164_));
  OAI21_X1   g2788(.A1(new_n2971_), .A2(new_n2966_), .B(\shift[6] ), .ZN(new_n3165_));
  NAND2_X1   g2789(.A1(new_n3165_), .A2(new_n3164_), .ZN(\result[127] ));
endmodule


