// Benchmark "adder" written by ABC on Thu Sep 14 18:32:01 2023

module adder ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n387_, new_n388_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1712_, new_n1713_;
  XOR2_X1    g0000(.A1(\a[0] ), .A2(\b[0] ), .Z(\f[0] ));
  NAND2_X1   g0001(.A1(\a[1] ), .A2(\b[1] ), .ZN(new_n387_));
  XNOR2_X1   g0002(.A1(new_n387_), .A2(\a[0] ), .ZN(new_n388_));
  XOR2_X1    g0003(.A1(new_n388_), .A2(\b[0] ), .Z(\f[1] ));
  AND2_X2    g0004(.A1(\a[1] ), .A2(\b[1] ), .Z(new_n390_));
  NOR2_X1    g0005(.A1(\a[1] ), .A2(\b[1] ), .ZN(new_n391_));
  INV_X1     g0006(.I(new_n391_), .ZN(new_n392_));
  AND2_X2    g0007(.A1(\a[0] ), .A2(\b[0] ), .Z(new_n393_));
  AOI21_X1   g0008(.A1(new_n392_), .A2(new_n393_), .B(new_n390_), .ZN(new_n394_));
  XNOR2_X1   g0009(.A1(\a[2] ), .A2(\b[2] ), .ZN(new_n395_));
  INV_X1     g0010(.I(\a[2] ), .ZN(new_n396_));
  INV_X1     g0011(.I(\b[2] ), .ZN(new_n397_));
  NOR2_X1    g0012(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1    g0013(.A1(\a[2] ), .A2(\b[2] ), .ZN(new_n399_));
  OAI21_X1   g0014(.A1(new_n398_), .A2(new_n399_), .B(new_n394_), .ZN(new_n400_));
  OAI21_X1   g0015(.A1(new_n394_), .A2(new_n395_), .B(new_n400_), .ZN(\f[2] ));
  NOR2_X1    g0016(.A1(new_n394_), .A2(new_n398_), .ZN(new_n402_));
  NOR2_X1    g0017(.A1(new_n402_), .A2(new_n399_), .ZN(new_n403_));
  XNOR2_X1   g0018(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n404_));
  NAND2_X1   g0019(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n405_));
  OR2_X2     g0020(.A1(\a[3] ), .A2(\b[3] ), .Z(new_n406_));
  NAND2_X1   g0021(.A1(new_n406_), .A2(new_n405_), .ZN(new_n407_));
  NAND2_X1   g0022(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1   g0023(.A1(new_n403_), .A2(new_n404_), .B(new_n408_), .ZN(\f[3] ));
  NAND2_X1   g0024(.A1(\a[0] ), .A2(\b[0] ), .ZN(new_n410_));
  OAI21_X1   g0025(.A1(new_n391_), .A2(new_n410_), .B(new_n387_), .ZN(new_n411_));
  OAI21_X1   g0026(.A1(new_n406_), .A2(new_n397_), .B(new_n396_), .ZN(new_n412_));
  OAI21_X1   g0027(.A1(\a[3] ), .A2(\b[3] ), .B(new_n397_), .ZN(new_n413_));
  NAND3_X1   g0028(.A1(new_n412_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1   g0029(.A1(\a[4] ), .A2(\b[4] ), .ZN(new_n415_));
  INV_X1     g0030(.I(new_n415_), .ZN(new_n416_));
  XOR2_X1    g0031(.A1(new_n414_), .A2(new_n416_), .Z(new_n417_));
  XOR2_X1    g0032(.A1(new_n417_), .A2(new_n405_), .Z(\f[4] ));
  NOR2_X1    g0033(.A1(\a[4] ), .A2(\b[4] ), .ZN(new_n419_));
  OR2_X2     g0034(.A1(new_n419_), .A2(new_n405_), .Z(new_n420_));
  OAI21_X1   g0035(.A1(new_n414_), .A2(new_n420_), .B(new_n415_), .ZN(new_n421_));
  XOR2_X1    g0036(.A1(\a[5] ), .A2(\b[5] ), .Z(new_n422_));
  NAND2_X1   g0037(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XOR2_X1    g0038(.A1(\a[5] ), .A2(\b[5] ), .Z(new_n424_));
  OAI21_X1   g0039(.A1(new_n421_), .A2(new_n424_), .B(new_n423_), .ZN(\f[5] ));
  NAND2_X1   g0040(.A1(\a[5] ), .A2(\b[5] ), .ZN(new_n426_));
  NOR2_X1    g0041(.A1(\a[5] ), .A2(\b[5] ), .ZN(new_n427_));
  AOI21_X1   g0042(.A1(new_n421_), .A2(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1   g0043(.A1(\a[6] ), .A2(\b[6] ), .ZN(new_n429_));
  INV_X1     g0044(.I(\a[6] ), .ZN(new_n430_));
  INV_X1     g0045(.I(\b[6] ), .ZN(new_n431_));
  NOR2_X1    g0046(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1    g0047(.A1(\a[6] ), .A2(\b[6] ), .ZN(new_n433_));
  OAI21_X1   g0048(.A1(new_n432_), .A2(new_n433_), .B(new_n428_), .ZN(new_n434_));
  OAI21_X1   g0049(.A1(new_n428_), .A2(new_n429_), .B(new_n434_), .ZN(\f[6] ));
  NOR2_X1    g0050(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n436_));
  AOI21_X1   g0051(.A1(new_n436_), .A2(\b[2] ), .B(\a[2] ), .ZN(new_n437_));
  NOR2_X1    g0052(.A1(new_n436_), .A2(\b[2] ), .ZN(new_n438_));
  NOR4_X1    g0053(.A1(new_n394_), .A2(new_n437_), .A3(new_n420_), .A4(new_n438_), .ZN(new_n439_));
  NOR2_X1    g0054(.A1(new_n433_), .A2(\b[5] ), .ZN(new_n440_));
  AOI21_X1   g0055(.A1(new_n433_), .A2(\b[5] ), .B(\a[5] ), .ZN(new_n441_));
  NOR2_X1    g0056(.A1(new_n441_), .A2(new_n440_), .ZN(new_n442_));
  OAI21_X1   g0057(.A1(new_n439_), .A2(new_n416_), .B(new_n442_), .ZN(new_n443_));
  NAND2_X1   g0058(.A1(\a[7] ), .A2(\b[7] ), .ZN(new_n444_));
  XOR2_X1    g0059(.A1(new_n443_), .A2(new_n444_), .Z(new_n445_));
  XOR2_X1    g0060(.A1(new_n445_), .A2(new_n432_), .Z(\f[7] ));
  INV_X1     g0061(.I(new_n432_), .ZN(new_n447_));
  NOR2_X1    g0062(.A1(\a[7] ), .A2(\b[7] ), .ZN(new_n448_));
  NOR2_X1    g0063(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1     g0064(.I(new_n449_), .ZN(new_n450_));
  OAI21_X1   g0065(.A1(new_n443_), .A2(new_n450_), .B(new_n444_), .ZN(new_n451_));
  XOR2_X1    g0066(.A1(\a[8] ), .A2(\b[8] ), .Z(new_n452_));
  NAND2_X1   g0067(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1    g0068(.A1(\a[8] ), .A2(\b[8] ), .Z(new_n454_));
  OAI21_X1   g0069(.A1(new_n451_), .A2(new_n454_), .B(new_n453_), .ZN(\f[8] ));
  NAND2_X1   g0070(.A1(\a[8] ), .A2(\b[8] ), .ZN(new_n456_));
  NOR2_X1    g0071(.A1(\a[8] ), .A2(\b[8] ), .ZN(new_n457_));
  AOI21_X1   g0072(.A1(new_n451_), .A2(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1   g0073(.A1(\a[9] ), .A2(\b[9] ), .ZN(new_n459_));
  NAND2_X1   g0074(.A1(\a[9] ), .A2(\b[9] ), .ZN(new_n460_));
  OR2_X2     g0075(.A1(\a[9] ), .A2(\b[9] ), .Z(new_n461_));
  NAND2_X1   g0076(.A1(new_n461_), .A2(new_n460_), .ZN(new_n462_));
  NAND2_X1   g0077(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1   g0078(.A1(new_n458_), .A2(new_n459_), .B(new_n463_), .ZN(\f[9] ));
  NAND3_X1   g0079(.A1(new_n421_), .A2(new_n442_), .A3(new_n449_), .ZN(new_n465_));
  INV_X1     g0080(.I(\b[8] ), .ZN(new_n466_));
  NOR2_X1    g0081(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  NOR2_X1    g0082(.A1(new_n467_), .A2(\a[8] ), .ZN(new_n468_));
  AOI21_X1   g0083(.A1(new_n466_), .A2(new_n461_), .B(new_n468_), .ZN(new_n469_));
  INV_X1     g0084(.I(new_n469_), .ZN(new_n470_));
  AOI21_X1   g0085(.A1(new_n465_), .A2(new_n444_), .B(new_n470_), .ZN(new_n471_));
  INV_X1     g0086(.I(\a[10] ), .ZN(new_n472_));
  INV_X1     g0087(.I(\b[10] ), .ZN(new_n473_));
  NOR2_X1    g0088(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1     g0089(.I(new_n474_), .ZN(new_n475_));
  XOR2_X1    g0090(.A1(new_n471_), .A2(new_n475_), .Z(new_n476_));
  XOR2_X1    g0091(.A1(new_n476_), .A2(new_n460_), .Z(\f[10] ));
  AOI21_X1   g0092(.A1(new_n472_), .A2(new_n473_), .B(new_n460_), .ZN(new_n478_));
  AOI21_X1   g0093(.A1(new_n471_), .A2(new_n478_), .B(new_n474_), .ZN(new_n479_));
  XNOR2_X1   g0094(.A1(\a[11] ), .A2(\b[11] ), .ZN(new_n480_));
  NAND2_X1   g0095(.A1(\a[11] ), .A2(\b[11] ), .ZN(new_n481_));
  NOR2_X1    g0096(.A1(\a[11] ), .A2(\b[11] ), .ZN(new_n482_));
  INV_X1     g0097(.I(new_n482_), .ZN(new_n483_));
  NAND2_X1   g0098(.A1(new_n483_), .A2(new_n481_), .ZN(new_n484_));
  NAND2_X1   g0099(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1   g0100(.A1(new_n479_), .A2(new_n480_), .B(new_n485_), .ZN(\f[11] ));
  INV_X1     g0101(.I(new_n479_), .ZN(new_n487_));
  AOI21_X1   g0102(.A1(new_n487_), .A2(new_n481_), .B(new_n482_), .ZN(new_n488_));
  XNOR2_X1   g0103(.A1(\a[12] ), .A2(\b[12] ), .ZN(new_n489_));
  AND2_X2    g0104(.A1(\a[12] ), .A2(\b[12] ), .Z(new_n490_));
  NOR2_X1    g0105(.A1(\a[12] ), .A2(\b[12] ), .ZN(new_n491_));
  OAI21_X1   g0106(.A1(new_n490_), .A2(new_n491_), .B(new_n488_), .ZN(new_n492_));
  OAI21_X1   g0107(.A1(new_n488_), .A2(new_n489_), .B(new_n492_), .ZN(\f[12] ));
  NAND3_X1   g0108(.A1(new_n451_), .A2(new_n469_), .A3(new_n478_), .ZN(new_n494_));
  INV_X1     g0109(.I(\b[11] ), .ZN(new_n495_));
  INV_X1     g0110(.I(new_n491_), .ZN(new_n496_));
  NAND2_X1   g0111(.A1(new_n496_), .A2(new_n495_), .ZN(new_n497_));
  NOR2_X1    g0112(.A1(new_n496_), .A2(new_n495_), .ZN(new_n498_));
  OAI21_X1   g0113(.A1(\a[11] ), .A2(new_n498_), .B(new_n497_), .ZN(new_n499_));
  AOI21_X1   g0114(.A1(new_n494_), .A2(new_n475_), .B(new_n499_), .ZN(new_n500_));
  INV_X1     g0115(.I(\a[13] ), .ZN(new_n501_));
  INV_X1     g0116(.I(\b[13] ), .ZN(new_n502_));
  NOR2_X1    g0117(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1    g0118(.A1(new_n500_), .A2(new_n503_), .Z(new_n504_));
  XOR2_X1    g0119(.A1(new_n504_), .A2(new_n490_), .Z(\f[13] ));
  INV_X1     g0120(.I(new_n490_), .ZN(new_n506_));
  AOI21_X1   g0121(.A1(new_n501_), .A2(new_n502_), .B(new_n506_), .ZN(new_n507_));
  AOI21_X1   g0122(.A1(new_n500_), .A2(new_n507_), .B(new_n503_), .ZN(new_n508_));
  XNOR2_X1   g0123(.A1(\a[14] ), .A2(\b[14] ), .ZN(new_n509_));
  NAND2_X1   g0124(.A1(\a[14] ), .A2(\b[14] ), .ZN(new_n510_));
  NOR2_X1    g0125(.A1(\a[14] ), .A2(\b[14] ), .ZN(new_n511_));
  INV_X1     g0126(.I(new_n511_), .ZN(new_n512_));
  NAND2_X1   g0127(.A1(new_n512_), .A2(new_n510_), .ZN(new_n513_));
  NAND2_X1   g0128(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1   g0129(.A1(new_n508_), .A2(new_n509_), .B(new_n514_), .ZN(\f[14] ));
  INV_X1     g0130(.I(new_n508_), .ZN(new_n516_));
  AOI21_X1   g0131(.A1(new_n516_), .A2(new_n510_), .B(new_n511_), .ZN(new_n517_));
  XNOR2_X1   g0132(.A1(\a[15] ), .A2(\b[15] ), .ZN(new_n518_));
  AND2_X2    g0133(.A1(\a[15] ), .A2(\b[15] ), .Z(new_n519_));
  NOR2_X1    g0134(.A1(\a[15] ), .A2(\b[15] ), .ZN(new_n520_));
  OAI21_X1   g0135(.A1(new_n519_), .A2(new_n520_), .B(new_n517_), .ZN(new_n521_));
  OAI21_X1   g0136(.A1(new_n517_), .A2(new_n518_), .B(new_n521_), .ZN(\f[15] ));
  INV_X1     g0137(.I(new_n519_), .ZN(new_n523_));
  INV_X1     g0138(.I(new_n507_), .ZN(new_n524_));
  NOR3_X1    g0139(.A1(new_n479_), .A2(new_n499_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1     g0140(.I(\b[14] ), .ZN(new_n526_));
  INV_X1     g0141(.I(new_n520_), .ZN(new_n527_));
  AOI21_X1   g0142(.A1(new_n520_), .A2(\b[14] ), .B(\a[14] ), .ZN(new_n528_));
  AOI21_X1   g0143(.A1(new_n526_), .A2(new_n527_), .B(new_n528_), .ZN(new_n529_));
  OAI21_X1   g0144(.A1(new_n525_), .A2(new_n503_), .B(new_n529_), .ZN(new_n530_));
  INV_X1     g0145(.I(\a[16] ), .ZN(new_n531_));
  INV_X1     g0146(.I(\b[16] ), .ZN(new_n532_));
  NOR2_X1    g0147(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1    g0148(.A1(new_n530_), .A2(new_n533_), .Z(new_n534_));
  XOR2_X1    g0149(.A1(new_n534_), .A2(new_n523_), .Z(\f[16] ));
  INV_X1     g0150(.I(new_n533_), .ZN(new_n536_));
  AOI21_X1   g0151(.A1(new_n531_), .A2(new_n532_), .B(new_n523_), .ZN(new_n537_));
  INV_X1     g0152(.I(new_n537_), .ZN(new_n538_));
  OAI21_X1   g0153(.A1(new_n530_), .A2(new_n538_), .B(new_n536_), .ZN(new_n539_));
  INV_X1     g0154(.I(new_n539_), .ZN(new_n540_));
  XNOR2_X1   g0155(.A1(\a[17] ), .A2(\b[17] ), .ZN(new_n541_));
  INV_X1     g0156(.I(\a[17] ), .ZN(new_n542_));
  INV_X1     g0157(.I(\b[17] ), .ZN(new_n543_));
  NOR2_X1    g0158(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1    g0159(.A1(\a[17] ), .A2(\b[17] ), .ZN(new_n545_));
  OAI21_X1   g0160(.A1(new_n544_), .A2(new_n545_), .B(new_n540_), .ZN(new_n546_));
  OAI21_X1   g0161(.A1(new_n540_), .A2(new_n541_), .B(new_n546_), .ZN(\f[17] ));
  NAND2_X1   g0162(.A1(new_n542_), .A2(new_n543_), .ZN(new_n548_));
  OAI21_X1   g0163(.A1(new_n540_), .A2(new_n544_), .B(new_n548_), .ZN(new_n549_));
  XOR2_X1    g0164(.A1(\a[18] ), .A2(\b[18] ), .Z(new_n550_));
  NAND2_X1   g0165(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1     g0166(.I(\a[18] ), .ZN(new_n552_));
  INV_X1     g0167(.I(\b[18] ), .ZN(new_n553_));
  NOR2_X1    g0168(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1    g0169(.A1(\a[18] ), .A2(\b[18] ), .ZN(new_n555_));
  NOR2_X1    g0170(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1   g0171(.A1(new_n549_), .A2(new_n556_), .B(new_n551_), .ZN(\f[18] ));
  INV_X1     g0172(.I(new_n554_), .ZN(new_n558_));
  INV_X1     g0173(.I(new_n529_), .ZN(new_n559_));
  NOR3_X1    g0174(.A1(new_n508_), .A2(new_n559_), .A3(new_n538_), .ZN(new_n560_));
  NOR2_X1    g0175(.A1(new_n555_), .A2(\b[17] ), .ZN(new_n561_));
  AOI21_X1   g0176(.A1(new_n555_), .A2(\b[17] ), .B(\a[17] ), .ZN(new_n562_));
  NOR2_X1    g0177(.A1(new_n562_), .A2(new_n561_), .ZN(new_n563_));
  OAI21_X1   g0178(.A1(new_n560_), .A2(new_n533_), .B(new_n563_), .ZN(new_n564_));
  INV_X1     g0179(.I(\a[19] ), .ZN(new_n565_));
  INV_X1     g0180(.I(\b[19] ), .ZN(new_n566_));
  NOR2_X1    g0181(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1    g0182(.A1(new_n564_), .A2(new_n567_), .Z(new_n568_));
  XOR2_X1    g0183(.A1(new_n568_), .A2(new_n558_), .Z(\f[19] ));
  INV_X1     g0184(.I(new_n567_), .ZN(new_n570_));
  AOI21_X1   g0185(.A1(new_n565_), .A2(new_n566_), .B(new_n558_), .ZN(new_n571_));
  INV_X1     g0186(.I(new_n571_), .ZN(new_n572_));
  OAI21_X1   g0187(.A1(new_n564_), .A2(new_n572_), .B(new_n570_), .ZN(new_n573_));
  INV_X1     g0188(.I(new_n573_), .ZN(new_n574_));
  XNOR2_X1   g0189(.A1(\a[20] ), .A2(\b[20] ), .ZN(new_n575_));
  INV_X1     g0190(.I(\a[20] ), .ZN(new_n576_));
  INV_X1     g0191(.I(\b[20] ), .ZN(new_n577_));
  NOR2_X1    g0192(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1    g0193(.A1(\a[20] ), .A2(\b[20] ), .ZN(new_n579_));
  OAI21_X1   g0194(.A1(new_n578_), .A2(new_n579_), .B(new_n574_), .ZN(new_n580_));
  OAI21_X1   g0195(.A1(new_n574_), .A2(new_n575_), .B(new_n580_), .ZN(\f[20] ));
  NAND2_X1   g0196(.A1(new_n576_), .A2(new_n577_), .ZN(new_n582_));
  OAI21_X1   g0197(.A1(new_n574_), .A2(new_n578_), .B(new_n582_), .ZN(new_n583_));
  XOR2_X1    g0198(.A1(\a[21] ), .A2(\b[21] ), .Z(new_n584_));
  NAND2_X1   g0199(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1     g0200(.I(\a[21] ), .ZN(new_n586_));
  INV_X1     g0201(.I(\b[21] ), .ZN(new_n587_));
  NOR2_X1    g0202(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1    g0203(.A1(\a[21] ), .A2(\b[21] ), .ZN(new_n589_));
  NOR2_X1    g0204(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1   g0205(.A1(new_n583_), .A2(new_n590_), .B(new_n585_), .ZN(\f[21] ));
  INV_X1     g0206(.I(new_n588_), .ZN(new_n592_));
  NAND3_X1   g0207(.A1(new_n539_), .A2(new_n563_), .A3(new_n571_), .ZN(new_n593_));
  INV_X1     g0208(.I(new_n589_), .ZN(new_n594_));
  AOI21_X1   g0209(.A1(new_n589_), .A2(\b[20] ), .B(\a[20] ), .ZN(new_n595_));
  AOI21_X1   g0210(.A1(new_n577_), .A2(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1     g0211(.I(new_n596_), .ZN(new_n597_));
  AOI21_X1   g0212(.A1(new_n593_), .A2(new_n570_), .B(new_n597_), .ZN(new_n598_));
  INV_X1     g0213(.I(\a[22] ), .ZN(new_n599_));
  INV_X1     g0214(.I(\b[22] ), .ZN(new_n600_));
  NOR2_X1    g0215(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1     g0216(.I(new_n601_), .ZN(new_n602_));
  XOR2_X1    g0217(.A1(new_n598_), .A2(new_n602_), .Z(new_n603_));
  XOR2_X1    g0218(.A1(new_n603_), .A2(new_n592_), .Z(\f[22] ));
  AOI21_X1   g0219(.A1(new_n599_), .A2(new_n600_), .B(new_n592_), .ZN(new_n605_));
  AOI21_X1   g0220(.A1(new_n598_), .A2(new_n605_), .B(new_n601_), .ZN(new_n606_));
  XNOR2_X1   g0221(.A1(\a[23] ), .A2(\b[23] ), .ZN(new_n607_));
  NAND2_X1   g0222(.A1(\a[23] ), .A2(\b[23] ), .ZN(new_n608_));
  NOR2_X1    g0223(.A1(\a[23] ), .A2(\b[23] ), .ZN(new_n609_));
  INV_X1     g0224(.I(new_n609_), .ZN(new_n610_));
  NAND2_X1   g0225(.A1(new_n610_), .A2(new_n608_), .ZN(new_n611_));
  NAND2_X1   g0226(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1   g0227(.A1(new_n606_), .A2(new_n607_), .B(new_n612_), .ZN(\f[23] ));
  INV_X1     g0228(.I(new_n606_), .ZN(new_n614_));
  AOI21_X1   g0229(.A1(new_n614_), .A2(new_n608_), .B(new_n609_), .ZN(new_n615_));
  XNOR2_X1   g0230(.A1(\a[24] ), .A2(\b[24] ), .ZN(new_n616_));
  AND2_X2    g0231(.A1(\a[24] ), .A2(\b[24] ), .Z(new_n617_));
  NOR2_X1    g0232(.A1(\a[24] ), .A2(\b[24] ), .ZN(new_n618_));
  OAI21_X1   g0233(.A1(new_n617_), .A2(new_n618_), .B(new_n615_), .ZN(new_n619_));
  OAI21_X1   g0234(.A1(new_n615_), .A2(new_n616_), .B(new_n619_), .ZN(\f[24] ));
  NAND3_X1   g0235(.A1(new_n573_), .A2(new_n596_), .A3(new_n605_), .ZN(new_n621_));
  NOR2_X1    g0236(.A1(new_n618_), .A2(\b[23] ), .ZN(new_n622_));
  AOI21_X1   g0237(.A1(new_n618_), .A2(\b[23] ), .B(\a[23] ), .ZN(new_n623_));
  NOR2_X1    g0238(.A1(new_n623_), .A2(new_n622_), .ZN(new_n624_));
  INV_X1     g0239(.I(new_n624_), .ZN(new_n625_));
  AOI21_X1   g0240(.A1(new_n621_), .A2(new_n602_), .B(new_n625_), .ZN(new_n626_));
  INV_X1     g0241(.I(\a[25] ), .ZN(new_n627_));
  INV_X1     g0242(.I(\b[25] ), .ZN(new_n628_));
  NOR2_X1    g0243(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1    g0244(.A1(new_n626_), .A2(new_n629_), .Z(new_n630_));
  XOR2_X1    g0245(.A1(new_n630_), .A2(new_n617_), .Z(\f[25] ));
  INV_X1     g0246(.I(new_n617_), .ZN(new_n632_));
  AOI21_X1   g0247(.A1(new_n627_), .A2(new_n628_), .B(new_n632_), .ZN(new_n633_));
  AOI21_X1   g0248(.A1(new_n626_), .A2(new_n633_), .B(new_n629_), .ZN(new_n634_));
  XNOR2_X1   g0249(.A1(\a[26] ), .A2(\b[26] ), .ZN(new_n635_));
  NAND2_X1   g0250(.A1(\a[26] ), .A2(\b[26] ), .ZN(new_n636_));
  NOR2_X1    g0251(.A1(\a[26] ), .A2(\b[26] ), .ZN(new_n637_));
  INV_X1     g0252(.I(new_n637_), .ZN(new_n638_));
  NAND2_X1   g0253(.A1(new_n638_), .A2(new_n636_), .ZN(new_n639_));
  NAND2_X1   g0254(.A1(new_n634_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1   g0255(.A1(new_n634_), .A2(new_n635_), .B(new_n640_), .ZN(\f[26] ));
  INV_X1     g0256(.I(new_n634_), .ZN(new_n642_));
  AOI21_X1   g0257(.A1(new_n642_), .A2(new_n636_), .B(new_n637_), .ZN(new_n643_));
  XNOR2_X1   g0258(.A1(\a[27] ), .A2(\b[27] ), .ZN(new_n644_));
  AND2_X2    g0259(.A1(\a[27] ), .A2(\b[27] ), .Z(new_n645_));
  NOR2_X1    g0260(.A1(\a[27] ), .A2(\b[27] ), .ZN(new_n646_));
  OAI21_X1   g0261(.A1(new_n645_), .A2(new_n646_), .B(new_n643_), .ZN(new_n647_));
  OAI21_X1   g0262(.A1(new_n643_), .A2(new_n644_), .B(new_n647_), .ZN(\f[27] ));
  INV_X1     g0263(.I(new_n645_), .ZN(new_n649_));
  INV_X1     g0264(.I(new_n633_), .ZN(new_n650_));
  NOR3_X1    g0265(.A1(new_n606_), .A2(new_n625_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1     g0266(.I(\b[26] ), .ZN(new_n652_));
  INV_X1     g0267(.I(new_n646_), .ZN(new_n653_));
  AOI21_X1   g0268(.A1(new_n646_), .A2(\b[26] ), .B(\a[26] ), .ZN(new_n654_));
  AOI21_X1   g0269(.A1(new_n652_), .A2(new_n653_), .B(new_n654_), .ZN(new_n655_));
  OAI21_X1   g0270(.A1(new_n651_), .A2(new_n629_), .B(new_n655_), .ZN(new_n656_));
  INV_X1     g0271(.I(\a[28] ), .ZN(new_n657_));
  INV_X1     g0272(.I(\b[28] ), .ZN(new_n658_));
  NOR2_X1    g0273(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  XOR2_X1    g0274(.A1(new_n656_), .A2(new_n659_), .Z(new_n660_));
  XOR2_X1    g0275(.A1(new_n660_), .A2(new_n649_), .Z(\f[28] ));
  INV_X1     g0276(.I(new_n659_), .ZN(new_n662_));
  AOI21_X1   g0277(.A1(new_n657_), .A2(new_n658_), .B(new_n649_), .ZN(new_n663_));
  INV_X1     g0278(.I(new_n663_), .ZN(new_n664_));
  OAI21_X1   g0279(.A1(new_n656_), .A2(new_n664_), .B(new_n662_), .ZN(new_n665_));
  INV_X1     g0280(.I(new_n665_), .ZN(new_n666_));
  XNOR2_X1   g0281(.A1(\a[29] ), .A2(\b[29] ), .ZN(new_n667_));
  INV_X1     g0282(.I(\a[29] ), .ZN(new_n668_));
  INV_X1     g0283(.I(\b[29] ), .ZN(new_n669_));
  NOR2_X1    g0284(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1    g0285(.A1(\a[29] ), .A2(\b[29] ), .ZN(new_n671_));
  OAI21_X1   g0286(.A1(new_n670_), .A2(new_n671_), .B(new_n666_), .ZN(new_n672_));
  OAI21_X1   g0287(.A1(new_n666_), .A2(new_n667_), .B(new_n672_), .ZN(\f[29] ));
  NAND2_X1   g0288(.A1(new_n668_), .A2(new_n669_), .ZN(new_n674_));
  OAI21_X1   g0289(.A1(new_n666_), .A2(new_n670_), .B(new_n674_), .ZN(new_n675_));
  XOR2_X1    g0290(.A1(\a[30] ), .A2(\b[30] ), .Z(new_n676_));
  NAND2_X1   g0291(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1     g0292(.I(\a[30] ), .ZN(new_n678_));
  INV_X1     g0293(.I(\b[30] ), .ZN(new_n679_));
  NOR2_X1    g0294(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NOR2_X1    g0295(.A1(\a[30] ), .A2(\b[30] ), .ZN(new_n681_));
  NOR2_X1    g0296(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1   g0297(.A1(new_n675_), .A2(new_n682_), .B(new_n677_), .ZN(\f[30] ));
  INV_X1     g0298(.I(new_n680_), .ZN(new_n684_));
  INV_X1     g0299(.I(new_n655_), .ZN(new_n685_));
  NOR3_X1    g0300(.A1(new_n634_), .A2(new_n685_), .A3(new_n664_), .ZN(new_n686_));
  NOR2_X1    g0301(.A1(new_n681_), .A2(\b[29] ), .ZN(new_n687_));
  AOI21_X1   g0302(.A1(new_n681_), .A2(\b[29] ), .B(\a[29] ), .ZN(new_n688_));
  NOR2_X1    g0303(.A1(new_n688_), .A2(new_n687_), .ZN(new_n689_));
  OAI21_X1   g0304(.A1(new_n686_), .A2(new_n659_), .B(new_n689_), .ZN(new_n690_));
  INV_X1     g0305(.I(\a[31] ), .ZN(new_n691_));
  INV_X1     g0306(.I(\b[31] ), .ZN(new_n692_));
  NOR2_X1    g0307(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  XOR2_X1    g0308(.A1(new_n690_), .A2(new_n693_), .Z(new_n694_));
  XOR2_X1    g0309(.A1(new_n694_), .A2(new_n684_), .Z(\f[31] ));
  INV_X1     g0310(.I(new_n693_), .ZN(new_n696_));
  AOI21_X1   g0311(.A1(new_n691_), .A2(new_n692_), .B(new_n684_), .ZN(new_n697_));
  INV_X1     g0312(.I(new_n697_), .ZN(new_n698_));
  OAI21_X1   g0313(.A1(new_n690_), .A2(new_n698_), .B(new_n696_), .ZN(new_n699_));
  INV_X1     g0314(.I(new_n699_), .ZN(new_n700_));
  XNOR2_X1   g0315(.A1(\a[32] ), .A2(\b[32] ), .ZN(new_n701_));
  INV_X1     g0316(.I(\a[32] ), .ZN(new_n702_));
  INV_X1     g0317(.I(\b[32] ), .ZN(new_n703_));
  NOR2_X1    g0318(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1    g0319(.A1(\a[32] ), .A2(\b[32] ), .ZN(new_n705_));
  OAI21_X1   g0320(.A1(new_n704_), .A2(new_n705_), .B(new_n700_), .ZN(new_n706_));
  OAI21_X1   g0321(.A1(new_n700_), .A2(new_n701_), .B(new_n706_), .ZN(\f[32] ));
  NAND2_X1   g0322(.A1(new_n702_), .A2(new_n703_), .ZN(new_n708_));
  OAI21_X1   g0323(.A1(new_n700_), .A2(new_n704_), .B(new_n708_), .ZN(new_n709_));
  XOR2_X1    g0324(.A1(\a[33] ), .A2(\b[33] ), .Z(new_n710_));
  NAND2_X1   g0325(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1     g0326(.I(\a[33] ), .ZN(new_n712_));
  INV_X1     g0327(.I(\b[33] ), .ZN(new_n713_));
  NOR2_X1    g0328(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1    g0329(.A1(\a[33] ), .A2(\b[33] ), .ZN(new_n715_));
  NOR2_X1    g0330(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI21_X1   g0331(.A1(new_n709_), .A2(new_n716_), .B(new_n711_), .ZN(\f[33] ));
  INV_X1     g0332(.I(new_n714_), .ZN(new_n718_));
  NAND3_X1   g0333(.A1(new_n665_), .A2(new_n689_), .A3(new_n697_), .ZN(new_n719_));
  INV_X1     g0334(.I(new_n715_), .ZN(new_n720_));
  AOI21_X1   g0335(.A1(new_n715_), .A2(\b[32] ), .B(\a[32] ), .ZN(new_n721_));
  AOI21_X1   g0336(.A1(new_n703_), .A2(new_n720_), .B(new_n721_), .ZN(new_n722_));
  INV_X1     g0337(.I(new_n722_), .ZN(new_n723_));
  AOI21_X1   g0338(.A1(new_n719_), .A2(new_n696_), .B(new_n723_), .ZN(new_n724_));
  INV_X1     g0339(.I(\a[34] ), .ZN(new_n725_));
  INV_X1     g0340(.I(\b[34] ), .ZN(new_n726_));
  NOR2_X1    g0341(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1     g0342(.I(new_n727_), .ZN(new_n728_));
  XOR2_X1    g0343(.A1(new_n724_), .A2(new_n728_), .Z(new_n729_));
  XOR2_X1    g0344(.A1(new_n729_), .A2(new_n718_), .Z(\f[34] ));
  AOI21_X1   g0345(.A1(new_n725_), .A2(new_n726_), .B(new_n718_), .ZN(new_n731_));
  AOI21_X1   g0346(.A1(new_n724_), .A2(new_n731_), .B(new_n727_), .ZN(new_n732_));
  XNOR2_X1   g0347(.A1(\a[35] ), .A2(\b[35] ), .ZN(new_n733_));
  NAND2_X1   g0348(.A1(\a[35] ), .A2(\b[35] ), .ZN(new_n734_));
  NOR2_X1    g0349(.A1(\a[35] ), .A2(\b[35] ), .ZN(new_n735_));
  INV_X1     g0350(.I(new_n735_), .ZN(new_n736_));
  NAND2_X1   g0351(.A1(new_n736_), .A2(new_n734_), .ZN(new_n737_));
  NAND2_X1   g0352(.A1(new_n732_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1   g0353(.A1(new_n732_), .A2(new_n733_), .B(new_n738_), .ZN(\f[35] ));
  INV_X1     g0354(.I(new_n732_), .ZN(new_n740_));
  AOI21_X1   g0355(.A1(new_n740_), .A2(new_n734_), .B(new_n735_), .ZN(new_n741_));
  XNOR2_X1   g0356(.A1(\a[36] ), .A2(\b[36] ), .ZN(new_n742_));
  AND2_X2    g0357(.A1(\a[36] ), .A2(\b[36] ), .Z(new_n743_));
  NOR2_X1    g0358(.A1(\a[36] ), .A2(\b[36] ), .ZN(new_n744_));
  OAI21_X1   g0359(.A1(new_n743_), .A2(new_n744_), .B(new_n741_), .ZN(new_n745_));
  OAI21_X1   g0360(.A1(new_n741_), .A2(new_n742_), .B(new_n745_), .ZN(\f[36] ));
  NAND3_X1   g0361(.A1(new_n699_), .A2(new_n722_), .A3(new_n731_), .ZN(new_n747_));
  NOR2_X1    g0362(.A1(new_n744_), .A2(\b[35] ), .ZN(new_n748_));
  AOI21_X1   g0363(.A1(new_n744_), .A2(\b[35] ), .B(\a[35] ), .ZN(new_n749_));
  NOR2_X1    g0364(.A1(new_n749_), .A2(new_n748_), .ZN(new_n750_));
  INV_X1     g0365(.I(new_n750_), .ZN(new_n751_));
  AOI21_X1   g0366(.A1(new_n747_), .A2(new_n728_), .B(new_n751_), .ZN(new_n752_));
  INV_X1     g0367(.I(\a[37] ), .ZN(new_n753_));
  INV_X1     g0368(.I(\b[37] ), .ZN(new_n754_));
  NOR2_X1    g0369(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  XOR2_X1    g0370(.A1(new_n752_), .A2(new_n755_), .Z(new_n756_));
  XOR2_X1    g0371(.A1(new_n756_), .A2(new_n743_), .Z(\f[37] ));
  INV_X1     g0372(.I(new_n743_), .ZN(new_n758_));
  AOI21_X1   g0373(.A1(new_n753_), .A2(new_n754_), .B(new_n758_), .ZN(new_n759_));
  AOI21_X1   g0374(.A1(new_n752_), .A2(new_n759_), .B(new_n755_), .ZN(new_n760_));
  XNOR2_X1   g0375(.A1(\a[38] ), .A2(\b[38] ), .ZN(new_n761_));
  NAND2_X1   g0376(.A1(\a[38] ), .A2(\b[38] ), .ZN(new_n762_));
  NOR2_X1    g0377(.A1(\a[38] ), .A2(\b[38] ), .ZN(new_n763_));
  INV_X1     g0378(.I(new_n763_), .ZN(new_n764_));
  NAND2_X1   g0379(.A1(new_n764_), .A2(new_n762_), .ZN(new_n765_));
  NAND2_X1   g0380(.A1(new_n760_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1   g0381(.A1(new_n760_), .A2(new_n761_), .B(new_n766_), .ZN(\f[38] ));
  INV_X1     g0382(.I(new_n760_), .ZN(new_n768_));
  AOI21_X1   g0383(.A1(new_n768_), .A2(new_n762_), .B(new_n763_), .ZN(new_n769_));
  XNOR2_X1   g0384(.A1(\a[39] ), .A2(\b[39] ), .ZN(new_n770_));
  AND2_X2    g0385(.A1(\a[39] ), .A2(\b[39] ), .Z(new_n771_));
  NOR2_X1    g0386(.A1(\a[39] ), .A2(\b[39] ), .ZN(new_n772_));
  OAI21_X1   g0387(.A1(new_n771_), .A2(new_n772_), .B(new_n769_), .ZN(new_n773_));
  OAI21_X1   g0388(.A1(new_n769_), .A2(new_n770_), .B(new_n773_), .ZN(\f[39] ));
  INV_X1     g0389(.I(new_n771_), .ZN(new_n775_));
  INV_X1     g0390(.I(new_n759_), .ZN(new_n776_));
  NOR3_X1    g0391(.A1(new_n732_), .A2(new_n751_), .A3(new_n776_), .ZN(new_n777_));
  INV_X1     g0392(.I(\b[38] ), .ZN(new_n778_));
  INV_X1     g0393(.I(new_n772_), .ZN(new_n779_));
  AOI21_X1   g0394(.A1(new_n772_), .A2(\b[38] ), .B(\a[38] ), .ZN(new_n780_));
  AOI21_X1   g0395(.A1(new_n778_), .A2(new_n779_), .B(new_n780_), .ZN(new_n781_));
  OAI21_X1   g0396(.A1(new_n777_), .A2(new_n755_), .B(new_n781_), .ZN(new_n782_));
  INV_X1     g0397(.I(\a[40] ), .ZN(new_n783_));
  INV_X1     g0398(.I(\b[40] ), .ZN(new_n784_));
  NOR2_X1    g0399(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  XOR2_X1    g0400(.A1(new_n782_), .A2(new_n785_), .Z(new_n786_));
  XOR2_X1    g0401(.A1(new_n786_), .A2(new_n775_), .Z(\f[40] ));
  INV_X1     g0402(.I(new_n785_), .ZN(new_n788_));
  AOI21_X1   g0403(.A1(new_n783_), .A2(new_n784_), .B(new_n775_), .ZN(new_n789_));
  INV_X1     g0404(.I(new_n789_), .ZN(new_n790_));
  OAI21_X1   g0405(.A1(new_n782_), .A2(new_n790_), .B(new_n788_), .ZN(new_n791_));
  INV_X1     g0406(.I(new_n791_), .ZN(new_n792_));
  XNOR2_X1   g0407(.A1(\a[41] ), .A2(\b[41] ), .ZN(new_n793_));
  INV_X1     g0408(.I(\a[41] ), .ZN(new_n794_));
  INV_X1     g0409(.I(\b[41] ), .ZN(new_n795_));
  NOR2_X1    g0410(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1    g0411(.A1(\a[41] ), .A2(\b[41] ), .ZN(new_n797_));
  OAI21_X1   g0412(.A1(new_n796_), .A2(new_n797_), .B(new_n792_), .ZN(new_n798_));
  OAI21_X1   g0413(.A1(new_n792_), .A2(new_n793_), .B(new_n798_), .ZN(\f[41] ));
  NAND2_X1   g0414(.A1(new_n794_), .A2(new_n795_), .ZN(new_n800_));
  OAI21_X1   g0415(.A1(new_n792_), .A2(new_n796_), .B(new_n800_), .ZN(new_n801_));
  XOR2_X1    g0416(.A1(\a[42] ), .A2(\b[42] ), .Z(new_n802_));
  NAND2_X1   g0417(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1     g0418(.I(\a[42] ), .ZN(new_n804_));
  INV_X1     g0419(.I(\b[42] ), .ZN(new_n805_));
  NOR2_X1    g0420(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1    g0421(.A1(\a[42] ), .A2(\b[42] ), .ZN(new_n807_));
  NOR2_X1    g0422(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1   g0423(.A1(new_n801_), .A2(new_n808_), .B(new_n803_), .ZN(\f[42] ));
  INV_X1     g0424(.I(new_n806_), .ZN(new_n810_));
  INV_X1     g0425(.I(new_n781_), .ZN(new_n811_));
  NOR3_X1    g0426(.A1(new_n760_), .A2(new_n811_), .A3(new_n790_), .ZN(new_n812_));
  NOR2_X1    g0427(.A1(new_n807_), .A2(\b[41] ), .ZN(new_n813_));
  AOI21_X1   g0428(.A1(new_n807_), .A2(\b[41] ), .B(\a[41] ), .ZN(new_n814_));
  NOR2_X1    g0429(.A1(new_n814_), .A2(new_n813_), .ZN(new_n815_));
  OAI21_X1   g0430(.A1(new_n812_), .A2(new_n785_), .B(new_n815_), .ZN(new_n816_));
  INV_X1     g0431(.I(\a[43] ), .ZN(new_n817_));
  INV_X1     g0432(.I(\b[43] ), .ZN(new_n818_));
  NOR2_X1    g0433(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  XOR2_X1    g0434(.A1(new_n816_), .A2(new_n819_), .Z(new_n820_));
  XOR2_X1    g0435(.A1(new_n820_), .A2(new_n810_), .Z(\f[43] ));
  INV_X1     g0436(.I(new_n819_), .ZN(new_n822_));
  AOI21_X1   g0437(.A1(new_n817_), .A2(new_n818_), .B(new_n810_), .ZN(new_n823_));
  INV_X1     g0438(.I(new_n823_), .ZN(new_n824_));
  OAI21_X1   g0439(.A1(new_n816_), .A2(new_n824_), .B(new_n822_), .ZN(new_n825_));
  INV_X1     g0440(.I(new_n825_), .ZN(new_n826_));
  XNOR2_X1   g0441(.A1(\a[44] ), .A2(\b[44] ), .ZN(new_n827_));
  INV_X1     g0442(.I(\a[44] ), .ZN(new_n828_));
  INV_X1     g0443(.I(\b[44] ), .ZN(new_n829_));
  NOR2_X1    g0444(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NOR2_X1    g0445(.A1(\a[44] ), .A2(\b[44] ), .ZN(new_n831_));
  OAI21_X1   g0446(.A1(new_n830_), .A2(new_n831_), .B(new_n826_), .ZN(new_n832_));
  OAI21_X1   g0447(.A1(new_n826_), .A2(new_n827_), .B(new_n832_), .ZN(\f[44] ));
  NAND2_X1   g0448(.A1(new_n828_), .A2(new_n829_), .ZN(new_n834_));
  OAI21_X1   g0449(.A1(new_n826_), .A2(new_n830_), .B(new_n834_), .ZN(new_n835_));
  XOR2_X1    g0450(.A1(\a[45] ), .A2(\b[45] ), .Z(new_n836_));
  NAND2_X1   g0451(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1     g0452(.I(\a[45] ), .ZN(new_n838_));
  INV_X1     g0453(.I(\b[45] ), .ZN(new_n839_));
  NOR2_X1    g0454(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1    g0455(.A1(\a[45] ), .A2(\b[45] ), .ZN(new_n841_));
  NOR2_X1    g0456(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI21_X1   g0457(.A1(new_n835_), .A2(new_n842_), .B(new_n837_), .ZN(\f[45] ));
  INV_X1     g0458(.I(new_n840_), .ZN(new_n844_));
  NAND3_X1   g0459(.A1(new_n791_), .A2(new_n815_), .A3(new_n823_), .ZN(new_n845_));
  INV_X1     g0460(.I(new_n841_), .ZN(new_n846_));
  AOI21_X1   g0461(.A1(new_n841_), .A2(\b[44] ), .B(\a[44] ), .ZN(new_n847_));
  AOI21_X1   g0462(.A1(new_n829_), .A2(new_n846_), .B(new_n847_), .ZN(new_n848_));
  INV_X1     g0463(.I(new_n848_), .ZN(new_n849_));
  AOI21_X1   g0464(.A1(new_n845_), .A2(new_n822_), .B(new_n849_), .ZN(new_n850_));
  INV_X1     g0465(.I(\a[46] ), .ZN(new_n851_));
  INV_X1     g0466(.I(\b[46] ), .ZN(new_n852_));
  NOR2_X1    g0467(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1     g0468(.I(new_n853_), .ZN(new_n854_));
  XOR2_X1    g0469(.A1(new_n850_), .A2(new_n854_), .Z(new_n855_));
  XOR2_X1    g0470(.A1(new_n855_), .A2(new_n844_), .Z(\f[46] ));
  AOI21_X1   g0471(.A1(new_n851_), .A2(new_n852_), .B(new_n844_), .ZN(new_n857_));
  AOI21_X1   g0472(.A1(new_n850_), .A2(new_n857_), .B(new_n853_), .ZN(new_n858_));
  XNOR2_X1   g0473(.A1(\a[47] ), .A2(\b[47] ), .ZN(new_n859_));
  NAND2_X1   g0474(.A1(\a[47] ), .A2(\b[47] ), .ZN(new_n860_));
  NOR2_X1    g0475(.A1(\a[47] ), .A2(\b[47] ), .ZN(new_n861_));
  INV_X1     g0476(.I(new_n861_), .ZN(new_n862_));
  NAND2_X1   g0477(.A1(new_n862_), .A2(new_n860_), .ZN(new_n863_));
  NAND2_X1   g0478(.A1(new_n858_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1   g0479(.A1(new_n858_), .A2(new_n859_), .B(new_n864_), .ZN(\f[47] ));
  INV_X1     g0480(.I(new_n858_), .ZN(new_n866_));
  AOI21_X1   g0481(.A1(new_n866_), .A2(new_n860_), .B(new_n861_), .ZN(new_n867_));
  XNOR2_X1   g0482(.A1(\a[48] ), .A2(\b[48] ), .ZN(new_n868_));
  AND2_X2    g0483(.A1(\a[48] ), .A2(\b[48] ), .Z(new_n869_));
  NOR2_X1    g0484(.A1(\a[48] ), .A2(\b[48] ), .ZN(new_n870_));
  OAI21_X1   g0485(.A1(new_n869_), .A2(new_n870_), .B(new_n867_), .ZN(new_n871_));
  OAI21_X1   g0486(.A1(new_n867_), .A2(new_n868_), .B(new_n871_), .ZN(\f[48] ));
  NAND3_X1   g0487(.A1(new_n825_), .A2(new_n848_), .A3(new_n857_), .ZN(new_n873_));
  NOR2_X1    g0488(.A1(new_n870_), .A2(\b[47] ), .ZN(new_n874_));
  AOI21_X1   g0489(.A1(new_n870_), .A2(\b[47] ), .B(\a[47] ), .ZN(new_n875_));
  NOR2_X1    g0490(.A1(new_n875_), .A2(new_n874_), .ZN(new_n876_));
  INV_X1     g0491(.I(new_n876_), .ZN(new_n877_));
  AOI21_X1   g0492(.A1(new_n873_), .A2(new_n854_), .B(new_n877_), .ZN(new_n878_));
  INV_X1     g0493(.I(\a[49] ), .ZN(new_n879_));
  INV_X1     g0494(.I(\b[49] ), .ZN(new_n880_));
  NOR2_X1    g0495(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  XOR2_X1    g0496(.A1(new_n878_), .A2(new_n881_), .Z(new_n882_));
  XOR2_X1    g0497(.A1(new_n882_), .A2(new_n869_), .Z(\f[49] ));
  INV_X1     g0498(.I(new_n869_), .ZN(new_n884_));
  AOI21_X1   g0499(.A1(new_n879_), .A2(new_n880_), .B(new_n884_), .ZN(new_n885_));
  AOI21_X1   g0500(.A1(new_n878_), .A2(new_n885_), .B(new_n881_), .ZN(new_n886_));
  XNOR2_X1   g0501(.A1(\a[50] ), .A2(\b[50] ), .ZN(new_n887_));
  NAND2_X1   g0502(.A1(\a[50] ), .A2(\b[50] ), .ZN(new_n888_));
  NOR2_X1    g0503(.A1(\a[50] ), .A2(\b[50] ), .ZN(new_n889_));
  INV_X1     g0504(.I(new_n889_), .ZN(new_n890_));
  NAND2_X1   g0505(.A1(new_n890_), .A2(new_n888_), .ZN(new_n891_));
  NAND2_X1   g0506(.A1(new_n886_), .A2(new_n891_), .ZN(new_n892_));
  OAI21_X1   g0507(.A1(new_n886_), .A2(new_n887_), .B(new_n892_), .ZN(\f[50] ));
  INV_X1     g0508(.I(new_n886_), .ZN(new_n894_));
  AOI21_X1   g0509(.A1(new_n894_), .A2(new_n888_), .B(new_n889_), .ZN(new_n895_));
  XNOR2_X1   g0510(.A1(\a[51] ), .A2(\b[51] ), .ZN(new_n896_));
  AND2_X2    g0511(.A1(\a[51] ), .A2(\b[51] ), .Z(new_n897_));
  NOR2_X1    g0512(.A1(\a[51] ), .A2(\b[51] ), .ZN(new_n898_));
  OAI21_X1   g0513(.A1(new_n897_), .A2(new_n898_), .B(new_n895_), .ZN(new_n899_));
  OAI21_X1   g0514(.A1(new_n895_), .A2(new_n896_), .B(new_n899_), .ZN(\f[51] ));
  INV_X1     g0515(.I(new_n897_), .ZN(new_n901_));
  INV_X1     g0516(.I(new_n885_), .ZN(new_n902_));
  NOR3_X1    g0517(.A1(new_n858_), .A2(new_n877_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1     g0518(.I(\b[50] ), .ZN(new_n904_));
  INV_X1     g0519(.I(new_n898_), .ZN(new_n905_));
  AOI21_X1   g0520(.A1(new_n898_), .A2(\b[50] ), .B(\a[50] ), .ZN(new_n906_));
  AOI21_X1   g0521(.A1(new_n904_), .A2(new_n905_), .B(new_n906_), .ZN(new_n907_));
  OAI21_X1   g0522(.A1(new_n903_), .A2(new_n881_), .B(new_n907_), .ZN(new_n908_));
  INV_X1     g0523(.I(\a[52] ), .ZN(new_n909_));
  INV_X1     g0524(.I(\b[52] ), .ZN(new_n910_));
  NOR2_X1    g0525(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  XOR2_X1    g0526(.A1(new_n908_), .A2(new_n911_), .Z(new_n912_));
  XOR2_X1    g0527(.A1(new_n912_), .A2(new_n901_), .Z(\f[52] ));
  INV_X1     g0528(.I(new_n911_), .ZN(new_n914_));
  AOI21_X1   g0529(.A1(new_n909_), .A2(new_n910_), .B(new_n901_), .ZN(new_n915_));
  INV_X1     g0530(.I(new_n915_), .ZN(new_n916_));
  OAI21_X1   g0531(.A1(new_n908_), .A2(new_n916_), .B(new_n914_), .ZN(new_n917_));
  INV_X1     g0532(.I(new_n917_), .ZN(new_n918_));
  XNOR2_X1   g0533(.A1(\a[53] ), .A2(\b[53] ), .ZN(new_n919_));
  INV_X1     g0534(.I(\a[53] ), .ZN(new_n920_));
  INV_X1     g0535(.I(\b[53] ), .ZN(new_n921_));
  NOR2_X1    g0536(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NOR2_X1    g0537(.A1(\a[53] ), .A2(\b[53] ), .ZN(new_n923_));
  OAI21_X1   g0538(.A1(new_n922_), .A2(new_n923_), .B(new_n918_), .ZN(new_n924_));
  OAI21_X1   g0539(.A1(new_n918_), .A2(new_n919_), .B(new_n924_), .ZN(\f[53] ));
  NAND2_X1   g0540(.A1(new_n920_), .A2(new_n921_), .ZN(new_n926_));
  OAI21_X1   g0541(.A1(new_n918_), .A2(new_n922_), .B(new_n926_), .ZN(new_n927_));
  XOR2_X1    g0542(.A1(\a[54] ), .A2(\b[54] ), .Z(new_n928_));
  NAND2_X1   g0543(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1     g0544(.I(\a[54] ), .ZN(new_n930_));
  INV_X1     g0545(.I(\b[54] ), .ZN(new_n931_));
  NOR2_X1    g0546(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1    g0547(.A1(\a[54] ), .A2(\b[54] ), .ZN(new_n933_));
  NOR2_X1    g0548(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  OAI21_X1   g0549(.A1(new_n927_), .A2(new_n934_), .B(new_n929_), .ZN(\f[54] ));
  INV_X1     g0550(.I(new_n932_), .ZN(new_n936_));
  INV_X1     g0551(.I(new_n907_), .ZN(new_n937_));
  NOR3_X1    g0552(.A1(new_n886_), .A2(new_n937_), .A3(new_n916_), .ZN(new_n938_));
  NOR2_X1    g0553(.A1(new_n933_), .A2(\b[53] ), .ZN(new_n939_));
  AOI21_X1   g0554(.A1(new_n933_), .A2(\b[53] ), .B(\a[53] ), .ZN(new_n940_));
  NOR2_X1    g0555(.A1(new_n940_), .A2(new_n939_), .ZN(new_n941_));
  OAI21_X1   g0556(.A1(new_n938_), .A2(new_n911_), .B(new_n941_), .ZN(new_n942_));
  INV_X1     g0557(.I(\a[55] ), .ZN(new_n943_));
  INV_X1     g0558(.I(\b[55] ), .ZN(new_n944_));
  NOR2_X1    g0559(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  XOR2_X1    g0560(.A1(new_n942_), .A2(new_n945_), .Z(new_n946_));
  XOR2_X1    g0561(.A1(new_n946_), .A2(new_n936_), .Z(\f[55] ));
  INV_X1     g0562(.I(new_n945_), .ZN(new_n948_));
  AOI21_X1   g0563(.A1(new_n943_), .A2(new_n944_), .B(new_n936_), .ZN(new_n949_));
  INV_X1     g0564(.I(new_n949_), .ZN(new_n950_));
  OAI21_X1   g0565(.A1(new_n942_), .A2(new_n950_), .B(new_n948_), .ZN(new_n951_));
  INV_X1     g0566(.I(new_n951_), .ZN(new_n952_));
  XNOR2_X1   g0567(.A1(\a[56] ), .A2(\b[56] ), .ZN(new_n953_));
  INV_X1     g0568(.I(\a[56] ), .ZN(new_n954_));
  INV_X1     g0569(.I(\b[56] ), .ZN(new_n955_));
  NOR2_X1    g0570(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  NOR2_X1    g0571(.A1(\a[56] ), .A2(\b[56] ), .ZN(new_n957_));
  OAI21_X1   g0572(.A1(new_n956_), .A2(new_n957_), .B(new_n952_), .ZN(new_n958_));
  OAI21_X1   g0573(.A1(new_n952_), .A2(new_n953_), .B(new_n958_), .ZN(\f[56] ));
  NAND2_X1   g0574(.A1(new_n954_), .A2(new_n955_), .ZN(new_n960_));
  OAI21_X1   g0575(.A1(new_n952_), .A2(new_n956_), .B(new_n960_), .ZN(new_n961_));
  XOR2_X1    g0576(.A1(\a[57] ), .A2(\b[57] ), .Z(new_n962_));
  NAND2_X1   g0577(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  INV_X1     g0578(.I(\a[57] ), .ZN(new_n964_));
  INV_X1     g0579(.I(\b[57] ), .ZN(new_n965_));
  NOR2_X1    g0580(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  NOR2_X1    g0581(.A1(\a[57] ), .A2(\b[57] ), .ZN(new_n967_));
  NOR2_X1    g0582(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  OAI21_X1   g0583(.A1(new_n961_), .A2(new_n968_), .B(new_n963_), .ZN(\f[57] ));
  INV_X1     g0584(.I(new_n966_), .ZN(new_n970_));
  NAND3_X1   g0585(.A1(new_n917_), .A2(new_n941_), .A3(new_n949_), .ZN(new_n971_));
  INV_X1     g0586(.I(new_n967_), .ZN(new_n972_));
  AOI21_X1   g0587(.A1(new_n967_), .A2(\b[56] ), .B(\a[56] ), .ZN(new_n973_));
  AOI21_X1   g0588(.A1(new_n955_), .A2(new_n972_), .B(new_n973_), .ZN(new_n974_));
  INV_X1     g0589(.I(new_n974_), .ZN(new_n975_));
  AOI21_X1   g0590(.A1(new_n971_), .A2(new_n948_), .B(new_n975_), .ZN(new_n976_));
  INV_X1     g0591(.I(\a[58] ), .ZN(new_n977_));
  INV_X1     g0592(.I(\b[58] ), .ZN(new_n978_));
  NOR2_X1    g0593(.A1(new_n977_), .A2(new_n978_), .ZN(new_n979_));
  INV_X1     g0594(.I(new_n979_), .ZN(new_n980_));
  XOR2_X1    g0595(.A1(new_n976_), .A2(new_n980_), .Z(new_n981_));
  XOR2_X1    g0596(.A1(new_n981_), .A2(new_n970_), .Z(\f[58] ));
  AOI21_X1   g0597(.A1(new_n977_), .A2(new_n978_), .B(new_n970_), .ZN(new_n983_));
  AOI21_X1   g0598(.A1(new_n976_), .A2(new_n983_), .B(new_n979_), .ZN(new_n984_));
  XNOR2_X1   g0599(.A1(\a[59] ), .A2(\b[59] ), .ZN(new_n985_));
  NAND2_X1   g0600(.A1(\a[59] ), .A2(\b[59] ), .ZN(new_n986_));
  NOR2_X1    g0601(.A1(\a[59] ), .A2(\b[59] ), .ZN(new_n987_));
  INV_X1     g0602(.I(new_n987_), .ZN(new_n988_));
  NAND2_X1   g0603(.A1(new_n988_), .A2(new_n986_), .ZN(new_n989_));
  NAND2_X1   g0604(.A1(new_n984_), .A2(new_n989_), .ZN(new_n990_));
  OAI21_X1   g0605(.A1(new_n984_), .A2(new_n985_), .B(new_n990_), .ZN(\f[59] ));
  INV_X1     g0606(.I(new_n984_), .ZN(new_n992_));
  AOI21_X1   g0607(.A1(new_n992_), .A2(new_n986_), .B(new_n987_), .ZN(new_n993_));
  XNOR2_X1   g0608(.A1(\a[60] ), .A2(\b[60] ), .ZN(new_n994_));
  AND2_X2    g0609(.A1(\a[60] ), .A2(\b[60] ), .Z(new_n995_));
  NOR2_X1    g0610(.A1(\a[60] ), .A2(\b[60] ), .ZN(new_n996_));
  OAI21_X1   g0611(.A1(new_n995_), .A2(new_n996_), .B(new_n993_), .ZN(new_n997_));
  OAI21_X1   g0612(.A1(new_n993_), .A2(new_n994_), .B(new_n997_), .ZN(\f[60] ));
  NAND3_X1   g0613(.A1(new_n951_), .A2(new_n974_), .A3(new_n983_), .ZN(new_n999_));
  NOR2_X1    g0614(.A1(new_n996_), .A2(\b[59] ), .ZN(new_n1000_));
  AOI21_X1   g0615(.A1(new_n996_), .A2(\b[59] ), .B(\a[59] ), .ZN(new_n1001_));
  NOR2_X1    g0616(.A1(new_n1001_), .A2(new_n1000_), .ZN(new_n1002_));
  INV_X1     g0617(.I(new_n1002_), .ZN(new_n1003_));
  AOI21_X1   g0618(.A1(new_n999_), .A2(new_n980_), .B(new_n1003_), .ZN(new_n1004_));
  INV_X1     g0619(.I(\a[61] ), .ZN(new_n1005_));
  INV_X1     g0620(.I(\b[61] ), .ZN(new_n1006_));
  NOR2_X1    g0621(.A1(new_n1005_), .A2(new_n1006_), .ZN(new_n1007_));
  XOR2_X1    g0622(.A1(new_n1004_), .A2(new_n1007_), .Z(new_n1008_));
  XOR2_X1    g0623(.A1(new_n1008_), .A2(new_n995_), .Z(\f[61] ));
  INV_X1     g0624(.I(new_n995_), .ZN(new_n1010_));
  AOI21_X1   g0625(.A1(new_n1005_), .A2(new_n1006_), .B(new_n1010_), .ZN(new_n1011_));
  AOI21_X1   g0626(.A1(new_n1004_), .A2(new_n1011_), .B(new_n1007_), .ZN(new_n1012_));
  XNOR2_X1   g0627(.A1(\a[62] ), .A2(\b[62] ), .ZN(new_n1013_));
  NAND2_X1   g0628(.A1(\a[62] ), .A2(\b[62] ), .ZN(new_n1014_));
  NOR2_X1    g0629(.A1(\a[62] ), .A2(\b[62] ), .ZN(new_n1015_));
  INV_X1     g0630(.I(new_n1015_), .ZN(new_n1016_));
  NAND2_X1   g0631(.A1(new_n1016_), .A2(new_n1014_), .ZN(new_n1017_));
  NAND2_X1   g0632(.A1(new_n1012_), .A2(new_n1017_), .ZN(new_n1018_));
  OAI21_X1   g0633(.A1(new_n1012_), .A2(new_n1013_), .B(new_n1018_), .ZN(\f[62] ));
  INV_X1     g0634(.I(new_n1012_), .ZN(new_n1020_));
  AOI21_X1   g0635(.A1(new_n1020_), .A2(new_n1014_), .B(new_n1015_), .ZN(new_n1021_));
  XNOR2_X1   g0636(.A1(\a[63] ), .A2(\b[63] ), .ZN(new_n1022_));
  AND2_X2    g0637(.A1(\a[63] ), .A2(\b[63] ), .Z(new_n1023_));
  NOR2_X1    g0638(.A1(\a[63] ), .A2(\b[63] ), .ZN(new_n1024_));
  OAI21_X1   g0639(.A1(new_n1023_), .A2(new_n1024_), .B(new_n1021_), .ZN(new_n1025_));
  OAI21_X1   g0640(.A1(new_n1021_), .A2(new_n1022_), .B(new_n1025_), .ZN(\f[63] ));
  INV_X1     g0641(.I(new_n1023_), .ZN(new_n1027_));
  INV_X1     g0642(.I(new_n1011_), .ZN(new_n1028_));
  NOR3_X1    g0643(.A1(new_n984_), .A2(new_n1003_), .A3(new_n1028_), .ZN(new_n1029_));
  INV_X1     g0644(.I(\b[62] ), .ZN(new_n1030_));
  INV_X1     g0645(.I(new_n1024_), .ZN(new_n1031_));
  AOI21_X1   g0646(.A1(new_n1024_), .A2(\b[62] ), .B(\a[62] ), .ZN(new_n1032_));
  AOI21_X1   g0647(.A1(new_n1030_), .A2(new_n1031_), .B(new_n1032_), .ZN(new_n1033_));
  OAI21_X1   g0648(.A1(new_n1029_), .A2(new_n1007_), .B(new_n1033_), .ZN(new_n1034_));
  INV_X1     g0649(.I(\a[64] ), .ZN(new_n1035_));
  INV_X1     g0650(.I(\b[64] ), .ZN(new_n1036_));
  NOR2_X1    g0651(.A1(new_n1035_), .A2(new_n1036_), .ZN(new_n1037_));
  XOR2_X1    g0652(.A1(new_n1034_), .A2(new_n1037_), .Z(new_n1038_));
  XOR2_X1    g0653(.A1(new_n1038_), .A2(new_n1027_), .Z(\f[64] ));
  INV_X1     g0654(.I(new_n1037_), .ZN(new_n1040_));
  AOI21_X1   g0655(.A1(new_n1035_), .A2(new_n1036_), .B(new_n1027_), .ZN(new_n1041_));
  INV_X1     g0656(.I(new_n1041_), .ZN(new_n1042_));
  OAI21_X1   g0657(.A1(new_n1034_), .A2(new_n1042_), .B(new_n1040_), .ZN(new_n1043_));
  INV_X1     g0658(.I(new_n1043_), .ZN(new_n1044_));
  XNOR2_X1   g0659(.A1(\a[65] ), .A2(\b[65] ), .ZN(new_n1045_));
  INV_X1     g0660(.I(\a[65] ), .ZN(new_n1046_));
  INV_X1     g0661(.I(\b[65] ), .ZN(new_n1047_));
  NOR2_X1    g0662(.A1(new_n1046_), .A2(new_n1047_), .ZN(new_n1048_));
  NOR2_X1    g0663(.A1(\a[65] ), .A2(\b[65] ), .ZN(new_n1049_));
  OAI21_X1   g0664(.A1(new_n1048_), .A2(new_n1049_), .B(new_n1044_), .ZN(new_n1050_));
  OAI21_X1   g0665(.A1(new_n1044_), .A2(new_n1045_), .B(new_n1050_), .ZN(\f[65] ));
  NAND2_X1   g0666(.A1(new_n1046_), .A2(new_n1047_), .ZN(new_n1052_));
  OAI21_X1   g0667(.A1(new_n1044_), .A2(new_n1048_), .B(new_n1052_), .ZN(new_n1053_));
  XOR2_X1    g0668(.A1(\a[66] ), .A2(\b[66] ), .Z(new_n1054_));
  NAND2_X1   g0669(.A1(new_n1053_), .A2(new_n1054_), .ZN(new_n1055_));
  INV_X1     g0670(.I(\a[66] ), .ZN(new_n1056_));
  INV_X1     g0671(.I(\b[66] ), .ZN(new_n1057_));
  NOR2_X1    g0672(.A1(new_n1056_), .A2(new_n1057_), .ZN(new_n1058_));
  NOR2_X1    g0673(.A1(\a[66] ), .A2(\b[66] ), .ZN(new_n1059_));
  NOR2_X1    g0674(.A1(new_n1058_), .A2(new_n1059_), .ZN(new_n1060_));
  OAI21_X1   g0675(.A1(new_n1053_), .A2(new_n1060_), .B(new_n1055_), .ZN(\f[66] ));
  INV_X1     g0676(.I(new_n1058_), .ZN(new_n1062_));
  INV_X1     g0677(.I(new_n1033_), .ZN(new_n1063_));
  NOR3_X1    g0678(.A1(new_n1012_), .A2(new_n1063_), .A3(new_n1042_), .ZN(new_n1064_));
  NOR2_X1    g0679(.A1(new_n1059_), .A2(\b[65] ), .ZN(new_n1065_));
  AOI21_X1   g0680(.A1(new_n1059_), .A2(\b[65] ), .B(\a[65] ), .ZN(new_n1066_));
  NOR2_X1    g0681(.A1(new_n1066_), .A2(new_n1065_), .ZN(new_n1067_));
  OAI21_X1   g0682(.A1(new_n1064_), .A2(new_n1037_), .B(new_n1067_), .ZN(new_n1068_));
  INV_X1     g0683(.I(\a[67] ), .ZN(new_n1069_));
  INV_X1     g0684(.I(\b[67] ), .ZN(new_n1070_));
  NOR2_X1    g0685(.A1(new_n1069_), .A2(new_n1070_), .ZN(new_n1071_));
  XOR2_X1    g0686(.A1(new_n1068_), .A2(new_n1071_), .Z(new_n1072_));
  XOR2_X1    g0687(.A1(new_n1072_), .A2(new_n1062_), .Z(\f[67] ));
  INV_X1     g0688(.I(new_n1071_), .ZN(new_n1074_));
  AOI21_X1   g0689(.A1(new_n1069_), .A2(new_n1070_), .B(new_n1062_), .ZN(new_n1075_));
  INV_X1     g0690(.I(new_n1075_), .ZN(new_n1076_));
  OAI21_X1   g0691(.A1(new_n1068_), .A2(new_n1076_), .B(new_n1074_), .ZN(new_n1077_));
  INV_X1     g0692(.I(new_n1077_), .ZN(new_n1078_));
  XNOR2_X1   g0693(.A1(\a[68] ), .A2(\b[68] ), .ZN(new_n1079_));
  INV_X1     g0694(.I(\a[68] ), .ZN(new_n1080_));
  INV_X1     g0695(.I(\b[68] ), .ZN(new_n1081_));
  NOR2_X1    g0696(.A1(new_n1080_), .A2(new_n1081_), .ZN(new_n1082_));
  NOR2_X1    g0697(.A1(\a[68] ), .A2(\b[68] ), .ZN(new_n1083_));
  OAI21_X1   g0698(.A1(new_n1082_), .A2(new_n1083_), .B(new_n1078_), .ZN(new_n1084_));
  OAI21_X1   g0699(.A1(new_n1078_), .A2(new_n1079_), .B(new_n1084_), .ZN(\f[68] ));
  NAND2_X1   g0700(.A1(new_n1080_), .A2(new_n1081_), .ZN(new_n1086_));
  OAI21_X1   g0701(.A1(new_n1078_), .A2(new_n1082_), .B(new_n1086_), .ZN(new_n1087_));
  XOR2_X1    g0702(.A1(\a[69] ), .A2(\b[69] ), .Z(new_n1088_));
  NAND2_X1   g0703(.A1(new_n1087_), .A2(new_n1088_), .ZN(new_n1089_));
  INV_X1     g0704(.I(\a[69] ), .ZN(new_n1090_));
  INV_X1     g0705(.I(\b[69] ), .ZN(new_n1091_));
  NOR2_X1    g0706(.A1(new_n1090_), .A2(new_n1091_), .ZN(new_n1092_));
  NOR2_X1    g0707(.A1(\a[69] ), .A2(\b[69] ), .ZN(new_n1093_));
  NOR2_X1    g0708(.A1(new_n1092_), .A2(new_n1093_), .ZN(new_n1094_));
  OAI21_X1   g0709(.A1(new_n1087_), .A2(new_n1094_), .B(new_n1089_), .ZN(\f[69] ));
  INV_X1     g0710(.I(new_n1092_), .ZN(new_n1096_));
  NAND3_X1   g0711(.A1(new_n1043_), .A2(new_n1067_), .A3(new_n1075_), .ZN(new_n1097_));
  INV_X1     g0712(.I(new_n1093_), .ZN(new_n1098_));
  AOI21_X1   g0713(.A1(new_n1093_), .A2(\b[68] ), .B(\a[68] ), .ZN(new_n1099_));
  AOI21_X1   g0714(.A1(new_n1081_), .A2(new_n1098_), .B(new_n1099_), .ZN(new_n1100_));
  INV_X1     g0715(.I(new_n1100_), .ZN(new_n1101_));
  AOI21_X1   g0716(.A1(new_n1097_), .A2(new_n1074_), .B(new_n1101_), .ZN(new_n1102_));
  INV_X1     g0717(.I(\a[70] ), .ZN(new_n1103_));
  INV_X1     g0718(.I(\b[70] ), .ZN(new_n1104_));
  NOR2_X1    g0719(.A1(new_n1103_), .A2(new_n1104_), .ZN(new_n1105_));
  INV_X1     g0720(.I(new_n1105_), .ZN(new_n1106_));
  XOR2_X1    g0721(.A1(new_n1102_), .A2(new_n1106_), .Z(new_n1107_));
  XOR2_X1    g0722(.A1(new_n1107_), .A2(new_n1096_), .Z(\f[70] ));
  AOI21_X1   g0723(.A1(new_n1103_), .A2(new_n1104_), .B(new_n1096_), .ZN(new_n1109_));
  AOI21_X1   g0724(.A1(new_n1102_), .A2(new_n1109_), .B(new_n1105_), .ZN(new_n1110_));
  XNOR2_X1   g0725(.A1(\a[71] ), .A2(\b[71] ), .ZN(new_n1111_));
  NAND2_X1   g0726(.A1(\a[71] ), .A2(\b[71] ), .ZN(new_n1112_));
  NOR2_X1    g0727(.A1(\a[71] ), .A2(\b[71] ), .ZN(new_n1113_));
  INV_X1     g0728(.I(new_n1113_), .ZN(new_n1114_));
  NAND2_X1   g0729(.A1(new_n1114_), .A2(new_n1112_), .ZN(new_n1115_));
  NAND2_X1   g0730(.A1(new_n1110_), .A2(new_n1115_), .ZN(new_n1116_));
  OAI21_X1   g0731(.A1(new_n1110_), .A2(new_n1111_), .B(new_n1116_), .ZN(\f[71] ));
  INV_X1     g0732(.I(new_n1110_), .ZN(new_n1118_));
  AOI21_X1   g0733(.A1(new_n1118_), .A2(new_n1112_), .B(new_n1113_), .ZN(new_n1119_));
  XNOR2_X1   g0734(.A1(\a[72] ), .A2(\b[72] ), .ZN(new_n1120_));
  AND2_X2    g0735(.A1(\a[72] ), .A2(\b[72] ), .Z(new_n1121_));
  NOR2_X1    g0736(.A1(\a[72] ), .A2(\b[72] ), .ZN(new_n1122_));
  OAI21_X1   g0737(.A1(new_n1121_), .A2(new_n1122_), .B(new_n1119_), .ZN(new_n1123_));
  OAI21_X1   g0738(.A1(new_n1119_), .A2(new_n1120_), .B(new_n1123_), .ZN(\f[72] ));
  NAND3_X1   g0739(.A1(new_n1077_), .A2(new_n1100_), .A3(new_n1109_), .ZN(new_n1125_));
  NOR2_X1    g0740(.A1(new_n1122_), .A2(\b[71] ), .ZN(new_n1126_));
  AOI21_X1   g0741(.A1(new_n1122_), .A2(\b[71] ), .B(\a[71] ), .ZN(new_n1127_));
  NOR2_X1    g0742(.A1(new_n1127_), .A2(new_n1126_), .ZN(new_n1128_));
  INV_X1     g0743(.I(new_n1128_), .ZN(new_n1129_));
  AOI21_X1   g0744(.A1(new_n1125_), .A2(new_n1106_), .B(new_n1129_), .ZN(new_n1130_));
  INV_X1     g0745(.I(\a[73] ), .ZN(new_n1131_));
  INV_X1     g0746(.I(\b[73] ), .ZN(new_n1132_));
  NOR2_X1    g0747(.A1(new_n1131_), .A2(new_n1132_), .ZN(new_n1133_));
  XOR2_X1    g0748(.A1(new_n1130_), .A2(new_n1133_), .Z(new_n1134_));
  XOR2_X1    g0749(.A1(new_n1134_), .A2(new_n1121_), .Z(\f[73] ));
  INV_X1     g0750(.I(new_n1121_), .ZN(new_n1136_));
  AOI21_X1   g0751(.A1(new_n1131_), .A2(new_n1132_), .B(new_n1136_), .ZN(new_n1137_));
  AOI21_X1   g0752(.A1(new_n1130_), .A2(new_n1137_), .B(new_n1133_), .ZN(new_n1138_));
  XNOR2_X1   g0753(.A1(\a[74] ), .A2(\b[74] ), .ZN(new_n1139_));
  NAND2_X1   g0754(.A1(\a[74] ), .A2(\b[74] ), .ZN(new_n1140_));
  NOR2_X1    g0755(.A1(\a[74] ), .A2(\b[74] ), .ZN(new_n1141_));
  INV_X1     g0756(.I(new_n1141_), .ZN(new_n1142_));
  NAND2_X1   g0757(.A1(new_n1142_), .A2(new_n1140_), .ZN(new_n1143_));
  NAND2_X1   g0758(.A1(new_n1138_), .A2(new_n1143_), .ZN(new_n1144_));
  OAI21_X1   g0759(.A1(new_n1138_), .A2(new_n1139_), .B(new_n1144_), .ZN(\f[74] ));
  INV_X1     g0760(.I(new_n1138_), .ZN(new_n1146_));
  AOI21_X1   g0761(.A1(new_n1146_), .A2(new_n1140_), .B(new_n1141_), .ZN(new_n1147_));
  XNOR2_X1   g0762(.A1(\a[75] ), .A2(\b[75] ), .ZN(new_n1148_));
  AND2_X2    g0763(.A1(\a[75] ), .A2(\b[75] ), .Z(new_n1149_));
  NOR2_X1    g0764(.A1(\a[75] ), .A2(\b[75] ), .ZN(new_n1150_));
  OAI21_X1   g0765(.A1(new_n1149_), .A2(new_n1150_), .B(new_n1147_), .ZN(new_n1151_));
  OAI21_X1   g0766(.A1(new_n1147_), .A2(new_n1148_), .B(new_n1151_), .ZN(\f[75] ));
  INV_X1     g0767(.I(new_n1149_), .ZN(new_n1153_));
  INV_X1     g0768(.I(new_n1137_), .ZN(new_n1154_));
  NOR3_X1    g0769(.A1(new_n1110_), .A2(new_n1129_), .A3(new_n1154_), .ZN(new_n1155_));
  INV_X1     g0770(.I(\b[74] ), .ZN(new_n1156_));
  INV_X1     g0771(.I(new_n1150_), .ZN(new_n1157_));
  AOI21_X1   g0772(.A1(new_n1150_), .A2(\b[74] ), .B(\a[74] ), .ZN(new_n1158_));
  AOI21_X1   g0773(.A1(new_n1156_), .A2(new_n1157_), .B(new_n1158_), .ZN(new_n1159_));
  OAI21_X1   g0774(.A1(new_n1155_), .A2(new_n1133_), .B(new_n1159_), .ZN(new_n1160_));
  INV_X1     g0775(.I(\a[76] ), .ZN(new_n1161_));
  INV_X1     g0776(.I(\b[76] ), .ZN(new_n1162_));
  NOR2_X1    g0777(.A1(new_n1161_), .A2(new_n1162_), .ZN(new_n1163_));
  XOR2_X1    g0778(.A1(new_n1160_), .A2(new_n1163_), .Z(new_n1164_));
  XOR2_X1    g0779(.A1(new_n1164_), .A2(new_n1153_), .Z(\f[76] ));
  INV_X1     g0780(.I(new_n1163_), .ZN(new_n1166_));
  AOI21_X1   g0781(.A1(new_n1161_), .A2(new_n1162_), .B(new_n1153_), .ZN(new_n1167_));
  INV_X1     g0782(.I(new_n1167_), .ZN(new_n1168_));
  OAI21_X1   g0783(.A1(new_n1160_), .A2(new_n1168_), .B(new_n1166_), .ZN(new_n1169_));
  INV_X1     g0784(.I(new_n1169_), .ZN(new_n1170_));
  XNOR2_X1   g0785(.A1(\a[77] ), .A2(\b[77] ), .ZN(new_n1171_));
  INV_X1     g0786(.I(\a[77] ), .ZN(new_n1172_));
  INV_X1     g0787(.I(\b[77] ), .ZN(new_n1173_));
  NOR2_X1    g0788(.A1(new_n1172_), .A2(new_n1173_), .ZN(new_n1174_));
  NOR2_X1    g0789(.A1(\a[77] ), .A2(\b[77] ), .ZN(new_n1175_));
  OAI21_X1   g0790(.A1(new_n1174_), .A2(new_n1175_), .B(new_n1170_), .ZN(new_n1176_));
  OAI21_X1   g0791(.A1(new_n1170_), .A2(new_n1171_), .B(new_n1176_), .ZN(\f[77] ));
  NAND2_X1   g0792(.A1(new_n1172_), .A2(new_n1173_), .ZN(new_n1178_));
  OAI21_X1   g0793(.A1(new_n1170_), .A2(new_n1174_), .B(new_n1178_), .ZN(new_n1179_));
  XOR2_X1    g0794(.A1(\a[78] ), .A2(\b[78] ), .Z(new_n1180_));
  NAND2_X1   g0795(.A1(new_n1179_), .A2(new_n1180_), .ZN(new_n1181_));
  INV_X1     g0796(.I(\a[78] ), .ZN(new_n1182_));
  INV_X1     g0797(.I(\b[78] ), .ZN(new_n1183_));
  NOR2_X1    g0798(.A1(new_n1182_), .A2(new_n1183_), .ZN(new_n1184_));
  NOR2_X1    g0799(.A1(\a[78] ), .A2(\b[78] ), .ZN(new_n1185_));
  NOR2_X1    g0800(.A1(new_n1184_), .A2(new_n1185_), .ZN(new_n1186_));
  OAI21_X1   g0801(.A1(new_n1179_), .A2(new_n1186_), .B(new_n1181_), .ZN(\f[78] ));
  INV_X1     g0802(.I(new_n1184_), .ZN(new_n1188_));
  INV_X1     g0803(.I(new_n1159_), .ZN(new_n1189_));
  NOR3_X1    g0804(.A1(new_n1138_), .A2(new_n1189_), .A3(new_n1168_), .ZN(new_n1190_));
  NOR2_X1    g0805(.A1(new_n1185_), .A2(\b[77] ), .ZN(new_n1191_));
  AOI21_X1   g0806(.A1(new_n1185_), .A2(\b[77] ), .B(\a[77] ), .ZN(new_n1192_));
  NOR2_X1    g0807(.A1(new_n1192_), .A2(new_n1191_), .ZN(new_n1193_));
  OAI21_X1   g0808(.A1(new_n1190_), .A2(new_n1163_), .B(new_n1193_), .ZN(new_n1194_));
  INV_X1     g0809(.I(\a[79] ), .ZN(new_n1195_));
  INV_X1     g0810(.I(\b[79] ), .ZN(new_n1196_));
  NOR2_X1    g0811(.A1(new_n1195_), .A2(new_n1196_), .ZN(new_n1197_));
  XOR2_X1    g0812(.A1(new_n1194_), .A2(new_n1197_), .Z(new_n1198_));
  XOR2_X1    g0813(.A1(new_n1198_), .A2(new_n1188_), .Z(\f[79] ));
  INV_X1     g0814(.I(new_n1197_), .ZN(new_n1200_));
  AOI21_X1   g0815(.A1(new_n1195_), .A2(new_n1196_), .B(new_n1188_), .ZN(new_n1201_));
  INV_X1     g0816(.I(new_n1201_), .ZN(new_n1202_));
  OAI21_X1   g0817(.A1(new_n1194_), .A2(new_n1202_), .B(new_n1200_), .ZN(new_n1203_));
  INV_X1     g0818(.I(new_n1203_), .ZN(new_n1204_));
  XNOR2_X1   g0819(.A1(\a[80] ), .A2(\b[80] ), .ZN(new_n1205_));
  INV_X1     g0820(.I(\a[80] ), .ZN(new_n1206_));
  INV_X1     g0821(.I(\b[80] ), .ZN(new_n1207_));
  NOR2_X1    g0822(.A1(new_n1206_), .A2(new_n1207_), .ZN(new_n1208_));
  NOR2_X1    g0823(.A1(\a[80] ), .A2(\b[80] ), .ZN(new_n1209_));
  OAI21_X1   g0824(.A1(new_n1208_), .A2(new_n1209_), .B(new_n1204_), .ZN(new_n1210_));
  OAI21_X1   g0825(.A1(new_n1204_), .A2(new_n1205_), .B(new_n1210_), .ZN(\f[80] ));
  NAND2_X1   g0826(.A1(new_n1206_), .A2(new_n1207_), .ZN(new_n1212_));
  OAI21_X1   g0827(.A1(new_n1204_), .A2(new_n1208_), .B(new_n1212_), .ZN(new_n1213_));
  XOR2_X1    g0828(.A1(\a[81] ), .A2(\b[81] ), .Z(new_n1214_));
  NAND2_X1   g0829(.A1(new_n1213_), .A2(new_n1214_), .ZN(new_n1215_));
  INV_X1     g0830(.I(\a[81] ), .ZN(new_n1216_));
  INV_X1     g0831(.I(\b[81] ), .ZN(new_n1217_));
  NOR2_X1    g0832(.A1(new_n1216_), .A2(new_n1217_), .ZN(new_n1218_));
  NOR2_X1    g0833(.A1(\a[81] ), .A2(\b[81] ), .ZN(new_n1219_));
  NOR2_X1    g0834(.A1(new_n1218_), .A2(new_n1219_), .ZN(new_n1220_));
  OAI21_X1   g0835(.A1(new_n1213_), .A2(new_n1220_), .B(new_n1215_), .ZN(\f[81] ));
  INV_X1     g0836(.I(new_n1218_), .ZN(new_n1222_));
  NAND3_X1   g0837(.A1(new_n1169_), .A2(new_n1193_), .A3(new_n1201_), .ZN(new_n1223_));
  INV_X1     g0838(.I(new_n1219_), .ZN(new_n1224_));
  AOI21_X1   g0839(.A1(new_n1219_), .A2(\b[80] ), .B(\a[80] ), .ZN(new_n1225_));
  AOI21_X1   g0840(.A1(new_n1207_), .A2(new_n1224_), .B(new_n1225_), .ZN(new_n1226_));
  INV_X1     g0841(.I(new_n1226_), .ZN(new_n1227_));
  AOI21_X1   g0842(.A1(new_n1223_), .A2(new_n1200_), .B(new_n1227_), .ZN(new_n1228_));
  INV_X1     g0843(.I(\a[82] ), .ZN(new_n1229_));
  INV_X1     g0844(.I(\b[82] ), .ZN(new_n1230_));
  NOR2_X1    g0845(.A1(new_n1229_), .A2(new_n1230_), .ZN(new_n1231_));
  INV_X1     g0846(.I(new_n1231_), .ZN(new_n1232_));
  XOR2_X1    g0847(.A1(new_n1228_), .A2(new_n1232_), .Z(new_n1233_));
  XOR2_X1    g0848(.A1(new_n1233_), .A2(new_n1222_), .Z(\f[82] ));
  AOI21_X1   g0849(.A1(new_n1229_), .A2(new_n1230_), .B(new_n1222_), .ZN(new_n1235_));
  AOI21_X1   g0850(.A1(new_n1228_), .A2(new_n1235_), .B(new_n1231_), .ZN(new_n1236_));
  XNOR2_X1   g0851(.A1(\a[83] ), .A2(\b[83] ), .ZN(new_n1237_));
  NAND2_X1   g0852(.A1(\a[83] ), .A2(\b[83] ), .ZN(new_n1238_));
  NOR2_X1    g0853(.A1(\a[83] ), .A2(\b[83] ), .ZN(new_n1239_));
  INV_X1     g0854(.I(new_n1239_), .ZN(new_n1240_));
  NAND2_X1   g0855(.A1(new_n1240_), .A2(new_n1238_), .ZN(new_n1241_));
  NAND2_X1   g0856(.A1(new_n1236_), .A2(new_n1241_), .ZN(new_n1242_));
  OAI21_X1   g0857(.A1(new_n1236_), .A2(new_n1237_), .B(new_n1242_), .ZN(\f[83] ));
  INV_X1     g0858(.I(new_n1236_), .ZN(new_n1244_));
  AOI21_X1   g0859(.A1(new_n1244_), .A2(new_n1238_), .B(new_n1239_), .ZN(new_n1245_));
  XNOR2_X1   g0860(.A1(\a[84] ), .A2(\b[84] ), .ZN(new_n1246_));
  AND2_X2    g0861(.A1(\a[84] ), .A2(\b[84] ), .Z(new_n1247_));
  NOR2_X1    g0862(.A1(\a[84] ), .A2(\b[84] ), .ZN(new_n1248_));
  OAI21_X1   g0863(.A1(new_n1247_), .A2(new_n1248_), .B(new_n1245_), .ZN(new_n1249_));
  OAI21_X1   g0864(.A1(new_n1245_), .A2(new_n1246_), .B(new_n1249_), .ZN(\f[84] ));
  NAND3_X1   g0865(.A1(new_n1203_), .A2(new_n1226_), .A3(new_n1235_), .ZN(new_n1251_));
  NOR2_X1    g0866(.A1(new_n1248_), .A2(\b[83] ), .ZN(new_n1252_));
  AOI21_X1   g0867(.A1(new_n1248_), .A2(\b[83] ), .B(\a[83] ), .ZN(new_n1253_));
  NOR2_X1    g0868(.A1(new_n1253_), .A2(new_n1252_), .ZN(new_n1254_));
  INV_X1     g0869(.I(new_n1254_), .ZN(new_n1255_));
  AOI21_X1   g0870(.A1(new_n1251_), .A2(new_n1232_), .B(new_n1255_), .ZN(new_n1256_));
  INV_X1     g0871(.I(\a[85] ), .ZN(new_n1257_));
  INV_X1     g0872(.I(\b[85] ), .ZN(new_n1258_));
  NOR2_X1    g0873(.A1(new_n1257_), .A2(new_n1258_), .ZN(new_n1259_));
  XOR2_X1    g0874(.A1(new_n1256_), .A2(new_n1259_), .Z(new_n1260_));
  XOR2_X1    g0875(.A1(new_n1260_), .A2(new_n1247_), .Z(\f[85] ));
  INV_X1     g0876(.I(new_n1247_), .ZN(new_n1262_));
  AOI21_X1   g0877(.A1(new_n1257_), .A2(new_n1258_), .B(new_n1262_), .ZN(new_n1263_));
  AOI21_X1   g0878(.A1(new_n1256_), .A2(new_n1263_), .B(new_n1259_), .ZN(new_n1264_));
  XNOR2_X1   g0879(.A1(\a[86] ), .A2(\b[86] ), .ZN(new_n1265_));
  NAND2_X1   g0880(.A1(\a[86] ), .A2(\b[86] ), .ZN(new_n1266_));
  NOR2_X1    g0881(.A1(\a[86] ), .A2(\b[86] ), .ZN(new_n1267_));
  INV_X1     g0882(.I(new_n1267_), .ZN(new_n1268_));
  NAND2_X1   g0883(.A1(new_n1268_), .A2(new_n1266_), .ZN(new_n1269_));
  NAND2_X1   g0884(.A1(new_n1264_), .A2(new_n1269_), .ZN(new_n1270_));
  OAI21_X1   g0885(.A1(new_n1264_), .A2(new_n1265_), .B(new_n1270_), .ZN(\f[86] ));
  INV_X1     g0886(.I(new_n1264_), .ZN(new_n1272_));
  AOI21_X1   g0887(.A1(new_n1272_), .A2(new_n1266_), .B(new_n1267_), .ZN(new_n1273_));
  XNOR2_X1   g0888(.A1(\a[87] ), .A2(\b[87] ), .ZN(new_n1274_));
  AND2_X2    g0889(.A1(\a[87] ), .A2(\b[87] ), .Z(new_n1275_));
  NOR2_X1    g0890(.A1(\a[87] ), .A2(\b[87] ), .ZN(new_n1276_));
  OAI21_X1   g0891(.A1(new_n1275_), .A2(new_n1276_), .B(new_n1273_), .ZN(new_n1277_));
  OAI21_X1   g0892(.A1(new_n1273_), .A2(new_n1274_), .B(new_n1277_), .ZN(\f[87] ));
  INV_X1     g0893(.I(new_n1275_), .ZN(new_n1279_));
  INV_X1     g0894(.I(new_n1263_), .ZN(new_n1280_));
  NOR3_X1    g0895(.A1(new_n1236_), .A2(new_n1255_), .A3(new_n1280_), .ZN(new_n1281_));
  INV_X1     g0896(.I(\b[86] ), .ZN(new_n1282_));
  INV_X1     g0897(.I(new_n1276_), .ZN(new_n1283_));
  AOI21_X1   g0898(.A1(new_n1276_), .A2(\b[86] ), .B(\a[86] ), .ZN(new_n1284_));
  AOI21_X1   g0899(.A1(new_n1282_), .A2(new_n1283_), .B(new_n1284_), .ZN(new_n1285_));
  OAI21_X1   g0900(.A1(new_n1281_), .A2(new_n1259_), .B(new_n1285_), .ZN(new_n1286_));
  INV_X1     g0901(.I(\a[88] ), .ZN(new_n1287_));
  INV_X1     g0902(.I(\b[88] ), .ZN(new_n1288_));
  NOR2_X1    g0903(.A1(new_n1287_), .A2(new_n1288_), .ZN(new_n1289_));
  XOR2_X1    g0904(.A1(new_n1286_), .A2(new_n1289_), .Z(new_n1290_));
  XOR2_X1    g0905(.A1(new_n1290_), .A2(new_n1279_), .Z(\f[88] ));
  INV_X1     g0906(.I(new_n1289_), .ZN(new_n1292_));
  AOI21_X1   g0907(.A1(new_n1287_), .A2(new_n1288_), .B(new_n1279_), .ZN(new_n1293_));
  INV_X1     g0908(.I(new_n1293_), .ZN(new_n1294_));
  OAI21_X1   g0909(.A1(new_n1286_), .A2(new_n1294_), .B(new_n1292_), .ZN(new_n1295_));
  INV_X1     g0910(.I(new_n1295_), .ZN(new_n1296_));
  XNOR2_X1   g0911(.A1(\a[89] ), .A2(\b[89] ), .ZN(new_n1297_));
  INV_X1     g0912(.I(\a[89] ), .ZN(new_n1298_));
  INV_X1     g0913(.I(\b[89] ), .ZN(new_n1299_));
  NOR2_X1    g0914(.A1(new_n1298_), .A2(new_n1299_), .ZN(new_n1300_));
  NOR2_X1    g0915(.A1(\a[89] ), .A2(\b[89] ), .ZN(new_n1301_));
  OAI21_X1   g0916(.A1(new_n1300_), .A2(new_n1301_), .B(new_n1296_), .ZN(new_n1302_));
  OAI21_X1   g0917(.A1(new_n1296_), .A2(new_n1297_), .B(new_n1302_), .ZN(\f[89] ));
  NAND2_X1   g0918(.A1(new_n1298_), .A2(new_n1299_), .ZN(new_n1304_));
  OAI21_X1   g0919(.A1(new_n1296_), .A2(new_n1300_), .B(new_n1304_), .ZN(new_n1305_));
  XOR2_X1    g0920(.A1(\a[90] ), .A2(\b[90] ), .Z(new_n1306_));
  NAND2_X1   g0921(.A1(new_n1305_), .A2(new_n1306_), .ZN(new_n1307_));
  INV_X1     g0922(.I(\a[90] ), .ZN(new_n1308_));
  INV_X1     g0923(.I(\b[90] ), .ZN(new_n1309_));
  NOR2_X1    g0924(.A1(new_n1308_), .A2(new_n1309_), .ZN(new_n1310_));
  NOR2_X1    g0925(.A1(\a[90] ), .A2(\b[90] ), .ZN(new_n1311_));
  NOR2_X1    g0926(.A1(new_n1310_), .A2(new_n1311_), .ZN(new_n1312_));
  OAI21_X1   g0927(.A1(new_n1305_), .A2(new_n1312_), .B(new_n1307_), .ZN(\f[90] ));
  INV_X1     g0928(.I(new_n1310_), .ZN(new_n1314_));
  INV_X1     g0929(.I(new_n1285_), .ZN(new_n1315_));
  NOR3_X1    g0930(.A1(new_n1264_), .A2(new_n1315_), .A3(new_n1294_), .ZN(new_n1316_));
  NOR2_X1    g0931(.A1(new_n1311_), .A2(\b[89] ), .ZN(new_n1317_));
  AOI21_X1   g0932(.A1(new_n1311_), .A2(\b[89] ), .B(\a[89] ), .ZN(new_n1318_));
  NOR2_X1    g0933(.A1(new_n1318_), .A2(new_n1317_), .ZN(new_n1319_));
  OAI21_X1   g0934(.A1(new_n1316_), .A2(new_n1289_), .B(new_n1319_), .ZN(new_n1320_));
  INV_X1     g0935(.I(\a[91] ), .ZN(new_n1321_));
  INV_X1     g0936(.I(\b[91] ), .ZN(new_n1322_));
  NOR2_X1    g0937(.A1(new_n1321_), .A2(new_n1322_), .ZN(new_n1323_));
  XOR2_X1    g0938(.A1(new_n1320_), .A2(new_n1323_), .Z(new_n1324_));
  XOR2_X1    g0939(.A1(new_n1324_), .A2(new_n1314_), .Z(\f[91] ));
  INV_X1     g0940(.I(new_n1323_), .ZN(new_n1326_));
  AOI21_X1   g0941(.A1(new_n1321_), .A2(new_n1322_), .B(new_n1314_), .ZN(new_n1327_));
  INV_X1     g0942(.I(new_n1327_), .ZN(new_n1328_));
  OAI21_X1   g0943(.A1(new_n1320_), .A2(new_n1328_), .B(new_n1326_), .ZN(new_n1329_));
  INV_X1     g0944(.I(new_n1329_), .ZN(new_n1330_));
  XNOR2_X1   g0945(.A1(\a[92] ), .A2(\b[92] ), .ZN(new_n1331_));
  INV_X1     g0946(.I(\a[92] ), .ZN(new_n1332_));
  INV_X1     g0947(.I(\b[92] ), .ZN(new_n1333_));
  NOR2_X1    g0948(.A1(new_n1332_), .A2(new_n1333_), .ZN(new_n1334_));
  NOR2_X1    g0949(.A1(\a[92] ), .A2(\b[92] ), .ZN(new_n1335_));
  OAI21_X1   g0950(.A1(new_n1334_), .A2(new_n1335_), .B(new_n1330_), .ZN(new_n1336_));
  OAI21_X1   g0951(.A1(new_n1330_), .A2(new_n1331_), .B(new_n1336_), .ZN(\f[92] ));
  NAND2_X1   g0952(.A1(new_n1332_), .A2(new_n1333_), .ZN(new_n1338_));
  OAI21_X1   g0953(.A1(new_n1330_), .A2(new_n1334_), .B(new_n1338_), .ZN(new_n1339_));
  XOR2_X1    g0954(.A1(\a[93] ), .A2(\b[93] ), .Z(new_n1340_));
  NAND2_X1   g0955(.A1(new_n1339_), .A2(new_n1340_), .ZN(new_n1341_));
  INV_X1     g0956(.I(\a[93] ), .ZN(new_n1342_));
  INV_X1     g0957(.I(\b[93] ), .ZN(new_n1343_));
  NOR2_X1    g0958(.A1(new_n1342_), .A2(new_n1343_), .ZN(new_n1344_));
  NOR2_X1    g0959(.A1(\a[93] ), .A2(\b[93] ), .ZN(new_n1345_));
  NOR2_X1    g0960(.A1(new_n1344_), .A2(new_n1345_), .ZN(new_n1346_));
  OAI21_X1   g0961(.A1(new_n1339_), .A2(new_n1346_), .B(new_n1341_), .ZN(\f[93] ));
  INV_X1     g0962(.I(new_n1344_), .ZN(new_n1348_));
  NAND3_X1   g0963(.A1(new_n1295_), .A2(new_n1319_), .A3(new_n1327_), .ZN(new_n1349_));
  INV_X1     g0964(.I(new_n1345_), .ZN(new_n1350_));
  AOI21_X1   g0965(.A1(new_n1345_), .A2(\b[92] ), .B(\a[92] ), .ZN(new_n1351_));
  AOI21_X1   g0966(.A1(new_n1333_), .A2(new_n1350_), .B(new_n1351_), .ZN(new_n1352_));
  INV_X1     g0967(.I(new_n1352_), .ZN(new_n1353_));
  AOI21_X1   g0968(.A1(new_n1349_), .A2(new_n1326_), .B(new_n1353_), .ZN(new_n1354_));
  INV_X1     g0969(.I(\a[94] ), .ZN(new_n1355_));
  INV_X1     g0970(.I(\b[94] ), .ZN(new_n1356_));
  NOR2_X1    g0971(.A1(new_n1355_), .A2(new_n1356_), .ZN(new_n1357_));
  INV_X1     g0972(.I(new_n1357_), .ZN(new_n1358_));
  XOR2_X1    g0973(.A1(new_n1354_), .A2(new_n1358_), .Z(new_n1359_));
  XOR2_X1    g0974(.A1(new_n1359_), .A2(new_n1348_), .Z(\f[94] ));
  AOI21_X1   g0975(.A1(new_n1355_), .A2(new_n1356_), .B(new_n1348_), .ZN(new_n1361_));
  AOI21_X1   g0976(.A1(new_n1354_), .A2(new_n1361_), .B(new_n1357_), .ZN(new_n1362_));
  XNOR2_X1   g0977(.A1(\a[95] ), .A2(\b[95] ), .ZN(new_n1363_));
  NAND2_X1   g0978(.A1(\a[95] ), .A2(\b[95] ), .ZN(new_n1364_));
  NOR2_X1    g0979(.A1(\a[95] ), .A2(\b[95] ), .ZN(new_n1365_));
  INV_X1     g0980(.I(new_n1365_), .ZN(new_n1366_));
  NAND2_X1   g0981(.A1(new_n1366_), .A2(new_n1364_), .ZN(new_n1367_));
  NAND2_X1   g0982(.A1(new_n1362_), .A2(new_n1367_), .ZN(new_n1368_));
  OAI21_X1   g0983(.A1(new_n1362_), .A2(new_n1363_), .B(new_n1368_), .ZN(\f[95] ));
  INV_X1     g0984(.I(new_n1362_), .ZN(new_n1370_));
  AOI21_X1   g0985(.A1(new_n1370_), .A2(new_n1364_), .B(new_n1365_), .ZN(new_n1371_));
  XNOR2_X1   g0986(.A1(\a[96] ), .A2(\b[96] ), .ZN(new_n1372_));
  AND2_X2    g0987(.A1(\a[96] ), .A2(\b[96] ), .Z(new_n1373_));
  NOR2_X1    g0988(.A1(\a[96] ), .A2(\b[96] ), .ZN(new_n1374_));
  OAI21_X1   g0989(.A1(new_n1373_), .A2(new_n1374_), .B(new_n1371_), .ZN(new_n1375_));
  OAI21_X1   g0990(.A1(new_n1371_), .A2(new_n1372_), .B(new_n1375_), .ZN(\f[96] ));
  NAND3_X1   g0991(.A1(new_n1329_), .A2(new_n1352_), .A3(new_n1361_), .ZN(new_n1377_));
  NOR2_X1    g0992(.A1(new_n1374_), .A2(\b[95] ), .ZN(new_n1378_));
  AOI21_X1   g0993(.A1(new_n1374_), .A2(\b[95] ), .B(\a[95] ), .ZN(new_n1379_));
  NOR2_X1    g0994(.A1(new_n1379_), .A2(new_n1378_), .ZN(new_n1380_));
  INV_X1     g0995(.I(new_n1380_), .ZN(new_n1381_));
  AOI21_X1   g0996(.A1(new_n1377_), .A2(new_n1358_), .B(new_n1381_), .ZN(new_n1382_));
  INV_X1     g0997(.I(\a[97] ), .ZN(new_n1383_));
  INV_X1     g0998(.I(\b[97] ), .ZN(new_n1384_));
  NOR2_X1    g0999(.A1(new_n1383_), .A2(new_n1384_), .ZN(new_n1385_));
  XOR2_X1    g1000(.A1(new_n1382_), .A2(new_n1385_), .Z(new_n1386_));
  XOR2_X1    g1001(.A1(new_n1386_), .A2(new_n1373_), .Z(\f[97] ));
  INV_X1     g1002(.I(new_n1373_), .ZN(new_n1388_));
  AOI21_X1   g1003(.A1(new_n1383_), .A2(new_n1384_), .B(new_n1388_), .ZN(new_n1389_));
  AOI21_X1   g1004(.A1(new_n1382_), .A2(new_n1389_), .B(new_n1385_), .ZN(new_n1390_));
  XNOR2_X1   g1005(.A1(\a[98] ), .A2(\b[98] ), .ZN(new_n1391_));
  NAND2_X1   g1006(.A1(\a[98] ), .A2(\b[98] ), .ZN(new_n1392_));
  NOR2_X1    g1007(.A1(\a[98] ), .A2(\b[98] ), .ZN(new_n1393_));
  INV_X1     g1008(.I(new_n1393_), .ZN(new_n1394_));
  NAND2_X1   g1009(.A1(new_n1394_), .A2(new_n1392_), .ZN(new_n1395_));
  NAND2_X1   g1010(.A1(new_n1390_), .A2(new_n1395_), .ZN(new_n1396_));
  OAI21_X1   g1011(.A1(new_n1390_), .A2(new_n1391_), .B(new_n1396_), .ZN(\f[98] ));
  INV_X1     g1012(.I(new_n1390_), .ZN(new_n1398_));
  AOI21_X1   g1013(.A1(new_n1398_), .A2(new_n1392_), .B(new_n1393_), .ZN(new_n1399_));
  XNOR2_X1   g1014(.A1(\a[99] ), .A2(\b[99] ), .ZN(new_n1400_));
  AND2_X2    g1015(.A1(\a[99] ), .A2(\b[99] ), .Z(new_n1401_));
  NOR2_X1    g1016(.A1(\a[99] ), .A2(\b[99] ), .ZN(new_n1402_));
  OAI21_X1   g1017(.A1(new_n1401_), .A2(new_n1402_), .B(new_n1399_), .ZN(new_n1403_));
  OAI21_X1   g1018(.A1(new_n1399_), .A2(new_n1400_), .B(new_n1403_), .ZN(\f[99] ));
  INV_X1     g1019(.I(new_n1401_), .ZN(new_n1405_));
  INV_X1     g1020(.I(new_n1389_), .ZN(new_n1406_));
  NOR3_X1    g1021(.A1(new_n1362_), .A2(new_n1381_), .A3(new_n1406_), .ZN(new_n1407_));
  INV_X1     g1022(.I(\b[98] ), .ZN(new_n1408_));
  INV_X1     g1023(.I(new_n1402_), .ZN(new_n1409_));
  AOI21_X1   g1024(.A1(new_n1402_), .A2(\b[98] ), .B(\a[98] ), .ZN(new_n1410_));
  AOI21_X1   g1025(.A1(new_n1408_), .A2(new_n1409_), .B(new_n1410_), .ZN(new_n1411_));
  OAI21_X1   g1026(.A1(new_n1407_), .A2(new_n1385_), .B(new_n1411_), .ZN(new_n1412_));
  INV_X1     g1027(.I(\a[100] ), .ZN(new_n1413_));
  INV_X1     g1028(.I(\b[100] ), .ZN(new_n1414_));
  NOR2_X1    g1029(.A1(new_n1413_), .A2(new_n1414_), .ZN(new_n1415_));
  XOR2_X1    g1030(.A1(new_n1412_), .A2(new_n1415_), .Z(new_n1416_));
  XOR2_X1    g1031(.A1(new_n1416_), .A2(new_n1405_), .Z(\f[100] ));
  INV_X1     g1032(.I(new_n1415_), .ZN(new_n1418_));
  AOI21_X1   g1033(.A1(new_n1413_), .A2(new_n1414_), .B(new_n1405_), .ZN(new_n1419_));
  INV_X1     g1034(.I(new_n1419_), .ZN(new_n1420_));
  OAI21_X1   g1035(.A1(new_n1412_), .A2(new_n1420_), .B(new_n1418_), .ZN(new_n1421_));
  INV_X1     g1036(.I(new_n1421_), .ZN(new_n1422_));
  XNOR2_X1   g1037(.A1(\a[101] ), .A2(\b[101] ), .ZN(new_n1423_));
  INV_X1     g1038(.I(\a[101] ), .ZN(new_n1424_));
  INV_X1     g1039(.I(\b[101] ), .ZN(new_n1425_));
  NOR2_X1    g1040(.A1(new_n1424_), .A2(new_n1425_), .ZN(new_n1426_));
  NOR2_X1    g1041(.A1(\a[101] ), .A2(\b[101] ), .ZN(new_n1427_));
  OAI21_X1   g1042(.A1(new_n1426_), .A2(new_n1427_), .B(new_n1422_), .ZN(new_n1428_));
  OAI21_X1   g1043(.A1(new_n1422_), .A2(new_n1423_), .B(new_n1428_), .ZN(\f[101] ));
  NAND2_X1   g1044(.A1(new_n1424_), .A2(new_n1425_), .ZN(new_n1430_));
  OAI21_X1   g1045(.A1(new_n1422_), .A2(new_n1426_), .B(new_n1430_), .ZN(new_n1431_));
  XOR2_X1    g1046(.A1(\a[102] ), .A2(\b[102] ), .Z(new_n1432_));
  NAND2_X1   g1047(.A1(new_n1431_), .A2(new_n1432_), .ZN(new_n1433_));
  INV_X1     g1048(.I(\a[102] ), .ZN(new_n1434_));
  INV_X1     g1049(.I(\b[102] ), .ZN(new_n1435_));
  NOR2_X1    g1050(.A1(new_n1434_), .A2(new_n1435_), .ZN(new_n1436_));
  NOR2_X1    g1051(.A1(\a[102] ), .A2(\b[102] ), .ZN(new_n1437_));
  NOR2_X1    g1052(.A1(new_n1436_), .A2(new_n1437_), .ZN(new_n1438_));
  OAI21_X1   g1053(.A1(new_n1431_), .A2(new_n1438_), .B(new_n1433_), .ZN(\f[102] ));
  INV_X1     g1054(.I(new_n1436_), .ZN(new_n1440_));
  INV_X1     g1055(.I(new_n1411_), .ZN(new_n1441_));
  NOR3_X1    g1056(.A1(new_n1390_), .A2(new_n1441_), .A3(new_n1420_), .ZN(new_n1442_));
  NOR2_X1    g1057(.A1(new_n1437_), .A2(\b[101] ), .ZN(new_n1443_));
  AOI21_X1   g1058(.A1(new_n1437_), .A2(\b[101] ), .B(\a[101] ), .ZN(new_n1444_));
  NOR2_X1    g1059(.A1(new_n1444_), .A2(new_n1443_), .ZN(new_n1445_));
  OAI21_X1   g1060(.A1(new_n1442_), .A2(new_n1415_), .B(new_n1445_), .ZN(new_n1446_));
  INV_X1     g1061(.I(\a[103] ), .ZN(new_n1447_));
  INV_X1     g1062(.I(\b[103] ), .ZN(new_n1448_));
  NOR2_X1    g1063(.A1(new_n1447_), .A2(new_n1448_), .ZN(new_n1449_));
  XOR2_X1    g1064(.A1(new_n1446_), .A2(new_n1449_), .Z(new_n1450_));
  XOR2_X1    g1065(.A1(new_n1450_), .A2(new_n1440_), .Z(\f[103] ));
  INV_X1     g1066(.I(new_n1449_), .ZN(new_n1452_));
  AOI21_X1   g1067(.A1(new_n1447_), .A2(new_n1448_), .B(new_n1440_), .ZN(new_n1453_));
  INV_X1     g1068(.I(new_n1453_), .ZN(new_n1454_));
  OAI21_X1   g1069(.A1(new_n1446_), .A2(new_n1454_), .B(new_n1452_), .ZN(new_n1455_));
  INV_X1     g1070(.I(new_n1455_), .ZN(new_n1456_));
  XNOR2_X1   g1071(.A1(\a[104] ), .A2(\b[104] ), .ZN(new_n1457_));
  INV_X1     g1072(.I(\a[104] ), .ZN(new_n1458_));
  INV_X1     g1073(.I(\b[104] ), .ZN(new_n1459_));
  NOR2_X1    g1074(.A1(new_n1458_), .A2(new_n1459_), .ZN(new_n1460_));
  NOR2_X1    g1075(.A1(\a[104] ), .A2(\b[104] ), .ZN(new_n1461_));
  OAI21_X1   g1076(.A1(new_n1460_), .A2(new_n1461_), .B(new_n1456_), .ZN(new_n1462_));
  OAI21_X1   g1077(.A1(new_n1456_), .A2(new_n1457_), .B(new_n1462_), .ZN(\f[104] ));
  NAND2_X1   g1078(.A1(new_n1458_), .A2(new_n1459_), .ZN(new_n1464_));
  OAI21_X1   g1079(.A1(new_n1456_), .A2(new_n1460_), .B(new_n1464_), .ZN(new_n1465_));
  XOR2_X1    g1080(.A1(\a[105] ), .A2(\b[105] ), .Z(new_n1466_));
  NAND2_X1   g1081(.A1(new_n1465_), .A2(new_n1466_), .ZN(new_n1467_));
  INV_X1     g1082(.I(\a[105] ), .ZN(new_n1468_));
  INV_X1     g1083(.I(\b[105] ), .ZN(new_n1469_));
  NOR2_X1    g1084(.A1(new_n1468_), .A2(new_n1469_), .ZN(new_n1470_));
  NOR2_X1    g1085(.A1(\a[105] ), .A2(\b[105] ), .ZN(new_n1471_));
  NOR2_X1    g1086(.A1(new_n1470_), .A2(new_n1471_), .ZN(new_n1472_));
  OAI21_X1   g1087(.A1(new_n1465_), .A2(new_n1472_), .B(new_n1467_), .ZN(\f[105] ));
  INV_X1     g1088(.I(new_n1470_), .ZN(new_n1474_));
  NAND3_X1   g1089(.A1(new_n1421_), .A2(new_n1445_), .A3(new_n1453_), .ZN(new_n1475_));
  INV_X1     g1090(.I(new_n1471_), .ZN(new_n1476_));
  AOI21_X1   g1091(.A1(new_n1471_), .A2(\b[104] ), .B(\a[104] ), .ZN(new_n1477_));
  AOI21_X1   g1092(.A1(new_n1459_), .A2(new_n1476_), .B(new_n1477_), .ZN(new_n1478_));
  INV_X1     g1093(.I(new_n1478_), .ZN(new_n1479_));
  AOI21_X1   g1094(.A1(new_n1475_), .A2(new_n1452_), .B(new_n1479_), .ZN(new_n1480_));
  INV_X1     g1095(.I(\a[106] ), .ZN(new_n1481_));
  INV_X1     g1096(.I(\b[106] ), .ZN(new_n1482_));
  NOR2_X1    g1097(.A1(new_n1481_), .A2(new_n1482_), .ZN(new_n1483_));
  INV_X1     g1098(.I(new_n1483_), .ZN(new_n1484_));
  XOR2_X1    g1099(.A1(new_n1480_), .A2(new_n1484_), .Z(new_n1485_));
  XOR2_X1    g1100(.A1(new_n1485_), .A2(new_n1474_), .Z(\f[106] ));
  AOI21_X1   g1101(.A1(new_n1481_), .A2(new_n1482_), .B(new_n1474_), .ZN(new_n1487_));
  AOI21_X1   g1102(.A1(new_n1480_), .A2(new_n1487_), .B(new_n1483_), .ZN(new_n1488_));
  XNOR2_X1   g1103(.A1(\a[107] ), .A2(\b[107] ), .ZN(new_n1489_));
  NAND2_X1   g1104(.A1(\a[107] ), .A2(\b[107] ), .ZN(new_n1490_));
  NOR2_X1    g1105(.A1(\a[107] ), .A2(\b[107] ), .ZN(new_n1491_));
  INV_X1     g1106(.I(new_n1491_), .ZN(new_n1492_));
  NAND2_X1   g1107(.A1(new_n1492_), .A2(new_n1490_), .ZN(new_n1493_));
  NAND2_X1   g1108(.A1(new_n1488_), .A2(new_n1493_), .ZN(new_n1494_));
  OAI21_X1   g1109(.A1(new_n1488_), .A2(new_n1489_), .B(new_n1494_), .ZN(\f[107] ));
  INV_X1     g1110(.I(new_n1488_), .ZN(new_n1496_));
  AOI21_X1   g1111(.A1(new_n1496_), .A2(new_n1490_), .B(new_n1491_), .ZN(new_n1497_));
  XNOR2_X1   g1112(.A1(\a[108] ), .A2(\b[108] ), .ZN(new_n1498_));
  AND2_X2    g1113(.A1(\a[108] ), .A2(\b[108] ), .Z(new_n1499_));
  NOR2_X1    g1114(.A1(\a[108] ), .A2(\b[108] ), .ZN(new_n1500_));
  OAI21_X1   g1115(.A1(new_n1499_), .A2(new_n1500_), .B(new_n1497_), .ZN(new_n1501_));
  OAI21_X1   g1116(.A1(new_n1497_), .A2(new_n1498_), .B(new_n1501_), .ZN(\f[108] ));
  NAND3_X1   g1117(.A1(new_n1455_), .A2(new_n1478_), .A3(new_n1487_), .ZN(new_n1503_));
  NOR2_X1    g1118(.A1(new_n1500_), .A2(\b[107] ), .ZN(new_n1504_));
  AOI21_X1   g1119(.A1(new_n1500_), .A2(\b[107] ), .B(\a[107] ), .ZN(new_n1505_));
  NOR2_X1    g1120(.A1(new_n1505_), .A2(new_n1504_), .ZN(new_n1506_));
  INV_X1     g1121(.I(new_n1506_), .ZN(new_n1507_));
  AOI21_X1   g1122(.A1(new_n1503_), .A2(new_n1484_), .B(new_n1507_), .ZN(new_n1508_));
  INV_X1     g1123(.I(\a[109] ), .ZN(new_n1509_));
  INV_X1     g1124(.I(\b[109] ), .ZN(new_n1510_));
  NOR2_X1    g1125(.A1(new_n1509_), .A2(new_n1510_), .ZN(new_n1511_));
  XOR2_X1    g1126(.A1(new_n1508_), .A2(new_n1511_), .Z(new_n1512_));
  XOR2_X1    g1127(.A1(new_n1512_), .A2(new_n1499_), .Z(\f[109] ));
  INV_X1     g1128(.I(new_n1499_), .ZN(new_n1514_));
  AOI21_X1   g1129(.A1(new_n1509_), .A2(new_n1510_), .B(new_n1514_), .ZN(new_n1515_));
  AOI21_X1   g1130(.A1(new_n1508_), .A2(new_n1515_), .B(new_n1511_), .ZN(new_n1516_));
  XNOR2_X1   g1131(.A1(\a[110] ), .A2(\b[110] ), .ZN(new_n1517_));
  NAND2_X1   g1132(.A1(\a[110] ), .A2(\b[110] ), .ZN(new_n1518_));
  NOR2_X1    g1133(.A1(\a[110] ), .A2(\b[110] ), .ZN(new_n1519_));
  INV_X1     g1134(.I(new_n1519_), .ZN(new_n1520_));
  NAND2_X1   g1135(.A1(new_n1520_), .A2(new_n1518_), .ZN(new_n1521_));
  NAND2_X1   g1136(.A1(new_n1516_), .A2(new_n1521_), .ZN(new_n1522_));
  OAI21_X1   g1137(.A1(new_n1516_), .A2(new_n1517_), .B(new_n1522_), .ZN(\f[110] ));
  INV_X1     g1138(.I(new_n1516_), .ZN(new_n1524_));
  AOI21_X1   g1139(.A1(new_n1524_), .A2(new_n1518_), .B(new_n1519_), .ZN(new_n1525_));
  XNOR2_X1   g1140(.A1(\a[111] ), .A2(\b[111] ), .ZN(new_n1526_));
  AND2_X2    g1141(.A1(\a[111] ), .A2(\b[111] ), .Z(new_n1527_));
  NOR2_X1    g1142(.A1(\a[111] ), .A2(\b[111] ), .ZN(new_n1528_));
  OAI21_X1   g1143(.A1(new_n1527_), .A2(new_n1528_), .B(new_n1525_), .ZN(new_n1529_));
  OAI21_X1   g1144(.A1(new_n1525_), .A2(new_n1526_), .B(new_n1529_), .ZN(\f[111] ));
  INV_X1     g1145(.I(new_n1527_), .ZN(new_n1531_));
  INV_X1     g1146(.I(new_n1515_), .ZN(new_n1532_));
  NOR3_X1    g1147(.A1(new_n1488_), .A2(new_n1507_), .A3(new_n1532_), .ZN(new_n1533_));
  INV_X1     g1148(.I(\b[110] ), .ZN(new_n1534_));
  INV_X1     g1149(.I(new_n1528_), .ZN(new_n1535_));
  AOI21_X1   g1150(.A1(new_n1528_), .A2(\b[110] ), .B(\a[110] ), .ZN(new_n1536_));
  AOI21_X1   g1151(.A1(new_n1534_), .A2(new_n1535_), .B(new_n1536_), .ZN(new_n1537_));
  OAI21_X1   g1152(.A1(new_n1533_), .A2(new_n1511_), .B(new_n1537_), .ZN(new_n1538_));
  INV_X1     g1153(.I(\a[112] ), .ZN(new_n1539_));
  INV_X1     g1154(.I(\b[112] ), .ZN(new_n1540_));
  NOR2_X1    g1155(.A1(new_n1539_), .A2(new_n1540_), .ZN(new_n1541_));
  XOR2_X1    g1156(.A1(new_n1538_), .A2(new_n1541_), .Z(new_n1542_));
  XOR2_X1    g1157(.A1(new_n1542_), .A2(new_n1531_), .Z(\f[112] ));
  INV_X1     g1158(.I(new_n1541_), .ZN(new_n1544_));
  AOI21_X1   g1159(.A1(new_n1539_), .A2(new_n1540_), .B(new_n1531_), .ZN(new_n1545_));
  INV_X1     g1160(.I(new_n1545_), .ZN(new_n1546_));
  OAI21_X1   g1161(.A1(new_n1538_), .A2(new_n1546_), .B(new_n1544_), .ZN(new_n1547_));
  INV_X1     g1162(.I(new_n1547_), .ZN(new_n1548_));
  XNOR2_X1   g1163(.A1(\a[113] ), .A2(\b[113] ), .ZN(new_n1549_));
  INV_X1     g1164(.I(\a[113] ), .ZN(new_n1550_));
  INV_X1     g1165(.I(\b[113] ), .ZN(new_n1551_));
  NOR2_X1    g1166(.A1(new_n1550_), .A2(new_n1551_), .ZN(new_n1552_));
  NOR2_X1    g1167(.A1(\a[113] ), .A2(\b[113] ), .ZN(new_n1553_));
  OAI21_X1   g1168(.A1(new_n1552_), .A2(new_n1553_), .B(new_n1548_), .ZN(new_n1554_));
  OAI21_X1   g1169(.A1(new_n1548_), .A2(new_n1549_), .B(new_n1554_), .ZN(\f[113] ));
  NAND2_X1   g1170(.A1(new_n1550_), .A2(new_n1551_), .ZN(new_n1556_));
  OAI21_X1   g1171(.A1(new_n1548_), .A2(new_n1552_), .B(new_n1556_), .ZN(new_n1557_));
  XOR2_X1    g1172(.A1(\a[114] ), .A2(\b[114] ), .Z(new_n1558_));
  NAND2_X1   g1173(.A1(new_n1557_), .A2(new_n1558_), .ZN(new_n1559_));
  INV_X1     g1174(.I(\a[114] ), .ZN(new_n1560_));
  INV_X1     g1175(.I(\b[114] ), .ZN(new_n1561_));
  NOR2_X1    g1176(.A1(new_n1560_), .A2(new_n1561_), .ZN(new_n1562_));
  NOR2_X1    g1177(.A1(\a[114] ), .A2(\b[114] ), .ZN(new_n1563_));
  NOR2_X1    g1178(.A1(new_n1562_), .A2(new_n1563_), .ZN(new_n1564_));
  OAI21_X1   g1179(.A1(new_n1557_), .A2(new_n1564_), .B(new_n1559_), .ZN(\f[114] ));
  INV_X1     g1180(.I(new_n1562_), .ZN(new_n1566_));
  INV_X1     g1181(.I(new_n1537_), .ZN(new_n1567_));
  NOR3_X1    g1182(.A1(new_n1516_), .A2(new_n1567_), .A3(new_n1546_), .ZN(new_n1568_));
  NOR2_X1    g1183(.A1(new_n1563_), .A2(\b[113] ), .ZN(new_n1569_));
  AOI21_X1   g1184(.A1(new_n1563_), .A2(\b[113] ), .B(\a[113] ), .ZN(new_n1570_));
  NOR2_X1    g1185(.A1(new_n1570_), .A2(new_n1569_), .ZN(new_n1571_));
  OAI21_X1   g1186(.A1(new_n1568_), .A2(new_n1541_), .B(new_n1571_), .ZN(new_n1572_));
  INV_X1     g1187(.I(\a[115] ), .ZN(new_n1573_));
  INV_X1     g1188(.I(\b[115] ), .ZN(new_n1574_));
  NOR2_X1    g1189(.A1(new_n1573_), .A2(new_n1574_), .ZN(new_n1575_));
  XOR2_X1    g1190(.A1(new_n1572_), .A2(new_n1575_), .Z(new_n1576_));
  XOR2_X1    g1191(.A1(new_n1576_), .A2(new_n1566_), .Z(\f[115] ));
  INV_X1     g1192(.I(new_n1575_), .ZN(new_n1578_));
  AOI21_X1   g1193(.A1(new_n1573_), .A2(new_n1574_), .B(new_n1566_), .ZN(new_n1579_));
  INV_X1     g1194(.I(new_n1579_), .ZN(new_n1580_));
  OAI21_X1   g1195(.A1(new_n1572_), .A2(new_n1580_), .B(new_n1578_), .ZN(new_n1581_));
  INV_X1     g1196(.I(new_n1581_), .ZN(new_n1582_));
  XNOR2_X1   g1197(.A1(\a[116] ), .A2(\b[116] ), .ZN(new_n1583_));
  INV_X1     g1198(.I(\a[116] ), .ZN(new_n1584_));
  INV_X1     g1199(.I(\b[116] ), .ZN(new_n1585_));
  NOR2_X1    g1200(.A1(new_n1584_), .A2(new_n1585_), .ZN(new_n1586_));
  NOR2_X1    g1201(.A1(\a[116] ), .A2(\b[116] ), .ZN(new_n1587_));
  OAI21_X1   g1202(.A1(new_n1586_), .A2(new_n1587_), .B(new_n1582_), .ZN(new_n1588_));
  OAI21_X1   g1203(.A1(new_n1582_), .A2(new_n1583_), .B(new_n1588_), .ZN(\f[116] ));
  NAND2_X1   g1204(.A1(new_n1584_), .A2(new_n1585_), .ZN(new_n1590_));
  OAI21_X1   g1205(.A1(new_n1582_), .A2(new_n1586_), .B(new_n1590_), .ZN(new_n1591_));
  XOR2_X1    g1206(.A1(\a[117] ), .A2(\b[117] ), .Z(new_n1592_));
  NAND2_X1   g1207(.A1(new_n1591_), .A2(new_n1592_), .ZN(new_n1593_));
  NAND2_X1   g1208(.A1(\a[117] ), .A2(\b[117] ), .ZN(new_n1594_));
  NOR2_X1    g1209(.A1(\a[117] ), .A2(\b[117] ), .ZN(new_n1595_));
  INV_X1     g1210(.I(new_n1595_), .ZN(new_n1596_));
  AND2_X2    g1211(.A1(new_n1596_), .A2(new_n1594_), .Z(new_n1597_));
  OAI21_X1   g1212(.A1(new_n1591_), .A2(new_n1597_), .B(new_n1593_), .ZN(\f[117] ));
  NAND3_X1   g1213(.A1(new_n1547_), .A2(new_n1571_), .A3(new_n1579_), .ZN(new_n1599_));
  AOI21_X1   g1214(.A1(new_n1595_), .A2(\b[116] ), .B(\a[116] ), .ZN(new_n1600_));
  AOI21_X1   g1215(.A1(new_n1585_), .A2(new_n1596_), .B(new_n1600_), .ZN(new_n1601_));
  INV_X1     g1216(.I(new_n1601_), .ZN(new_n1602_));
  AOI21_X1   g1217(.A1(new_n1599_), .A2(new_n1578_), .B(new_n1602_), .ZN(new_n1603_));
  INV_X1     g1218(.I(\a[118] ), .ZN(new_n1604_));
  INV_X1     g1219(.I(\b[118] ), .ZN(new_n1605_));
  NOR2_X1    g1220(.A1(new_n1604_), .A2(new_n1605_), .ZN(new_n1606_));
  INV_X1     g1221(.I(new_n1606_), .ZN(new_n1607_));
  XOR2_X1    g1222(.A1(new_n1603_), .A2(new_n1607_), .Z(new_n1608_));
  XOR2_X1    g1223(.A1(new_n1608_), .A2(new_n1594_), .Z(\f[118] ));
  AOI21_X1   g1224(.A1(new_n1604_), .A2(new_n1605_), .B(new_n1594_), .ZN(new_n1610_));
  AOI21_X1   g1225(.A1(new_n1603_), .A2(new_n1610_), .B(new_n1606_), .ZN(new_n1611_));
  XNOR2_X1   g1226(.A1(\a[119] ), .A2(\b[119] ), .ZN(new_n1612_));
  NAND2_X1   g1227(.A1(\a[119] ), .A2(\b[119] ), .ZN(new_n1613_));
  NOR2_X1    g1228(.A1(\a[119] ), .A2(\b[119] ), .ZN(new_n1614_));
  INV_X1     g1229(.I(new_n1614_), .ZN(new_n1615_));
  NAND2_X1   g1230(.A1(new_n1615_), .A2(new_n1613_), .ZN(new_n1616_));
  NAND2_X1   g1231(.A1(new_n1611_), .A2(new_n1616_), .ZN(new_n1617_));
  OAI21_X1   g1232(.A1(new_n1611_), .A2(new_n1612_), .B(new_n1617_), .ZN(\f[119] ));
  NAND3_X1   g1233(.A1(new_n1581_), .A2(new_n1601_), .A3(new_n1610_), .ZN(new_n1619_));
  NAND2_X1   g1234(.A1(new_n1619_), .A2(new_n1607_), .ZN(new_n1620_));
  AOI21_X1   g1235(.A1(new_n1620_), .A2(new_n1613_), .B(new_n1614_), .ZN(new_n1621_));
  XNOR2_X1   g1236(.A1(\a[120] ), .A2(\b[120] ), .ZN(new_n1622_));
  AND2_X2    g1237(.A1(\a[120] ), .A2(\b[120] ), .Z(new_n1623_));
  NOR2_X1    g1238(.A1(\a[120] ), .A2(\b[120] ), .ZN(new_n1624_));
  OAI21_X1   g1239(.A1(new_n1623_), .A2(new_n1624_), .B(new_n1621_), .ZN(new_n1625_));
  OAI21_X1   g1240(.A1(new_n1621_), .A2(new_n1622_), .B(new_n1625_), .ZN(\f[120] ));
  INV_X1     g1241(.I(new_n1623_), .ZN(new_n1627_));
  INV_X1     g1242(.I(\b[119] ), .ZN(new_n1628_));
  INV_X1     g1243(.I(new_n1624_), .ZN(new_n1629_));
  AOI21_X1   g1244(.A1(new_n1624_), .A2(\b[119] ), .B(\a[119] ), .ZN(new_n1630_));
  AOI21_X1   g1245(.A1(new_n1628_), .A2(new_n1629_), .B(new_n1630_), .ZN(new_n1631_));
  INV_X1     g1246(.I(new_n1631_), .ZN(new_n1632_));
  NOR2_X1    g1247(.A1(new_n1611_), .A2(new_n1632_), .ZN(new_n1633_));
  INV_X1     g1248(.I(\a[121] ), .ZN(new_n1634_));
  INV_X1     g1249(.I(\b[121] ), .ZN(new_n1635_));
  NOR2_X1    g1250(.A1(new_n1634_), .A2(new_n1635_), .ZN(new_n1636_));
  INV_X1     g1251(.I(new_n1636_), .ZN(new_n1637_));
  XOR2_X1    g1252(.A1(new_n1633_), .A2(new_n1637_), .Z(new_n1638_));
  XOR2_X1    g1253(.A1(new_n1638_), .A2(new_n1627_), .Z(\f[121] ));
  AOI21_X1   g1254(.A1(new_n1634_), .A2(new_n1635_), .B(new_n1627_), .ZN(new_n1640_));
  NAND3_X1   g1255(.A1(new_n1620_), .A2(new_n1631_), .A3(new_n1640_), .ZN(new_n1641_));
  NAND2_X1   g1256(.A1(new_n1641_), .A2(new_n1637_), .ZN(new_n1642_));
  XOR2_X1    g1257(.A1(\a[122] ), .A2(\b[122] ), .Z(new_n1643_));
  NAND2_X1   g1258(.A1(new_n1642_), .A2(new_n1643_), .ZN(new_n1644_));
  XOR2_X1    g1259(.A1(\a[122] ), .A2(\b[122] ), .Z(new_n1645_));
  OAI21_X1   g1260(.A1(new_n1642_), .A2(new_n1645_), .B(new_n1644_), .ZN(\f[122] ));
  NAND2_X1   g1261(.A1(\a[122] ), .A2(\b[122] ), .ZN(new_n1647_));
  NOR2_X1    g1262(.A1(\a[122] ), .A2(\b[122] ), .ZN(new_n1648_));
  AOI21_X1   g1263(.A1(new_n1642_), .A2(new_n1647_), .B(new_n1648_), .ZN(new_n1649_));
  XNOR2_X1   g1264(.A1(\a[123] ), .A2(\b[123] ), .ZN(new_n1650_));
  INV_X1     g1265(.I(\a[123] ), .ZN(new_n1651_));
  INV_X1     g1266(.I(\b[123] ), .ZN(new_n1652_));
  NOR2_X1    g1267(.A1(new_n1651_), .A2(new_n1652_), .ZN(new_n1653_));
  NOR2_X1    g1268(.A1(\a[123] ), .A2(\b[123] ), .ZN(new_n1654_));
  OAI21_X1   g1269(.A1(new_n1653_), .A2(new_n1654_), .B(new_n1649_), .ZN(new_n1655_));
  OAI21_X1   g1270(.A1(new_n1649_), .A2(new_n1650_), .B(new_n1655_), .ZN(\f[123] ));
  INV_X1     g1271(.I(new_n1640_), .ZN(new_n1657_));
  NOR3_X1    g1272(.A1(new_n1611_), .A2(new_n1632_), .A3(new_n1657_), .ZN(new_n1658_));
  INV_X1     g1273(.I(\b[122] ), .ZN(new_n1659_));
  INV_X1     g1274(.I(new_n1654_), .ZN(new_n1660_));
  AOI21_X1   g1275(.A1(new_n1654_), .A2(\b[122] ), .B(\a[122] ), .ZN(new_n1661_));
  AOI21_X1   g1276(.A1(new_n1659_), .A2(new_n1660_), .B(new_n1661_), .ZN(new_n1662_));
  OAI21_X1   g1277(.A1(new_n1658_), .A2(new_n1636_), .B(new_n1662_), .ZN(new_n1663_));
  INV_X1     g1278(.I(\a[124] ), .ZN(new_n1664_));
  INV_X1     g1279(.I(\b[124] ), .ZN(new_n1665_));
  NOR2_X1    g1280(.A1(new_n1664_), .A2(new_n1665_), .ZN(new_n1666_));
  NAND2_X1   g1281(.A1(new_n1663_), .A2(new_n1666_), .ZN(new_n1667_));
  INV_X1     g1282(.I(new_n1662_), .ZN(new_n1668_));
  AOI21_X1   g1283(.A1(new_n1641_), .A2(new_n1637_), .B(new_n1668_), .ZN(new_n1669_));
  INV_X1     g1284(.I(new_n1666_), .ZN(new_n1670_));
  NAND2_X1   g1285(.A1(new_n1669_), .A2(new_n1670_), .ZN(new_n1671_));
  NAND2_X1   g1286(.A1(new_n1671_), .A2(new_n1667_), .ZN(new_n1672_));
  XOR2_X1    g1287(.A1(new_n1672_), .A2(new_n1653_), .Z(\f[124] ));
  INV_X1     g1288(.I(new_n1653_), .ZN(new_n1674_));
  AOI21_X1   g1289(.A1(new_n1664_), .A2(new_n1665_), .B(new_n1674_), .ZN(new_n1675_));
  AOI21_X1   g1290(.A1(new_n1669_), .A2(new_n1675_), .B(new_n1666_), .ZN(new_n1676_));
  XNOR2_X1   g1291(.A1(\a[125] ), .A2(\b[125] ), .ZN(new_n1677_));
  NAND2_X1   g1292(.A1(\a[125] ), .A2(\b[125] ), .ZN(new_n1678_));
  NOR2_X1    g1293(.A1(\a[125] ), .A2(\b[125] ), .ZN(new_n1679_));
  INV_X1     g1294(.I(new_n1679_), .ZN(new_n1680_));
  NAND2_X1   g1295(.A1(new_n1680_), .A2(new_n1678_), .ZN(new_n1681_));
  NAND2_X1   g1296(.A1(new_n1676_), .A2(new_n1681_), .ZN(new_n1682_));
  OAI21_X1   g1297(.A1(new_n1676_), .A2(new_n1677_), .B(new_n1682_), .ZN(\f[125] ));
  INV_X1     g1298(.I(new_n1675_), .ZN(new_n1684_));
  OAI21_X1   g1299(.A1(new_n1663_), .A2(new_n1684_), .B(new_n1670_), .ZN(new_n1685_));
  AOI21_X1   g1300(.A1(new_n1685_), .A2(new_n1678_), .B(new_n1679_), .ZN(new_n1686_));
  XNOR2_X1   g1301(.A1(\a[126] ), .A2(\b[126] ), .ZN(new_n1687_));
  INV_X1     g1302(.I(\a[126] ), .ZN(new_n1688_));
  INV_X1     g1303(.I(\b[126] ), .ZN(new_n1689_));
  NOR2_X1    g1304(.A1(new_n1688_), .A2(new_n1689_), .ZN(new_n1690_));
  INV_X1     g1305(.I(new_n1690_), .ZN(new_n1691_));
  NOR2_X1    g1306(.A1(\a[126] ), .A2(\b[126] ), .ZN(new_n1692_));
  INV_X1     g1307(.I(new_n1692_), .ZN(new_n1693_));
  NAND2_X1   g1308(.A1(new_n1691_), .A2(new_n1693_), .ZN(new_n1694_));
  NAND2_X1   g1309(.A1(new_n1686_), .A2(new_n1694_), .ZN(new_n1695_));
  OAI21_X1   g1310(.A1(new_n1686_), .A2(new_n1687_), .B(new_n1695_), .ZN(\f[126] ));
  INV_X1     g1311(.I(\b[125] ), .ZN(new_n1697_));
  AOI21_X1   g1312(.A1(new_n1692_), .A2(\b[125] ), .B(\a[125] ), .ZN(new_n1698_));
  AOI21_X1   g1313(.A1(new_n1697_), .A2(new_n1693_), .B(new_n1698_), .ZN(new_n1699_));
  INV_X1     g1314(.I(\a[127] ), .ZN(new_n1700_));
  INV_X1     g1315(.I(\b[127] ), .ZN(new_n1701_));
  NOR2_X1    g1316(.A1(new_n1700_), .A2(new_n1701_), .ZN(new_n1702_));
  INV_X1     g1317(.I(new_n1702_), .ZN(new_n1703_));
  AOI21_X1   g1318(.A1(new_n1685_), .A2(new_n1699_), .B(new_n1703_), .ZN(new_n1704_));
  INV_X1     g1319(.I(new_n1699_), .ZN(new_n1705_));
  NOR3_X1    g1320(.A1(new_n1676_), .A2(new_n1705_), .A3(new_n1702_), .ZN(new_n1706_));
  OAI21_X1   g1321(.A1(new_n1706_), .A2(new_n1704_), .B(new_n1691_), .ZN(new_n1707_));
  OAI21_X1   g1322(.A1(new_n1676_), .A2(new_n1705_), .B(new_n1702_), .ZN(new_n1708_));
  NAND3_X1   g1323(.A1(new_n1685_), .A2(new_n1699_), .A3(new_n1703_), .ZN(new_n1709_));
  NAND3_X1   g1324(.A1(new_n1708_), .A2(new_n1690_), .A3(new_n1709_), .ZN(new_n1710_));
  NAND2_X1   g1325(.A1(new_n1707_), .A2(new_n1710_), .ZN(\f[127] ));
  NAND2_X1   g1326(.A1(new_n1685_), .A2(new_n1699_), .ZN(new_n1712_));
  OAI21_X1   g1327(.A1(\a[127] ), .A2(\b[127] ), .B(new_n1690_), .ZN(new_n1713_));
  OAI21_X1   g1328(.A1(new_n1712_), .A2(new_n1713_), .B(new_n1703_), .ZN(cOut));
endmodule


